`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: lirc572
// Engineer: lirc572
// 
// Create Date: 
// Design Name: NECPU
// Module Name: InstMem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module instMem (
    input  [31:0]  address,
    output reg [31:0] inst
  );
  always @ (address) begin
    inst = 32'd0;
    case (address)
      0: inst = 32'd268468224;
      1: inst = 32'd201342944;
      2: inst = 32'd203484854;
      3: inst = 32'd471859200;
      4: inst = 32'd136314880;
      5: inst = 32'd268468224;
      6: inst = 32'd201342945;
      7: inst = 32'd203484854;
      8: inst = 32'd471859200;
      9: inst = 32'd136314880;
      10: inst = 32'd268468224;
      11: inst = 32'd201342946;
      12: inst = 32'd203484854;
      13: inst = 32'd471859200;
      14: inst = 32'd136314880;
      15: inst = 32'd268468224;
      16: inst = 32'd201342947;
      17: inst = 32'd203484854;
      18: inst = 32'd471859200;
      19: inst = 32'd136314880;
      20: inst = 32'd268468224;
      21: inst = 32'd201342948;
      22: inst = 32'd203484854;
      23: inst = 32'd471859200;
      24: inst = 32'd136314880;
      25: inst = 32'd268468224;
      26: inst = 32'd201342949;
      27: inst = 32'd203484854;
      28: inst = 32'd471859200;
      29: inst = 32'd136314880;
      30: inst = 32'd268468224;
      31: inst = 32'd201342950;
      32: inst = 32'd203484854;
      33: inst = 32'd471859200;
      34: inst = 32'd136314880;
      35: inst = 32'd268468224;
      36: inst = 32'd201342951;
      37: inst = 32'd203484854;
      38: inst = 32'd471859200;
      39: inst = 32'd136314880;
      40: inst = 32'd268468224;
      41: inst = 32'd201342952;
      42: inst = 32'd203484854;
      43: inst = 32'd471859200;
      44: inst = 32'd136314880;
      45: inst = 32'd268468224;
      46: inst = 32'd201342953;
      47: inst = 32'd203484854;
      48: inst = 32'd471859200;
      49: inst = 32'd136314880;
      50: inst = 32'd268468224;
      51: inst = 32'd201342954;
      52: inst = 32'd203484854;
      53: inst = 32'd471859200;
      54: inst = 32'd136314880;
      55: inst = 32'd268468224;
      56: inst = 32'd201342955;
      57: inst = 32'd203461810;
      58: inst = 32'd471859200;
      59: inst = 32'd136314880;
      60: inst = 32'd268468224;
      61: inst = 32'd201342956;
      62: inst = 32'd203484854;
      63: inst = 32'd471859200;
      64: inst = 32'd136314880;
      65: inst = 32'd268468224;
      66: inst = 32'd201342957;
      67: inst = 32'd203484854;
      68: inst = 32'd471859200;
      69: inst = 32'd136314880;
      70: inst = 32'd268468224;
      71: inst = 32'd201342958;
      72: inst = 32'd203484854;
      73: inst = 32'd471859200;
      74: inst = 32'd136314880;
      75: inst = 32'd268468224;
      76: inst = 32'd201342959;
      77: inst = 32'd203484854;
      78: inst = 32'd471859200;
      79: inst = 32'd136314880;
      80: inst = 32'd268468224;
      81: inst = 32'd201342960;
      82: inst = 32'd203484854;
      83: inst = 32'd471859200;
      84: inst = 32'd136314880;
      85: inst = 32'd268468224;
      86: inst = 32'd201342961;
      87: inst = 32'd203484854;
      88: inst = 32'd471859200;
      89: inst = 32'd136314880;
      90: inst = 32'd268468224;
      91: inst = 32'd201342962;
      92: inst = 32'd203484854;
      93: inst = 32'd471859200;
      94: inst = 32'd136314880;
      95: inst = 32'd268468224;
      96: inst = 32'd201342963;
      97: inst = 32'd203484854;
      98: inst = 32'd471859200;
      99: inst = 32'd136314880;
      100: inst = 32'd268468224;
      101: inst = 32'd201342964;
      102: inst = 32'd203484854;
      103: inst = 32'd471859200;
      104: inst = 32'd136314880;
      105: inst = 32'd268468224;
      106: inst = 32'd201342965;
      107: inst = 32'd203484854;
      108: inst = 32'd471859200;
      109: inst = 32'd136314880;
      110: inst = 32'd268468224;
      111: inst = 32'd201342966;
      112: inst = 32'd203484854;
      113: inst = 32'd471859200;
      114: inst = 32'd136314880;
      115: inst = 32'd268468224;
      116: inst = 32'd201342967;
      117: inst = 32'd203484854;
      118: inst = 32'd471859200;
      119: inst = 32'd136314880;
      120: inst = 32'd268468224;
      121: inst = 32'd201342968;
      122: inst = 32'd203484854;
      123: inst = 32'd471859200;
      124: inst = 32'd136314880;
      125: inst = 32'd268468224;
      126: inst = 32'd201342969;
      127: inst = 32'd203484854;
      128: inst = 32'd471859200;
      129: inst = 32'd136314880;
      130: inst = 32'd268468224;
      131: inst = 32'd201342970;
      132: inst = 32'd203484854;
      133: inst = 32'd471859200;
      134: inst = 32'd136314880;
      135: inst = 32'd268468224;
      136: inst = 32'd201342971;
      137: inst = 32'd203484854;
      138: inst = 32'd471859200;
      139: inst = 32'd136314880;
      140: inst = 32'd268468224;
      141: inst = 32'd201342972;
      142: inst = 32'd203484854;
      143: inst = 32'd471859200;
      144: inst = 32'd136314880;
      145: inst = 32'd268468224;
      146: inst = 32'd201342973;
      147: inst = 32'd203484854;
      148: inst = 32'd471859200;
      149: inst = 32'd136314880;
      150: inst = 32'd268468224;
      151: inst = 32'd201342974;
      152: inst = 32'd203484854;
      153: inst = 32'd471859200;
      154: inst = 32'd136314880;
      155: inst = 32'd268468224;
      156: inst = 32'd201342975;
      157: inst = 32'd203484854;
      158: inst = 32'd471859200;
      159: inst = 32'd136314880;
      160: inst = 32'd268468224;
      161: inst = 32'd201342976;
      162: inst = 32'd203484854;
      163: inst = 32'd471859200;
      164: inst = 32'd136314880;
      165: inst = 32'd268468224;
      166: inst = 32'd201342977;
      167: inst = 32'd203484854;
      168: inst = 32'd471859200;
      169: inst = 32'd136314880;
      170: inst = 32'd268468224;
      171: inst = 32'd201342978;
      172: inst = 32'd203484854;
      173: inst = 32'd471859200;
      174: inst = 32'd136314880;
      175: inst = 32'd268468224;
      176: inst = 32'd201342979;
      177: inst = 32'd203484854;
      178: inst = 32'd471859200;
      179: inst = 32'd136314880;
      180: inst = 32'd268468224;
      181: inst = 32'd201342980;
      182: inst = 32'd203484854;
      183: inst = 32'd471859200;
      184: inst = 32'd136314880;
      185: inst = 32'd268468224;
      186: inst = 32'd201342981;
      187: inst = 32'd203484854;
      188: inst = 32'd471859200;
      189: inst = 32'd136314880;
      190: inst = 32'd268468224;
      191: inst = 32'd201342982;
      192: inst = 32'd203484854;
      193: inst = 32'd471859200;
      194: inst = 32'd136314880;
      195: inst = 32'd268468224;
      196: inst = 32'd201342983;
      197: inst = 32'd203484854;
      198: inst = 32'd471859200;
      199: inst = 32'd136314880;
      200: inst = 32'd268468224;
      201: inst = 32'd201342984;
      202: inst = 32'd203484854;
      203: inst = 32'd471859200;
      204: inst = 32'd136314880;
      205: inst = 32'd268468224;
      206: inst = 32'd201342985;
      207: inst = 32'd203484854;
      208: inst = 32'd471859200;
      209: inst = 32'd136314880;
      210: inst = 32'd268468224;
      211: inst = 32'd201342986;
      212: inst = 32'd203484854;
      213: inst = 32'd471859200;
      214: inst = 32'd136314880;
      215: inst = 32'd268468224;
      216: inst = 32'd201342987;
      217: inst = 32'd203484854;
      218: inst = 32'd471859200;
      219: inst = 32'd136314880;
      220: inst = 32'd268468224;
      221: inst = 32'd201342988;
      222: inst = 32'd203484854;
      223: inst = 32'd471859200;
      224: inst = 32'd136314880;
      225: inst = 32'd268468224;
      226: inst = 32'd201342989;
      227: inst = 32'd203484854;
      228: inst = 32'd471859200;
      229: inst = 32'd136314880;
      230: inst = 32'd268468224;
      231: inst = 32'd201342990;
      232: inst = 32'd203484854;
      233: inst = 32'd471859200;
      234: inst = 32'd136314880;
      235: inst = 32'd268468224;
      236: inst = 32'd201342991;
      237: inst = 32'd203484854;
      238: inst = 32'd471859200;
      239: inst = 32'd136314880;
      240: inst = 32'd268468224;
      241: inst = 32'd201342992;
      242: inst = 32'd203484854;
      243: inst = 32'd471859200;
      244: inst = 32'd136314880;
      245: inst = 32'd268468224;
      246: inst = 32'd201342993;
      247: inst = 32'd203484854;
      248: inst = 32'd471859200;
      249: inst = 32'd136314880;
      250: inst = 32'd268468224;
      251: inst = 32'd201342994;
      252: inst = 32'd203484854;
      253: inst = 32'd471859200;
      254: inst = 32'd136314880;
      255: inst = 32'd268468224;
      256: inst = 32'd201342995;
      257: inst = 32'd203484854;
      258: inst = 32'd471859200;
      259: inst = 32'd136314880;
      260: inst = 32'd268468224;
      261: inst = 32'd201342996;
      262: inst = 32'd203484854;
      263: inst = 32'd471859200;
      264: inst = 32'd136314880;
      265: inst = 32'd268468224;
      266: inst = 32'd201342997;
      267: inst = 32'd203484854;
      268: inst = 32'd471859200;
      269: inst = 32'd136314880;
      270: inst = 32'd268468224;
      271: inst = 32'd201342998;
      272: inst = 32'd203484854;
      273: inst = 32'd471859200;
      274: inst = 32'd136314880;
      275: inst = 32'd268468224;
      276: inst = 32'd201342999;
      277: inst = 32'd203484854;
      278: inst = 32'd471859200;
      279: inst = 32'd136314880;
      280: inst = 32'd268468224;
      281: inst = 32'd201343000;
      282: inst = 32'd203484854;
      283: inst = 32'd471859200;
      284: inst = 32'd136314880;
      285: inst = 32'd268468224;
      286: inst = 32'd201343001;
      287: inst = 32'd203484854;
      288: inst = 32'd471859200;
      289: inst = 32'd136314880;
      290: inst = 32'd268468224;
      291: inst = 32'd201343002;
      292: inst = 32'd203484854;
      293: inst = 32'd471859200;
      294: inst = 32'd136314880;
      295: inst = 32'd268468224;
      296: inst = 32'd201343003;
      297: inst = 32'd203484854;
      298: inst = 32'd471859200;
      299: inst = 32'd136314880;
      300: inst = 32'd268468224;
      301: inst = 32'd201343004;
      302: inst = 32'd203484854;
      303: inst = 32'd471859200;
      304: inst = 32'd136314880;
      305: inst = 32'd268468224;
      306: inst = 32'd201343005;
      307: inst = 32'd203484854;
      308: inst = 32'd471859200;
      309: inst = 32'd136314880;
      310: inst = 32'd268468224;
      311: inst = 32'd201343006;
      312: inst = 32'd203484854;
      313: inst = 32'd471859200;
      314: inst = 32'd136314880;
      315: inst = 32'd268468224;
      316: inst = 32'd201343007;
      317: inst = 32'd203484854;
      318: inst = 32'd471859200;
      319: inst = 32'd136314880;
      320: inst = 32'd268468224;
      321: inst = 32'd201343008;
      322: inst = 32'd203484854;
      323: inst = 32'd471859200;
      324: inst = 32'd136314880;
      325: inst = 32'd268468224;
      326: inst = 32'd201343009;
      327: inst = 32'd203484854;
      328: inst = 32'd471859200;
      329: inst = 32'd136314880;
      330: inst = 32'd268468224;
      331: inst = 32'd201343010;
      332: inst = 32'd203484854;
      333: inst = 32'd471859200;
      334: inst = 32'd136314880;
      335: inst = 32'd268468224;
      336: inst = 32'd201343011;
      337: inst = 32'd203484854;
      338: inst = 32'd471859200;
      339: inst = 32'd136314880;
      340: inst = 32'd268468224;
      341: inst = 32'd201343012;
      342: inst = 32'd203484854;
      343: inst = 32'd471859200;
      344: inst = 32'd136314880;
      345: inst = 32'd268468224;
      346: inst = 32'd201343013;
      347: inst = 32'd203484854;
      348: inst = 32'd471859200;
      349: inst = 32'd136314880;
      350: inst = 32'd268468224;
      351: inst = 32'd201343014;
      352: inst = 32'd203484854;
      353: inst = 32'd471859200;
      354: inst = 32'd136314880;
      355: inst = 32'd268468224;
      356: inst = 32'd201343015;
      357: inst = 32'd203484854;
      358: inst = 32'd471859200;
      359: inst = 32'd136314880;
      360: inst = 32'd268468224;
      361: inst = 32'd201343016;
      362: inst = 32'd203484854;
      363: inst = 32'd471859200;
      364: inst = 32'd136314880;
      365: inst = 32'd268468224;
      366: inst = 32'd201343017;
      367: inst = 32'd203484854;
      368: inst = 32'd471859200;
      369: inst = 32'd136314880;
      370: inst = 32'd268468224;
      371: inst = 32'd201343018;
      372: inst = 32'd203484854;
      373: inst = 32'd471859200;
      374: inst = 32'd136314880;
      375: inst = 32'd268468224;
      376: inst = 32'd201343019;
      377: inst = 32'd203484854;
      378: inst = 32'd471859200;
      379: inst = 32'd136314880;
      380: inst = 32'd268468224;
      381: inst = 32'd201343020;
      382: inst = 32'd203484854;
      383: inst = 32'd471859200;
      384: inst = 32'd136314880;
      385: inst = 32'd268468224;
      386: inst = 32'd201343021;
      387: inst = 32'd203484854;
      388: inst = 32'd471859200;
      389: inst = 32'd136314880;
      390: inst = 32'd268468224;
      391: inst = 32'd201343022;
      392: inst = 32'd203484854;
      393: inst = 32'd471859200;
      394: inst = 32'd136314880;
      395: inst = 32'd268468224;
      396: inst = 32'd201343023;
      397: inst = 32'd203484854;
      398: inst = 32'd471859200;
      399: inst = 32'd136314880;
      400: inst = 32'd268468224;
      401: inst = 32'd201343024;
      402: inst = 32'd203484854;
      403: inst = 32'd471859200;
      404: inst = 32'd136314880;
      405: inst = 32'd268468224;
      406: inst = 32'd201343025;
      407: inst = 32'd203484854;
      408: inst = 32'd471859200;
      409: inst = 32'd136314880;
      410: inst = 32'd268468224;
      411: inst = 32'd201343026;
      412: inst = 32'd203484854;
      413: inst = 32'd471859200;
      414: inst = 32'd136314880;
      415: inst = 32'd268468224;
      416: inst = 32'd201343027;
      417: inst = 32'd203484854;
      418: inst = 32'd471859200;
      419: inst = 32'd136314880;
      420: inst = 32'd268468224;
      421: inst = 32'd201343028;
      422: inst = 32'd203484854;
      423: inst = 32'd471859200;
      424: inst = 32'd136314880;
      425: inst = 32'd268468224;
      426: inst = 32'd201343029;
      427: inst = 32'd203484854;
      428: inst = 32'd471859200;
      429: inst = 32'd136314880;
      430: inst = 32'd268468224;
      431: inst = 32'd201343030;
      432: inst = 32'd203484854;
      433: inst = 32'd471859200;
      434: inst = 32'd136314880;
      435: inst = 32'd268468224;
      436: inst = 32'd201343031;
      437: inst = 32'd203484854;
      438: inst = 32'd471859200;
      439: inst = 32'd136314880;
      440: inst = 32'd268468224;
      441: inst = 32'd201343032;
      442: inst = 32'd203484854;
      443: inst = 32'd471859200;
      444: inst = 32'd136314880;
      445: inst = 32'd268468224;
      446: inst = 32'd201343033;
      447: inst = 32'd203484854;
      448: inst = 32'd471859200;
      449: inst = 32'd136314880;
      450: inst = 32'd268468224;
      451: inst = 32'd201343034;
      452: inst = 32'd203484854;
      453: inst = 32'd471859200;
      454: inst = 32'd136314880;
      455: inst = 32'd268468224;
      456: inst = 32'd201343035;
      457: inst = 32'd203484854;
      458: inst = 32'd471859200;
      459: inst = 32'd136314880;
      460: inst = 32'd268468224;
      461: inst = 32'd201343036;
      462: inst = 32'd203484854;
      463: inst = 32'd471859200;
      464: inst = 32'd136314880;
      465: inst = 32'd268468224;
      466: inst = 32'd201343037;
      467: inst = 32'd203484854;
      468: inst = 32'd471859200;
      469: inst = 32'd136314880;
      470: inst = 32'd268468224;
      471: inst = 32'd201343038;
      472: inst = 32'd203484854;
      473: inst = 32'd471859200;
      474: inst = 32'd136314880;
      475: inst = 32'd268468224;
      476: inst = 32'd201343039;
      477: inst = 32'd203484854;
      478: inst = 32'd471859200;
      479: inst = 32'd136314880;
      480: inst = 32'd268468224;
      481: inst = 32'd201343040;
      482: inst = 32'd203484854;
      483: inst = 32'd471859200;
      484: inst = 32'd136314880;
      485: inst = 32'd268468224;
      486: inst = 32'd201343041;
      487: inst = 32'd203484854;
      488: inst = 32'd471859200;
      489: inst = 32'd136314880;
      490: inst = 32'd268468224;
      491: inst = 32'd201343042;
      492: inst = 32'd203484854;
      493: inst = 32'd471859200;
      494: inst = 32'd136314880;
      495: inst = 32'd268468224;
      496: inst = 32'd201343043;
      497: inst = 32'd203484854;
      498: inst = 32'd471859200;
      499: inst = 32'd136314880;
      500: inst = 32'd268468224;
      501: inst = 32'd201343044;
      502: inst = 32'd203484854;
      503: inst = 32'd471859200;
      504: inst = 32'd136314880;
      505: inst = 32'd268468224;
      506: inst = 32'd201343045;
      507: inst = 32'd203484854;
      508: inst = 32'd471859200;
      509: inst = 32'd136314880;
      510: inst = 32'd268468224;
      511: inst = 32'd201343046;
      512: inst = 32'd203484854;
      513: inst = 32'd471859200;
      514: inst = 32'd136314880;
      515: inst = 32'd268468224;
      516: inst = 32'd201343047;
      517: inst = 32'd203484854;
      518: inst = 32'd471859200;
      519: inst = 32'd136314880;
      520: inst = 32'd268468224;
      521: inst = 32'd201343048;
      522: inst = 32'd203484854;
      523: inst = 32'd471859200;
      524: inst = 32'd136314880;
      525: inst = 32'd268468224;
      526: inst = 32'd201343049;
      527: inst = 32'd203484854;
      528: inst = 32'd471859200;
      529: inst = 32'd136314880;
      530: inst = 32'd268468224;
      531: inst = 32'd201343050;
      532: inst = 32'd203484854;
      533: inst = 32'd471859200;
      534: inst = 32'd136314880;
      535: inst = 32'd268468224;
      536: inst = 32'd201343051;
      537: inst = 32'd203461810;
      538: inst = 32'd471859200;
      539: inst = 32'd136314880;
      540: inst = 32'd268468224;
      541: inst = 32'd201343052;
      542: inst = 32'd203484854;
      543: inst = 32'd471859200;
      544: inst = 32'd136314880;
      545: inst = 32'd268468224;
      546: inst = 32'd201343053;
      547: inst = 32'd203484854;
      548: inst = 32'd471859200;
      549: inst = 32'd136314880;
      550: inst = 32'd268468224;
      551: inst = 32'd201343054;
      552: inst = 32'd203484854;
      553: inst = 32'd471859200;
      554: inst = 32'd136314880;
      555: inst = 32'd268468224;
      556: inst = 32'd201343055;
      557: inst = 32'd203484854;
      558: inst = 32'd471859200;
      559: inst = 32'd136314880;
      560: inst = 32'd268468224;
      561: inst = 32'd201343056;
      562: inst = 32'd203484854;
      563: inst = 32'd471859200;
      564: inst = 32'd136314880;
      565: inst = 32'd268468224;
      566: inst = 32'd201343057;
      567: inst = 32'd203484854;
      568: inst = 32'd471859200;
      569: inst = 32'd136314880;
      570: inst = 32'd268468224;
      571: inst = 32'd201343058;
      572: inst = 32'd203484854;
      573: inst = 32'd471859200;
      574: inst = 32'd136314880;
      575: inst = 32'd268468224;
      576: inst = 32'd201343059;
      577: inst = 32'd203484854;
      578: inst = 32'd471859200;
      579: inst = 32'd136314880;
      580: inst = 32'd268468224;
      581: inst = 32'd201343060;
      582: inst = 32'd203484854;
      583: inst = 32'd471859200;
      584: inst = 32'd136314880;
      585: inst = 32'd268468224;
      586: inst = 32'd201343061;
      587: inst = 32'd203484854;
      588: inst = 32'd471859200;
      589: inst = 32'd136314880;
      590: inst = 32'd268468224;
      591: inst = 32'd201343062;
      592: inst = 32'd203484854;
      593: inst = 32'd471859200;
      594: inst = 32'd136314880;
      595: inst = 32'd268468224;
      596: inst = 32'd201343063;
      597: inst = 32'd203484854;
      598: inst = 32'd471859200;
      599: inst = 32'd136314880;
      600: inst = 32'd268468224;
      601: inst = 32'd201343064;
      602: inst = 32'd203484854;
      603: inst = 32'd471859200;
      604: inst = 32'd136314880;
      605: inst = 32'd268468224;
      606: inst = 32'd201343065;
      607: inst = 32'd203484854;
      608: inst = 32'd471859200;
      609: inst = 32'd136314880;
      610: inst = 32'd268468224;
      611: inst = 32'd201343066;
      612: inst = 32'd203484854;
      613: inst = 32'd471859200;
      614: inst = 32'd136314880;
      615: inst = 32'd268468224;
      616: inst = 32'd201343067;
      617: inst = 32'd203484854;
      618: inst = 32'd471859200;
      619: inst = 32'd136314880;
      620: inst = 32'd268468224;
      621: inst = 32'd201343068;
      622: inst = 32'd203484854;
      623: inst = 32'd471859200;
      624: inst = 32'd136314880;
      625: inst = 32'd268468224;
      626: inst = 32'd201343069;
      627: inst = 32'd203484854;
      628: inst = 32'd471859200;
      629: inst = 32'd136314880;
      630: inst = 32'd268468224;
      631: inst = 32'd201343070;
      632: inst = 32'd203484854;
      633: inst = 32'd471859200;
      634: inst = 32'd136314880;
      635: inst = 32'd268468224;
      636: inst = 32'd201343071;
      637: inst = 32'd203484854;
      638: inst = 32'd471859200;
      639: inst = 32'd136314880;
      640: inst = 32'd268468224;
      641: inst = 32'd201343072;
      642: inst = 32'd203484854;
      643: inst = 32'd471859200;
      644: inst = 32'd136314880;
      645: inst = 32'd268468224;
      646: inst = 32'd201343073;
      647: inst = 32'd203484854;
      648: inst = 32'd471859200;
      649: inst = 32'd136314880;
      650: inst = 32'd268468224;
      651: inst = 32'd201343074;
      652: inst = 32'd203484854;
      653: inst = 32'd471859200;
      654: inst = 32'd136314880;
      655: inst = 32'd268468224;
      656: inst = 32'd201343075;
      657: inst = 32'd203484854;
      658: inst = 32'd471859200;
      659: inst = 32'd136314880;
      660: inst = 32'd268468224;
      661: inst = 32'd201343076;
      662: inst = 32'd203484854;
      663: inst = 32'd471859200;
      664: inst = 32'd136314880;
      665: inst = 32'd268468224;
      666: inst = 32'd201343077;
      667: inst = 32'd203484854;
      668: inst = 32'd471859200;
      669: inst = 32'd136314880;
      670: inst = 32'd268468224;
      671: inst = 32'd201343078;
      672: inst = 32'd203484854;
      673: inst = 32'd471859200;
      674: inst = 32'd136314880;
      675: inst = 32'd268468224;
      676: inst = 32'd201343079;
      677: inst = 32'd203484854;
      678: inst = 32'd471859200;
      679: inst = 32'd136314880;
      680: inst = 32'd268468224;
      681: inst = 32'd201343080;
      682: inst = 32'd203484854;
      683: inst = 32'd471859200;
      684: inst = 32'd136314880;
      685: inst = 32'd268468224;
      686: inst = 32'd201343081;
      687: inst = 32'd203484854;
      688: inst = 32'd471859200;
      689: inst = 32'd136314880;
      690: inst = 32'd268468224;
      691: inst = 32'd201343082;
      692: inst = 32'd203484854;
      693: inst = 32'd471859200;
      694: inst = 32'd136314880;
      695: inst = 32'd268468224;
      696: inst = 32'd201343083;
      697: inst = 32'd203484854;
      698: inst = 32'd471859200;
      699: inst = 32'd136314880;
      700: inst = 32'd268468224;
      701: inst = 32'd201343084;
      702: inst = 32'd203484854;
      703: inst = 32'd471859200;
      704: inst = 32'd136314880;
      705: inst = 32'd268468224;
      706: inst = 32'd201343085;
      707: inst = 32'd203484854;
      708: inst = 32'd471859200;
      709: inst = 32'd136314880;
      710: inst = 32'd268468224;
      711: inst = 32'd201343086;
      712: inst = 32'd203484854;
      713: inst = 32'd471859200;
      714: inst = 32'd136314880;
      715: inst = 32'd268468224;
      716: inst = 32'd201343087;
      717: inst = 32'd203484854;
      718: inst = 32'd471859200;
      719: inst = 32'd136314880;
      720: inst = 32'd268468224;
      721: inst = 32'd201343088;
      722: inst = 32'd203484854;
      723: inst = 32'd471859200;
      724: inst = 32'd136314880;
      725: inst = 32'd268468224;
      726: inst = 32'd201343089;
      727: inst = 32'd203484854;
      728: inst = 32'd471859200;
      729: inst = 32'd136314880;
      730: inst = 32'd268468224;
      731: inst = 32'd201343090;
      732: inst = 32'd203484854;
      733: inst = 32'd471859200;
      734: inst = 32'd136314880;
      735: inst = 32'd268468224;
      736: inst = 32'd201343091;
      737: inst = 32'd203484854;
      738: inst = 32'd471859200;
      739: inst = 32'd136314880;
      740: inst = 32'd268468224;
      741: inst = 32'd201343092;
      742: inst = 32'd203484854;
      743: inst = 32'd471859200;
      744: inst = 32'd136314880;
      745: inst = 32'd268468224;
      746: inst = 32'd201343093;
      747: inst = 32'd203484854;
      748: inst = 32'd471859200;
      749: inst = 32'd136314880;
      750: inst = 32'd268468224;
      751: inst = 32'd201343094;
      752: inst = 32'd203484854;
      753: inst = 32'd471859200;
      754: inst = 32'd136314880;
      755: inst = 32'd268468224;
      756: inst = 32'd201343095;
      757: inst = 32'd203484854;
      758: inst = 32'd471859200;
      759: inst = 32'd136314880;
      760: inst = 32'd268468224;
      761: inst = 32'd201343096;
      762: inst = 32'd203484854;
      763: inst = 32'd471859200;
      764: inst = 32'd136314880;
      765: inst = 32'd268468224;
      766: inst = 32'd201343097;
      767: inst = 32'd203484854;
      768: inst = 32'd471859200;
      769: inst = 32'd136314880;
      770: inst = 32'd268468224;
      771: inst = 32'd201343098;
      772: inst = 32'd203484854;
      773: inst = 32'd471859200;
      774: inst = 32'd136314880;
      775: inst = 32'd268468224;
      776: inst = 32'd201343099;
      777: inst = 32'd203484854;
      778: inst = 32'd471859200;
      779: inst = 32'd136314880;
      780: inst = 32'd268468224;
      781: inst = 32'd201343100;
      782: inst = 32'd203484854;
      783: inst = 32'd471859200;
      784: inst = 32'd136314880;
      785: inst = 32'd268468224;
      786: inst = 32'd201343101;
      787: inst = 32'd203484854;
      788: inst = 32'd471859200;
      789: inst = 32'd136314880;
      790: inst = 32'd268468224;
      791: inst = 32'd201343102;
      792: inst = 32'd203484854;
      793: inst = 32'd471859200;
      794: inst = 32'd136314880;
      795: inst = 32'd268468224;
      796: inst = 32'd201343103;
      797: inst = 32'd203484854;
      798: inst = 32'd471859200;
      799: inst = 32'd136314880;
      800: inst = 32'd268468224;
      801: inst = 32'd201343104;
      802: inst = 32'd203484854;
      803: inst = 32'd471859200;
      804: inst = 32'd136314880;
      805: inst = 32'd268468224;
      806: inst = 32'd201343105;
      807: inst = 32'd203484854;
      808: inst = 32'd471859200;
      809: inst = 32'd136314880;
      810: inst = 32'd268468224;
      811: inst = 32'd201343106;
      812: inst = 32'd203484854;
      813: inst = 32'd471859200;
      814: inst = 32'd136314880;
      815: inst = 32'd268468224;
      816: inst = 32'd201343107;
      817: inst = 32'd203484854;
      818: inst = 32'd471859200;
      819: inst = 32'd136314880;
      820: inst = 32'd268468224;
      821: inst = 32'd201343108;
      822: inst = 32'd203484854;
      823: inst = 32'd471859200;
      824: inst = 32'd136314880;
      825: inst = 32'd268468224;
      826: inst = 32'd201343109;
      827: inst = 32'd203484854;
      828: inst = 32'd471859200;
      829: inst = 32'd136314880;
      830: inst = 32'd268468224;
      831: inst = 32'd201343110;
      832: inst = 32'd203484854;
      833: inst = 32'd471859200;
      834: inst = 32'd136314880;
      835: inst = 32'd268468224;
      836: inst = 32'd201343111;
      837: inst = 32'd203484854;
      838: inst = 32'd471859200;
      839: inst = 32'd136314880;
      840: inst = 32'd268468224;
      841: inst = 32'd201343112;
      842: inst = 32'd203484854;
      843: inst = 32'd471859200;
      844: inst = 32'd136314880;
      845: inst = 32'd268468224;
      846: inst = 32'd201343113;
      847: inst = 32'd203484854;
      848: inst = 32'd471859200;
      849: inst = 32'd136314880;
      850: inst = 32'd268468224;
      851: inst = 32'd201343114;
      852: inst = 32'd203484854;
      853: inst = 32'd471859200;
      854: inst = 32'd136314880;
      855: inst = 32'd268468224;
      856: inst = 32'd201343115;
      857: inst = 32'd203484854;
      858: inst = 32'd471859200;
      859: inst = 32'd136314880;
      860: inst = 32'd268468224;
      861: inst = 32'd201343116;
      862: inst = 32'd203484854;
      863: inst = 32'd471859200;
      864: inst = 32'd136314880;
      865: inst = 32'd268468224;
      866: inst = 32'd201343117;
      867: inst = 32'd203484854;
      868: inst = 32'd471859200;
      869: inst = 32'd136314880;
      870: inst = 32'd268468224;
      871: inst = 32'd201343118;
      872: inst = 32'd203484854;
      873: inst = 32'd471859200;
      874: inst = 32'd136314880;
      875: inst = 32'd268468224;
      876: inst = 32'd201343119;
      877: inst = 32'd203484854;
      878: inst = 32'd471859200;
      879: inst = 32'd136314880;
      880: inst = 32'd268468224;
      881: inst = 32'd201343120;
      882: inst = 32'd203484854;
      883: inst = 32'd471859200;
      884: inst = 32'd136314880;
      885: inst = 32'd268468224;
      886: inst = 32'd201343121;
      887: inst = 32'd203484854;
      888: inst = 32'd471859200;
      889: inst = 32'd136314880;
      890: inst = 32'd268468224;
      891: inst = 32'd201343122;
      892: inst = 32'd203484854;
      893: inst = 32'd471859200;
      894: inst = 32'd136314880;
      895: inst = 32'd268468224;
      896: inst = 32'd201343123;
      897: inst = 32'd203484854;
      898: inst = 32'd471859200;
      899: inst = 32'd136314880;
      900: inst = 32'd268468224;
      901: inst = 32'd201343124;
      902: inst = 32'd203484854;
      903: inst = 32'd471859200;
      904: inst = 32'd136314880;
      905: inst = 32'd268468224;
      906: inst = 32'd201343125;
      907: inst = 32'd203484854;
      908: inst = 32'd471859200;
      909: inst = 32'd136314880;
      910: inst = 32'd268468224;
      911: inst = 32'd201343126;
      912: inst = 32'd203484854;
      913: inst = 32'd471859200;
      914: inst = 32'd136314880;
      915: inst = 32'd268468224;
      916: inst = 32'd201343127;
      917: inst = 32'd203484854;
      918: inst = 32'd471859200;
      919: inst = 32'd136314880;
      920: inst = 32'd268468224;
      921: inst = 32'd201343128;
      922: inst = 32'd203484854;
      923: inst = 32'd471859200;
      924: inst = 32'd136314880;
      925: inst = 32'd268468224;
      926: inst = 32'd201343129;
      927: inst = 32'd203484854;
      928: inst = 32'd471859200;
      929: inst = 32'd136314880;
      930: inst = 32'd268468224;
      931: inst = 32'd201343130;
      932: inst = 32'd203484854;
      933: inst = 32'd471859200;
      934: inst = 32'd136314880;
      935: inst = 32'd268468224;
      936: inst = 32'd201343131;
      937: inst = 32'd203484854;
      938: inst = 32'd471859200;
      939: inst = 32'd136314880;
      940: inst = 32'd268468224;
      941: inst = 32'd201343132;
      942: inst = 32'd203484854;
      943: inst = 32'd471859200;
      944: inst = 32'd136314880;
      945: inst = 32'd268468224;
      946: inst = 32'd201343133;
      947: inst = 32'd203484854;
      948: inst = 32'd471859200;
      949: inst = 32'd136314880;
      950: inst = 32'd268468224;
      951: inst = 32'd201343134;
      952: inst = 32'd203484854;
      953: inst = 32'd471859200;
      954: inst = 32'd136314880;
      955: inst = 32'd268468224;
      956: inst = 32'd201343135;
      957: inst = 32'd203484854;
      958: inst = 32'd471859200;
      959: inst = 32'd136314880;
      960: inst = 32'd268468224;
      961: inst = 32'd201343136;
      962: inst = 32'd203484854;
      963: inst = 32'd471859200;
      964: inst = 32'd136314880;
      965: inst = 32'd268468224;
      966: inst = 32'd201343137;
      967: inst = 32'd203484854;
      968: inst = 32'd471859200;
      969: inst = 32'd136314880;
      970: inst = 32'd268468224;
      971: inst = 32'd201343138;
      972: inst = 32'd203484854;
      973: inst = 32'd471859200;
      974: inst = 32'd136314880;
      975: inst = 32'd268468224;
      976: inst = 32'd201343139;
      977: inst = 32'd203484854;
      978: inst = 32'd471859200;
      979: inst = 32'd136314880;
      980: inst = 32'd268468224;
      981: inst = 32'd201343140;
      982: inst = 32'd203484854;
      983: inst = 32'd471859200;
      984: inst = 32'd136314880;
      985: inst = 32'd268468224;
      986: inst = 32'd201343141;
      987: inst = 32'd203484854;
      988: inst = 32'd471859200;
      989: inst = 32'd136314880;
      990: inst = 32'd268468224;
      991: inst = 32'd201343142;
      992: inst = 32'd203484854;
      993: inst = 32'd471859200;
      994: inst = 32'd136314880;
      995: inst = 32'd268468224;
      996: inst = 32'd201343143;
      997: inst = 32'd203484854;
      998: inst = 32'd471859200;
      999: inst = 32'd136314880;
      1000: inst = 32'd268468224;
      1001: inst = 32'd201343144;
      1002: inst = 32'd203484854;
      1003: inst = 32'd471859200;
      1004: inst = 32'd136314880;
      1005: inst = 32'd268468224;
      1006: inst = 32'd201343145;
      1007: inst = 32'd203484854;
      1008: inst = 32'd471859200;
      1009: inst = 32'd136314880;
      1010: inst = 32'd268468224;
      1011: inst = 32'd201343146;
      1012: inst = 32'd203484854;
      1013: inst = 32'd471859200;
      1014: inst = 32'd136314880;
      1015: inst = 32'd268468224;
      1016: inst = 32'd201343147;
      1017: inst = 32'd203461810;
      1018: inst = 32'd471859200;
      1019: inst = 32'd136314880;
      1020: inst = 32'd268468224;
      1021: inst = 32'd201343148;
      1022: inst = 32'd203484854;
      1023: inst = 32'd471859200;
      1024: inst = 32'd136314880;
      1025: inst = 32'd268468224;
      1026: inst = 32'd201343149;
      1027: inst = 32'd203484854;
      1028: inst = 32'd471859200;
      1029: inst = 32'd136314880;
      1030: inst = 32'd268468224;
      1031: inst = 32'd201343150;
      1032: inst = 32'd203484854;
      1033: inst = 32'd471859200;
      1034: inst = 32'd136314880;
      1035: inst = 32'd268468224;
      1036: inst = 32'd201343151;
      1037: inst = 32'd203484854;
      1038: inst = 32'd471859200;
      1039: inst = 32'd136314880;
      1040: inst = 32'd268468224;
      1041: inst = 32'd201343152;
      1042: inst = 32'd203484854;
      1043: inst = 32'd471859200;
      1044: inst = 32'd136314880;
      1045: inst = 32'd268468224;
      1046: inst = 32'd201343153;
      1047: inst = 32'd203484854;
      1048: inst = 32'd471859200;
      1049: inst = 32'd136314880;
      1050: inst = 32'd268468224;
      1051: inst = 32'd201343154;
      1052: inst = 32'd203484854;
      1053: inst = 32'd471859200;
      1054: inst = 32'd136314880;
      1055: inst = 32'd268468224;
      1056: inst = 32'd201343155;
      1057: inst = 32'd203484854;
      1058: inst = 32'd471859200;
      1059: inst = 32'd136314880;
      1060: inst = 32'd268468224;
      1061: inst = 32'd201343156;
      1062: inst = 32'd203484854;
      1063: inst = 32'd471859200;
      1064: inst = 32'd136314880;
      1065: inst = 32'd268468224;
      1066: inst = 32'd201343157;
      1067: inst = 32'd203484854;
      1068: inst = 32'd471859200;
      1069: inst = 32'd136314880;
      1070: inst = 32'd268468224;
      1071: inst = 32'd201343158;
      1072: inst = 32'd203484854;
      1073: inst = 32'd471859200;
      1074: inst = 32'd136314880;
      1075: inst = 32'd268468224;
      1076: inst = 32'd201343159;
      1077: inst = 32'd203484854;
      1078: inst = 32'd471859200;
      1079: inst = 32'd136314880;
      1080: inst = 32'd268468224;
      1081: inst = 32'd201343160;
      1082: inst = 32'd203484854;
      1083: inst = 32'd471859200;
      1084: inst = 32'd136314880;
      1085: inst = 32'd268468224;
      1086: inst = 32'd201343161;
      1087: inst = 32'd203484854;
      1088: inst = 32'd471859200;
      1089: inst = 32'd136314880;
      1090: inst = 32'd268468224;
      1091: inst = 32'd201343162;
      1092: inst = 32'd203484854;
      1093: inst = 32'd471859200;
      1094: inst = 32'd136314880;
      1095: inst = 32'd268468224;
      1096: inst = 32'd201343163;
      1097: inst = 32'd203484854;
      1098: inst = 32'd471859200;
      1099: inst = 32'd136314880;
      1100: inst = 32'd268468224;
      1101: inst = 32'd201343164;
      1102: inst = 32'd203484854;
      1103: inst = 32'd471859200;
      1104: inst = 32'd136314880;
      1105: inst = 32'd268468224;
      1106: inst = 32'd201343165;
      1107: inst = 32'd203484854;
      1108: inst = 32'd471859200;
      1109: inst = 32'd136314880;
      1110: inst = 32'd268468224;
      1111: inst = 32'd201343166;
      1112: inst = 32'd203484854;
      1113: inst = 32'd471859200;
      1114: inst = 32'd136314880;
      1115: inst = 32'd268468224;
      1116: inst = 32'd201343167;
      1117: inst = 32'd203484854;
      1118: inst = 32'd471859200;
      1119: inst = 32'd136314880;
      1120: inst = 32'd268468224;
      1121: inst = 32'd201343168;
      1122: inst = 32'd203484854;
      1123: inst = 32'd471859200;
      1124: inst = 32'd136314880;
      1125: inst = 32'd268468224;
      1126: inst = 32'd201343169;
      1127: inst = 32'd203484854;
      1128: inst = 32'd471859200;
      1129: inst = 32'd136314880;
      1130: inst = 32'd268468224;
      1131: inst = 32'd201343170;
      1132: inst = 32'd203484854;
      1133: inst = 32'd471859200;
      1134: inst = 32'd136314880;
      1135: inst = 32'd268468224;
      1136: inst = 32'd201343171;
      1137: inst = 32'd203484854;
      1138: inst = 32'd471859200;
      1139: inst = 32'd136314880;
      1140: inst = 32'd268468224;
      1141: inst = 32'd201343172;
      1142: inst = 32'd203484854;
      1143: inst = 32'd471859200;
      1144: inst = 32'd136314880;
      1145: inst = 32'd268468224;
      1146: inst = 32'd201343173;
      1147: inst = 32'd203484854;
      1148: inst = 32'd471859200;
      1149: inst = 32'd136314880;
      1150: inst = 32'd268468224;
      1151: inst = 32'd201343174;
      1152: inst = 32'd203484854;
      1153: inst = 32'd471859200;
      1154: inst = 32'd136314880;
      1155: inst = 32'd268468224;
      1156: inst = 32'd201343175;
      1157: inst = 32'd203484854;
      1158: inst = 32'd471859200;
      1159: inst = 32'd136314880;
      1160: inst = 32'd268468224;
      1161: inst = 32'd201343176;
      1162: inst = 32'd203484854;
      1163: inst = 32'd471859200;
      1164: inst = 32'd136314880;
      1165: inst = 32'd268468224;
      1166: inst = 32'd201343177;
      1167: inst = 32'd203484854;
      1168: inst = 32'd471859200;
      1169: inst = 32'd136314880;
      1170: inst = 32'd268468224;
      1171: inst = 32'd201343178;
      1172: inst = 32'd203484854;
      1173: inst = 32'd471859200;
      1174: inst = 32'd136314880;
      1175: inst = 32'd268468224;
      1176: inst = 32'd201343179;
      1177: inst = 32'd203484854;
      1178: inst = 32'd471859200;
      1179: inst = 32'd136314880;
      1180: inst = 32'd268468224;
      1181: inst = 32'd201343180;
      1182: inst = 32'd203484854;
      1183: inst = 32'd471859200;
      1184: inst = 32'd136314880;
      1185: inst = 32'd268468224;
      1186: inst = 32'd201343181;
      1187: inst = 32'd203484854;
      1188: inst = 32'd471859200;
      1189: inst = 32'd136314880;
      1190: inst = 32'd268468224;
      1191: inst = 32'd201343182;
      1192: inst = 32'd203484854;
      1193: inst = 32'd471859200;
      1194: inst = 32'd136314880;
      1195: inst = 32'd268468224;
      1196: inst = 32'd201343183;
      1197: inst = 32'd203484854;
      1198: inst = 32'd471859200;
      1199: inst = 32'd136314880;
      1200: inst = 32'd268468224;
      1201: inst = 32'd201343184;
      1202: inst = 32'd203484854;
      1203: inst = 32'd471859200;
      1204: inst = 32'd136314880;
      1205: inst = 32'd268468224;
      1206: inst = 32'd201343185;
      1207: inst = 32'd203484854;
      1208: inst = 32'd471859200;
      1209: inst = 32'd136314880;
      1210: inst = 32'd268468224;
      1211: inst = 32'd201343186;
      1212: inst = 32'd203484854;
      1213: inst = 32'd471859200;
      1214: inst = 32'd136314880;
      1215: inst = 32'd268468224;
      1216: inst = 32'd201343187;
      1217: inst = 32'd203484854;
      1218: inst = 32'd471859200;
      1219: inst = 32'd136314880;
      1220: inst = 32'd268468224;
      1221: inst = 32'd201343188;
      1222: inst = 32'd203484854;
      1223: inst = 32'd471859200;
      1224: inst = 32'd136314880;
      1225: inst = 32'd268468224;
      1226: inst = 32'd201343189;
      1227: inst = 32'd203484854;
      1228: inst = 32'd471859200;
      1229: inst = 32'd136314880;
      1230: inst = 32'd268468224;
      1231: inst = 32'd201343190;
      1232: inst = 32'd203484854;
      1233: inst = 32'd471859200;
      1234: inst = 32'd136314880;
      1235: inst = 32'd268468224;
      1236: inst = 32'd201343191;
      1237: inst = 32'd203484854;
      1238: inst = 32'd471859200;
      1239: inst = 32'd136314880;
      1240: inst = 32'd268468224;
      1241: inst = 32'd201343192;
      1242: inst = 32'd203484854;
      1243: inst = 32'd471859200;
      1244: inst = 32'd136314880;
      1245: inst = 32'd268468224;
      1246: inst = 32'd201343193;
      1247: inst = 32'd203484854;
      1248: inst = 32'd471859200;
      1249: inst = 32'd136314880;
      1250: inst = 32'd268468224;
      1251: inst = 32'd201343194;
      1252: inst = 32'd203484854;
      1253: inst = 32'd471859200;
      1254: inst = 32'd136314880;
      1255: inst = 32'd268468224;
      1256: inst = 32'd201343195;
      1257: inst = 32'd203484854;
      1258: inst = 32'd471859200;
      1259: inst = 32'd136314880;
      1260: inst = 32'd268468224;
      1261: inst = 32'd201343196;
      1262: inst = 32'd203484854;
      1263: inst = 32'd471859200;
      1264: inst = 32'd136314880;
      1265: inst = 32'd268468224;
      1266: inst = 32'd201343197;
      1267: inst = 32'd203484854;
      1268: inst = 32'd471859200;
      1269: inst = 32'd136314880;
      1270: inst = 32'd268468224;
      1271: inst = 32'd201343198;
      1272: inst = 32'd203484854;
      1273: inst = 32'd471859200;
      1274: inst = 32'd136314880;
      1275: inst = 32'd268468224;
      1276: inst = 32'd201343199;
      1277: inst = 32'd203484854;
      1278: inst = 32'd471859200;
      1279: inst = 32'd136314880;
      1280: inst = 32'd268468224;
      1281: inst = 32'd201343200;
      1282: inst = 32'd203484854;
      1283: inst = 32'd471859200;
      1284: inst = 32'd136314880;
      1285: inst = 32'd268468224;
      1286: inst = 32'd201343201;
      1287: inst = 32'd203484854;
      1288: inst = 32'd471859200;
      1289: inst = 32'd136314880;
      1290: inst = 32'd268468224;
      1291: inst = 32'd201343202;
      1292: inst = 32'd203484854;
      1293: inst = 32'd471859200;
      1294: inst = 32'd136314880;
      1295: inst = 32'd268468224;
      1296: inst = 32'd201343203;
      1297: inst = 32'd203484854;
      1298: inst = 32'd471859200;
      1299: inst = 32'd136314880;
      1300: inst = 32'd268468224;
      1301: inst = 32'd201343204;
      1302: inst = 32'd203484854;
      1303: inst = 32'd471859200;
      1304: inst = 32'd136314880;
      1305: inst = 32'd268468224;
      1306: inst = 32'd201343205;
      1307: inst = 32'd203484854;
      1308: inst = 32'd471859200;
      1309: inst = 32'd136314880;
      1310: inst = 32'd268468224;
      1311: inst = 32'd201343206;
      1312: inst = 32'd203484854;
      1313: inst = 32'd471859200;
      1314: inst = 32'd136314880;
      1315: inst = 32'd268468224;
      1316: inst = 32'd201343207;
      1317: inst = 32'd203484854;
      1318: inst = 32'd471859200;
      1319: inst = 32'd136314880;
      1320: inst = 32'd268468224;
      1321: inst = 32'd201343208;
      1322: inst = 32'd203484854;
      1323: inst = 32'd471859200;
      1324: inst = 32'd136314880;
      1325: inst = 32'd268468224;
      1326: inst = 32'd201343209;
      1327: inst = 32'd203484854;
      1328: inst = 32'd471859200;
      1329: inst = 32'd136314880;
      1330: inst = 32'd268468224;
      1331: inst = 32'd201343210;
      1332: inst = 32'd203484854;
      1333: inst = 32'd471859200;
      1334: inst = 32'd136314880;
      1335: inst = 32'd268468224;
      1336: inst = 32'd201343211;
      1337: inst = 32'd203484854;
      1338: inst = 32'd471859200;
      1339: inst = 32'd136314880;
      1340: inst = 32'd268468224;
      1341: inst = 32'd201343212;
      1342: inst = 32'd203484854;
      1343: inst = 32'd471859200;
      1344: inst = 32'd136314880;
      1345: inst = 32'd268468224;
      1346: inst = 32'd201343213;
      1347: inst = 32'd203484854;
      1348: inst = 32'd471859200;
      1349: inst = 32'd136314880;
      1350: inst = 32'd268468224;
      1351: inst = 32'd201343214;
      1352: inst = 32'd203484854;
      1353: inst = 32'd471859200;
      1354: inst = 32'd136314880;
      1355: inst = 32'd268468224;
      1356: inst = 32'd201343215;
      1357: inst = 32'd203484854;
      1358: inst = 32'd471859200;
      1359: inst = 32'd136314880;
      1360: inst = 32'd268468224;
      1361: inst = 32'd201343216;
      1362: inst = 32'd203484854;
      1363: inst = 32'd471859200;
      1364: inst = 32'd136314880;
      1365: inst = 32'd268468224;
      1366: inst = 32'd201343217;
      1367: inst = 32'd203484854;
      1368: inst = 32'd471859200;
      1369: inst = 32'd136314880;
      1370: inst = 32'd268468224;
      1371: inst = 32'd201343218;
      1372: inst = 32'd203484854;
      1373: inst = 32'd471859200;
      1374: inst = 32'd136314880;
      1375: inst = 32'd268468224;
      1376: inst = 32'd201343219;
      1377: inst = 32'd203484854;
      1378: inst = 32'd471859200;
      1379: inst = 32'd136314880;
      1380: inst = 32'd268468224;
      1381: inst = 32'd201343220;
      1382: inst = 32'd203484854;
      1383: inst = 32'd471859200;
      1384: inst = 32'd136314880;
      1385: inst = 32'd268468224;
      1386: inst = 32'd201343221;
      1387: inst = 32'd203484854;
      1388: inst = 32'd471859200;
      1389: inst = 32'd136314880;
      1390: inst = 32'd268468224;
      1391: inst = 32'd201343222;
      1392: inst = 32'd203484854;
      1393: inst = 32'd471859200;
      1394: inst = 32'd136314880;
      1395: inst = 32'd268468224;
      1396: inst = 32'd201343223;
      1397: inst = 32'd203484854;
      1398: inst = 32'd471859200;
      1399: inst = 32'd136314880;
      1400: inst = 32'd268468224;
      1401: inst = 32'd201343224;
      1402: inst = 32'd203484854;
      1403: inst = 32'd471859200;
      1404: inst = 32'd136314880;
      1405: inst = 32'd268468224;
      1406: inst = 32'd201343225;
      1407: inst = 32'd203484854;
      1408: inst = 32'd471859200;
      1409: inst = 32'd136314880;
      1410: inst = 32'd268468224;
      1411: inst = 32'd201343226;
      1412: inst = 32'd203484854;
      1413: inst = 32'd471859200;
      1414: inst = 32'd136314880;
      1415: inst = 32'd268468224;
      1416: inst = 32'd201343227;
      1417: inst = 32'd203484854;
      1418: inst = 32'd471859200;
      1419: inst = 32'd136314880;
      1420: inst = 32'd268468224;
      1421: inst = 32'd201343228;
      1422: inst = 32'd203484854;
      1423: inst = 32'd471859200;
      1424: inst = 32'd136314880;
      1425: inst = 32'd268468224;
      1426: inst = 32'd201343229;
      1427: inst = 32'd203484854;
      1428: inst = 32'd471859200;
      1429: inst = 32'd136314880;
      1430: inst = 32'd268468224;
      1431: inst = 32'd201343230;
      1432: inst = 32'd203484854;
      1433: inst = 32'd471859200;
      1434: inst = 32'd136314880;
      1435: inst = 32'd268468224;
      1436: inst = 32'd201343231;
      1437: inst = 32'd203484854;
      1438: inst = 32'd471859200;
      1439: inst = 32'd136314880;
      1440: inst = 32'd268468224;
      1441: inst = 32'd201343232;
      1442: inst = 32'd203484854;
      1443: inst = 32'd471859200;
      1444: inst = 32'd136314880;
      1445: inst = 32'd268468224;
      1446: inst = 32'd201343233;
      1447: inst = 32'd203484854;
      1448: inst = 32'd471859200;
      1449: inst = 32'd136314880;
      1450: inst = 32'd268468224;
      1451: inst = 32'd201343234;
      1452: inst = 32'd203484854;
      1453: inst = 32'd471859200;
      1454: inst = 32'd136314880;
      1455: inst = 32'd268468224;
      1456: inst = 32'd201343235;
      1457: inst = 32'd203484854;
      1458: inst = 32'd471859200;
      1459: inst = 32'd136314880;
      1460: inst = 32'd268468224;
      1461: inst = 32'd201343236;
      1462: inst = 32'd203484854;
      1463: inst = 32'd471859200;
      1464: inst = 32'd136314880;
      1465: inst = 32'd268468224;
      1466: inst = 32'd201343237;
      1467: inst = 32'd203484854;
      1468: inst = 32'd471859200;
      1469: inst = 32'd136314880;
      1470: inst = 32'd268468224;
      1471: inst = 32'd201343238;
      1472: inst = 32'd203484854;
      1473: inst = 32'd471859200;
      1474: inst = 32'd136314880;
      1475: inst = 32'd268468224;
      1476: inst = 32'd201343239;
      1477: inst = 32'd203484854;
      1478: inst = 32'd471859200;
      1479: inst = 32'd136314880;
      1480: inst = 32'd268468224;
      1481: inst = 32'd201343240;
      1482: inst = 32'd203484854;
      1483: inst = 32'd471859200;
      1484: inst = 32'd136314880;
      1485: inst = 32'd268468224;
      1486: inst = 32'd201343241;
      1487: inst = 32'd203484854;
      1488: inst = 32'd471859200;
      1489: inst = 32'd136314880;
      1490: inst = 32'd268468224;
      1491: inst = 32'd201343242;
      1492: inst = 32'd203484854;
      1493: inst = 32'd471859200;
      1494: inst = 32'd136314880;
      1495: inst = 32'd268468224;
      1496: inst = 32'd201343243;
      1497: inst = 32'd203461810;
      1498: inst = 32'd471859200;
      1499: inst = 32'd136314880;
      1500: inst = 32'd268468224;
      1501: inst = 32'd201343244;
      1502: inst = 32'd203484854;
      1503: inst = 32'd471859200;
      1504: inst = 32'd136314880;
      1505: inst = 32'd268468224;
      1506: inst = 32'd201343245;
      1507: inst = 32'd203484854;
      1508: inst = 32'd471859200;
      1509: inst = 32'd136314880;
      1510: inst = 32'd268468224;
      1511: inst = 32'd201343246;
      1512: inst = 32'd203484854;
      1513: inst = 32'd471859200;
      1514: inst = 32'd136314880;
      1515: inst = 32'd268468224;
      1516: inst = 32'd201343247;
      1517: inst = 32'd203484854;
      1518: inst = 32'd471859200;
      1519: inst = 32'd136314880;
      1520: inst = 32'd268468224;
      1521: inst = 32'd201343248;
      1522: inst = 32'd203484854;
      1523: inst = 32'd471859200;
      1524: inst = 32'd136314880;
      1525: inst = 32'd268468224;
      1526: inst = 32'd201343249;
      1527: inst = 32'd203484854;
      1528: inst = 32'd471859200;
      1529: inst = 32'd136314880;
      1530: inst = 32'd268468224;
      1531: inst = 32'd201343250;
      1532: inst = 32'd203484854;
      1533: inst = 32'd471859200;
      1534: inst = 32'd136314880;
      1535: inst = 32'd268468224;
      1536: inst = 32'd201343251;
      1537: inst = 32'd203484854;
      1538: inst = 32'd471859200;
      1539: inst = 32'd136314880;
      1540: inst = 32'd268468224;
      1541: inst = 32'd201343252;
      1542: inst = 32'd203484854;
      1543: inst = 32'd471859200;
      1544: inst = 32'd136314880;
      1545: inst = 32'd268468224;
      1546: inst = 32'd201343253;
      1547: inst = 32'd203484854;
      1548: inst = 32'd471859200;
      1549: inst = 32'd136314880;
      1550: inst = 32'd268468224;
      1551: inst = 32'd201343254;
      1552: inst = 32'd203484854;
      1553: inst = 32'd471859200;
      1554: inst = 32'd136314880;
      1555: inst = 32'd268468224;
      1556: inst = 32'd201343255;
      1557: inst = 32'd203484854;
      1558: inst = 32'd471859200;
      1559: inst = 32'd136314880;
      1560: inst = 32'd268468224;
      1561: inst = 32'd201343256;
      1562: inst = 32'd203484854;
      1563: inst = 32'd471859200;
      1564: inst = 32'd136314880;
      1565: inst = 32'd268468224;
      1566: inst = 32'd201343257;
      1567: inst = 32'd203484854;
      1568: inst = 32'd471859200;
      1569: inst = 32'd136314880;
      1570: inst = 32'd268468224;
      1571: inst = 32'd201343258;
      1572: inst = 32'd203484854;
      1573: inst = 32'd471859200;
      1574: inst = 32'd136314880;
      1575: inst = 32'd268468224;
      1576: inst = 32'd201343259;
      1577: inst = 32'd203484854;
      1578: inst = 32'd471859200;
      1579: inst = 32'd136314880;
      1580: inst = 32'd268468224;
      1581: inst = 32'd201343260;
      1582: inst = 32'd203484854;
      1583: inst = 32'd471859200;
      1584: inst = 32'd136314880;
      1585: inst = 32'd268468224;
      1586: inst = 32'd201343261;
      1587: inst = 32'd203484854;
      1588: inst = 32'd471859200;
      1589: inst = 32'd136314880;
      1590: inst = 32'd268468224;
      1591: inst = 32'd201343262;
      1592: inst = 32'd203484854;
      1593: inst = 32'd471859200;
      1594: inst = 32'd136314880;
      1595: inst = 32'd268468224;
      1596: inst = 32'd201343263;
      1597: inst = 32'd203484854;
      1598: inst = 32'd471859200;
      1599: inst = 32'd136314880;
      1600: inst = 32'd268468224;
      1601: inst = 32'd201343264;
      1602: inst = 32'd203484854;
      1603: inst = 32'd471859200;
      1604: inst = 32'd136314880;
      1605: inst = 32'd268468224;
      1606: inst = 32'd201343265;
      1607: inst = 32'd203484854;
      1608: inst = 32'd471859200;
      1609: inst = 32'd136314880;
      1610: inst = 32'd268468224;
      1611: inst = 32'd201343266;
      1612: inst = 32'd203484854;
      1613: inst = 32'd471859200;
      1614: inst = 32'd136314880;
      1615: inst = 32'd268468224;
      1616: inst = 32'd201343267;
      1617: inst = 32'd203484854;
      1618: inst = 32'd471859200;
      1619: inst = 32'd136314880;
      1620: inst = 32'd268468224;
      1621: inst = 32'd201343268;
      1622: inst = 32'd203484854;
      1623: inst = 32'd471859200;
      1624: inst = 32'd136314880;
      1625: inst = 32'd268468224;
      1626: inst = 32'd201343269;
      1627: inst = 32'd203484854;
      1628: inst = 32'd471859200;
      1629: inst = 32'd136314880;
      1630: inst = 32'd268468224;
      1631: inst = 32'd201343270;
      1632: inst = 32'd203484854;
      1633: inst = 32'd471859200;
      1634: inst = 32'd136314880;
      1635: inst = 32'd268468224;
      1636: inst = 32'd201343271;
      1637: inst = 32'd203484854;
      1638: inst = 32'd471859200;
      1639: inst = 32'd136314880;
      1640: inst = 32'd268468224;
      1641: inst = 32'd201343272;
      1642: inst = 32'd203484854;
      1643: inst = 32'd471859200;
      1644: inst = 32'd136314880;
      1645: inst = 32'd268468224;
      1646: inst = 32'd201343273;
      1647: inst = 32'd203484854;
      1648: inst = 32'd471859200;
      1649: inst = 32'd136314880;
      1650: inst = 32'd268468224;
      1651: inst = 32'd201343274;
      1652: inst = 32'd203484854;
      1653: inst = 32'd471859200;
      1654: inst = 32'd136314880;
      1655: inst = 32'd268468224;
      1656: inst = 32'd201343275;
      1657: inst = 32'd203484854;
      1658: inst = 32'd471859200;
      1659: inst = 32'd136314880;
      1660: inst = 32'd268468224;
      1661: inst = 32'd201343276;
      1662: inst = 32'd203484854;
      1663: inst = 32'd471859200;
      1664: inst = 32'd136314880;
      1665: inst = 32'd268468224;
      1666: inst = 32'd201343277;
      1667: inst = 32'd203484854;
      1668: inst = 32'd471859200;
      1669: inst = 32'd136314880;
      1670: inst = 32'd268468224;
      1671: inst = 32'd201343278;
      1672: inst = 32'd203484854;
      1673: inst = 32'd471859200;
      1674: inst = 32'd136314880;
      1675: inst = 32'd268468224;
      1676: inst = 32'd201343279;
      1677: inst = 32'd203484854;
      1678: inst = 32'd471859200;
      1679: inst = 32'd136314880;
      1680: inst = 32'd268468224;
      1681: inst = 32'd201343280;
      1682: inst = 32'd203484854;
      1683: inst = 32'd471859200;
      1684: inst = 32'd136314880;
      1685: inst = 32'd268468224;
      1686: inst = 32'd201343281;
      1687: inst = 32'd203484854;
      1688: inst = 32'd471859200;
      1689: inst = 32'd136314880;
      1690: inst = 32'd268468224;
      1691: inst = 32'd201343282;
      1692: inst = 32'd203484854;
      1693: inst = 32'd471859200;
      1694: inst = 32'd136314880;
      1695: inst = 32'd268468224;
      1696: inst = 32'd201343283;
      1697: inst = 32'd203484854;
      1698: inst = 32'd471859200;
      1699: inst = 32'd136314880;
      1700: inst = 32'd268468224;
      1701: inst = 32'd201343284;
      1702: inst = 32'd203484854;
      1703: inst = 32'd471859200;
      1704: inst = 32'd136314880;
      1705: inst = 32'd268468224;
      1706: inst = 32'd201343285;
      1707: inst = 32'd203484854;
      1708: inst = 32'd471859200;
      1709: inst = 32'd136314880;
      1710: inst = 32'd268468224;
      1711: inst = 32'd201343286;
      1712: inst = 32'd203484854;
      1713: inst = 32'd471859200;
      1714: inst = 32'd136314880;
      1715: inst = 32'd268468224;
      1716: inst = 32'd201343287;
      1717: inst = 32'd203484854;
      1718: inst = 32'd471859200;
      1719: inst = 32'd136314880;
      1720: inst = 32'd268468224;
      1721: inst = 32'd201343288;
      1722: inst = 32'd203484854;
      1723: inst = 32'd471859200;
      1724: inst = 32'd136314880;
      1725: inst = 32'd268468224;
      1726: inst = 32'd201343289;
      1727: inst = 32'd203484854;
      1728: inst = 32'd471859200;
      1729: inst = 32'd136314880;
      1730: inst = 32'd268468224;
      1731: inst = 32'd201343290;
      1732: inst = 32'd203484854;
      1733: inst = 32'd471859200;
      1734: inst = 32'd136314880;
      1735: inst = 32'd268468224;
      1736: inst = 32'd201343291;
      1737: inst = 32'd203484854;
      1738: inst = 32'd471859200;
      1739: inst = 32'd136314880;
      1740: inst = 32'd268468224;
      1741: inst = 32'd201343292;
      1742: inst = 32'd203484854;
      1743: inst = 32'd471859200;
      1744: inst = 32'd136314880;
      1745: inst = 32'd268468224;
      1746: inst = 32'd201343293;
      1747: inst = 32'd203484854;
      1748: inst = 32'd471859200;
      1749: inst = 32'd136314880;
      1750: inst = 32'd268468224;
      1751: inst = 32'd201343294;
      1752: inst = 32'd203484854;
      1753: inst = 32'd471859200;
      1754: inst = 32'd136314880;
      1755: inst = 32'd268468224;
      1756: inst = 32'd201343295;
      1757: inst = 32'd203484854;
      1758: inst = 32'd471859200;
      1759: inst = 32'd136314880;
      1760: inst = 32'd268468224;
      1761: inst = 32'd201343296;
      1762: inst = 32'd203484854;
      1763: inst = 32'd471859200;
      1764: inst = 32'd136314880;
      1765: inst = 32'd268468224;
      1766: inst = 32'd201343297;
      1767: inst = 32'd203484854;
      1768: inst = 32'd471859200;
      1769: inst = 32'd136314880;
      1770: inst = 32'd268468224;
      1771: inst = 32'd201343298;
      1772: inst = 32'd203484854;
      1773: inst = 32'd471859200;
      1774: inst = 32'd136314880;
      1775: inst = 32'd268468224;
      1776: inst = 32'd201343299;
      1777: inst = 32'd203484854;
      1778: inst = 32'd471859200;
      1779: inst = 32'd136314880;
      1780: inst = 32'd268468224;
      1781: inst = 32'd201343300;
      1782: inst = 32'd203484854;
      1783: inst = 32'd471859200;
      1784: inst = 32'd136314880;
      1785: inst = 32'd268468224;
      1786: inst = 32'd201343301;
      1787: inst = 32'd203484854;
      1788: inst = 32'd471859200;
      1789: inst = 32'd136314880;
      1790: inst = 32'd268468224;
      1791: inst = 32'd201343302;
      1792: inst = 32'd203484854;
      1793: inst = 32'd471859200;
      1794: inst = 32'd136314880;
      1795: inst = 32'd268468224;
      1796: inst = 32'd201343303;
      1797: inst = 32'd203484854;
      1798: inst = 32'd471859200;
      1799: inst = 32'd136314880;
      1800: inst = 32'd268468224;
      1801: inst = 32'd201343304;
      1802: inst = 32'd203484854;
      1803: inst = 32'd471859200;
      1804: inst = 32'd136314880;
      1805: inst = 32'd268468224;
      1806: inst = 32'd201343305;
      1807: inst = 32'd203484854;
      1808: inst = 32'd471859200;
      1809: inst = 32'd136314880;
      1810: inst = 32'd268468224;
      1811: inst = 32'd201343306;
      1812: inst = 32'd203484854;
      1813: inst = 32'd471859200;
      1814: inst = 32'd136314880;
      1815: inst = 32'd268468224;
      1816: inst = 32'd201343307;
      1817: inst = 32'd203484854;
      1818: inst = 32'd471859200;
      1819: inst = 32'd136314880;
      1820: inst = 32'd268468224;
      1821: inst = 32'd201343308;
      1822: inst = 32'd203484854;
      1823: inst = 32'd471859200;
      1824: inst = 32'd136314880;
      1825: inst = 32'd268468224;
      1826: inst = 32'd201343309;
      1827: inst = 32'd203484854;
      1828: inst = 32'd471859200;
      1829: inst = 32'd136314880;
      1830: inst = 32'd268468224;
      1831: inst = 32'd201343310;
      1832: inst = 32'd203484854;
      1833: inst = 32'd471859200;
      1834: inst = 32'd136314880;
      1835: inst = 32'd268468224;
      1836: inst = 32'd201343311;
      1837: inst = 32'd203484854;
      1838: inst = 32'd471859200;
      1839: inst = 32'd136314880;
      1840: inst = 32'd268468224;
      1841: inst = 32'd201343312;
      1842: inst = 32'd203484854;
      1843: inst = 32'd471859200;
      1844: inst = 32'd136314880;
      1845: inst = 32'd268468224;
      1846: inst = 32'd201343313;
      1847: inst = 32'd203484854;
      1848: inst = 32'd471859200;
      1849: inst = 32'd136314880;
      1850: inst = 32'd268468224;
      1851: inst = 32'd201343314;
      1852: inst = 32'd203484854;
      1853: inst = 32'd471859200;
      1854: inst = 32'd136314880;
      1855: inst = 32'd268468224;
      1856: inst = 32'd201343315;
      1857: inst = 32'd203484854;
      1858: inst = 32'd471859200;
      1859: inst = 32'd136314880;
      1860: inst = 32'd268468224;
      1861: inst = 32'd201343316;
      1862: inst = 32'd203484854;
      1863: inst = 32'd471859200;
      1864: inst = 32'd136314880;
      1865: inst = 32'd268468224;
      1866: inst = 32'd201343317;
      1867: inst = 32'd203484854;
      1868: inst = 32'd471859200;
      1869: inst = 32'd136314880;
      1870: inst = 32'd268468224;
      1871: inst = 32'd201343318;
      1872: inst = 32'd203484854;
      1873: inst = 32'd471859200;
      1874: inst = 32'd136314880;
      1875: inst = 32'd268468224;
      1876: inst = 32'd201343319;
      1877: inst = 32'd203484854;
      1878: inst = 32'd471859200;
      1879: inst = 32'd136314880;
      1880: inst = 32'd268468224;
      1881: inst = 32'd201343320;
      1882: inst = 32'd203484854;
      1883: inst = 32'd471859200;
      1884: inst = 32'd136314880;
      1885: inst = 32'd268468224;
      1886: inst = 32'd201343321;
      1887: inst = 32'd203484854;
      1888: inst = 32'd471859200;
      1889: inst = 32'd136314880;
      1890: inst = 32'd268468224;
      1891: inst = 32'd201343322;
      1892: inst = 32'd203484854;
      1893: inst = 32'd471859200;
      1894: inst = 32'd136314880;
      1895: inst = 32'd268468224;
      1896: inst = 32'd201343323;
      1897: inst = 32'd203484854;
      1898: inst = 32'd471859200;
      1899: inst = 32'd136314880;
      1900: inst = 32'd268468224;
      1901: inst = 32'd201343324;
      1902: inst = 32'd203484854;
      1903: inst = 32'd471859200;
      1904: inst = 32'd136314880;
      1905: inst = 32'd268468224;
      1906: inst = 32'd201343325;
      1907: inst = 32'd203484854;
      1908: inst = 32'd471859200;
      1909: inst = 32'd136314880;
      1910: inst = 32'd268468224;
      1911: inst = 32'd201343326;
      1912: inst = 32'd203484854;
      1913: inst = 32'd471859200;
      1914: inst = 32'd136314880;
      1915: inst = 32'd268468224;
      1916: inst = 32'd201343327;
      1917: inst = 32'd203484854;
      1918: inst = 32'd471859200;
      1919: inst = 32'd136314880;
      1920: inst = 32'd268468224;
      1921: inst = 32'd201343328;
      1922: inst = 32'd203484854;
      1923: inst = 32'd471859200;
      1924: inst = 32'd136314880;
      1925: inst = 32'd268468224;
      1926: inst = 32'd201343329;
      1927: inst = 32'd203484854;
      1928: inst = 32'd471859200;
      1929: inst = 32'd136314880;
      1930: inst = 32'd268468224;
      1931: inst = 32'd201343330;
      1932: inst = 32'd203484854;
      1933: inst = 32'd471859200;
      1934: inst = 32'd136314880;
      1935: inst = 32'd268468224;
      1936: inst = 32'd201343331;
      1937: inst = 32'd203484854;
      1938: inst = 32'd471859200;
      1939: inst = 32'd136314880;
      1940: inst = 32'd268468224;
      1941: inst = 32'd201343332;
      1942: inst = 32'd203484854;
      1943: inst = 32'd471859200;
      1944: inst = 32'd136314880;
      1945: inst = 32'd268468224;
      1946: inst = 32'd201343333;
      1947: inst = 32'd203484854;
      1948: inst = 32'd471859200;
      1949: inst = 32'd136314880;
      1950: inst = 32'd268468224;
      1951: inst = 32'd201343334;
      1952: inst = 32'd203484854;
      1953: inst = 32'd471859200;
      1954: inst = 32'd136314880;
      1955: inst = 32'd268468224;
      1956: inst = 32'd201343335;
      1957: inst = 32'd203484854;
      1958: inst = 32'd471859200;
      1959: inst = 32'd136314880;
      1960: inst = 32'd268468224;
      1961: inst = 32'd201343336;
      1962: inst = 32'd203484854;
      1963: inst = 32'd471859200;
      1964: inst = 32'd136314880;
      1965: inst = 32'd268468224;
      1966: inst = 32'd201343337;
      1967: inst = 32'd203484854;
      1968: inst = 32'd471859200;
      1969: inst = 32'd136314880;
      1970: inst = 32'd268468224;
      1971: inst = 32'd201343338;
      1972: inst = 32'd203484854;
      1973: inst = 32'd471859200;
      1974: inst = 32'd136314880;
      1975: inst = 32'd268468224;
      1976: inst = 32'd201343339;
      1977: inst = 32'd203461810;
      1978: inst = 32'd471859200;
      1979: inst = 32'd136314880;
      1980: inst = 32'd268468224;
      1981: inst = 32'd201343340;
      1982: inst = 32'd203484854;
      1983: inst = 32'd471859200;
      1984: inst = 32'd136314880;
      1985: inst = 32'd268468224;
      1986: inst = 32'd201343341;
      1987: inst = 32'd203484854;
      1988: inst = 32'd471859200;
      1989: inst = 32'd136314880;
      1990: inst = 32'd268468224;
      1991: inst = 32'd201343342;
      1992: inst = 32'd203484854;
      1993: inst = 32'd471859200;
      1994: inst = 32'd136314880;
      1995: inst = 32'd268468224;
      1996: inst = 32'd201343343;
      1997: inst = 32'd203484854;
      1998: inst = 32'd471859200;
      1999: inst = 32'd136314880;
      2000: inst = 32'd268468224;
      2001: inst = 32'd201343344;
      2002: inst = 32'd203484854;
      2003: inst = 32'd471859200;
      2004: inst = 32'd136314880;
      2005: inst = 32'd268468224;
      2006: inst = 32'd201343345;
      2007: inst = 32'd203484854;
      2008: inst = 32'd471859200;
      2009: inst = 32'd136314880;
      2010: inst = 32'd268468224;
      2011: inst = 32'd201343346;
      2012: inst = 32'd203484854;
      2013: inst = 32'd471859200;
      2014: inst = 32'd136314880;
      2015: inst = 32'd268468224;
      2016: inst = 32'd201343347;
      2017: inst = 32'd203484854;
      2018: inst = 32'd471859200;
      2019: inst = 32'd136314880;
      2020: inst = 32'd268468224;
      2021: inst = 32'd201343348;
      2022: inst = 32'd203484854;
      2023: inst = 32'd471859200;
      2024: inst = 32'd136314880;
      2025: inst = 32'd268468224;
      2026: inst = 32'd201343349;
      2027: inst = 32'd203484854;
      2028: inst = 32'd471859200;
      2029: inst = 32'd136314880;
      2030: inst = 32'd268468224;
      2031: inst = 32'd201343350;
      2032: inst = 32'd203484854;
      2033: inst = 32'd471859200;
      2034: inst = 32'd136314880;
      2035: inst = 32'd268468224;
      2036: inst = 32'd201343351;
      2037: inst = 32'd203484854;
      2038: inst = 32'd471859200;
      2039: inst = 32'd136314880;
      2040: inst = 32'd268468224;
      2041: inst = 32'd201343352;
      2042: inst = 32'd203484854;
      2043: inst = 32'd471859200;
      2044: inst = 32'd136314880;
      2045: inst = 32'd268468224;
      2046: inst = 32'd201343353;
      2047: inst = 32'd203484854;
      2048: inst = 32'd471859200;
      2049: inst = 32'd136314880;
      2050: inst = 32'd268468224;
      2051: inst = 32'd201343354;
      2052: inst = 32'd203484854;
      2053: inst = 32'd471859200;
      2054: inst = 32'd136314880;
      2055: inst = 32'd268468224;
      2056: inst = 32'd201343355;
      2057: inst = 32'd203484854;
      2058: inst = 32'd471859200;
      2059: inst = 32'd136314880;
      2060: inst = 32'd268468224;
      2061: inst = 32'd201343356;
      2062: inst = 32'd203484854;
      2063: inst = 32'd471859200;
      2064: inst = 32'd136314880;
      2065: inst = 32'd268468224;
      2066: inst = 32'd201343357;
      2067: inst = 32'd203484854;
      2068: inst = 32'd471859200;
      2069: inst = 32'd136314880;
      2070: inst = 32'd268468224;
      2071: inst = 32'd201343358;
      2072: inst = 32'd203484854;
      2073: inst = 32'd471859200;
      2074: inst = 32'd136314880;
      2075: inst = 32'd268468224;
      2076: inst = 32'd201343359;
      2077: inst = 32'd203484854;
      2078: inst = 32'd471859200;
      2079: inst = 32'd136314880;
      2080: inst = 32'd268468224;
      2081: inst = 32'd201343360;
      2082: inst = 32'd203484854;
      2083: inst = 32'd471859200;
      2084: inst = 32'd136314880;
      2085: inst = 32'd268468224;
      2086: inst = 32'd201343361;
      2087: inst = 32'd203484854;
      2088: inst = 32'd471859200;
      2089: inst = 32'd136314880;
      2090: inst = 32'd268468224;
      2091: inst = 32'd201343362;
      2092: inst = 32'd203484854;
      2093: inst = 32'd471859200;
      2094: inst = 32'd136314880;
      2095: inst = 32'd268468224;
      2096: inst = 32'd201343363;
      2097: inst = 32'd203484854;
      2098: inst = 32'd471859200;
      2099: inst = 32'd136314880;
      2100: inst = 32'd268468224;
      2101: inst = 32'd201343364;
      2102: inst = 32'd203484854;
      2103: inst = 32'd471859200;
      2104: inst = 32'd136314880;
      2105: inst = 32'd268468224;
      2106: inst = 32'd201343365;
      2107: inst = 32'd203484854;
      2108: inst = 32'd471859200;
      2109: inst = 32'd136314880;
      2110: inst = 32'd268468224;
      2111: inst = 32'd201343366;
      2112: inst = 32'd203484854;
      2113: inst = 32'd471859200;
      2114: inst = 32'd136314880;
      2115: inst = 32'd268468224;
      2116: inst = 32'd201343367;
      2117: inst = 32'd203484854;
      2118: inst = 32'd471859200;
      2119: inst = 32'd136314880;
      2120: inst = 32'd268468224;
      2121: inst = 32'd201343368;
      2122: inst = 32'd203484854;
      2123: inst = 32'd471859200;
      2124: inst = 32'd136314880;
      2125: inst = 32'd268468224;
      2126: inst = 32'd201343369;
      2127: inst = 32'd203484854;
      2128: inst = 32'd471859200;
      2129: inst = 32'd136314880;
      2130: inst = 32'd268468224;
      2131: inst = 32'd201343370;
      2132: inst = 32'd203484854;
      2133: inst = 32'd471859200;
      2134: inst = 32'd136314880;
      2135: inst = 32'd268468224;
      2136: inst = 32'd201343371;
      2137: inst = 32'd203484854;
      2138: inst = 32'd471859200;
      2139: inst = 32'd136314880;
      2140: inst = 32'd268468224;
      2141: inst = 32'd201343372;
      2142: inst = 32'd203484854;
      2143: inst = 32'd471859200;
      2144: inst = 32'd136314880;
      2145: inst = 32'd268468224;
      2146: inst = 32'd201343373;
      2147: inst = 32'd203484854;
      2148: inst = 32'd471859200;
      2149: inst = 32'd136314880;
      2150: inst = 32'd268468224;
      2151: inst = 32'd201343374;
      2152: inst = 32'd203484854;
      2153: inst = 32'd471859200;
      2154: inst = 32'd136314880;
      2155: inst = 32'd268468224;
      2156: inst = 32'd201343375;
      2157: inst = 32'd203484854;
      2158: inst = 32'd471859200;
      2159: inst = 32'd136314880;
      2160: inst = 32'd268468224;
      2161: inst = 32'd201343376;
      2162: inst = 32'd203484854;
      2163: inst = 32'd471859200;
      2164: inst = 32'd136314880;
      2165: inst = 32'd268468224;
      2166: inst = 32'd201343377;
      2167: inst = 32'd203484854;
      2168: inst = 32'd471859200;
      2169: inst = 32'd136314880;
      2170: inst = 32'd268468224;
      2171: inst = 32'd201343378;
      2172: inst = 32'd203484854;
      2173: inst = 32'd471859200;
      2174: inst = 32'd136314880;
      2175: inst = 32'd268468224;
      2176: inst = 32'd201343379;
      2177: inst = 32'd203484854;
      2178: inst = 32'd471859200;
      2179: inst = 32'd136314880;
      2180: inst = 32'd268468224;
      2181: inst = 32'd201343380;
      2182: inst = 32'd203484854;
      2183: inst = 32'd471859200;
      2184: inst = 32'd136314880;
      2185: inst = 32'd268468224;
      2186: inst = 32'd201343381;
      2187: inst = 32'd203484854;
      2188: inst = 32'd471859200;
      2189: inst = 32'd136314880;
      2190: inst = 32'd268468224;
      2191: inst = 32'd201343382;
      2192: inst = 32'd203484854;
      2193: inst = 32'd471859200;
      2194: inst = 32'd136314880;
      2195: inst = 32'd268468224;
      2196: inst = 32'd201343383;
      2197: inst = 32'd203484854;
      2198: inst = 32'd471859200;
      2199: inst = 32'd136314880;
      2200: inst = 32'd268468224;
      2201: inst = 32'd201343384;
      2202: inst = 32'd203484854;
      2203: inst = 32'd471859200;
      2204: inst = 32'd136314880;
      2205: inst = 32'd268468224;
      2206: inst = 32'd201343385;
      2207: inst = 32'd203484854;
      2208: inst = 32'd471859200;
      2209: inst = 32'd136314880;
      2210: inst = 32'd268468224;
      2211: inst = 32'd201343386;
      2212: inst = 32'd203484854;
      2213: inst = 32'd471859200;
      2214: inst = 32'd136314880;
      2215: inst = 32'd268468224;
      2216: inst = 32'd201343387;
      2217: inst = 32'd203484854;
      2218: inst = 32'd471859200;
      2219: inst = 32'd136314880;
      2220: inst = 32'd268468224;
      2221: inst = 32'd201343388;
      2222: inst = 32'd203484854;
      2223: inst = 32'd471859200;
      2224: inst = 32'd136314880;
      2225: inst = 32'd268468224;
      2226: inst = 32'd201343389;
      2227: inst = 32'd203484854;
      2228: inst = 32'd471859200;
      2229: inst = 32'd136314880;
      2230: inst = 32'd268468224;
      2231: inst = 32'd201343390;
      2232: inst = 32'd203484854;
      2233: inst = 32'd471859200;
      2234: inst = 32'd136314880;
      2235: inst = 32'd268468224;
      2236: inst = 32'd201343391;
      2237: inst = 32'd203484854;
      2238: inst = 32'd471859200;
      2239: inst = 32'd136314880;
      2240: inst = 32'd268468224;
      2241: inst = 32'd201343392;
      2242: inst = 32'd203484854;
      2243: inst = 32'd471859200;
      2244: inst = 32'd136314880;
      2245: inst = 32'd268468224;
      2246: inst = 32'd201343393;
      2247: inst = 32'd203484854;
      2248: inst = 32'd471859200;
      2249: inst = 32'd136314880;
      2250: inst = 32'd268468224;
      2251: inst = 32'd201343394;
      2252: inst = 32'd203484854;
      2253: inst = 32'd471859200;
      2254: inst = 32'd136314880;
      2255: inst = 32'd268468224;
      2256: inst = 32'd201343395;
      2257: inst = 32'd203484854;
      2258: inst = 32'd471859200;
      2259: inst = 32'd136314880;
      2260: inst = 32'd268468224;
      2261: inst = 32'd201343396;
      2262: inst = 32'd203484854;
      2263: inst = 32'd471859200;
      2264: inst = 32'd136314880;
      2265: inst = 32'd268468224;
      2266: inst = 32'd201343397;
      2267: inst = 32'd203484854;
      2268: inst = 32'd471859200;
      2269: inst = 32'd136314880;
      2270: inst = 32'd268468224;
      2271: inst = 32'd201343398;
      2272: inst = 32'd203484854;
      2273: inst = 32'd471859200;
      2274: inst = 32'd136314880;
      2275: inst = 32'd268468224;
      2276: inst = 32'd201343399;
      2277: inst = 32'd203484854;
      2278: inst = 32'd471859200;
      2279: inst = 32'd136314880;
      2280: inst = 32'd268468224;
      2281: inst = 32'd201343400;
      2282: inst = 32'd203484854;
      2283: inst = 32'd471859200;
      2284: inst = 32'd136314880;
      2285: inst = 32'd268468224;
      2286: inst = 32'd201343401;
      2287: inst = 32'd203484854;
      2288: inst = 32'd471859200;
      2289: inst = 32'd136314880;
      2290: inst = 32'd268468224;
      2291: inst = 32'd201343402;
      2292: inst = 32'd203484854;
      2293: inst = 32'd471859200;
      2294: inst = 32'd136314880;
      2295: inst = 32'd268468224;
      2296: inst = 32'd201343403;
      2297: inst = 32'd203484854;
      2298: inst = 32'd471859200;
      2299: inst = 32'd136314880;
      2300: inst = 32'd268468224;
      2301: inst = 32'd201343404;
      2302: inst = 32'd203484854;
      2303: inst = 32'd471859200;
      2304: inst = 32'd136314880;
      2305: inst = 32'd268468224;
      2306: inst = 32'd201343405;
      2307: inst = 32'd203484854;
      2308: inst = 32'd471859200;
      2309: inst = 32'd136314880;
      2310: inst = 32'd268468224;
      2311: inst = 32'd201343406;
      2312: inst = 32'd203484854;
      2313: inst = 32'd471859200;
      2314: inst = 32'd136314880;
      2315: inst = 32'd268468224;
      2316: inst = 32'd201343407;
      2317: inst = 32'd203484854;
      2318: inst = 32'd471859200;
      2319: inst = 32'd136314880;
      2320: inst = 32'd268468224;
      2321: inst = 32'd201343408;
      2322: inst = 32'd203484854;
      2323: inst = 32'd471859200;
      2324: inst = 32'd136314880;
      2325: inst = 32'd268468224;
      2326: inst = 32'd201343409;
      2327: inst = 32'd203484854;
      2328: inst = 32'd471859200;
      2329: inst = 32'd136314880;
      2330: inst = 32'd268468224;
      2331: inst = 32'd201343410;
      2332: inst = 32'd203484854;
      2333: inst = 32'd471859200;
      2334: inst = 32'd136314880;
      2335: inst = 32'd268468224;
      2336: inst = 32'd201343411;
      2337: inst = 32'd203484854;
      2338: inst = 32'd471859200;
      2339: inst = 32'd136314880;
      2340: inst = 32'd268468224;
      2341: inst = 32'd201343412;
      2342: inst = 32'd203484854;
      2343: inst = 32'd471859200;
      2344: inst = 32'd136314880;
      2345: inst = 32'd268468224;
      2346: inst = 32'd201343413;
      2347: inst = 32'd203484854;
      2348: inst = 32'd471859200;
      2349: inst = 32'd136314880;
      2350: inst = 32'd268468224;
      2351: inst = 32'd201343414;
      2352: inst = 32'd203484854;
      2353: inst = 32'd471859200;
      2354: inst = 32'd136314880;
      2355: inst = 32'd268468224;
      2356: inst = 32'd201343415;
      2357: inst = 32'd203484854;
      2358: inst = 32'd471859200;
      2359: inst = 32'd136314880;
      2360: inst = 32'd268468224;
      2361: inst = 32'd201343416;
      2362: inst = 32'd203484854;
      2363: inst = 32'd471859200;
      2364: inst = 32'd136314880;
      2365: inst = 32'd268468224;
      2366: inst = 32'd201343417;
      2367: inst = 32'd203484854;
      2368: inst = 32'd471859200;
      2369: inst = 32'd136314880;
      2370: inst = 32'd268468224;
      2371: inst = 32'd201343418;
      2372: inst = 32'd203484854;
      2373: inst = 32'd471859200;
      2374: inst = 32'd136314880;
      2375: inst = 32'd268468224;
      2376: inst = 32'd201343419;
      2377: inst = 32'd203484854;
      2378: inst = 32'd471859200;
      2379: inst = 32'd136314880;
      2380: inst = 32'd268468224;
      2381: inst = 32'd201343420;
      2382: inst = 32'd203484854;
      2383: inst = 32'd471859200;
      2384: inst = 32'd136314880;
      2385: inst = 32'd268468224;
      2386: inst = 32'd201343421;
      2387: inst = 32'd203484854;
      2388: inst = 32'd471859200;
      2389: inst = 32'd136314880;
      2390: inst = 32'd268468224;
      2391: inst = 32'd201343422;
      2392: inst = 32'd203484854;
      2393: inst = 32'd471859200;
      2394: inst = 32'd136314880;
      2395: inst = 32'd268468224;
      2396: inst = 32'd201343423;
      2397: inst = 32'd203484854;
      2398: inst = 32'd471859200;
      2399: inst = 32'd136314880;
      2400: inst = 32'd268468224;
      2401: inst = 32'd201343424;
      2402: inst = 32'd203484854;
      2403: inst = 32'd471859200;
      2404: inst = 32'd136314880;
      2405: inst = 32'd268468224;
      2406: inst = 32'd201343425;
      2407: inst = 32'd203484854;
      2408: inst = 32'd471859200;
      2409: inst = 32'd136314880;
      2410: inst = 32'd268468224;
      2411: inst = 32'd201343426;
      2412: inst = 32'd203484854;
      2413: inst = 32'd471859200;
      2414: inst = 32'd136314880;
      2415: inst = 32'd268468224;
      2416: inst = 32'd201343427;
      2417: inst = 32'd203484854;
      2418: inst = 32'd471859200;
      2419: inst = 32'd136314880;
      2420: inst = 32'd268468224;
      2421: inst = 32'd201343428;
      2422: inst = 32'd203484854;
      2423: inst = 32'd471859200;
      2424: inst = 32'd136314880;
      2425: inst = 32'd268468224;
      2426: inst = 32'd201343429;
      2427: inst = 32'd203484854;
      2428: inst = 32'd471859200;
      2429: inst = 32'd136314880;
      2430: inst = 32'd268468224;
      2431: inst = 32'd201343430;
      2432: inst = 32'd203484854;
      2433: inst = 32'd471859200;
      2434: inst = 32'd136314880;
      2435: inst = 32'd268468224;
      2436: inst = 32'd201343431;
      2437: inst = 32'd203484854;
      2438: inst = 32'd471859200;
      2439: inst = 32'd136314880;
      2440: inst = 32'd268468224;
      2441: inst = 32'd201343432;
      2442: inst = 32'd203484854;
      2443: inst = 32'd471859200;
      2444: inst = 32'd136314880;
      2445: inst = 32'd268468224;
      2446: inst = 32'd201343433;
      2447: inst = 32'd203484854;
      2448: inst = 32'd471859200;
      2449: inst = 32'd136314880;
      2450: inst = 32'd268468224;
      2451: inst = 32'd201343434;
      2452: inst = 32'd203484854;
      2453: inst = 32'd471859200;
      2454: inst = 32'd136314880;
      2455: inst = 32'd268468224;
      2456: inst = 32'd201343435;
      2457: inst = 32'd203461810;
      2458: inst = 32'd471859200;
      2459: inst = 32'd136314880;
      2460: inst = 32'd268468224;
      2461: inst = 32'd201343436;
      2462: inst = 32'd203484854;
      2463: inst = 32'd471859200;
      2464: inst = 32'd136314880;
      2465: inst = 32'd268468224;
      2466: inst = 32'd201343437;
      2467: inst = 32'd203484854;
      2468: inst = 32'd471859200;
      2469: inst = 32'd136314880;
      2470: inst = 32'd268468224;
      2471: inst = 32'd201343438;
      2472: inst = 32'd203484854;
      2473: inst = 32'd471859200;
      2474: inst = 32'd136314880;
      2475: inst = 32'd268468224;
      2476: inst = 32'd201343439;
      2477: inst = 32'd203484854;
      2478: inst = 32'd471859200;
      2479: inst = 32'd136314880;
      2480: inst = 32'd268468224;
      2481: inst = 32'd201343440;
      2482: inst = 32'd203484854;
      2483: inst = 32'd471859200;
      2484: inst = 32'd136314880;
      2485: inst = 32'd268468224;
      2486: inst = 32'd201343441;
      2487: inst = 32'd203484854;
      2488: inst = 32'd471859200;
      2489: inst = 32'd136314880;
      2490: inst = 32'd268468224;
      2491: inst = 32'd201343442;
      2492: inst = 32'd203484854;
      2493: inst = 32'd471859200;
      2494: inst = 32'd136314880;
      2495: inst = 32'd268468224;
      2496: inst = 32'd201343443;
      2497: inst = 32'd203484854;
      2498: inst = 32'd471859200;
      2499: inst = 32'd136314880;
      2500: inst = 32'd268468224;
      2501: inst = 32'd201343444;
      2502: inst = 32'd203484854;
      2503: inst = 32'd471859200;
      2504: inst = 32'd136314880;
      2505: inst = 32'd268468224;
      2506: inst = 32'd201343445;
      2507: inst = 32'd203484854;
      2508: inst = 32'd471859200;
      2509: inst = 32'd136314880;
      2510: inst = 32'd268468224;
      2511: inst = 32'd201343446;
      2512: inst = 32'd203484854;
      2513: inst = 32'd471859200;
      2514: inst = 32'd136314880;
      2515: inst = 32'd268468224;
      2516: inst = 32'd201343447;
      2517: inst = 32'd203484854;
      2518: inst = 32'd471859200;
      2519: inst = 32'd136314880;
      2520: inst = 32'd268468224;
      2521: inst = 32'd201343448;
      2522: inst = 32'd203484854;
      2523: inst = 32'd471859200;
      2524: inst = 32'd136314880;
      2525: inst = 32'd268468224;
      2526: inst = 32'd201343449;
      2527: inst = 32'd203484854;
      2528: inst = 32'd471859200;
      2529: inst = 32'd136314880;
      2530: inst = 32'd268468224;
      2531: inst = 32'd201343450;
      2532: inst = 32'd203470230;
      2533: inst = 32'd471859200;
      2534: inst = 32'd136314880;
      2535: inst = 32'd268468224;
      2536: inst = 32'd201343451;
      2537: inst = 32'd203470230;
      2538: inst = 32'd471859200;
      2539: inst = 32'd136314880;
      2540: inst = 32'd268468224;
      2541: inst = 32'd201343452;
      2542: inst = 32'd203470230;
      2543: inst = 32'd471859200;
      2544: inst = 32'd136314880;
      2545: inst = 32'd268468224;
      2546: inst = 32'd201343453;
      2547: inst = 32'd203470230;
      2548: inst = 32'd471859200;
      2549: inst = 32'd136314880;
      2550: inst = 32'd268468224;
      2551: inst = 32'd201343454;
      2552: inst = 32'd203470230;
      2553: inst = 32'd471859200;
      2554: inst = 32'd136314880;
      2555: inst = 32'd268468224;
      2556: inst = 32'd201343455;
      2557: inst = 32'd203470230;
      2558: inst = 32'd471859200;
      2559: inst = 32'd136314880;
      2560: inst = 32'd268468224;
      2561: inst = 32'd201343456;
      2562: inst = 32'd203470230;
      2563: inst = 32'd471859200;
      2564: inst = 32'd136314880;
      2565: inst = 32'd268468224;
      2566: inst = 32'd201343457;
      2567: inst = 32'd203470230;
      2568: inst = 32'd471859200;
      2569: inst = 32'd136314880;
      2570: inst = 32'd268468224;
      2571: inst = 32'd201343458;
      2572: inst = 32'd203470230;
      2573: inst = 32'd471859200;
      2574: inst = 32'd136314880;
      2575: inst = 32'd268468224;
      2576: inst = 32'd201343459;
      2577: inst = 32'd203470230;
      2578: inst = 32'd471859200;
      2579: inst = 32'd136314880;
      2580: inst = 32'd268468224;
      2581: inst = 32'd201343460;
      2582: inst = 32'd203470230;
      2583: inst = 32'd471859200;
      2584: inst = 32'd136314880;
      2585: inst = 32'd268468224;
      2586: inst = 32'd201343461;
      2587: inst = 32'd203470230;
      2588: inst = 32'd471859200;
      2589: inst = 32'd136314880;
      2590: inst = 32'd268468224;
      2591: inst = 32'd201343462;
      2592: inst = 32'd203470230;
      2593: inst = 32'd471859200;
      2594: inst = 32'd136314880;
      2595: inst = 32'd268468224;
      2596: inst = 32'd201343463;
      2597: inst = 32'd203470230;
      2598: inst = 32'd471859200;
      2599: inst = 32'd136314880;
      2600: inst = 32'd268468224;
      2601: inst = 32'd201343464;
      2602: inst = 32'd203470230;
      2603: inst = 32'd471859200;
      2604: inst = 32'd136314880;
      2605: inst = 32'd268468224;
      2606: inst = 32'd201343465;
      2607: inst = 32'd203470230;
      2608: inst = 32'd471859200;
      2609: inst = 32'd136314880;
      2610: inst = 32'd268468224;
      2611: inst = 32'd201343466;
      2612: inst = 32'd203470230;
      2613: inst = 32'd471859200;
      2614: inst = 32'd136314880;
      2615: inst = 32'd268468224;
      2616: inst = 32'd201343467;
      2617: inst = 32'd203470230;
      2618: inst = 32'd471859200;
      2619: inst = 32'd136314880;
      2620: inst = 32'd268468224;
      2621: inst = 32'd201343468;
      2622: inst = 32'd203470230;
      2623: inst = 32'd471859200;
      2624: inst = 32'd136314880;
      2625: inst = 32'd268468224;
      2626: inst = 32'd201343469;
      2627: inst = 32'd203470230;
      2628: inst = 32'd471859200;
      2629: inst = 32'd136314880;
      2630: inst = 32'd268468224;
      2631: inst = 32'd201343470;
      2632: inst = 32'd203470230;
      2633: inst = 32'd471859200;
      2634: inst = 32'd136314880;
      2635: inst = 32'd268468224;
      2636: inst = 32'd201343471;
      2637: inst = 32'd203470230;
      2638: inst = 32'd471859200;
      2639: inst = 32'd136314880;
      2640: inst = 32'd268468224;
      2641: inst = 32'd201343472;
      2642: inst = 32'd203470230;
      2643: inst = 32'd471859200;
      2644: inst = 32'd136314880;
      2645: inst = 32'd268468224;
      2646: inst = 32'd201343473;
      2647: inst = 32'd203470230;
      2648: inst = 32'd471859200;
      2649: inst = 32'd136314880;
      2650: inst = 32'd268468224;
      2651: inst = 32'd201343474;
      2652: inst = 32'd203470230;
      2653: inst = 32'd471859200;
      2654: inst = 32'd136314880;
      2655: inst = 32'd268468224;
      2656: inst = 32'd201343475;
      2657: inst = 32'd203470230;
      2658: inst = 32'd471859200;
      2659: inst = 32'd136314880;
      2660: inst = 32'd268468224;
      2661: inst = 32'd201343476;
      2662: inst = 32'd203470230;
      2663: inst = 32'd471859200;
      2664: inst = 32'd136314880;
      2665: inst = 32'd268468224;
      2666: inst = 32'd201343477;
      2667: inst = 32'd203470230;
      2668: inst = 32'd471859200;
      2669: inst = 32'd136314880;
      2670: inst = 32'd268468224;
      2671: inst = 32'd201343478;
      2672: inst = 32'd203470230;
      2673: inst = 32'd471859200;
      2674: inst = 32'd136314880;
      2675: inst = 32'd268468224;
      2676: inst = 32'd201343479;
      2677: inst = 32'd203470230;
      2678: inst = 32'd471859200;
      2679: inst = 32'd136314880;
      2680: inst = 32'd268468224;
      2681: inst = 32'd201343480;
      2682: inst = 32'd203470230;
      2683: inst = 32'd471859200;
      2684: inst = 32'd136314880;
      2685: inst = 32'd268468224;
      2686: inst = 32'd201343481;
      2687: inst = 32'd203470230;
      2688: inst = 32'd471859200;
      2689: inst = 32'd136314880;
      2690: inst = 32'd268468224;
      2691: inst = 32'd201343482;
      2692: inst = 32'd203470230;
      2693: inst = 32'd471859200;
      2694: inst = 32'd136314880;
      2695: inst = 32'd268468224;
      2696: inst = 32'd201343483;
      2697: inst = 32'd203470230;
      2698: inst = 32'd471859200;
      2699: inst = 32'd136314880;
      2700: inst = 32'd268468224;
      2701: inst = 32'd201343484;
      2702: inst = 32'd203470230;
      2703: inst = 32'd471859200;
      2704: inst = 32'd136314880;
      2705: inst = 32'd268468224;
      2706: inst = 32'd201343485;
      2707: inst = 32'd203470230;
      2708: inst = 32'd471859200;
      2709: inst = 32'd136314880;
      2710: inst = 32'd268468224;
      2711: inst = 32'd201343486;
      2712: inst = 32'd203470230;
      2713: inst = 32'd471859200;
      2714: inst = 32'd136314880;
      2715: inst = 32'd268468224;
      2716: inst = 32'd201343487;
      2717: inst = 32'd203470230;
      2718: inst = 32'd471859200;
      2719: inst = 32'd136314880;
      2720: inst = 32'd268468224;
      2721: inst = 32'd201343488;
      2722: inst = 32'd203470230;
      2723: inst = 32'd471859200;
      2724: inst = 32'd136314880;
      2725: inst = 32'd268468224;
      2726: inst = 32'd201343489;
      2727: inst = 32'd203470230;
      2728: inst = 32'd471859200;
      2729: inst = 32'd136314880;
      2730: inst = 32'd268468224;
      2731: inst = 32'd201343490;
      2732: inst = 32'd203470230;
      2733: inst = 32'd471859200;
      2734: inst = 32'd136314880;
      2735: inst = 32'd268468224;
      2736: inst = 32'd201343491;
      2737: inst = 32'd203470230;
      2738: inst = 32'd471859200;
      2739: inst = 32'd136314880;
      2740: inst = 32'd268468224;
      2741: inst = 32'd201343492;
      2742: inst = 32'd203470230;
      2743: inst = 32'd471859200;
      2744: inst = 32'd136314880;
      2745: inst = 32'd268468224;
      2746: inst = 32'd201343493;
      2747: inst = 32'd203470230;
      2748: inst = 32'd471859200;
      2749: inst = 32'd136314880;
      2750: inst = 32'd268468224;
      2751: inst = 32'd201343494;
      2752: inst = 32'd203484854;
      2753: inst = 32'd471859200;
      2754: inst = 32'd136314880;
      2755: inst = 32'd268468224;
      2756: inst = 32'd201343495;
      2757: inst = 32'd203484854;
      2758: inst = 32'd471859200;
      2759: inst = 32'd136314880;
      2760: inst = 32'd268468224;
      2761: inst = 32'd201343496;
      2762: inst = 32'd203484854;
      2763: inst = 32'd471859200;
      2764: inst = 32'd136314880;
      2765: inst = 32'd268468224;
      2766: inst = 32'd201343497;
      2767: inst = 32'd203484854;
      2768: inst = 32'd471859200;
      2769: inst = 32'd136314880;
      2770: inst = 32'd268468224;
      2771: inst = 32'd201343498;
      2772: inst = 32'd203484854;
      2773: inst = 32'd471859200;
      2774: inst = 32'd136314880;
      2775: inst = 32'd268468224;
      2776: inst = 32'd201343499;
      2777: inst = 32'd203484854;
      2778: inst = 32'd471859200;
      2779: inst = 32'd136314880;
      2780: inst = 32'd268468224;
      2781: inst = 32'd201343500;
      2782: inst = 32'd203484854;
      2783: inst = 32'd471859200;
      2784: inst = 32'd136314880;
      2785: inst = 32'd268468224;
      2786: inst = 32'd201343501;
      2787: inst = 32'd203484854;
      2788: inst = 32'd471859200;
      2789: inst = 32'd136314880;
      2790: inst = 32'd268468224;
      2791: inst = 32'd201343502;
      2792: inst = 32'd203484854;
      2793: inst = 32'd471859200;
      2794: inst = 32'd136314880;
      2795: inst = 32'd268468224;
      2796: inst = 32'd201343503;
      2797: inst = 32'd203484854;
      2798: inst = 32'd471859200;
      2799: inst = 32'd136314880;
      2800: inst = 32'd268468224;
      2801: inst = 32'd201343504;
      2802: inst = 32'd203484854;
      2803: inst = 32'd471859200;
      2804: inst = 32'd136314880;
      2805: inst = 32'd268468224;
      2806: inst = 32'd201343505;
      2807: inst = 32'd203484854;
      2808: inst = 32'd471859200;
      2809: inst = 32'd136314880;
      2810: inst = 32'd268468224;
      2811: inst = 32'd201343506;
      2812: inst = 32'd203484854;
      2813: inst = 32'd471859200;
      2814: inst = 32'd136314880;
      2815: inst = 32'd268468224;
      2816: inst = 32'd201343507;
      2817: inst = 32'd203484854;
      2818: inst = 32'd471859200;
      2819: inst = 32'd136314880;
      2820: inst = 32'd268468224;
      2821: inst = 32'd201343508;
      2822: inst = 32'd203484854;
      2823: inst = 32'd471859200;
      2824: inst = 32'd136314880;
      2825: inst = 32'd268468224;
      2826: inst = 32'd201343509;
      2827: inst = 32'd203484854;
      2828: inst = 32'd471859200;
      2829: inst = 32'd136314880;
      2830: inst = 32'd268468224;
      2831: inst = 32'd201343510;
      2832: inst = 32'd203484854;
      2833: inst = 32'd471859200;
      2834: inst = 32'd136314880;
      2835: inst = 32'd268468224;
      2836: inst = 32'd201343511;
      2837: inst = 32'd203484854;
      2838: inst = 32'd471859200;
      2839: inst = 32'd136314880;
      2840: inst = 32'd268468224;
      2841: inst = 32'd201343512;
      2842: inst = 32'd203484854;
      2843: inst = 32'd471859200;
      2844: inst = 32'd136314880;
      2845: inst = 32'd268468224;
      2846: inst = 32'd201343513;
      2847: inst = 32'd203484854;
      2848: inst = 32'd471859200;
      2849: inst = 32'd136314880;
      2850: inst = 32'd268468224;
      2851: inst = 32'd201343514;
      2852: inst = 32'd203484854;
      2853: inst = 32'd471859200;
      2854: inst = 32'd136314880;
      2855: inst = 32'd268468224;
      2856: inst = 32'd201343515;
      2857: inst = 32'd203484854;
      2858: inst = 32'd471859200;
      2859: inst = 32'd136314880;
      2860: inst = 32'd268468224;
      2861: inst = 32'd201343516;
      2862: inst = 32'd203484854;
      2863: inst = 32'd471859200;
      2864: inst = 32'd136314880;
      2865: inst = 32'd268468224;
      2866: inst = 32'd201343517;
      2867: inst = 32'd203484854;
      2868: inst = 32'd471859200;
      2869: inst = 32'd136314880;
      2870: inst = 32'd268468224;
      2871: inst = 32'd201343518;
      2872: inst = 32'd203484854;
      2873: inst = 32'd471859200;
      2874: inst = 32'd136314880;
      2875: inst = 32'd268468224;
      2876: inst = 32'd201343519;
      2877: inst = 32'd203484854;
      2878: inst = 32'd471859200;
      2879: inst = 32'd136314880;
      2880: inst = 32'd268468224;
      2881: inst = 32'd201343520;
      2882: inst = 32'd203484854;
      2883: inst = 32'd471859200;
      2884: inst = 32'd136314880;
      2885: inst = 32'd268468224;
      2886: inst = 32'd201343521;
      2887: inst = 32'd203484854;
      2888: inst = 32'd471859200;
      2889: inst = 32'd136314880;
      2890: inst = 32'd268468224;
      2891: inst = 32'd201343522;
      2892: inst = 32'd203484854;
      2893: inst = 32'd471859200;
      2894: inst = 32'd136314880;
      2895: inst = 32'd268468224;
      2896: inst = 32'd201343523;
      2897: inst = 32'd203484854;
      2898: inst = 32'd471859200;
      2899: inst = 32'd136314880;
      2900: inst = 32'd268468224;
      2901: inst = 32'd201343524;
      2902: inst = 32'd203484854;
      2903: inst = 32'd471859200;
      2904: inst = 32'd136314880;
      2905: inst = 32'd268468224;
      2906: inst = 32'd201343525;
      2907: inst = 32'd203484854;
      2908: inst = 32'd471859200;
      2909: inst = 32'd136314880;
      2910: inst = 32'd268468224;
      2911: inst = 32'd201343526;
      2912: inst = 32'd203484854;
      2913: inst = 32'd471859200;
      2914: inst = 32'd136314880;
      2915: inst = 32'd268468224;
      2916: inst = 32'd201343527;
      2917: inst = 32'd203484854;
      2918: inst = 32'd471859200;
      2919: inst = 32'd136314880;
      2920: inst = 32'd268468224;
      2921: inst = 32'd201343528;
      2922: inst = 32'd203484854;
      2923: inst = 32'd471859200;
      2924: inst = 32'd136314880;
      2925: inst = 32'd268468224;
      2926: inst = 32'd201343529;
      2927: inst = 32'd203484854;
      2928: inst = 32'd471859200;
      2929: inst = 32'd136314880;
      2930: inst = 32'd268468224;
      2931: inst = 32'd201343530;
      2932: inst = 32'd203484854;
      2933: inst = 32'd471859200;
      2934: inst = 32'd136314880;
      2935: inst = 32'd268468224;
      2936: inst = 32'd201343531;
      2937: inst = 32'd203461810;
      2938: inst = 32'd471859200;
      2939: inst = 32'd136314880;
      2940: inst = 32'd268468224;
      2941: inst = 32'd201343532;
      2942: inst = 32'd203484854;
      2943: inst = 32'd471859200;
      2944: inst = 32'd136314880;
      2945: inst = 32'd268468224;
      2946: inst = 32'd201343533;
      2947: inst = 32'd203484854;
      2948: inst = 32'd471859200;
      2949: inst = 32'd136314880;
      2950: inst = 32'd268468224;
      2951: inst = 32'd201343534;
      2952: inst = 32'd203484854;
      2953: inst = 32'd471859200;
      2954: inst = 32'd136314880;
      2955: inst = 32'd268468224;
      2956: inst = 32'd201343535;
      2957: inst = 32'd203484854;
      2958: inst = 32'd471859200;
      2959: inst = 32'd136314880;
      2960: inst = 32'd268468224;
      2961: inst = 32'd201343536;
      2962: inst = 32'd203484854;
      2963: inst = 32'd471859200;
      2964: inst = 32'd136314880;
      2965: inst = 32'd268468224;
      2966: inst = 32'd201343537;
      2967: inst = 32'd203484854;
      2968: inst = 32'd471859200;
      2969: inst = 32'd136314880;
      2970: inst = 32'd268468224;
      2971: inst = 32'd201343538;
      2972: inst = 32'd203484854;
      2973: inst = 32'd471859200;
      2974: inst = 32'd136314880;
      2975: inst = 32'd268468224;
      2976: inst = 32'd201343539;
      2977: inst = 32'd203484854;
      2978: inst = 32'd471859200;
      2979: inst = 32'd136314880;
      2980: inst = 32'd268468224;
      2981: inst = 32'd201343540;
      2982: inst = 32'd203484854;
      2983: inst = 32'd471859200;
      2984: inst = 32'd136314880;
      2985: inst = 32'd268468224;
      2986: inst = 32'd201343541;
      2987: inst = 32'd203484854;
      2988: inst = 32'd471859200;
      2989: inst = 32'd136314880;
      2990: inst = 32'd268468224;
      2991: inst = 32'd201343542;
      2992: inst = 32'd203484854;
      2993: inst = 32'd471859200;
      2994: inst = 32'd136314880;
      2995: inst = 32'd268468224;
      2996: inst = 32'd201343543;
      2997: inst = 32'd203484854;
      2998: inst = 32'd471859200;
      2999: inst = 32'd136314880;
      3000: inst = 32'd268468224;
      3001: inst = 32'd201343544;
      3002: inst = 32'd203484854;
      3003: inst = 32'd471859200;
      3004: inst = 32'd136314880;
      3005: inst = 32'd268468224;
      3006: inst = 32'd201343545;
      3007: inst = 32'd203484854;
      3008: inst = 32'd471859200;
      3009: inst = 32'd136314880;
      3010: inst = 32'd268468224;
      3011: inst = 32'd201343546;
      3012: inst = 32'd203484854;
      3013: inst = 32'd471859200;
      3014: inst = 32'd136314880;
      3015: inst = 32'd268468224;
      3016: inst = 32'd201343547;
      3017: inst = 32'd203484854;
      3018: inst = 32'd471859200;
      3019: inst = 32'd136314880;
      3020: inst = 32'd268468224;
      3021: inst = 32'd201343548;
      3022: inst = 32'd203489279;
      3023: inst = 32'd471859200;
      3024: inst = 32'd136314880;
      3025: inst = 32'd268468224;
      3026: inst = 32'd201343549;
      3027: inst = 32'd203489279;
      3028: inst = 32'd471859200;
      3029: inst = 32'd136314880;
      3030: inst = 32'd268468224;
      3031: inst = 32'd201343550;
      3032: inst = 32'd203489279;
      3033: inst = 32'd471859200;
      3034: inst = 32'd136314880;
      3035: inst = 32'd268468224;
      3036: inst = 32'd201343551;
      3037: inst = 32'd203489279;
      3038: inst = 32'd471859200;
      3039: inst = 32'd136314880;
      3040: inst = 32'd268468224;
      3041: inst = 32'd201343552;
      3042: inst = 32'd203489279;
      3043: inst = 32'd471859200;
      3044: inst = 32'd136314880;
      3045: inst = 32'd268468224;
      3046: inst = 32'd201343553;
      3047: inst = 32'd203489279;
      3048: inst = 32'd471859200;
      3049: inst = 32'd136314880;
      3050: inst = 32'd268468224;
      3051: inst = 32'd201343554;
      3052: inst = 32'd203489279;
      3053: inst = 32'd471859200;
      3054: inst = 32'd136314880;
      3055: inst = 32'd268468224;
      3056: inst = 32'd201343555;
      3057: inst = 32'd203489279;
      3058: inst = 32'd471859200;
      3059: inst = 32'd136314880;
      3060: inst = 32'd268468224;
      3061: inst = 32'd201343556;
      3062: inst = 32'd203489279;
      3063: inst = 32'd471859200;
      3064: inst = 32'd136314880;
      3065: inst = 32'd268468224;
      3066: inst = 32'd201343557;
      3067: inst = 32'd203489279;
      3068: inst = 32'd471859200;
      3069: inst = 32'd136314880;
      3070: inst = 32'd268468224;
      3071: inst = 32'd201343558;
      3072: inst = 32'd203489279;
      3073: inst = 32'd471859200;
      3074: inst = 32'd136314880;
      3075: inst = 32'd268468224;
      3076: inst = 32'd201343559;
      3077: inst = 32'd203489279;
      3078: inst = 32'd471859200;
      3079: inst = 32'd136314880;
      3080: inst = 32'd268468224;
      3081: inst = 32'd201343560;
      3082: inst = 32'd203489279;
      3083: inst = 32'd471859200;
      3084: inst = 32'd136314880;
      3085: inst = 32'd268468224;
      3086: inst = 32'd201343561;
      3087: inst = 32'd203489279;
      3088: inst = 32'd471859200;
      3089: inst = 32'd136314880;
      3090: inst = 32'd268468224;
      3091: inst = 32'd201343562;
      3092: inst = 32'd203489279;
      3093: inst = 32'd471859200;
      3094: inst = 32'd136314880;
      3095: inst = 32'd268468224;
      3096: inst = 32'd201343563;
      3097: inst = 32'd203489279;
      3098: inst = 32'd471859200;
      3099: inst = 32'd136314880;
      3100: inst = 32'd268468224;
      3101: inst = 32'd201343564;
      3102: inst = 32'd203489279;
      3103: inst = 32'd471859200;
      3104: inst = 32'd136314880;
      3105: inst = 32'd268468224;
      3106: inst = 32'd201343565;
      3107: inst = 32'd203489279;
      3108: inst = 32'd471859200;
      3109: inst = 32'd136314880;
      3110: inst = 32'd268468224;
      3111: inst = 32'd201343566;
      3112: inst = 32'd203489279;
      3113: inst = 32'd471859200;
      3114: inst = 32'd136314880;
      3115: inst = 32'd268468224;
      3116: inst = 32'd201343567;
      3117: inst = 32'd203489279;
      3118: inst = 32'd471859200;
      3119: inst = 32'd136314880;
      3120: inst = 32'd268468224;
      3121: inst = 32'd201343568;
      3122: inst = 32'd203489279;
      3123: inst = 32'd471859200;
      3124: inst = 32'd136314880;
      3125: inst = 32'd268468224;
      3126: inst = 32'd201343569;
      3127: inst = 32'd203489279;
      3128: inst = 32'd471859200;
      3129: inst = 32'd136314880;
      3130: inst = 32'd268468224;
      3131: inst = 32'd201343570;
      3132: inst = 32'd203489279;
      3133: inst = 32'd471859200;
      3134: inst = 32'd136314880;
      3135: inst = 32'd268468224;
      3136: inst = 32'd201343571;
      3137: inst = 32'd203489279;
      3138: inst = 32'd471859200;
      3139: inst = 32'd136314880;
      3140: inst = 32'd268468224;
      3141: inst = 32'd201343572;
      3142: inst = 32'd203489279;
      3143: inst = 32'd471859200;
      3144: inst = 32'd136314880;
      3145: inst = 32'd268468224;
      3146: inst = 32'd201343573;
      3147: inst = 32'd203489279;
      3148: inst = 32'd471859200;
      3149: inst = 32'd136314880;
      3150: inst = 32'd268468224;
      3151: inst = 32'd201343574;
      3152: inst = 32'd203489279;
      3153: inst = 32'd471859200;
      3154: inst = 32'd136314880;
      3155: inst = 32'd268468224;
      3156: inst = 32'd201343575;
      3157: inst = 32'd203489279;
      3158: inst = 32'd471859200;
      3159: inst = 32'd136314880;
      3160: inst = 32'd268468224;
      3161: inst = 32'd201343576;
      3162: inst = 32'd203489279;
      3163: inst = 32'd471859200;
      3164: inst = 32'd136314880;
      3165: inst = 32'd268468224;
      3166: inst = 32'd201343577;
      3167: inst = 32'd203489279;
      3168: inst = 32'd471859200;
      3169: inst = 32'd136314880;
      3170: inst = 32'd268468224;
      3171: inst = 32'd201343578;
      3172: inst = 32'd203489279;
      3173: inst = 32'd471859200;
      3174: inst = 32'd136314880;
      3175: inst = 32'd268468224;
      3176: inst = 32'd201343579;
      3177: inst = 32'd203489279;
      3178: inst = 32'd471859200;
      3179: inst = 32'd136314880;
      3180: inst = 32'd268468224;
      3181: inst = 32'd201343580;
      3182: inst = 32'd203489279;
      3183: inst = 32'd471859200;
      3184: inst = 32'd136314880;
      3185: inst = 32'd268468224;
      3186: inst = 32'd201343581;
      3187: inst = 32'd203489279;
      3188: inst = 32'd471859200;
      3189: inst = 32'd136314880;
      3190: inst = 32'd268468224;
      3191: inst = 32'd201343582;
      3192: inst = 32'd203489279;
      3193: inst = 32'd471859200;
      3194: inst = 32'd136314880;
      3195: inst = 32'd268468224;
      3196: inst = 32'd201343583;
      3197: inst = 32'd203489279;
      3198: inst = 32'd471859200;
      3199: inst = 32'd136314880;
      3200: inst = 32'd268468224;
      3201: inst = 32'd201343584;
      3202: inst = 32'd203489279;
      3203: inst = 32'd471859200;
      3204: inst = 32'd136314880;
      3205: inst = 32'd268468224;
      3206: inst = 32'd201343585;
      3207: inst = 32'd203489279;
      3208: inst = 32'd471859200;
      3209: inst = 32'd136314880;
      3210: inst = 32'd268468224;
      3211: inst = 32'd201343586;
      3212: inst = 32'd203489279;
      3213: inst = 32'd471859200;
      3214: inst = 32'd136314880;
      3215: inst = 32'd268468224;
      3216: inst = 32'd201343587;
      3217: inst = 32'd203489279;
      3218: inst = 32'd471859200;
      3219: inst = 32'd136314880;
      3220: inst = 32'd268468224;
      3221: inst = 32'd201343588;
      3222: inst = 32'd203484854;
      3223: inst = 32'd471859200;
      3224: inst = 32'd136314880;
      3225: inst = 32'd268468224;
      3226: inst = 32'd201343589;
      3227: inst = 32'd203484854;
      3228: inst = 32'd471859200;
      3229: inst = 32'd136314880;
      3230: inst = 32'd268468224;
      3231: inst = 32'd201343590;
      3232: inst = 32'd203484854;
      3233: inst = 32'd471859200;
      3234: inst = 32'd136314880;
      3235: inst = 32'd268468224;
      3236: inst = 32'd201343591;
      3237: inst = 32'd203484854;
      3238: inst = 32'd471859200;
      3239: inst = 32'd136314880;
      3240: inst = 32'd268468224;
      3241: inst = 32'd201343592;
      3242: inst = 32'd203484854;
      3243: inst = 32'd471859200;
      3244: inst = 32'd136314880;
      3245: inst = 32'd268468224;
      3246: inst = 32'd201343593;
      3247: inst = 32'd203484854;
      3248: inst = 32'd471859200;
      3249: inst = 32'd136314880;
      3250: inst = 32'd268468224;
      3251: inst = 32'd201343594;
      3252: inst = 32'd203484854;
      3253: inst = 32'd471859200;
      3254: inst = 32'd136314880;
      3255: inst = 32'd268468224;
      3256: inst = 32'd201343595;
      3257: inst = 32'd203484854;
      3258: inst = 32'd471859200;
      3259: inst = 32'd136314880;
      3260: inst = 32'd268468224;
      3261: inst = 32'd201343596;
      3262: inst = 32'd203484854;
      3263: inst = 32'd471859200;
      3264: inst = 32'd136314880;
      3265: inst = 32'd268468224;
      3266: inst = 32'd201343597;
      3267: inst = 32'd203484854;
      3268: inst = 32'd471859200;
      3269: inst = 32'd136314880;
      3270: inst = 32'd268468224;
      3271: inst = 32'd201343598;
      3272: inst = 32'd203484854;
      3273: inst = 32'd471859200;
      3274: inst = 32'd136314880;
      3275: inst = 32'd268468224;
      3276: inst = 32'd201343599;
      3277: inst = 32'd203484854;
      3278: inst = 32'd471859200;
      3279: inst = 32'd136314880;
      3280: inst = 32'd268468224;
      3281: inst = 32'd201343600;
      3282: inst = 32'd203484854;
      3283: inst = 32'd471859200;
      3284: inst = 32'd136314880;
      3285: inst = 32'd268468224;
      3286: inst = 32'd201343601;
      3287: inst = 32'd203484854;
      3288: inst = 32'd471859200;
      3289: inst = 32'd136314880;
      3290: inst = 32'd268468224;
      3291: inst = 32'd201343602;
      3292: inst = 32'd203484854;
      3293: inst = 32'd471859200;
      3294: inst = 32'd136314880;
      3295: inst = 32'd268468224;
      3296: inst = 32'd201343603;
      3297: inst = 32'd203484854;
      3298: inst = 32'd471859200;
      3299: inst = 32'd136314880;
      3300: inst = 32'd268468224;
      3301: inst = 32'd201343604;
      3302: inst = 32'd203484854;
      3303: inst = 32'd471859200;
      3304: inst = 32'd136314880;
      3305: inst = 32'd268468224;
      3306: inst = 32'd201343605;
      3307: inst = 32'd203484854;
      3308: inst = 32'd471859200;
      3309: inst = 32'd136314880;
      3310: inst = 32'd268468224;
      3311: inst = 32'd201343606;
      3312: inst = 32'd203484854;
      3313: inst = 32'd471859200;
      3314: inst = 32'd136314880;
      3315: inst = 32'd268468224;
      3316: inst = 32'd201343607;
      3317: inst = 32'd203484854;
      3318: inst = 32'd471859200;
      3319: inst = 32'd136314880;
      3320: inst = 32'd268468224;
      3321: inst = 32'd201343608;
      3322: inst = 32'd203484854;
      3323: inst = 32'd471859200;
      3324: inst = 32'd136314880;
      3325: inst = 32'd268468224;
      3326: inst = 32'd201343609;
      3327: inst = 32'd203484854;
      3328: inst = 32'd471859200;
      3329: inst = 32'd136314880;
      3330: inst = 32'd268468224;
      3331: inst = 32'd201343610;
      3332: inst = 32'd203484854;
      3333: inst = 32'd471859200;
      3334: inst = 32'd136314880;
      3335: inst = 32'd268468224;
      3336: inst = 32'd201343611;
      3337: inst = 32'd203484854;
      3338: inst = 32'd471859200;
      3339: inst = 32'd136314880;
      3340: inst = 32'd268468224;
      3341: inst = 32'd201343612;
      3342: inst = 32'd203484854;
      3343: inst = 32'd471859200;
      3344: inst = 32'd136314880;
      3345: inst = 32'd268468224;
      3346: inst = 32'd201343613;
      3347: inst = 32'd203484854;
      3348: inst = 32'd471859200;
      3349: inst = 32'd136314880;
      3350: inst = 32'd268468224;
      3351: inst = 32'd201343614;
      3352: inst = 32'd203484854;
      3353: inst = 32'd471859200;
      3354: inst = 32'd136314880;
      3355: inst = 32'd268468224;
      3356: inst = 32'd201343615;
      3357: inst = 32'd203484854;
      3358: inst = 32'd471859200;
      3359: inst = 32'd136314880;
      3360: inst = 32'd268468224;
      3361: inst = 32'd201343616;
      3362: inst = 32'd203484854;
      3363: inst = 32'd471859200;
      3364: inst = 32'd136314880;
      3365: inst = 32'd268468224;
      3366: inst = 32'd201343617;
      3367: inst = 32'd203484854;
      3368: inst = 32'd471859200;
      3369: inst = 32'd136314880;
      3370: inst = 32'd268468224;
      3371: inst = 32'd201343618;
      3372: inst = 32'd203484854;
      3373: inst = 32'd471859200;
      3374: inst = 32'd136314880;
      3375: inst = 32'd268468224;
      3376: inst = 32'd201343619;
      3377: inst = 32'd203484854;
      3378: inst = 32'd471859200;
      3379: inst = 32'd136314880;
      3380: inst = 32'd268468224;
      3381: inst = 32'd201343620;
      3382: inst = 32'd203484854;
      3383: inst = 32'd471859200;
      3384: inst = 32'd136314880;
      3385: inst = 32'd268468224;
      3386: inst = 32'd201343621;
      3387: inst = 32'd203484854;
      3388: inst = 32'd471859200;
      3389: inst = 32'd136314880;
      3390: inst = 32'd268468224;
      3391: inst = 32'd201343622;
      3392: inst = 32'd203484854;
      3393: inst = 32'd471859200;
      3394: inst = 32'd136314880;
      3395: inst = 32'd268468224;
      3396: inst = 32'd201343623;
      3397: inst = 32'd203484854;
      3398: inst = 32'd471859200;
      3399: inst = 32'd136314880;
      3400: inst = 32'd268468224;
      3401: inst = 32'd201343624;
      3402: inst = 32'd203484854;
      3403: inst = 32'd471859200;
      3404: inst = 32'd136314880;
      3405: inst = 32'd268468224;
      3406: inst = 32'd201343625;
      3407: inst = 32'd203484854;
      3408: inst = 32'd471859200;
      3409: inst = 32'd136314880;
      3410: inst = 32'd268468224;
      3411: inst = 32'd201343626;
      3412: inst = 32'd203484854;
      3413: inst = 32'd471859200;
      3414: inst = 32'd136314880;
      3415: inst = 32'd268468224;
      3416: inst = 32'd201343627;
      3417: inst = 32'd203461810;
      3418: inst = 32'd471859200;
      3419: inst = 32'd136314880;
      3420: inst = 32'd268468224;
      3421: inst = 32'd201343628;
      3422: inst = 32'd203484854;
      3423: inst = 32'd471859200;
      3424: inst = 32'd136314880;
      3425: inst = 32'd268468224;
      3426: inst = 32'd201343629;
      3427: inst = 32'd203484854;
      3428: inst = 32'd471859200;
      3429: inst = 32'd136314880;
      3430: inst = 32'd268468224;
      3431: inst = 32'd201343630;
      3432: inst = 32'd203484854;
      3433: inst = 32'd471859200;
      3434: inst = 32'd136314880;
      3435: inst = 32'd268468224;
      3436: inst = 32'd201343631;
      3437: inst = 32'd203484854;
      3438: inst = 32'd471859200;
      3439: inst = 32'd136314880;
      3440: inst = 32'd268468224;
      3441: inst = 32'd201343632;
      3442: inst = 32'd203484854;
      3443: inst = 32'd471859200;
      3444: inst = 32'd136314880;
      3445: inst = 32'd268468224;
      3446: inst = 32'd201343633;
      3447: inst = 32'd203484854;
      3448: inst = 32'd471859200;
      3449: inst = 32'd136314880;
      3450: inst = 32'd268468224;
      3451: inst = 32'd201343634;
      3452: inst = 32'd203484854;
      3453: inst = 32'd471859200;
      3454: inst = 32'd136314880;
      3455: inst = 32'd268468224;
      3456: inst = 32'd201343635;
      3457: inst = 32'd203484854;
      3458: inst = 32'd471859200;
      3459: inst = 32'd136314880;
      3460: inst = 32'd268468224;
      3461: inst = 32'd201343636;
      3462: inst = 32'd203484854;
      3463: inst = 32'd471859200;
      3464: inst = 32'd136314880;
      3465: inst = 32'd268468224;
      3466: inst = 32'd201343637;
      3467: inst = 32'd203484854;
      3468: inst = 32'd471859200;
      3469: inst = 32'd136314880;
      3470: inst = 32'd268468224;
      3471: inst = 32'd201343638;
      3472: inst = 32'd203484854;
      3473: inst = 32'd471859200;
      3474: inst = 32'd136314880;
      3475: inst = 32'd268468224;
      3476: inst = 32'd201343639;
      3477: inst = 32'd203484854;
      3478: inst = 32'd471859200;
      3479: inst = 32'd136314880;
      3480: inst = 32'd268468224;
      3481: inst = 32'd201343640;
      3482: inst = 32'd203484854;
      3483: inst = 32'd471859200;
      3484: inst = 32'd136314880;
      3485: inst = 32'd268468224;
      3486: inst = 32'd201343641;
      3487: inst = 32'd203484854;
      3488: inst = 32'd471859200;
      3489: inst = 32'd136314880;
      3490: inst = 32'd268468224;
      3491: inst = 32'd201343642;
      3492: inst = 32'd203484854;
      3493: inst = 32'd471859200;
      3494: inst = 32'd136314880;
      3495: inst = 32'd268468224;
      3496: inst = 32'd201343643;
      3497: inst = 32'd203484854;
      3498: inst = 32'd471859200;
      3499: inst = 32'd136314880;
      3500: inst = 32'd268468224;
      3501: inst = 32'd201343644;
      3502: inst = 32'd203489279;
      3503: inst = 32'd471859200;
      3504: inst = 32'd136314880;
      3505: inst = 32'd268468224;
      3506: inst = 32'd201343645;
      3507: inst = 32'd203489279;
      3508: inst = 32'd471859200;
      3509: inst = 32'd136314880;
      3510: inst = 32'd268468224;
      3511: inst = 32'd201343646;
      3512: inst = 32'd203489279;
      3513: inst = 32'd471859200;
      3514: inst = 32'd136314880;
      3515: inst = 32'd268468224;
      3516: inst = 32'd201343647;
      3517: inst = 32'd203489279;
      3518: inst = 32'd471859200;
      3519: inst = 32'd136314880;
      3520: inst = 32'd268468224;
      3521: inst = 32'd201343648;
      3522: inst = 32'd203489279;
      3523: inst = 32'd471859200;
      3524: inst = 32'd136314880;
      3525: inst = 32'd268468224;
      3526: inst = 32'd201343649;
      3527: inst = 32'd203489279;
      3528: inst = 32'd471859200;
      3529: inst = 32'd136314880;
      3530: inst = 32'd268468224;
      3531: inst = 32'd201343650;
      3532: inst = 32'd203489279;
      3533: inst = 32'd471859200;
      3534: inst = 32'd136314880;
      3535: inst = 32'd268468224;
      3536: inst = 32'd201343651;
      3537: inst = 32'd203489279;
      3538: inst = 32'd471859200;
      3539: inst = 32'd136314880;
      3540: inst = 32'd268468224;
      3541: inst = 32'd201343652;
      3542: inst = 32'd203489279;
      3543: inst = 32'd471859200;
      3544: inst = 32'd136314880;
      3545: inst = 32'd268468224;
      3546: inst = 32'd201343653;
      3547: inst = 32'd203489279;
      3548: inst = 32'd471859200;
      3549: inst = 32'd136314880;
      3550: inst = 32'd268468224;
      3551: inst = 32'd201343654;
      3552: inst = 32'd203489279;
      3553: inst = 32'd471859200;
      3554: inst = 32'd136314880;
      3555: inst = 32'd268468224;
      3556: inst = 32'd201343655;
      3557: inst = 32'd203489279;
      3558: inst = 32'd471859200;
      3559: inst = 32'd136314880;
      3560: inst = 32'd268468224;
      3561: inst = 32'd201343656;
      3562: inst = 32'd203489279;
      3563: inst = 32'd471859200;
      3564: inst = 32'd136314880;
      3565: inst = 32'd268468224;
      3566: inst = 32'd201343657;
      3567: inst = 32'd203489279;
      3568: inst = 32'd471859200;
      3569: inst = 32'd136314880;
      3570: inst = 32'd268468224;
      3571: inst = 32'd201343658;
      3572: inst = 32'd203489279;
      3573: inst = 32'd471859200;
      3574: inst = 32'd136314880;
      3575: inst = 32'd268468224;
      3576: inst = 32'd201343659;
      3577: inst = 32'd203489279;
      3578: inst = 32'd471859200;
      3579: inst = 32'd136314880;
      3580: inst = 32'd268468224;
      3581: inst = 32'd201343660;
      3582: inst = 32'd203489279;
      3583: inst = 32'd471859200;
      3584: inst = 32'd136314880;
      3585: inst = 32'd268468224;
      3586: inst = 32'd201343661;
      3587: inst = 32'd203489279;
      3588: inst = 32'd471859200;
      3589: inst = 32'd136314880;
      3590: inst = 32'd268468224;
      3591: inst = 32'd201343662;
      3592: inst = 32'd203489279;
      3593: inst = 32'd471859200;
      3594: inst = 32'd136314880;
      3595: inst = 32'd268468224;
      3596: inst = 32'd201343663;
      3597: inst = 32'd203489279;
      3598: inst = 32'd471859200;
      3599: inst = 32'd136314880;
      3600: inst = 32'd268468224;
      3601: inst = 32'd201343664;
      3602: inst = 32'd203489279;
      3603: inst = 32'd471859200;
      3604: inst = 32'd136314880;
      3605: inst = 32'd268468224;
      3606: inst = 32'd201343665;
      3607: inst = 32'd203489279;
      3608: inst = 32'd471859200;
      3609: inst = 32'd136314880;
      3610: inst = 32'd268468224;
      3611: inst = 32'd201343666;
      3612: inst = 32'd203489279;
      3613: inst = 32'd471859200;
      3614: inst = 32'd136314880;
      3615: inst = 32'd268468224;
      3616: inst = 32'd201343667;
      3617: inst = 32'd203489279;
      3618: inst = 32'd471859200;
      3619: inst = 32'd136314880;
      3620: inst = 32'd268468224;
      3621: inst = 32'd201343668;
      3622: inst = 32'd203489279;
      3623: inst = 32'd471859200;
      3624: inst = 32'd136314880;
      3625: inst = 32'd268468224;
      3626: inst = 32'd201343669;
      3627: inst = 32'd203489279;
      3628: inst = 32'd471859200;
      3629: inst = 32'd136314880;
      3630: inst = 32'd268468224;
      3631: inst = 32'd201343670;
      3632: inst = 32'd203489279;
      3633: inst = 32'd471859200;
      3634: inst = 32'd136314880;
      3635: inst = 32'd268468224;
      3636: inst = 32'd201343671;
      3637: inst = 32'd203489279;
      3638: inst = 32'd471859200;
      3639: inst = 32'd136314880;
      3640: inst = 32'd268468224;
      3641: inst = 32'd201343672;
      3642: inst = 32'd203489279;
      3643: inst = 32'd471859200;
      3644: inst = 32'd136314880;
      3645: inst = 32'd268468224;
      3646: inst = 32'd201343673;
      3647: inst = 32'd203489279;
      3648: inst = 32'd471859200;
      3649: inst = 32'd136314880;
      3650: inst = 32'd268468224;
      3651: inst = 32'd201343674;
      3652: inst = 32'd203489279;
      3653: inst = 32'd471859200;
      3654: inst = 32'd136314880;
      3655: inst = 32'd268468224;
      3656: inst = 32'd201343675;
      3657: inst = 32'd203489279;
      3658: inst = 32'd471859200;
      3659: inst = 32'd136314880;
      3660: inst = 32'd268468224;
      3661: inst = 32'd201343676;
      3662: inst = 32'd203489279;
      3663: inst = 32'd471859200;
      3664: inst = 32'd136314880;
      3665: inst = 32'd268468224;
      3666: inst = 32'd201343677;
      3667: inst = 32'd203489279;
      3668: inst = 32'd471859200;
      3669: inst = 32'd136314880;
      3670: inst = 32'd268468224;
      3671: inst = 32'd201343678;
      3672: inst = 32'd203489279;
      3673: inst = 32'd471859200;
      3674: inst = 32'd136314880;
      3675: inst = 32'd268468224;
      3676: inst = 32'd201343679;
      3677: inst = 32'd203489279;
      3678: inst = 32'd471859200;
      3679: inst = 32'd136314880;
      3680: inst = 32'd268468224;
      3681: inst = 32'd201343680;
      3682: inst = 32'd203489279;
      3683: inst = 32'd471859200;
      3684: inst = 32'd136314880;
      3685: inst = 32'd268468224;
      3686: inst = 32'd201343681;
      3687: inst = 32'd203489279;
      3688: inst = 32'd471859200;
      3689: inst = 32'd136314880;
      3690: inst = 32'd268468224;
      3691: inst = 32'd201343682;
      3692: inst = 32'd203489279;
      3693: inst = 32'd471859200;
      3694: inst = 32'd136314880;
      3695: inst = 32'd268468224;
      3696: inst = 32'd201343683;
      3697: inst = 32'd203489279;
      3698: inst = 32'd471859200;
      3699: inst = 32'd136314880;
      3700: inst = 32'd268468224;
      3701: inst = 32'd201343684;
      3702: inst = 32'd203484854;
      3703: inst = 32'd471859200;
      3704: inst = 32'd136314880;
      3705: inst = 32'd268468224;
      3706: inst = 32'd201343685;
      3707: inst = 32'd203484854;
      3708: inst = 32'd471859200;
      3709: inst = 32'd136314880;
      3710: inst = 32'd268468224;
      3711: inst = 32'd201343686;
      3712: inst = 32'd203484854;
      3713: inst = 32'd471859200;
      3714: inst = 32'd136314880;
      3715: inst = 32'd268468224;
      3716: inst = 32'd201343687;
      3717: inst = 32'd203484854;
      3718: inst = 32'd471859200;
      3719: inst = 32'd136314880;
      3720: inst = 32'd268468224;
      3721: inst = 32'd201343688;
      3722: inst = 32'd203484854;
      3723: inst = 32'd471859200;
      3724: inst = 32'd136314880;
      3725: inst = 32'd268468224;
      3726: inst = 32'd201343689;
      3727: inst = 32'd203484854;
      3728: inst = 32'd471859200;
      3729: inst = 32'd136314880;
      3730: inst = 32'd268468224;
      3731: inst = 32'd201343690;
      3732: inst = 32'd203484854;
      3733: inst = 32'd471859200;
      3734: inst = 32'd136314880;
      3735: inst = 32'd268468224;
      3736: inst = 32'd201343691;
      3737: inst = 32'd203484854;
      3738: inst = 32'd471859200;
      3739: inst = 32'd136314880;
      3740: inst = 32'd268468224;
      3741: inst = 32'd201343692;
      3742: inst = 32'd203484854;
      3743: inst = 32'd471859200;
      3744: inst = 32'd136314880;
      3745: inst = 32'd268468224;
      3746: inst = 32'd201343693;
      3747: inst = 32'd203484854;
      3748: inst = 32'd471859200;
      3749: inst = 32'd136314880;
      3750: inst = 32'd268468224;
      3751: inst = 32'd201343694;
      3752: inst = 32'd203484854;
      3753: inst = 32'd471859200;
      3754: inst = 32'd136314880;
      3755: inst = 32'd268468224;
      3756: inst = 32'd201343695;
      3757: inst = 32'd203484854;
      3758: inst = 32'd471859200;
      3759: inst = 32'd136314880;
      3760: inst = 32'd268468224;
      3761: inst = 32'd201343696;
      3762: inst = 32'd203484854;
      3763: inst = 32'd471859200;
      3764: inst = 32'd136314880;
      3765: inst = 32'd268468224;
      3766: inst = 32'd201343697;
      3767: inst = 32'd203484854;
      3768: inst = 32'd471859200;
      3769: inst = 32'd136314880;
      3770: inst = 32'd268468224;
      3771: inst = 32'd201343698;
      3772: inst = 32'd203484854;
      3773: inst = 32'd471859200;
      3774: inst = 32'd136314880;
      3775: inst = 32'd268468224;
      3776: inst = 32'd201343699;
      3777: inst = 32'd203484854;
      3778: inst = 32'd471859200;
      3779: inst = 32'd136314880;
      3780: inst = 32'd268468224;
      3781: inst = 32'd201343700;
      3782: inst = 32'd203484854;
      3783: inst = 32'd471859200;
      3784: inst = 32'd136314880;
      3785: inst = 32'd268468224;
      3786: inst = 32'd201343701;
      3787: inst = 32'd203484854;
      3788: inst = 32'd471859200;
      3789: inst = 32'd136314880;
      3790: inst = 32'd268468224;
      3791: inst = 32'd201343702;
      3792: inst = 32'd203484854;
      3793: inst = 32'd471859200;
      3794: inst = 32'd136314880;
      3795: inst = 32'd268468224;
      3796: inst = 32'd201343703;
      3797: inst = 32'd203484854;
      3798: inst = 32'd471859200;
      3799: inst = 32'd136314880;
      3800: inst = 32'd268468224;
      3801: inst = 32'd201343704;
      3802: inst = 32'd203484854;
      3803: inst = 32'd471859200;
      3804: inst = 32'd136314880;
      3805: inst = 32'd268468224;
      3806: inst = 32'd201343705;
      3807: inst = 32'd203484854;
      3808: inst = 32'd471859200;
      3809: inst = 32'd136314880;
      3810: inst = 32'd268468224;
      3811: inst = 32'd201343706;
      3812: inst = 32'd203484854;
      3813: inst = 32'd471859200;
      3814: inst = 32'd136314880;
      3815: inst = 32'd268468224;
      3816: inst = 32'd201343707;
      3817: inst = 32'd203484854;
      3818: inst = 32'd471859200;
      3819: inst = 32'd136314880;
      3820: inst = 32'd268468224;
      3821: inst = 32'd201343708;
      3822: inst = 32'd203484854;
      3823: inst = 32'd471859200;
      3824: inst = 32'd136314880;
      3825: inst = 32'd268468224;
      3826: inst = 32'd201343709;
      3827: inst = 32'd203484854;
      3828: inst = 32'd471859200;
      3829: inst = 32'd136314880;
      3830: inst = 32'd268468224;
      3831: inst = 32'd201343710;
      3832: inst = 32'd203484854;
      3833: inst = 32'd471859200;
      3834: inst = 32'd136314880;
      3835: inst = 32'd268468224;
      3836: inst = 32'd201343711;
      3837: inst = 32'd203484854;
      3838: inst = 32'd471859200;
      3839: inst = 32'd136314880;
      3840: inst = 32'd268468224;
      3841: inst = 32'd201343712;
      3842: inst = 32'd203484854;
      3843: inst = 32'd471859200;
      3844: inst = 32'd136314880;
      3845: inst = 32'd268468224;
      3846: inst = 32'd201343713;
      3847: inst = 32'd203484854;
      3848: inst = 32'd471859200;
      3849: inst = 32'd136314880;
      3850: inst = 32'd268468224;
      3851: inst = 32'd201343714;
      3852: inst = 32'd203484854;
      3853: inst = 32'd471859200;
      3854: inst = 32'd136314880;
      3855: inst = 32'd268468224;
      3856: inst = 32'd201343715;
      3857: inst = 32'd203484854;
      3858: inst = 32'd471859200;
      3859: inst = 32'd136314880;
      3860: inst = 32'd268468224;
      3861: inst = 32'd201343716;
      3862: inst = 32'd203484854;
      3863: inst = 32'd471859200;
      3864: inst = 32'd136314880;
      3865: inst = 32'd268468224;
      3866: inst = 32'd201343717;
      3867: inst = 32'd203484854;
      3868: inst = 32'd471859200;
      3869: inst = 32'd136314880;
      3870: inst = 32'd268468224;
      3871: inst = 32'd201343718;
      3872: inst = 32'd203484854;
      3873: inst = 32'd471859200;
      3874: inst = 32'd136314880;
      3875: inst = 32'd268468224;
      3876: inst = 32'd201343719;
      3877: inst = 32'd203484854;
      3878: inst = 32'd471859200;
      3879: inst = 32'd136314880;
      3880: inst = 32'd268468224;
      3881: inst = 32'd201343720;
      3882: inst = 32'd203484854;
      3883: inst = 32'd471859200;
      3884: inst = 32'd136314880;
      3885: inst = 32'd268468224;
      3886: inst = 32'd201343721;
      3887: inst = 32'd203484854;
      3888: inst = 32'd471859200;
      3889: inst = 32'd136314880;
      3890: inst = 32'd268468224;
      3891: inst = 32'd201343722;
      3892: inst = 32'd203484789;
      3893: inst = 32'd471859200;
      3894: inst = 32'd136314880;
      3895: inst = 32'd268468224;
      3896: inst = 32'd201343723;
      3897: inst = 32'd203478060;
      3898: inst = 32'd471859200;
      3899: inst = 32'd136314880;
      3900: inst = 32'd268468224;
      3901: inst = 32'd201343724;
      3902: inst = 32'd203478060;
      3903: inst = 32'd471859200;
      3904: inst = 32'd136314880;
      3905: inst = 32'd268468224;
      3906: inst = 32'd201343725;
      3907: inst = 32'd203484757;
      3908: inst = 32'd471859200;
      3909: inst = 32'd136314880;
      3910: inst = 32'd268468224;
      3911: inst = 32'd201343726;
      3912: inst = 32'd203484854;
      3913: inst = 32'd471859200;
      3914: inst = 32'd136314880;
      3915: inst = 32'd268468224;
      3916: inst = 32'd201343727;
      3917: inst = 32'd203484854;
      3918: inst = 32'd471859200;
      3919: inst = 32'd136314880;
      3920: inst = 32'd268468224;
      3921: inst = 32'd201343728;
      3922: inst = 32'd203484854;
      3923: inst = 32'd471859200;
      3924: inst = 32'd136314880;
      3925: inst = 32'd268468224;
      3926: inst = 32'd201343729;
      3927: inst = 32'd203484854;
      3928: inst = 32'd471859200;
      3929: inst = 32'd136314880;
      3930: inst = 32'd268468224;
      3931: inst = 32'd201343730;
      3932: inst = 32'd203484854;
      3933: inst = 32'd471859200;
      3934: inst = 32'd136314880;
      3935: inst = 32'd268468224;
      3936: inst = 32'd201343731;
      3937: inst = 32'd203484854;
      3938: inst = 32'd471859200;
      3939: inst = 32'd136314880;
      3940: inst = 32'd268468224;
      3941: inst = 32'd201343732;
      3942: inst = 32'd203484854;
      3943: inst = 32'd471859200;
      3944: inst = 32'd136314880;
      3945: inst = 32'd268468224;
      3946: inst = 32'd201343733;
      3947: inst = 32'd203484854;
      3948: inst = 32'd471859200;
      3949: inst = 32'd136314880;
      3950: inst = 32'd268468224;
      3951: inst = 32'd201343734;
      3952: inst = 32'd203484854;
      3953: inst = 32'd471859200;
      3954: inst = 32'd136314880;
      3955: inst = 32'd268468224;
      3956: inst = 32'd201343735;
      3957: inst = 32'd203484854;
      3958: inst = 32'd471859200;
      3959: inst = 32'd136314880;
      3960: inst = 32'd268468224;
      3961: inst = 32'd201343736;
      3962: inst = 32'd203484854;
      3963: inst = 32'd471859200;
      3964: inst = 32'd136314880;
      3965: inst = 32'd268468224;
      3966: inst = 32'd201343737;
      3967: inst = 32'd203484854;
      3968: inst = 32'd471859200;
      3969: inst = 32'd136314880;
      3970: inst = 32'd268468224;
      3971: inst = 32'd201343738;
      3972: inst = 32'd203484854;
      3973: inst = 32'd471859200;
      3974: inst = 32'd136314880;
      3975: inst = 32'd268468224;
      3976: inst = 32'd201343739;
      3977: inst = 32'd203484854;
      3978: inst = 32'd471859200;
      3979: inst = 32'd136314880;
      3980: inst = 32'd268468224;
      3981: inst = 32'd201343740;
      3982: inst = 32'd203489279;
      3983: inst = 32'd471859200;
      3984: inst = 32'd136314880;
      3985: inst = 32'd268468224;
      3986: inst = 32'd201343741;
      3987: inst = 32'd203489279;
      3988: inst = 32'd471859200;
      3989: inst = 32'd136314880;
      3990: inst = 32'd268468224;
      3991: inst = 32'd201343742;
      3992: inst = 32'd203489279;
      3993: inst = 32'd471859200;
      3994: inst = 32'd136314880;
      3995: inst = 32'd268468224;
      3996: inst = 32'd201343743;
      3997: inst = 32'd203489279;
      3998: inst = 32'd471859200;
      3999: inst = 32'd136314880;
      4000: inst = 32'd268468224;
      4001: inst = 32'd201343744;
      4002: inst = 32'd203489279;
      4003: inst = 32'd471859200;
      4004: inst = 32'd136314880;
      4005: inst = 32'd268468224;
      4006: inst = 32'd201343745;
      4007: inst = 32'd203489279;
      4008: inst = 32'd471859200;
      4009: inst = 32'd136314880;
      4010: inst = 32'd268468224;
      4011: inst = 32'd201343746;
      4012: inst = 32'd203489279;
      4013: inst = 32'd471859200;
      4014: inst = 32'd136314880;
      4015: inst = 32'd268468224;
      4016: inst = 32'd201343747;
      4017: inst = 32'd203489279;
      4018: inst = 32'd471859200;
      4019: inst = 32'd136314880;
      4020: inst = 32'd268468224;
      4021: inst = 32'd201343748;
      4022: inst = 32'd203489279;
      4023: inst = 32'd471859200;
      4024: inst = 32'd136314880;
      4025: inst = 32'd268468224;
      4026: inst = 32'd201343749;
      4027: inst = 32'd203489279;
      4028: inst = 32'd471859200;
      4029: inst = 32'd136314880;
      4030: inst = 32'd268468224;
      4031: inst = 32'd201343750;
      4032: inst = 32'd203489279;
      4033: inst = 32'd471859200;
      4034: inst = 32'd136314880;
      4035: inst = 32'd268468224;
      4036: inst = 32'd201343751;
      4037: inst = 32'd203489279;
      4038: inst = 32'd471859200;
      4039: inst = 32'd136314880;
      4040: inst = 32'd268468224;
      4041: inst = 32'd201343752;
      4042: inst = 32'd203489279;
      4043: inst = 32'd471859200;
      4044: inst = 32'd136314880;
      4045: inst = 32'd268468224;
      4046: inst = 32'd201343753;
      4047: inst = 32'd203489279;
      4048: inst = 32'd471859200;
      4049: inst = 32'd136314880;
      4050: inst = 32'd268468224;
      4051: inst = 32'd201343754;
      4052: inst = 32'd203489279;
      4053: inst = 32'd471859200;
      4054: inst = 32'd136314880;
      4055: inst = 32'd268468224;
      4056: inst = 32'd201343755;
      4057: inst = 32'd203489279;
      4058: inst = 32'd471859200;
      4059: inst = 32'd136314880;
      4060: inst = 32'd268468224;
      4061: inst = 32'd201343756;
      4062: inst = 32'd203489279;
      4063: inst = 32'd471859200;
      4064: inst = 32'd136314880;
      4065: inst = 32'd268468224;
      4066: inst = 32'd201343757;
      4067: inst = 32'd203489279;
      4068: inst = 32'd471859200;
      4069: inst = 32'd136314880;
      4070: inst = 32'd268468224;
      4071: inst = 32'd201343758;
      4072: inst = 32'd203489279;
      4073: inst = 32'd471859200;
      4074: inst = 32'd136314880;
      4075: inst = 32'd268468224;
      4076: inst = 32'd201343759;
      4077: inst = 32'd203489279;
      4078: inst = 32'd471859200;
      4079: inst = 32'd136314880;
      4080: inst = 32'd268468224;
      4081: inst = 32'd201343760;
      4082: inst = 32'd203489279;
      4083: inst = 32'd471859200;
      4084: inst = 32'd136314880;
      4085: inst = 32'd268468224;
      4086: inst = 32'd201343761;
      4087: inst = 32'd203489279;
      4088: inst = 32'd471859200;
      4089: inst = 32'd136314880;
      4090: inst = 32'd268468224;
      4091: inst = 32'd201343762;
      4092: inst = 32'd203489279;
      4093: inst = 32'd471859200;
      4094: inst = 32'd136314880;
      4095: inst = 32'd268468224;
      4096: inst = 32'd201343763;
      4097: inst = 32'd203489279;
      4098: inst = 32'd471859200;
      4099: inst = 32'd136314880;
      4100: inst = 32'd268468224;
      4101: inst = 32'd201343764;
      4102: inst = 32'd203489279;
      4103: inst = 32'd471859200;
      4104: inst = 32'd136314880;
      4105: inst = 32'd268468224;
      4106: inst = 32'd201343765;
      4107: inst = 32'd203489279;
      4108: inst = 32'd471859200;
      4109: inst = 32'd136314880;
      4110: inst = 32'd268468224;
      4111: inst = 32'd201343766;
      4112: inst = 32'd203489279;
      4113: inst = 32'd471859200;
      4114: inst = 32'd136314880;
      4115: inst = 32'd268468224;
      4116: inst = 32'd201343767;
      4117: inst = 32'd203489279;
      4118: inst = 32'd471859200;
      4119: inst = 32'd136314880;
      4120: inst = 32'd268468224;
      4121: inst = 32'd201343768;
      4122: inst = 32'd203489279;
      4123: inst = 32'd471859200;
      4124: inst = 32'd136314880;
      4125: inst = 32'd268468224;
      4126: inst = 32'd201343769;
      4127: inst = 32'd203489279;
      4128: inst = 32'd471859200;
      4129: inst = 32'd136314880;
      4130: inst = 32'd268468224;
      4131: inst = 32'd201343770;
      4132: inst = 32'd203489279;
      4133: inst = 32'd471859200;
      4134: inst = 32'd136314880;
      4135: inst = 32'd268468224;
      4136: inst = 32'd201343771;
      4137: inst = 32'd203489279;
      4138: inst = 32'd471859200;
      4139: inst = 32'd136314880;
      4140: inst = 32'd268468224;
      4141: inst = 32'd201343772;
      4142: inst = 32'd203489279;
      4143: inst = 32'd471859200;
      4144: inst = 32'd136314880;
      4145: inst = 32'd268468224;
      4146: inst = 32'd201343773;
      4147: inst = 32'd203489279;
      4148: inst = 32'd471859200;
      4149: inst = 32'd136314880;
      4150: inst = 32'd268468224;
      4151: inst = 32'd201343774;
      4152: inst = 32'd203489279;
      4153: inst = 32'd471859200;
      4154: inst = 32'd136314880;
      4155: inst = 32'd268468224;
      4156: inst = 32'd201343775;
      4157: inst = 32'd203489279;
      4158: inst = 32'd471859200;
      4159: inst = 32'd136314880;
      4160: inst = 32'd268468224;
      4161: inst = 32'd201343776;
      4162: inst = 32'd203489279;
      4163: inst = 32'd471859200;
      4164: inst = 32'd136314880;
      4165: inst = 32'd268468224;
      4166: inst = 32'd201343777;
      4167: inst = 32'd203489279;
      4168: inst = 32'd471859200;
      4169: inst = 32'd136314880;
      4170: inst = 32'd268468224;
      4171: inst = 32'd201343778;
      4172: inst = 32'd203489279;
      4173: inst = 32'd471859200;
      4174: inst = 32'd136314880;
      4175: inst = 32'd268468224;
      4176: inst = 32'd201343779;
      4177: inst = 32'd203489279;
      4178: inst = 32'd471859200;
      4179: inst = 32'd136314880;
      4180: inst = 32'd268468224;
      4181: inst = 32'd201343780;
      4182: inst = 32'd203484854;
      4183: inst = 32'd471859200;
      4184: inst = 32'd136314880;
      4185: inst = 32'd268468224;
      4186: inst = 32'd201343781;
      4187: inst = 32'd203484854;
      4188: inst = 32'd471859200;
      4189: inst = 32'd136314880;
      4190: inst = 32'd268468224;
      4191: inst = 32'd201343782;
      4192: inst = 32'd203484854;
      4193: inst = 32'd471859200;
      4194: inst = 32'd136314880;
      4195: inst = 32'd268468224;
      4196: inst = 32'd201343783;
      4197: inst = 32'd203484854;
      4198: inst = 32'd471859200;
      4199: inst = 32'd136314880;
      4200: inst = 32'd268468224;
      4201: inst = 32'd201343784;
      4202: inst = 32'd203484854;
      4203: inst = 32'd471859200;
      4204: inst = 32'd136314880;
      4205: inst = 32'd268468224;
      4206: inst = 32'd201343785;
      4207: inst = 32'd203484854;
      4208: inst = 32'd471859200;
      4209: inst = 32'd136314880;
      4210: inst = 32'd268468224;
      4211: inst = 32'd201343786;
      4212: inst = 32'd203484854;
      4213: inst = 32'd471859200;
      4214: inst = 32'd136314880;
      4215: inst = 32'd268468224;
      4216: inst = 32'd201343787;
      4217: inst = 32'd203484854;
      4218: inst = 32'd471859200;
      4219: inst = 32'd136314880;
      4220: inst = 32'd268468224;
      4221: inst = 32'd201343788;
      4222: inst = 32'd203484854;
      4223: inst = 32'd471859200;
      4224: inst = 32'd136314880;
      4225: inst = 32'd268468224;
      4226: inst = 32'd201343789;
      4227: inst = 32'd203484854;
      4228: inst = 32'd471859200;
      4229: inst = 32'd136314880;
      4230: inst = 32'd268468224;
      4231: inst = 32'd201343790;
      4232: inst = 32'd203484854;
      4233: inst = 32'd471859200;
      4234: inst = 32'd136314880;
      4235: inst = 32'd268468224;
      4236: inst = 32'd201343791;
      4237: inst = 32'd203484854;
      4238: inst = 32'd471859200;
      4239: inst = 32'd136314880;
      4240: inst = 32'd268468224;
      4241: inst = 32'd201343792;
      4242: inst = 32'd203484854;
      4243: inst = 32'd471859200;
      4244: inst = 32'd136314880;
      4245: inst = 32'd268468224;
      4246: inst = 32'd201343793;
      4247: inst = 32'd203484854;
      4248: inst = 32'd471859200;
      4249: inst = 32'd136314880;
      4250: inst = 32'd268468224;
      4251: inst = 32'd201343794;
      4252: inst = 32'd203484854;
      4253: inst = 32'd471859200;
      4254: inst = 32'd136314880;
      4255: inst = 32'd268468224;
      4256: inst = 32'd201343795;
      4257: inst = 32'd203484854;
      4258: inst = 32'd471859200;
      4259: inst = 32'd136314880;
      4260: inst = 32'd268468224;
      4261: inst = 32'd201343796;
      4262: inst = 32'd203484854;
      4263: inst = 32'd471859200;
      4264: inst = 32'd136314880;
      4265: inst = 32'd268468224;
      4266: inst = 32'd201343797;
      4267: inst = 32'd203484854;
      4268: inst = 32'd471859200;
      4269: inst = 32'd136314880;
      4270: inst = 32'd268468224;
      4271: inst = 32'd201343798;
      4272: inst = 32'd203484854;
      4273: inst = 32'd471859200;
      4274: inst = 32'd136314880;
      4275: inst = 32'd268468224;
      4276: inst = 32'd201343799;
      4277: inst = 32'd203484854;
      4278: inst = 32'd471859200;
      4279: inst = 32'd136314880;
      4280: inst = 32'd268468224;
      4281: inst = 32'd201343800;
      4282: inst = 32'd203484854;
      4283: inst = 32'd471859200;
      4284: inst = 32'd136314880;
      4285: inst = 32'd268468224;
      4286: inst = 32'd201343801;
      4287: inst = 32'd203484854;
      4288: inst = 32'd471859200;
      4289: inst = 32'd136314880;
      4290: inst = 32'd268468224;
      4291: inst = 32'd201343802;
      4292: inst = 32'd203484854;
      4293: inst = 32'd471859200;
      4294: inst = 32'd136314880;
      4295: inst = 32'd268468224;
      4296: inst = 32'd201343803;
      4297: inst = 32'd203484854;
      4298: inst = 32'd471859200;
      4299: inst = 32'd136314880;
      4300: inst = 32'd268468224;
      4301: inst = 32'd201343804;
      4302: inst = 32'd203484854;
      4303: inst = 32'd471859200;
      4304: inst = 32'd136314880;
      4305: inst = 32'd268468224;
      4306: inst = 32'd201343805;
      4307: inst = 32'd203484854;
      4308: inst = 32'd471859200;
      4309: inst = 32'd136314880;
      4310: inst = 32'd268468224;
      4311: inst = 32'd201343806;
      4312: inst = 32'd203484854;
      4313: inst = 32'd471859200;
      4314: inst = 32'd136314880;
      4315: inst = 32'd268468224;
      4316: inst = 32'd201343807;
      4317: inst = 32'd203484854;
      4318: inst = 32'd471859200;
      4319: inst = 32'd136314880;
      4320: inst = 32'd268468224;
      4321: inst = 32'd201343808;
      4322: inst = 32'd203484854;
      4323: inst = 32'd471859200;
      4324: inst = 32'd136314880;
      4325: inst = 32'd268468224;
      4326: inst = 32'd201343809;
      4327: inst = 32'd203484854;
      4328: inst = 32'd471859200;
      4329: inst = 32'd136314880;
      4330: inst = 32'd268468224;
      4331: inst = 32'd201343810;
      4332: inst = 32'd203484854;
      4333: inst = 32'd471859200;
      4334: inst = 32'd136314880;
      4335: inst = 32'd268468224;
      4336: inst = 32'd201343811;
      4337: inst = 32'd203484854;
      4338: inst = 32'd471859200;
      4339: inst = 32'd136314880;
      4340: inst = 32'd268468224;
      4341: inst = 32'd201343812;
      4342: inst = 32'd203484854;
      4343: inst = 32'd471859200;
      4344: inst = 32'd136314880;
      4345: inst = 32'd268468224;
      4346: inst = 32'd201343813;
      4347: inst = 32'd203484854;
      4348: inst = 32'd471859200;
      4349: inst = 32'd136314880;
      4350: inst = 32'd268468224;
      4351: inst = 32'd201343814;
      4352: inst = 32'd203484854;
      4353: inst = 32'd471859200;
      4354: inst = 32'd136314880;
      4355: inst = 32'd268468224;
      4356: inst = 32'd201343815;
      4357: inst = 32'd203484854;
      4358: inst = 32'd471859200;
      4359: inst = 32'd136314880;
      4360: inst = 32'd268468224;
      4361: inst = 32'd201343816;
      4362: inst = 32'd203484854;
      4363: inst = 32'd471859200;
      4364: inst = 32'd136314880;
      4365: inst = 32'd268468224;
      4366: inst = 32'd201343817;
      4367: inst = 32'd203482481;
      4368: inst = 32'd471859200;
      4369: inst = 32'd136314880;
      4370: inst = 32'd268468224;
      4371: inst = 32'd201343818;
      4372: inst = 32'd203475752;
      4373: inst = 32'd471859200;
      4374: inst = 32'd136314880;
      4375: inst = 32'd268468224;
      4376: inst = 32'd201343819;
      4377: inst = 32'd203475655;
      4378: inst = 32'd471859200;
      4379: inst = 32'd136314880;
      4380: inst = 32'd268468224;
      4381: inst = 32'd201343820;
      4382: inst = 32'd203475655;
      4383: inst = 32'd471859200;
      4384: inst = 32'd136314880;
      4385: inst = 32'd268468224;
      4386: inst = 32'd201343821;
      4387: inst = 32'd203475752;
      4388: inst = 32'd471859200;
      4389: inst = 32'd136314880;
      4390: inst = 32'd268468224;
      4391: inst = 32'd201343822;
      4392: inst = 32'd203482481;
      4393: inst = 32'd471859200;
      4394: inst = 32'd136314880;
      4395: inst = 32'd268468224;
      4396: inst = 32'd201343823;
      4397: inst = 32'd203484854;
      4398: inst = 32'd471859200;
      4399: inst = 32'd136314880;
      4400: inst = 32'd268468224;
      4401: inst = 32'd201343824;
      4402: inst = 32'd203484854;
      4403: inst = 32'd471859200;
      4404: inst = 32'd136314880;
      4405: inst = 32'd268468224;
      4406: inst = 32'd201343825;
      4407: inst = 32'd203484854;
      4408: inst = 32'd471859200;
      4409: inst = 32'd136314880;
      4410: inst = 32'd268468224;
      4411: inst = 32'd201343826;
      4412: inst = 32'd203484854;
      4413: inst = 32'd471859200;
      4414: inst = 32'd136314880;
      4415: inst = 32'd268468224;
      4416: inst = 32'd201343827;
      4417: inst = 32'd203484854;
      4418: inst = 32'd471859200;
      4419: inst = 32'd136314880;
      4420: inst = 32'd268468224;
      4421: inst = 32'd201343828;
      4422: inst = 32'd203484854;
      4423: inst = 32'd471859200;
      4424: inst = 32'd136314880;
      4425: inst = 32'd268468224;
      4426: inst = 32'd201343829;
      4427: inst = 32'd203484854;
      4428: inst = 32'd471859200;
      4429: inst = 32'd136314880;
      4430: inst = 32'd268468224;
      4431: inst = 32'd201343830;
      4432: inst = 32'd203484854;
      4433: inst = 32'd471859200;
      4434: inst = 32'd136314880;
      4435: inst = 32'd268468224;
      4436: inst = 32'd201343831;
      4437: inst = 32'd203484854;
      4438: inst = 32'd471859200;
      4439: inst = 32'd136314880;
      4440: inst = 32'd268468224;
      4441: inst = 32'd201343832;
      4442: inst = 32'd203484854;
      4443: inst = 32'd471859200;
      4444: inst = 32'd136314880;
      4445: inst = 32'd268468224;
      4446: inst = 32'd201343833;
      4447: inst = 32'd203484854;
      4448: inst = 32'd471859200;
      4449: inst = 32'd136314880;
      4450: inst = 32'd268468224;
      4451: inst = 32'd201343834;
      4452: inst = 32'd203484854;
      4453: inst = 32'd471859200;
      4454: inst = 32'd136314880;
      4455: inst = 32'd268468224;
      4456: inst = 32'd201343835;
      4457: inst = 32'd203484854;
      4458: inst = 32'd471859200;
      4459: inst = 32'd136314880;
      4460: inst = 32'd268468224;
      4461: inst = 32'd201343836;
      4462: inst = 32'd203489279;
      4463: inst = 32'd471859200;
      4464: inst = 32'd136314880;
      4465: inst = 32'd268468224;
      4466: inst = 32'd201343837;
      4467: inst = 32'd203489279;
      4468: inst = 32'd471859200;
      4469: inst = 32'd136314880;
      4470: inst = 32'd268468224;
      4471: inst = 32'd201343838;
      4472: inst = 32'd203489279;
      4473: inst = 32'd471859200;
      4474: inst = 32'd136314880;
      4475: inst = 32'd268468224;
      4476: inst = 32'd201343839;
      4477: inst = 32'd203489279;
      4478: inst = 32'd471859200;
      4479: inst = 32'd136314880;
      4480: inst = 32'd268468224;
      4481: inst = 32'd201343840;
      4482: inst = 32'd203489279;
      4483: inst = 32'd471859200;
      4484: inst = 32'd136314880;
      4485: inst = 32'd268468224;
      4486: inst = 32'd201343841;
      4487: inst = 32'd203489279;
      4488: inst = 32'd471859200;
      4489: inst = 32'd136314880;
      4490: inst = 32'd268468224;
      4491: inst = 32'd201343842;
      4492: inst = 32'd203489279;
      4493: inst = 32'd471859200;
      4494: inst = 32'd136314880;
      4495: inst = 32'd268468224;
      4496: inst = 32'd201343843;
      4497: inst = 32'd203489279;
      4498: inst = 32'd471859200;
      4499: inst = 32'd136314880;
      4500: inst = 32'd268468224;
      4501: inst = 32'd201343844;
      4502: inst = 32'd203489279;
      4503: inst = 32'd471859200;
      4504: inst = 32'd136314880;
      4505: inst = 32'd268468224;
      4506: inst = 32'd201343845;
      4507: inst = 32'd203489279;
      4508: inst = 32'd471859200;
      4509: inst = 32'd136314880;
      4510: inst = 32'd268468224;
      4511: inst = 32'd201343846;
      4512: inst = 32'd203489279;
      4513: inst = 32'd471859200;
      4514: inst = 32'd136314880;
      4515: inst = 32'd268468224;
      4516: inst = 32'd201343847;
      4517: inst = 32'd203489279;
      4518: inst = 32'd471859200;
      4519: inst = 32'd136314880;
      4520: inst = 32'd268468224;
      4521: inst = 32'd201343848;
      4522: inst = 32'd203489279;
      4523: inst = 32'd471859200;
      4524: inst = 32'd136314880;
      4525: inst = 32'd268468224;
      4526: inst = 32'd201343849;
      4527: inst = 32'd203489279;
      4528: inst = 32'd471859200;
      4529: inst = 32'd136314880;
      4530: inst = 32'd268468224;
      4531: inst = 32'd201343850;
      4532: inst = 32'd203489279;
      4533: inst = 32'd471859200;
      4534: inst = 32'd136314880;
      4535: inst = 32'd268468224;
      4536: inst = 32'd201343851;
      4537: inst = 32'd203489279;
      4538: inst = 32'd471859200;
      4539: inst = 32'd136314880;
      4540: inst = 32'd268468224;
      4541: inst = 32'd201343852;
      4542: inst = 32'd203489279;
      4543: inst = 32'd471859200;
      4544: inst = 32'd136314880;
      4545: inst = 32'd268468224;
      4546: inst = 32'd201343853;
      4547: inst = 32'd203489279;
      4548: inst = 32'd471859200;
      4549: inst = 32'd136314880;
      4550: inst = 32'd268468224;
      4551: inst = 32'd201343854;
      4552: inst = 32'd203489279;
      4553: inst = 32'd471859200;
      4554: inst = 32'd136314880;
      4555: inst = 32'd268468224;
      4556: inst = 32'd201343855;
      4557: inst = 32'd203489279;
      4558: inst = 32'd471859200;
      4559: inst = 32'd136314880;
      4560: inst = 32'd268468224;
      4561: inst = 32'd201343856;
      4562: inst = 32'd203489279;
      4563: inst = 32'd471859200;
      4564: inst = 32'd136314880;
      4565: inst = 32'd268468224;
      4566: inst = 32'd201343857;
      4567: inst = 32'd203489279;
      4568: inst = 32'd471859200;
      4569: inst = 32'd136314880;
      4570: inst = 32'd268468224;
      4571: inst = 32'd201343858;
      4572: inst = 32'd203489279;
      4573: inst = 32'd471859200;
      4574: inst = 32'd136314880;
      4575: inst = 32'd268468224;
      4576: inst = 32'd201343859;
      4577: inst = 32'd203489279;
      4578: inst = 32'd471859200;
      4579: inst = 32'd136314880;
      4580: inst = 32'd268468224;
      4581: inst = 32'd201343860;
      4582: inst = 32'd203489279;
      4583: inst = 32'd471859200;
      4584: inst = 32'd136314880;
      4585: inst = 32'd268468224;
      4586: inst = 32'd201343861;
      4587: inst = 32'd203489279;
      4588: inst = 32'd471859200;
      4589: inst = 32'd136314880;
      4590: inst = 32'd268468224;
      4591: inst = 32'd201343862;
      4592: inst = 32'd203489279;
      4593: inst = 32'd471859200;
      4594: inst = 32'd136314880;
      4595: inst = 32'd268468224;
      4596: inst = 32'd201343863;
      4597: inst = 32'd203489279;
      4598: inst = 32'd471859200;
      4599: inst = 32'd136314880;
      4600: inst = 32'd268468224;
      4601: inst = 32'd201343864;
      4602: inst = 32'd203489279;
      4603: inst = 32'd471859200;
      4604: inst = 32'd136314880;
      4605: inst = 32'd268468224;
      4606: inst = 32'd201343865;
      4607: inst = 32'd203489279;
      4608: inst = 32'd471859200;
      4609: inst = 32'd136314880;
      4610: inst = 32'd268468224;
      4611: inst = 32'd201343866;
      4612: inst = 32'd203489279;
      4613: inst = 32'd471859200;
      4614: inst = 32'd136314880;
      4615: inst = 32'd268468224;
      4616: inst = 32'd201343867;
      4617: inst = 32'd203489279;
      4618: inst = 32'd471859200;
      4619: inst = 32'd136314880;
      4620: inst = 32'd268468224;
      4621: inst = 32'd201343868;
      4622: inst = 32'd203489279;
      4623: inst = 32'd471859200;
      4624: inst = 32'd136314880;
      4625: inst = 32'd268468224;
      4626: inst = 32'd201343869;
      4627: inst = 32'd203489279;
      4628: inst = 32'd471859200;
      4629: inst = 32'd136314880;
      4630: inst = 32'd268468224;
      4631: inst = 32'd201343870;
      4632: inst = 32'd203489279;
      4633: inst = 32'd471859200;
      4634: inst = 32'd136314880;
      4635: inst = 32'd268468224;
      4636: inst = 32'd201343871;
      4637: inst = 32'd203489279;
      4638: inst = 32'd471859200;
      4639: inst = 32'd136314880;
      4640: inst = 32'd268468224;
      4641: inst = 32'd201343872;
      4642: inst = 32'd203489279;
      4643: inst = 32'd471859200;
      4644: inst = 32'd136314880;
      4645: inst = 32'd268468224;
      4646: inst = 32'd201343873;
      4647: inst = 32'd203489279;
      4648: inst = 32'd471859200;
      4649: inst = 32'd136314880;
      4650: inst = 32'd268468224;
      4651: inst = 32'd201343874;
      4652: inst = 32'd203489279;
      4653: inst = 32'd471859200;
      4654: inst = 32'd136314880;
      4655: inst = 32'd268468224;
      4656: inst = 32'd201343875;
      4657: inst = 32'd203489279;
      4658: inst = 32'd471859200;
      4659: inst = 32'd136314880;
      4660: inst = 32'd268468224;
      4661: inst = 32'd201343876;
      4662: inst = 32'd203484854;
      4663: inst = 32'd471859200;
      4664: inst = 32'd136314880;
      4665: inst = 32'd268468224;
      4666: inst = 32'd201343877;
      4667: inst = 32'd203484854;
      4668: inst = 32'd471859200;
      4669: inst = 32'd136314880;
      4670: inst = 32'd268468224;
      4671: inst = 32'd201343878;
      4672: inst = 32'd203484854;
      4673: inst = 32'd471859200;
      4674: inst = 32'd136314880;
      4675: inst = 32'd268468224;
      4676: inst = 32'd201343879;
      4677: inst = 32'd203484854;
      4678: inst = 32'd471859200;
      4679: inst = 32'd136314880;
      4680: inst = 32'd268468224;
      4681: inst = 32'd201343880;
      4682: inst = 32'd203484854;
      4683: inst = 32'd471859200;
      4684: inst = 32'd136314880;
      4685: inst = 32'd268468224;
      4686: inst = 32'd201343881;
      4687: inst = 32'd203484854;
      4688: inst = 32'd471859200;
      4689: inst = 32'd136314880;
      4690: inst = 32'd268468224;
      4691: inst = 32'd201343882;
      4692: inst = 32'd203484854;
      4693: inst = 32'd471859200;
      4694: inst = 32'd136314880;
      4695: inst = 32'd268468224;
      4696: inst = 32'd201343883;
      4697: inst = 32'd203484854;
      4698: inst = 32'd471859200;
      4699: inst = 32'd136314880;
      4700: inst = 32'd268468224;
      4701: inst = 32'd201343884;
      4702: inst = 32'd203484854;
      4703: inst = 32'd471859200;
      4704: inst = 32'd136314880;
      4705: inst = 32'd268468224;
      4706: inst = 32'd201343885;
      4707: inst = 32'd203484854;
      4708: inst = 32'd471859200;
      4709: inst = 32'd136314880;
      4710: inst = 32'd268468224;
      4711: inst = 32'd201343886;
      4712: inst = 32'd203484854;
      4713: inst = 32'd471859200;
      4714: inst = 32'd136314880;
      4715: inst = 32'd268468224;
      4716: inst = 32'd201343887;
      4717: inst = 32'd203484854;
      4718: inst = 32'd471859200;
      4719: inst = 32'd136314880;
      4720: inst = 32'd268468224;
      4721: inst = 32'd201343888;
      4722: inst = 32'd203484854;
      4723: inst = 32'd471859200;
      4724: inst = 32'd136314880;
      4725: inst = 32'd268468224;
      4726: inst = 32'd201343889;
      4727: inst = 32'd203484854;
      4728: inst = 32'd471859200;
      4729: inst = 32'd136314880;
      4730: inst = 32'd268468224;
      4731: inst = 32'd201343890;
      4732: inst = 32'd203484854;
      4733: inst = 32'd471859200;
      4734: inst = 32'd136314880;
      4735: inst = 32'd268468224;
      4736: inst = 32'd201343891;
      4737: inst = 32'd203484854;
      4738: inst = 32'd471859200;
      4739: inst = 32'd136314880;
      4740: inst = 32'd268468224;
      4741: inst = 32'd201343892;
      4742: inst = 32'd203484854;
      4743: inst = 32'd471859200;
      4744: inst = 32'd136314880;
      4745: inst = 32'd268468224;
      4746: inst = 32'd201343893;
      4747: inst = 32'd203484854;
      4748: inst = 32'd471859200;
      4749: inst = 32'd136314880;
      4750: inst = 32'd268468224;
      4751: inst = 32'd201343894;
      4752: inst = 32'd203484854;
      4753: inst = 32'd471859200;
      4754: inst = 32'd136314880;
      4755: inst = 32'd268468224;
      4756: inst = 32'd201343895;
      4757: inst = 32'd203484854;
      4758: inst = 32'd471859200;
      4759: inst = 32'd136314880;
      4760: inst = 32'd268468224;
      4761: inst = 32'd201343896;
      4762: inst = 32'd203484854;
      4763: inst = 32'd471859200;
      4764: inst = 32'd136314880;
      4765: inst = 32'd268468224;
      4766: inst = 32'd201343897;
      4767: inst = 32'd203484854;
      4768: inst = 32'd471859200;
      4769: inst = 32'd136314880;
      4770: inst = 32'd268468224;
      4771: inst = 32'd201343898;
      4772: inst = 32'd203484854;
      4773: inst = 32'd471859200;
      4774: inst = 32'd136314880;
      4775: inst = 32'd268468224;
      4776: inst = 32'd201343899;
      4777: inst = 32'd203484854;
      4778: inst = 32'd471859200;
      4779: inst = 32'd136314880;
      4780: inst = 32'd268468224;
      4781: inst = 32'd201343900;
      4782: inst = 32'd203484854;
      4783: inst = 32'd471859200;
      4784: inst = 32'd136314880;
      4785: inst = 32'd268468224;
      4786: inst = 32'd201343901;
      4787: inst = 32'd203484854;
      4788: inst = 32'd471859200;
      4789: inst = 32'd136314880;
      4790: inst = 32'd268468224;
      4791: inst = 32'd201343902;
      4792: inst = 32'd203484854;
      4793: inst = 32'd471859200;
      4794: inst = 32'd136314880;
      4795: inst = 32'd268468224;
      4796: inst = 32'd201343903;
      4797: inst = 32'd203484854;
      4798: inst = 32'd471859200;
      4799: inst = 32'd136314880;
      4800: inst = 32'd268468224;
      4801: inst = 32'd201343904;
      4802: inst = 32'd203484854;
      4803: inst = 32'd471859200;
      4804: inst = 32'd136314880;
      4805: inst = 32'd268468224;
      4806: inst = 32'd201343905;
      4807: inst = 32'd203484854;
      4808: inst = 32'd471859200;
      4809: inst = 32'd136314880;
      4810: inst = 32'd268468224;
      4811: inst = 32'd201343906;
      4812: inst = 32'd203484854;
      4813: inst = 32'd471859200;
      4814: inst = 32'd136314880;
      4815: inst = 32'd268468224;
      4816: inst = 32'd201343907;
      4817: inst = 32'd203484854;
      4818: inst = 32'd471859200;
      4819: inst = 32'd136314880;
      4820: inst = 32'd268468224;
      4821: inst = 32'd201343908;
      4822: inst = 32'd203484854;
      4823: inst = 32'd471859200;
      4824: inst = 32'd136314880;
      4825: inst = 32'd268468224;
      4826: inst = 32'd201343909;
      4827: inst = 32'd203484854;
      4828: inst = 32'd471859200;
      4829: inst = 32'd136314880;
      4830: inst = 32'd268468224;
      4831: inst = 32'd201343910;
      4832: inst = 32'd203484854;
      4833: inst = 32'd471859200;
      4834: inst = 32'd136314880;
      4835: inst = 32'd268468224;
      4836: inst = 32'd201343911;
      4837: inst = 32'd203484789;
      4838: inst = 32'd471859200;
      4839: inst = 32'd136314880;
      4840: inst = 32'd268468224;
      4841: inst = 32'd201343912;
      4842: inst = 32'd203478060;
      4843: inst = 32'd471859200;
      4844: inst = 32'd136314880;
      4845: inst = 32'd268468224;
      4846: inst = 32'd201343913;
      4847: inst = 32'd203475655;
      4848: inst = 32'd471859200;
      4849: inst = 32'd136314880;
      4850: inst = 32'd268468224;
      4851: inst = 32'd201343914;
      4852: inst = 32'd203475655;
      4853: inst = 32'd471859200;
      4854: inst = 32'd136314880;
      4855: inst = 32'd268468224;
      4856: inst = 32'd201343915;
      4857: inst = 32'd203475655;
      4858: inst = 32'd471859200;
      4859: inst = 32'd136314880;
      4860: inst = 32'd268468224;
      4861: inst = 32'd201343916;
      4862: inst = 32'd203475655;
      4863: inst = 32'd471859200;
      4864: inst = 32'd136314880;
      4865: inst = 32'd268468224;
      4866: inst = 32'd201343917;
      4867: inst = 32'd203475655;
      4868: inst = 32'd471859200;
      4869: inst = 32'd136314880;
      4870: inst = 32'd268468224;
      4871: inst = 32'd201343918;
      4872: inst = 32'd203475655;
      4873: inst = 32'd471859200;
      4874: inst = 32'd136314880;
      4875: inst = 32'd268468224;
      4876: inst = 32'd201343919;
      4877: inst = 32'd203478028;
      4878: inst = 32'd471859200;
      4879: inst = 32'd136314880;
      4880: inst = 32'd268468224;
      4881: inst = 32'd201343920;
      4882: inst = 32'd203484757;
      4883: inst = 32'd471859200;
      4884: inst = 32'd136314880;
      4885: inst = 32'd268468224;
      4886: inst = 32'd201343921;
      4887: inst = 32'd203484854;
      4888: inst = 32'd471859200;
      4889: inst = 32'd136314880;
      4890: inst = 32'd268468224;
      4891: inst = 32'd201343922;
      4892: inst = 32'd203484854;
      4893: inst = 32'd471859200;
      4894: inst = 32'd136314880;
      4895: inst = 32'd268468224;
      4896: inst = 32'd201343923;
      4897: inst = 32'd203484854;
      4898: inst = 32'd471859200;
      4899: inst = 32'd136314880;
      4900: inst = 32'd268468224;
      4901: inst = 32'd201343924;
      4902: inst = 32'd203484854;
      4903: inst = 32'd471859200;
      4904: inst = 32'd136314880;
      4905: inst = 32'd268468224;
      4906: inst = 32'd201343925;
      4907: inst = 32'd203484854;
      4908: inst = 32'd471859200;
      4909: inst = 32'd136314880;
      4910: inst = 32'd268468224;
      4911: inst = 32'd201343926;
      4912: inst = 32'd203484854;
      4913: inst = 32'd471859200;
      4914: inst = 32'd136314880;
      4915: inst = 32'd268468224;
      4916: inst = 32'd201343927;
      4917: inst = 32'd203484854;
      4918: inst = 32'd471859200;
      4919: inst = 32'd136314880;
      4920: inst = 32'd268468224;
      4921: inst = 32'd201343928;
      4922: inst = 32'd203484854;
      4923: inst = 32'd471859200;
      4924: inst = 32'd136314880;
      4925: inst = 32'd268468224;
      4926: inst = 32'd201343929;
      4927: inst = 32'd203484854;
      4928: inst = 32'd471859200;
      4929: inst = 32'd136314880;
      4930: inst = 32'd268468224;
      4931: inst = 32'd201343930;
      4932: inst = 32'd203484854;
      4933: inst = 32'd471859200;
      4934: inst = 32'd136314880;
      4935: inst = 32'd268468224;
      4936: inst = 32'd201343931;
      4937: inst = 32'd203484854;
      4938: inst = 32'd471859200;
      4939: inst = 32'd136314880;
      4940: inst = 32'd268468224;
      4941: inst = 32'd201343932;
      4942: inst = 32'd203489279;
      4943: inst = 32'd471859200;
      4944: inst = 32'd136314880;
      4945: inst = 32'd268468224;
      4946: inst = 32'd201343933;
      4947: inst = 32'd203489279;
      4948: inst = 32'd471859200;
      4949: inst = 32'd136314880;
      4950: inst = 32'd268468224;
      4951: inst = 32'd201343934;
      4952: inst = 32'd203489279;
      4953: inst = 32'd471859200;
      4954: inst = 32'd136314880;
      4955: inst = 32'd268468224;
      4956: inst = 32'd201343935;
      4957: inst = 32'd203489279;
      4958: inst = 32'd471859200;
      4959: inst = 32'd136314880;
      4960: inst = 32'd268468224;
      4961: inst = 32'd201343936;
      4962: inst = 32'd203489279;
      4963: inst = 32'd471859200;
      4964: inst = 32'd136314880;
      4965: inst = 32'd268468224;
      4966: inst = 32'd201343937;
      4967: inst = 32'd203489279;
      4968: inst = 32'd471859200;
      4969: inst = 32'd136314880;
      4970: inst = 32'd268468224;
      4971: inst = 32'd201343938;
      4972: inst = 32'd203489279;
      4973: inst = 32'd471859200;
      4974: inst = 32'd136314880;
      4975: inst = 32'd268468224;
      4976: inst = 32'd201343939;
      4977: inst = 32'd203489279;
      4978: inst = 32'd471859200;
      4979: inst = 32'd136314880;
      4980: inst = 32'd268468224;
      4981: inst = 32'd201343940;
      4982: inst = 32'd203489279;
      4983: inst = 32'd471859200;
      4984: inst = 32'd136314880;
      4985: inst = 32'd268468224;
      4986: inst = 32'd201343941;
      4987: inst = 32'd203489279;
      4988: inst = 32'd471859200;
      4989: inst = 32'd136314880;
      4990: inst = 32'd268468224;
      4991: inst = 32'd201343942;
      4992: inst = 32'd203489279;
      4993: inst = 32'd471859200;
      4994: inst = 32'd136314880;
      4995: inst = 32'd268468224;
      4996: inst = 32'd201343943;
      4997: inst = 32'd203489279;
      4998: inst = 32'd471859200;
      4999: inst = 32'd136314880;
      5000: inst = 32'd268468224;
      5001: inst = 32'd201343944;
      5002: inst = 32'd203489279;
      5003: inst = 32'd471859200;
      5004: inst = 32'd136314880;
      5005: inst = 32'd268468224;
      5006: inst = 32'd201343945;
      5007: inst = 32'd203489279;
      5008: inst = 32'd471859200;
      5009: inst = 32'd136314880;
      5010: inst = 32'd268468224;
      5011: inst = 32'd201343946;
      5012: inst = 32'd203489279;
      5013: inst = 32'd471859200;
      5014: inst = 32'd136314880;
      5015: inst = 32'd268468224;
      5016: inst = 32'd201343947;
      5017: inst = 32'd203489279;
      5018: inst = 32'd471859200;
      5019: inst = 32'd136314880;
      5020: inst = 32'd268468224;
      5021: inst = 32'd201343948;
      5022: inst = 32'd203489279;
      5023: inst = 32'd471859200;
      5024: inst = 32'd136314880;
      5025: inst = 32'd268468224;
      5026: inst = 32'd201343949;
      5027: inst = 32'd203489279;
      5028: inst = 32'd471859200;
      5029: inst = 32'd136314880;
      5030: inst = 32'd268468224;
      5031: inst = 32'd201343950;
      5032: inst = 32'd203489279;
      5033: inst = 32'd471859200;
      5034: inst = 32'd136314880;
      5035: inst = 32'd268468224;
      5036: inst = 32'd201343951;
      5037: inst = 32'd203489279;
      5038: inst = 32'd471859200;
      5039: inst = 32'd136314880;
      5040: inst = 32'd268468224;
      5041: inst = 32'd201343952;
      5042: inst = 32'd203489279;
      5043: inst = 32'd471859200;
      5044: inst = 32'd136314880;
      5045: inst = 32'd268468224;
      5046: inst = 32'd201343953;
      5047: inst = 32'd203489279;
      5048: inst = 32'd471859200;
      5049: inst = 32'd136314880;
      5050: inst = 32'd268468224;
      5051: inst = 32'd201343954;
      5052: inst = 32'd203489279;
      5053: inst = 32'd471859200;
      5054: inst = 32'd136314880;
      5055: inst = 32'd268468224;
      5056: inst = 32'd201343955;
      5057: inst = 32'd203489279;
      5058: inst = 32'd471859200;
      5059: inst = 32'd136314880;
      5060: inst = 32'd268468224;
      5061: inst = 32'd201343956;
      5062: inst = 32'd203489279;
      5063: inst = 32'd471859200;
      5064: inst = 32'd136314880;
      5065: inst = 32'd268468224;
      5066: inst = 32'd201343957;
      5067: inst = 32'd203489279;
      5068: inst = 32'd471859200;
      5069: inst = 32'd136314880;
      5070: inst = 32'd268468224;
      5071: inst = 32'd201343958;
      5072: inst = 32'd203489279;
      5073: inst = 32'd471859200;
      5074: inst = 32'd136314880;
      5075: inst = 32'd268468224;
      5076: inst = 32'd201343959;
      5077: inst = 32'd203489279;
      5078: inst = 32'd471859200;
      5079: inst = 32'd136314880;
      5080: inst = 32'd268468224;
      5081: inst = 32'd201343960;
      5082: inst = 32'd203489279;
      5083: inst = 32'd471859200;
      5084: inst = 32'd136314880;
      5085: inst = 32'd268468224;
      5086: inst = 32'd201343961;
      5087: inst = 32'd203489279;
      5088: inst = 32'd471859200;
      5089: inst = 32'd136314880;
      5090: inst = 32'd268468224;
      5091: inst = 32'd201343962;
      5092: inst = 32'd203489279;
      5093: inst = 32'd471859200;
      5094: inst = 32'd136314880;
      5095: inst = 32'd268468224;
      5096: inst = 32'd201343963;
      5097: inst = 32'd203489279;
      5098: inst = 32'd471859200;
      5099: inst = 32'd136314880;
      5100: inst = 32'd268468224;
      5101: inst = 32'd201343964;
      5102: inst = 32'd203489279;
      5103: inst = 32'd471859200;
      5104: inst = 32'd136314880;
      5105: inst = 32'd268468224;
      5106: inst = 32'd201343965;
      5107: inst = 32'd203489279;
      5108: inst = 32'd471859200;
      5109: inst = 32'd136314880;
      5110: inst = 32'd268468224;
      5111: inst = 32'd201343966;
      5112: inst = 32'd203489279;
      5113: inst = 32'd471859200;
      5114: inst = 32'd136314880;
      5115: inst = 32'd268468224;
      5116: inst = 32'd201343967;
      5117: inst = 32'd203489279;
      5118: inst = 32'd471859200;
      5119: inst = 32'd136314880;
      5120: inst = 32'd268468224;
      5121: inst = 32'd201343968;
      5122: inst = 32'd203489279;
      5123: inst = 32'd471859200;
      5124: inst = 32'd136314880;
      5125: inst = 32'd268468224;
      5126: inst = 32'd201343969;
      5127: inst = 32'd203489279;
      5128: inst = 32'd471859200;
      5129: inst = 32'd136314880;
      5130: inst = 32'd268468224;
      5131: inst = 32'd201343970;
      5132: inst = 32'd203489279;
      5133: inst = 32'd471859200;
      5134: inst = 32'd136314880;
      5135: inst = 32'd268468224;
      5136: inst = 32'd201343971;
      5137: inst = 32'd203489279;
      5138: inst = 32'd471859200;
      5139: inst = 32'd136314880;
      5140: inst = 32'd268468224;
      5141: inst = 32'd201343972;
      5142: inst = 32'd203484854;
      5143: inst = 32'd471859200;
      5144: inst = 32'd136314880;
      5145: inst = 32'd268468224;
      5146: inst = 32'd201343973;
      5147: inst = 32'd203484854;
      5148: inst = 32'd471859200;
      5149: inst = 32'd136314880;
      5150: inst = 32'd268468224;
      5151: inst = 32'd201343974;
      5152: inst = 32'd203484854;
      5153: inst = 32'd471859200;
      5154: inst = 32'd136314880;
      5155: inst = 32'd268468224;
      5156: inst = 32'd201343975;
      5157: inst = 32'd203484854;
      5158: inst = 32'd471859200;
      5159: inst = 32'd136314880;
      5160: inst = 32'd268468224;
      5161: inst = 32'd201343976;
      5162: inst = 32'd203484854;
      5163: inst = 32'd471859200;
      5164: inst = 32'd136314880;
      5165: inst = 32'd268468224;
      5166: inst = 32'd201343977;
      5167: inst = 32'd203484854;
      5168: inst = 32'd471859200;
      5169: inst = 32'd136314880;
      5170: inst = 32'd268468224;
      5171: inst = 32'd201343978;
      5172: inst = 32'd203484854;
      5173: inst = 32'd471859200;
      5174: inst = 32'd136314880;
      5175: inst = 32'd268468224;
      5176: inst = 32'd201343979;
      5177: inst = 32'd203484854;
      5178: inst = 32'd471859200;
      5179: inst = 32'd136314880;
      5180: inst = 32'd268468224;
      5181: inst = 32'd201343980;
      5182: inst = 32'd203484854;
      5183: inst = 32'd471859200;
      5184: inst = 32'd136314880;
      5185: inst = 32'd268468224;
      5186: inst = 32'd201343981;
      5187: inst = 32'd203484854;
      5188: inst = 32'd471859200;
      5189: inst = 32'd136314880;
      5190: inst = 32'd268468224;
      5191: inst = 32'd201343982;
      5192: inst = 32'd203484854;
      5193: inst = 32'd471859200;
      5194: inst = 32'd136314880;
      5195: inst = 32'd268468224;
      5196: inst = 32'd201343983;
      5197: inst = 32'd203484854;
      5198: inst = 32'd471859200;
      5199: inst = 32'd136314880;
      5200: inst = 32'd268468224;
      5201: inst = 32'd201343984;
      5202: inst = 32'd203484854;
      5203: inst = 32'd471859200;
      5204: inst = 32'd136314880;
      5205: inst = 32'd268468224;
      5206: inst = 32'd201343985;
      5207: inst = 32'd203484854;
      5208: inst = 32'd471859200;
      5209: inst = 32'd136314880;
      5210: inst = 32'd268468224;
      5211: inst = 32'd201343986;
      5212: inst = 32'd203484854;
      5213: inst = 32'd471859200;
      5214: inst = 32'd136314880;
      5215: inst = 32'd268468224;
      5216: inst = 32'd201343987;
      5217: inst = 32'd203484854;
      5218: inst = 32'd471859200;
      5219: inst = 32'd136314880;
      5220: inst = 32'd268468224;
      5221: inst = 32'd201343988;
      5222: inst = 32'd203484854;
      5223: inst = 32'd471859200;
      5224: inst = 32'd136314880;
      5225: inst = 32'd268468224;
      5226: inst = 32'd201343989;
      5227: inst = 32'd203484854;
      5228: inst = 32'd471859200;
      5229: inst = 32'd136314880;
      5230: inst = 32'd268468224;
      5231: inst = 32'd201343990;
      5232: inst = 32'd203484854;
      5233: inst = 32'd471859200;
      5234: inst = 32'd136314880;
      5235: inst = 32'd268468224;
      5236: inst = 32'd201343991;
      5237: inst = 32'd203484854;
      5238: inst = 32'd471859200;
      5239: inst = 32'd136314880;
      5240: inst = 32'd268468224;
      5241: inst = 32'd201343992;
      5242: inst = 32'd203484854;
      5243: inst = 32'd471859200;
      5244: inst = 32'd136314880;
      5245: inst = 32'd268468224;
      5246: inst = 32'd201343993;
      5247: inst = 32'd203484854;
      5248: inst = 32'd471859200;
      5249: inst = 32'd136314880;
      5250: inst = 32'd268468224;
      5251: inst = 32'd201343994;
      5252: inst = 32'd203484854;
      5253: inst = 32'd471859200;
      5254: inst = 32'd136314880;
      5255: inst = 32'd268468224;
      5256: inst = 32'd201343995;
      5257: inst = 32'd203484854;
      5258: inst = 32'd471859200;
      5259: inst = 32'd136314880;
      5260: inst = 32'd268468224;
      5261: inst = 32'd201343996;
      5262: inst = 32'd203484854;
      5263: inst = 32'd471859200;
      5264: inst = 32'd136314880;
      5265: inst = 32'd268468224;
      5266: inst = 32'd201343997;
      5267: inst = 32'd203484854;
      5268: inst = 32'd471859200;
      5269: inst = 32'd136314880;
      5270: inst = 32'd268468224;
      5271: inst = 32'd201343998;
      5272: inst = 32'd203484854;
      5273: inst = 32'd471859200;
      5274: inst = 32'd136314880;
      5275: inst = 32'd268468224;
      5276: inst = 32'd201343999;
      5277: inst = 32'd203484854;
      5278: inst = 32'd471859200;
      5279: inst = 32'd136314880;
      5280: inst = 32'd268468224;
      5281: inst = 32'd201344000;
      5282: inst = 32'd203484854;
      5283: inst = 32'd471859200;
      5284: inst = 32'd136314880;
      5285: inst = 32'd268468224;
      5286: inst = 32'd201344001;
      5287: inst = 32'd203484854;
      5288: inst = 32'd471859200;
      5289: inst = 32'd136314880;
      5290: inst = 32'd268468224;
      5291: inst = 32'd201344002;
      5292: inst = 32'd203484854;
      5293: inst = 32'd471859200;
      5294: inst = 32'd136314880;
      5295: inst = 32'd268468224;
      5296: inst = 32'd201344003;
      5297: inst = 32'd203484854;
      5298: inst = 32'd471859200;
      5299: inst = 32'd136314880;
      5300: inst = 32'd268468224;
      5301: inst = 32'd201344004;
      5302: inst = 32'd203484854;
      5303: inst = 32'd471859200;
      5304: inst = 32'd136314880;
      5305: inst = 32'd268468224;
      5306: inst = 32'd201344005;
      5307: inst = 32'd203484854;
      5308: inst = 32'd471859200;
      5309: inst = 32'd136314880;
      5310: inst = 32'd268468224;
      5311: inst = 32'd201344006;
      5312: inst = 32'd203482481;
      5313: inst = 32'd471859200;
      5314: inst = 32'd136314880;
      5315: inst = 32'd268468224;
      5316: inst = 32'd201344007;
      5317: inst = 32'd203475752;
      5318: inst = 32'd471859200;
      5319: inst = 32'd136314880;
      5320: inst = 32'd268468224;
      5321: inst = 32'd201344008;
      5322: inst = 32'd203475655;
      5323: inst = 32'd471859200;
      5324: inst = 32'd136314880;
      5325: inst = 32'd268468224;
      5326: inst = 32'd201344009;
      5327: inst = 32'd203475655;
      5328: inst = 32'd471859200;
      5329: inst = 32'd136314880;
      5330: inst = 32'd268468224;
      5331: inst = 32'd201344010;
      5332: inst = 32'd203475655;
      5333: inst = 32'd471859200;
      5334: inst = 32'd136314880;
      5335: inst = 32'd268468224;
      5336: inst = 32'd201344011;
      5337: inst = 32'd203475655;
      5338: inst = 32'd471859200;
      5339: inst = 32'd136314880;
      5340: inst = 32'd268468224;
      5341: inst = 32'd201344012;
      5342: inst = 32'd203475655;
      5343: inst = 32'd471859200;
      5344: inst = 32'd136314880;
      5345: inst = 32'd268468224;
      5346: inst = 32'd201344013;
      5347: inst = 32'd203475655;
      5348: inst = 32'd471859200;
      5349: inst = 32'd136314880;
      5350: inst = 32'd268468224;
      5351: inst = 32'd201344014;
      5352: inst = 32'd203475655;
      5353: inst = 32'd471859200;
      5354: inst = 32'd136314880;
      5355: inst = 32'd268468224;
      5356: inst = 32'd201344015;
      5357: inst = 32'd203475655;
      5358: inst = 32'd471859200;
      5359: inst = 32'd136314880;
      5360: inst = 32'd268468224;
      5361: inst = 32'd201344016;
      5362: inst = 32'd203475752;
      5363: inst = 32'd471859200;
      5364: inst = 32'd136314880;
      5365: inst = 32'd268468224;
      5366: inst = 32'd201344017;
      5367: inst = 32'd203482481;
      5368: inst = 32'd471859200;
      5369: inst = 32'd136314880;
      5370: inst = 32'd268468224;
      5371: inst = 32'd201344018;
      5372: inst = 32'd203484854;
      5373: inst = 32'd471859200;
      5374: inst = 32'd136314880;
      5375: inst = 32'd268468224;
      5376: inst = 32'd201344019;
      5377: inst = 32'd203484854;
      5378: inst = 32'd471859200;
      5379: inst = 32'd136314880;
      5380: inst = 32'd268468224;
      5381: inst = 32'd201344020;
      5382: inst = 32'd203484854;
      5383: inst = 32'd471859200;
      5384: inst = 32'd136314880;
      5385: inst = 32'd268468224;
      5386: inst = 32'd201344021;
      5387: inst = 32'd203484854;
      5388: inst = 32'd471859200;
      5389: inst = 32'd136314880;
      5390: inst = 32'd268468224;
      5391: inst = 32'd201344022;
      5392: inst = 32'd203484854;
      5393: inst = 32'd471859200;
      5394: inst = 32'd136314880;
      5395: inst = 32'd268468224;
      5396: inst = 32'd201344023;
      5397: inst = 32'd203484854;
      5398: inst = 32'd471859200;
      5399: inst = 32'd136314880;
      5400: inst = 32'd268468224;
      5401: inst = 32'd201344024;
      5402: inst = 32'd203484854;
      5403: inst = 32'd471859200;
      5404: inst = 32'd136314880;
      5405: inst = 32'd268468224;
      5406: inst = 32'd201344025;
      5407: inst = 32'd203484854;
      5408: inst = 32'd471859200;
      5409: inst = 32'd136314880;
      5410: inst = 32'd268468224;
      5411: inst = 32'd201344026;
      5412: inst = 32'd203484854;
      5413: inst = 32'd471859200;
      5414: inst = 32'd136314880;
      5415: inst = 32'd268468224;
      5416: inst = 32'd201344027;
      5417: inst = 32'd203484854;
      5418: inst = 32'd471859200;
      5419: inst = 32'd136314880;
      5420: inst = 32'd268468224;
      5421: inst = 32'd201344028;
      5422: inst = 32'd203489279;
      5423: inst = 32'd471859200;
      5424: inst = 32'd136314880;
      5425: inst = 32'd268468224;
      5426: inst = 32'd201344029;
      5427: inst = 32'd203489279;
      5428: inst = 32'd471859200;
      5429: inst = 32'd136314880;
      5430: inst = 32'd268468224;
      5431: inst = 32'd201344030;
      5432: inst = 32'd203489279;
      5433: inst = 32'd471859200;
      5434: inst = 32'd136314880;
      5435: inst = 32'd268468224;
      5436: inst = 32'd201344031;
      5437: inst = 32'd203489279;
      5438: inst = 32'd471859200;
      5439: inst = 32'd136314880;
      5440: inst = 32'd268468224;
      5441: inst = 32'd201344032;
      5442: inst = 32'd203489279;
      5443: inst = 32'd471859200;
      5444: inst = 32'd136314880;
      5445: inst = 32'd268468224;
      5446: inst = 32'd201344033;
      5447: inst = 32'd203489279;
      5448: inst = 32'd471859200;
      5449: inst = 32'd136314880;
      5450: inst = 32'd268468224;
      5451: inst = 32'd201344034;
      5452: inst = 32'd203489279;
      5453: inst = 32'd471859200;
      5454: inst = 32'd136314880;
      5455: inst = 32'd268468224;
      5456: inst = 32'd201344035;
      5457: inst = 32'd203489279;
      5458: inst = 32'd471859200;
      5459: inst = 32'd136314880;
      5460: inst = 32'd268468224;
      5461: inst = 32'd201344036;
      5462: inst = 32'd203489279;
      5463: inst = 32'd471859200;
      5464: inst = 32'd136314880;
      5465: inst = 32'd268468224;
      5466: inst = 32'd201344037;
      5467: inst = 32'd203489279;
      5468: inst = 32'd471859200;
      5469: inst = 32'd136314880;
      5470: inst = 32'd268468224;
      5471: inst = 32'd201344038;
      5472: inst = 32'd203489279;
      5473: inst = 32'd471859200;
      5474: inst = 32'd136314880;
      5475: inst = 32'd268468224;
      5476: inst = 32'd201344039;
      5477: inst = 32'd203489279;
      5478: inst = 32'd471859200;
      5479: inst = 32'd136314880;
      5480: inst = 32'd268468224;
      5481: inst = 32'd201344040;
      5482: inst = 32'd203489279;
      5483: inst = 32'd471859200;
      5484: inst = 32'd136314880;
      5485: inst = 32'd268468224;
      5486: inst = 32'd201344041;
      5487: inst = 32'd203489279;
      5488: inst = 32'd471859200;
      5489: inst = 32'd136314880;
      5490: inst = 32'd268468224;
      5491: inst = 32'd201344042;
      5492: inst = 32'd203489279;
      5493: inst = 32'd471859200;
      5494: inst = 32'd136314880;
      5495: inst = 32'd268468224;
      5496: inst = 32'd201344043;
      5497: inst = 32'd203489279;
      5498: inst = 32'd471859200;
      5499: inst = 32'd136314880;
      5500: inst = 32'd268468224;
      5501: inst = 32'd201344044;
      5502: inst = 32'd203489279;
      5503: inst = 32'd471859200;
      5504: inst = 32'd136314880;
      5505: inst = 32'd268468224;
      5506: inst = 32'd201344045;
      5507: inst = 32'd203489279;
      5508: inst = 32'd471859200;
      5509: inst = 32'd136314880;
      5510: inst = 32'd268468224;
      5511: inst = 32'd201344046;
      5512: inst = 32'd203489279;
      5513: inst = 32'd471859200;
      5514: inst = 32'd136314880;
      5515: inst = 32'd268468224;
      5516: inst = 32'd201344047;
      5517: inst = 32'd203489279;
      5518: inst = 32'd471859200;
      5519: inst = 32'd136314880;
      5520: inst = 32'd268468224;
      5521: inst = 32'd201344048;
      5522: inst = 32'd203489279;
      5523: inst = 32'd471859200;
      5524: inst = 32'd136314880;
      5525: inst = 32'd268468224;
      5526: inst = 32'd201344049;
      5527: inst = 32'd203489279;
      5528: inst = 32'd471859200;
      5529: inst = 32'd136314880;
      5530: inst = 32'd268468224;
      5531: inst = 32'd201344050;
      5532: inst = 32'd203489279;
      5533: inst = 32'd471859200;
      5534: inst = 32'd136314880;
      5535: inst = 32'd268468224;
      5536: inst = 32'd201344051;
      5537: inst = 32'd203489279;
      5538: inst = 32'd471859200;
      5539: inst = 32'd136314880;
      5540: inst = 32'd268468224;
      5541: inst = 32'd201344052;
      5542: inst = 32'd203489279;
      5543: inst = 32'd471859200;
      5544: inst = 32'd136314880;
      5545: inst = 32'd268468224;
      5546: inst = 32'd201344053;
      5547: inst = 32'd203489279;
      5548: inst = 32'd471859200;
      5549: inst = 32'd136314880;
      5550: inst = 32'd268468224;
      5551: inst = 32'd201344054;
      5552: inst = 32'd203489279;
      5553: inst = 32'd471859200;
      5554: inst = 32'd136314880;
      5555: inst = 32'd268468224;
      5556: inst = 32'd201344055;
      5557: inst = 32'd203489279;
      5558: inst = 32'd471859200;
      5559: inst = 32'd136314880;
      5560: inst = 32'd268468224;
      5561: inst = 32'd201344056;
      5562: inst = 32'd203489279;
      5563: inst = 32'd471859200;
      5564: inst = 32'd136314880;
      5565: inst = 32'd268468224;
      5566: inst = 32'd201344057;
      5567: inst = 32'd203489279;
      5568: inst = 32'd471859200;
      5569: inst = 32'd136314880;
      5570: inst = 32'd268468224;
      5571: inst = 32'd201344058;
      5572: inst = 32'd203489279;
      5573: inst = 32'd471859200;
      5574: inst = 32'd136314880;
      5575: inst = 32'd268468224;
      5576: inst = 32'd201344059;
      5577: inst = 32'd203489279;
      5578: inst = 32'd471859200;
      5579: inst = 32'd136314880;
      5580: inst = 32'd268468224;
      5581: inst = 32'd201344060;
      5582: inst = 32'd203489279;
      5583: inst = 32'd471859200;
      5584: inst = 32'd136314880;
      5585: inst = 32'd268468224;
      5586: inst = 32'd201344061;
      5587: inst = 32'd203489279;
      5588: inst = 32'd471859200;
      5589: inst = 32'd136314880;
      5590: inst = 32'd268468224;
      5591: inst = 32'd201344062;
      5592: inst = 32'd203489279;
      5593: inst = 32'd471859200;
      5594: inst = 32'd136314880;
      5595: inst = 32'd268468224;
      5596: inst = 32'd201344063;
      5597: inst = 32'd203489279;
      5598: inst = 32'd471859200;
      5599: inst = 32'd136314880;
      5600: inst = 32'd268468224;
      5601: inst = 32'd201344064;
      5602: inst = 32'd203489279;
      5603: inst = 32'd471859200;
      5604: inst = 32'd136314880;
      5605: inst = 32'd268468224;
      5606: inst = 32'd201344065;
      5607: inst = 32'd203489279;
      5608: inst = 32'd471859200;
      5609: inst = 32'd136314880;
      5610: inst = 32'd268468224;
      5611: inst = 32'd201344066;
      5612: inst = 32'd203489279;
      5613: inst = 32'd471859200;
      5614: inst = 32'd136314880;
      5615: inst = 32'd268468224;
      5616: inst = 32'd201344067;
      5617: inst = 32'd203489279;
      5618: inst = 32'd471859200;
      5619: inst = 32'd136314880;
      5620: inst = 32'd268468224;
      5621: inst = 32'd201344068;
      5622: inst = 32'd203484854;
      5623: inst = 32'd471859200;
      5624: inst = 32'd136314880;
      5625: inst = 32'd268468224;
      5626: inst = 32'd201344069;
      5627: inst = 32'd203484854;
      5628: inst = 32'd471859200;
      5629: inst = 32'd136314880;
      5630: inst = 32'd268468224;
      5631: inst = 32'd201344070;
      5632: inst = 32'd203484854;
      5633: inst = 32'd471859200;
      5634: inst = 32'd136314880;
      5635: inst = 32'd268468224;
      5636: inst = 32'd201344071;
      5637: inst = 32'd203484854;
      5638: inst = 32'd471859200;
      5639: inst = 32'd136314880;
      5640: inst = 32'd268468224;
      5641: inst = 32'd201344072;
      5642: inst = 32'd203484854;
      5643: inst = 32'd471859200;
      5644: inst = 32'd136314880;
      5645: inst = 32'd268468224;
      5646: inst = 32'd201344073;
      5647: inst = 32'd203484854;
      5648: inst = 32'd471859200;
      5649: inst = 32'd136314880;
      5650: inst = 32'd268468224;
      5651: inst = 32'd201344074;
      5652: inst = 32'd203484854;
      5653: inst = 32'd471859200;
      5654: inst = 32'd136314880;
      5655: inst = 32'd268468224;
      5656: inst = 32'd201344075;
      5657: inst = 32'd203484854;
      5658: inst = 32'd471859200;
      5659: inst = 32'd136314880;
      5660: inst = 32'd268468224;
      5661: inst = 32'd201344076;
      5662: inst = 32'd203484854;
      5663: inst = 32'd471859200;
      5664: inst = 32'd136314880;
      5665: inst = 32'd268468224;
      5666: inst = 32'd201344077;
      5667: inst = 32'd203484854;
      5668: inst = 32'd471859200;
      5669: inst = 32'd136314880;
      5670: inst = 32'd268468224;
      5671: inst = 32'd201344078;
      5672: inst = 32'd203484854;
      5673: inst = 32'd471859200;
      5674: inst = 32'd136314880;
      5675: inst = 32'd268468224;
      5676: inst = 32'd201344079;
      5677: inst = 32'd203484854;
      5678: inst = 32'd471859200;
      5679: inst = 32'd136314880;
      5680: inst = 32'd268468224;
      5681: inst = 32'd201344080;
      5682: inst = 32'd203484854;
      5683: inst = 32'd471859200;
      5684: inst = 32'd136314880;
      5685: inst = 32'd268468224;
      5686: inst = 32'd201344081;
      5687: inst = 32'd203484854;
      5688: inst = 32'd471859200;
      5689: inst = 32'd136314880;
      5690: inst = 32'd268468224;
      5691: inst = 32'd201344082;
      5692: inst = 32'd203484854;
      5693: inst = 32'd471859200;
      5694: inst = 32'd136314880;
      5695: inst = 32'd268468224;
      5696: inst = 32'd201344083;
      5697: inst = 32'd203484854;
      5698: inst = 32'd471859200;
      5699: inst = 32'd136314880;
      5700: inst = 32'd268468224;
      5701: inst = 32'd201344084;
      5702: inst = 32'd203484854;
      5703: inst = 32'd471859200;
      5704: inst = 32'd136314880;
      5705: inst = 32'd268468224;
      5706: inst = 32'd201344085;
      5707: inst = 32'd203484854;
      5708: inst = 32'd471859200;
      5709: inst = 32'd136314880;
      5710: inst = 32'd268468224;
      5711: inst = 32'd201344086;
      5712: inst = 32'd203484854;
      5713: inst = 32'd471859200;
      5714: inst = 32'd136314880;
      5715: inst = 32'd268468224;
      5716: inst = 32'd201344087;
      5717: inst = 32'd203484854;
      5718: inst = 32'd471859200;
      5719: inst = 32'd136314880;
      5720: inst = 32'd268468224;
      5721: inst = 32'd201344088;
      5722: inst = 32'd203484854;
      5723: inst = 32'd471859200;
      5724: inst = 32'd136314880;
      5725: inst = 32'd268468224;
      5726: inst = 32'd201344089;
      5727: inst = 32'd203484854;
      5728: inst = 32'd471859200;
      5729: inst = 32'd136314880;
      5730: inst = 32'd268468224;
      5731: inst = 32'd201344090;
      5732: inst = 32'd203484854;
      5733: inst = 32'd471859200;
      5734: inst = 32'd136314880;
      5735: inst = 32'd268468224;
      5736: inst = 32'd201344091;
      5737: inst = 32'd203484854;
      5738: inst = 32'd471859200;
      5739: inst = 32'd136314880;
      5740: inst = 32'd268468224;
      5741: inst = 32'd201344092;
      5742: inst = 32'd203484854;
      5743: inst = 32'd471859200;
      5744: inst = 32'd136314880;
      5745: inst = 32'd268468224;
      5746: inst = 32'd201344093;
      5747: inst = 32'd203484854;
      5748: inst = 32'd471859200;
      5749: inst = 32'd136314880;
      5750: inst = 32'd268468224;
      5751: inst = 32'd201344094;
      5752: inst = 32'd203484854;
      5753: inst = 32'd471859200;
      5754: inst = 32'd136314880;
      5755: inst = 32'd268468224;
      5756: inst = 32'd201344095;
      5757: inst = 32'd203484854;
      5758: inst = 32'd471859200;
      5759: inst = 32'd136314880;
      5760: inst = 32'd268468224;
      5761: inst = 32'd201344096;
      5762: inst = 32'd203484854;
      5763: inst = 32'd471859200;
      5764: inst = 32'd136314880;
      5765: inst = 32'd268468224;
      5766: inst = 32'd201344097;
      5767: inst = 32'd203484854;
      5768: inst = 32'd471859200;
      5769: inst = 32'd136314880;
      5770: inst = 32'd268468224;
      5771: inst = 32'd201344098;
      5772: inst = 32'd203484854;
      5773: inst = 32'd471859200;
      5774: inst = 32'd136314880;
      5775: inst = 32'd268468224;
      5776: inst = 32'd201344099;
      5777: inst = 32'd203484854;
      5778: inst = 32'd471859200;
      5779: inst = 32'd136314880;
      5780: inst = 32'd268468224;
      5781: inst = 32'd201344100;
      5782: inst = 32'd203484854;
      5783: inst = 32'd471859200;
      5784: inst = 32'd136314880;
      5785: inst = 32'd268468224;
      5786: inst = 32'd201344101;
      5787: inst = 32'd203484854;
      5788: inst = 32'd471859200;
      5789: inst = 32'd136314880;
      5790: inst = 32'd268468224;
      5791: inst = 32'd201344102;
      5792: inst = 32'd203484854;
      5793: inst = 32'd471859200;
      5794: inst = 32'd136314880;
      5795: inst = 32'd268468224;
      5796: inst = 32'd201344103;
      5797: inst = 32'd203484854;
      5798: inst = 32'd471859200;
      5799: inst = 32'd136314880;
      5800: inst = 32'd268468224;
      5801: inst = 32'd201344104;
      5802: inst = 32'd203484854;
      5803: inst = 32'd471859200;
      5804: inst = 32'd136314880;
      5805: inst = 32'd268468224;
      5806: inst = 32'd201344105;
      5807: inst = 32'd203484854;
      5808: inst = 32'd471859200;
      5809: inst = 32'd136314880;
      5810: inst = 32'd268468224;
      5811: inst = 32'd201344106;
      5812: inst = 32'd203484814;
      5813: inst = 32'd471859200;
      5814: inst = 32'd136314880;
      5815: inst = 32'd268468224;
      5816: inst = 32'd201344107;
      5817: inst = 32'd203484744;
      5818: inst = 32'd471859200;
      5819: inst = 32'd136314880;
      5820: inst = 32'd268468224;
      5821: inst = 32'd201344108;
      5822: inst = 32'd203484744;
      5823: inst = 32'd471859200;
      5824: inst = 32'd136314880;
      5825: inst = 32'd268468224;
      5826: inst = 32'd201344109;
      5827: inst = 32'd203484816;
      5828: inst = 32'd471859200;
      5829: inst = 32'd136314880;
      5830: inst = 32'd268468224;
      5831: inst = 32'd201344110;
      5832: inst = 32'd203484854;
      5833: inst = 32'd471859200;
      5834: inst = 32'd136314880;
      5835: inst = 32'd268468224;
      5836: inst = 32'd201344111;
      5837: inst = 32'd203484854;
      5838: inst = 32'd471859200;
      5839: inst = 32'd136314880;
      5840: inst = 32'd268468224;
      5841: inst = 32'd201344112;
      5842: inst = 32'd203484854;
      5843: inst = 32'd471859200;
      5844: inst = 32'd136314880;
      5845: inst = 32'd268468224;
      5846: inst = 32'd201344113;
      5847: inst = 32'd203484854;
      5848: inst = 32'd471859200;
      5849: inst = 32'd136314880;
      5850: inst = 32'd268468224;
      5851: inst = 32'd201344114;
      5852: inst = 32'd203484854;
      5853: inst = 32'd471859200;
      5854: inst = 32'd136314880;
      5855: inst = 32'd268468224;
      5856: inst = 32'd201344115;
      5857: inst = 32'd203484854;
      5858: inst = 32'd471859200;
      5859: inst = 32'd136314880;
      5860: inst = 32'd268468224;
      5861: inst = 32'd201344116;
      5862: inst = 32'd203484854;
      5863: inst = 32'd471859200;
      5864: inst = 32'd136314880;
      5865: inst = 32'd268468224;
      5866: inst = 32'd201344117;
      5867: inst = 32'd203484854;
      5868: inst = 32'd471859200;
      5869: inst = 32'd136314880;
      5870: inst = 32'd268468224;
      5871: inst = 32'd201344118;
      5872: inst = 32'd203484854;
      5873: inst = 32'd471859200;
      5874: inst = 32'd136314880;
      5875: inst = 32'd268468224;
      5876: inst = 32'd201344119;
      5877: inst = 32'd203484854;
      5878: inst = 32'd471859200;
      5879: inst = 32'd136314880;
      5880: inst = 32'd268468224;
      5881: inst = 32'd201344120;
      5882: inst = 32'd203484854;
      5883: inst = 32'd471859200;
      5884: inst = 32'd136314880;
      5885: inst = 32'd268468224;
      5886: inst = 32'd201344121;
      5887: inst = 32'd203484854;
      5888: inst = 32'd471859200;
      5889: inst = 32'd136314880;
      5890: inst = 32'd268468224;
      5891: inst = 32'd201344122;
      5892: inst = 32'd203484854;
      5893: inst = 32'd471859200;
      5894: inst = 32'd136314880;
      5895: inst = 32'd268468224;
      5896: inst = 32'd201344123;
      5897: inst = 32'd203484854;
      5898: inst = 32'd471859200;
      5899: inst = 32'd136314880;
      5900: inst = 32'd268468224;
      5901: inst = 32'd201344124;
      5902: inst = 32'd203489279;
      5903: inst = 32'd471859200;
      5904: inst = 32'd136314880;
      5905: inst = 32'd268468224;
      5906: inst = 32'd201344125;
      5907: inst = 32'd203489279;
      5908: inst = 32'd471859200;
      5909: inst = 32'd136314880;
      5910: inst = 32'd268468224;
      5911: inst = 32'd201344126;
      5912: inst = 32'd203489279;
      5913: inst = 32'd471859200;
      5914: inst = 32'd136314880;
      5915: inst = 32'd268468224;
      5916: inst = 32'd201344127;
      5917: inst = 32'd203489279;
      5918: inst = 32'd471859200;
      5919: inst = 32'd136314880;
      5920: inst = 32'd268468224;
      5921: inst = 32'd201344128;
      5922: inst = 32'd203489279;
      5923: inst = 32'd471859200;
      5924: inst = 32'd136314880;
      5925: inst = 32'd268468224;
      5926: inst = 32'd201344129;
      5927: inst = 32'd203489279;
      5928: inst = 32'd471859200;
      5929: inst = 32'd136314880;
      5930: inst = 32'd268468224;
      5931: inst = 32'd201344130;
      5932: inst = 32'd203489279;
      5933: inst = 32'd471859200;
      5934: inst = 32'd136314880;
      5935: inst = 32'd268468224;
      5936: inst = 32'd201344131;
      5937: inst = 32'd203489279;
      5938: inst = 32'd471859200;
      5939: inst = 32'd136314880;
      5940: inst = 32'd268468224;
      5941: inst = 32'd201344132;
      5942: inst = 32'd203489279;
      5943: inst = 32'd471859200;
      5944: inst = 32'd136314880;
      5945: inst = 32'd268468224;
      5946: inst = 32'd201344133;
      5947: inst = 32'd203489279;
      5948: inst = 32'd471859200;
      5949: inst = 32'd136314880;
      5950: inst = 32'd268468224;
      5951: inst = 32'd201344134;
      5952: inst = 32'd203489279;
      5953: inst = 32'd471859200;
      5954: inst = 32'd136314880;
      5955: inst = 32'd268468224;
      5956: inst = 32'd201344135;
      5957: inst = 32'd203489279;
      5958: inst = 32'd471859200;
      5959: inst = 32'd136314880;
      5960: inst = 32'd268468224;
      5961: inst = 32'd201344136;
      5962: inst = 32'd203489279;
      5963: inst = 32'd471859200;
      5964: inst = 32'd136314880;
      5965: inst = 32'd268468224;
      5966: inst = 32'd201344137;
      5967: inst = 32'd203489279;
      5968: inst = 32'd471859200;
      5969: inst = 32'd136314880;
      5970: inst = 32'd268468224;
      5971: inst = 32'd201344138;
      5972: inst = 32'd203489279;
      5973: inst = 32'd471859200;
      5974: inst = 32'd136314880;
      5975: inst = 32'd268468224;
      5976: inst = 32'd201344139;
      5977: inst = 32'd203489279;
      5978: inst = 32'd471859200;
      5979: inst = 32'd136314880;
      5980: inst = 32'd268468224;
      5981: inst = 32'd201344140;
      5982: inst = 32'd203489279;
      5983: inst = 32'd471859200;
      5984: inst = 32'd136314880;
      5985: inst = 32'd268468224;
      5986: inst = 32'd201344141;
      5987: inst = 32'd203489279;
      5988: inst = 32'd471859200;
      5989: inst = 32'd136314880;
      5990: inst = 32'd268468224;
      5991: inst = 32'd201344142;
      5992: inst = 32'd203489279;
      5993: inst = 32'd471859200;
      5994: inst = 32'd136314880;
      5995: inst = 32'd268468224;
      5996: inst = 32'd201344143;
      5997: inst = 32'd203489279;
      5998: inst = 32'd471859200;
      5999: inst = 32'd136314880;
      6000: inst = 32'd268468224;
      6001: inst = 32'd201344144;
      6002: inst = 32'd203489279;
      6003: inst = 32'd471859200;
      6004: inst = 32'd136314880;
      6005: inst = 32'd268468224;
      6006: inst = 32'd201344145;
      6007: inst = 32'd203489279;
      6008: inst = 32'd471859200;
      6009: inst = 32'd136314880;
      6010: inst = 32'd268468224;
      6011: inst = 32'd201344146;
      6012: inst = 32'd203489279;
      6013: inst = 32'd471859200;
      6014: inst = 32'd136314880;
      6015: inst = 32'd268468224;
      6016: inst = 32'd201344147;
      6017: inst = 32'd203489279;
      6018: inst = 32'd471859200;
      6019: inst = 32'd136314880;
      6020: inst = 32'd268468224;
      6021: inst = 32'd201344148;
      6022: inst = 32'd203489279;
      6023: inst = 32'd471859200;
      6024: inst = 32'd136314880;
      6025: inst = 32'd268468224;
      6026: inst = 32'd201344149;
      6027: inst = 32'd203489279;
      6028: inst = 32'd471859200;
      6029: inst = 32'd136314880;
      6030: inst = 32'd268468224;
      6031: inst = 32'd201344150;
      6032: inst = 32'd203489279;
      6033: inst = 32'd471859200;
      6034: inst = 32'd136314880;
      6035: inst = 32'd268468224;
      6036: inst = 32'd201344151;
      6037: inst = 32'd203489279;
      6038: inst = 32'd471859200;
      6039: inst = 32'd136314880;
      6040: inst = 32'd268468224;
      6041: inst = 32'd201344152;
      6042: inst = 32'd203489279;
      6043: inst = 32'd471859200;
      6044: inst = 32'd136314880;
      6045: inst = 32'd268468224;
      6046: inst = 32'd201344153;
      6047: inst = 32'd203489279;
      6048: inst = 32'd471859200;
      6049: inst = 32'd136314880;
      6050: inst = 32'd268468224;
      6051: inst = 32'd201344154;
      6052: inst = 32'd203489279;
      6053: inst = 32'd471859200;
      6054: inst = 32'd136314880;
      6055: inst = 32'd268468224;
      6056: inst = 32'd201344155;
      6057: inst = 32'd203489279;
      6058: inst = 32'd471859200;
      6059: inst = 32'd136314880;
      6060: inst = 32'd268468224;
      6061: inst = 32'd201344156;
      6062: inst = 32'd203489279;
      6063: inst = 32'd471859200;
      6064: inst = 32'd136314880;
      6065: inst = 32'd268468224;
      6066: inst = 32'd201344157;
      6067: inst = 32'd203489279;
      6068: inst = 32'd471859200;
      6069: inst = 32'd136314880;
      6070: inst = 32'd268468224;
      6071: inst = 32'd201344158;
      6072: inst = 32'd203489279;
      6073: inst = 32'd471859200;
      6074: inst = 32'd136314880;
      6075: inst = 32'd268468224;
      6076: inst = 32'd201344159;
      6077: inst = 32'd203489279;
      6078: inst = 32'd471859200;
      6079: inst = 32'd136314880;
      6080: inst = 32'd268468224;
      6081: inst = 32'd201344160;
      6082: inst = 32'd203489279;
      6083: inst = 32'd471859200;
      6084: inst = 32'd136314880;
      6085: inst = 32'd268468224;
      6086: inst = 32'd201344161;
      6087: inst = 32'd203489279;
      6088: inst = 32'd471859200;
      6089: inst = 32'd136314880;
      6090: inst = 32'd268468224;
      6091: inst = 32'd201344162;
      6092: inst = 32'd203489279;
      6093: inst = 32'd471859200;
      6094: inst = 32'd136314880;
      6095: inst = 32'd268468224;
      6096: inst = 32'd201344163;
      6097: inst = 32'd203489279;
      6098: inst = 32'd471859200;
      6099: inst = 32'd136314880;
      6100: inst = 32'd268468224;
      6101: inst = 32'd201344164;
      6102: inst = 32'd203484854;
      6103: inst = 32'd471859200;
      6104: inst = 32'd136314880;
      6105: inst = 32'd268468224;
      6106: inst = 32'd201344165;
      6107: inst = 32'd203484854;
      6108: inst = 32'd471859200;
      6109: inst = 32'd136314880;
      6110: inst = 32'd268468224;
      6111: inst = 32'd201344166;
      6112: inst = 32'd203484854;
      6113: inst = 32'd471859200;
      6114: inst = 32'd136314880;
      6115: inst = 32'd268468224;
      6116: inst = 32'd201344167;
      6117: inst = 32'd203484854;
      6118: inst = 32'd471859200;
      6119: inst = 32'd136314880;
      6120: inst = 32'd268468224;
      6121: inst = 32'd201344168;
      6122: inst = 32'd203484854;
      6123: inst = 32'd471859200;
      6124: inst = 32'd136314880;
      6125: inst = 32'd268468224;
      6126: inst = 32'd201344169;
      6127: inst = 32'd203484854;
      6128: inst = 32'd471859200;
      6129: inst = 32'd136314880;
      6130: inst = 32'd268468224;
      6131: inst = 32'd201344170;
      6132: inst = 32'd203484854;
      6133: inst = 32'd471859200;
      6134: inst = 32'd136314880;
      6135: inst = 32'd268468224;
      6136: inst = 32'd201344171;
      6137: inst = 32'd203484854;
      6138: inst = 32'd471859200;
      6139: inst = 32'd136314880;
      6140: inst = 32'd268468224;
      6141: inst = 32'd201344172;
      6142: inst = 32'd203484854;
      6143: inst = 32'd471859200;
      6144: inst = 32'd136314880;
      6145: inst = 32'd268468224;
      6146: inst = 32'd201344173;
      6147: inst = 32'd203484854;
      6148: inst = 32'd471859200;
      6149: inst = 32'd136314880;
      6150: inst = 32'd268468224;
      6151: inst = 32'd201344174;
      6152: inst = 32'd203484854;
      6153: inst = 32'd471859200;
      6154: inst = 32'd136314880;
      6155: inst = 32'd268468224;
      6156: inst = 32'd201344175;
      6157: inst = 32'd203484854;
      6158: inst = 32'd471859200;
      6159: inst = 32'd136314880;
      6160: inst = 32'd268468224;
      6161: inst = 32'd201344176;
      6162: inst = 32'd203484854;
      6163: inst = 32'd471859200;
      6164: inst = 32'd136314880;
      6165: inst = 32'd268468224;
      6166: inst = 32'd201344177;
      6167: inst = 32'd203484854;
      6168: inst = 32'd471859200;
      6169: inst = 32'd136314880;
      6170: inst = 32'd268468224;
      6171: inst = 32'd201344178;
      6172: inst = 32'd203484816;
      6173: inst = 32'd471859200;
      6174: inst = 32'd136314880;
      6175: inst = 32'd268468224;
      6176: inst = 32'd201344179;
      6177: inst = 32'd203484744;
      6178: inst = 32'd471859200;
      6179: inst = 32'd136314880;
      6180: inst = 32'd268468224;
      6181: inst = 32'd201344180;
      6182: inst = 32'd203484744;
      6183: inst = 32'd471859200;
      6184: inst = 32'd136314880;
      6185: inst = 32'd268468224;
      6186: inst = 32'd201344181;
      6187: inst = 32'd203484814;
      6188: inst = 32'd471859200;
      6189: inst = 32'd136314880;
      6190: inst = 32'd268468224;
      6191: inst = 32'd201344182;
      6192: inst = 32'd203484854;
      6193: inst = 32'd471859200;
      6194: inst = 32'd136314880;
      6195: inst = 32'd268468224;
      6196: inst = 32'd201344183;
      6197: inst = 32'd203484854;
      6198: inst = 32'd471859200;
      6199: inst = 32'd136314880;
      6200: inst = 32'd268468224;
      6201: inst = 32'd201344184;
      6202: inst = 32'd203484854;
      6203: inst = 32'd471859200;
      6204: inst = 32'd136314880;
      6205: inst = 32'd268468224;
      6206: inst = 32'd201344185;
      6207: inst = 32'd203484854;
      6208: inst = 32'd471859200;
      6209: inst = 32'd136314880;
      6210: inst = 32'd268468224;
      6211: inst = 32'd201344186;
      6212: inst = 32'd203484854;
      6213: inst = 32'd471859200;
      6214: inst = 32'd136314880;
      6215: inst = 32'd268468224;
      6216: inst = 32'd201344187;
      6217: inst = 32'd203484854;
      6218: inst = 32'd471859200;
      6219: inst = 32'd136314880;
      6220: inst = 32'd268468224;
      6221: inst = 32'd201344188;
      6222: inst = 32'd203484854;
      6223: inst = 32'd471859200;
      6224: inst = 32'd136314880;
      6225: inst = 32'd268468224;
      6226: inst = 32'd201344189;
      6227: inst = 32'd203484854;
      6228: inst = 32'd471859200;
      6229: inst = 32'd136314880;
      6230: inst = 32'd268468224;
      6231: inst = 32'd201344190;
      6232: inst = 32'd203484854;
      6233: inst = 32'd471859200;
      6234: inst = 32'd136314880;
      6235: inst = 32'd268468224;
      6236: inst = 32'd201344191;
      6237: inst = 32'd203484854;
      6238: inst = 32'd471859200;
      6239: inst = 32'd136314880;
      6240: inst = 32'd268468224;
      6241: inst = 32'd201344192;
      6242: inst = 32'd203484854;
      6243: inst = 32'd471859200;
      6244: inst = 32'd136314880;
      6245: inst = 32'd268468224;
      6246: inst = 32'd201344193;
      6247: inst = 32'd203484854;
      6248: inst = 32'd471859200;
      6249: inst = 32'd136314880;
      6250: inst = 32'd268468224;
      6251: inst = 32'd201344194;
      6252: inst = 32'd203484854;
      6253: inst = 32'd471859200;
      6254: inst = 32'd136314880;
      6255: inst = 32'd268468224;
      6256: inst = 32'd201344195;
      6257: inst = 32'd203484854;
      6258: inst = 32'd471859200;
      6259: inst = 32'd136314880;
      6260: inst = 32'd268468224;
      6261: inst = 32'd201344196;
      6262: inst = 32'd203484854;
      6263: inst = 32'd471859200;
      6264: inst = 32'd136314880;
      6265: inst = 32'd268468224;
      6266: inst = 32'd201344197;
      6267: inst = 32'd203484854;
      6268: inst = 32'd471859200;
      6269: inst = 32'd136314880;
      6270: inst = 32'd268468224;
      6271: inst = 32'd201344198;
      6272: inst = 32'd203484854;
      6273: inst = 32'd471859200;
      6274: inst = 32'd136314880;
      6275: inst = 32'd268468224;
      6276: inst = 32'd201344199;
      6277: inst = 32'd203484854;
      6278: inst = 32'd471859200;
      6279: inst = 32'd136314880;
      6280: inst = 32'd268468224;
      6281: inst = 32'd201344200;
      6282: inst = 32'd203484854;
      6283: inst = 32'd471859200;
      6284: inst = 32'd136314880;
      6285: inst = 32'd268468224;
      6286: inst = 32'd201344201;
      6287: inst = 32'd203484854;
      6288: inst = 32'd471859200;
      6289: inst = 32'd136314880;
      6290: inst = 32'd268468224;
      6291: inst = 32'd201344202;
      6292: inst = 32'd203484854;
      6293: inst = 32'd471859200;
      6294: inst = 32'd136314880;
      6295: inst = 32'd268468224;
      6296: inst = 32'd201344203;
      6297: inst = 32'd203484853;
      6298: inst = 32'd471859200;
      6299: inst = 32'd136314880;
      6300: inst = 32'd268468224;
      6301: inst = 32'd201344204;
      6302: inst = 32'd203484853;
      6303: inst = 32'd471859200;
      6304: inst = 32'd136314880;
      6305: inst = 32'd268468224;
      6306: inst = 32'd201344205;
      6307: inst = 32'd203484854;
      6308: inst = 32'd471859200;
      6309: inst = 32'd136314880;
      6310: inst = 32'd268468224;
      6311: inst = 32'd201344206;
      6312: inst = 32'd203484854;
      6313: inst = 32'd471859200;
      6314: inst = 32'd136314880;
      6315: inst = 32'd268468224;
      6316: inst = 32'd201344207;
      6317: inst = 32'd203484854;
      6318: inst = 32'd471859200;
      6319: inst = 32'd136314880;
      6320: inst = 32'd268468224;
      6321: inst = 32'd201344208;
      6322: inst = 32'd203484854;
      6323: inst = 32'd471859200;
      6324: inst = 32'd136314880;
      6325: inst = 32'd268468224;
      6326: inst = 32'd201344209;
      6327: inst = 32'd203484854;
      6328: inst = 32'd471859200;
      6329: inst = 32'd136314880;
      6330: inst = 32'd268468224;
      6331: inst = 32'd201344210;
      6332: inst = 32'd203484854;
      6333: inst = 32'd471859200;
      6334: inst = 32'd136314880;
      6335: inst = 32'd268468224;
      6336: inst = 32'd201344211;
      6337: inst = 32'd203484854;
      6338: inst = 32'd471859200;
      6339: inst = 32'd136314880;
      6340: inst = 32'd268468224;
      6341: inst = 32'd201344212;
      6342: inst = 32'd203484854;
      6343: inst = 32'd471859200;
      6344: inst = 32'd136314880;
      6345: inst = 32'd268468224;
      6346: inst = 32'd201344213;
      6347: inst = 32'd203484854;
      6348: inst = 32'd471859200;
      6349: inst = 32'd136314880;
      6350: inst = 32'd268468224;
      6351: inst = 32'd201344214;
      6352: inst = 32'd203484854;
      6353: inst = 32'd471859200;
      6354: inst = 32'd136314880;
      6355: inst = 32'd268468224;
      6356: inst = 32'd201344215;
      6357: inst = 32'd203484854;
      6358: inst = 32'd471859200;
      6359: inst = 32'd136314880;
      6360: inst = 32'd268468224;
      6361: inst = 32'd201344216;
      6362: inst = 32'd203484854;
      6363: inst = 32'd471859200;
      6364: inst = 32'd136314880;
      6365: inst = 32'd268468224;
      6366: inst = 32'd201344217;
      6367: inst = 32'd203484854;
      6368: inst = 32'd471859200;
      6369: inst = 32'd136314880;
      6370: inst = 32'd268468224;
      6371: inst = 32'd201344218;
      6372: inst = 32'd203484854;
      6373: inst = 32'd471859200;
      6374: inst = 32'd136314880;
      6375: inst = 32'd268468224;
      6376: inst = 32'd201344219;
      6377: inst = 32'd203484854;
      6378: inst = 32'd471859200;
      6379: inst = 32'd136314880;
      6380: inst = 32'd268468224;
      6381: inst = 32'd201344220;
      6382: inst = 32'd203489279;
      6383: inst = 32'd471859200;
      6384: inst = 32'd136314880;
      6385: inst = 32'd268468224;
      6386: inst = 32'd201344221;
      6387: inst = 32'd203489279;
      6388: inst = 32'd471859200;
      6389: inst = 32'd136314880;
      6390: inst = 32'd268468224;
      6391: inst = 32'd201344222;
      6392: inst = 32'd203489279;
      6393: inst = 32'd471859200;
      6394: inst = 32'd136314880;
      6395: inst = 32'd268468224;
      6396: inst = 32'd201344223;
      6397: inst = 32'd203489279;
      6398: inst = 32'd471859200;
      6399: inst = 32'd136314880;
      6400: inst = 32'd268468224;
      6401: inst = 32'd201344224;
      6402: inst = 32'd203489279;
      6403: inst = 32'd471859200;
      6404: inst = 32'd136314880;
      6405: inst = 32'd268468224;
      6406: inst = 32'd201344225;
      6407: inst = 32'd203489279;
      6408: inst = 32'd471859200;
      6409: inst = 32'd136314880;
      6410: inst = 32'd268468224;
      6411: inst = 32'd201344226;
      6412: inst = 32'd203489279;
      6413: inst = 32'd471859200;
      6414: inst = 32'd136314880;
      6415: inst = 32'd268468224;
      6416: inst = 32'd201344227;
      6417: inst = 32'd203489279;
      6418: inst = 32'd471859200;
      6419: inst = 32'd136314880;
      6420: inst = 32'd268468224;
      6421: inst = 32'd201344228;
      6422: inst = 32'd203489279;
      6423: inst = 32'd471859200;
      6424: inst = 32'd136314880;
      6425: inst = 32'd268468224;
      6426: inst = 32'd201344229;
      6427: inst = 32'd203489279;
      6428: inst = 32'd471859200;
      6429: inst = 32'd136314880;
      6430: inst = 32'd268468224;
      6431: inst = 32'd201344230;
      6432: inst = 32'd203489279;
      6433: inst = 32'd471859200;
      6434: inst = 32'd136314880;
      6435: inst = 32'd268468224;
      6436: inst = 32'd201344231;
      6437: inst = 32'd203489279;
      6438: inst = 32'd471859200;
      6439: inst = 32'd136314880;
      6440: inst = 32'd268468224;
      6441: inst = 32'd201344232;
      6442: inst = 32'd203489279;
      6443: inst = 32'd471859200;
      6444: inst = 32'd136314880;
      6445: inst = 32'd268468224;
      6446: inst = 32'd201344233;
      6447: inst = 32'd203489279;
      6448: inst = 32'd471859200;
      6449: inst = 32'd136314880;
      6450: inst = 32'd268468224;
      6451: inst = 32'd201344234;
      6452: inst = 32'd203489279;
      6453: inst = 32'd471859200;
      6454: inst = 32'd136314880;
      6455: inst = 32'd268468224;
      6456: inst = 32'd201344235;
      6457: inst = 32'd203489279;
      6458: inst = 32'd471859200;
      6459: inst = 32'd136314880;
      6460: inst = 32'd268468224;
      6461: inst = 32'd201344236;
      6462: inst = 32'd203489279;
      6463: inst = 32'd471859200;
      6464: inst = 32'd136314880;
      6465: inst = 32'd268468224;
      6466: inst = 32'd201344237;
      6467: inst = 32'd203489279;
      6468: inst = 32'd471859200;
      6469: inst = 32'd136314880;
      6470: inst = 32'd268468224;
      6471: inst = 32'd201344238;
      6472: inst = 32'd203489279;
      6473: inst = 32'd471859200;
      6474: inst = 32'd136314880;
      6475: inst = 32'd268468224;
      6476: inst = 32'd201344239;
      6477: inst = 32'd203489279;
      6478: inst = 32'd471859200;
      6479: inst = 32'd136314880;
      6480: inst = 32'd268468224;
      6481: inst = 32'd201344240;
      6482: inst = 32'd203489279;
      6483: inst = 32'd471859200;
      6484: inst = 32'd136314880;
      6485: inst = 32'd268468224;
      6486: inst = 32'd201344241;
      6487: inst = 32'd203489279;
      6488: inst = 32'd471859200;
      6489: inst = 32'd136314880;
      6490: inst = 32'd268468224;
      6491: inst = 32'd201344242;
      6492: inst = 32'd203489279;
      6493: inst = 32'd471859200;
      6494: inst = 32'd136314880;
      6495: inst = 32'd268468224;
      6496: inst = 32'd201344243;
      6497: inst = 32'd203489279;
      6498: inst = 32'd471859200;
      6499: inst = 32'd136314880;
      6500: inst = 32'd268468224;
      6501: inst = 32'd201344244;
      6502: inst = 32'd203489279;
      6503: inst = 32'd471859200;
      6504: inst = 32'd136314880;
      6505: inst = 32'd268468224;
      6506: inst = 32'd201344245;
      6507: inst = 32'd203489279;
      6508: inst = 32'd471859200;
      6509: inst = 32'd136314880;
      6510: inst = 32'd268468224;
      6511: inst = 32'd201344246;
      6512: inst = 32'd203489279;
      6513: inst = 32'd471859200;
      6514: inst = 32'd136314880;
      6515: inst = 32'd268468224;
      6516: inst = 32'd201344247;
      6517: inst = 32'd203489279;
      6518: inst = 32'd471859200;
      6519: inst = 32'd136314880;
      6520: inst = 32'd268468224;
      6521: inst = 32'd201344248;
      6522: inst = 32'd203489279;
      6523: inst = 32'd471859200;
      6524: inst = 32'd136314880;
      6525: inst = 32'd268468224;
      6526: inst = 32'd201344249;
      6527: inst = 32'd203489279;
      6528: inst = 32'd471859200;
      6529: inst = 32'd136314880;
      6530: inst = 32'd268468224;
      6531: inst = 32'd201344250;
      6532: inst = 32'd203489279;
      6533: inst = 32'd471859200;
      6534: inst = 32'd136314880;
      6535: inst = 32'd268468224;
      6536: inst = 32'd201344251;
      6537: inst = 32'd203489279;
      6538: inst = 32'd471859200;
      6539: inst = 32'd136314880;
      6540: inst = 32'd268468224;
      6541: inst = 32'd201344252;
      6542: inst = 32'd203489279;
      6543: inst = 32'd471859200;
      6544: inst = 32'd136314880;
      6545: inst = 32'd268468224;
      6546: inst = 32'd201344253;
      6547: inst = 32'd203489279;
      6548: inst = 32'd471859200;
      6549: inst = 32'd136314880;
      6550: inst = 32'd268468224;
      6551: inst = 32'd201344254;
      6552: inst = 32'd203489279;
      6553: inst = 32'd471859200;
      6554: inst = 32'd136314880;
      6555: inst = 32'd268468224;
      6556: inst = 32'd201344255;
      6557: inst = 32'd203489279;
      6558: inst = 32'd471859200;
      6559: inst = 32'd136314880;
      6560: inst = 32'd268468224;
      6561: inst = 32'd201344256;
      6562: inst = 32'd203489279;
      6563: inst = 32'd471859200;
      6564: inst = 32'd136314880;
      6565: inst = 32'd268468224;
      6566: inst = 32'd201344257;
      6567: inst = 32'd203489279;
      6568: inst = 32'd471859200;
      6569: inst = 32'd136314880;
      6570: inst = 32'd268468224;
      6571: inst = 32'd201344258;
      6572: inst = 32'd203489279;
      6573: inst = 32'd471859200;
      6574: inst = 32'd136314880;
      6575: inst = 32'd268468224;
      6576: inst = 32'd201344259;
      6577: inst = 32'd203489279;
      6578: inst = 32'd471859200;
      6579: inst = 32'd136314880;
      6580: inst = 32'd268468224;
      6581: inst = 32'd201344260;
      6582: inst = 32'd203484854;
      6583: inst = 32'd471859200;
      6584: inst = 32'd136314880;
      6585: inst = 32'd268468224;
      6586: inst = 32'd201344261;
      6587: inst = 32'd203484854;
      6588: inst = 32'd471859200;
      6589: inst = 32'd136314880;
      6590: inst = 32'd268468224;
      6591: inst = 32'd201344262;
      6592: inst = 32'd203484854;
      6593: inst = 32'd471859200;
      6594: inst = 32'd136314880;
      6595: inst = 32'd268468224;
      6596: inst = 32'd201344263;
      6597: inst = 32'd203484854;
      6598: inst = 32'd471859200;
      6599: inst = 32'd136314880;
      6600: inst = 32'd268468224;
      6601: inst = 32'd201344264;
      6602: inst = 32'd203484854;
      6603: inst = 32'd471859200;
      6604: inst = 32'd136314880;
      6605: inst = 32'd268468224;
      6606: inst = 32'd201344265;
      6607: inst = 32'd203484854;
      6608: inst = 32'd471859200;
      6609: inst = 32'd136314880;
      6610: inst = 32'd268468224;
      6611: inst = 32'd201344266;
      6612: inst = 32'd203484854;
      6613: inst = 32'd471859200;
      6614: inst = 32'd136314880;
      6615: inst = 32'd268468224;
      6616: inst = 32'd201344267;
      6617: inst = 32'd203484854;
      6618: inst = 32'd471859200;
      6619: inst = 32'd136314880;
      6620: inst = 32'd268468224;
      6621: inst = 32'd201344268;
      6622: inst = 32'd203484854;
      6623: inst = 32'd471859200;
      6624: inst = 32'd136314880;
      6625: inst = 32'd268468224;
      6626: inst = 32'd201344269;
      6627: inst = 32'd203484854;
      6628: inst = 32'd471859200;
      6629: inst = 32'd136314880;
      6630: inst = 32'd268468224;
      6631: inst = 32'd201344270;
      6632: inst = 32'd203484854;
      6633: inst = 32'd471859200;
      6634: inst = 32'd136314880;
      6635: inst = 32'd268468224;
      6636: inst = 32'd201344271;
      6637: inst = 32'd203484854;
      6638: inst = 32'd471859200;
      6639: inst = 32'd136314880;
      6640: inst = 32'd268468224;
      6641: inst = 32'd201344272;
      6642: inst = 32'd203484854;
      6643: inst = 32'd471859200;
      6644: inst = 32'd136314880;
      6645: inst = 32'd268468224;
      6646: inst = 32'd201344273;
      6647: inst = 32'd203484854;
      6648: inst = 32'd471859200;
      6649: inst = 32'd136314880;
      6650: inst = 32'd268468224;
      6651: inst = 32'd201344274;
      6652: inst = 32'd203484854;
      6653: inst = 32'd471859200;
      6654: inst = 32'd136314880;
      6655: inst = 32'd268468224;
      6656: inst = 32'd201344275;
      6657: inst = 32'd203484853;
      6658: inst = 32'd471859200;
      6659: inst = 32'd136314880;
      6660: inst = 32'd268468224;
      6661: inst = 32'd201344276;
      6662: inst = 32'd203484853;
      6663: inst = 32'd471859200;
      6664: inst = 32'd136314880;
      6665: inst = 32'd268468224;
      6666: inst = 32'd201344277;
      6667: inst = 32'd203484854;
      6668: inst = 32'd471859200;
      6669: inst = 32'd136314880;
      6670: inst = 32'd268468224;
      6671: inst = 32'd201344278;
      6672: inst = 32'd203484854;
      6673: inst = 32'd471859200;
      6674: inst = 32'd136314880;
      6675: inst = 32'd268468224;
      6676: inst = 32'd201344279;
      6677: inst = 32'd203484854;
      6678: inst = 32'd471859200;
      6679: inst = 32'd136314880;
      6680: inst = 32'd268468224;
      6681: inst = 32'd201344280;
      6682: inst = 32'd203484854;
      6683: inst = 32'd471859200;
      6684: inst = 32'd136314880;
      6685: inst = 32'd268468224;
      6686: inst = 32'd201344281;
      6687: inst = 32'd203484854;
      6688: inst = 32'd471859200;
      6689: inst = 32'd136314880;
      6690: inst = 32'd268468224;
      6691: inst = 32'd201344282;
      6692: inst = 32'd203484854;
      6693: inst = 32'd471859200;
      6694: inst = 32'd136314880;
      6695: inst = 32'd268468224;
      6696: inst = 32'd201344283;
      6697: inst = 32'd203484854;
      6698: inst = 32'd471859200;
      6699: inst = 32'd136314880;
      6700: inst = 32'd268468224;
      6701: inst = 32'd201344284;
      6702: inst = 32'd203484854;
      6703: inst = 32'd471859200;
      6704: inst = 32'd136314880;
      6705: inst = 32'd268468224;
      6706: inst = 32'd201344285;
      6707: inst = 32'd203484854;
      6708: inst = 32'd471859200;
      6709: inst = 32'd136314880;
      6710: inst = 32'd268468224;
      6711: inst = 32'd201344286;
      6712: inst = 32'd203484854;
      6713: inst = 32'd471859200;
      6714: inst = 32'd136314880;
      6715: inst = 32'd268468224;
      6716: inst = 32'd201344287;
      6717: inst = 32'd203484854;
      6718: inst = 32'd471859200;
      6719: inst = 32'd136314880;
      6720: inst = 32'd268468224;
      6721: inst = 32'd201344288;
      6722: inst = 32'd203484854;
      6723: inst = 32'd471859200;
      6724: inst = 32'd136314880;
      6725: inst = 32'd268468224;
      6726: inst = 32'd201344289;
      6727: inst = 32'd203484854;
      6728: inst = 32'd471859200;
      6729: inst = 32'd136314880;
      6730: inst = 32'd268468224;
      6731: inst = 32'd201344290;
      6732: inst = 32'd203484854;
      6733: inst = 32'd471859200;
      6734: inst = 32'd136314880;
      6735: inst = 32'd268468224;
      6736: inst = 32'd201344291;
      6737: inst = 32'd203484854;
      6738: inst = 32'd471859200;
      6739: inst = 32'd136314880;
      6740: inst = 32'd268468224;
      6741: inst = 32'd201344292;
      6742: inst = 32'd203484854;
      6743: inst = 32'd471859200;
      6744: inst = 32'd136314880;
      6745: inst = 32'd268468224;
      6746: inst = 32'd201344293;
      6747: inst = 32'd203484854;
      6748: inst = 32'd471859200;
      6749: inst = 32'd136314880;
      6750: inst = 32'd268468224;
      6751: inst = 32'd201344294;
      6752: inst = 32'd203484854;
      6753: inst = 32'd471859200;
      6754: inst = 32'd136314880;
      6755: inst = 32'd268468224;
      6756: inst = 32'd201344295;
      6757: inst = 32'd203484854;
      6758: inst = 32'd471859200;
      6759: inst = 32'd136314880;
      6760: inst = 32'd268468224;
      6761: inst = 32'd201344296;
      6762: inst = 32'd203484854;
      6763: inst = 32'd471859200;
      6764: inst = 32'd136314880;
      6765: inst = 32'd268468224;
      6766: inst = 32'd201344297;
      6767: inst = 32'd203484854;
      6768: inst = 32'd471859200;
      6769: inst = 32'd136314880;
      6770: inst = 32'd268468224;
      6771: inst = 32'd201344298;
      6772: inst = 32'd203484854;
      6773: inst = 32'd471859200;
      6774: inst = 32'd136314880;
      6775: inst = 32'd268468224;
      6776: inst = 32'd201344299;
      6777: inst = 32'd203484854;
      6778: inst = 32'd471859200;
      6779: inst = 32'd136314880;
      6780: inst = 32'd268468224;
      6781: inst = 32'd201344300;
      6782: inst = 32'd203484854;
      6783: inst = 32'd471859200;
      6784: inst = 32'd136314880;
      6785: inst = 32'd268468224;
      6786: inst = 32'd201344301;
      6787: inst = 32'd203484854;
      6788: inst = 32'd471859200;
      6789: inst = 32'd136314880;
      6790: inst = 32'd268468224;
      6791: inst = 32'd201344302;
      6792: inst = 32'd203484854;
      6793: inst = 32'd471859200;
      6794: inst = 32'd136314880;
      6795: inst = 32'd268468224;
      6796: inst = 32'd201344303;
      6797: inst = 32'd203484854;
      6798: inst = 32'd471859200;
      6799: inst = 32'd136314880;
      6800: inst = 32'd268468224;
      6801: inst = 32'd201344304;
      6802: inst = 32'd203484854;
      6803: inst = 32'd471859200;
      6804: inst = 32'd136314880;
      6805: inst = 32'd268468224;
      6806: inst = 32'd201344305;
      6807: inst = 32'd203484854;
      6808: inst = 32'd471859200;
      6809: inst = 32'd136314880;
      6810: inst = 32'd268468224;
      6811: inst = 32'd201344306;
      6812: inst = 32'd203484854;
      6813: inst = 32'd471859200;
      6814: inst = 32'd136314880;
      6815: inst = 32'd268468224;
      6816: inst = 32'd201344307;
      6817: inst = 32'd203484854;
      6818: inst = 32'd471859200;
      6819: inst = 32'd136314880;
      6820: inst = 32'd268468224;
      6821: inst = 32'd201344308;
      6822: inst = 32'd203484854;
      6823: inst = 32'd471859200;
      6824: inst = 32'd136314880;
      6825: inst = 32'd268468224;
      6826: inst = 32'd201344309;
      6827: inst = 32'd203484854;
      6828: inst = 32'd471859200;
      6829: inst = 32'd136314880;
      6830: inst = 32'd268468224;
      6831: inst = 32'd201344310;
      6832: inst = 32'd203484854;
      6833: inst = 32'd471859200;
      6834: inst = 32'd136314880;
      6835: inst = 32'd268468224;
      6836: inst = 32'd201344311;
      6837: inst = 32'd203484854;
      6838: inst = 32'd471859200;
      6839: inst = 32'd136314880;
      6840: inst = 32'd268468224;
      6841: inst = 32'd201344312;
      6842: inst = 32'd203484854;
      6843: inst = 32'd471859200;
      6844: inst = 32'd136314880;
      6845: inst = 32'd268468224;
      6846: inst = 32'd201344313;
      6847: inst = 32'd203484854;
      6848: inst = 32'd471859200;
      6849: inst = 32'd136314880;
      6850: inst = 32'd268468224;
      6851: inst = 32'd201344314;
      6852: inst = 32'd203484854;
      6853: inst = 32'd471859200;
      6854: inst = 32'd136314880;
      6855: inst = 32'd268468224;
      6856: inst = 32'd201344315;
      6857: inst = 32'd203484854;
      6858: inst = 32'd471859200;
      6859: inst = 32'd136314880;
      6860: inst = 32'd268468224;
      6861: inst = 32'd201344316;
      6862: inst = 32'd203489279;
      6863: inst = 32'd471859200;
      6864: inst = 32'd136314880;
      6865: inst = 32'd268468224;
      6866: inst = 32'd201344317;
      6867: inst = 32'd203489279;
      6868: inst = 32'd471859200;
      6869: inst = 32'd136314880;
      6870: inst = 32'd268468224;
      6871: inst = 32'd201344318;
      6872: inst = 32'd203489279;
      6873: inst = 32'd471859200;
      6874: inst = 32'd136314880;
      6875: inst = 32'd268468224;
      6876: inst = 32'd201344319;
      6877: inst = 32'd203489279;
      6878: inst = 32'd471859200;
      6879: inst = 32'd136314880;
      6880: inst = 32'd268468224;
      6881: inst = 32'd201344320;
      6882: inst = 32'd203489279;
      6883: inst = 32'd471859200;
      6884: inst = 32'd136314880;
      6885: inst = 32'd268468224;
      6886: inst = 32'd201344321;
      6887: inst = 32'd203489279;
      6888: inst = 32'd471859200;
      6889: inst = 32'd136314880;
      6890: inst = 32'd268468224;
      6891: inst = 32'd201344322;
      6892: inst = 32'd203489279;
      6893: inst = 32'd471859200;
      6894: inst = 32'd136314880;
      6895: inst = 32'd268468224;
      6896: inst = 32'd201344323;
      6897: inst = 32'd203489279;
      6898: inst = 32'd471859200;
      6899: inst = 32'd136314880;
      6900: inst = 32'd268468224;
      6901: inst = 32'd201344324;
      6902: inst = 32'd203489279;
      6903: inst = 32'd471859200;
      6904: inst = 32'd136314880;
      6905: inst = 32'd268468224;
      6906: inst = 32'd201344325;
      6907: inst = 32'd203489279;
      6908: inst = 32'd471859200;
      6909: inst = 32'd136314880;
      6910: inst = 32'd268468224;
      6911: inst = 32'd201344326;
      6912: inst = 32'd203489279;
      6913: inst = 32'd471859200;
      6914: inst = 32'd136314880;
      6915: inst = 32'd268468224;
      6916: inst = 32'd201344327;
      6917: inst = 32'd203489279;
      6918: inst = 32'd471859200;
      6919: inst = 32'd136314880;
      6920: inst = 32'd268468224;
      6921: inst = 32'd201344328;
      6922: inst = 32'd203489279;
      6923: inst = 32'd471859200;
      6924: inst = 32'd136314880;
      6925: inst = 32'd268468224;
      6926: inst = 32'd201344329;
      6927: inst = 32'd203489279;
      6928: inst = 32'd471859200;
      6929: inst = 32'd136314880;
      6930: inst = 32'd268468224;
      6931: inst = 32'd201344330;
      6932: inst = 32'd203489279;
      6933: inst = 32'd471859200;
      6934: inst = 32'd136314880;
      6935: inst = 32'd268468224;
      6936: inst = 32'd201344331;
      6937: inst = 32'd203489279;
      6938: inst = 32'd471859200;
      6939: inst = 32'd136314880;
      6940: inst = 32'd268468224;
      6941: inst = 32'd201344332;
      6942: inst = 32'd203489279;
      6943: inst = 32'd471859200;
      6944: inst = 32'd136314880;
      6945: inst = 32'd268468224;
      6946: inst = 32'd201344333;
      6947: inst = 32'd203489279;
      6948: inst = 32'd471859200;
      6949: inst = 32'd136314880;
      6950: inst = 32'd268468224;
      6951: inst = 32'd201344334;
      6952: inst = 32'd203489279;
      6953: inst = 32'd471859200;
      6954: inst = 32'd136314880;
      6955: inst = 32'd268468224;
      6956: inst = 32'd201344335;
      6957: inst = 32'd203489279;
      6958: inst = 32'd471859200;
      6959: inst = 32'd136314880;
      6960: inst = 32'd268468224;
      6961: inst = 32'd201344336;
      6962: inst = 32'd203489279;
      6963: inst = 32'd471859200;
      6964: inst = 32'd136314880;
      6965: inst = 32'd268468224;
      6966: inst = 32'd201344337;
      6967: inst = 32'd203489279;
      6968: inst = 32'd471859200;
      6969: inst = 32'd136314880;
      6970: inst = 32'd268468224;
      6971: inst = 32'd201344338;
      6972: inst = 32'd203489279;
      6973: inst = 32'd471859200;
      6974: inst = 32'd136314880;
      6975: inst = 32'd268468224;
      6976: inst = 32'd201344339;
      6977: inst = 32'd203489279;
      6978: inst = 32'd471859200;
      6979: inst = 32'd136314880;
      6980: inst = 32'd268468224;
      6981: inst = 32'd201344340;
      6982: inst = 32'd203489279;
      6983: inst = 32'd471859200;
      6984: inst = 32'd136314880;
      6985: inst = 32'd268468224;
      6986: inst = 32'd201344341;
      6987: inst = 32'd203489279;
      6988: inst = 32'd471859200;
      6989: inst = 32'd136314880;
      6990: inst = 32'd268468224;
      6991: inst = 32'd201344342;
      6992: inst = 32'd203489279;
      6993: inst = 32'd471859200;
      6994: inst = 32'd136314880;
      6995: inst = 32'd268468224;
      6996: inst = 32'd201344343;
      6997: inst = 32'd203489279;
      6998: inst = 32'd471859200;
      6999: inst = 32'd136314880;
      7000: inst = 32'd268468224;
      7001: inst = 32'd201344344;
      7002: inst = 32'd203489279;
      7003: inst = 32'd471859200;
      7004: inst = 32'd136314880;
      7005: inst = 32'd268468224;
      7006: inst = 32'd201344345;
      7007: inst = 32'd203489279;
      7008: inst = 32'd471859200;
      7009: inst = 32'd136314880;
      7010: inst = 32'd268468224;
      7011: inst = 32'd201344346;
      7012: inst = 32'd203489279;
      7013: inst = 32'd471859200;
      7014: inst = 32'd136314880;
      7015: inst = 32'd268468224;
      7016: inst = 32'd201344347;
      7017: inst = 32'd203489279;
      7018: inst = 32'd471859200;
      7019: inst = 32'd136314880;
      7020: inst = 32'd268468224;
      7021: inst = 32'd201344348;
      7022: inst = 32'd203489279;
      7023: inst = 32'd471859200;
      7024: inst = 32'd136314880;
      7025: inst = 32'd268468224;
      7026: inst = 32'd201344349;
      7027: inst = 32'd203489279;
      7028: inst = 32'd471859200;
      7029: inst = 32'd136314880;
      7030: inst = 32'd268468224;
      7031: inst = 32'd201344350;
      7032: inst = 32'd203489279;
      7033: inst = 32'd471859200;
      7034: inst = 32'd136314880;
      7035: inst = 32'd268468224;
      7036: inst = 32'd201344351;
      7037: inst = 32'd203489279;
      7038: inst = 32'd471859200;
      7039: inst = 32'd136314880;
      7040: inst = 32'd268468224;
      7041: inst = 32'd201344352;
      7042: inst = 32'd203489279;
      7043: inst = 32'd471859200;
      7044: inst = 32'd136314880;
      7045: inst = 32'd268468224;
      7046: inst = 32'd201344353;
      7047: inst = 32'd203489279;
      7048: inst = 32'd471859200;
      7049: inst = 32'd136314880;
      7050: inst = 32'd268468224;
      7051: inst = 32'd201344354;
      7052: inst = 32'd203489279;
      7053: inst = 32'd471859200;
      7054: inst = 32'd136314880;
      7055: inst = 32'd268468224;
      7056: inst = 32'd201344355;
      7057: inst = 32'd203489279;
      7058: inst = 32'd471859200;
      7059: inst = 32'd136314880;
      7060: inst = 32'd268468224;
      7061: inst = 32'd201344356;
      7062: inst = 32'd203484854;
      7063: inst = 32'd471859200;
      7064: inst = 32'd136314880;
      7065: inst = 32'd268468224;
      7066: inst = 32'd201344357;
      7067: inst = 32'd203484854;
      7068: inst = 32'd471859200;
      7069: inst = 32'd136314880;
      7070: inst = 32'd268468224;
      7071: inst = 32'd201344358;
      7072: inst = 32'd203484854;
      7073: inst = 32'd471859200;
      7074: inst = 32'd136314880;
      7075: inst = 32'd268468224;
      7076: inst = 32'd201344359;
      7077: inst = 32'd203484854;
      7078: inst = 32'd471859200;
      7079: inst = 32'd136314880;
      7080: inst = 32'd268468224;
      7081: inst = 32'd201344360;
      7082: inst = 32'd203484854;
      7083: inst = 32'd471859200;
      7084: inst = 32'd136314880;
      7085: inst = 32'd268468224;
      7086: inst = 32'd201344361;
      7087: inst = 32'd203484854;
      7088: inst = 32'd471859200;
      7089: inst = 32'd136314880;
      7090: inst = 32'd268468224;
      7091: inst = 32'd201344362;
      7092: inst = 32'd203484854;
      7093: inst = 32'd471859200;
      7094: inst = 32'd136314880;
      7095: inst = 32'd268468224;
      7096: inst = 32'd201344363;
      7097: inst = 32'd203484854;
      7098: inst = 32'd471859200;
      7099: inst = 32'd136314880;
      7100: inst = 32'd268468224;
      7101: inst = 32'd201344364;
      7102: inst = 32'd203484854;
      7103: inst = 32'd471859200;
      7104: inst = 32'd136314880;
      7105: inst = 32'd268468224;
      7106: inst = 32'd201344365;
      7107: inst = 32'd203484854;
      7108: inst = 32'd471859200;
      7109: inst = 32'd136314880;
      7110: inst = 32'd268468224;
      7111: inst = 32'd201344366;
      7112: inst = 32'd203484854;
      7113: inst = 32'd471859200;
      7114: inst = 32'd136314880;
      7115: inst = 32'd268468224;
      7116: inst = 32'd201344367;
      7117: inst = 32'd203484854;
      7118: inst = 32'd471859200;
      7119: inst = 32'd136314880;
      7120: inst = 32'd268468224;
      7121: inst = 32'd201344368;
      7122: inst = 32'd203484854;
      7123: inst = 32'd471859200;
      7124: inst = 32'd136314880;
      7125: inst = 32'd268468224;
      7126: inst = 32'd201344369;
      7127: inst = 32'd203484854;
      7128: inst = 32'd471859200;
      7129: inst = 32'd136314880;
      7130: inst = 32'd268468224;
      7131: inst = 32'd201344370;
      7132: inst = 32'd203484854;
      7133: inst = 32'd471859200;
      7134: inst = 32'd136314880;
      7135: inst = 32'd268468224;
      7136: inst = 32'd201344371;
      7137: inst = 32'd203484854;
      7138: inst = 32'd471859200;
      7139: inst = 32'd136314880;
      7140: inst = 32'd268468224;
      7141: inst = 32'd201344372;
      7142: inst = 32'd203484854;
      7143: inst = 32'd471859200;
      7144: inst = 32'd136314880;
      7145: inst = 32'd268468224;
      7146: inst = 32'd201344373;
      7147: inst = 32'd203484854;
      7148: inst = 32'd471859200;
      7149: inst = 32'd136314880;
      7150: inst = 32'd268468224;
      7151: inst = 32'd201344374;
      7152: inst = 32'd203484854;
      7153: inst = 32'd471859200;
      7154: inst = 32'd136314880;
      7155: inst = 32'd268468224;
      7156: inst = 32'd201344375;
      7157: inst = 32'd203484854;
      7158: inst = 32'd471859200;
      7159: inst = 32'd136314880;
      7160: inst = 32'd268468224;
      7161: inst = 32'd201344376;
      7162: inst = 32'd203484854;
      7163: inst = 32'd471859200;
      7164: inst = 32'd136314880;
      7165: inst = 32'd268468224;
      7166: inst = 32'd201344377;
      7167: inst = 32'd203484854;
      7168: inst = 32'd471859200;
      7169: inst = 32'd136314880;
      7170: inst = 32'd268468224;
      7171: inst = 32'd201344378;
      7172: inst = 32'd203484854;
      7173: inst = 32'd471859200;
      7174: inst = 32'd136314880;
      7175: inst = 32'd268468224;
      7176: inst = 32'd201344379;
      7177: inst = 32'd203484854;
      7178: inst = 32'd471859200;
      7179: inst = 32'd136314880;
      7180: inst = 32'd268468224;
      7181: inst = 32'd201344380;
      7182: inst = 32'd203484854;
      7183: inst = 32'd471859200;
      7184: inst = 32'd136314880;
      7185: inst = 32'd268468224;
      7186: inst = 32'd201344381;
      7187: inst = 32'd203484854;
      7188: inst = 32'd471859200;
      7189: inst = 32'd136314880;
      7190: inst = 32'd268468224;
      7191: inst = 32'd201344382;
      7192: inst = 32'd203484854;
      7193: inst = 32'd471859200;
      7194: inst = 32'd136314880;
      7195: inst = 32'd268468224;
      7196: inst = 32'd201344383;
      7197: inst = 32'd203484854;
      7198: inst = 32'd471859200;
      7199: inst = 32'd136314880;
      7200: inst = 32'd268468224;
      7201: inst = 32'd201344384;
      7202: inst = 32'd203484854;
      7203: inst = 32'd471859200;
      7204: inst = 32'd136314880;
      7205: inst = 32'd268468224;
      7206: inst = 32'd201344385;
      7207: inst = 32'd203484854;
      7208: inst = 32'd471859200;
      7209: inst = 32'd136314880;
      7210: inst = 32'd268468224;
      7211: inst = 32'd201344386;
      7212: inst = 32'd203484854;
      7213: inst = 32'd471859200;
      7214: inst = 32'd136314880;
      7215: inst = 32'd268468224;
      7216: inst = 32'd201344387;
      7217: inst = 32'd203484854;
      7218: inst = 32'd471859200;
      7219: inst = 32'd136314880;
      7220: inst = 32'd268468224;
      7221: inst = 32'd201344388;
      7222: inst = 32'd203484854;
      7223: inst = 32'd471859200;
      7224: inst = 32'd136314880;
      7225: inst = 32'd268468224;
      7226: inst = 32'd201344389;
      7227: inst = 32'd203484854;
      7228: inst = 32'd471859200;
      7229: inst = 32'd136314880;
      7230: inst = 32'd268468224;
      7231: inst = 32'd201344390;
      7232: inst = 32'd203484854;
      7233: inst = 32'd471859200;
      7234: inst = 32'd136314880;
      7235: inst = 32'd268468224;
      7236: inst = 32'd201344391;
      7237: inst = 32'd203484854;
      7238: inst = 32'd471859200;
      7239: inst = 32'd136314880;
      7240: inst = 32'd268468224;
      7241: inst = 32'd201344392;
      7242: inst = 32'd203484854;
      7243: inst = 32'd471859200;
      7244: inst = 32'd136314880;
      7245: inst = 32'd268468224;
      7246: inst = 32'd201344393;
      7247: inst = 32'd203484854;
      7248: inst = 32'd471859200;
      7249: inst = 32'd136314880;
      7250: inst = 32'd268468224;
      7251: inst = 32'd201344394;
      7252: inst = 32'd203484854;
      7253: inst = 32'd471859200;
      7254: inst = 32'd136314880;
      7255: inst = 32'd268468224;
      7256: inst = 32'd201344395;
      7257: inst = 32'd203484854;
      7258: inst = 32'd471859200;
      7259: inst = 32'd136314880;
      7260: inst = 32'd268468224;
      7261: inst = 32'd201344396;
      7262: inst = 32'd203484854;
      7263: inst = 32'd471859200;
      7264: inst = 32'd136314880;
      7265: inst = 32'd268468224;
      7266: inst = 32'd201344397;
      7267: inst = 32'd203484854;
      7268: inst = 32'd471859200;
      7269: inst = 32'd136314880;
      7270: inst = 32'd268468224;
      7271: inst = 32'd201344398;
      7272: inst = 32'd203484854;
      7273: inst = 32'd471859200;
      7274: inst = 32'd136314880;
      7275: inst = 32'd268468224;
      7276: inst = 32'd201344399;
      7277: inst = 32'd203484854;
      7278: inst = 32'd471859200;
      7279: inst = 32'd136314880;
      7280: inst = 32'd268468224;
      7281: inst = 32'd201344400;
      7282: inst = 32'd203484854;
      7283: inst = 32'd471859200;
      7284: inst = 32'd136314880;
      7285: inst = 32'd268468224;
      7286: inst = 32'd201344401;
      7287: inst = 32'd203484854;
      7288: inst = 32'd471859200;
      7289: inst = 32'd136314880;
      7290: inst = 32'd268468224;
      7291: inst = 32'd201344402;
      7292: inst = 32'd203484854;
      7293: inst = 32'd471859200;
      7294: inst = 32'd136314880;
      7295: inst = 32'd268468224;
      7296: inst = 32'd201344403;
      7297: inst = 32'd203484854;
      7298: inst = 32'd471859200;
      7299: inst = 32'd136314880;
      7300: inst = 32'd268468224;
      7301: inst = 32'd201344404;
      7302: inst = 32'd203484854;
      7303: inst = 32'd471859200;
      7304: inst = 32'd136314880;
      7305: inst = 32'd268468224;
      7306: inst = 32'd201344405;
      7307: inst = 32'd203484854;
      7308: inst = 32'd471859200;
      7309: inst = 32'd136314880;
      7310: inst = 32'd268468224;
      7311: inst = 32'd201344406;
      7312: inst = 32'd203484854;
      7313: inst = 32'd471859200;
      7314: inst = 32'd136314880;
      7315: inst = 32'd268468224;
      7316: inst = 32'd201344407;
      7317: inst = 32'd203484854;
      7318: inst = 32'd471859200;
      7319: inst = 32'd136314880;
      7320: inst = 32'd268468224;
      7321: inst = 32'd201344408;
      7322: inst = 32'd203484854;
      7323: inst = 32'd471859200;
      7324: inst = 32'd136314880;
      7325: inst = 32'd268468224;
      7326: inst = 32'd201344409;
      7327: inst = 32'd203484854;
      7328: inst = 32'd471859200;
      7329: inst = 32'd136314880;
      7330: inst = 32'd268468224;
      7331: inst = 32'd201344410;
      7332: inst = 32'd203484854;
      7333: inst = 32'd471859200;
      7334: inst = 32'd136314880;
      7335: inst = 32'd268468224;
      7336: inst = 32'd201344411;
      7337: inst = 32'd203484854;
      7338: inst = 32'd471859200;
      7339: inst = 32'd136314880;
      7340: inst = 32'd268468224;
      7341: inst = 32'd201344412;
      7342: inst = 32'd203489279;
      7343: inst = 32'd471859200;
      7344: inst = 32'd136314880;
      7345: inst = 32'd268468224;
      7346: inst = 32'd201344413;
      7347: inst = 32'd203489279;
      7348: inst = 32'd471859200;
      7349: inst = 32'd136314880;
      7350: inst = 32'd268468224;
      7351: inst = 32'd201344414;
      7352: inst = 32'd203489279;
      7353: inst = 32'd471859200;
      7354: inst = 32'd136314880;
      7355: inst = 32'd268468224;
      7356: inst = 32'd201344415;
      7357: inst = 32'd203489279;
      7358: inst = 32'd471859200;
      7359: inst = 32'd136314880;
      7360: inst = 32'd268468224;
      7361: inst = 32'd201344416;
      7362: inst = 32'd203489279;
      7363: inst = 32'd471859200;
      7364: inst = 32'd136314880;
      7365: inst = 32'd268468224;
      7366: inst = 32'd201344417;
      7367: inst = 32'd203489279;
      7368: inst = 32'd471859200;
      7369: inst = 32'd136314880;
      7370: inst = 32'd268468224;
      7371: inst = 32'd201344418;
      7372: inst = 32'd203489279;
      7373: inst = 32'd471859200;
      7374: inst = 32'd136314880;
      7375: inst = 32'd268468224;
      7376: inst = 32'd201344419;
      7377: inst = 32'd203489279;
      7378: inst = 32'd471859200;
      7379: inst = 32'd136314880;
      7380: inst = 32'd268468224;
      7381: inst = 32'd201344420;
      7382: inst = 32'd203489279;
      7383: inst = 32'd471859200;
      7384: inst = 32'd136314880;
      7385: inst = 32'd268468224;
      7386: inst = 32'd201344421;
      7387: inst = 32'd203489279;
      7388: inst = 32'd471859200;
      7389: inst = 32'd136314880;
      7390: inst = 32'd268468224;
      7391: inst = 32'd201344422;
      7392: inst = 32'd203489279;
      7393: inst = 32'd471859200;
      7394: inst = 32'd136314880;
      7395: inst = 32'd268468224;
      7396: inst = 32'd201344423;
      7397: inst = 32'd203489279;
      7398: inst = 32'd471859200;
      7399: inst = 32'd136314880;
      7400: inst = 32'd268468224;
      7401: inst = 32'd201344424;
      7402: inst = 32'd203489279;
      7403: inst = 32'd471859200;
      7404: inst = 32'd136314880;
      7405: inst = 32'd268468224;
      7406: inst = 32'd201344425;
      7407: inst = 32'd203489279;
      7408: inst = 32'd471859200;
      7409: inst = 32'd136314880;
      7410: inst = 32'd268468224;
      7411: inst = 32'd201344426;
      7412: inst = 32'd203489279;
      7413: inst = 32'd471859200;
      7414: inst = 32'd136314880;
      7415: inst = 32'd268468224;
      7416: inst = 32'd201344427;
      7417: inst = 32'd203489279;
      7418: inst = 32'd471859200;
      7419: inst = 32'd136314880;
      7420: inst = 32'd268468224;
      7421: inst = 32'd201344428;
      7422: inst = 32'd203489279;
      7423: inst = 32'd471859200;
      7424: inst = 32'd136314880;
      7425: inst = 32'd268468224;
      7426: inst = 32'd201344429;
      7427: inst = 32'd203489279;
      7428: inst = 32'd471859200;
      7429: inst = 32'd136314880;
      7430: inst = 32'd268468224;
      7431: inst = 32'd201344430;
      7432: inst = 32'd203489279;
      7433: inst = 32'd471859200;
      7434: inst = 32'd136314880;
      7435: inst = 32'd268468224;
      7436: inst = 32'd201344431;
      7437: inst = 32'd203489279;
      7438: inst = 32'd471859200;
      7439: inst = 32'd136314880;
      7440: inst = 32'd268468224;
      7441: inst = 32'd201344432;
      7442: inst = 32'd203489279;
      7443: inst = 32'd471859200;
      7444: inst = 32'd136314880;
      7445: inst = 32'd268468224;
      7446: inst = 32'd201344433;
      7447: inst = 32'd203489279;
      7448: inst = 32'd471859200;
      7449: inst = 32'd136314880;
      7450: inst = 32'd268468224;
      7451: inst = 32'd201344434;
      7452: inst = 32'd203489279;
      7453: inst = 32'd471859200;
      7454: inst = 32'd136314880;
      7455: inst = 32'd268468224;
      7456: inst = 32'd201344435;
      7457: inst = 32'd203489279;
      7458: inst = 32'd471859200;
      7459: inst = 32'd136314880;
      7460: inst = 32'd268468224;
      7461: inst = 32'd201344436;
      7462: inst = 32'd203489279;
      7463: inst = 32'd471859200;
      7464: inst = 32'd136314880;
      7465: inst = 32'd268468224;
      7466: inst = 32'd201344437;
      7467: inst = 32'd203489279;
      7468: inst = 32'd471859200;
      7469: inst = 32'd136314880;
      7470: inst = 32'd268468224;
      7471: inst = 32'd201344438;
      7472: inst = 32'd203489279;
      7473: inst = 32'd471859200;
      7474: inst = 32'd136314880;
      7475: inst = 32'd268468224;
      7476: inst = 32'd201344439;
      7477: inst = 32'd203489279;
      7478: inst = 32'd471859200;
      7479: inst = 32'd136314880;
      7480: inst = 32'd268468224;
      7481: inst = 32'd201344440;
      7482: inst = 32'd203489279;
      7483: inst = 32'd471859200;
      7484: inst = 32'd136314880;
      7485: inst = 32'd268468224;
      7486: inst = 32'd201344441;
      7487: inst = 32'd203489279;
      7488: inst = 32'd471859200;
      7489: inst = 32'd136314880;
      7490: inst = 32'd268468224;
      7491: inst = 32'd201344442;
      7492: inst = 32'd203489279;
      7493: inst = 32'd471859200;
      7494: inst = 32'd136314880;
      7495: inst = 32'd268468224;
      7496: inst = 32'd201344443;
      7497: inst = 32'd203489279;
      7498: inst = 32'd471859200;
      7499: inst = 32'd136314880;
      7500: inst = 32'd268468224;
      7501: inst = 32'd201344444;
      7502: inst = 32'd203489279;
      7503: inst = 32'd471859200;
      7504: inst = 32'd136314880;
      7505: inst = 32'd268468224;
      7506: inst = 32'd201344445;
      7507: inst = 32'd203489279;
      7508: inst = 32'd471859200;
      7509: inst = 32'd136314880;
      7510: inst = 32'd268468224;
      7511: inst = 32'd201344446;
      7512: inst = 32'd203489279;
      7513: inst = 32'd471859200;
      7514: inst = 32'd136314880;
      7515: inst = 32'd268468224;
      7516: inst = 32'd201344447;
      7517: inst = 32'd203489279;
      7518: inst = 32'd471859200;
      7519: inst = 32'd136314880;
      7520: inst = 32'd268468224;
      7521: inst = 32'd201344448;
      7522: inst = 32'd203489279;
      7523: inst = 32'd471859200;
      7524: inst = 32'd136314880;
      7525: inst = 32'd268468224;
      7526: inst = 32'd201344449;
      7527: inst = 32'd203489279;
      7528: inst = 32'd471859200;
      7529: inst = 32'd136314880;
      7530: inst = 32'd268468224;
      7531: inst = 32'd201344450;
      7532: inst = 32'd203489279;
      7533: inst = 32'd471859200;
      7534: inst = 32'd136314880;
      7535: inst = 32'd268468224;
      7536: inst = 32'd201344451;
      7537: inst = 32'd203489279;
      7538: inst = 32'd471859200;
      7539: inst = 32'd136314880;
      7540: inst = 32'd268468224;
      7541: inst = 32'd201344452;
      7542: inst = 32'd203484854;
      7543: inst = 32'd471859200;
      7544: inst = 32'd136314880;
      7545: inst = 32'd268468224;
      7546: inst = 32'd201344453;
      7547: inst = 32'd203484854;
      7548: inst = 32'd471859200;
      7549: inst = 32'd136314880;
      7550: inst = 32'd268468224;
      7551: inst = 32'd201344454;
      7552: inst = 32'd203484854;
      7553: inst = 32'd471859200;
      7554: inst = 32'd136314880;
      7555: inst = 32'd268468224;
      7556: inst = 32'd201344455;
      7557: inst = 32'd203484854;
      7558: inst = 32'd471859200;
      7559: inst = 32'd136314880;
      7560: inst = 32'd268468224;
      7561: inst = 32'd201344456;
      7562: inst = 32'd203484854;
      7563: inst = 32'd471859200;
      7564: inst = 32'd136314880;
      7565: inst = 32'd268468224;
      7566: inst = 32'd201344457;
      7567: inst = 32'd203484854;
      7568: inst = 32'd471859200;
      7569: inst = 32'd136314880;
      7570: inst = 32'd268468224;
      7571: inst = 32'd201344458;
      7572: inst = 32'd203484854;
      7573: inst = 32'd471859200;
      7574: inst = 32'd136314880;
      7575: inst = 32'd268468224;
      7576: inst = 32'd201344459;
      7577: inst = 32'd203484854;
      7578: inst = 32'd471859200;
      7579: inst = 32'd136314880;
      7580: inst = 32'd268468224;
      7581: inst = 32'd201344460;
      7582: inst = 32'd203484854;
      7583: inst = 32'd471859200;
      7584: inst = 32'd136314880;
      7585: inst = 32'd268468224;
      7586: inst = 32'd201344461;
      7587: inst = 32'd203484854;
      7588: inst = 32'd471859200;
      7589: inst = 32'd136314880;
      7590: inst = 32'd268468224;
      7591: inst = 32'd201344462;
      7592: inst = 32'd203484854;
      7593: inst = 32'd471859200;
      7594: inst = 32'd136314880;
      7595: inst = 32'd268468224;
      7596: inst = 32'd201344463;
      7597: inst = 32'd203484854;
      7598: inst = 32'd471859200;
      7599: inst = 32'd136314880;
      7600: inst = 32'd268468224;
      7601: inst = 32'd201344464;
      7602: inst = 32'd203484854;
      7603: inst = 32'd471859200;
      7604: inst = 32'd136314880;
      7605: inst = 32'd268468224;
      7606: inst = 32'd201344465;
      7607: inst = 32'd203484854;
      7608: inst = 32'd471859200;
      7609: inst = 32'd136314880;
      7610: inst = 32'd268468224;
      7611: inst = 32'd201344466;
      7612: inst = 32'd203484854;
      7613: inst = 32'd471859200;
      7614: inst = 32'd136314880;
      7615: inst = 32'd268468224;
      7616: inst = 32'd201344467;
      7617: inst = 32'd203484854;
      7618: inst = 32'd471859200;
      7619: inst = 32'd136314880;
      7620: inst = 32'd268468224;
      7621: inst = 32'd201344468;
      7622: inst = 32'd203484854;
      7623: inst = 32'd471859200;
      7624: inst = 32'd136314880;
      7625: inst = 32'd268468224;
      7626: inst = 32'd201344469;
      7627: inst = 32'd203484854;
      7628: inst = 32'd471859200;
      7629: inst = 32'd136314880;
      7630: inst = 32'd268468224;
      7631: inst = 32'd201344470;
      7632: inst = 32'd203484854;
      7633: inst = 32'd471859200;
      7634: inst = 32'd136314880;
      7635: inst = 32'd268468224;
      7636: inst = 32'd201344471;
      7637: inst = 32'd203484854;
      7638: inst = 32'd471859200;
      7639: inst = 32'd136314880;
      7640: inst = 32'd268468224;
      7641: inst = 32'd201344472;
      7642: inst = 32'd203484854;
      7643: inst = 32'd471859200;
      7644: inst = 32'd136314880;
      7645: inst = 32'd268468224;
      7646: inst = 32'd201344473;
      7647: inst = 32'd203484854;
      7648: inst = 32'd471859200;
      7649: inst = 32'd136314880;
      7650: inst = 32'd268468224;
      7651: inst = 32'd201344474;
      7652: inst = 32'd203484854;
      7653: inst = 32'd471859200;
      7654: inst = 32'd136314880;
      7655: inst = 32'd268468224;
      7656: inst = 32'd201344475;
      7657: inst = 32'd203484854;
      7658: inst = 32'd471859200;
      7659: inst = 32'd136314880;
      7660: inst = 32'd268468224;
      7661: inst = 32'd201344476;
      7662: inst = 32'd203484854;
      7663: inst = 32'd471859200;
      7664: inst = 32'd136314880;
      7665: inst = 32'd268468224;
      7666: inst = 32'd201344477;
      7667: inst = 32'd203484854;
      7668: inst = 32'd471859200;
      7669: inst = 32'd136314880;
      7670: inst = 32'd268468224;
      7671: inst = 32'd201344478;
      7672: inst = 32'd203484854;
      7673: inst = 32'd471859200;
      7674: inst = 32'd136314880;
      7675: inst = 32'd268468224;
      7676: inst = 32'd201344479;
      7677: inst = 32'd203484854;
      7678: inst = 32'd471859200;
      7679: inst = 32'd136314880;
      7680: inst = 32'd268468224;
      7681: inst = 32'd201344480;
      7682: inst = 32'd203484854;
      7683: inst = 32'd471859200;
      7684: inst = 32'd136314880;
      7685: inst = 32'd268468224;
      7686: inst = 32'd201344481;
      7687: inst = 32'd203484854;
      7688: inst = 32'd471859200;
      7689: inst = 32'd136314880;
      7690: inst = 32'd268468224;
      7691: inst = 32'd201344482;
      7692: inst = 32'd203484854;
      7693: inst = 32'd471859200;
      7694: inst = 32'd136314880;
      7695: inst = 32'd268468224;
      7696: inst = 32'd201344483;
      7697: inst = 32'd203484854;
      7698: inst = 32'd471859200;
      7699: inst = 32'd136314880;
      7700: inst = 32'd268468224;
      7701: inst = 32'd201344484;
      7702: inst = 32'd203484854;
      7703: inst = 32'd471859200;
      7704: inst = 32'd136314880;
      7705: inst = 32'd268468224;
      7706: inst = 32'd201344485;
      7707: inst = 32'd203484854;
      7708: inst = 32'd471859200;
      7709: inst = 32'd136314880;
      7710: inst = 32'd268468224;
      7711: inst = 32'd201344486;
      7712: inst = 32'd203484854;
      7713: inst = 32'd471859200;
      7714: inst = 32'd136314880;
      7715: inst = 32'd268468224;
      7716: inst = 32'd201344487;
      7717: inst = 32'd203484854;
      7718: inst = 32'd471859200;
      7719: inst = 32'd136314880;
      7720: inst = 32'd268468224;
      7721: inst = 32'd201344488;
      7722: inst = 32'd203484854;
      7723: inst = 32'd471859200;
      7724: inst = 32'd136314880;
      7725: inst = 32'd268468224;
      7726: inst = 32'd201344489;
      7727: inst = 32'd203484854;
      7728: inst = 32'd471859200;
      7729: inst = 32'd136314880;
      7730: inst = 32'd268468224;
      7731: inst = 32'd201344490;
      7732: inst = 32'd203484854;
      7733: inst = 32'd471859200;
      7734: inst = 32'd136314880;
      7735: inst = 32'd268468224;
      7736: inst = 32'd201344491;
      7737: inst = 32'd203484854;
      7738: inst = 32'd471859200;
      7739: inst = 32'd136314880;
      7740: inst = 32'd268468224;
      7741: inst = 32'd201344492;
      7742: inst = 32'd203484854;
      7743: inst = 32'd471859200;
      7744: inst = 32'd136314880;
      7745: inst = 32'd268468224;
      7746: inst = 32'd201344493;
      7747: inst = 32'd203484854;
      7748: inst = 32'd471859200;
      7749: inst = 32'd136314880;
      7750: inst = 32'd268468224;
      7751: inst = 32'd201344494;
      7752: inst = 32'd203484854;
      7753: inst = 32'd471859200;
      7754: inst = 32'd136314880;
      7755: inst = 32'd268468224;
      7756: inst = 32'd201344495;
      7757: inst = 32'd203484854;
      7758: inst = 32'd471859200;
      7759: inst = 32'd136314880;
      7760: inst = 32'd268468224;
      7761: inst = 32'd201344496;
      7762: inst = 32'd203484854;
      7763: inst = 32'd471859200;
      7764: inst = 32'd136314880;
      7765: inst = 32'd268468224;
      7766: inst = 32'd201344497;
      7767: inst = 32'd203484854;
      7768: inst = 32'd471859200;
      7769: inst = 32'd136314880;
      7770: inst = 32'd268468224;
      7771: inst = 32'd201344498;
      7772: inst = 32'd203484854;
      7773: inst = 32'd471859200;
      7774: inst = 32'd136314880;
      7775: inst = 32'd268468224;
      7776: inst = 32'd201344499;
      7777: inst = 32'd203484854;
      7778: inst = 32'd471859200;
      7779: inst = 32'd136314880;
      7780: inst = 32'd268468224;
      7781: inst = 32'd201344500;
      7782: inst = 32'd203484854;
      7783: inst = 32'd471859200;
      7784: inst = 32'd136314880;
      7785: inst = 32'd268468224;
      7786: inst = 32'd201344501;
      7787: inst = 32'd203484854;
      7788: inst = 32'd471859200;
      7789: inst = 32'd136314880;
      7790: inst = 32'd268468224;
      7791: inst = 32'd201344502;
      7792: inst = 32'd203484854;
      7793: inst = 32'd471859200;
      7794: inst = 32'd136314880;
      7795: inst = 32'd268468224;
      7796: inst = 32'd201344503;
      7797: inst = 32'd203484854;
      7798: inst = 32'd471859200;
      7799: inst = 32'd136314880;
      7800: inst = 32'd268468224;
      7801: inst = 32'd201344504;
      7802: inst = 32'd203484854;
      7803: inst = 32'd471859200;
      7804: inst = 32'd136314880;
      7805: inst = 32'd268468224;
      7806: inst = 32'd201344505;
      7807: inst = 32'd203484854;
      7808: inst = 32'd471859200;
      7809: inst = 32'd136314880;
      7810: inst = 32'd268468224;
      7811: inst = 32'd201344506;
      7812: inst = 32'd203484854;
      7813: inst = 32'd471859200;
      7814: inst = 32'd136314880;
      7815: inst = 32'd268468224;
      7816: inst = 32'd201344507;
      7817: inst = 32'd203484854;
      7818: inst = 32'd471859200;
      7819: inst = 32'd136314880;
      7820: inst = 32'd268468224;
      7821: inst = 32'd201344508;
      7822: inst = 32'd203489279;
      7823: inst = 32'd471859200;
      7824: inst = 32'd136314880;
      7825: inst = 32'd268468224;
      7826: inst = 32'd201344509;
      7827: inst = 32'd203489279;
      7828: inst = 32'd471859200;
      7829: inst = 32'd136314880;
      7830: inst = 32'd268468224;
      7831: inst = 32'd201344510;
      7832: inst = 32'd203489279;
      7833: inst = 32'd471859200;
      7834: inst = 32'd136314880;
      7835: inst = 32'd268468224;
      7836: inst = 32'd201344511;
      7837: inst = 32'd203489279;
      7838: inst = 32'd471859200;
      7839: inst = 32'd136314880;
      7840: inst = 32'd268468224;
      7841: inst = 32'd201344512;
      7842: inst = 32'd203489279;
      7843: inst = 32'd471859200;
      7844: inst = 32'd136314880;
      7845: inst = 32'd268468224;
      7846: inst = 32'd201344513;
      7847: inst = 32'd203489279;
      7848: inst = 32'd471859200;
      7849: inst = 32'd136314880;
      7850: inst = 32'd268468224;
      7851: inst = 32'd201344514;
      7852: inst = 32'd203489279;
      7853: inst = 32'd471859200;
      7854: inst = 32'd136314880;
      7855: inst = 32'd268468224;
      7856: inst = 32'd201344515;
      7857: inst = 32'd203489279;
      7858: inst = 32'd471859200;
      7859: inst = 32'd136314880;
      7860: inst = 32'd268468224;
      7861: inst = 32'd201344516;
      7862: inst = 32'd203489279;
      7863: inst = 32'd471859200;
      7864: inst = 32'd136314880;
      7865: inst = 32'd268468224;
      7866: inst = 32'd201344517;
      7867: inst = 32'd203489279;
      7868: inst = 32'd471859200;
      7869: inst = 32'd136314880;
      7870: inst = 32'd268468224;
      7871: inst = 32'd201344518;
      7872: inst = 32'd203489279;
      7873: inst = 32'd471859200;
      7874: inst = 32'd136314880;
      7875: inst = 32'd268468224;
      7876: inst = 32'd201344519;
      7877: inst = 32'd203489279;
      7878: inst = 32'd471859200;
      7879: inst = 32'd136314880;
      7880: inst = 32'd268468224;
      7881: inst = 32'd201344520;
      7882: inst = 32'd203489279;
      7883: inst = 32'd471859200;
      7884: inst = 32'd136314880;
      7885: inst = 32'd268468224;
      7886: inst = 32'd201344521;
      7887: inst = 32'd203489279;
      7888: inst = 32'd471859200;
      7889: inst = 32'd136314880;
      7890: inst = 32'd268468224;
      7891: inst = 32'd201344522;
      7892: inst = 32'd203489279;
      7893: inst = 32'd471859200;
      7894: inst = 32'd136314880;
      7895: inst = 32'd268468224;
      7896: inst = 32'd201344523;
      7897: inst = 32'd203489279;
      7898: inst = 32'd471859200;
      7899: inst = 32'd136314880;
      7900: inst = 32'd268468224;
      7901: inst = 32'd201344524;
      7902: inst = 32'd203489279;
      7903: inst = 32'd471859200;
      7904: inst = 32'd136314880;
      7905: inst = 32'd268468224;
      7906: inst = 32'd201344525;
      7907: inst = 32'd203489279;
      7908: inst = 32'd471859200;
      7909: inst = 32'd136314880;
      7910: inst = 32'd268468224;
      7911: inst = 32'd201344526;
      7912: inst = 32'd203489279;
      7913: inst = 32'd471859200;
      7914: inst = 32'd136314880;
      7915: inst = 32'd268468224;
      7916: inst = 32'd201344527;
      7917: inst = 32'd203489279;
      7918: inst = 32'd471859200;
      7919: inst = 32'd136314880;
      7920: inst = 32'd268468224;
      7921: inst = 32'd201344528;
      7922: inst = 32'd203489279;
      7923: inst = 32'd471859200;
      7924: inst = 32'd136314880;
      7925: inst = 32'd268468224;
      7926: inst = 32'd201344529;
      7927: inst = 32'd203489279;
      7928: inst = 32'd471859200;
      7929: inst = 32'd136314880;
      7930: inst = 32'd268468224;
      7931: inst = 32'd201344530;
      7932: inst = 32'd203489279;
      7933: inst = 32'd471859200;
      7934: inst = 32'd136314880;
      7935: inst = 32'd268468224;
      7936: inst = 32'd201344531;
      7937: inst = 32'd203489279;
      7938: inst = 32'd471859200;
      7939: inst = 32'd136314880;
      7940: inst = 32'd268468224;
      7941: inst = 32'd201344532;
      7942: inst = 32'd203489279;
      7943: inst = 32'd471859200;
      7944: inst = 32'd136314880;
      7945: inst = 32'd268468224;
      7946: inst = 32'd201344533;
      7947: inst = 32'd203489279;
      7948: inst = 32'd471859200;
      7949: inst = 32'd136314880;
      7950: inst = 32'd268468224;
      7951: inst = 32'd201344534;
      7952: inst = 32'd203489279;
      7953: inst = 32'd471859200;
      7954: inst = 32'd136314880;
      7955: inst = 32'd268468224;
      7956: inst = 32'd201344535;
      7957: inst = 32'd203489279;
      7958: inst = 32'd471859200;
      7959: inst = 32'd136314880;
      7960: inst = 32'd268468224;
      7961: inst = 32'd201344536;
      7962: inst = 32'd203489279;
      7963: inst = 32'd471859200;
      7964: inst = 32'd136314880;
      7965: inst = 32'd268468224;
      7966: inst = 32'd201344537;
      7967: inst = 32'd203489279;
      7968: inst = 32'd471859200;
      7969: inst = 32'd136314880;
      7970: inst = 32'd268468224;
      7971: inst = 32'd201344538;
      7972: inst = 32'd203489279;
      7973: inst = 32'd471859200;
      7974: inst = 32'd136314880;
      7975: inst = 32'd268468224;
      7976: inst = 32'd201344539;
      7977: inst = 32'd203489279;
      7978: inst = 32'd471859200;
      7979: inst = 32'd136314880;
      7980: inst = 32'd268468224;
      7981: inst = 32'd201344540;
      7982: inst = 32'd203489279;
      7983: inst = 32'd471859200;
      7984: inst = 32'd136314880;
      7985: inst = 32'd268468224;
      7986: inst = 32'd201344541;
      7987: inst = 32'd203489279;
      7988: inst = 32'd471859200;
      7989: inst = 32'd136314880;
      7990: inst = 32'd268468224;
      7991: inst = 32'd201344542;
      7992: inst = 32'd203489279;
      7993: inst = 32'd471859200;
      7994: inst = 32'd136314880;
      7995: inst = 32'd268468224;
      7996: inst = 32'd201344543;
      7997: inst = 32'd203489279;
      7998: inst = 32'd471859200;
      7999: inst = 32'd136314880;
      8000: inst = 32'd268468224;
      8001: inst = 32'd201344544;
      8002: inst = 32'd203489279;
      8003: inst = 32'd471859200;
      8004: inst = 32'd136314880;
      8005: inst = 32'd268468224;
      8006: inst = 32'd201344545;
      8007: inst = 32'd203489279;
      8008: inst = 32'd471859200;
      8009: inst = 32'd136314880;
      8010: inst = 32'd268468224;
      8011: inst = 32'd201344546;
      8012: inst = 32'd203489279;
      8013: inst = 32'd471859200;
      8014: inst = 32'd136314880;
      8015: inst = 32'd268468224;
      8016: inst = 32'd201344547;
      8017: inst = 32'd203489279;
      8018: inst = 32'd471859200;
      8019: inst = 32'd136314880;
      8020: inst = 32'd268468224;
      8021: inst = 32'd201344548;
      8022: inst = 32'd203484854;
      8023: inst = 32'd471859200;
      8024: inst = 32'd136314880;
      8025: inst = 32'd268468224;
      8026: inst = 32'd201344549;
      8027: inst = 32'd203484854;
      8028: inst = 32'd471859200;
      8029: inst = 32'd136314880;
      8030: inst = 32'd268468224;
      8031: inst = 32'd201344550;
      8032: inst = 32'd203484854;
      8033: inst = 32'd471859200;
      8034: inst = 32'd136314880;
      8035: inst = 32'd268468224;
      8036: inst = 32'd201344551;
      8037: inst = 32'd203484854;
      8038: inst = 32'd471859200;
      8039: inst = 32'd136314880;
      8040: inst = 32'd268468224;
      8041: inst = 32'd201344552;
      8042: inst = 32'd203484854;
      8043: inst = 32'd471859200;
      8044: inst = 32'd136314880;
      8045: inst = 32'd268468224;
      8046: inst = 32'd201344553;
      8047: inst = 32'd203484854;
      8048: inst = 32'd471859200;
      8049: inst = 32'd136314880;
      8050: inst = 32'd268468224;
      8051: inst = 32'd201344554;
      8052: inst = 32'd203484854;
      8053: inst = 32'd471859200;
      8054: inst = 32'd136314880;
      8055: inst = 32'd268468224;
      8056: inst = 32'd201344555;
      8057: inst = 32'd203484854;
      8058: inst = 32'd471859200;
      8059: inst = 32'd136314880;
      8060: inst = 32'd268468224;
      8061: inst = 32'd201344556;
      8062: inst = 32'd203484854;
      8063: inst = 32'd471859200;
      8064: inst = 32'd136314880;
      8065: inst = 32'd268468224;
      8066: inst = 32'd201344557;
      8067: inst = 32'd203484854;
      8068: inst = 32'd471859200;
      8069: inst = 32'd136314880;
      8070: inst = 32'd268468224;
      8071: inst = 32'd201344558;
      8072: inst = 32'd203484854;
      8073: inst = 32'd471859200;
      8074: inst = 32'd136314880;
      8075: inst = 32'd268468224;
      8076: inst = 32'd201344559;
      8077: inst = 32'd203484854;
      8078: inst = 32'd471859200;
      8079: inst = 32'd136314880;
      8080: inst = 32'd268468224;
      8081: inst = 32'd201344560;
      8082: inst = 32'd203484854;
      8083: inst = 32'd471859200;
      8084: inst = 32'd136314880;
      8085: inst = 32'd268468224;
      8086: inst = 32'd201344561;
      8087: inst = 32'd203484854;
      8088: inst = 32'd471859200;
      8089: inst = 32'd136314880;
      8090: inst = 32'd268468224;
      8091: inst = 32'd201344562;
      8092: inst = 32'd203484854;
      8093: inst = 32'd471859200;
      8094: inst = 32'd136314880;
      8095: inst = 32'd268468224;
      8096: inst = 32'd201344563;
      8097: inst = 32'd203484854;
      8098: inst = 32'd471859200;
      8099: inst = 32'd136314880;
      8100: inst = 32'd268468224;
      8101: inst = 32'd201344564;
      8102: inst = 32'd203484854;
      8103: inst = 32'd471859200;
      8104: inst = 32'd136314880;
      8105: inst = 32'd268468224;
      8106: inst = 32'd201344565;
      8107: inst = 32'd203484854;
      8108: inst = 32'd471859200;
      8109: inst = 32'd136314880;
      8110: inst = 32'd268468224;
      8111: inst = 32'd201344566;
      8112: inst = 32'd203484854;
      8113: inst = 32'd471859200;
      8114: inst = 32'd136314880;
      8115: inst = 32'd268468224;
      8116: inst = 32'd201344567;
      8117: inst = 32'd203484854;
      8118: inst = 32'd471859200;
      8119: inst = 32'd136314880;
      8120: inst = 32'd268468224;
      8121: inst = 32'd201344568;
      8122: inst = 32'd203484854;
      8123: inst = 32'd471859200;
      8124: inst = 32'd136314880;
      8125: inst = 32'd268468224;
      8126: inst = 32'd201344569;
      8127: inst = 32'd203484854;
      8128: inst = 32'd471859200;
      8129: inst = 32'd136314880;
      8130: inst = 32'd268468224;
      8131: inst = 32'd201344570;
      8132: inst = 32'd203484854;
      8133: inst = 32'd471859200;
      8134: inst = 32'd136314880;
      8135: inst = 32'd268468224;
      8136: inst = 32'd201344571;
      8137: inst = 32'd203484854;
      8138: inst = 32'd471859200;
      8139: inst = 32'd136314880;
      8140: inst = 32'd268468224;
      8141: inst = 32'd201344572;
      8142: inst = 32'd203484854;
      8143: inst = 32'd471859200;
      8144: inst = 32'd136314880;
      8145: inst = 32'd268468224;
      8146: inst = 32'd201344573;
      8147: inst = 32'd203484854;
      8148: inst = 32'd471859200;
      8149: inst = 32'd136314880;
      8150: inst = 32'd268468224;
      8151: inst = 32'd201344574;
      8152: inst = 32'd203484854;
      8153: inst = 32'd471859200;
      8154: inst = 32'd136314880;
      8155: inst = 32'd268468224;
      8156: inst = 32'd201344575;
      8157: inst = 32'd203484854;
      8158: inst = 32'd471859200;
      8159: inst = 32'd136314880;
      8160: inst = 32'd268468224;
      8161: inst = 32'd201344576;
      8162: inst = 32'd203484854;
      8163: inst = 32'd471859200;
      8164: inst = 32'd136314880;
      8165: inst = 32'd268468224;
      8166: inst = 32'd201344577;
      8167: inst = 32'd203484854;
      8168: inst = 32'd471859200;
      8169: inst = 32'd136314880;
      8170: inst = 32'd268468224;
      8171: inst = 32'd201344578;
      8172: inst = 32'd203484854;
      8173: inst = 32'd471859200;
      8174: inst = 32'd136314880;
      8175: inst = 32'd268468224;
      8176: inst = 32'd201344579;
      8177: inst = 32'd203484854;
      8178: inst = 32'd471859200;
      8179: inst = 32'd136314880;
      8180: inst = 32'd268468224;
      8181: inst = 32'd201344580;
      8182: inst = 32'd203484854;
      8183: inst = 32'd471859200;
      8184: inst = 32'd136314880;
      8185: inst = 32'd268468224;
      8186: inst = 32'd201344581;
      8187: inst = 32'd203484854;
      8188: inst = 32'd471859200;
      8189: inst = 32'd136314880;
      8190: inst = 32'd268468224;
      8191: inst = 32'd201344582;
      8192: inst = 32'd203484854;
      8193: inst = 32'd471859200;
      8194: inst = 32'd136314880;
      8195: inst = 32'd268468224;
      8196: inst = 32'd201344583;
      8197: inst = 32'd203484854;
      8198: inst = 32'd471859200;
      8199: inst = 32'd136314880;
      8200: inst = 32'd268468224;
      8201: inst = 32'd201344584;
      8202: inst = 32'd203484854;
      8203: inst = 32'd471859200;
      8204: inst = 32'd136314880;
      8205: inst = 32'd268468224;
      8206: inst = 32'd201344585;
      8207: inst = 32'd203484854;
      8208: inst = 32'd471859200;
      8209: inst = 32'd136314880;
      8210: inst = 32'd268468224;
      8211: inst = 32'd201344586;
      8212: inst = 32'd203484854;
      8213: inst = 32'd471859200;
      8214: inst = 32'd136314880;
      8215: inst = 32'd268468224;
      8216: inst = 32'd201344587;
      8217: inst = 32'd203484854;
      8218: inst = 32'd471859200;
      8219: inst = 32'd136314880;
      8220: inst = 32'd268468224;
      8221: inst = 32'd201344588;
      8222: inst = 32'd203484854;
      8223: inst = 32'd471859200;
      8224: inst = 32'd136314880;
      8225: inst = 32'd268468224;
      8226: inst = 32'd201344589;
      8227: inst = 32'd203484854;
      8228: inst = 32'd471859200;
      8229: inst = 32'd136314880;
      8230: inst = 32'd268468224;
      8231: inst = 32'd201344590;
      8232: inst = 32'd203484854;
      8233: inst = 32'd471859200;
      8234: inst = 32'd136314880;
      8235: inst = 32'd268468224;
      8236: inst = 32'd201344591;
      8237: inst = 32'd203484854;
      8238: inst = 32'd471859200;
      8239: inst = 32'd136314880;
      8240: inst = 32'd268468224;
      8241: inst = 32'd201344592;
      8242: inst = 32'd203484854;
      8243: inst = 32'd471859200;
      8244: inst = 32'd136314880;
      8245: inst = 32'd268468224;
      8246: inst = 32'd201344593;
      8247: inst = 32'd203484854;
      8248: inst = 32'd471859200;
      8249: inst = 32'd136314880;
      8250: inst = 32'd268468224;
      8251: inst = 32'd201344594;
      8252: inst = 32'd203484854;
      8253: inst = 32'd471859200;
      8254: inst = 32'd136314880;
      8255: inst = 32'd268468224;
      8256: inst = 32'd201344595;
      8257: inst = 32'd203484854;
      8258: inst = 32'd471859200;
      8259: inst = 32'd136314880;
      8260: inst = 32'd268468224;
      8261: inst = 32'd201344596;
      8262: inst = 32'd203484854;
      8263: inst = 32'd471859200;
      8264: inst = 32'd136314880;
      8265: inst = 32'd268468224;
      8266: inst = 32'd201344597;
      8267: inst = 32'd203484854;
      8268: inst = 32'd471859200;
      8269: inst = 32'd136314880;
      8270: inst = 32'd268468224;
      8271: inst = 32'd201344598;
      8272: inst = 32'd203484854;
      8273: inst = 32'd471859200;
      8274: inst = 32'd136314880;
      8275: inst = 32'd268468224;
      8276: inst = 32'd201344599;
      8277: inst = 32'd203484854;
      8278: inst = 32'd471859200;
      8279: inst = 32'd136314880;
      8280: inst = 32'd268468224;
      8281: inst = 32'd201344600;
      8282: inst = 32'd203484854;
      8283: inst = 32'd471859200;
      8284: inst = 32'd136314880;
      8285: inst = 32'd268468224;
      8286: inst = 32'd201344601;
      8287: inst = 32'd203484854;
      8288: inst = 32'd471859200;
      8289: inst = 32'd136314880;
      8290: inst = 32'd268468224;
      8291: inst = 32'd201344602;
      8292: inst = 32'd203484854;
      8293: inst = 32'd471859200;
      8294: inst = 32'd136314880;
      8295: inst = 32'd268468224;
      8296: inst = 32'd201344603;
      8297: inst = 32'd203484854;
      8298: inst = 32'd471859200;
      8299: inst = 32'd136314880;
      8300: inst = 32'd268468224;
      8301: inst = 32'd201344604;
      8302: inst = 32'd203489279;
      8303: inst = 32'd471859200;
      8304: inst = 32'd136314880;
      8305: inst = 32'd268468224;
      8306: inst = 32'd201344605;
      8307: inst = 32'd203489279;
      8308: inst = 32'd471859200;
      8309: inst = 32'd136314880;
      8310: inst = 32'd268468224;
      8311: inst = 32'd201344606;
      8312: inst = 32'd203489279;
      8313: inst = 32'd471859200;
      8314: inst = 32'd136314880;
      8315: inst = 32'd268468224;
      8316: inst = 32'd201344607;
      8317: inst = 32'd203489279;
      8318: inst = 32'd471859200;
      8319: inst = 32'd136314880;
      8320: inst = 32'd268468224;
      8321: inst = 32'd201344608;
      8322: inst = 32'd203489279;
      8323: inst = 32'd471859200;
      8324: inst = 32'd136314880;
      8325: inst = 32'd268468224;
      8326: inst = 32'd201344609;
      8327: inst = 32'd203489279;
      8328: inst = 32'd471859200;
      8329: inst = 32'd136314880;
      8330: inst = 32'd268468224;
      8331: inst = 32'd201344610;
      8332: inst = 32'd203489279;
      8333: inst = 32'd471859200;
      8334: inst = 32'd136314880;
      8335: inst = 32'd268468224;
      8336: inst = 32'd201344611;
      8337: inst = 32'd203489279;
      8338: inst = 32'd471859200;
      8339: inst = 32'd136314880;
      8340: inst = 32'd268468224;
      8341: inst = 32'd201344612;
      8342: inst = 32'd203489279;
      8343: inst = 32'd471859200;
      8344: inst = 32'd136314880;
      8345: inst = 32'd268468224;
      8346: inst = 32'd201344613;
      8347: inst = 32'd203489279;
      8348: inst = 32'd471859200;
      8349: inst = 32'd136314880;
      8350: inst = 32'd268468224;
      8351: inst = 32'd201344614;
      8352: inst = 32'd203489279;
      8353: inst = 32'd471859200;
      8354: inst = 32'd136314880;
      8355: inst = 32'd268468224;
      8356: inst = 32'd201344615;
      8357: inst = 32'd203489279;
      8358: inst = 32'd471859200;
      8359: inst = 32'd136314880;
      8360: inst = 32'd268468224;
      8361: inst = 32'd201344616;
      8362: inst = 32'd203489279;
      8363: inst = 32'd471859200;
      8364: inst = 32'd136314880;
      8365: inst = 32'd268468224;
      8366: inst = 32'd201344617;
      8367: inst = 32'd203489279;
      8368: inst = 32'd471859200;
      8369: inst = 32'd136314880;
      8370: inst = 32'd268468224;
      8371: inst = 32'd201344618;
      8372: inst = 32'd203489279;
      8373: inst = 32'd471859200;
      8374: inst = 32'd136314880;
      8375: inst = 32'd268468224;
      8376: inst = 32'd201344619;
      8377: inst = 32'd203489279;
      8378: inst = 32'd471859200;
      8379: inst = 32'd136314880;
      8380: inst = 32'd268468224;
      8381: inst = 32'd201344620;
      8382: inst = 32'd203489279;
      8383: inst = 32'd471859200;
      8384: inst = 32'd136314880;
      8385: inst = 32'd268468224;
      8386: inst = 32'd201344621;
      8387: inst = 32'd203489279;
      8388: inst = 32'd471859200;
      8389: inst = 32'd136314880;
      8390: inst = 32'd268468224;
      8391: inst = 32'd201344622;
      8392: inst = 32'd203489279;
      8393: inst = 32'd471859200;
      8394: inst = 32'd136314880;
      8395: inst = 32'd268468224;
      8396: inst = 32'd201344623;
      8397: inst = 32'd203489279;
      8398: inst = 32'd471859200;
      8399: inst = 32'd136314880;
      8400: inst = 32'd268468224;
      8401: inst = 32'd201344624;
      8402: inst = 32'd203489279;
      8403: inst = 32'd471859200;
      8404: inst = 32'd136314880;
      8405: inst = 32'd268468224;
      8406: inst = 32'd201344625;
      8407: inst = 32'd203489279;
      8408: inst = 32'd471859200;
      8409: inst = 32'd136314880;
      8410: inst = 32'd268468224;
      8411: inst = 32'd201344626;
      8412: inst = 32'd203489279;
      8413: inst = 32'd471859200;
      8414: inst = 32'd136314880;
      8415: inst = 32'd268468224;
      8416: inst = 32'd201344627;
      8417: inst = 32'd203489279;
      8418: inst = 32'd471859200;
      8419: inst = 32'd136314880;
      8420: inst = 32'd268468224;
      8421: inst = 32'd201344628;
      8422: inst = 32'd203489279;
      8423: inst = 32'd471859200;
      8424: inst = 32'd136314880;
      8425: inst = 32'd268468224;
      8426: inst = 32'd201344629;
      8427: inst = 32'd203489279;
      8428: inst = 32'd471859200;
      8429: inst = 32'd136314880;
      8430: inst = 32'd268468224;
      8431: inst = 32'd201344630;
      8432: inst = 32'd203489279;
      8433: inst = 32'd471859200;
      8434: inst = 32'd136314880;
      8435: inst = 32'd268468224;
      8436: inst = 32'd201344631;
      8437: inst = 32'd203489279;
      8438: inst = 32'd471859200;
      8439: inst = 32'd136314880;
      8440: inst = 32'd268468224;
      8441: inst = 32'd201344632;
      8442: inst = 32'd203489279;
      8443: inst = 32'd471859200;
      8444: inst = 32'd136314880;
      8445: inst = 32'd268468224;
      8446: inst = 32'd201344633;
      8447: inst = 32'd203489279;
      8448: inst = 32'd471859200;
      8449: inst = 32'd136314880;
      8450: inst = 32'd268468224;
      8451: inst = 32'd201344634;
      8452: inst = 32'd203489279;
      8453: inst = 32'd471859200;
      8454: inst = 32'd136314880;
      8455: inst = 32'd268468224;
      8456: inst = 32'd201344635;
      8457: inst = 32'd203489279;
      8458: inst = 32'd471859200;
      8459: inst = 32'd136314880;
      8460: inst = 32'd268468224;
      8461: inst = 32'd201344636;
      8462: inst = 32'd203489279;
      8463: inst = 32'd471859200;
      8464: inst = 32'd136314880;
      8465: inst = 32'd268468224;
      8466: inst = 32'd201344637;
      8467: inst = 32'd203489279;
      8468: inst = 32'd471859200;
      8469: inst = 32'd136314880;
      8470: inst = 32'd268468224;
      8471: inst = 32'd201344638;
      8472: inst = 32'd203489279;
      8473: inst = 32'd471859200;
      8474: inst = 32'd136314880;
      8475: inst = 32'd268468224;
      8476: inst = 32'd201344639;
      8477: inst = 32'd203489279;
      8478: inst = 32'd471859200;
      8479: inst = 32'd136314880;
      8480: inst = 32'd268468224;
      8481: inst = 32'd201344640;
      8482: inst = 32'd203489279;
      8483: inst = 32'd471859200;
      8484: inst = 32'd136314880;
      8485: inst = 32'd268468224;
      8486: inst = 32'd201344641;
      8487: inst = 32'd203489279;
      8488: inst = 32'd471859200;
      8489: inst = 32'd136314880;
      8490: inst = 32'd268468224;
      8491: inst = 32'd201344642;
      8492: inst = 32'd203489279;
      8493: inst = 32'd471859200;
      8494: inst = 32'd136314880;
      8495: inst = 32'd268468224;
      8496: inst = 32'd201344643;
      8497: inst = 32'd203489279;
      8498: inst = 32'd471859200;
      8499: inst = 32'd136314880;
      8500: inst = 32'd268468224;
      8501: inst = 32'd201344644;
      8502: inst = 32'd203484854;
      8503: inst = 32'd471859200;
      8504: inst = 32'd136314880;
      8505: inst = 32'd268468224;
      8506: inst = 32'd201344645;
      8507: inst = 32'd203484854;
      8508: inst = 32'd471859200;
      8509: inst = 32'd136314880;
      8510: inst = 32'd268468224;
      8511: inst = 32'd201344646;
      8512: inst = 32'd203484854;
      8513: inst = 32'd471859200;
      8514: inst = 32'd136314880;
      8515: inst = 32'd268468224;
      8516: inst = 32'd201344647;
      8517: inst = 32'd203484854;
      8518: inst = 32'd471859200;
      8519: inst = 32'd136314880;
      8520: inst = 32'd268468224;
      8521: inst = 32'd201344648;
      8522: inst = 32'd203484854;
      8523: inst = 32'd471859200;
      8524: inst = 32'd136314880;
      8525: inst = 32'd268468224;
      8526: inst = 32'd201344649;
      8527: inst = 32'd203484854;
      8528: inst = 32'd471859200;
      8529: inst = 32'd136314880;
      8530: inst = 32'd268468224;
      8531: inst = 32'd201344650;
      8532: inst = 32'd203484854;
      8533: inst = 32'd471859200;
      8534: inst = 32'd136314880;
      8535: inst = 32'd268468224;
      8536: inst = 32'd201344651;
      8537: inst = 32'd203484854;
      8538: inst = 32'd471859200;
      8539: inst = 32'd136314880;
      8540: inst = 32'd268468224;
      8541: inst = 32'd201344652;
      8542: inst = 32'd203484854;
      8543: inst = 32'd471859200;
      8544: inst = 32'd136314880;
      8545: inst = 32'd268468224;
      8546: inst = 32'd201344653;
      8547: inst = 32'd203484854;
      8548: inst = 32'd471859200;
      8549: inst = 32'd136314880;
      8550: inst = 32'd268468224;
      8551: inst = 32'd201344654;
      8552: inst = 32'd203484854;
      8553: inst = 32'd471859200;
      8554: inst = 32'd136314880;
      8555: inst = 32'd268468224;
      8556: inst = 32'd201344655;
      8557: inst = 32'd203484854;
      8558: inst = 32'd471859200;
      8559: inst = 32'd136314880;
      8560: inst = 32'd268468224;
      8561: inst = 32'd201344656;
      8562: inst = 32'd203484854;
      8563: inst = 32'd471859200;
      8564: inst = 32'd136314880;
      8565: inst = 32'd268468224;
      8566: inst = 32'd201344657;
      8567: inst = 32'd203484854;
      8568: inst = 32'd471859200;
      8569: inst = 32'd136314880;
      8570: inst = 32'd268468224;
      8571: inst = 32'd201344658;
      8572: inst = 32'd203484854;
      8573: inst = 32'd471859200;
      8574: inst = 32'd136314880;
      8575: inst = 32'd268468224;
      8576: inst = 32'd201344659;
      8577: inst = 32'd203484854;
      8578: inst = 32'd471859200;
      8579: inst = 32'd136314880;
      8580: inst = 32'd268468224;
      8581: inst = 32'd201344660;
      8582: inst = 32'd203484854;
      8583: inst = 32'd471859200;
      8584: inst = 32'd136314880;
      8585: inst = 32'd268468224;
      8586: inst = 32'd201344661;
      8587: inst = 32'd203484854;
      8588: inst = 32'd471859200;
      8589: inst = 32'd136314880;
      8590: inst = 32'd268468224;
      8591: inst = 32'd201344662;
      8592: inst = 32'd203484854;
      8593: inst = 32'd471859200;
      8594: inst = 32'd136314880;
      8595: inst = 32'd268468224;
      8596: inst = 32'd201344663;
      8597: inst = 32'd203484854;
      8598: inst = 32'd471859200;
      8599: inst = 32'd136314880;
      8600: inst = 32'd268468224;
      8601: inst = 32'd201344664;
      8602: inst = 32'd203484854;
      8603: inst = 32'd471859200;
      8604: inst = 32'd136314880;
      8605: inst = 32'd268468224;
      8606: inst = 32'd201344665;
      8607: inst = 32'd203484854;
      8608: inst = 32'd471859200;
      8609: inst = 32'd136314880;
      8610: inst = 32'd268468224;
      8611: inst = 32'd201344666;
      8612: inst = 32'd203484854;
      8613: inst = 32'd471859200;
      8614: inst = 32'd136314880;
      8615: inst = 32'd268468224;
      8616: inst = 32'd201344667;
      8617: inst = 32'd203484854;
      8618: inst = 32'd471859200;
      8619: inst = 32'd136314880;
      8620: inst = 32'd268468224;
      8621: inst = 32'd201344668;
      8622: inst = 32'd203484854;
      8623: inst = 32'd471859200;
      8624: inst = 32'd136314880;
      8625: inst = 32'd268468224;
      8626: inst = 32'd201344669;
      8627: inst = 32'd203484854;
      8628: inst = 32'd471859200;
      8629: inst = 32'd136314880;
      8630: inst = 32'd268468224;
      8631: inst = 32'd201344670;
      8632: inst = 32'd203484854;
      8633: inst = 32'd471859200;
      8634: inst = 32'd136314880;
      8635: inst = 32'd268468224;
      8636: inst = 32'd201344671;
      8637: inst = 32'd203484854;
      8638: inst = 32'd471859200;
      8639: inst = 32'd136314880;
      8640: inst = 32'd268468224;
      8641: inst = 32'd201344672;
      8642: inst = 32'd203484854;
      8643: inst = 32'd471859200;
      8644: inst = 32'd136314880;
      8645: inst = 32'd268468224;
      8646: inst = 32'd201344673;
      8647: inst = 32'd203484854;
      8648: inst = 32'd471859200;
      8649: inst = 32'd136314880;
      8650: inst = 32'd268468224;
      8651: inst = 32'd201344674;
      8652: inst = 32'd203484854;
      8653: inst = 32'd471859200;
      8654: inst = 32'd136314880;
      8655: inst = 32'd268468224;
      8656: inst = 32'd201344675;
      8657: inst = 32'd203484854;
      8658: inst = 32'd471859200;
      8659: inst = 32'd136314880;
      8660: inst = 32'd268468224;
      8661: inst = 32'd201344676;
      8662: inst = 32'd203484854;
      8663: inst = 32'd471859200;
      8664: inst = 32'd136314880;
      8665: inst = 32'd268468224;
      8666: inst = 32'd201344677;
      8667: inst = 32'd203484854;
      8668: inst = 32'd471859200;
      8669: inst = 32'd136314880;
      8670: inst = 32'd268468224;
      8671: inst = 32'd201344678;
      8672: inst = 32'd203484854;
      8673: inst = 32'd471859200;
      8674: inst = 32'd136314880;
      8675: inst = 32'd268468224;
      8676: inst = 32'd201344679;
      8677: inst = 32'd203484854;
      8678: inst = 32'd471859200;
      8679: inst = 32'd136314880;
      8680: inst = 32'd268468224;
      8681: inst = 32'd201344680;
      8682: inst = 32'd203484854;
      8683: inst = 32'd471859200;
      8684: inst = 32'd136314880;
      8685: inst = 32'd268468224;
      8686: inst = 32'd201344681;
      8687: inst = 32'd203484854;
      8688: inst = 32'd471859200;
      8689: inst = 32'd136314880;
      8690: inst = 32'd268468224;
      8691: inst = 32'd201344682;
      8692: inst = 32'd203484854;
      8693: inst = 32'd471859200;
      8694: inst = 32'd136314880;
      8695: inst = 32'd268468224;
      8696: inst = 32'd201344683;
      8697: inst = 32'd203484854;
      8698: inst = 32'd471859200;
      8699: inst = 32'd136314880;
      8700: inst = 32'd268468224;
      8701: inst = 32'd201344684;
      8702: inst = 32'd203484854;
      8703: inst = 32'd471859200;
      8704: inst = 32'd136314880;
      8705: inst = 32'd268468224;
      8706: inst = 32'd201344685;
      8707: inst = 32'd203484854;
      8708: inst = 32'd471859200;
      8709: inst = 32'd136314880;
      8710: inst = 32'd268468224;
      8711: inst = 32'd201344686;
      8712: inst = 32'd203484854;
      8713: inst = 32'd471859200;
      8714: inst = 32'd136314880;
      8715: inst = 32'd268468224;
      8716: inst = 32'd201344687;
      8717: inst = 32'd203484854;
      8718: inst = 32'd471859200;
      8719: inst = 32'd136314880;
      8720: inst = 32'd268468224;
      8721: inst = 32'd201344688;
      8722: inst = 32'd203484854;
      8723: inst = 32'd471859200;
      8724: inst = 32'd136314880;
      8725: inst = 32'd268468224;
      8726: inst = 32'd201344689;
      8727: inst = 32'd203484854;
      8728: inst = 32'd471859200;
      8729: inst = 32'd136314880;
      8730: inst = 32'd268468224;
      8731: inst = 32'd201344690;
      8732: inst = 32'd203484854;
      8733: inst = 32'd471859200;
      8734: inst = 32'd136314880;
      8735: inst = 32'd268468224;
      8736: inst = 32'd201344691;
      8737: inst = 32'd203484854;
      8738: inst = 32'd471859200;
      8739: inst = 32'd136314880;
      8740: inst = 32'd268468224;
      8741: inst = 32'd201344692;
      8742: inst = 32'd203484854;
      8743: inst = 32'd471859200;
      8744: inst = 32'd136314880;
      8745: inst = 32'd268468224;
      8746: inst = 32'd201344693;
      8747: inst = 32'd203484854;
      8748: inst = 32'd471859200;
      8749: inst = 32'd136314880;
      8750: inst = 32'd268468224;
      8751: inst = 32'd201344694;
      8752: inst = 32'd203484854;
      8753: inst = 32'd471859200;
      8754: inst = 32'd136314880;
      8755: inst = 32'd268468224;
      8756: inst = 32'd201344695;
      8757: inst = 32'd203484854;
      8758: inst = 32'd471859200;
      8759: inst = 32'd136314880;
      8760: inst = 32'd268468224;
      8761: inst = 32'd201344696;
      8762: inst = 32'd203484854;
      8763: inst = 32'd471859200;
      8764: inst = 32'd136314880;
      8765: inst = 32'd268468224;
      8766: inst = 32'd201344697;
      8767: inst = 32'd203484854;
      8768: inst = 32'd471859200;
      8769: inst = 32'd136314880;
      8770: inst = 32'd268468224;
      8771: inst = 32'd201344698;
      8772: inst = 32'd203484854;
      8773: inst = 32'd471859200;
      8774: inst = 32'd136314880;
      8775: inst = 32'd268468224;
      8776: inst = 32'd201344699;
      8777: inst = 32'd203484854;
      8778: inst = 32'd471859200;
      8779: inst = 32'd136314880;
      8780: inst = 32'd268468224;
      8781: inst = 32'd201344700;
      8782: inst = 32'd203489279;
      8783: inst = 32'd471859200;
      8784: inst = 32'd136314880;
      8785: inst = 32'd268468224;
      8786: inst = 32'd201344701;
      8787: inst = 32'd203489279;
      8788: inst = 32'd471859200;
      8789: inst = 32'd136314880;
      8790: inst = 32'd268468224;
      8791: inst = 32'd201344702;
      8792: inst = 32'd203489279;
      8793: inst = 32'd471859200;
      8794: inst = 32'd136314880;
      8795: inst = 32'd268468224;
      8796: inst = 32'd201344703;
      8797: inst = 32'd203489279;
      8798: inst = 32'd471859200;
      8799: inst = 32'd136314880;
      8800: inst = 32'd268468224;
      8801: inst = 32'd201344704;
      8802: inst = 32'd203489279;
      8803: inst = 32'd471859200;
      8804: inst = 32'd136314880;
      8805: inst = 32'd268468224;
      8806: inst = 32'd201344705;
      8807: inst = 32'd203489279;
      8808: inst = 32'd471859200;
      8809: inst = 32'd136314880;
      8810: inst = 32'd268468224;
      8811: inst = 32'd201344706;
      8812: inst = 32'd203489279;
      8813: inst = 32'd471859200;
      8814: inst = 32'd136314880;
      8815: inst = 32'd268468224;
      8816: inst = 32'd201344707;
      8817: inst = 32'd203489279;
      8818: inst = 32'd471859200;
      8819: inst = 32'd136314880;
      8820: inst = 32'd268468224;
      8821: inst = 32'd201344708;
      8822: inst = 32'd203489279;
      8823: inst = 32'd471859200;
      8824: inst = 32'd136314880;
      8825: inst = 32'd268468224;
      8826: inst = 32'd201344709;
      8827: inst = 32'd203489279;
      8828: inst = 32'd471859200;
      8829: inst = 32'd136314880;
      8830: inst = 32'd268468224;
      8831: inst = 32'd201344710;
      8832: inst = 32'd203489279;
      8833: inst = 32'd471859200;
      8834: inst = 32'd136314880;
      8835: inst = 32'd268468224;
      8836: inst = 32'd201344711;
      8837: inst = 32'd203489279;
      8838: inst = 32'd471859200;
      8839: inst = 32'd136314880;
      8840: inst = 32'd268468224;
      8841: inst = 32'd201344712;
      8842: inst = 32'd203489279;
      8843: inst = 32'd471859200;
      8844: inst = 32'd136314880;
      8845: inst = 32'd268468224;
      8846: inst = 32'd201344713;
      8847: inst = 32'd203489279;
      8848: inst = 32'd471859200;
      8849: inst = 32'd136314880;
      8850: inst = 32'd268468224;
      8851: inst = 32'd201344714;
      8852: inst = 32'd203489279;
      8853: inst = 32'd471859200;
      8854: inst = 32'd136314880;
      8855: inst = 32'd268468224;
      8856: inst = 32'd201344715;
      8857: inst = 32'd203489279;
      8858: inst = 32'd471859200;
      8859: inst = 32'd136314880;
      8860: inst = 32'd268468224;
      8861: inst = 32'd201344716;
      8862: inst = 32'd203489279;
      8863: inst = 32'd471859200;
      8864: inst = 32'd136314880;
      8865: inst = 32'd268468224;
      8866: inst = 32'd201344717;
      8867: inst = 32'd203489279;
      8868: inst = 32'd471859200;
      8869: inst = 32'd136314880;
      8870: inst = 32'd268468224;
      8871: inst = 32'd201344718;
      8872: inst = 32'd203489279;
      8873: inst = 32'd471859200;
      8874: inst = 32'd136314880;
      8875: inst = 32'd268468224;
      8876: inst = 32'd201344719;
      8877: inst = 32'd203489279;
      8878: inst = 32'd471859200;
      8879: inst = 32'd136314880;
      8880: inst = 32'd268468224;
      8881: inst = 32'd201344720;
      8882: inst = 32'd203489279;
      8883: inst = 32'd471859200;
      8884: inst = 32'd136314880;
      8885: inst = 32'd268468224;
      8886: inst = 32'd201344721;
      8887: inst = 32'd203489279;
      8888: inst = 32'd471859200;
      8889: inst = 32'd136314880;
      8890: inst = 32'd268468224;
      8891: inst = 32'd201344722;
      8892: inst = 32'd203489279;
      8893: inst = 32'd471859200;
      8894: inst = 32'd136314880;
      8895: inst = 32'd268468224;
      8896: inst = 32'd201344723;
      8897: inst = 32'd203489279;
      8898: inst = 32'd471859200;
      8899: inst = 32'd136314880;
      8900: inst = 32'd268468224;
      8901: inst = 32'd201344724;
      8902: inst = 32'd203489279;
      8903: inst = 32'd471859200;
      8904: inst = 32'd136314880;
      8905: inst = 32'd268468224;
      8906: inst = 32'd201344725;
      8907: inst = 32'd203489279;
      8908: inst = 32'd471859200;
      8909: inst = 32'd136314880;
      8910: inst = 32'd268468224;
      8911: inst = 32'd201344726;
      8912: inst = 32'd203489279;
      8913: inst = 32'd471859200;
      8914: inst = 32'd136314880;
      8915: inst = 32'd268468224;
      8916: inst = 32'd201344727;
      8917: inst = 32'd203489279;
      8918: inst = 32'd471859200;
      8919: inst = 32'd136314880;
      8920: inst = 32'd268468224;
      8921: inst = 32'd201344728;
      8922: inst = 32'd203489279;
      8923: inst = 32'd471859200;
      8924: inst = 32'd136314880;
      8925: inst = 32'd268468224;
      8926: inst = 32'd201344729;
      8927: inst = 32'd203489279;
      8928: inst = 32'd471859200;
      8929: inst = 32'd136314880;
      8930: inst = 32'd268468224;
      8931: inst = 32'd201344730;
      8932: inst = 32'd203489279;
      8933: inst = 32'd471859200;
      8934: inst = 32'd136314880;
      8935: inst = 32'd268468224;
      8936: inst = 32'd201344731;
      8937: inst = 32'd203489279;
      8938: inst = 32'd471859200;
      8939: inst = 32'd136314880;
      8940: inst = 32'd268468224;
      8941: inst = 32'd201344732;
      8942: inst = 32'd203489279;
      8943: inst = 32'd471859200;
      8944: inst = 32'd136314880;
      8945: inst = 32'd268468224;
      8946: inst = 32'd201344733;
      8947: inst = 32'd203489279;
      8948: inst = 32'd471859200;
      8949: inst = 32'd136314880;
      8950: inst = 32'd268468224;
      8951: inst = 32'd201344734;
      8952: inst = 32'd203489279;
      8953: inst = 32'd471859200;
      8954: inst = 32'd136314880;
      8955: inst = 32'd268468224;
      8956: inst = 32'd201344735;
      8957: inst = 32'd203489279;
      8958: inst = 32'd471859200;
      8959: inst = 32'd136314880;
      8960: inst = 32'd268468224;
      8961: inst = 32'd201344736;
      8962: inst = 32'd203489279;
      8963: inst = 32'd471859200;
      8964: inst = 32'd136314880;
      8965: inst = 32'd268468224;
      8966: inst = 32'd201344737;
      8967: inst = 32'd203489279;
      8968: inst = 32'd471859200;
      8969: inst = 32'd136314880;
      8970: inst = 32'd268468224;
      8971: inst = 32'd201344738;
      8972: inst = 32'd203489279;
      8973: inst = 32'd471859200;
      8974: inst = 32'd136314880;
      8975: inst = 32'd268468224;
      8976: inst = 32'd201344739;
      8977: inst = 32'd203489279;
      8978: inst = 32'd471859200;
      8979: inst = 32'd136314880;
      8980: inst = 32'd268468224;
      8981: inst = 32'd201344740;
      8982: inst = 32'd203484854;
      8983: inst = 32'd471859200;
      8984: inst = 32'd136314880;
      8985: inst = 32'd268468224;
      8986: inst = 32'd201344741;
      8987: inst = 32'd203484854;
      8988: inst = 32'd471859200;
      8989: inst = 32'd136314880;
      8990: inst = 32'd268468224;
      8991: inst = 32'd201344742;
      8992: inst = 32'd203484854;
      8993: inst = 32'd471859200;
      8994: inst = 32'd136314880;
      8995: inst = 32'd268468224;
      8996: inst = 32'd201344743;
      8997: inst = 32'd203484854;
      8998: inst = 32'd471859200;
      8999: inst = 32'd136314880;
      9000: inst = 32'd268468224;
      9001: inst = 32'd201344744;
      9002: inst = 32'd203484854;
      9003: inst = 32'd471859200;
      9004: inst = 32'd136314880;
      9005: inst = 32'd268468224;
      9006: inst = 32'd201344745;
      9007: inst = 32'd203484854;
      9008: inst = 32'd471859200;
      9009: inst = 32'd136314880;
      9010: inst = 32'd268468224;
      9011: inst = 32'd201344746;
      9012: inst = 32'd203484854;
      9013: inst = 32'd471859200;
      9014: inst = 32'd136314880;
      9015: inst = 32'd268468224;
      9016: inst = 32'd201344747;
      9017: inst = 32'd203484854;
      9018: inst = 32'd471859200;
      9019: inst = 32'd136314880;
      9020: inst = 32'd268468224;
      9021: inst = 32'd201344748;
      9022: inst = 32'd203484854;
      9023: inst = 32'd471859200;
      9024: inst = 32'd136314880;
      9025: inst = 32'd268468224;
      9026: inst = 32'd201344749;
      9027: inst = 32'd203484854;
      9028: inst = 32'd471859200;
      9029: inst = 32'd136314880;
      9030: inst = 32'd268468224;
      9031: inst = 32'd201344750;
      9032: inst = 32'd203484854;
      9033: inst = 32'd471859200;
      9034: inst = 32'd136314880;
      9035: inst = 32'd268468224;
      9036: inst = 32'd201344751;
      9037: inst = 32'd203473634;
      9038: inst = 32'd471859200;
      9039: inst = 32'd136314880;
      9040: inst = 32'd268468224;
      9041: inst = 32'd201344752;
      9042: inst = 32'd203473634;
      9043: inst = 32'd471859200;
      9044: inst = 32'd136314880;
      9045: inst = 32'd268468224;
      9046: inst = 32'd201344753;
      9047: inst = 32'd203473634;
      9048: inst = 32'd471859200;
      9049: inst = 32'd136314880;
      9050: inst = 32'd268468224;
      9051: inst = 32'd201344754;
      9052: inst = 32'd203473634;
      9053: inst = 32'd471859200;
      9054: inst = 32'd136314880;
      9055: inst = 32'd268468224;
      9056: inst = 32'd201344755;
      9057: inst = 32'd203473634;
      9058: inst = 32'd471859200;
      9059: inst = 32'd136314880;
      9060: inst = 32'd268468224;
      9061: inst = 32'd201344756;
      9062: inst = 32'd203473634;
      9063: inst = 32'd471859200;
      9064: inst = 32'd136314880;
      9065: inst = 32'd268468224;
      9066: inst = 32'd201344757;
      9067: inst = 32'd203473634;
      9068: inst = 32'd471859200;
      9069: inst = 32'd136314880;
      9070: inst = 32'd268468224;
      9071: inst = 32'd201344758;
      9072: inst = 32'd203473634;
      9073: inst = 32'd471859200;
      9074: inst = 32'd136314880;
      9075: inst = 32'd268468224;
      9076: inst = 32'd201344759;
      9077: inst = 32'd203473634;
      9078: inst = 32'd471859200;
      9079: inst = 32'd136314880;
      9080: inst = 32'd268468224;
      9081: inst = 32'd201344760;
      9082: inst = 32'd203473634;
      9083: inst = 32'd471859200;
      9084: inst = 32'd136314880;
      9085: inst = 32'd268468224;
      9086: inst = 32'd201344761;
      9087: inst = 32'd203473634;
      9088: inst = 32'd471859200;
      9089: inst = 32'd136314880;
      9090: inst = 32'd268468224;
      9091: inst = 32'd201344762;
      9092: inst = 32'd203473634;
      9093: inst = 32'd471859200;
      9094: inst = 32'd136314880;
      9095: inst = 32'd268468224;
      9096: inst = 32'd201344763;
      9097: inst = 32'd203473634;
      9098: inst = 32'd471859200;
      9099: inst = 32'd136314880;
      9100: inst = 32'd268468224;
      9101: inst = 32'd201344764;
      9102: inst = 32'd203473634;
      9103: inst = 32'd471859200;
      9104: inst = 32'd136314880;
      9105: inst = 32'd268468224;
      9106: inst = 32'd201344765;
      9107: inst = 32'd203473634;
      9108: inst = 32'd471859200;
      9109: inst = 32'd136314880;
      9110: inst = 32'd268468224;
      9111: inst = 32'd201344766;
      9112: inst = 32'd203473634;
      9113: inst = 32'd471859200;
      9114: inst = 32'd136314880;
      9115: inst = 32'd268468224;
      9116: inst = 32'd201344767;
      9117: inst = 32'd203473634;
      9118: inst = 32'd471859200;
      9119: inst = 32'd136314880;
      9120: inst = 32'd268468224;
      9121: inst = 32'd201344768;
      9122: inst = 32'd203484854;
      9123: inst = 32'd471859200;
      9124: inst = 32'd136314880;
      9125: inst = 32'd268468224;
      9126: inst = 32'd201344769;
      9127: inst = 32'd203484854;
      9128: inst = 32'd471859200;
      9129: inst = 32'd136314880;
      9130: inst = 32'd268468224;
      9131: inst = 32'd201344770;
      9132: inst = 32'd203484854;
      9133: inst = 32'd471859200;
      9134: inst = 32'd136314880;
      9135: inst = 32'd268468224;
      9136: inst = 32'd201344771;
      9137: inst = 32'd203484854;
      9138: inst = 32'd471859200;
      9139: inst = 32'd136314880;
      9140: inst = 32'd268468224;
      9141: inst = 32'd201344772;
      9142: inst = 32'd203484854;
      9143: inst = 32'd471859200;
      9144: inst = 32'd136314880;
      9145: inst = 32'd268468224;
      9146: inst = 32'd201344773;
      9147: inst = 32'd203484854;
      9148: inst = 32'd471859200;
      9149: inst = 32'd136314880;
      9150: inst = 32'd268468224;
      9151: inst = 32'd201344774;
      9152: inst = 32'd203484854;
      9153: inst = 32'd471859200;
      9154: inst = 32'd136314880;
      9155: inst = 32'd268468224;
      9156: inst = 32'd201344775;
      9157: inst = 32'd203484854;
      9158: inst = 32'd471859200;
      9159: inst = 32'd136314880;
      9160: inst = 32'd268468224;
      9161: inst = 32'd201344776;
      9162: inst = 32'd203484854;
      9163: inst = 32'd471859200;
      9164: inst = 32'd136314880;
      9165: inst = 32'd268468224;
      9166: inst = 32'd201344777;
      9167: inst = 32'd203484854;
      9168: inst = 32'd471859200;
      9169: inst = 32'd136314880;
      9170: inst = 32'd268468224;
      9171: inst = 32'd201344778;
      9172: inst = 32'd203484854;
      9173: inst = 32'd471859200;
      9174: inst = 32'd136314880;
      9175: inst = 32'd268468224;
      9176: inst = 32'd201344779;
      9177: inst = 32'd203484854;
      9178: inst = 32'd471859200;
      9179: inst = 32'd136314880;
      9180: inst = 32'd268468224;
      9181: inst = 32'd201344780;
      9182: inst = 32'd203484854;
      9183: inst = 32'd471859200;
      9184: inst = 32'd136314880;
      9185: inst = 32'd268468224;
      9186: inst = 32'd201344781;
      9187: inst = 32'd203484854;
      9188: inst = 32'd471859200;
      9189: inst = 32'd136314880;
      9190: inst = 32'd268468224;
      9191: inst = 32'd201344782;
      9192: inst = 32'd203484854;
      9193: inst = 32'd471859200;
      9194: inst = 32'd136314880;
      9195: inst = 32'd268468224;
      9196: inst = 32'd201344783;
      9197: inst = 32'd203484854;
      9198: inst = 32'd471859200;
      9199: inst = 32'd136314880;
      9200: inst = 32'd268468224;
      9201: inst = 32'd201344784;
      9202: inst = 32'd203484854;
      9203: inst = 32'd471859200;
      9204: inst = 32'd136314880;
      9205: inst = 32'd268468224;
      9206: inst = 32'd201344785;
      9207: inst = 32'd203484854;
      9208: inst = 32'd471859200;
      9209: inst = 32'd136314880;
      9210: inst = 32'd268468224;
      9211: inst = 32'd201344786;
      9212: inst = 32'd203484854;
      9213: inst = 32'd471859200;
      9214: inst = 32'd136314880;
      9215: inst = 32'd268468224;
      9216: inst = 32'd201344787;
      9217: inst = 32'd203484854;
      9218: inst = 32'd471859200;
      9219: inst = 32'd136314880;
      9220: inst = 32'd268468224;
      9221: inst = 32'd201344788;
      9222: inst = 32'd203484854;
      9223: inst = 32'd471859200;
      9224: inst = 32'd136314880;
      9225: inst = 32'd268468224;
      9226: inst = 32'd201344789;
      9227: inst = 32'd203484854;
      9228: inst = 32'd471859200;
      9229: inst = 32'd136314880;
      9230: inst = 32'd268468224;
      9231: inst = 32'd201344790;
      9232: inst = 32'd203484854;
      9233: inst = 32'd471859200;
      9234: inst = 32'd136314880;
      9235: inst = 32'd268468224;
      9236: inst = 32'd201344791;
      9237: inst = 32'd203484854;
      9238: inst = 32'd471859200;
      9239: inst = 32'd136314880;
      9240: inst = 32'd268468224;
      9241: inst = 32'd201344792;
      9242: inst = 32'd203484854;
      9243: inst = 32'd471859200;
      9244: inst = 32'd136314880;
      9245: inst = 32'd268468224;
      9246: inst = 32'd201344793;
      9247: inst = 32'd203484854;
      9248: inst = 32'd471859200;
      9249: inst = 32'd136314880;
      9250: inst = 32'd268468224;
      9251: inst = 32'd201344794;
      9252: inst = 32'd203484854;
      9253: inst = 32'd471859200;
      9254: inst = 32'd136314880;
      9255: inst = 32'd268468224;
      9256: inst = 32'd201344795;
      9257: inst = 32'd203484854;
      9258: inst = 32'd471859200;
      9259: inst = 32'd136314880;
      9260: inst = 32'd268468224;
      9261: inst = 32'd201344796;
      9262: inst = 32'd203489279;
      9263: inst = 32'd471859200;
      9264: inst = 32'd136314880;
      9265: inst = 32'd268468224;
      9266: inst = 32'd201344797;
      9267: inst = 32'd203489279;
      9268: inst = 32'd471859200;
      9269: inst = 32'd136314880;
      9270: inst = 32'd268468224;
      9271: inst = 32'd201344798;
      9272: inst = 32'd203489279;
      9273: inst = 32'd471859200;
      9274: inst = 32'd136314880;
      9275: inst = 32'd268468224;
      9276: inst = 32'd201344799;
      9277: inst = 32'd203489279;
      9278: inst = 32'd471859200;
      9279: inst = 32'd136314880;
      9280: inst = 32'd268468224;
      9281: inst = 32'd201344800;
      9282: inst = 32'd203489279;
      9283: inst = 32'd471859200;
      9284: inst = 32'd136314880;
      9285: inst = 32'd268468224;
      9286: inst = 32'd201344801;
      9287: inst = 32'd203489279;
      9288: inst = 32'd471859200;
      9289: inst = 32'd136314880;
      9290: inst = 32'd268468224;
      9291: inst = 32'd201344802;
      9292: inst = 32'd203489279;
      9293: inst = 32'd471859200;
      9294: inst = 32'd136314880;
      9295: inst = 32'd268468224;
      9296: inst = 32'd201344803;
      9297: inst = 32'd203489279;
      9298: inst = 32'd471859200;
      9299: inst = 32'd136314880;
      9300: inst = 32'd268468224;
      9301: inst = 32'd201344804;
      9302: inst = 32'd203489279;
      9303: inst = 32'd471859200;
      9304: inst = 32'd136314880;
      9305: inst = 32'd268468224;
      9306: inst = 32'd201344805;
      9307: inst = 32'd203489279;
      9308: inst = 32'd471859200;
      9309: inst = 32'd136314880;
      9310: inst = 32'd268468224;
      9311: inst = 32'd201344806;
      9312: inst = 32'd203489279;
      9313: inst = 32'd471859200;
      9314: inst = 32'd136314880;
      9315: inst = 32'd268468224;
      9316: inst = 32'd201344807;
      9317: inst = 32'd203489279;
      9318: inst = 32'd471859200;
      9319: inst = 32'd136314880;
      9320: inst = 32'd268468224;
      9321: inst = 32'd201344808;
      9322: inst = 32'd203489279;
      9323: inst = 32'd471859200;
      9324: inst = 32'd136314880;
      9325: inst = 32'd268468224;
      9326: inst = 32'd201344809;
      9327: inst = 32'd203489279;
      9328: inst = 32'd471859200;
      9329: inst = 32'd136314880;
      9330: inst = 32'd268468224;
      9331: inst = 32'd201344810;
      9332: inst = 32'd203489279;
      9333: inst = 32'd471859200;
      9334: inst = 32'd136314880;
      9335: inst = 32'd268468224;
      9336: inst = 32'd201344811;
      9337: inst = 32'd203489279;
      9338: inst = 32'd471859200;
      9339: inst = 32'd136314880;
      9340: inst = 32'd268468224;
      9341: inst = 32'd201344812;
      9342: inst = 32'd203489279;
      9343: inst = 32'd471859200;
      9344: inst = 32'd136314880;
      9345: inst = 32'd268468224;
      9346: inst = 32'd201344813;
      9347: inst = 32'd203489279;
      9348: inst = 32'd471859200;
      9349: inst = 32'd136314880;
      9350: inst = 32'd268468224;
      9351: inst = 32'd201344814;
      9352: inst = 32'd203489279;
      9353: inst = 32'd471859200;
      9354: inst = 32'd136314880;
      9355: inst = 32'd268468224;
      9356: inst = 32'd201344815;
      9357: inst = 32'd203489279;
      9358: inst = 32'd471859200;
      9359: inst = 32'd136314880;
      9360: inst = 32'd268468224;
      9361: inst = 32'd201344816;
      9362: inst = 32'd203489279;
      9363: inst = 32'd471859200;
      9364: inst = 32'd136314880;
      9365: inst = 32'd268468224;
      9366: inst = 32'd201344817;
      9367: inst = 32'd203489279;
      9368: inst = 32'd471859200;
      9369: inst = 32'd136314880;
      9370: inst = 32'd268468224;
      9371: inst = 32'd201344818;
      9372: inst = 32'd203489279;
      9373: inst = 32'd471859200;
      9374: inst = 32'd136314880;
      9375: inst = 32'd268468224;
      9376: inst = 32'd201344819;
      9377: inst = 32'd203489279;
      9378: inst = 32'd471859200;
      9379: inst = 32'd136314880;
      9380: inst = 32'd268468224;
      9381: inst = 32'd201344820;
      9382: inst = 32'd203489279;
      9383: inst = 32'd471859200;
      9384: inst = 32'd136314880;
      9385: inst = 32'd268468224;
      9386: inst = 32'd201344821;
      9387: inst = 32'd203489279;
      9388: inst = 32'd471859200;
      9389: inst = 32'd136314880;
      9390: inst = 32'd268468224;
      9391: inst = 32'd201344822;
      9392: inst = 32'd203489279;
      9393: inst = 32'd471859200;
      9394: inst = 32'd136314880;
      9395: inst = 32'd268468224;
      9396: inst = 32'd201344823;
      9397: inst = 32'd203489279;
      9398: inst = 32'd471859200;
      9399: inst = 32'd136314880;
      9400: inst = 32'd268468224;
      9401: inst = 32'd201344824;
      9402: inst = 32'd203489279;
      9403: inst = 32'd471859200;
      9404: inst = 32'd136314880;
      9405: inst = 32'd268468224;
      9406: inst = 32'd201344825;
      9407: inst = 32'd203489279;
      9408: inst = 32'd471859200;
      9409: inst = 32'd136314880;
      9410: inst = 32'd268468224;
      9411: inst = 32'd201344826;
      9412: inst = 32'd203489279;
      9413: inst = 32'd471859200;
      9414: inst = 32'd136314880;
      9415: inst = 32'd268468224;
      9416: inst = 32'd201344827;
      9417: inst = 32'd203489279;
      9418: inst = 32'd471859200;
      9419: inst = 32'd136314880;
      9420: inst = 32'd268468224;
      9421: inst = 32'd201344828;
      9422: inst = 32'd203489279;
      9423: inst = 32'd471859200;
      9424: inst = 32'd136314880;
      9425: inst = 32'd268468224;
      9426: inst = 32'd201344829;
      9427: inst = 32'd203489279;
      9428: inst = 32'd471859200;
      9429: inst = 32'd136314880;
      9430: inst = 32'd268468224;
      9431: inst = 32'd201344830;
      9432: inst = 32'd203489279;
      9433: inst = 32'd471859200;
      9434: inst = 32'd136314880;
      9435: inst = 32'd268468224;
      9436: inst = 32'd201344831;
      9437: inst = 32'd203489279;
      9438: inst = 32'd471859200;
      9439: inst = 32'd136314880;
      9440: inst = 32'd268468224;
      9441: inst = 32'd201344832;
      9442: inst = 32'd203489279;
      9443: inst = 32'd471859200;
      9444: inst = 32'd136314880;
      9445: inst = 32'd268468224;
      9446: inst = 32'd201344833;
      9447: inst = 32'd203489279;
      9448: inst = 32'd471859200;
      9449: inst = 32'd136314880;
      9450: inst = 32'd268468224;
      9451: inst = 32'd201344834;
      9452: inst = 32'd203489279;
      9453: inst = 32'd471859200;
      9454: inst = 32'd136314880;
      9455: inst = 32'd268468224;
      9456: inst = 32'd201344835;
      9457: inst = 32'd203489279;
      9458: inst = 32'd471859200;
      9459: inst = 32'd136314880;
      9460: inst = 32'd268468224;
      9461: inst = 32'd201344836;
      9462: inst = 32'd203484854;
      9463: inst = 32'd471859200;
      9464: inst = 32'd136314880;
      9465: inst = 32'd268468224;
      9466: inst = 32'd201344837;
      9467: inst = 32'd203484854;
      9468: inst = 32'd471859200;
      9469: inst = 32'd136314880;
      9470: inst = 32'd268468224;
      9471: inst = 32'd201344838;
      9472: inst = 32'd203484854;
      9473: inst = 32'd471859200;
      9474: inst = 32'd136314880;
      9475: inst = 32'd268468224;
      9476: inst = 32'd201344839;
      9477: inst = 32'd203484854;
      9478: inst = 32'd471859200;
      9479: inst = 32'd136314880;
      9480: inst = 32'd268468224;
      9481: inst = 32'd201344840;
      9482: inst = 32'd203484854;
      9483: inst = 32'd471859200;
      9484: inst = 32'd136314880;
      9485: inst = 32'd268468224;
      9486: inst = 32'd201344841;
      9487: inst = 32'd203484854;
      9488: inst = 32'd471859200;
      9489: inst = 32'd136314880;
      9490: inst = 32'd268468224;
      9491: inst = 32'd201344842;
      9492: inst = 32'd203484854;
      9493: inst = 32'd471859200;
      9494: inst = 32'd136314880;
      9495: inst = 32'd268468224;
      9496: inst = 32'd201344843;
      9497: inst = 32'd203484854;
      9498: inst = 32'd471859200;
      9499: inst = 32'd136314880;
      9500: inst = 32'd268468224;
      9501: inst = 32'd201344844;
      9502: inst = 32'd203484854;
      9503: inst = 32'd471859200;
      9504: inst = 32'd136314880;
      9505: inst = 32'd268468224;
      9506: inst = 32'd201344845;
      9507: inst = 32'd203484854;
      9508: inst = 32'd471859200;
      9509: inst = 32'd136314880;
      9510: inst = 32'd268468224;
      9511: inst = 32'd201344846;
      9512: inst = 32'd203484854;
      9513: inst = 32'd471859200;
      9514: inst = 32'd136314880;
      9515: inst = 32'd268468224;
      9516: inst = 32'd201344847;
      9517: inst = 32'd203473634;
      9518: inst = 32'd471859200;
      9519: inst = 32'd136314880;
      9520: inst = 32'd268468224;
      9521: inst = 32'd201344848;
      9522: inst = 32'd203480005;
      9523: inst = 32'd471859200;
      9524: inst = 32'd136314880;
      9525: inst = 32'd268468224;
      9526: inst = 32'd201344849;
      9527: inst = 32'd203480005;
      9528: inst = 32'd471859200;
      9529: inst = 32'd136314880;
      9530: inst = 32'd268468224;
      9531: inst = 32'd201344850;
      9532: inst = 32'd203480005;
      9533: inst = 32'd471859200;
      9534: inst = 32'd136314880;
      9535: inst = 32'd268468224;
      9536: inst = 32'd201344851;
      9537: inst = 32'd203480005;
      9538: inst = 32'd471859200;
      9539: inst = 32'd136314880;
      9540: inst = 32'd268468224;
      9541: inst = 32'd201344852;
      9542: inst = 32'd203480005;
      9543: inst = 32'd471859200;
      9544: inst = 32'd136314880;
      9545: inst = 32'd268468224;
      9546: inst = 32'd201344853;
      9547: inst = 32'd203480005;
      9548: inst = 32'd471859200;
      9549: inst = 32'd136314880;
      9550: inst = 32'd268468224;
      9551: inst = 32'd201344854;
      9552: inst = 32'd203480005;
      9553: inst = 32'd471859200;
      9554: inst = 32'd136314880;
      9555: inst = 32'd268468224;
      9556: inst = 32'd201344855;
      9557: inst = 32'd203480005;
      9558: inst = 32'd471859200;
      9559: inst = 32'd136314880;
      9560: inst = 32'd268468224;
      9561: inst = 32'd201344856;
      9562: inst = 32'd203480005;
      9563: inst = 32'd471859200;
      9564: inst = 32'd136314880;
      9565: inst = 32'd268468224;
      9566: inst = 32'd201344857;
      9567: inst = 32'd203480005;
      9568: inst = 32'd471859200;
      9569: inst = 32'd136314880;
      9570: inst = 32'd268468224;
      9571: inst = 32'd201344858;
      9572: inst = 32'd203480005;
      9573: inst = 32'd471859200;
      9574: inst = 32'd136314880;
      9575: inst = 32'd268468224;
      9576: inst = 32'd201344859;
      9577: inst = 32'd203480005;
      9578: inst = 32'd471859200;
      9579: inst = 32'd136314880;
      9580: inst = 32'd268468224;
      9581: inst = 32'd201344860;
      9582: inst = 32'd203480005;
      9583: inst = 32'd471859200;
      9584: inst = 32'd136314880;
      9585: inst = 32'd268468224;
      9586: inst = 32'd201344861;
      9587: inst = 32'd203480005;
      9588: inst = 32'd471859200;
      9589: inst = 32'd136314880;
      9590: inst = 32'd268468224;
      9591: inst = 32'd201344862;
      9592: inst = 32'd203480005;
      9593: inst = 32'd471859200;
      9594: inst = 32'd136314880;
      9595: inst = 32'd268468224;
      9596: inst = 32'd201344863;
      9597: inst = 32'd203473634;
      9598: inst = 32'd471859200;
      9599: inst = 32'd136314880;
      9600: inst = 32'd268468224;
      9601: inst = 32'd201344864;
      9602: inst = 32'd203484854;
      9603: inst = 32'd471859200;
      9604: inst = 32'd136314880;
      9605: inst = 32'd268468224;
      9606: inst = 32'd201344865;
      9607: inst = 32'd203484854;
      9608: inst = 32'd471859200;
      9609: inst = 32'd136314880;
      9610: inst = 32'd268468224;
      9611: inst = 32'd201344866;
      9612: inst = 32'd203484854;
      9613: inst = 32'd471859200;
      9614: inst = 32'd136314880;
      9615: inst = 32'd268468224;
      9616: inst = 32'd201344867;
      9617: inst = 32'd203484854;
      9618: inst = 32'd471859200;
      9619: inst = 32'd136314880;
      9620: inst = 32'd268468224;
      9621: inst = 32'd201344868;
      9622: inst = 32'd203484854;
      9623: inst = 32'd471859200;
      9624: inst = 32'd136314880;
      9625: inst = 32'd268468224;
      9626: inst = 32'd201344869;
      9627: inst = 32'd203484854;
      9628: inst = 32'd471859200;
      9629: inst = 32'd136314880;
      9630: inst = 32'd268468224;
      9631: inst = 32'd201344870;
      9632: inst = 32'd203484854;
      9633: inst = 32'd471859200;
      9634: inst = 32'd136314880;
      9635: inst = 32'd268468224;
      9636: inst = 32'd201344871;
      9637: inst = 32'd203484854;
      9638: inst = 32'd471859200;
      9639: inst = 32'd136314880;
      9640: inst = 32'd268468224;
      9641: inst = 32'd201344872;
      9642: inst = 32'd203484854;
      9643: inst = 32'd471859200;
      9644: inst = 32'd136314880;
      9645: inst = 32'd268468224;
      9646: inst = 32'd201344873;
      9647: inst = 32'd203484854;
      9648: inst = 32'd471859200;
      9649: inst = 32'd136314880;
      9650: inst = 32'd268468224;
      9651: inst = 32'd201344874;
      9652: inst = 32'd203484854;
      9653: inst = 32'd471859200;
      9654: inst = 32'd136314880;
      9655: inst = 32'd268468224;
      9656: inst = 32'd201344875;
      9657: inst = 32'd203484854;
      9658: inst = 32'd471859200;
      9659: inst = 32'd136314880;
      9660: inst = 32'd268468224;
      9661: inst = 32'd201344876;
      9662: inst = 32'd203484854;
      9663: inst = 32'd471859200;
      9664: inst = 32'd136314880;
      9665: inst = 32'd268468224;
      9666: inst = 32'd201344877;
      9667: inst = 32'd203484854;
      9668: inst = 32'd471859200;
      9669: inst = 32'd136314880;
      9670: inst = 32'd268468224;
      9671: inst = 32'd201344878;
      9672: inst = 32'd203484854;
      9673: inst = 32'd471859200;
      9674: inst = 32'd136314880;
      9675: inst = 32'd268468224;
      9676: inst = 32'd201344879;
      9677: inst = 32'd203484854;
      9678: inst = 32'd471859200;
      9679: inst = 32'd136314880;
      9680: inst = 32'd268468224;
      9681: inst = 32'd201344880;
      9682: inst = 32'd203484854;
      9683: inst = 32'd471859200;
      9684: inst = 32'd136314880;
      9685: inst = 32'd268468224;
      9686: inst = 32'd201344881;
      9687: inst = 32'd203484854;
      9688: inst = 32'd471859200;
      9689: inst = 32'd136314880;
      9690: inst = 32'd268468224;
      9691: inst = 32'd201344882;
      9692: inst = 32'd203484854;
      9693: inst = 32'd471859200;
      9694: inst = 32'd136314880;
      9695: inst = 32'd268468224;
      9696: inst = 32'd201344883;
      9697: inst = 32'd203484854;
      9698: inst = 32'd471859200;
      9699: inst = 32'd136314880;
      9700: inst = 32'd268468224;
      9701: inst = 32'd201344884;
      9702: inst = 32'd203484854;
      9703: inst = 32'd471859200;
      9704: inst = 32'd136314880;
      9705: inst = 32'd268468224;
      9706: inst = 32'd201344885;
      9707: inst = 32'd203484854;
      9708: inst = 32'd471859200;
      9709: inst = 32'd136314880;
      9710: inst = 32'd268468224;
      9711: inst = 32'd201344886;
      9712: inst = 32'd203484854;
      9713: inst = 32'd471859200;
      9714: inst = 32'd136314880;
      9715: inst = 32'd268468224;
      9716: inst = 32'd201344887;
      9717: inst = 32'd203484854;
      9718: inst = 32'd471859200;
      9719: inst = 32'd136314880;
      9720: inst = 32'd268468224;
      9721: inst = 32'd201344888;
      9722: inst = 32'd203484854;
      9723: inst = 32'd471859200;
      9724: inst = 32'd136314880;
      9725: inst = 32'd268468224;
      9726: inst = 32'd201344889;
      9727: inst = 32'd203484854;
      9728: inst = 32'd471859200;
      9729: inst = 32'd136314880;
      9730: inst = 32'd268468224;
      9731: inst = 32'd201344890;
      9732: inst = 32'd203484854;
      9733: inst = 32'd471859200;
      9734: inst = 32'd136314880;
      9735: inst = 32'd268468224;
      9736: inst = 32'd201344891;
      9737: inst = 32'd203484854;
      9738: inst = 32'd471859200;
      9739: inst = 32'd136314880;
      9740: inst = 32'd268468224;
      9741: inst = 32'd201344892;
      9742: inst = 32'd203489279;
      9743: inst = 32'd471859200;
      9744: inst = 32'd136314880;
      9745: inst = 32'd268468224;
      9746: inst = 32'd201344893;
      9747: inst = 32'd203489279;
      9748: inst = 32'd471859200;
      9749: inst = 32'd136314880;
      9750: inst = 32'd268468224;
      9751: inst = 32'd201344894;
      9752: inst = 32'd203489279;
      9753: inst = 32'd471859200;
      9754: inst = 32'd136314880;
      9755: inst = 32'd268468224;
      9756: inst = 32'd201344895;
      9757: inst = 32'd203489279;
      9758: inst = 32'd471859200;
      9759: inst = 32'd136314880;
      9760: inst = 32'd268468224;
      9761: inst = 32'd201344896;
      9762: inst = 32'd203489279;
      9763: inst = 32'd471859200;
      9764: inst = 32'd136314880;
      9765: inst = 32'd268468224;
      9766: inst = 32'd201344897;
      9767: inst = 32'd203489279;
      9768: inst = 32'd471859200;
      9769: inst = 32'd136314880;
      9770: inst = 32'd268468224;
      9771: inst = 32'd201344898;
      9772: inst = 32'd203489279;
      9773: inst = 32'd471859200;
      9774: inst = 32'd136314880;
      9775: inst = 32'd268468224;
      9776: inst = 32'd201344899;
      9777: inst = 32'd203489279;
      9778: inst = 32'd471859200;
      9779: inst = 32'd136314880;
      9780: inst = 32'd268468224;
      9781: inst = 32'd201344900;
      9782: inst = 32'd203489279;
      9783: inst = 32'd471859200;
      9784: inst = 32'd136314880;
      9785: inst = 32'd268468224;
      9786: inst = 32'd201344901;
      9787: inst = 32'd203489279;
      9788: inst = 32'd471859200;
      9789: inst = 32'd136314880;
      9790: inst = 32'd268468224;
      9791: inst = 32'd201344902;
      9792: inst = 32'd203489279;
      9793: inst = 32'd471859200;
      9794: inst = 32'd136314880;
      9795: inst = 32'd268468224;
      9796: inst = 32'd201344903;
      9797: inst = 32'd203489279;
      9798: inst = 32'd471859200;
      9799: inst = 32'd136314880;
      9800: inst = 32'd268468224;
      9801: inst = 32'd201344904;
      9802: inst = 32'd203489279;
      9803: inst = 32'd471859200;
      9804: inst = 32'd136314880;
      9805: inst = 32'd268468224;
      9806: inst = 32'd201344905;
      9807: inst = 32'd203489279;
      9808: inst = 32'd471859200;
      9809: inst = 32'd136314880;
      9810: inst = 32'd268468224;
      9811: inst = 32'd201344906;
      9812: inst = 32'd203489279;
      9813: inst = 32'd471859200;
      9814: inst = 32'd136314880;
      9815: inst = 32'd268468224;
      9816: inst = 32'd201344907;
      9817: inst = 32'd203489279;
      9818: inst = 32'd471859200;
      9819: inst = 32'd136314880;
      9820: inst = 32'd268468224;
      9821: inst = 32'd201344908;
      9822: inst = 32'd203489279;
      9823: inst = 32'd471859200;
      9824: inst = 32'd136314880;
      9825: inst = 32'd268468224;
      9826: inst = 32'd201344909;
      9827: inst = 32'd203489279;
      9828: inst = 32'd471859200;
      9829: inst = 32'd136314880;
      9830: inst = 32'd268468224;
      9831: inst = 32'd201344910;
      9832: inst = 32'd203489279;
      9833: inst = 32'd471859200;
      9834: inst = 32'd136314880;
      9835: inst = 32'd268468224;
      9836: inst = 32'd201344911;
      9837: inst = 32'd203489279;
      9838: inst = 32'd471859200;
      9839: inst = 32'd136314880;
      9840: inst = 32'd268468224;
      9841: inst = 32'd201344912;
      9842: inst = 32'd203489279;
      9843: inst = 32'd471859200;
      9844: inst = 32'd136314880;
      9845: inst = 32'd268468224;
      9846: inst = 32'd201344913;
      9847: inst = 32'd203489279;
      9848: inst = 32'd471859200;
      9849: inst = 32'd136314880;
      9850: inst = 32'd268468224;
      9851: inst = 32'd201344914;
      9852: inst = 32'd203489279;
      9853: inst = 32'd471859200;
      9854: inst = 32'd136314880;
      9855: inst = 32'd268468224;
      9856: inst = 32'd201344915;
      9857: inst = 32'd203489279;
      9858: inst = 32'd471859200;
      9859: inst = 32'd136314880;
      9860: inst = 32'd268468224;
      9861: inst = 32'd201344916;
      9862: inst = 32'd203489279;
      9863: inst = 32'd471859200;
      9864: inst = 32'd136314880;
      9865: inst = 32'd268468224;
      9866: inst = 32'd201344917;
      9867: inst = 32'd203489279;
      9868: inst = 32'd471859200;
      9869: inst = 32'd136314880;
      9870: inst = 32'd268468224;
      9871: inst = 32'd201344918;
      9872: inst = 32'd203489279;
      9873: inst = 32'd471859200;
      9874: inst = 32'd136314880;
      9875: inst = 32'd268468224;
      9876: inst = 32'd201344919;
      9877: inst = 32'd203489279;
      9878: inst = 32'd471859200;
      9879: inst = 32'd136314880;
      9880: inst = 32'd268468224;
      9881: inst = 32'd201344920;
      9882: inst = 32'd203489279;
      9883: inst = 32'd471859200;
      9884: inst = 32'd136314880;
      9885: inst = 32'd268468224;
      9886: inst = 32'd201344921;
      9887: inst = 32'd203489279;
      9888: inst = 32'd471859200;
      9889: inst = 32'd136314880;
      9890: inst = 32'd268468224;
      9891: inst = 32'd201344922;
      9892: inst = 32'd203489279;
      9893: inst = 32'd471859200;
      9894: inst = 32'd136314880;
      9895: inst = 32'd268468224;
      9896: inst = 32'd201344923;
      9897: inst = 32'd203489279;
      9898: inst = 32'd471859200;
      9899: inst = 32'd136314880;
      9900: inst = 32'd268468224;
      9901: inst = 32'd201344924;
      9902: inst = 32'd203489279;
      9903: inst = 32'd471859200;
      9904: inst = 32'd136314880;
      9905: inst = 32'd268468224;
      9906: inst = 32'd201344925;
      9907: inst = 32'd203489279;
      9908: inst = 32'd471859200;
      9909: inst = 32'd136314880;
      9910: inst = 32'd268468224;
      9911: inst = 32'd201344926;
      9912: inst = 32'd203489279;
      9913: inst = 32'd471859200;
      9914: inst = 32'd136314880;
      9915: inst = 32'd268468224;
      9916: inst = 32'd201344927;
      9917: inst = 32'd203489279;
      9918: inst = 32'd471859200;
      9919: inst = 32'd136314880;
      9920: inst = 32'd268468224;
      9921: inst = 32'd201344928;
      9922: inst = 32'd203489279;
      9923: inst = 32'd471859200;
      9924: inst = 32'd136314880;
      9925: inst = 32'd268468224;
      9926: inst = 32'd201344929;
      9927: inst = 32'd203489279;
      9928: inst = 32'd471859200;
      9929: inst = 32'd136314880;
      9930: inst = 32'd268468224;
      9931: inst = 32'd201344930;
      9932: inst = 32'd203489279;
      9933: inst = 32'd471859200;
      9934: inst = 32'd136314880;
      9935: inst = 32'd268468224;
      9936: inst = 32'd201344931;
      9937: inst = 32'd203489279;
      9938: inst = 32'd471859200;
      9939: inst = 32'd136314880;
      9940: inst = 32'd268468224;
      9941: inst = 32'd201344932;
      9942: inst = 32'd203484854;
      9943: inst = 32'd471859200;
      9944: inst = 32'd136314880;
      9945: inst = 32'd268468224;
      9946: inst = 32'd201344933;
      9947: inst = 32'd203484854;
      9948: inst = 32'd471859200;
      9949: inst = 32'd136314880;
      9950: inst = 32'd268468224;
      9951: inst = 32'd201344934;
      9952: inst = 32'd203484854;
      9953: inst = 32'd471859200;
      9954: inst = 32'd136314880;
      9955: inst = 32'd268468224;
      9956: inst = 32'd201344935;
      9957: inst = 32'd203484854;
      9958: inst = 32'd471859200;
      9959: inst = 32'd136314880;
      9960: inst = 32'd268468224;
      9961: inst = 32'd201344936;
      9962: inst = 32'd203484854;
      9963: inst = 32'd471859200;
      9964: inst = 32'd136314880;
      9965: inst = 32'd268468224;
      9966: inst = 32'd201344937;
      9967: inst = 32'd203484854;
      9968: inst = 32'd471859200;
      9969: inst = 32'd136314880;
      9970: inst = 32'd268468224;
      9971: inst = 32'd201344938;
      9972: inst = 32'd203484854;
      9973: inst = 32'd471859200;
      9974: inst = 32'd136314880;
      9975: inst = 32'd268468224;
      9976: inst = 32'd201344939;
      9977: inst = 32'd203484854;
      9978: inst = 32'd471859200;
      9979: inst = 32'd136314880;
      9980: inst = 32'd268468224;
      9981: inst = 32'd201344940;
      9982: inst = 32'd203484854;
      9983: inst = 32'd471859200;
      9984: inst = 32'd136314880;
      9985: inst = 32'd268468224;
      9986: inst = 32'd201344941;
      9987: inst = 32'd203484854;
      9988: inst = 32'd471859200;
      9989: inst = 32'd136314880;
      9990: inst = 32'd268468224;
      9991: inst = 32'd201344942;
      9992: inst = 32'd203484854;
      9993: inst = 32'd471859200;
      9994: inst = 32'd136314880;
      9995: inst = 32'd268468224;
      9996: inst = 32'd201344943;
      9997: inst = 32'd203473634;
      9998: inst = 32'd471859200;
      9999: inst = 32'd136314880;
      10000: inst = 32'd268468224;
      10001: inst = 32'd201344944;
      10002: inst = 32'd203480005;
      10003: inst = 32'd471859200;
      10004: inst = 32'd136314880;
      10005: inst = 32'd268468224;
      10006: inst = 32'd201344945;
      10007: inst = 32'd203480005;
      10008: inst = 32'd471859200;
      10009: inst = 32'd136314880;
      10010: inst = 32'd268468224;
      10011: inst = 32'd201344946;
      10012: inst = 32'd203480005;
      10013: inst = 32'd471859200;
      10014: inst = 32'd136314880;
      10015: inst = 32'd268468224;
      10016: inst = 32'd201344947;
      10017: inst = 32'd203480005;
      10018: inst = 32'd471859200;
      10019: inst = 32'd136314880;
      10020: inst = 32'd268468224;
      10021: inst = 32'd201344948;
      10022: inst = 32'd203480005;
      10023: inst = 32'd471859200;
      10024: inst = 32'd136314880;
      10025: inst = 32'd268468224;
      10026: inst = 32'd201344949;
      10027: inst = 32'd203480005;
      10028: inst = 32'd471859200;
      10029: inst = 32'd136314880;
      10030: inst = 32'd268468224;
      10031: inst = 32'd201344950;
      10032: inst = 32'd203480005;
      10033: inst = 32'd471859200;
      10034: inst = 32'd136314880;
      10035: inst = 32'd268468224;
      10036: inst = 32'd201344951;
      10037: inst = 32'd203480005;
      10038: inst = 32'd471859200;
      10039: inst = 32'd136314880;
      10040: inst = 32'd268468224;
      10041: inst = 32'd201344952;
      10042: inst = 32'd203480005;
      10043: inst = 32'd471859200;
      10044: inst = 32'd136314880;
      10045: inst = 32'd268468224;
      10046: inst = 32'd201344953;
      10047: inst = 32'd203480005;
      10048: inst = 32'd471859200;
      10049: inst = 32'd136314880;
      10050: inst = 32'd268468224;
      10051: inst = 32'd201344954;
      10052: inst = 32'd203480005;
      10053: inst = 32'd471859200;
      10054: inst = 32'd136314880;
      10055: inst = 32'd268468224;
      10056: inst = 32'd201344955;
      10057: inst = 32'd203480005;
      10058: inst = 32'd471859200;
      10059: inst = 32'd136314880;
      10060: inst = 32'd268468224;
      10061: inst = 32'd201344956;
      10062: inst = 32'd203480005;
      10063: inst = 32'd471859200;
      10064: inst = 32'd136314880;
      10065: inst = 32'd268468224;
      10066: inst = 32'd201344957;
      10067: inst = 32'd203480005;
      10068: inst = 32'd471859200;
      10069: inst = 32'd136314880;
      10070: inst = 32'd268468224;
      10071: inst = 32'd201344958;
      10072: inst = 32'd203480005;
      10073: inst = 32'd471859200;
      10074: inst = 32'd136314880;
      10075: inst = 32'd268468224;
      10076: inst = 32'd201344959;
      10077: inst = 32'd203473634;
      10078: inst = 32'd471859200;
      10079: inst = 32'd136314880;
      10080: inst = 32'd268468224;
      10081: inst = 32'd201344960;
      10082: inst = 32'd203484854;
      10083: inst = 32'd471859200;
      10084: inst = 32'd136314880;
      10085: inst = 32'd268468224;
      10086: inst = 32'd201344961;
      10087: inst = 32'd203484854;
      10088: inst = 32'd471859200;
      10089: inst = 32'd136314880;
      10090: inst = 32'd268468224;
      10091: inst = 32'd201344962;
      10092: inst = 32'd203484854;
      10093: inst = 32'd471859200;
      10094: inst = 32'd136314880;
      10095: inst = 32'd268468224;
      10096: inst = 32'd201344963;
      10097: inst = 32'd203484854;
      10098: inst = 32'd471859200;
      10099: inst = 32'd136314880;
      10100: inst = 32'd268468224;
      10101: inst = 32'd201344964;
      10102: inst = 32'd203484854;
      10103: inst = 32'd471859200;
      10104: inst = 32'd136314880;
      10105: inst = 32'd268468224;
      10106: inst = 32'd201344965;
      10107: inst = 32'd203484854;
      10108: inst = 32'd471859200;
      10109: inst = 32'd136314880;
      10110: inst = 32'd268468224;
      10111: inst = 32'd201344966;
      10112: inst = 32'd203484854;
      10113: inst = 32'd471859200;
      10114: inst = 32'd136314880;
      10115: inst = 32'd268468224;
      10116: inst = 32'd201344967;
      10117: inst = 32'd203484854;
      10118: inst = 32'd471859200;
      10119: inst = 32'd136314880;
      10120: inst = 32'd268468224;
      10121: inst = 32'd201344968;
      10122: inst = 32'd203484854;
      10123: inst = 32'd471859200;
      10124: inst = 32'd136314880;
      10125: inst = 32'd268468224;
      10126: inst = 32'd201344969;
      10127: inst = 32'd203484854;
      10128: inst = 32'd471859200;
      10129: inst = 32'd136314880;
      10130: inst = 32'd268468224;
      10131: inst = 32'd201344970;
      10132: inst = 32'd203484854;
      10133: inst = 32'd471859200;
      10134: inst = 32'd136314880;
      10135: inst = 32'd268468224;
      10136: inst = 32'd201344971;
      10137: inst = 32'd203484854;
      10138: inst = 32'd471859200;
      10139: inst = 32'd136314880;
      10140: inst = 32'd268468224;
      10141: inst = 32'd201344972;
      10142: inst = 32'd203484854;
      10143: inst = 32'd471859200;
      10144: inst = 32'd136314880;
      10145: inst = 32'd268468224;
      10146: inst = 32'd201344973;
      10147: inst = 32'd203484854;
      10148: inst = 32'd471859200;
      10149: inst = 32'd136314880;
      10150: inst = 32'd268468224;
      10151: inst = 32'd201344974;
      10152: inst = 32'd203484854;
      10153: inst = 32'd471859200;
      10154: inst = 32'd136314880;
      10155: inst = 32'd268468224;
      10156: inst = 32'd201344975;
      10157: inst = 32'd203484854;
      10158: inst = 32'd471859200;
      10159: inst = 32'd136314880;
      10160: inst = 32'd268468224;
      10161: inst = 32'd201344976;
      10162: inst = 32'd203484854;
      10163: inst = 32'd471859200;
      10164: inst = 32'd136314880;
      10165: inst = 32'd268468224;
      10166: inst = 32'd201344977;
      10167: inst = 32'd203484854;
      10168: inst = 32'd471859200;
      10169: inst = 32'd136314880;
      10170: inst = 32'd268468224;
      10171: inst = 32'd201344978;
      10172: inst = 32'd203484854;
      10173: inst = 32'd471859200;
      10174: inst = 32'd136314880;
      10175: inst = 32'd268468224;
      10176: inst = 32'd201344979;
      10177: inst = 32'd203484854;
      10178: inst = 32'd471859200;
      10179: inst = 32'd136314880;
      10180: inst = 32'd268468224;
      10181: inst = 32'd201344980;
      10182: inst = 32'd203484854;
      10183: inst = 32'd471859200;
      10184: inst = 32'd136314880;
      10185: inst = 32'd268468224;
      10186: inst = 32'd201344981;
      10187: inst = 32'd203484854;
      10188: inst = 32'd471859200;
      10189: inst = 32'd136314880;
      10190: inst = 32'd268468224;
      10191: inst = 32'd201344982;
      10192: inst = 32'd203484854;
      10193: inst = 32'd471859200;
      10194: inst = 32'd136314880;
      10195: inst = 32'd268468224;
      10196: inst = 32'd201344983;
      10197: inst = 32'd203484854;
      10198: inst = 32'd471859200;
      10199: inst = 32'd136314880;
      10200: inst = 32'd268468224;
      10201: inst = 32'd201344984;
      10202: inst = 32'd203484854;
      10203: inst = 32'd471859200;
      10204: inst = 32'd136314880;
      10205: inst = 32'd268468224;
      10206: inst = 32'd201344985;
      10207: inst = 32'd203484854;
      10208: inst = 32'd471859200;
      10209: inst = 32'd136314880;
      10210: inst = 32'd268468224;
      10211: inst = 32'd201344986;
      10212: inst = 32'd203484854;
      10213: inst = 32'd471859200;
      10214: inst = 32'd136314880;
      10215: inst = 32'd268468224;
      10216: inst = 32'd201344987;
      10217: inst = 32'd203484854;
      10218: inst = 32'd471859200;
      10219: inst = 32'd136314880;
      10220: inst = 32'd268468224;
      10221: inst = 32'd201344988;
      10222: inst = 32'd203489279;
      10223: inst = 32'd471859200;
      10224: inst = 32'd136314880;
      10225: inst = 32'd268468224;
      10226: inst = 32'd201344989;
      10227: inst = 32'd203489279;
      10228: inst = 32'd471859200;
      10229: inst = 32'd136314880;
      10230: inst = 32'd268468224;
      10231: inst = 32'd201344990;
      10232: inst = 32'd203489279;
      10233: inst = 32'd471859200;
      10234: inst = 32'd136314880;
      10235: inst = 32'd268468224;
      10236: inst = 32'd201344991;
      10237: inst = 32'd203489279;
      10238: inst = 32'd471859200;
      10239: inst = 32'd136314880;
      10240: inst = 32'd268468224;
      10241: inst = 32'd201344992;
      10242: inst = 32'd203489279;
      10243: inst = 32'd471859200;
      10244: inst = 32'd136314880;
      10245: inst = 32'd268468224;
      10246: inst = 32'd201344993;
      10247: inst = 32'd203489279;
      10248: inst = 32'd471859200;
      10249: inst = 32'd136314880;
      10250: inst = 32'd268468224;
      10251: inst = 32'd201344994;
      10252: inst = 32'd203489279;
      10253: inst = 32'd471859200;
      10254: inst = 32'd136314880;
      10255: inst = 32'd268468224;
      10256: inst = 32'd201344995;
      10257: inst = 32'd203489279;
      10258: inst = 32'd471859200;
      10259: inst = 32'd136314880;
      10260: inst = 32'd268468224;
      10261: inst = 32'd201344996;
      10262: inst = 32'd203489279;
      10263: inst = 32'd471859200;
      10264: inst = 32'd136314880;
      10265: inst = 32'd268468224;
      10266: inst = 32'd201344997;
      10267: inst = 32'd203489279;
      10268: inst = 32'd471859200;
      10269: inst = 32'd136314880;
      10270: inst = 32'd268468224;
      10271: inst = 32'd201344998;
      10272: inst = 32'd203489279;
      10273: inst = 32'd471859200;
      10274: inst = 32'd136314880;
      10275: inst = 32'd268468224;
      10276: inst = 32'd201344999;
      10277: inst = 32'd203489279;
      10278: inst = 32'd471859200;
      10279: inst = 32'd136314880;
      10280: inst = 32'd268468224;
      10281: inst = 32'd201345000;
      10282: inst = 32'd203489279;
      10283: inst = 32'd471859200;
      10284: inst = 32'd136314880;
      10285: inst = 32'd268468224;
      10286: inst = 32'd201345001;
      10287: inst = 32'd203489279;
      10288: inst = 32'd471859200;
      10289: inst = 32'd136314880;
      10290: inst = 32'd268468224;
      10291: inst = 32'd201345002;
      10292: inst = 32'd203489279;
      10293: inst = 32'd471859200;
      10294: inst = 32'd136314880;
      10295: inst = 32'd268468224;
      10296: inst = 32'd201345003;
      10297: inst = 32'd203489279;
      10298: inst = 32'd471859200;
      10299: inst = 32'd136314880;
      10300: inst = 32'd268468224;
      10301: inst = 32'd201345004;
      10302: inst = 32'd203489279;
      10303: inst = 32'd471859200;
      10304: inst = 32'd136314880;
      10305: inst = 32'd268468224;
      10306: inst = 32'd201345005;
      10307: inst = 32'd203489279;
      10308: inst = 32'd471859200;
      10309: inst = 32'd136314880;
      10310: inst = 32'd268468224;
      10311: inst = 32'd201345006;
      10312: inst = 32'd203489279;
      10313: inst = 32'd471859200;
      10314: inst = 32'd136314880;
      10315: inst = 32'd268468224;
      10316: inst = 32'd201345007;
      10317: inst = 32'd203489279;
      10318: inst = 32'd471859200;
      10319: inst = 32'd136314880;
      10320: inst = 32'd268468224;
      10321: inst = 32'd201345008;
      10322: inst = 32'd203489279;
      10323: inst = 32'd471859200;
      10324: inst = 32'd136314880;
      10325: inst = 32'd268468224;
      10326: inst = 32'd201345009;
      10327: inst = 32'd203489279;
      10328: inst = 32'd471859200;
      10329: inst = 32'd136314880;
      10330: inst = 32'd268468224;
      10331: inst = 32'd201345010;
      10332: inst = 32'd203489279;
      10333: inst = 32'd471859200;
      10334: inst = 32'd136314880;
      10335: inst = 32'd268468224;
      10336: inst = 32'd201345011;
      10337: inst = 32'd203489279;
      10338: inst = 32'd471859200;
      10339: inst = 32'd136314880;
      10340: inst = 32'd268468224;
      10341: inst = 32'd201345012;
      10342: inst = 32'd203489279;
      10343: inst = 32'd471859200;
      10344: inst = 32'd136314880;
      10345: inst = 32'd268468224;
      10346: inst = 32'd201345013;
      10347: inst = 32'd203489279;
      10348: inst = 32'd471859200;
      10349: inst = 32'd136314880;
      10350: inst = 32'd268468224;
      10351: inst = 32'd201345014;
      10352: inst = 32'd203489279;
      10353: inst = 32'd471859200;
      10354: inst = 32'd136314880;
      10355: inst = 32'd268468224;
      10356: inst = 32'd201345015;
      10357: inst = 32'd203489279;
      10358: inst = 32'd471859200;
      10359: inst = 32'd136314880;
      10360: inst = 32'd268468224;
      10361: inst = 32'd201345016;
      10362: inst = 32'd203489279;
      10363: inst = 32'd471859200;
      10364: inst = 32'd136314880;
      10365: inst = 32'd268468224;
      10366: inst = 32'd201345017;
      10367: inst = 32'd203489279;
      10368: inst = 32'd471859200;
      10369: inst = 32'd136314880;
      10370: inst = 32'd268468224;
      10371: inst = 32'd201345018;
      10372: inst = 32'd203489279;
      10373: inst = 32'd471859200;
      10374: inst = 32'd136314880;
      10375: inst = 32'd268468224;
      10376: inst = 32'd201345019;
      10377: inst = 32'd203489279;
      10378: inst = 32'd471859200;
      10379: inst = 32'd136314880;
      10380: inst = 32'd268468224;
      10381: inst = 32'd201345020;
      10382: inst = 32'd203489279;
      10383: inst = 32'd471859200;
      10384: inst = 32'd136314880;
      10385: inst = 32'd268468224;
      10386: inst = 32'd201345021;
      10387: inst = 32'd203489279;
      10388: inst = 32'd471859200;
      10389: inst = 32'd136314880;
      10390: inst = 32'd268468224;
      10391: inst = 32'd201345022;
      10392: inst = 32'd203489279;
      10393: inst = 32'd471859200;
      10394: inst = 32'd136314880;
      10395: inst = 32'd268468224;
      10396: inst = 32'd201345023;
      10397: inst = 32'd203489279;
      10398: inst = 32'd471859200;
      10399: inst = 32'd136314880;
      10400: inst = 32'd268468224;
      10401: inst = 32'd201345024;
      10402: inst = 32'd203489279;
      10403: inst = 32'd471859200;
      10404: inst = 32'd136314880;
      10405: inst = 32'd268468224;
      10406: inst = 32'd201345025;
      10407: inst = 32'd203489279;
      10408: inst = 32'd471859200;
      10409: inst = 32'd136314880;
      10410: inst = 32'd268468224;
      10411: inst = 32'd201345026;
      10412: inst = 32'd203489279;
      10413: inst = 32'd471859200;
      10414: inst = 32'd136314880;
      10415: inst = 32'd268468224;
      10416: inst = 32'd201345027;
      10417: inst = 32'd203489279;
      10418: inst = 32'd471859200;
      10419: inst = 32'd136314880;
      10420: inst = 32'd268468224;
      10421: inst = 32'd201345028;
      10422: inst = 32'd203484854;
      10423: inst = 32'd471859200;
      10424: inst = 32'd136314880;
      10425: inst = 32'd268468224;
      10426: inst = 32'd201345029;
      10427: inst = 32'd203484854;
      10428: inst = 32'd471859200;
      10429: inst = 32'd136314880;
      10430: inst = 32'd268468224;
      10431: inst = 32'd201345030;
      10432: inst = 32'd203484854;
      10433: inst = 32'd471859200;
      10434: inst = 32'd136314880;
      10435: inst = 32'd268468224;
      10436: inst = 32'd201345031;
      10437: inst = 32'd203484854;
      10438: inst = 32'd471859200;
      10439: inst = 32'd136314880;
      10440: inst = 32'd268468224;
      10441: inst = 32'd201345032;
      10442: inst = 32'd203484854;
      10443: inst = 32'd471859200;
      10444: inst = 32'd136314880;
      10445: inst = 32'd268468224;
      10446: inst = 32'd201345033;
      10447: inst = 32'd203484854;
      10448: inst = 32'd471859200;
      10449: inst = 32'd136314880;
      10450: inst = 32'd268468224;
      10451: inst = 32'd201345034;
      10452: inst = 32'd203484854;
      10453: inst = 32'd471859200;
      10454: inst = 32'd136314880;
      10455: inst = 32'd268468224;
      10456: inst = 32'd201345035;
      10457: inst = 32'd203484854;
      10458: inst = 32'd471859200;
      10459: inst = 32'd136314880;
      10460: inst = 32'd268468224;
      10461: inst = 32'd201345036;
      10462: inst = 32'd203484854;
      10463: inst = 32'd471859200;
      10464: inst = 32'd136314880;
      10465: inst = 32'd268468224;
      10466: inst = 32'd201345037;
      10467: inst = 32'd203484854;
      10468: inst = 32'd471859200;
      10469: inst = 32'd136314880;
      10470: inst = 32'd268468224;
      10471: inst = 32'd201345038;
      10472: inst = 32'd203484854;
      10473: inst = 32'd471859200;
      10474: inst = 32'd136314880;
      10475: inst = 32'd268468224;
      10476: inst = 32'd201345039;
      10477: inst = 32'd203473634;
      10478: inst = 32'd471859200;
      10479: inst = 32'd136314880;
      10480: inst = 32'd268468224;
      10481: inst = 32'd201345040;
      10482: inst = 32'd203480005;
      10483: inst = 32'd471859200;
      10484: inst = 32'd136314880;
      10485: inst = 32'd268468224;
      10486: inst = 32'd201345041;
      10487: inst = 32'd203480005;
      10488: inst = 32'd471859200;
      10489: inst = 32'd136314880;
      10490: inst = 32'd268468224;
      10491: inst = 32'd201345042;
      10492: inst = 32'd203480005;
      10493: inst = 32'd471859200;
      10494: inst = 32'd136314880;
      10495: inst = 32'd268468224;
      10496: inst = 32'd201345043;
      10497: inst = 32'd203480005;
      10498: inst = 32'd471859200;
      10499: inst = 32'd136314880;
      10500: inst = 32'd268468224;
      10501: inst = 32'd201345044;
      10502: inst = 32'd203480005;
      10503: inst = 32'd471859200;
      10504: inst = 32'd136314880;
      10505: inst = 32'd268468224;
      10506: inst = 32'd201345045;
      10507: inst = 32'd203480005;
      10508: inst = 32'd471859200;
      10509: inst = 32'd136314880;
      10510: inst = 32'd268468224;
      10511: inst = 32'd201345046;
      10512: inst = 32'd203480005;
      10513: inst = 32'd471859200;
      10514: inst = 32'd136314880;
      10515: inst = 32'd268468224;
      10516: inst = 32'd201345047;
      10517: inst = 32'd203480005;
      10518: inst = 32'd471859200;
      10519: inst = 32'd136314880;
      10520: inst = 32'd268468224;
      10521: inst = 32'd201345048;
      10522: inst = 32'd203480005;
      10523: inst = 32'd471859200;
      10524: inst = 32'd136314880;
      10525: inst = 32'd268468224;
      10526: inst = 32'd201345049;
      10527: inst = 32'd203480005;
      10528: inst = 32'd471859200;
      10529: inst = 32'd136314880;
      10530: inst = 32'd268468224;
      10531: inst = 32'd201345050;
      10532: inst = 32'd203480005;
      10533: inst = 32'd471859200;
      10534: inst = 32'd136314880;
      10535: inst = 32'd268468224;
      10536: inst = 32'd201345051;
      10537: inst = 32'd203480005;
      10538: inst = 32'd471859200;
      10539: inst = 32'd136314880;
      10540: inst = 32'd268468224;
      10541: inst = 32'd201345052;
      10542: inst = 32'd203480005;
      10543: inst = 32'd471859200;
      10544: inst = 32'd136314880;
      10545: inst = 32'd268468224;
      10546: inst = 32'd201345053;
      10547: inst = 32'd203480005;
      10548: inst = 32'd471859200;
      10549: inst = 32'd136314880;
      10550: inst = 32'd268468224;
      10551: inst = 32'd201345054;
      10552: inst = 32'd203480005;
      10553: inst = 32'd471859200;
      10554: inst = 32'd136314880;
      10555: inst = 32'd268468224;
      10556: inst = 32'd201345055;
      10557: inst = 32'd203473634;
      10558: inst = 32'd471859200;
      10559: inst = 32'd136314880;
      10560: inst = 32'd268468224;
      10561: inst = 32'd201345056;
      10562: inst = 32'd203484854;
      10563: inst = 32'd471859200;
      10564: inst = 32'd136314880;
      10565: inst = 32'd268468224;
      10566: inst = 32'd201345057;
      10567: inst = 32'd203484854;
      10568: inst = 32'd471859200;
      10569: inst = 32'd136314880;
      10570: inst = 32'd268468224;
      10571: inst = 32'd201345058;
      10572: inst = 32'd203484854;
      10573: inst = 32'd471859200;
      10574: inst = 32'd136314880;
      10575: inst = 32'd268468224;
      10576: inst = 32'd201345059;
      10577: inst = 32'd203484854;
      10578: inst = 32'd471859200;
      10579: inst = 32'd136314880;
      10580: inst = 32'd268468224;
      10581: inst = 32'd201345060;
      10582: inst = 32'd203484854;
      10583: inst = 32'd471859200;
      10584: inst = 32'd136314880;
      10585: inst = 32'd268468224;
      10586: inst = 32'd201345061;
      10587: inst = 32'd203484854;
      10588: inst = 32'd471859200;
      10589: inst = 32'd136314880;
      10590: inst = 32'd268468224;
      10591: inst = 32'd201345062;
      10592: inst = 32'd203484854;
      10593: inst = 32'd471859200;
      10594: inst = 32'd136314880;
      10595: inst = 32'd268468224;
      10596: inst = 32'd201345063;
      10597: inst = 32'd203484854;
      10598: inst = 32'd471859200;
      10599: inst = 32'd136314880;
      10600: inst = 32'd268468224;
      10601: inst = 32'd201345064;
      10602: inst = 32'd203484854;
      10603: inst = 32'd471859200;
      10604: inst = 32'd136314880;
      10605: inst = 32'd268468224;
      10606: inst = 32'd201345065;
      10607: inst = 32'd203484854;
      10608: inst = 32'd471859200;
      10609: inst = 32'd136314880;
      10610: inst = 32'd268468224;
      10611: inst = 32'd201345066;
      10612: inst = 32'd203484854;
      10613: inst = 32'd471859200;
      10614: inst = 32'd136314880;
      10615: inst = 32'd268468224;
      10616: inst = 32'd201345067;
      10617: inst = 32'd203484854;
      10618: inst = 32'd471859200;
      10619: inst = 32'd136314880;
      10620: inst = 32'd268468224;
      10621: inst = 32'd201345068;
      10622: inst = 32'd203484854;
      10623: inst = 32'd471859200;
      10624: inst = 32'd136314880;
      10625: inst = 32'd268468224;
      10626: inst = 32'd201345069;
      10627: inst = 32'd203484854;
      10628: inst = 32'd471859200;
      10629: inst = 32'd136314880;
      10630: inst = 32'd268468224;
      10631: inst = 32'd201345070;
      10632: inst = 32'd203484854;
      10633: inst = 32'd471859200;
      10634: inst = 32'd136314880;
      10635: inst = 32'd268468224;
      10636: inst = 32'd201345071;
      10637: inst = 32'd203484854;
      10638: inst = 32'd471859200;
      10639: inst = 32'd136314880;
      10640: inst = 32'd268468224;
      10641: inst = 32'd201345072;
      10642: inst = 32'd203484854;
      10643: inst = 32'd471859200;
      10644: inst = 32'd136314880;
      10645: inst = 32'd268468224;
      10646: inst = 32'd201345073;
      10647: inst = 32'd203484854;
      10648: inst = 32'd471859200;
      10649: inst = 32'd136314880;
      10650: inst = 32'd268468224;
      10651: inst = 32'd201345074;
      10652: inst = 32'd203484854;
      10653: inst = 32'd471859200;
      10654: inst = 32'd136314880;
      10655: inst = 32'd268468224;
      10656: inst = 32'd201345075;
      10657: inst = 32'd203484854;
      10658: inst = 32'd471859200;
      10659: inst = 32'd136314880;
      10660: inst = 32'd268468224;
      10661: inst = 32'd201345076;
      10662: inst = 32'd203484854;
      10663: inst = 32'd471859200;
      10664: inst = 32'd136314880;
      10665: inst = 32'd268468224;
      10666: inst = 32'd201345077;
      10667: inst = 32'd203484854;
      10668: inst = 32'd471859200;
      10669: inst = 32'd136314880;
      10670: inst = 32'd268468224;
      10671: inst = 32'd201345078;
      10672: inst = 32'd203484854;
      10673: inst = 32'd471859200;
      10674: inst = 32'd136314880;
      10675: inst = 32'd268468224;
      10676: inst = 32'd201345079;
      10677: inst = 32'd203484854;
      10678: inst = 32'd471859200;
      10679: inst = 32'd136314880;
      10680: inst = 32'd268468224;
      10681: inst = 32'd201345080;
      10682: inst = 32'd203484854;
      10683: inst = 32'd471859200;
      10684: inst = 32'd136314880;
      10685: inst = 32'd268468224;
      10686: inst = 32'd201345081;
      10687: inst = 32'd203484854;
      10688: inst = 32'd471859200;
      10689: inst = 32'd136314880;
      10690: inst = 32'd268468224;
      10691: inst = 32'd201345082;
      10692: inst = 32'd203484854;
      10693: inst = 32'd471859200;
      10694: inst = 32'd136314880;
      10695: inst = 32'd268468224;
      10696: inst = 32'd201345083;
      10697: inst = 32'd203484854;
      10698: inst = 32'd471859200;
      10699: inst = 32'd136314880;
      10700: inst = 32'd268468224;
      10701: inst = 32'd201345084;
      10702: inst = 32'd203489279;
      10703: inst = 32'd471859200;
      10704: inst = 32'd136314880;
      10705: inst = 32'd268468224;
      10706: inst = 32'd201345085;
      10707: inst = 32'd203489279;
      10708: inst = 32'd471859200;
      10709: inst = 32'd136314880;
      10710: inst = 32'd268468224;
      10711: inst = 32'd201345086;
      10712: inst = 32'd203489279;
      10713: inst = 32'd471859200;
      10714: inst = 32'd136314880;
      10715: inst = 32'd268468224;
      10716: inst = 32'd201345087;
      10717: inst = 32'd203489279;
      10718: inst = 32'd471859200;
      10719: inst = 32'd136314880;
      10720: inst = 32'd268468224;
      10721: inst = 32'd201345088;
      10722: inst = 32'd203489279;
      10723: inst = 32'd471859200;
      10724: inst = 32'd136314880;
      10725: inst = 32'd268468224;
      10726: inst = 32'd201345089;
      10727: inst = 32'd203489279;
      10728: inst = 32'd471859200;
      10729: inst = 32'd136314880;
      10730: inst = 32'd268468224;
      10731: inst = 32'd201345090;
      10732: inst = 32'd203489279;
      10733: inst = 32'd471859200;
      10734: inst = 32'd136314880;
      10735: inst = 32'd268468224;
      10736: inst = 32'd201345091;
      10737: inst = 32'd203489279;
      10738: inst = 32'd471859200;
      10739: inst = 32'd136314880;
      10740: inst = 32'd268468224;
      10741: inst = 32'd201345092;
      10742: inst = 32'd203489279;
      10743: inst = 32'd471859200;
      10744: inst = 32'd136314880;
      10745: inst = 32'd268468224;
      10746: inst = 32'd201345093;
      10747: inst = 32'd203489279;
      10748: inst = 32'd471859200;
      10749: inst = 32'd136314880;
      10750: inst = 32'd268468224;
      10751: inst = 32'd201345094;
      10752: inst = 32'd203489279;
      10753: inst = 32'd471859200;
      10754: inst = 32'd136314880;
      10755: inst = 32'd268468224;
      10756: inst = 32'd201345095;
      10757: inst = 32'd203489279;
      10758: inst = 32'd471859200;
      10759: inst = 32'd136314880;
      10760: inst = 32'd268468224;
      10761: inst = 32'd201345096;
      10762: inst = 32'd203489279;
      10763: inst = 32'd471859200;
      10764: inst = 32'd136314880;
      10765: inst = 32'd268468224;
      10766: inst = 32'd201345097;
      10767: inst = 32'd203489279;
      10768: inst = 32'd471859200;
      10769: inst = 32'd136314880;
      10770: inst = 32'd268468224;
      10771: inst = 32'd201345098;
      10772: inst = 32'd203489279;
      10773: inst = 32'd471859200;
      10774: inst = 32'd136314880;
      10775: inst = 32'd268468224;
      10776: inst = 32'd201345099;
      10777: inst = 32'd203489279;
      10778: inst = 32'd471859200;
      10779: inst = 32'd136314880;
      10780: inst = 32'd268468224;
      10781: inst = 32'd201345100;
      10782: inst = 32'd203489279;
      10783: inst = 32'd471859200;
      10784: inst = 32'd136314880;
      10785: inst = 32'd268468224;
      10786: inst = 32'd201345101;
      10787: inst = 32'd203489279;
      10788: inst = 32'd471859200;
      10789: inst = 32'd136314880;
      10790: inst = 32'd268468224;
      10791: inst = 32'd201345102;
      10792: inst = 32'd203489279;
      10793: inst = 32'd471859200;
      10794: inst = 32'd136314880;
      10795: inst = 32'd268468224;
      10796: inst = 32'd201345103;
      10797: inst = 32'd203489279;
      10798: inst = 32'd471859200;
      10799: inst = 32'd136314880;
      10800: inst = 32'd268468224;
      10801: inst = 32'd201345104;
      10802: inst = 32'd203489279;
      10803: inst = 32'd471859200;
      10804: inst = 32'd136314880;
      10805: inst = 32'd268468224;
      10806: inst = 32'd201345105;
      10807: inst = 32'd203489279;
      10808: inst = 32'd471859200;
      10809: inst = 32'd136314880;
      10810: inst = 32'd268468224;
      10811: inst = 32'd201345106;
      10812: inst = 32'd203489279;
      10813: inst = 32'd471859200;
      10814: inst = 32'd136314880;
      10815: inst = 32'd268468224;
      10816: inst = 32'd201345107;
      10817: inst = 32'd203489279;
      10818: inst = 32'd471859200;
      10819: inst = 32'd136314880;
      10820: inst = 32'd268468224;
      10821: inst = 32'd201345108;
      10822: inst = 32'd203489279;
      10823: inst = 32'd471859200;
      10824: inst = 32'd136314880;
      10825: inst = 32'd268468224;
      10826: inst = 32'd201345109;
      10827: inst = 32'd203489279;
      10828: inst = 32'd471859200;
      10829: inst = 32'd136314880;
      10830: inst = 32'd268468224;
      10831: inst = 32'd201345110;
      10832: inst = 32'd203489279;
      10833: inst = 32'd471859200;
      10834: inst = 32'd136314880;
      10835: inst = 32'd268468224;
      10836: inst = 32'd201345111;
      10837: inst = 32'd203489279;
      10838: inst = 32'd471859200;
      10839: inst = 32'd136314880;
      10840: inst = 32'd268468224;
      10841: inst = 32'd201345112;
      10842: inst = 32'd203489279;
      10843: inst = 32'd471859200;
      10844: inst = 32'd136314880;
      10845: inst = 32'd268468224;
      10846: inst = 32'd201345113;
      10847: inst = 32'd203489279;
      10848: inst = 32'd471859200;
      10849: inst = 32'd136314880;
      10850: inst = 32'd268468224;
      10851: inst = 32'd201345114;
      10852: inst = 32'd203489279;
      10853: inst = 32'd471859200;
      10854: inst = 32'd136314880;
      10855: inst = 32'd268468224;
      10856: inst = 32'd201345115;
      10857: inst = 32'd203489279;
      10858: inst = 32'd471859200;
      10859: inst = 32'd136314880;
      10860: inst = 32'd268468224;
      10861: inst = 32'd201345116;
      10862: inst = 32'd203489279;
      10863: inst = 32'd471859200;
      10864: inst = 32'd136314880;
      10865: inst = 32'd268468224;
      10866: inst = 32'd201345117;
      10867: inst = 32'd203489279;
      10868: inst = 32'd471859200;
      10869: inst = 32'd136314880;
      10870: inst = 32'd268468224;
      10871: inst = 32'd201345118;
      10872: inst = 32'd203489279;
      10873: inst = 32'd471859200;
      10874: inst = 32'd136314880;
      10875: inst = 32'd268468224;
      10876: inst = 32'd201345119;
      10877: inst = 32'd203489279;
      10878: inst = 32'd471859200;
      10879: inst = 32'd136314880;
      10880: inst = 32'd268468224;
      10881: inst = 32'd201345120;
      10882: inst = 32'd203489279;
      10883: inst = 32'd471859200;
      10884: inst = 32'd136314880;
      10885: inst = 32'd268468224;
      10886: inst = 32'd201345121;
      10887: inst = 32'd203489279;
      10888: inst = 32'd471859200;
      10889: inst = 32'd136314880;
      10890: inst = 32'd268468224;
      10891: inst = 32'd201345122;
      10892: inst = 32'd203489279;
      10893: inst = 32'd471859200;
      10894: inst = 32'd136314880;
      10895: inst = 32'd268468224;
      10896: inst = 32'd201345123;
      10897: inst = 32'd203489279;
      10898: inst = 32'd471859200;
      10899: inst = 32'd136314880;
      10900: inst = 32'd268468224;
      10901: inst = 32'd201345124;
      10902: inst = 32'd203484854;
      10903: inst = 32'd471859200;
      10904: inst = 32'd136314880;
      10905: inst = 32'd268468224;
      10906: inst = 32'd201345125;
      10907: inst = 32'd203484854;
      10908: inst = 32'd471859200;
      10909: inst = 32'd136314880;
      10910: inst = 32'd268468224;
      10911: inst = 32'd201345126;
      10912: inst = 32'd203484854;
      10913: inst = 32'd471859200;
      10914: inst = 32'd136314880;
      10915: inst = 32'd268468224;
      10916: inst = 32'd201345127;
      10917: inst = 32'd203484854;
      10918: inst = 32'd471859200;
      10919: inst = 32'd136314880;
      10920: inst = 32'd268468224;
      10921: inst = 32'd201345128;
      10922: inst = 32'd203484854;
      10923: inst = 32'd471859200;
      10924: inst = 32'd136314880;
      10925: inst = 32'd268468224;
      10926: inst = 32'd201345129;
      10927: inst = 32'd203484854;
      10928: inst = 32'd471859200;
      10929: inst = 32'd136314880;
      10930: inst = 32'd268468224;
      10931: inst = 32'd201345130;
      10932: inst = 32'd203484854;
      10933: inst = 32'd471859200;
      10934: inst = 32'd136314880;
      10935: inst = 32'd268468224;
      10936: inst = 32'd201345131;
      10937: inst = 32'd203484854;
      10938: inst = 32'd471859200;
      10939: inst = 32'd136314880;
      10940: inst = 32'd268468224;
      10941: inst = 32'd201345132;
      10942: inst = 32'd203484854;
      10943: inst = 32'd471859200;
      10944: inst = 32'd136314880;
      10945: inst = 32'd268468224;
      10946: inst = 32'd201345133;
      10947: inst = 32'd203484854;
      10948: inst = 32'd471859200;
      10949: inst = 32'd136314880;
      10950: inst = 32'd268468224;
      10951: inst = 32'd201345134;
      10952: inst = 32'd203484854;
      10953: inst = 32'd471859200;
      10954: inst = 32'd136314880;
      10955: inst = 32'd268468224;
      10956: inst = 32'd201345135;
      10957: inst = 32'd203473634;
      10958: inst = 32'd471859200;
      10959: inst = 32'd136314880;
      10960: inst = 32'd268468224;
      10961: inst = 32'd201345136;
      10962: inst = 32'd203480005;
      10963: inst = 32'd471859200;
      10964: inst = 32'd136314880;
      10965: inst = 32'd268468224;
      10966: inst = 32'd201345137;
      10967: inst = 32'd203480005;
      10968: inst = 32'd471859200;
      10969: inst = 32'd136314880;
      10970: inst = 32'd268468224;
      10971: inst = 32'd201345138;
      10972: inst = 32'd203480005;
      10973: inst = 32'd471859200;
      10974: inst = 32'd136314880;
      10975: inst = 32'd268468224;
      10976: inst = 32'd201345139;
      10977: inst = 32'd203480005;
      10978: inst = 32'd471859200;
      10979: inst = 32'd136314880;
      10980: inst = 32'd268468224;
      10981: inst = 32'd201345140;
      10982: inst = 32'd203480005;
      10983: inst = 32'd471859200;
      10984: inst = 32'd136314880;
      10985: inst = 32'd268468224;
      10986: inst = 32'd201345141;
      10987: inst = 32'd203480005;
      10988: inst = 32'd471859200;
      10989: inst = 32'd136314880;
      10990: inst = 32'd268468224;
      10991: inst = 32'd201345142;
      10992: inst = 32'd203480005;
      10993: inst = 32'd471859200;
      10994: inst = 32'd136314880;
      10995: inst = 32'd268468224;
      10996: inst = 32'd201345143;
      10997: inst = 32'd203480005;
      10998: inst = 32'd471859200;
      10999: inst = 32'd136314880;
      11000: inst = 32'd268468224;
      11001: inst = 32'd201345144;
      11002: inst = 32'd203480005;
      11003: inst = 32'd471859200;
      11004: inst = 32'd136314880;
      11005: inst = 32'd268468224;
      11006: inst = 32'd201345145;
      11007: inst = 32'd203480005;
      11008: inst = 32'd471859200;
      11009: inst = 32'd136314880;
      11010: inst = 32'd268468224;
      11011: inst = 32'd201345146;
      11012: inst = 32'd203480005;
      11013: inst = 32'd471859200;
      11014: inst = 32'd136314880;
      11015: inst = 32'd268468224;
      11016: inst = 32'd201345147;
      11017: inst = 32'd203480005;
      11018: inst = 32'd471859200;
      11019: inst = 32'd136314880;
      11020: inst = 32'd268468224;
      11021: inst = 32'd201345148;
      11022: inst = 32'd203480005;
      11023: inst = 32'd471859200;
      11024: inst = 32'd136314880;
      11025: inst = 32'd268468224;
      11026: inst = 32'd201345149;
      11027: inst = 32'd203480005;
      11028: inst = 32'd471859200;
      11029: inst = 32'd136314880;
      11030: inst = 32'd268468224;
      11031: inst = 32'd201345150;
      11032: inst = 32'd203480005;
      11033: inst = 32'd471859200;
      11034: inst = 32'd136314880;
      11035: inst = 32'd268468224;
      11036: inst = 32'd201345151;
      11037: inst = 32'd203473634;
      11038: inst = 32'd471859200;
      11039: inst = 32'd136314880;
      11040: inst = 32'd268468224;
      11041: inst = 32'd201345152;
      11042: inst = 32'd203484854;
      11043: inst = 32'd471859200;
      11044: inst = 32'd136314880;
      11045: inst = 32'd268468224;
      11046: inst = 32'd201345153;
      11047: inst = 32'd203484854;
      11048: inst = 32'd471859200;
      11049: inst = 32'd136314880;
      11050: inst = 32'd268468224;
      11051: inst = 32'd201345154;
      11052: inst = 32'd203484854;
      11053: inst = 32'd471859200;
      11054: inst = 32'd136314880;
      11055: inst = 32'd268468224;
      11056: inst = 32'd201345155;
      11057: inst = 32'd203484854;
      11058: inst = 32'd471859200;
      11059: inst = 32'd136314880;
      11060: inst = 32'd268468224;
      11061: inst = 32'd201345156;
      11062: inst = 32'd203484854;
      11063: inst = 32'd471859200;
      11064: inst = 32'd136314880;
      11065: inst = 32'd268468224;
      11066: inst = 32'd201345157;
      11067: inst = 32'd203484854;
      11068: inst = 32'd471859200;
      11069: inst = 32'd136314880;
      11070: inst = 32'd268468224;
      11071: inst = 32'd201345158;
      11072: inst = 32'd203484854;
      11073: inst = 32'd471859200;
      11074: inst = 32'd136314880;
      11075: inst = 32'd268468224;
      11076: inst = 32'd201345159;
      11077: inst = 32'd203484854;
      11078: inst = 32'd471859200;
      11079: inst = 32'd136314880;
      11080: inst = 32'd268468224;
      11081: inst = 32'd201345160;
      11082: inst = 32'd203484854;
      11083: inst = 32'd471859200;
      11084: inst = 32'd136314880;
      11085: inst = 32'd268468224;
      11086: inst = 32'd201345161;
      11087: inst = 32'd203484854;
      11088: inst = 32'd471859200;
      11089: inst = 32'd136314880;
      11090: inst = 32'd268468224;
      11091: inst = 32'd201345162;
      11092: inst = 32'd203484854;
      11093: inst = 32'd471859200;
      11094: inst = 32'd136314880;
      11095: inst = 32'd268468224;
      11096: inst = 32'd201345163;
      11097: inst = 32'd203484854;
      11098: inst = 32'd471859200;
      11099: inst = 32'd136314880;
      11100: inst = 32'd268468224;
      11101: inst = 32'd201345164;
      11102: inst = 32'd203484854;
      11103: inst = 32'd471859200;
      11104: inst = 32'd136314880;
      11105: inst = 32'd268468224;
      11106: inst = 32'd201345165;
      11107: inst = 32'd203484854;
      11108: inst = 32'd471859200;
      11109: inst = 32'd136314880;
      11110: inst = 32'd268468224;
      11111: inst = 32'd201345166;
      11112: inst = 32'd203484854;
      11113: inst = 32'd471859200;
      11114: inst = 32'd136314880;
      11115: inst = 32'd268468224;
      11116: inst = 32'd201345167;
      11117: inst = 32'd203484854;
      11118: inst = 32'd471859200;
      11119: inst = 32'd136314880;
      11120: inst = 32'd268468224;
      11121: inst = 32'd201345168;
      11122: inst = 32'd203484854;
      11123: inst = 32'd471859200;
      11124: inst = 32'd136314880;
      11125: inst = 32'd268468224;
      11126: inst = 32'd201345169;
      11127: inst = 32'd203484854;
      11128: inst = 32'd471859200;
      11129: inst = 32'd136314880;
      11130: inst = 32'd268468224;
      11131: inst = 32'd201345170;
      11132: inst = 32'd203484854;
      11133: inst = 32'd471859200;
      11134: inst = 32'd136314880;
      11135: inst = 32'd268468224;
      11136: inst = 32'd201345171;
      11137: inst = 32'd203484854;
      11138: inst = 32'd471859200;
      11139: inst = 32'd136314880;
      11140: inst = 32'd268468224;
      11141: inst = 32'd201345172;
      11142: inst = 32'd203484854;
      11143: inst = 32'd471859200;
      11144: inst = 32'd136314880;
      11145: inst = 32'd268468224;
      11146: inst = 32'd201345173;
      11147: inst = 32'd203484854;
      11148: inst = 32'd471859200;
      11149: inst = 32'd136314880;
      11150: inst = 32'd268468224;
      11151: inst = 32'd201345174;
      11152: inst = 32'd203484854;
      11153: inst = 32'd471859200;
      11154: inst = 32'd136314880;
      11155: inst = 32'd268468224;
      11156: inst = 32'd201345175;
      11157: inst = 32'd203484854;
      11158: inst = 32'd471859200;
      11159: inst = 32'd136314880;
      11160: inst = 32'd268468224;
      11161: inst = 32'd201345176;
      11162: inst = 32'd203484854;
      11163: inst = 32'd471859200;
      11164: inst = 32'd136314880;
      11165: inst = 32'd268468224;
      11166: inst = 32'd201345177;
      11167: inst = 32'd203484854;
      11168: inst = 32'd471859200;
      11169: inst = 32'd136314880;
      11170: inst = 32'd268468224;
      11171: inst = 32'd201345178;
      11172: inst = 32'd203484854;
      11173: inst = 32'd471859200;
      11174: inst = 32'd136314880;
      11175: inst = 32'd268468224;
      11176: inst = 32'd201345179;
      11177: inst = 32'd203484854;
      11178: inst = 32'd471859200;
      11179: inst = 32'd136314880;
      11180: inst = 32'd268468224;
      11181: inst = 32'd201345180;
      11182: inst = 32'd203489279;
      11183: inst = 32'd471859200;
      11184: inst = 32'd136314880;
      11185: inst = 32'd268468224;
      11186: inst = 32'd201345181;
      11187: inst = 32'd203489279;
      11188: inst = 32'd471859200;
      11189: inst = 32'd136314880;
      11190: inst = 32'd268468224;
      11191: inst = 32'd201345182;
      11192: inst = 32'd203489279;
      11193: inst = 32'd471859200;
      11194: inst = 32'd136314880;
      11195: inst = 32'd268468224;
      11196: inst = 32'd201345183;
      11197: inst = 32'd203489279;
      11198: inst = 32'd471859200;
      11199: inst = 32'd136314880;
      11200: inst = 32'd268468224;
      11201: inst = 32'd201345184;
      11202: inst = 32'd203489279;
      11203: inst = 32'd471859200;
      11204: inst = 32'd136314880;
      11205: inst = 32'd268468224;
      11206: inst = 32'd201345185;
      11207: inst = 32'd203489279;
      11208: inst = 32'd471859200;
      11209: inst = 32'd136314880;
      11210: inst = 32'd268468224;
      11211: inst = 32'd201345186;
      11212: inst = 32'd203489279;
      11213: inst = 32'd471859200;
      11214: inst = 32'd136314880;
      11215: inst = 32'd268468224;
      11216: inst = 32'd201345187;
      11217: inst = 32'd203489279;
      11218: inst = 32'd471859200;
      11219: inst = 32'd136314880;
      11220: inst = 32'd268468224;
      11221: inst = 32'd201345188;
      11222: inst = 32'd203489279;
      11223: inst = 32'd471859200;
      11224: inst = 32'd136314880;
      11225: inst = 32'd268468224;
      11226: inst = 32'd201345189;
      11227: inst = 32'd203489279;
      11228: inst = 32'd471859200;
      11229: inst = 32'd136314880;
      11230: inst = 32'd268468224;
      11231: inst = 32'd201345190;
      11232: inst = 32'd203489279;
      11233: inst = 32'd471859200;
      11234: inst = 32'd136314880;
      11235: inst = 32'd268468224;
      11236: inst = 32'd201345191;
      11237: inst = 32'd203489279;
      11238: inst = 32'd471859200;
      11239: inst = 32'd136314880;
      11240: inst = 32'd268468224;
      11241: inst = 32'd201345192;
      11242: inst = 32'd203489279;
      11243: inst = 32'd471859200;
      11244: inst = 32'd136314880;
      11245: inst = 32'd268468224;
      11246: inst = 32'd201345193;
      11247: inst = 32'd203489279;
      11248: inst = 32'd471859200;
      11249: inst = 32'd136314880;
      11250: inst = 32'd268468224;
      11251: inst = 32'd201345194;
      11252: inst = 32'd203489279;
      11253: inst = 32'd471859200;
      11254: inst = 32'd136314880;
      11255: inst = 32'd268468224;
      11256: inst = 32'd201345195;
      11257: inst = 32'd203489279;
      11258: inst = 32'd471859200;
      11259: inst = 32'd136314880;
      11260: inst = 32'd268468224;
      11261: inst = 32'd201345196;
      11262: inst = 32'd203489279;
      11263: inst = 32'd471859200;
      11264: inst = 32'd136314880;
      11265: inst = 32'd268468224;
      11266: inst = 32'd201345197;
      11267: inst = 32'd203489279;
      11268: inst = 32'd471859200;
      11269: inst = 32'd136314880;
      11270: inst = 32'd268468224;
      11271: inst = 32'd201345198;
      11272: inst = 32'd203489279;
      11273: inst = 32'd471859200;
      11274: inst = 32'd136314880;
      11275: inst = 32'd268468224;
      11276: inst = 32'd201345199;
      11277: inst = 32'd203489279;
      11278: inst = 32'd471859200;
      11279: inst = 32'd136314880;
      11280: inst = 32'd268468224;
      11281: inst = 32'd201345200;
      11282: inst = 32'd203489279;
      11283: inst = 32'd471859200;
      11284: inst = 32'd136314880;
      11285: inst = 32'd268468224;
      11286: inst = 32'd201345201;
      11287: inst = 32'd203489279;
      11288: inst = 32'd471859200;
      11289: inst = 32'd136314880;
      11290: inst = 32'd268468224;
      11291: inst = 32'd201345202;
      11292: inst = 32'd203489279;
      11293: inst = 32'd471859200;
      11294: inst = 32'd136314880;
      11295: inst = 32'd268468224;
      11296: inst = 32'd201345203;
      11297: inst = 32'd203489279;
      11298: inst = 32'd471859200;
      11299: inst = 32'd136314880;
      11300: inst = 32'd268468224;
      11301: inst = 32'd201345204;
      11302: inst = 32'd203489279;
      11303: inst = 32'd471859200;
      11304: inst = 32'd136314880;
      11305: inst = 32'd268468224;
      11306: inst = 32'd201345205;
      11307: inst = 32'd203489279;
      11308: inst = 32'd471859200;
      11309: inst = 32'd136314880;
      11310: inst = 32'd268468224;
      11311: inst = 32'd201345206;
      11312: inst = 32'd203489279;
      11313: inst = 32'd471859200;
      11314: inst = 32'd136314880;
      11315: inst = 32'd268468224;
      11316: inst = 32'd201345207;
      11317: inst = 32'd203489279;
      11318: inst = 32'd471859200;
      11319: inst = 32'd136314880;
      11320: inst = 32'd268468224;
      11321: inst = 32'd201345208;
      11322: inst = 32'd203489279;
      11323: inst = 32'd471859200;
      11324: inst = 32'd136314880;
      11325: inst = 32'd268468224;
      11326: inst = 32'd201345209;
      11327: inst = 32'd203489279;
      11328: inst = 32'd471859200;
      11329: inst = 32'd136314880;
      11330: inst = 32'd268468224;
      11331: inst = 32'd201345210;
      11332: inst = 32'd203489279;
      11333: inst = 32'd471859200;
      11334: inst = 32'd136314880;
      11335: inst = 32'd268468224;
      11336: inst = 32'd201345211;
      11337: inst = 32'd203489279;
      11338: inst = 32'd471859200;
      11339: inst = 32'd136314880;
      11340: inst = 32'd268468224;
      11341: inst = 32'd201345212;
      11342: inst = 32'd203489279;
      11343: inst = 32'd471859200;
      11344: inst = 32'd136314880;
      11345: inst = 32'd268468224;
      11346: inst = 32'd201345213;
      11347: inst = 32'd203489279;
      11348: inst = 32'd471859200;
      11349: inst = 32'd136314880;
      11350: inst = 32'd268468224;
      11351: inst = 32'd201345214;
      11352: inst = 32'd203489279;
      11353: inst = 32'd471859200;
      11354: inst = 32'd136314880;
      11355: inst = 32'd268468224;
      11356: inst = 32'd201345215;
      11357: inst = 32'd203489279;
      11358: inst = 32'd471859200;
      11359: inst = 32'd136314880;
      11360: inst = 32'd268468224;
      11361: inst = 32'd201345216;
      11362: inst = 32'd203489279;
      11363: inst = 32'd471859200;
      11364: inst = 32'd136314880;
      11365: inst = 32'd268468224;
      11366: inst = 32'd201345217;
      11367: inst = 32'd203489279;
      11368: inst = 32'd471859200;
      11369: inst = 32'd136314880;
      11370: inst = 32'd268468224;
      11371: inst = 32'd201345218;
      11372: inst = 32'd203489279;
      11373: inst = 32'd471859200;
      11374: inst = 32'd136314880;
      11375: inst = 32'd268468224;
      11376: inst = 32'd201345219;
      11377: inst = 32'd203489279;
      11378: inst = 32'd471859200;
      11379: inst = 32'd136314880;
      11380: inst = 32'd268468224;
      11381: inst = 32'd201345220;
      11382: inst = 32'd203484854;
      11383: inst = 32'd471859200;
      11384: inst = 32'd136314880;
      11385: inst = 32'd268468224;
      11386: inst = 32'd201345221;
      11387: inst = 32'd203484854;
      11388: inst = 32'd471859200;
      11389: inst = 32'd136314880;
      11390: inst = 32'd268468224;
      11391: inst = 32'd201345222;
      11392: inst = 32'd203484854;
      11393: inst = 32'd471859200;
      11394: inst = 32'd136314880;
      11395: inst = 32'd268468224;
      11396: inst = 32'd201345223;
      11397: inst = 32'd203484854;
      11398: inst = 32'd471859200;
      11399: inst = 32'd136314880;
      11400: inst = 32'd268468224;
      11401: inst = 32'd201345224;
      11402: inst = 32'd203484854;
      11403: inst = 32'd471859200;
      11404: inst = 32'd136314880;
      11405: inst = 32'd268468224;
      11406: inst = 32'd201345225;
      11407: inst = 32'd203484854;
      11408: inst = 32'd471859200;
      11409: inst = 32'd136314880;
      11410: inst = 32'd268468224;
      11411: inst = 32'd201345226;
      11412: inst = 32'd203484854;
      11413: inst = 32'd471859200;
      11414: inst = 32'd136314880;
      11415: inst = 32'd268468224;
      11416: inst = 32'd201345227;
      11417: inst = 32'd203484854;
      11418: inst = 32'd471859200;
      11419: inst = 32'd136314880;
      11420: inst = 32'd268468224;
      11421: inst = 32'd201345228;
      11422: inst = 32'd203484854;
      11423: inst = 32'd471859200;
      11424: inst = 32'd136314880;
      11425: inst = 32'd268468224;
      11426: inst = 32'd201345229;
      11427: inst = 32'd203484854;
      11428: inst = 32'd471859200;
      11429: inst = 32'd136314880;
      11430: inst = 32'd268468224;
      11431: inst = 32'd201345230;
      11432: inst = 32'd203484854;
      11433: inst = 32'd471859200;
      11434: inst = 32'd136314880;
      11435: inst = 32'd268468224;
      11436: inst = 32'd201345231;
      11437: inst = 32'd203473634;
      11438: inst = 32'd471859200;
      11439: inst = 32'd136314880;
      11440: inst = 32'd268468224;
      11441: inst = 32'd201345232;
      11442: inst = 32'd203480005;
      11443: inst = 32'd471859200;
      11444: inst = 32'd136314880;
      11445: inst = 32'd268468224;
      11446: inst = 32'd201345233;
      11447: inst = 32'd203480005;
      11448: inst = 32'd471859200;
      11449: inst = 32'd136314880;
      11450: inst = 32'd268468224;
      11451: inst = 32'd201345234;
      11452: inst = 32'd203480005;
      11453: inst = 32'd471859200;
      11454: inst = 32'd136314880;
      11455: inst = 32'd268468224;
      11456: inst = 32'd201345235;
      11457: inst = 32'd203480005;
      11458: inst = 32'd471859200;
      11459: inst = 32'd136314880;
      11460: inst = 32'd268468224;
      11461: inst = 32'd201345236;
      11462: inst = 32'd203480005;
      11463: inst = 32'd471859200;
      11464: inst = 32'd136314880;
      11465: inst = 32'd268468224;
      11466: inst = 32'd201345237;
      11467: inst = 32'd203480005;
      11468: inst = 32'd471859200;
      11469: inst = 32'd136314880;
      11470: inst = 32'd268468224;
      11471: inst = 32'd201345238;
      11472: inst = 32'd203480005;
      11473: inst = 32'd471859200;
      11474: inst = 32'd136314880;
      11475: inst = 32'd268468224;
      11476: inst = 32'd201345239;
      11477: inst = 32'd203480005;
      11478: inst = 32'd471859200;
      11479: inst = 32'd136314880;
      11480: inst = 32'd268468224;
      11481: inst = 32'd201345240;
      11482: inst = 32'd203480005;
      11483: inst = 32'd471859200;
      11484: inst = 32'd136314880;
      11485: inst = 32'd268468224;
      11486: inst = 32'd201345241;
      11487: inst = 32'd203480005;
      11488: inst = 32'd471859200;
      11489: inst = 32'd136314880;
      11490: inst = 32'd268468224;
      11491: inst = 32'd201345242;
      11492: inst = 32'd203480005;
      11493: inst = 32'd471859200;
      11494: inst = 32'd136314880;
      11495: inst = 32'd268468224;
      11496: inst = 32'd201345243;
      11497: inst = 32'd203480005;
      11498: inst = 32'd471859200;
      11499: inst = 32'd136314880;
      11500: inst = 32'd268468224;
      11501: inst = 32'd201345244;
      11502: inst = 32'd203480005;
      11503: inst = 32'd471859200;
      11504: inst = 32'd136314880;
      11505: inst = 32'd268468224;
      11506: inst = 32'd201345245;
      11507: inst = 32'd203480005;
      11508: inst = 32'd471859200;
      11509: inst = 32'd136314880;
      11510: inst = 32'd268468224;
      11511: inst = 32'd201345246;
      11512: inst = 32'd203480005;
      11513: inst = 32'd471859200;
      11514: inst = 32'd136314880;
      11515: inst = 32'd268468224;
      11516: inst = 32'd201345247;
      11517: inst = 32'd203473634;
      11518: inst = 32'd471859200;
      11519: inst = 32'd136314880;
      11520: inst = 32'd268468224;
      11521: inst = 32'd201345248;
      11522: inst = 32'd203484854;
      11523: inst = 32'd471859200;
      11524: inst = 32'd136314880;
      11525: inst = 32'd268468224;
      11526: inst = 32'd201345249;
      11527: inst = 32'd203484854;
      11528: inst = 32'd471859200;
      11529: inst = 32'd136314880;
      11530: inst = 32'd268468224;
      11531: inst = 32'd201345250;
      11532: inst = 32'd203484854;
      11533: inst = 32'd471859200;
      11534: inst = 32'd136314880;
      11535: inst = 32'd268468224;
      11536: inst = 32'd201345251;
      11537: inst = 32'd203484854;
      11538: inst = 32'd471859200;
      11539: inst = 32'd136314880;
      11540: inst = 32'd268468224;
      11541: inst = 32'd201345252;
      11542: inst = 32'd203484854;
      11543: inst = 32'd471859200;
      11544: inst = 32'd136314880;
      11545: inst = 32'd268468224;
      11546: inst = 32'd201345253;
      11547: inst = 32'd203484854;
      11548: inst = 32'd471859200;
      11549: inst = 32'd136314880;
      11550: inst = 32'd268468224;
      11551: inst = 32'd201345254;
      11552: inst = 32'd203484854;
      11553: inst = 32'd471859200;
      11554: inst = 32'd136314880;
      11555: inst = 32'd268468224;
      11556: inst = 32'd201345255;
      11557: inst = 32'd203484854;
      11558: inst = 32'd471859200;
      11559: inst = 32'd136314880;
      11560: inst = 32'd268468224;
      11561: inst = 32'd201345256;
      11562: inst = 32'd203484854;
      11563: inst = 32'd471859200;
      11564: inst = 32'd136314880;
      11565: inst = 32'd268468224;
      11566: inst = 32'd201345257;
      11567: inst = 32'd203484854;
      11568: inst = 32'd471859200;
      11569: inst = 32'd136314880;
      11570: inst = 32'd268468224;
      11571: inst = 32'd201345258;
      11572: inst = 32'd203484854;
      11573: inst = 32'd471859200;
      11574: inst = 32'd136314880;
      11575: inst = 32'd268468224;
      11576: inst = 32'd201345259;
      11577: inst = 32'd203484854;
      11578: inst = 32'd471859200;
      11579: inst = 32'd136314880;
      11580: inst = 32'd268468224;
      11581: inst = 32'd201345260;
      11582: inst = 32'd203484854;
      11583: inst = 32'd471859200;
      11584: inst = 32'd136314880;
      11585: inst = 32'd268468224;
      11586: inst = 32'd201345261;
      11587: inst = 32'd203484854;
      11588: inst = 32'd471859200;
      11589: inst = 32'd136314880;
      11590: inst = 32'd268468224;
      11591: inst = 32'd201345262;
      11592: inst = 32'd203484854;
      11593: inst = 32'd471859200;
      11594: inst = 32'd136314880;
      11595: inst = 32'd268468224;
      11596: inst = 32'd201345263;
      11597: inst = 32'd203484854;
      11598: inst = 32'd471859200;
      11599: inst = 32'd136314880;
      11600: inst = 32'd268468224;
      11601: inst = 32'd201345264;
      11602: inst = 32'd203484854;
      11603: inst = 32'd471859200;
      11604: inst = 32'd136314880;
      11605: inst = 32'd268468224;
      11606: inst = 32'd201345265;
      11607: inst = 32'd203484854;
      11608: inst = 32'd471859200;
      11609: inst = 32'd136314880;
      11610: inst = 32'd268468224;
      11611: inst = 32'd201345266;
      11612: inst = 32'd203484854;
      11613: inst = 32'd471859200;
      11614: inst = 32'd136314880;
      11615: inst = 32'd268468224;
      11616: inst = 32'd201345267;
      11617: inst = 32'd203484854;
      11618: inst = 32'd471859200;
      11619: inst = 32'd136314880;
      11620: inst = 32'd268468224;
      11621: inst = 32'd201345268;
      11622: inst = 32'd203484854;
      11623: inst = 32'd471859200;
      11624: inst = 32'd136314880;
      11625: inst = 32'd268468224;
      11626: inst = 32'd201345269;
      11627: inst = 32'd203484854;
      11628: inst = 32'd471859200;
      11629: inst = 32'd136314880;
      11630: inst = 32'd268468224;
      11631: inst = 32'd201345270;
      11632: inst = 32'd203484854;
      11633: inst = 32'd471859200;
      11634: inst = 32'd136314880;
      11635: inst = 32'd268468224;
      11636: inst = 32'd201345271;
      11637: inst = 32'd203484854;
      11638: inst = 32'd471859200;
      11639: inst = 32'd136314880;
      11640: inst = 32'd268468224;
      11641: inst = 32'd201345272;
      11642: inst = 32'd203484854;
      11643: inst = 32'd471859200;
      11644: inst = 32'd136314880;
      11645: inst = 32'd268468224;
      11646: inst = 32'd201345273;
      11647: inst = 32'd203484854;
      11648: inst = 32'd471859200;
      11649: inst = 32'd136314880;
      11650: inst = 32'd268468224;
      11651: inst = 32'd201345274;
      11652: inst = 32'd203484854;
      11653: inst = 32'd471859200;
      11654: inst = 32'd136314880;
      11655: inst = 32'd268468224;
      11656: inst = 32'd201345275;
      11657: inst = 32'd203484854;
      11658: inst = 32'd471859200;
      11659: inst = 32'd136314880;
      11660: inst = 32'd268468224;
      11661: inst = 32'd201345276;
      11662: inst = 32'd203489279;
      11663: inst = 32'd471859200;
      11664: inst = 32'd136314880;
      11665: inst = 32'd268468224;
      11666: inst = 32'd201345277;
      11667: inst = 32'd203489279;
      11668: inst = 32'd471859200;
      11669: inst = 32'd136314880;
      11670: inst = 32'd268468224;
      11671: inst = 32'd201345278;
      11672: inst = 32'd203489279;
      11673: inst = 32'd471859200;
      11674: inst = 32'd136314880;
      11675: inst = 32'd268468224;
      11676: inst = 32'd201345279;
      11677: inst = 32'd203489279;
      11678: inst = 32'd471859200;
      11679: inst = 32'd136314880;
      11680: inst = 32'd268468224;
      11681: inst = 32'd201345280;
      11682: inst = 32'd203489279;
      11683: inst = 32'd471859200;
      11684: inst = 32'd136314880;
      11685: inst = 32'd268468224;
      11686: inst = 32'd201345281;
      11687: inst = 32'd203489279;
      11688: inst = 32'd471859200;
      11689: inst = 32'd136314880;
      11690: inst = 32'd268468224;
      11691: inst = 32'd201345282;
      11692: inst = 32'd203489279;
      11693: inst = 32'd471859200;
      11694: inst = 32'd136314880;
      11695: inst = 32'd268468224;
      11696: inst = 32'd201345283;
      11697: inst = 32'd203489279;
      11698: inst = 32'd471859200;
      11699: inst = 32'd136314880;
      11700: inst = 32'd268468224;
      11701: inst = 32'd201345284;
      11702: inst = 32'd203489279;
      11703: inst = 32'd471859200;
      11704: inst = 32'd136314880;
      11705: inst = 32'd268468224;
      11706: inst = 32'd201345285;
      11707: inst = 32'd203489279;
      11708: inst = 32'd471859200;
      11709: inst = 32'd136314880;
      11710: inst = 32'd268468224;
      11711: inst = 32'd201345286;
      11712: inst = 32'd203489279;
      11713: inst = 32'd471859200;
      11714: inst = 32'd136314880;
      11715: inst = 32'd268468224;
      11716: inst = 32'd201345287;
      11717: inst = 32'd203489279;
      11718: inst = 32'd471859200;
      11719: inst = 32'd136314880;
      11720: inst = 32'd268468224;
      11721: inst = 32'd201345288;
      11722: inst = 32'd203489279;
      11723: inst = 32'd471859200;
      11724: inst = 32'd136314880;
      11725: inst = 32'd268468224;
      11726: inst = 32'd201345289;
      11727: inst = 32'd203489279;
      11728: inst = 32'd471859200;
      11729: inst = 32'd136314880;
      11730: inst = 32'd268468224;
      11731: inst = 32'd201345290;
      11732: inst = 32'd203489279;
      11733: inst = 32'd471859200;
      11734: inst = 32'd136314880;
      11735: inst = 32'd268468224;
      11736: inst = 32'd201345291;
      11737: inst = 32'd203489279;
      11738: inst = 32'd471859200;
      11739: inst = 32'd136314880;
      11740: inst = 32'd268468224;
      11741: inst = 32'd201345292;
      11742: inst = 32'd203489279;
      11743: inst = 32'd471859200;
      11744: inst = 32'd136314880;
      11745: inst = 32'd268468224;
      11746: inst = 32'd201345293;
      11747: inst = 32'd203489279;
      11748: inst = 32'd471859200;
      11749: inst = 32'd136314880;
      11750: inst = 32'd268468224;
      11751: inst = 32'd201345294;
      11752: inst = 32'd203489279;
      11753: inst = 32'd471859200;
      11754: inst = 32'd136314880;
      11755: inst = 32'd268468224;
      11756: inst = 32'd201345295;
      11757: inst = 32'd203489279;
      11758: inst = 32'd471859200;
      11759: inst = 32'd136314880;
      11760: inst = 32'd268468224;
      11761: inst = 32'd201345296;
      11762: inst = 32'd203489279;
      11763: inst = 32'd471859200;
      11764: inst = 32'd136314880;
      11765: inst = 32'd268468224;
      11766: inst = 32'd201345297;
      11767: inst = 32'd203489279;
      11768: inst = 32'd471859200;
      11769: inst = 32'd136314880;
      11770: inst = 32'd268468224;
      11771: inst = 32'd201345298;
      11772: inst = 32'd203489279;
      11773: inst = 32'd471859200;
      11774: inst = 32'd136314880;
      11775: inst = 32'd268468224;
      11776: inst = 32'd201345299;
      11777: inst = 32'd203489279;
      11778: inst = 32'd471859200;
      11779: inst = 32'd136314880;
      11780: inst = 32'd268468224;
      11781: inst = 32'd201345300;
      11782: inst = 32'd203489279;
      11783: inst = 32'd471859200;
      11784: inst = 32'd136314880;
      11785: inst = 32'd268468224;
      11786: inst = 32'd201345301;
      11787: inst = 32'd203489279;
      11788: inst = 32'd471859200;
      11789: inst = 32'd136314880;
      11790: inst = 32'd268468224;
      11791: inst = 32'd201345302;
      11792: inst = 32'd203489279;
      11793: inst = 32'd471859200;
      11794: inst = 32'd136314880;
      11795: inst = 32'd268468224;
      11796: inst = 32'd201345303;
      11797: inst = 32'd203489279;
      11798: inst = 32'd471859200;
      11799: inst = 32'd136314880;
      11800: inst = 32'd268468224;
      11801: inst = 32'd201345304;
      11802: inst = 32'd203489279;
      11803: inst = 32'd471859200;
      11804: inst = 32'd136314880;
      11805: inst = 32'd268468224;
      11806: inst = 32'd201345305;
      11807: inst = 32'd203489279;
      11808: inst = 32'd471859200;
      11809: inst = 32'd136314880;
      11810: inst = 32'd268468224;
      11811: inst = 32'd201345306;
      11812: inst = 32'd203489279;
      11813: inst = 32'd471859200;
      11814: inst = 32'd136314880;
      11815: inst = 32'd268468224;
      11816: inst = 32'd201345307;
      11817: inst = 32'd203489279;
      11818: inst = 32'd471859200;
      11819: inst = 32'd136314880;
      11820: inst = 32'd268468224;
      11821: inst = 32'd201345308;
      11822: inst = 32'd203489279;
      11823: inst = 32'd471859200;
      11824: inst = 32'd136314880;
      11825: inst = 32'd268468224;
      11826: inst = 32'd201345309;
      11827: inst = 32'd203489279;
      11828: inst = 32'd471859200;
      11829: inst = 32'd136314880;
      11830: inst = 32'd268468224;
      11831: inst = 32'd201345310;
      11832: inst = 32'd203489279;
      11833: inst = 32'd471859200;
      11834: inst = 32'd136314880;
      11835: inst = 32'd268468224;
      11836: inst = 32'd201345311;
      11837: inst = 32'd203489279;
      11838: inst = 32'd471859200;
      11839: inst = 32'd136314880;
      11840: inst = 32'd268468224;
      11841: inst = 32'd201345312;
      11842: inst = 32'd203489279;
      11843: inst = 32'd471859200;
      11844: inst = 32'd136314880;
      11845: inst = 32'd268468224;
      11846: inst = 32'd201345313;
      11847: inst = 32'd203489279;
      11848: inst = 32'd471859200;
      11849: inst = 32'd136314880;
      11850: inst = 32'd268468224;
      11851: inst = 32'd201345314;
      11852: inst = 32'd203489279;
      11853: inst = 32'd471859200;
      11854: inst = 32'd136314880;
      11855: inst = 32'd268468224;
      11856: inst = 32'd201345315;
      11857: inst = 32'd203489279;
      11858: inst = 32'd471859200;
      11859: inst = 32'd136314880;
      11860: inst = 32'd268468224;
      11861: inst = 32'd201345316;
      11862: inst = 32'd203484854;
      11863: inst = 32'd471859200;
      11864: inst = 32'd136314880;
      11865: inst = 32'd268468224;
      11866: inst = 32'd201345317;
      11867: inst = 32'd203484854;
      11868: inst = 32'd471859200;
      11869: inst = 32'd136314880;
      11870: inst = 32'd268468224;
      11871: inst = 32'd201345318;
      11872: inst = 32'd203484854;
      11873: inst = 32'd471859200;
      11874: inst = 32'd136314880;
      11875: inst = 32'd268468224;
      11876: inst = 32'd201345319;
      11877: inst = 32'd203484854;
      11878: inst = 32'd471859200;
      11879: inst = 32'd136314880;
      11880: inst = 32'd268468224;
      11881: inst = 32'd201345320;
      11882: inst = 32'd203484854;
      11883: inst = 32'd471859200;
      11884: inst = 32'd136314880;
      11885: inst = 32'd268468224;
      11886: inst = 32'd201345321;
      11887: inst = 32'd203484854;
      11888: inst = 32'd471859200;
      11889: inst = 32'd136314880;
      11890: inst = 32'd268468224;
      11891: inst = 32'd201345322;
      11892: inst = 32'd203484854;
      11893: inst = 32'd471859200;
      11894: inst = 32'd136314880;
      11895: inst = 32'd268468224;
      11896: inst = 32'd201345323;
      11897: inst = 32'd203484854;
      11898: inst = 32'd471859200;
      11899: inst = 32'd136314880;
      11900: inst = 32'd268468224;
      11901: inst = 32'd201345324;
      11902: inst = 32'd203484854;
      11903: inst = 32'd471859200;
      11904: inst = 32'd136314880;
      11905: inst = 32'd268468224;
      11906: inst = 32'd201345325;
      11907: inst = 32'd203484854;
      11908: inst = 32'd471859200;
      11909: inst = 32'd136314880;
      11910: inst = 32'd268468224;
      11911: inst = 32'd201345326;
      11912: inst = 32'd203484854;
      11913: inst = 32'd471859200;
      11914: inst = 32'd136314880;
      11915: inst = 32'd268468224;
      11916: inst = 32'd201345327;
      11917: inst = 32'd203473634;
      11918: inst = 32'd471859200;
      11919: inst = 32'd136314880;
      11920: inst = 32'd268468224;
      11921: inst = 32'd201345328;
      11922: inst = 32'd203480005;
      11923: inst = 32'd471859200;
      11924: inst = 32'd136314880;
      11925: inst = 32'd268468224;
      11926: inst = 32'd201345329;
      11927: inst = 32'd203480005;
      11928: inst = 32'd471859200;
      11929: inst = 32'd136314880;
      11930: inst = 32'd268468224;
      11931: inst = 32'd201345330;
      11932: inst = 32'd203485052;
      11933: inst = 32'd471859200;
      11934: inst = 32'd136314880;
      11935: inst = 32'd268468224;
      11936: inst = 32'd201345331;
      11937: inst = 32'd203485052;
      11938: inst = 32'd471859200;
      11939: inst = 32'd136314880;
      11940: inst = 32'd268468224;
      11941: inst = 32'd201345332;
      11942: inst = 32'd203485052;
      11943: inst = 32'd471859200;
      11944: inst = 32'd136314880;
      11945: inst = 32'd268468224;
      11946: inst = 32'd201345333;
      11947: inst = 32'd203485052;
      11948: inst = 32'd471859200;
      11949: inst = 32'd136314880;
      11950: inst = 32'd268468224;
      11951: inst = 32'd201345334;
      11952: inst = 32'd203480005;
      11953: inst = 32'd471859200;
      11954: inst = 32'd136314880;
      11955: inst = 32'd268468224;
      11956: inst = 32'd201345335;
      11957: inst = 32'd203480005;
      11958: inst = 32'd471859200;
      11959: inst = 32'd136314880;
      11960: inst = 32'd268468224;
      11961: inst = 32'd201345336;
      11962: inst = 32'd203480005;
      11963: inst = 32'd471859200;
      11964: inst = 32'd136314880;
      11965: inst = 32'd268468224;
      11966: inst = 32'd201345337;
      11967: inst = 32'd203480005;
      11968: inst = 32'd471859200;
      11969: inst = 32'd136314880;
      11970: inst = 32'd268468224;
      11971: inst = 32'd201345338;
      11972: inst = 32'd203480005;
      11973: inst = 32'd471859200;
      11974: inst = 32'd136314880;
      11975: inst = 32'd268468224;
      11976: inst = 32'd201345339;
      11977: inst = 32'd203480005;
      11978: inst = 32'd471859200;
      11979: inst = 32'd136314880;
      11980: inst = 32'd268468224;
      11981: inst = 32'd201345340;
      11982: inst = 32'd203480005;
      11983: inst = 32'd471859200;
      11984: inst = 32'd136314880;
      11985: inst = 32'd268468224;
      11986: inst = 32'd201345341;
      11987: inst = 32'd203480005;
      11988: inst = 32'd471859200;
      11989: inst = 32'd136314880;
      11990: inst = 32'd268468224;
      11991: inst = 32'd201345342;
      11992: inst = 32'd203480005;
      11993: inst = 32'd471859200;
      11994: inst = 32'd136314880;
      11995: inst = 32'd268468224;
      11996: inst = 32'd201345343;
      11997: inst = 32'd203473634;
      11998: inst = 32'd471859200;
      11999: inst = 32'd136314880;
      12000: inst = 32'd268468224;
      12001: inst = 32'd201345344;
      12002: inst = 32'd203484854;
      12003: inst = 32'd471859200;
      12004: inst = 32'd136314880;
      12005: inst = 32'd268468224;
      12006: inst = 32'd201345345;
      12007: inst = 32'd203484854;
      12008: inst = 32'd471859200;
      12009: inst = 32'd136314880;
      12010: inst = 32'd268468224;
      12011: inst = 32'd201345346;
      12012: inst = 32'd203484854;
      12013: inst = 32'd471859200;
      12014: inst = 32'd136314880;
      12015: inst = 32'd268468224;
      12016: inst = 32'd201345347;
      12017: inst = 32'd203484854;
      12018: inst = 32'd471859200;
      12019: inst = 32'd136314880;
      12020: inst = 32'd268468224;
      12021: inst = 32'd201345348;
      12022: inst = 32'd203484854;
      12023: inst = 32'd471859200;
      12024: inst = 32'd136314880;
      12025: inst = 32'd268468224;
      12026: inst = 32'd201345349;
      12027: inst = 32'd203484854;
      12028: inst = 32'd471859200;
      12029: inst = 32'd136314880;
      12030: inst = 32'd268468224;
      12031: inst = 32'd201345350;
      12032: inst = 32'd203484854;
      12033: inst = 32'd471859200;
      12034: inst = 32'd136314880;
      12035: inst = 32'd268468224;
      12036: inst = 32'd201345351;
      12037: inst = 32'd203484854;
      12038: inst = 32'd471859200;
      12039: inst = 32'd136314880;
      12040: inst = 32'd268468224;
      12041: inst = 32'd201345352;
      12042: inst = 32'd203484854;
      12043: inst = 32'd471859200;
      12044: inst = 32'd136314880;
      12045: inst = 32'd268468224;
      12046: inst = 32'd201345353;
      12047: inst = 32'd203484854;
      12048: inst = 32'd471859200;
      12049: inst = 32'd136314880;
      12050: inst = 32'd268468224;
      12051: inst = 32'd201345354;
      12052: inst = 32'd203484854;
      12053: inst = 32'd471859200;
      12054: inst = 32'd136314880;
      12055: inst = 32'd268468224;
      12056: inst = 32'd201345355;
      12057: inst = 32'd203484854;
      12058: inst = 32'd471859200;
      12059: inst = 32'd136314880;
      12060: inst = 32'd268468224;
      12061: inst = 32'd201345356;
      12062: inst = 32'd203484854;
      12063: inst = 32'd471859200;
      12064: inst = 32'd136314880;
      12065: inst = 32'd268468224;
      12066: inst = 32'd201345357;
      12067: inst = 32'd203484854;
      12068: inst = 32'd471859200;
      12069: inst = 32'd136314880;
      12070: inst = 32'd268468224;
      12071: inst = 32'd201345358;
      12072: inst = 32'd203484854;
      12073: inst = 32'd471859200;
      12074: inst = 32'd136314880;
      12075: inst = 32'd268468224;
      12076: inst = 32'd201345359;
      12077: inst = 32'd203484854;
      12078: inst = 32'd471859200;
      12079: inst = 32'd136314880;
      12080: inst = 32'd268468224;
      12081: inst = 32'd201345360;
      12082: inst = 32'd203484854;
      12083: inst = 32'd471859200;
      12084: inst = 32'd136314880;
      12085: inst = 32'd268468224;
      12086: inst = 32'd201345361;
      12087: inst = 32'd203484854;
      12088: inst = 32'd471859200;
      12089: inst = 32'd136314880;
      12090: inst = 32'd268468224;
      12091: inst = 32'd201345362;
      12092: inst = 32'd203484854;
      12093: inst = 32'd471859200;
      12094: inst = 32'd136314880;
      12095: inst = 32'd268468224;
      12096: inst = 32'd201345363;
      12097: inst = 32'd203484854;
      12098: inst = 32'd471859200;
      12099: inst = 32'd136314880;
      12100: inst = 32'd268468224;
      12101: inst = 32'd201345364;
      12102: inst = 32'd203484854;
      12103: inst = 32'd471859200;
      12104: inst = 32'd136314880;
      12105: inst = 32'd268468224;
      12106: inst = 32'd201345365;
      12107: inst = 32'd203484854;
      12108: inst = 32'd471859200;
      12109: inst = 32'd136314880;
      12110: inst = 32'd268468224;
      12111: inst = 32'd201345366;
      12112: inst = 32'd203484854;
      12113: inst = 32'd471859200;
      12114: inst = 32'd136314880;
      12115: inst = 32'd268468224;
      12116: inst = 32'd201345367;
      12117: inst = 32'd203484854;
      12118: inst = 32'd471859200;
      12119: inst = 32'd136314880;
      12120: inst = 32'd268468224;
      12121: inst = 32'd201345368;
      12122: inst = 32'd203484854;
      12123: inst = 32'd471859200;
      12124: inst = 32'd136314880;
      12125: inst = 32'd268468224;
      12126: inst = 32'd201345369;
      12127: inst = 32'd203484854;
      12128: inst = 32'd471859200;
      12129: inst = 32'd136314880;
      12130: inst = 32'd268468224;
      12131: inst = 32'd201345370;
      12132: inst = 32'd203484854;
      12133: inst = 32'd471859200;
      12134: inst = 32'd136314880;
      12135: inst = 32'd268468224;
      12136: inst = 32'd201345371;
      12137: inst = 32'd203484854;
      12138: inst = 32'd471859200;
      12139: inst = 32'd136314880;
      12140: inst = 32'd268468224;
      12141: inst = 32'd201345372;
      12142: inst = 32'd203489279;
      12143: inst = 32'd471859200;
      12144: inst = 32'd136314880;
      12145: inst = 32'd268468224;
      12146: inst = 32'd201345373;
      12147: inst = 32'd203489279;
      12148: inst = 32'd471859200;
      12149: inst = 32'd136314880;
      12150: inst = 32'd268468224;
      12151: inst = 32'd201345374;
      12152: inst = 32'd203489279;
      12153: inst = 32'd471859200;
      12154: inst = 32'd136314880;
      12155: inst = 32'd268468224;
      12156: inst = 32'd201345375;
      12157: inst = 32'd203489279;
      12158: inst = 32'd471859200;
      12159: inst = 32'd136314880;
      12160: inst = 32'd268468224;
      12161: inst = 32'd201345376;
      12162: inst = 32'd203489279;
      12163: inst = 32'd471859200;
      12164: inst = 32'd136314880;
      12165: inst = 32'd268468224;
      12166: inst = 32'd201345377;
      12167: inst = 32'd203489279;
      12168: inst = 32'd471859200;
      12169: inst = 32'd136314880;
      12170: inst = 32'd268468224;
      12171: inst = 32'd201345378;
      12172: inst = 32'd203489279;
      12173: inst = 32'd471859200;
      12174: inst = 32'd136314880;
      12175: inst = 32'd268468224;
      12176: inst = 32'd201345379;
      12177: inst = 32'd203489279;
      12178: inst = 32'd471859200;
      12179: inst = 32'd136314880;
      12180: inst = 32'd268468224;
      12181: inst = 32'd201345380;
      12182: inst = 32'd203489279;
      12183: inst = 32'd471859200;
      12184: inst = 32'd136314880;
      12185: inst = 32'd268468224;
      12186: inst = 32'd201345381;
      12187: inst = 32'd203489279;
      12188: inst = 32'd471859200;
      12189: inst = 32'd136314880;
      12190: inst = 32'd268468224;
      12191: inst = 32'd201345382;
      12192: inst = 32'd203489279;
      12193: inst = 32'd471859200;
      12194: inst = 32'd136314880;
      12195: inst = 32'd268468224;
      12196: inst = 32'd201345383;
      12197: inst = 32'd203489279;
      12198: inst = 32'd471859200;
      12199: inst = 32'd136314880;
      12200: inst = 32'd268468224;
      12201: inst = 32'd201345384;
      12202: inst = 32'd203489279;
      12203: inst = 32'd471859200;
      12204: inst = 32'd136314880;
      12205: inst = 32'd268468224;
      12206: inst = 32'd201345385;
      12207: inst = 32'd203489279;
      12208: inst = 32'd471859200;
      12209: inst = 32'd136314880;
      12210: inst = 32'd268468224;
      12211: inst = 32'd201345386;
      12212: inst = 32'd203489279;
      12213: inst = 32'd471859200;
      12214: inst = 32'd136314880;
      12215: inst = 32'd268468224;
      12216: inst = 32'd201345387;
      12217: inst = 32'd203489279;
      12218: inst = 32'd471859200;
      12219: inst = 32'd136314880;
      12220: inst = 32'd268468224;
      12221: inst = 32'd201345388;
      12222: inst = 32'd203489279;
      12223: inst = 32'd471859200;
      12224: inst = 32'd136314880;
      12225: inst = 32'd268468224;
      12226: inst = 32'd201345389;
      12227: inst = 32'd203489279;
      12228: inst = 32'd471859200;
      12229: inst = 32'd136314880;
      12230: inst = 32'd268468224;
      12231: inst = 32'd201345390;
      12232: inst = 32'd203489279;
      12233: inst = 32'd471859200;
      12234: inst = 32'd136314880;
      12235: inst = 32'd268468224;
      12236: inst = 32'd201345391;
      12237: inst = 32'd203489279;
      12238: inst = 32'd471859200;
      12239: inst = 32'd136314880;
      12240: inst = 32'd268468224;
      12241: inst = 32'd201345392;
      12242: inst = 32'd203489279;
      12243: inst = 32'd471859200;
      12244: inst = 32'd136314880;
      12245: inst = 32'd268468224;
      12246: inst = 32'd201345393;
      12247: inst = 32'd203489279;
      12248: inst = 32'd471859200;
      12249: inst = 32'd136314880;
      12250: inst = 32'd268468224;
      12251: inst = 32'd201345394;
      12252: inst = 32'd203489279;
      12253: inst = 32'd471859200;
      12254: inst = 32'd136314880;
      12255: inst = 32'd268468224;
      12256: inst = 32'd201345395;
      12257: inst = 32'd203489279;
      12258: inst = 32'd471859200;
      12259: inst = 32'd136314880;
      12260: inst = 32'd268468224;
      12261: inst = 32'd201345396;
      12262: inst = 32'd203489279;
      12263: inst = 32'd471859200;
      12264: inst = 32'd136314880;
      12265: inst = 32'd268468224;
      12266: inst = 32'd201345397;
      12267: inst = 32'd203489279;
      12268: inst = 32'd471859200;
      12269: inst = 32'd136314880;
      12270: inst = 32'd268468224;
      12271: inst = 32'd201345398;
      12272: inst = 32'd203489279;
      12273: inst = 32'd471859200;
      12274: inst = 32'd136314880;
      12275: inst = 32'd268468224;
      12276: inst = 32'd201345399;
      12277: inst = 32'd203489279;
      12278: inst = 32'd471859200;
      12279: inst = 32'd136314880;
      12280: inst = 32'd268468224;
      12281: inst = 32'd201345400;
      12282: inst = 32'd203489279;
      12283: inst = 32'd471859200;
      12284: inst = 32'd136314880;
      12285: inst = 32'd268468224;
      12286: inst = 32'd201345401;
      12287: inst = 32'd203489279;
      12288: inst = 32'd471859200;
      12289: inst = 32'd136314880;
      12290: inst = 32'd268468224;
      12291: inst = 32'd201345402;
      12292: inst = 32'd203489279;
      12293: inst = 32'd471859200;
      12294: inst = 32'd136314880;
      12295: inst = 32'd268468224;
      12296: inst = 32'd201345403;
      12297: inst = 32'd203489279;
      12298: inst = 32'd471859200;
      12299: inst = 32'd136314880;
      12300: inst = 32'd268468224;
      12301: inst = 32'd201345404;
      12302: inst = 32'd203489279;
      12303: inst = 32'd471859200;
      12304: inst = 32'd136314880;
      12305: inst = 32'd268468224;
      12306: inst = 32'd201345405;
      12307: inst = 32'd203489279;
      12308: inst = 32'd471859200;
      12309: inst = 32'd136314880;
      12310: inst = 32'd268468224;
      12311: inst = 32'd201345406;
      12312: inst = 32'd203489279;
      12313: inst = 32'd471859200;
      12314: inst = 32'd136314880;
      12315: inst = 32'd268468224;
      12316: inst = 32'd201345407;
      12317: inst = 32'd203489279;
      12318: inst = 32'd471859200;
      12319: inst = 32'd136314880;
      12320: inst = 32'd268468224;
      12321: inst = 32'd201345408;
      12322: inst = 32'd203489279;
      12323: inst = 32'd471859200;
      12324: inst = 32'd136314880;
      12325: inst = 32'd268468224;
      12326: inst = 32'd201345409;
      12327: inst = 32'd203489279;
      12328: inst = 32'd471859200;
      12329: inst = 32'd136314880;
      12330: inst = 32'd268468224;
      12331: inst = 32'd201345410;
      12332: inst = 32'd203489279;
      12333: inst = 32'd471859200;
      12334: inst = 32'd136314880;
      12335: inst = 32'd268468224;
      12336: inst = 32'd201345411;
      12337: inst = 32'd203489279;
      12338: inst = 32'd471859200;
      12339: inst = 32'd136314880;
      12340: inst = 32'd268468224;
      12341: inst = 32'd201345412;
      12342: inst = 32'd203484854;
      12343: inst = 32'd471859200;
      12344: inst = 32'd136314880;
      12345: inst = 32'd268468224;
      12346: inst = 32'd201345413;
      12347: inst = 32'd203484854;
      12348: inst = 32'd471859200;
      12349: inst = 32'd136314880;
      12350: inst = 32'd268468224;
      12351: inst = 32'd201345414;
      12352: inst = 32'd203484854;
      12353: inst = 32'd471859200;
      12354: inst = 32'd136314880;
      12355: inst = 32'd268468224;
      12356: inst = 32'd201345415;
      12357: inst = 32'd203484854;
      12358: inst = 32'd471859200;
      12359: inst = 32'd136314880;
      12360: inst = 32'd268468224;
      12361: inst = 32'd201345416;
      12362: inst = 32'd203484854;
      12363: inst = 32'd471859200;
      12364: inst = 32'd136314880;
      12365: inst = 32'd268468224;
      12366: inst = 32'd201345417;
      12367: inst = 32'd203484854;
      12368: inst = 32'd471859200;
      12369: inst = 32'd136314880;
      12370: inst = 32'd268468224;
      12371: inst = 32'd201345418;
      12372: inst = 32'd203484854;
      12373: inst = 32'd471859200;
      12374: inst = 32'd136314880;
      12375: inst = 32'd268468224;
      12376: inst = 32'd201345419;
      12377: inst = 32'd203484854;
      12378: inst = 32'd471859200;
      12379: inst = 32'd136314880;
      12380: inst = 32'd268468224;
      12381: inst = 32'd201345420;
      12382: inst = 32'd203484854;
      12383: inst = 32'd471859200;
      12384: inst = 32'd136314880;
      12385: inst = 32'd268468224;
      12386: inst = 32'd201345421;
      12387: inst = 32'd203484854;
      12388: inst = 32'd471859200;
      12389: inst = 32'd136314880;
      12390: inst = 32'd268468224;
      12391: inst = 32'd201345422;
      12392: inst = 32'd203484854;
      12393: inst = 32'd471859200;
      12394: inst = 32'd136314880;
      12395: inst = 32'd268468224;
      12396: inst = 32'd201345423;
      12397: inst = 32'd203473634;
      12398: inst = 32'd471859200;
      12399: inst = 32'd136314880;
      12400: inst = 32'd268468224;
      12401: inst = 32'd201345424;
      12402: inst = 32'd203480005;
      12403: inst = 32'd471859200;
      12404: inst = 32'd136314880;
      12405: inst = 32'd268468224;
      12406: inst = 32'd201345425;
      12407: inst = 32'd203480005;
      12408: inst = 32'd471859200;
      12409: inst = 32'd136314880;
      12410: inst = 32'd268468224;
      12411: inst = 32'd201345426;
      12412: inst = 32'd203489279;
      12413: inst = 32'd471859200;
      12414: inst = 32'd136314880;
      12415: inst = 32'd268468224;
      12416: inst = 32'd201345427;
      12417: inst = 32'd203485052;
      12418: inst = 32'd471859200;
      12419: inst = 32'd136314880;
      12420: inst = 32'd268468224;
      12421: inst = 32'd201345428;
      12422: inst = 32'd203485052;
      12423: inst = 32'd471859200;
      12424: inst = 32'd136314880;
      12425: inst = 32'd268468224;
      12426: inst = 32'd201345429;
      12427: inst = 32'd203485052;
      12428: inst = 32'd471859200;
      12429: inst = 32'd136314880;
      12430: inst = 32'd268468224;
      12431: inst = 32'd201345430;
      12432: inst = 32'd203480005;
      12433: inst = 32'd471859200;
      12434: inst = 32'd136314880;
      12435: inst = 32'd268468224;
      12436: inst = 32'd201345431;
      12437: inst = 32'd203480005;
      12438: inst = 32'd471859200;
      12439: inst = 32'd136314880;
      12440: inst = 32'd268468224;
      12441: inst = 32'd201345432;
      12442: inst = 32'd203480005;
      12443: inst = 32'd471859200;
      12444: inst = 32'd136314880;
      12445: inst = 32'd268468224;
      12446: inst = 32'd201345433;
      12447: inst = 32'd203480005;
      12448: inst = 32'd471859200;
      12449: inst = 32'd136314880;
      12450: inst = 32'd268468224;
      12451: inst = 32'd201345434;
      12452: inst = 32'd203480005;
      12453: inst = 32'd471859200;
      12454: inst = 32'd136314880;
      12455: inst = 32'd268468224;
      12456: inst = 32'd201345435;
      12457: inst = 32'd203480005;
      12458: inst = 32'd471859200;
      12459: inst = 32'd136314880;
      12460: inst = 32'd268468224;
      12461: inst = 32'd201345436;
      12462: inst = 32'd203480005;
      12463: inst = 32'd471859200;
      12464: inst = 32'd136314880;
      12465: inst = 32'd268468224;
      12466: inst = 32'd201345437;
      12467: inst = 32'd203480005;
      12468: inst = 32'd471859200;
      12469: inst = 32'd136314880;
      12470: inst = 32'd268468224;
      12471: inst = 32'd201345438;
      12472: inst = 32'd203480005;
      12473: inst = 32'd471859200;
      12474: inst = 32'd136314880;
      12475: inst = 32'd268468224;
      12476: inst = 32'd201345439;
      12477: inst = 32'd203473634;
      12478: inst = 32'd471859200;
      12479: inst = 32'd136314880;
      12480: inst = 32'd268468224;
      12481: inst = 32'd201345440;
      12482: inst = 32'd203484854;
      12483: inst = 32'd471859200;
      12484: inst = 32'd136314880;
      12485: inst = 32'd268468224;
      12486: inst = 32'd201345441;
      12487: inst = 32'd203484854;
      12488: inst = 32'd471859200;
      12489: inst = 32'd136314880;
      12490: inst = 32'd268468224;
      12491: inst = 32'd201345442;
      12492: inst = 32'd203484854;
      12493: inst = 32'd471859200;
      12494: inst = 32'd136314880;
      12495: inst = 32'd268468224;
      12496: inst = 32'd201345443;
      12497: inst = 32'd203484854;
      12498: inst = 32'd471859200;
      12499: inst = 32'd136314880;
      12500: inst = 32'd268468224;
      12501: inst = 32'd201345444;
      12502: inst = 32'd203484854;
      12503: inst = 32'd471859200;
      12504: inst = 32'd136314880;
      12505: inst = 32'd268468224;
      12506: inst = 32'd201345445;
      12507: inst = 32'd203484854;
      12508: inst = 32'd471859200;
      12509: inst = 32'd136314880;
      12510: inst = 32'd268468224;
      12511: inst = 32'd201345446;
      12512: inst = 32'd203484854;
      12513: inst = 32'd471859200;
      12514: inst = 32'd136314880;
      12515: inst = 32'd268468224;
      12516: inst = 32'd201345447;
      12517: inst = 32'd203484854;
      12518: inst = 32'd471859200;
      12519: inst = 32'd136314880;
      12520: inst = 32'd268468224;
      12521: inst = 32'd201345448;
      12522: inst = 32'd203484854;
      12523: inst = 32'd471859200;
      12524: inst = 32'd136314880;
      12525: inst = 32'd268468224;
      12526: inst = 32'd201345449;
      12527: inst = 32'd203484854;
      12528: inst = 32'd471859200;
      12529: inst = 32'd136314880;
      12530: inst = 32'd268468224;
      12531: inst = 32'd201345450;
      12532: inst = 32'd203484854;
      12533: inst = 32'd471859200;
      12534: inst = 32'd136314880;
      12535: inst = 32'd268468224;
      12536: inst = 32'd201345451;
      12537: inst = 32'd203484854;
      12538: inst = 32'd471859200;
      12539: inst = 32'd136314880;
      12540: inst = 32'd268468224;
      12541: inst = 32'd201345452;
      12542: inst = 32'd203484854;
      12543: inst = 32'd471859200;
      12544: inst = 32'd136314880;
      12545: inst = 32'd268468224;
      12546: inst = 32'd201345453;
      12547: inst = 32'd203484854;
      12548: inst = 32'd471859200;
      12549: inst = 32'd136314880;
      12550: inst = 32'd268468224;
      12551: inst = 32'd201345454;
      12552: inst = 32'd203484854;
      12553: inst = 32'd471859200;
      12554: inst = 32'd136314880;
      12555: inst = 32'd268468224;
      12556: inst = 32'd201345455;
      12557: inst = 32'd203484854;
      12558: inst = 32'd471859200;
      12559: inst = 32'd136314880;
      12560: inst = 32'd268468224;
      12561: inst = 32'd201345456;
      12562: inst = 32'd203484854;
      12563: inst = 32'd471859200;
      12564: inst = 32'd136314880;
      12565: inst = 32'd268468224;
      12566: inst = 32'd201345457;
      12567: inst = 32'd203484854;
      12568: inst = 32'd471859200;
      12569: inst = 32'd136314880;
      12570: inst = 32'd268468224;
      12571: inst = 32'd201345458;
      12572: inst = 32'd203484854;
      12573: inst = 32'd471859200;
      12574: inst = 32'd136314880;
      12575: inst = 32'd268468224;
      12576: inst = 32'd201345459;
      12577: inst = 32'd203484854;
      12578: inst = 32'd471859200;
      12579: inst = 32'd136314880;
      12580: inst = 32'd268468224;
      12581: inst = 32'd201345460;
      12582: inst = 32'd203484854;
      12583: inst = 32'd471859200;
      12584: inst = 32'd136314880;
      12585: inst = 32'd268468224;
      12586: inst = 32'd201345461;
      12587: inst = 32'd203484854;
      12588: inst = 32'd471859200;
      12589: inst = 32'd136314880;
      12590: inst = 32'd268468224;
      12591: inst = 32'd201345462;
      12592: inst = 32'd203484854;
      12593: inst = 32'd471859200;
      12594: inst = 32'd136314880;
      12595: inst = 32'd268468224;
      12596: inst = 32'd201345463;
      12597: inst = 32'd203484854;
      12598: inst = 32'd471859200;
      12599: inst = 32'd136314880;
      12600: inst = 32'd268468224;
      12601: inst = 32'd201345464;
      12602: inst = 32'd203484854;
      12603: inst = 32'd471859200;
      12604: inst = 32'd136314880;
      12605: inst = 32'd268468224;
      12606: inst = 32'd201345465;
      12607: inst = 32'd203484854;
      12608: inst = 32'd471859200;
      12609: inst = 32'd136314880;
      12610: inst = 32'd268468224;
      12611: inst = 32'd201345466;
      12612: inst = 32'd203484854;
      12613: inst = 32'd471859200;
      12614: inst = 32'd136314880;
      12615: inst = 32'd268468224;
      12616: inst = 32'd201345467;
      12617: inst = 32'd203484854;
      12618: inst = 32'd471859200;
      12619: inst = 32'd136314880;
      12620: inst = 32'd268468224;
      12621: inst = 32'd201345468;
      12622: inst = 32'd203489279;
      12623: inst = 32'd471859200;
      12624: inst = 32'd136314880;
      12625: inst = 32'd268468224;
      12626: inst = 32'd201345469;
      12627: inst = 32'd203489279;
      12628: inst = 32'd471859200;
      12629: inst = 32'd136314880;
      12630: inst = 32'd268468224;
      12631: inst = 32'd201345470;
      12632: inst = 32'd203489279;
      12633: inst = 32'd471859200;
      12634: inst = 32'd136314880;
      12635: inst = 32'd268468224;
      12636: inst = 32'd201345471;
      12637: inst = 32'd203489279;
      12638: inst = 32'd471859200;
      12639: inst = 32'd136314880;
      12640: inst = 32'd268468224;
      12641: inst = 32'd201345472;
      12642: inst = 32'd203489279;
      12643: inst = 32'd471859200;
      12644: inst = 32'd136314880;
      12645: inst = 32'd268468224;
      12646: inst = 32'd201345473;
      12647: inst = 32'd203489279;
      12648: inst = 32'd471859200;
      12649: inst = 32'd136314880;
      12650: inst = 32'd268468224;
      12651: inst = 32'd201345474;
      12652: inst = 32'd203489279;
      12653: inst = 32'd471859200;
      12654: inst = 32'd136314880;
      12655: inst = 32'd268468224;
      12656: inst = 32'd201345475;
      12657: inst = 32'd203489279;
      12658: inst = 32'd471859200;
      12659: inst = 32'd136314880;
      12660: inst = 32'd268468224;
      12661: inst = 32'd201345476;
      12662: inst = 32'd203489279;
      12663: inst = 32'd471859200;
      12664: inst = 32'd136314880;
      12665: inst = 32'd268468224;
      12666: inst = 32'd201345477;
      12667: inst = 32'd203489279;
      12668: inst = 32'd471859200;
      12669: inst = 32'd136314880;
      12670: inst = 32'd268468224;
      12671: inst = 32'd201345478;
      12672: inst = 32'd203489279;
      12673: inst = 32'd471859200;
      12674: inst = 32'd136314880;
      12675: inst = 32'd268468224;
      12676: inst = 32'd201345479;
      12677: inst = 32'd203489279;
      12678: inst = 32'd471859200;
      12679: inst = 32'd136314880;
      12680: inst = 32'd268468224;
      12681: inst = 32'd201345480;
      12682: inst = 32'd203489279;
      12683: inst = 32'd471859200;
      12684: inst = 32'd136314880;
      12685: inst = 32'd268468224;
      12686: inst = 32'd201345481;
      12687: inst = 32'd203489279;
      12688: inst = 32'd471859200;
      12689: inst = 32'd136314880;
      12690: inst = 32'd268468224;
      12691: inst = 32'd201345482;
      12692: inst = 32'd203489279;
      12693: inst = 32'd471859200;
      12694: inst = 32'd136314880;
      12695: inst = 32'd268468224;
      12696: inst = 32'd201345483;
      12697: inst = 32'd203489279;
      12698: inst = 32'd471859200;
      12699: inst = 32'd136314880;
      12700: inst = 32'd268468224;
      12701: inst = 32'd201345484;
      12702: inst = 32'd203489279;
      12703: inst = 32'd471859200;
      12704: inst = 32'd136314880;
      12705: inst = 32'd268468224;
      12706: inst = 32'd201345485;
      12707: inst = 32'd203489279;
      12708: inst = 32'd471859200;
      12709: inst = 32'd136314880;
      12710: inst = 32'd268468224;
      12711: inst = 32'd201345486;
      12712: inst = 32'd203489279;
      12713: inst = 32'd471859200;
      12714: inst = 32'd136314880;
      12715: inst = 32'd268468224;
      12716: inst = 32'd201345487;
      12717: inst = 32'd203489279;
      12718: inst = 32'd471859200;
      12719: inst = 32'd136314880;
      12720: inst = 32'd268468224;
      12721: inst = 32'd201345488;
      12722: inst = 32'd203489279;
      12723: inst = 32'd471859200;
      12724: inst = 32'd136314880;
      12725: inst = 32'd268468224;
      12726: inst = 32'd201345489;
      12727: inst = 32'd203489279;
      12728: inst = 32'd471859200;
      12729: inst = 32'd136314880;
      12730: inst = 32'd268468224;
      12731: inst = 32'd201345490;
      12732: inst = 32'd203489279;
      12733: inst = 32'd471859200;
      12734: inst = 32'd136314880;
      12735: inst = 32'd268468224;
      12736: inst = 32'd201345491;
      12737: inst = 32'd203489279;
      12738: inst = 32'd471859200;
      12739: inst = 32'd136314880;
      12740: inst = 32'd268468224;
      12741: inst = 32'd201345492;
      12742: inst = 32'd203489279;
      12743: inst = 32'd471859200;
      12744: inst = 32'd136314880;
      12745: inst = 32'd268468224;
      12746: inst = 32'd201345493;
      12747: inst = 32'd203489279;
      12748: inst = 32'd471859200;
      12749: inst = 32'd136314880;
      12750: inst = 32'd268468224;
      12751: inst = 32'd201345494;
      12752: inst = 32'd203489279;
      12753: inst = 32'd471859200;
      12754: inst = 32'd136314880;
      12755: inst = 32'd268468224;
      12756: inst = 32'd201345495;
      12757: inst = 32'd203489279;
      12758: inst = 32'd471859200;
      12759: inst = 32'd136314880;
      12760: inst = 32'd268468224;
      12761: inst = 32'd201345496;
      12762: inst = 32'd203489279;
      12763: inst = 32'd471859200;
      12764: inst = 32'd136314880;
      12765: inst = 32'd268468224;
      12766: inst = 32'd201345497;
      12767: inst = 32'd203489279;
      12768: inst = 32'd471859200;
      12769: inst = 32'd136314880;
      12770: inst = 32'd268468224;
      12771: inst = 32'd201345498;
      12772: inst = 32'd203489279;
      12773: inst = 32'd471859200;
      12774: inst = 32'd136314880;
      12775: inst = 32'd268468224;
      12776: inst = 32'd201345499;
      12777: inst = 32'd203489279;
      12778: inst = 32'd471859200;
      12779: inst = 32'd136314880;
      12780: inst = 32'd268468224;
      12781: inst = 32'd201345500;
      12782: inst = 32'd203489279;
      12783: inst = 32'd471859200;
      12784: inst = 32'd136314880;
      12785: inst = 32'd268468224;
      12786: inst = 32'd201345501;
      12787: inst = 32'd203489279;
      12788: inst = 32'd471859200;
      12789: inst = 32'd136314880;
      12790: inst = 32'd268468224;
      12791: inst = 32'd201345502;
      12792: inst = 32'd203489279;
      12793: inst = 32'd471859200;
      12794: inst = 32'd136314880;
      12795: inst = 32'd268468224;
      12796: inst = 32'd201345503;
      12797: inst = 32'd203489279;
      12798: inst = 32'd471859200;
      12799: inst = 32'd136314880;
      12800: inst = 32'd268468224;
      12801: inst = 32'd201345504;
      12802: inst = 32'd203489279;
      12803: inst = 32'd471859200;
      12804: inst = 32'd136314880;
      12805: inst = 32'd268468224;
      12806: inst = 32'd201345505;
      12807: inst = 32'd203489279;
      12808: inst = 32'd471859200;
      12809: inst = 32'd136314880;
      12810: inst = 32'd268468224;
      12811: inst = 32'd201345506;
      12812: inst = 32'd203489279;
      12813: inst = 32'd471859200;
      12814: inst = 32'd136314880;
      12815: inst = 32'd268468224;
      12816: inst = 32'd201345507;
      12817: inst = 32'd203489279;
      12818: inst = 32'd471859200;
      12819: inst = 32'd136314880;
      12820: inst = 32'd268468224;
      12821: inst = 32'd201345508;
      12822: inst = 32'd203484854;
      12823: inst = 32'd471859200;
      12824: inst = 32'd136314880;
      12825: inst = 32'd268468224;
      12826: inst = 32'd201345509;
      12827: inst = 32'd203484854;
      12828: inst = 32'd471859200;
      12829: inst = 32'd136314880;
      12830: inst = 32'd268468224;
      12831: inst = 32'd201345510;
      12832: inst = 32'd203484854;
      12833: inst = 32'd471859200;
      12834: inst = 32'd136314880;
      12835: inst = 32'd268468224;
      12836: inst = 32'd201345511;
      12837: inst = 32'd203484854;
      12838: inst = 32'd471859200;
      12839: inst = 32'd136314880;
      12840: inst = 32'd268468224;
      12841: inst = 32'd201345512;
      12842: inst = 32'd203484854;
      12843: inst = 32'd471859200;
      12844: inst = 32'd136314880;
      12845: inst = 32'd268468224;
      12846: inst = 32'd201345513;
      12847: inst = 32'd203484854;
      12848: inst = 32'd471859200;
      12849: inst = 32'd136314880;
      12850: inst = 32'd268468224;
      12851: inst = 32'd201345514;
      12852: inst = 32'd203484854;
      12853: inst = 32'd471859200;
      12854: inst = 32'd136314880;
      12855: inst = 32'd268468224;
      12856: inst = 32'd201345515;
      12857: inst = 32'd203484854;
      12858: inst = 32'd471859200;
      12859: inst = 32'd136314880;
      12860: inst = 32'd268468224;
      12861: inst = 32'd201345516;
      12862: inst = 32'd203484854;
      12863: inst = 32'd471859200;
      12864: inst = 32'd136314880;
      12865: inst = 32'd268468224;
      12866: inst = 32'd201345517;
      12867: inst = 32'd203484854;
      12868: inst = 32'd471859200;
      12869: inst = 32'd136314880;
      12870: inst = 32'd268468224;
      12871: inst = 32'd201345518;
      12872: inst = 32'd203484854;
      12873: inst = 32'd471859200;
      12874: inst = 32'd136314880;
      12875: inst = 32'd268468224;
      12876: inst = 32'd201345519;
      12877: inst = 32'd203473634;
      12878: inst = 32'd471859200;
      12879: inst = 32'd136314880;
      12880: inst = 32'd268468224;
      12881: inst = 32'd201345520;
      12882: inst = 32'd203480005;
      12883: inst = 32'd471859200;
      12884: inst = 32'd136314880;
      12885: inst = 32'd268468224;
      12886: inst = 32'd201345521;
      12887: inst = 32'd203480005;
      12888: inst = 32'd471859200;
      12889: inst = 32'd136314880;
      12890: inst = 32'd268468224;
      12891: inst = 32'd201345522;
      12892: inst = 32'd203489279;
      12893: inst = 32'd471859200;
      12894: inst = 32'd136314880;
      12895: inst = 32'd268468224;
      12896: inst = 32'd201345523;
      12897: inst = 32'd203485052;
      12898: inst = 32'd471859200;
      12899: inst = 32'd136314880;
      12900: inst = 32'd268468224;
      12901: inst = 32'd201345524;
      12902: inst = 32'd203485052;
      12903: inst = 32'd471859200;
      12904: inst = 32'd136314880;
      12905: inst = 32'd268468224;
      12906: inst = 32'd201345525;
      12907: inst = 32'd203485052;
      12908: inst = 32'd471859200;
      12909: inst = 32'd136314880;
      12910: inst = 32'd268468224;
      12911: inst = 32'd201345526;
      12912: inst = 32'd203480005;
      12913: inst = 32'd471859200;
      12914: inst = 32'd136314880;
      12915: inst = 32'd268468224;
      12916: inst = 32'd201345527;
      12917: inst = 32'd203480005;
      12918: inst = 32'd471859200;
      12919: inst = 32'd136314880;
      12920: inst = 32'd268468224;
      12921: inst = 32'd201345528;
      12922: inst = 32'd203480005;
      12923: inst = 32'd471859200;
      12924: inst = 32'd136314880;
      12925: inst = 32'd268468224;
      12926: inst = 32'd201345529;
      12927: inst = 32'd203480005;
      12928: inst = 32'd471859200;
      12929: inst = 32'd136314880;
      12930: inst = 32'd268468224;
      12931: inst = 32'd201345530;
      12932: inst = 32'd203480005;
      12933: inst = 32'd471859200;
      12934: inst = 32'd136314880;
      12935: inst = 32'd268468224;
      12936: inst = 32'd201345531;
      12937: inst = 32'd203480005;
      12938: inst = 32'd471859200;
      12939: inst = 32'd136314880;
      12940: inst = 32'd268468224;
      12941: inst = 32'd201345532;
      12942: inst = 32'd203480005;
      12943: inst = 32'd471859200;
      12944: inst = 32'd136314880;
      12945: inst = 32'd268468224;
      12946: inst = 32'd201345533;
      12947: inst = 32'd203480005;
      12948: inst = 32'd471859200;
      12949: inst = 32'd136314880;
      12950: inst = 32'd268468224;
      12951: inst = 32'd201345534;
      12952: inst = 32'd203480005;
      12953: inst = 32'd471859200;
      12954: inst = 32'd136314880;
      12955: inst = 32'd268468224;
      12956: inst = 32'd201345535;
      12957: inst = 32'd203473634;
      12958: inst = 32'd471859200;
      12959: inst = 32'd136314880;
      12960: inst = 32'd268468224;
      12961: inst = 32'd201345536;
      12962: inst = 32'd203484854;
      12963: inst = 32'd471859200;
      12964: inst = 32'd136314880;
      12965: inst = 32'd268468224;
      12966: inst = 32'd201345537;
      12967: inst = 32'd203484854;
      12968: inst = 32'd471859200;
      12969: inst = 32'd136314880;
      12970: inst = 32'd268468224;
      12971: inst = 32'd201345538;
      12972: inst = 32'd203484854;
      12973: inst = 32'd471859200;
      12974: inst = 32'd136314880;
      12975: inst = 32'd268468224;
      12976: inst = 32'd201345539;
      12977: inst = 32'd203484854;
      12978: inst = 32'd471859200;
      12979: inst = 32'd136314880;
      12980: inst = 32'd268468224;
      12981: inst = 32'd201345540;
      12982: inst = 32'd203484854;
      12983: inst = 32'd471859200;
      12984: inst = 32'd136314880;
      12985: inst = 32'd268468224;
      12986: inst = 32'd201345541;
      12987: inst = 32'd203484854;
      12988: inst = 32'd471859200;
      12989: inst = 32'd136314880;
      12990: inst = 32'd268468224;
      12991: inst = 32'd201345542;
      12992: inst = 32'd203484854;
      12993: inst = 32'd471859200;
      12994: inst = 32'd136314880;
      12995: inst = 32'd268468224;
      12996: inst = 32'd201345543;
      12997: inst = 32'd203484854;
      12998: inst = 32'd471859200;
      12999: inst = 32'd136314880;
      13000: inst = 32'd268468224;
      13001: inst = 32'd201345544;
      13002: inst = 32'd203484887;
      13003: inst = 32'd471859200;
      13004: inst = 32'd136314880;
      13005: inst = 32'd268468224;
      13006: inst = 32'd201345545;
      13007: inst = 32'd203482874;
      13008: inst = 32'd471859200;
      13009: inst = 32'd136314880;
      13010: inst = 32'd268468224;
      13011: inst = 32'd201345546;
      13012: inst = 32'd203482875;
      13013: inst = 32'd471859200;
      13014: inst = 32'd136314880;
      13015: inst = 32'd268468224;
      13016: inst = 32'd201345547;
      13017: inst = 32'd203480827;
      13018: inst = 32'd471859200;
      13019: inst = 32'd136314880;
      13020: inst = 32'd268468224;
      13021: inst = 32'd201345548;
      13022: inst = 32'd203482875;
      13023: inst = 32'd471859200;
      13024: inst = 32'd136314880;
      13025: inst = 32'd268468224;
      13026: inst = 32'd201345549;
      13027: inst = 32'd203482874;
      13028: inst = 32'd471859200;
      13029: inst = 32'd136314880;
      13030: inst = 32'd268468224;
      13031: inst = 32'd201345550;
      13032: inst = 32'd203484887;
      13033: inst = 32'd471859200;
      13034: inst = 32'd136314880;
      13035: inst = 32'd268468224;
      13036: inst = 32'd201345551;
      13037: inst = 32'd203484854;
      13038: inst = 32'd471859200;
      13039: inst = 32'd136314880;
      13040: inst = 32'd268468224;
      13041: inst = 32'd201345552;
      13042: inst = 32'd203484854;
      13043: inst = 32'd471859200;
      13044: inst = 32'd136314880;
      13045: inst = 32'd268468224;
      13046: inst = 32'd201345553;
      13047: inst = 32'd203484854;
      13048: inst = 32'd471859200;
      13049: inst = 32'd136314880;
      13050: inst = 32'd268468224;
      13051: inst = 32'd201345554;
      13052: inst = 32'd203484854;
      13053: inst = 32'd471859200;
      13054: inst = 32'd136314880;
      13055: inst = 32'd268468224;
      13056: inst = 32'd201345555;
      13057: inst = 32'd203484854;
      13058: inst = 32'd471859200;
      13059: inst = 32'd136314880;
      13060: inst = 32'd268468224;
      13061: inst = 32'd201345556;
      13062: inst = 32'd203484854;
      13063: inst = 32'd471859200;
      13064: inst = 32'd136314880;
      13065: inst = 32'd268468224;
      13066: inst = 32'd201345557;
      13067: inst = 32'd203484854;
      13068: inst = 32'd471859200;
      13069: inst = 32'd136314880;
      13070: inst = 32'd268468224;
      13071: inst = 32'd201345558;
      13072: inst = 32'd203484854;
      13073: inst = 32'd471859200;
      13074: inst = 32'd136314880;
      13075: inst = 32'd268468224;
      13076: inst = 32'd201345559;
      13077: inst = 32'd203484854;
      13078: inst = 32'd471859200;
      13079: inst = 32'd136314880;
      13080: inst = 32'd268468224;
      13081: inst = 32'd201345560;
      13082: inst = 32'd203484854;
      13083: inst = 32'd471859200;
      13084: inst = 32'd136314880;
      13085: inst = 32'd268468224;
      13086: inst = 32'd201345561;
      13087: inst = 32'd203484854;
      13088: inst = 32'd471859200;
      13089: inst = 32'd136314880;
      13090: inst = 32'd268468224;
      13091: inst = 32'd201345562;
      13092: inst = 32'd203484854;
      13093: inst = 32'd471859200;
      13094: inst = 32'd136314880;
      13095: inst = 32'd268468224;
      13096: inst = 32'd201345563;
      13097: inst = 32'd203484854;
      13098: inst = 32'd471859200;
      13099: inst = 32'd136314880;
      13100: inst = 32'd268468224;
      13101: inst = 32'd201345564;
      13102: inst = 32'd203489279;
      13103: inst = 32'd471859200;
      13104: inst = 32'd136314880;
      13105: inst = 32'd268468224;
      13106: inst = 32'd201345565;
      13107: inst = 32'd203489279;
      13108: inst = 32'd471859200;
      13109: inst = 32'd136314880;
      13110: inst = 32'd268468224;
      13111: inst = 32'd201345566;
      13112: inst = 32'd203489279;
      13113: inst = 32'd471859200;
      13114: inst = 32'd136314880;
      13115: inst = 32'd268468224;
      13116: inst = 32'd201345567;
      13117: inst = 32'd203489279;
      13118: inst = 32'd471859200;
      13119: inst = 32'd136314880;
      13120: inst = 32'd268468224;
      13121: inst = 32'd201345568;
      13122: inst = 32'd203489279;
      13123: inst = 32'd471859200;
      13124: inst = 32'd136314880;
      13125: inst = 32'd268468224;
      13126: inst = 32'd201345569;
      13127: inst = 32'd203489279;
      13128: inst = 32'd471859200;
      13129: inst = 32'd136314880;
      13130: inst = 32'd268468224;
      13131: inst = 32'd201345570;
      13132: inst = 32'd203489279;
      13133: inst = 32'd471859200;
      13134: inst = 32'd136314880;
      13135: inst = 32'd268468224;
      13136: inst = 32'd201345571;
      13137: inst = 32'd203489279;
      13138: inst = 32'd471859200;
      13139: inst = 32'd136314880;
      13140: inst = 32'd268468224;
      13141: inst = 32'd201345572;
      13142: inst = 32'd203489279;
      13143: inst = 32'd471859200;
      13144: inst = 32'd136314880;
      13145: inst = 32'd268468224;
      13146: inst = 32'd201345573;
      13147: inst = 32'd203489279;
      13148: inst = 32'd471859200;
      13149: inst = 32'd136314880;
      13150: inst = 32'd268468224;
      13151: inst = 32'd201345574;
      13152: inst = 32'd203489279;
      13153: inst = 32'd471859200;
      13154: inst = 32'd136314880;
      13155: inst = 32'd268468224;
      13156: inst = 32'd201345575;
      13157: inst = 32'd203489279;
      13158: inst = 32'd471859200;
      13159: inst = 32'd136314880;
      13160: inst = 32'd268468224;
      13161: inst = 32'd201345576;
      13162: inst = 32'd203489279;
      13163: inst = 32'd471859200;
      13164: inst = 32'd136314880;
      13165: inst = 32'd268468224;
      13166: inst = 32'd201345577;
      13167: inst = 32'd203489279;
      13168: inst = 32'd471859200;
      13169: inst = 32'd136314880;
      13170: inst = 32'd268468224;
      13171: inst = 32'd201345578;
      13172: inst = 32'd203489279;
      13173: inst = 32'd471859200;
      13174: inst = 32'd136314880;
      13175: inst = 32'd268468224;
      13176: inst = 32'd201345579;
      13177: inst = 32'd203489279;
      13178: inst = 32'd471859200;
      13179: inst = 32'd136314880;
      13180: inst = 32'd268468224;
      13181: inst = 32'd201345580;
      13182: inst = 32'd203489279;
      13183: inst = 32'd471859200;
      13184: inst = 32'd136314880;
      13185: inst = 32'd268468224;
      13186: inst = 32'd201345581;
      13187: inst = 32'd203489279;
      13188: inst = 32'd471859200;
      13189: inst = 32'd136314880;
      13190: inst = 32'd268468224;
      13191: inst = 32'd201345582;
      13192: inst = 32'd203489279;
      13193: inst = 32'd471859200;
      13194: inst = 32'd136314880;
      13195: inst = 32'd268468224;
      13196: inst = 32'd201345583;
      13197: inst = 32'd203489279;
      13198: inst = 32'd471859200;
      13199: inst = 32'd136314880;
      13200: inst = 32'd268468224;
      13201: inst = 32'd201345584;
      13202: inst = 32'd203489279;
      13203: inst = 32'd471859200;
      13204: inst = 32'd136314880;
      13205: inst = 32'd268468224;
      13206: inst = 32'd201345585;
      13207: inst = 32'd203489279;
      13208: inst = 32'd471859200;
      13209: inst = 32'd136314880;
      13210: inst = 32'd268468224;
      13211: inst = 32'd201345586;
      13212: inst = 32'd203489279;
      13213: inst = 32'd471859200;
      13214: inst = 32'd136314880;
      13215: inst = 32'd268468224;
      13216: inst = 32'd201345587;
      13217: inst = 32'd203489279;
      13218: inst = 32'd471859200;
      13219: inst = 32'd136314880;
      13220: inst = 32'd268468224;
      13221: inst = 32'd201345588;
      13222: inst = 32'd203489279;
      13223: inst = 32'd471859200;
      13224: inst = 32'd136314880;
      13225: inst = 32'd268468224;
      13226: inst = 32'd201345589;
      13227: inst = 32'd203489279;
      13228: inst = 32'd471859200;
      13229: inst = 32'd136314880;
      13230: inst = 32'd268468224;
      13231: inst = 32'd201345590;
      13232: inst = 32'd203489279;
      13233: inst = 32'd471859200;
      13234: inst = 32'd136314880;
      13235: inst = 32'd268468224;
      13236: inst = 32'd201345591;
      13237: inst = 32'd203489279;
      13238: inst = 32'd471859200;
      13239: inst = 32'd136314880;
      13240: inst = 32'd268468224;
      13241: inst = 32'd201345592;
      13242: inst = 32'd203489279;
      13243: inst = 32'd471859200;
      13244: inst = 32'd136314880;
      13245: inst = 32'd268468224;
      13246: inst = 32'd201345593;
      13247: inst = 32'd203489279;
      13248: inst = 32'd471859200;
      13249: inst = 32'd136314880;
      13250: inst = 32'd268468224;
      13251: inst = 32'd201345594;
      13252: inst = 32'd203489279;
      13253: inst = 32'd471859200;
      13254: inst = 32'd136314880;
      13255: inst = 32'd268468224;
      13256: inst = 32'd201345595;
      13257: inst = 32'd203489279;
      13258: inst = 32'd471859200;
      13259: inst = 32'd136314880;
      13260: inst = 32'd268468224;
      13261: inst = 32'd201345596;
      13262: inst = 32'd203489279;
      13263: inst = 32'd471859200;
      13264: inst = 32'd136314880;
      13265: inst = 32'd268468224;
      13266: inst = 32'd201345597;
      13267: inst = 32'd203489279;
      13268: inst = 32'd471859200;
      13269: inst = 32'd136314880;
      13270: inst = 32'd268468224;
      13271: inst = 32'd201345598;
      13272: inst = 32'd203489279;
      13273: inst = 32'd471859200;
      13274: inst = 32'd136314880;
      13275: inst = 32'd268468224;
      13276: inst = 32'd201345599;
      13277: inst = 32'd203489279;
      13278: inst = 32'd471859200;
      13279: inst = 32'd136314880;
      13280: inst = 32'd268468224;
      13281: inst = 32'd201345600;
      13282: inst = 32'd203489279;
      13283: inst = 32'd471859200;
      13284: inst = 32'd136314880;
      13285: inst = 32'd268468224;
      13286: inst = 32'd201345601;
      13287: inst = 32'd203489279;
      13288: inst = 32'd471859200;
      13289: inst = 32'd136314880;
      13290: inst = 32'd268468224;
      13291: inst = 32'd201345602;
      13292: inst = 32'd203489279;
      13293: inst = 32'd471859200;
      13294: inst = 32'd136314880;
      13295: inst = 32'd268468224;
      13296: inst = 32'd201345603;
      13297: inst = 32'd203489279;
      13298: inst = 32'd471859200;
      13299: inst = 32'd136314880;
      13300: inst = 32'd268468224;
      13301: inst = 32'd201345604;
      13302: inst = 32'd203484854;
      13303: inst = 32'd471859200;
      13304: inst = 32'd136314880;
      13305: inst = 32'd268468224;
      13306: inst = 32'd201345605;
      13307: inst = 32'd203484854;
      13308: inst = 32'd471859200;
      13309: inst = 32'd136314880;
      13310: inst = 32'd268468224;
      13311: inst = 32'd201345606;
      13312: inst = 32'd203484854;
      13313: inst = 32'd471859200;
      13314: inst = 32'd136314880;
      13315: inst = 32'd268468224;
      13316: inst = 32'd201345607;
      13317: inst = 32'd203484854;
      13318: inst = 32'd471859200;
      13319: inst = 32'd136314880;
      13320: inst = 32'd268468224;
      13321: inst = 32'd201345608;
      13322: inst = 32'd203484854;
      13323: inst = 32'd471859200;
      13324: inst = 32'd136314880;
      13325: inst = 32'd268468224;
      13326: inst = 32'd201345609;
      13327: inst = 32'd203484854;
      13328: inst = 32'd471859200;
      13329: inst = 32'd136314880;
      13330: inst = 32'd268468224;
      13331: inst = 32'd201345610;
      13332: inst = 32'd203484854;
      13333: inst = 32'd471859200;
      13334: inst = 32'd136314880;
      13335: inst = 32'd268468224;
      13336: inst = 32'd201345611;
      13337: inst = 32'd203484854;
      13338: inst = 32'd471859200;
      13339: inst = 32'd136314880;
      13340: inst = 32'd268468224;
      13341: inst = 32'd201345612;
      13342: inst = 32'd203484854;
      13343: inst = 32'd471859200;
      13344: inst = 32'd136314880;
      13345: inst = 32'd268468224;
      13346: inst = 32'd201345613;
      13347: inst = 32'd203484854;
      13348: inst = 32'd471859200;
      13349: inst = 32'd136314880;
      13350: inst = 32'd268468224;
      13351: inst = 32'd201345614;
      13352: inst = 32'd203484854;
      13353: inst = 32'd471859200;
      13354: inst = 32'd136314880;
      13355: inst = 32'd268468224;
      13356: inst = 32'd201345615;
      13357: inst = 32'd203473634;
      13358: inst = 32'd471859200;
      13359: inst = 32'd136314880;
      13360: inst = 32'd268468224;
      13361: inst = 32'd201345616;
      13362: inst = 32'd203480005;
      13363: inst = 32'd471859200;
      13364: inst = 32'd136314880;
      13365: inst = 32'd268468224;
      13366: inst = 32'd201345617;
      13367: inst = 32'd203480005;
      13368: inst = 32'd471859200;
      13369: inst = 32'd136314880;
      13370: inst = 32'd268468224;
      13371: inst = 32'd201345618;
      13372: inst = 32'd203489279;
      13373: inst = 32'd471859200;
      13374: inst = 32'd136314880;
      13375: inst = 32'd268468224;
      13376: inst = 32'd201345619;
      13377: inst = 32'd203485052;
      13378: inst = 32'd471859200;
      13379: inst = 32'd136314880;
      13380: inst = 32'd268468224;
      13381: inst = 32'd201345620;
      13382: inst = 32'd203485052;
      13383: inst = 32'd471859200;
      13384: inst = 32'd136314880;
      13385: inst = 32'd268468224;
      13386: inst = 32'd201345621;
      13387: inst = 32'd203485052;
      13388: inst = 32'd471859200;
      13389: inst = 32'd136314880;
      13390: inst = 32'd268468224;
      13391: inst = 32'd201345622;
      13392: inst = 32'd203480005;
      13393: inst = 32'd471859200;
      13394: inst = 32'd136314880;
      13395: inst = 32'd268468224;
      13396: inst = 32'd201345623;
      13397: inst = 32'd203480005;
      13398: inst = 32'd471859200;
      13399: inst = 32'd136314880;
      13400: inst = 32'd268468224;
      13401: inst = 32'd201345624;
      13402: inst = 32'd203480005;
      13403: inst = 32'd471859200;
      13404: inst = 32'd136314880;
      13405: inst = 32'd268468224;
      13406: inst = 32'd201345625;
      13407: inst = 32'd203480005;
      13408: inst = 32'd471859200;
      13409: inst = 32'd136314880;
      13410: inst = 32'd268468224;
      13411: inst = 32'd201345626;
      13412: inst = 32'd203480005;
      13413: inst = 32'd471859200;
      13414: inst = 32'd136314880;
      13415: inst = 32'd268468224;
      13416: inst = 32'd201345627;
      13417: inst = 32'd203480005;
      13418: inst = 32'd471859200;
      13419: inst = 32'd136314880;
      13420: inst = 32'd268468224;
      13421: inst = 32'd201345628;
      13422: inst = 32'd203480005;
      13423: inst = 32'd471859200;
      13424: inst = 32'd136314880;
      13425: inst = 32'd268468224;
      13426: inst = 32'd201345629;
      13427: inst = 32'd203480005;
      13428: inst = 32'd471859200;
      13429: inst = 32'd136314880;
      13430: inst = 32'd268468224;
      13431: inst = 32'd201345630;
      13432: inst = 32'd203480005;
      13433: inst = 32'd471859200;
      13434: inst = 32'd136314880;
      13435: inst = 32'd268468224;
      13436: inst = 32'd201345631;
      13437: inst = 32'd203473634;
      13438: inst = 32'd471859200;
      13439: inst = 32'd136314880;
      13440: inst = 32'd268468224;
      13441: inst = 32'd201345632;
      13442: inst = 32'd203484854;
      13443: inst = 32'd471859200;
      13444: inst = 32'd136314880;
      13445: inst = 32'd268468224;
      13446: inst = 32'd201345633;
      13447: inst = 32'd203484854;
      13448: inst = 32'd471859200;
      13449: inst = 32'd136314880;
      13450: inst = 32'd268468224;
      13451: inst = 32'd201345634;
      13452: inst = 32'd203484854;
      13453: inst = 32'd471859200;
      13454: inst = 32'd136314880;
      13455: inst = 32'd268468224;
      13456: inst = 32'd201345635;
      13457: inst = 32'd203484854;
      13458: inst = 32'd471859200;
      13459: inst = 32'd136314880;
      13460: inst = 32'd268468224;
      13461: inst = 32'd201345636;
      13462: inst = 32'd203484854;
      13463: inst = 32'd471859200;
      13464: inst = 32'd136314880;
      13465: inst = 32'd268468224;
      13466: inst = 32'd201345637;
      13467: inst = 32'd203484854;
      13468: inst = 32'd471859200;
      13469: inst = 32'd136314880;
      13470: inst = 32'd268468224;
      13471: inst = 32'd201345638;
      13472: inst = 32'd203484854;
      13473: inst = 32'd471859200;
      13474: inst = 32'd136314880;
      13475: inst = 32'd268468224;
      13476: inst = 32'd201345639;
      13477: inst = 32'd203484888;
      13478: inst = 32'd471859200;
      13479: inst = 32'd136314880;
      13480: inst = 32'd268468224;
      13481: inst = 32'd201345640;
      13482: inst = 32'd203480827;
      13483: inst = 32'd471859200;
      13484: inst = 32'd136314880;
      13485: inst = 32'd268468224;
      13486: inst = 32'd201345641;
      13487: inst = 32'd203480827;
      13488: inst = 32'd471859200;
      13489: inst = 32'd136314880;
      13490: inst = 32'd268468224;
      13491: inst = 32'd201345642;
      13492: inst = 32'd203480827;
      13493: inst = 32'd471859200;
      13494: inst = 32'd136314880;
      13495: inst = 32'd268468224;
      13496: inst = 32'd201345643;
      13497: inst = 32'd203480827;
      13498: inst = 32'd471859200;
      13499: inst = 32'd136314880;
      13500: inst = 32'd268468224;
      13501: inst = 32'd201345644;
      13502: inst = 32'd203480827;
      13503: inst = 32'd471859200;
      13504: inst = 32'd136314880;
      13505: inst = 32'd268468224;
      13506: inst = 32'd201345645;
      13507: inst = 32'd203480827;
      13508: inst = 32'd471859200;
      13509: inst = 32'd136314880;
      13510: inst = 32'd268468224;
      13511: inst = 32'd201345646;
      13512: inst = 32'd203480827;
      13513: inst = 32'd471859200;
      13514: inst = 32'd136314880;
      13515: inst = 32'd268468224;
      13516: inst = 32'd201345647;
      13517: inst = 32'd203484888;
      13518: inst = 32'd471859200;
      13519: inst = 32'd136314880;
      13520: inst = 32'd268468224;
      13521: inst = 32'd201345648;
      13522: inst = 32'd203484854;
      13523: inst = 32'd471859200;
      13524: inst = 32'd136314880;
      13525: inst = 32'd268468224;
      13526: inst = 32'd201345649;
      13527: inst = 32'd203484854;
      13528: inst = 32'd471859200;
      13529: inst = 32'd136314880;
      13530: inst = 32'd268468224;
      13531: inst = 32'd201345650;
      13532: inst = 32'd203484854;
      13533: inst = 32'd471859200;
      13534: inst = 32'd136314880;
      13535: inst = 32'd268468224;
      13536: inst = 32'd201345651;
      13537: inst = 32'd203484854;
      13538: inst = 32'd471859200;
      13539: inst = 32'd136314880;
      13540: inst = 32'd268468224;
      13541: inst = 32'd201345652;
      13542: inst = 32'd203484854;
      13543: inst = 32'd471859200;
      13544: inst = 32'd136314880;
      13545: inst = 32'd268468224;
      13546: inst = 32'd201345653;
      13547: inst = 32'd203484854;
      13548: inst = 32'd471859200;
      13549: inst = 32'd136314880;
      13550: inst = 32'd268468224;
      13551: inst = 32'd201345654;
      13552: inst = 32'd203484854;
      13553: inst = 32'd471859200;
      13554: inst = 32'd136314880;
      13555: inst = 32'd268468224;
      13556: inst = 32'd201345655;
      13557: inst = 32'd203484854;
      13558: inst = 32'd471859200;
      13559: inst = 32'd136314880;
      13560: inst = 32'd268468224;
      13561: inst = 32'd201345656;
      13562: inst = 32'd203484854;
      13563: inst = 32'd471859200;
      13564: inst = 32'd136314880;
      13565: inst = 32'd268468224;
      13566: inst = 32'd201345657;
      13567: inst = 32'd203484854;
      13568: inst = 32'd471859200;
      13569: inst = 32'd136314880;
      13570: inst = 32'd268468224;
      13571: inst = 32'd201345658;
      13572: inst = 32'd203484854;
      13573: inst = 32'd471859200;
      13574: inst = 32'd136314880;
      13575: inst = 32'd268468224;
      13576: inst = 32'd201345659;
      13577: inst = 32'd203484854;
      13578: inst = 32'd471859200;
      13579: inst = 32'd136314880;
      13580: inst = 32'd268468224;
      13581: inst = 32'd201345660;
      13582: inst = 32'd203489279;
      13583: inst = 32'd471859200;
      13584: inst = 32'd136314880;
      13585: inst = 32'd268468224;
      13586: inst = 32'd201345661;
      13587: inst = 32'd203489279;
      13588: inst = 32'd471859200;
      13589: inst = 32'd136314880;
      13590: inst = 32'd268468224;
      13591: inst = 32'd201345662;
      13592: inst = 32'd203489279;
      13593: inst = 32'd471859200;
      13594: inst = 32'd136314880;
      13595: inst = 32'd268468224;
      13596: inst = 32'd201345663;
      13597: inst = 32'd203489279;
      13598: inst = 32'd471859200;
      13599: inst = 32'd136314880;
      13600: inst = 32'd268468224;
      13601: inst = 32'd201345664;
      13602: inst = 32'd203489279;
      13603: inst = 32'd471859200;
      13604: inst = 32'd136314880;
      13605: inst = 32'd268468224;
      13606: inst = 32'd201345665;
      13607: inst = 32'd203489279;
      13608: inst = 32'd471859200;
      13609: inst = 32'd136314880;
      13610: inst = 32'd268468224;
      13611: inst = 32'd201345666;
      13612: inst = 32'd203489279;
      13613: inst = 32'd471859200;
      13614: inst = 32'd136314880;
      13615: inst = 32'd268468224;
      13616: inst = 32'd201345667;
      13617: inst = 32'd203489279;
      13618: inst = 32'd471859200;
      13619: inst = 32'd136314880;
      13620: inst = 32'd268468224;
      13621: inst = 32'd201345668;
      13622: inst = 32'd203489279;
      13623: inst = 32'd471859200;
      13624: inst = 32'd136314880;
      13625: inst = 32'd268468224;
      13626: inst = 32'd201345669;
      13627: inst = 32'd203489279;
      13628: inst = 32'd471859200;
      13629: inst = 32'd136314880;
      13630: inst = 32'd268468224;
      13631: inst = 32'd201345670;
      13632: inst = 32'd203489279;
      13633: inst = 32'd471859200;
      13634: inst = 32'd136314880;
      13635: inst = 32'd268468224;
      13636: inst = 32'd201345671;
      13637: inst = 32'd203489279;
      13638: inst = 32'd471859200;
      13639: inst = 32'd136314880;
      13640: inst = 32'd268468224;
      13641: inst = 32'd201345672;
      13642: inst = 32'd203489279;
      13643: inst = 32'd471859200;
      13644: inst = 32'd136314880;
      13645: inst = 32'd268468224;
      13646: inst = 32'd201345673;
      13647: inst = 32'd203489279;
      13648: inst = 32'd471859200;
      13649: inst = 32'd136314880;
      13650: inst = 32'd268468224;
      13651: inst = 32'd201345674;
      13652: inst = 32'd203489279;
      13653: inst = 32'd471859200;
      13654: inst = 32'd136314880;
      13655: inst = 32'd268468224;
      13656: inst = 32'd201345675;
      13657: inst = 32'd203489279;
      13658: inst = 32'd471859200;
      13659: inst = 32'd136314880;
      13660: inst = 32'd268468224;
      13661: inst = 32'd201345676;
      13662: inst = 32'd203489279;
      13663: inst = 32'd471859200;
      13664: inst = 32'd136314880;
      13665: inst = 32'd268468224;
      13666: inst = 32'd201345677;
      13667: inst = 32'd203489279;
      13668: inst = 32'd471859200;
      13669: inst = 32'd136314880;
      13670: inst = 32'd268468224;
      13671: inst = 32'd201345678;
      13672: inst = 32'd203489279;
      13673: inst = 32'd471859200;
      13674: inst = 32'd136314880;
      13675: inst = 32'd268468224;
      13676: inst = 32'd201345679;
      13677: inst = 32'd203489279;
      13678: inst = 32'd471859200;
      13679: inst = 32'd136314880;
      13680: inst = 32'd268468224;
      13681: inst = 32'd201345680;
      13682: inst = 32'd203489279;
      13683: inst = 32'd471859200;
      13684: inst = 32'd136314880;
      13685: inst = 32'd268468224;
      13686: inst = 32'd201345681;
      13687: inst = 32'd203489279;
      13688: inst = 32'd471859200;
      13689: inst = 32'd136314880;
      13690: inst = 32'd268468224;
      13691: inst = 32'd201345682;
      13692: inst = 32'd203489279;
      13693: inst = 32'd471859200;
      13694: inst = 32'd136314880;
      13695: inst = 32'd268468224;
      13696: inst = 32'd201345683;
      13697: inst = 32'd203489279;
      13698: inst = 32'd471859200;
      13699: inst = 32'd136314880;
      13700: inst = 32'd268468224;
      13701: inst = 32'd201345684;
      13702: inst = 32'd203489279;
      13703: inst = 32'd471859200;
      13704: inst = 32'd136314880;
      13705: inst = 32'd268468224;
      13706: inst = 32'd201345685;
      13707: inst = 32'd203489279;
      13708: inst = 32'd471859200;
      13709: inst = 32'd136314880;
      13710: inst = 32'd268468224;
      13711: inst = 32'd201345686;
      13712: inst = 32'd203489279;
      13713: inst = 32'd471859200;
      13714: inst = 32'd136314880;
      13715: inst = 32'd268468224;
      13716: inst = 32'd201345687;
      13717: inst = 32'd203489279;
      13718: inst = 32'd471859200;
      13719: inst = 32'd136314880;
      13720: inst = 32'd268468224;
      13721: inst = 32'd201345688;
      13722: inst = 32'd203489279;
      13723: inst = 32'd471859200;
      13724: inst = 32'd136314880;
      13725: inst = 32'd268468224;
      13726: inst = 32'd201345689;
      13727: inst = 32'd203489279;
      13728: inst = 32'd471859200;
      13729: inst = 32'd136314880;
      13730: inst = 32'd268468224;
      13731: inst = 32'd201345690;
      13732: inst = 32'd203489279;
      13733: inst = 32'd471859200;
      13734: inst = 32'd136314880;
      13735: inst = 32'd268468224;
      13736: inst = 32'd201345691;
      13737: inst = 32'd203489279;
      13738: inst = 32'd471859200;
      13739: inst = 32'd136314880;
      13740: inst = 32'd268468224;
      13741: inst = 32'd201345692;
      13742: inst = 32'd203489279;
      13743: inst = 32'd471859200;
      13744: inst = 32'd136314880;
      13745: inst = 32'd268468224;
      13746: inst = 32'd201345693;
      13747: inst = 32'd203489279;
      13748: inst = 32'd471859200;
      13749: inst = 32'd136314880;
      13750: inst = 32'd268468224;
      13751: inst = 32'd201345694;
      13752: inst = 32'd203489279;
      13753: inst = 32'd471859200;
      13754: inst = 32'd136314880;
      13755: inst = 32'd268468224;
      13756: inst = 32'd201345695;
      13757: inst = 32'd203489279;
      13758: inst = 32'd471859200;
      13759: inst = 32'd136314880;
      13760: inst = 32'd268468224;
      13761: inst = 32'd201345696;
      13762: inst = 32'd203489279;
      13763: inst = 32'd471859200;
      13764: inst = 32'd136314880;
      13765: inst = 32'd268468224;
      13766: inst = 32'd201345697;
      13767: inst = 32'd203489279;
      13768: inst = 32'd471859200;
      13769: inst = 32'd136314880;
      13770: inst = 32'd268468224;
      13771: inst = 32'd201345698;
      13772: inst = 32'd203489279;
      13773: inst = 32'd471859200;
      13774: inst = 32'd136314880;
      13775: inst = 32'd268468224;
      13776: inst = 32'd201345699;
      13777: inst = 32'd203489279;
      13778: inst = 32'd471859200;
      13779: inst = 32'd136314880;
      13780: inst = 32'd268468224;
      13781: inst = 32'd201345700;
      13782: inst = 32'd203484854;
      13783: inst = 32'd471859200;
      13784: inst = 32'd136314880;
      13785: inst = 32'd268468224;
      13786: inst = 32'd201345701;
      13787: inst = 32'd203484854;
      13788: inst = 32'd471859200;
      13789: inst = 32'd136314880;
      13790: inst = 32'd268468224;
      13791: inst = 32'd201345702;
      13792: inst = 32'd203484854;
      13793: inst = 32'd471859200;
      13794: inst = 32'd136314880;
      13795: inst = 32'd268468224;
      13796: inst = 32'd201345703;
      13797: inst = 32'd203484854;
      13798: inst = 32'd471859200;
      13799: inst = 32'd136314880;
      13800: inst = 32'd268468224;
      13801: inst = 32'd201345704;
      13802: inst = 32'd203484854;
      13803: inst = 32'd471859200;
      13804: inst = 32'd136314880;
      13805: inst = 32'd268468224;
      13806: inst = 32'd201345705;
      13807: inst = 32'd203484854;
      13808: inst = 32'd471859200;
      13809: inst = 32'd136314880;
      13810: inst = 32'd268468224;
      13811: inst = 32'd201345706;
      13812: inst = 32'd203484854;
      13813: inst = 32'd471859200;
      13814: inst = 32'd136314880;
      13815: inst = 32'd268468224;
      13816: inst = 32'd201345707;
      13817: inst = 32'd203484854;
      13818: inst = 32'd471859200;
      13819: inst = 32'd136314880;
      13820: inst = 32'd268468224;
      13821: inst = 32'd201345708;
      13822: inst = 32'd203484854;
      13823: inst = 32'd471859200;
      13824: inst = 32'd136314880;
      13825: inst = 32'd268468224;
      13826: inst = 32'd201345709;
      13827: inst = 32'd203484854;
      13828: inst = 32'd471859200;
      13829: inst = 32'd136314880;
      13830: inst = 32'd268468224;
      13831: inst = 32'd201345710;
      13832: inst = 32'd203484854;
      13833: inst = 32'd471859200;
      13834: inst = 32'd136314880;
      13835: inst = 32'd268468224;
      13836: inst = 32'd201345711;
      13837: inst = 32'd203473634;
      13838: inst = 32'd471859200;
      13839: inst = 32'd136314880;
      13840: inst = 32'd268468224;
      13841: inst = 32'd201345712;
      13842: inst = 32'd203480005;
      13843: inst = 32'd471859200;
      13844: inst = 32'd136314880;
      13845: inst = 32'd268468224;
      13846: inst = 32'd201345713;
      13847: inst = 32'd203480005;
      13848: inst = 32'd471859200;
      13849: inst = 32'd136314880;
      13850: inst = 32'd268468224;
      13851: inst = 32'd201345714;
      13852: inst = 32'd203485052;
      13853: inst = 32'd471859200;
      13854: inst = 32'd136314880;
      13855: inst = 32'd268468224;
      13856: inst = 32'd201345715;
      13857: inst = 32'd203485052;
      13858: inst = 32'd471859200;
      13859: inst = 32'd136314880;
      13860: inst = 32'd268468224;
      13861: inst = 32'd201345716;
      13862: inst = 32'd203489279;
      13863: inst = 32'd471859200;
      13864: inst = 32'd136314880;
      13865: inst = 32'd268468224;
      13866: inst = 32'd201345717;
      13867: inst = 32'd203485052;
      13868: inst = 32'd471859200;
      13869: inst = 32'd136314880;
      13870: inst = 32'd268468224;
      13871: inst = 32'd201345718;
      13872: inst = 32'd203480005;
      13873: inst = 32'd471859200;
      13874: inst = 32'd136314880;
      13875: inst = 32'd268468224;
      13876: inst = 32'd201345719;
      13877: inst = 32'd203480005;
      13878: inst = 32'd471859200;
      13879: inst = 32'd136314880;
      13880: inst = 32'd268468224;
      13881: inst = 32'd201345720;
      13882: inst = 32'd203480005;
      13883: inst = 32'd471859200;
      13884: inst = 32'd136314880;
      13885: inst = 32'd268468224;
      13886: inst = 32'd201345721;
      13887: inst = 32'd203480005;
      13888: inst = 32'd471859200;
      13889: inst = 32'd136314880;
      13890: inst = 32'd268468224;
      13891: inst = 32'd201345722;
      13892: inst = 32'd203480005;
      13893: inst = 32'd471859200;
      13894: inst = 32'd136314880;
      13895: inst = 32'd268468224;
      13896: inst = 32'd201345723;
      13897: inst = 32'd203480005;
      13898: inst = 32'd471859200;
      13899: inst = 32'd136314880;
      13900: inst = 32'd268468224;
      13901: inst = 32'd201345724;
      13902: inst = 32'd203480005;
      13903: inst = 32'd471859200;
      13904: inst = 32'd136314880;
      13905: inst = 32'd268468224;
      13906: inst = 32'd201345725;
      13907: inst = 32'd203480005;
      13908: inst = 32'd471859200;
      13909: inst = 32'd136314880;
      13910: inst = 32'd268468224;
      13911: inst = 32'd201345726;
      13912: inst = 32'd203480005;
      13913: inst = 32'd471859200;
      13914: inst = 32'd136314880;
      13915: inst = 32'd268468224;
      13916: inst = 32'd201345727;
      13917: inst = 32'd203473634;
      13918: inst = 32'd471859200;
      13919: inst = 32'd136314880;
      13920: inst = 32'd268468224;
      13921: inst = 32'd201345728;
      13922: inst = 32'd203484854;
      13923: inst = 32'd471859200;
      13924: inst = 32'd136314880;
      13925: inst = 32'd268468224;
      13926: inst = 32'd201345729;
      13927: inst = 32'd203484854;
      13928: inst = 32'd471859200;
      13929: inst = 32'd136314880;
      13930: inst = 32'd268468224;
      13931: inst = 32'd201345730;
      13932: inst = 32'd203484854;
      13933: inst = 32'd471859200;
      13934: inst = 32'd136314880;
      13935: inst = 32'd268468224;
      13936: inst = 32'd201345731;
      13937: inst = 32'd203484854;
      13938: inst = 32'd471859200;
      13939: inst = 32'd136314880;
      13940: inst = 32'd268468224;
      13941: inst = 32'd201345732;
      13942: inst = 32'd203484854;
      13943: inst = 32'd471859200;
      13944: inst = 32'd136314880;
      13945: inst = 32'd268468224;
      13946: inst = 32'd201345733;
      13947: inst = 32'd203484854;
      13948: inst = 32'd471859200;
      13949: inst = 32'd136314880;
      13950: inst = 32'd268468224;
      13951: inst = 32'd201345734;
      13952: inst = 32'd203484854;
      13953: inst = 32'd471859200;
      13954: inst = 32'd136314880;
      13955: inst = 32'd268468224;
      13956: inst = 32'd201345735;
      13957: inst = 32'd203482875;
      13958: inst = 32'd471859200;
      13959: inst = 32'd136314880;
      13960: inst = 32'd268468224;
      13961: inst = 32'd201345736;
      13962: inst = 32'd203480827;
      13963: inst = 32'd471859200;
      13964: inst = 32'd136314880;
      13965: inst = 32'd268468224;
      13966: inst = 32'd201345737;
      13967: inst = 32'd203480827;
      13968: inst = 32'd471859200;
      13969: inst = 32'd136314880;
      13970: inst = 32'd268468224;
      13971: inst = 32'd201345738;
      13972: inst = 32'd203480827;
      13973: inst = 32'd471859200;
      13974: inst = 32'd136314880;
      13975: inst = 32'd268468224;
      13976: inst = 32'd201345739;
      13977: inst = 32'd203480827;
      13978: inst = 32'd471859200;
      13979: inst = 32'd136314880;
      13980: inst = 32'd268468224;
      13981: inst = 32'd201345740;
      13982: inst = 32'd203480827;
      13983: inst = 32'd471859200;
      13984: inst = 32'd136314880;
      13985: inst = 32'd268468224;
      13986: inst = 32'd201345741;
      13987: inst = 32'd203480827;
      13988: inst = 32'd471859200;
      13989: inst = 32'd136314880;
      13990: inst = 32'd268468224;
      13991: inst = 32'd201345742;
      13992: inst = 32'd203480827;
      13993: inst = 32'd471859200;
      13994: inst = 32'd136314880;
      13995: inst = 32'd268468224;
      13996: inst = 32'd201345743;
      13997: inst = 32'd203482875;
      13998: inst = 32'd471859200;
      13999: inst = 32'd136314880;
      14000: inst = 32'd268468224;
      14001: inst = 32'd201345744;
      14002: inst = 32'd203484854;
      14003: inst = 32'd471859200;
      14004: inst = 32'd136314880;
      14005: inst = 32'd268468224;
      14006: inst = 32'd201345745;
      14007: inst = 32'd203484854;
      14008: inst = 32'd471859200;
      14009: inst = 32'd136314880;
      14010: inst = 32'd268468224;
      14011: inst = 32'd201345746;
      14012: inst = 32'd203484854;
      14013: inst = 32'd471859200;
      14014: inst = 32'd136314880;
      14015: inst = 32'd268468224;
      14016: inst = 32'd201345747;
      14017: inst = 32'd203484854;
      14018: inst = 32'd471859200;
      14019: inst = 32'd136314880;
      14020: inst = 32'd268468224;
      14021: inst = 32'd201345748;
      14022: inst = 32'd203484854;
      14023: inst = 32'd471859200;
      14024: inst = 32'd136314880;
      14025: inst = 32'd268468224;
      14026: inst = 32'd201345749;
      14027: inst = 32'd203484854;
      14028: inst = 32'd471859200;
      14029: inst = 32'd136314880;
      14030: inst = 32'd268468224;
      14031: inst = 32'd201345750;
      14032: inst = 32'd203484854;
      14033: inst = 32'd471859200;
      14034: inst = 32'd136314880;
      14035: inst = 32'd268468224;
      14036: inst = 32'd201345751;
      14037: inst = 32'd203484854;
      14038: inst = 32'd471859200;
      14039: inst = 32'd136314880;
      14040: inst = 32'd268468224;
      14041: inst = 32'd201345752;
      14042: inst = 32'd203484854;
      14043: inst = 32'd471859200;
      14044: inst = 32'd136314880;
      14045: inst = 32'd268468224;
      14046: inst = 32'd201345753;
      14047: inst = 32'd203484854;
      14048: inst = 32'd471859200;
      14049: inst = 32'd136314880;
      14050: inst = 32'd268468224;
      14051: inst = 32'd201345754;
      14052: inst = 32'd203484854;
      14053: inst = 32'd471859200;
      14054: inst = 32'd136314880;
      14055: inst = 32'd268468224;
      14056: inst = 32'd201345755;
      14057: inst = 32'd203484854;
      14058: inst = 32'd471859200;
      14059: inst = 32'd136314880;
      14060: inst = 32'd268468224;
      14061: inst = 32'd201345756;
      14062: inst = 32'd203489279;
      14063: inst = 32'd471859200;
      14064: inst = 32'd136314880;
      14065: inst = 32'd268468224;
      14066: inst = 32'd201345757;
      14067: inst = 32'd203489279;
      14068: inst = 32'd471859200;
      14069: inst = 32'd136314880;
      14070: inst = 32'd268468224;
      14071: inst = 32'd201345758;
      14072: inst = 32'd203489279;
      14073: inst = 32'd471859200;
      14074: inst = 32'd136314880;
      14075: inst = 32'd268468224;
      14076: inst = 32'd201345759;
      14077: inst = 32'd203489279;
      14078: inst = 32'd471859200;
      14079: inst = 32'd136314880;
      14080: inst = 32'd268468224;
      14081: inst = 32'd201345760;
      14082: inst = 32'd203489279;
      14083: inst = 32'd471859200;
      14084: inst = 32'd136314880;
      14085: inst = 32'd268468224;
      14086: inst = 32'd201345761;
      14087: inst = 32'd203489279;
      14088: inst = 32'd471859200;
      14089: inst = 32'd136314880;
      14090: inst = 32'd268468224;
      14091: inst = 32'd201345762;
      14092: inst = 32'd203489279;
      14093: inst = 32'd471859200;
      14094: inst = 32'd136314880;
      14095: inst = 32'd268468224;
      14096: inst = 32'd201345763;
      14097: inst = 32'd203489279;
      14098: inst = 32'd471859200;
      14099: inst = 32'd136314880;
      14100: inst = 32'd268468224;
      14101: inst = 32'd201345764;
      14102: inst = 32'd203489279;
      14103: inst = 32'd471859200;
      14104: inst = 32'd136314880;
      14105: inst = 32'd268468224;
      14106: inst = 32'd201345765;
      14107: inst = 32'd203489279;
      14108: inst = 32'd471859200;
      14109: inst = 32'd136314880;
      14110: inst = 32'd268468224;
      14111: inst = 32'd201345766;
      14112: inst = 32'd203489279;
      14113: inst = 32'd471859200;
      14114: inst = 32'd136314880;
      14115: inst = 32'd268468224;
      14116: inst = 32'd201345767;
      14117: inst = 32'd203489279;
      14118: inst = 32'd471859200;
      14119: inst = 32'd136314880;
      14120: inst = 32'd268468224;
      14121: inst = 32'd201345768;
      14122: inst = 32'd203489279;
      14123: inst = 32'd471859200;
      14124: inst = 32'd136314880;
      14125: inst = 32'd268468224;
      14126: inst = 32'd201345769;
      14127: inst = 32'd203489279;
      14128: inst = 32'd471859200;
      14129: inst = 32'd136314880;
      14130: inst = 32'd268468224;
      14131: inst = 32'd201345770;
      14132: inst = 32'd203489279;
      14133: inst = 32'd471859200;
      14134: inst = 32'd136314880;
      14135: inst = 32'd268468224;
      14136: inst = 32'd201345771;
      14137: inst = 32'd203489279;
      14138: inst = 32'd471859200;
      14139: inst = 32'd136314880;
      14140: inst = 32'd268468224;
      14141: inst = 32'd201345772;
      14142: inst = 32'd203489279;
      14143: inst = 32'd471859200;
      14144: inst = 32'd136314880;
      14145: inst = 32'd268468224;
      14146: inst = 32'd201345773;
      14147: inst = 32'd203489279;
      14148: inst = 32'd471859200;
      14149: inst = 32'd136314880;
      14150: inst = 32'd268468224;
      14151: inst = 32'd201345774;
      14152: inst = 32'd203489279;
      14153: inst = 32'd471859200;
      14154: inst = 32'd136314880;
      14155: inst = 32'd268468224;
      14156: inst = 32'd201345775;
      14157: inst = 32'd203489279;
      14158: inst = 32'd471859200;
      14159: inst = 32'd136314880;
      14160: inst = 32'd268468224;
      14161: inst = 32'd201345776;
      14162: inst = 32'd203489279;
      14163: inst = 32'd471859200;
      14164: inst = 32'd136314880;
      14165: inst = 32'd268468224;
      14166: inst = 32'd201345777;
      14167: inst = 32'd203489279;
      14168: inst = 32'd471859200;
      14169: inst = 32'd136314880;
      14170: inst = 32'd268468224;
      14171: inst = 32'd201345778;
      14172: inst = 32'd203489279;
      14173: inst = 32'd471859200;
      14174: inst = 32'd136314880;
      14175: inst = 32'd268468224;
      14176: inst = 32'd201345779;
      14177: inst = 32'd203489279;
      14178: inst = 32'd471859200;
      14179: inst = 32'd136314880;
      14180: inst = 32'd268468224;
      14181: inst = 32'd201345780;
      14182: inst = 32'd203489279;
      14183: inst = 32'd471859200;
      14184: inst = 32'd136314880;
      14185: inst = 32'd268468224;
      14186: inst = 32'd201345781;
      14187: inst = 32'd203489279;
      14188: inst = 32'd471859200;
      14189: inst = 32'd136314880;
      14190: inst = 32'd268468224;
      14191: inst = 32'd201345782;
      14192: inst = 32'd203489279;
      14193: inst = 32'd471859200;
      14194: inst = 32'd136314880;
      14195: inst = 32'd268468224;
      14196: inst = 32'd201345783;
      14197: inst = 32'd203489279;
      14198: inst = 32'd471859200;
      14199: inst = 32'd136314880;
      14200: inst = 32'd268468224;
      14201: inst = 32'd201345784;
      14202: inst = 32'd203489279;
      14203: inst = 32'd471859200;
      14204: inst = 32'd136314880;
      14205: inst = 32'd268468224;
      14206: inst = 32'd201345785;
      14207: inst = 32'd203489279;
      14208: inst = 32'd471859200;
      14209: inst = 32'd136314880;
      14210: inst = 32'd268468224;
      14211: inst = 32'd201345786;
      14212: inst = 32'd203489279;
      14213: inst = 32'd471859200;
      14214: inst = 32'd136314880;
      14215: inst = 32'd268468224;
      14216: inst = 32'd201345787;
      14217: inst = 32'd203489279;
      14218: inst = 32'd471859200;
      14219: inst = 32'd136314880;
      14220: inst = 32'd268468224;
      14221: inst = 32'd201345788;
      14222: inst = 32'd203489279;
      14223: inst = 32'd471859200;
      14224: inst = 32'd136314880;
      14225: inst = 32'd268468224;
      14226: inst = 32'd201345789;
      14227: inst = 32'd203489279;
      14228: inst = 32'd471859200;
      14229: inst = 32'd136314880;
      14230: inst = 32'd268468224;
      14231: inst = 32'd201345790;
      14232: inst = 32'd203489279;
      14233: inst = 32'd471859200;
      14234: inst = 32'd136314880;
      14235: inst = 32'd268468224;
      14236: inst = 32'd201345791;
      14237: inst = 32'd203489279;
      14238: inst = 32'd471859200;
      14239: inst = 32'd136314880;
      14240: inst = 32'd268468224;
      14241: inst = 32'd201345792;
      14242: inst = 32'd203489279;
      14243: inst = 32'd471859200;
      14244: inst = 32'd136314880;
      14245: inst = 32'd268468224;
      14246: inst = 32'd201345793;
      14247: inst = 32'd203489279;
      14248: inst = 32'd471859200;
      14249: inst = 32'd136314880;
      14250: inst = 32'd268468224;
      14251: inst = 32'd201345794;
      14252: inst = 32'd203489279;
      14253: inst = 32'd471859200;
      14254: inst = 32'd136314880;
      14255: inst = 32'd268468224;
      14256: inst = 32'd201345795;
      14257: inst = 32'd203489279;
      14258: inst = 32'd471859200;
      14259: inst = 32'd136314880;
      14260: inst = 32'd268468224;
      14261: inst = 32'd201345796;
      14262: inst = 32'd203484854;
      14263: inst = 32'd471859200;
      14264: inst = 32'd136314880;
      14265: inst = 32'd268468224;
      14266: inst = 32'd201345797;
      14267: inst = 32'd203484854;
      14268: inst = 32'd471859200;
      14269: inst = 32'd136314880;
      14270: inst = 32'd268468224;
      14271: inst = 32'd201345798;
      14272: inst = 32'd203484854;
      14273: inst = 32'd471859200;
      14274: inst = 32'd136314880;
      14275: inst = 32'd268468224;
      14276: inst = 32'd201345799;
      14277: inst = 32'd203484854;
      14278: inst = 32'd471859200;
      14279: inst = 32'd136314880;
      14280: inst = 32'd268468224;
      14281: inst = 32'd201345800;
      14282: inst = 32'd203484854;
      14283: inst = 32'd471859200;
      14284: inst = 32'd136314880;
      14285: inst = 32'd268468224;
      14286: inst = 32'd201345801;
      14287: inst = 32'd203484854;
      14288: inst = 32'd471859200;
      14289: inst = 32'd136314880;
      14290: inst = 32'd268468224;
      14291: inst = 32'd201345802;
      14292: inst = 32'd203484854;
      14293: inst = 32'd471859200;
      14294: inst = 32'd136314880;
      14295: inst = 32'd268468224;
      14296: inst = 32'd201345803;
      14297: inst = 32'd203484854;
      14298: inst = 32'd471859200;
      14299: inst = 32'd136314880;
      14300: inst = 32'd268468224;
      14301: inst = 32'd201345804;
      14302: inst = 32'd203484854;
      14303: inst = 32'd471859200;
      14304: inst = 32'd136314880;
      14305: inst = 32'd268468224;
      14306: inst = 32'd201345805;
      14307: inst = 32'd203484854;
      14308: inst = 32'd471859200;
      14309: inst = 32'd136314880;
      14310: inst = 32'd268468224;
      14311: inst = 32'd201345806;
      14312: inst = 32'd203484854;
      14313: inst = 32'd471859200;
      14314: inst = 32'd136314880;
      14315: inst = 32'd268468224;
      14316: inst = 32'd201345807;
      14317: inst = 32'd203473634;
      14318: inst = 32'd471859200;
      14319: inst = 32'd136314880;
      14320: inst = 32'd268468224;
      14321: inst = 32'd201345808;
      14322: inst = 32'd203480005;
      14323: inst = 32'd471859200;
      14324: inst = 32'd136314880;
      14325: inst = 32'd268468224;
      14326: inst = 32'd201345809;
      14327: inst = 32'd203480005;
      14328: inst = 32'd471859200;
      14329: inst = 32'd136314880;
      14330: inst = 32'd268468224;
      14331: inst = 32'd201345810;
      14332: inst = 32'd203485052;
      14333: inst = 32'd471859200;
      14334: inst = 32'd136314880;
      14335: inst = 32'd268468224;
      14336: inst = 32'd201345811;
      14337: inst = 32'd203485052;
      14338: inst = 32'd471859200;
      14339: inst = 32'd136314880;
      14340: inst = 32'd268468224;
      14341: inst = 32'd201345812;
      14342: inst = 32'd203489279;
      14343: inst = 32'd471859200;
      14344: inst = 32'd136314880;
      14345: inst = 32'd268468224;
      14346: inst = 32'd201345813;
      14347: inst = 32'd203485052;
      14348: inst = 32'd471859200;
      14349: inst = 32'd136314880;
      14350: inst = 32'd268468224;
      14351: inst = 32'd201345814;
      14352: inst = 32'd203480005;
      14353: inst = 32'd471859200;
      14354: inst = 32'd136314880;
      14355: inst = 32'd268468224;
      14356: inst = 32'd201345815;
      14357: inst = 32'd203480005;
      14358: inst = 32'd471859200;
      14359: inst = 32'd136314880;
      14360: inst = 32'd268468224;
      14361: inst = 32'd201345816;
      14362: inst = 32'd203480005;
      14363: inst = 32'd471859200;
      14364: inst = 32'd136314880;
      14365: inst = 32'd268468224;
      14366: inst = 32'd201345817;
      14367: inst = 32'd203480005;
      14368: inst = 32'd471859200;
      14369: inst = 32'd136314880;
      14370: inst = 32'd268468224;
      14371: inst = 32'd201345818;
      14372: inst = 32'd203480005;
      14373: inst = 32'd471859200;
      14374: inst = 32'd136314880;
      14375: inst = 32'd268468224;
      14376: inst = 32'd201345819;
      14377: inst = 32'd203480005;
      14378: inst = 32'd471859200;
      14379: inst = 32'd136314880;
      14380: inst = 32'd268468224;
      14381: inst = 32'd201345820;
      14382: inst = 32'd203480005;
      14383: inst = 32'd471859200;
      14384: inst = 32'd136314880;
      14385: inst = 32'd268468224;
      14386: inst = 32'd201345821;
      14387: inst = 32'd203480005;
      14388: inst = 32'd471859200;
      14389: inst = 32'd136314880;
      14390: inst = 32'd268468224;
      14391: inst = 32'd201345822;
      14392: inst = 32'd203480005;
      14393: inst = 32'd471859200;
      14394: inst = 32'd136314880;
      14395: inst = 32'd268468224;
      14396: inst = 32'd201345823;
      14397: inst = 32'd203473634;
      14398: inst = 32'd471859200;
      14399: inst = 32'd136314880;
      14400: inst = 32'd268468224;
      14401: inst = 32'd201345824;
      14402: inst = 32'd203484854;
      14403: inst = 32'd471859200;
      14404: inst = 32'd136314880;
      14405: inst = 32'd268468224;
      14406: inst = 32'd201345825;
      14407: inst = 32'd203484854;
      14408: inst = 32'd471859200;
      14409: inst = 32'd136314880;
      14410: inst = 32'd268468224;
      14411: inst = 32'd201345826;
      14412: inst = 32'd203484854;
      14413: inst = 32'd471859200;
      14414: inst = 32'd136314880;
      14415: inst = 32'd268468224;
      14416: inst = 32'd201345827;
      14417: inst = 32'd203484854;
      14418: inst = 32'd471859200;
      14419: inst = 32'd136314880;
      14420: inst = 32'd268468224;
      14421: inst = 32'd201345828;
      14422: inst = 32'd203484854;
      14423: inst = 32'd471859200;
      14424: inst = 32'd136314880;
      14425: inst = 32'd268468224;
      14426: inst = 32'd201345829;
      14427: inst = 32'd203484854;
      14428: inst = 32'd471859200;
      14429: inst = 32'd136314880;
      14430: inst = 32'd268468224;
      14431: inst = 32'd201345830;
      14432: inst = 32'd203484854;
      14433: inst = 32'd471859200;
      14434: inst = 32'd136314880;
      14435: inst = 32'd268468224;
      14436: inst = 32'd201345831;
      14437: inst = 32'd203480827;
      14438: inst = 32'd471859200;
      14439: inst = 32'd136314880;
      14440: inst = 32'd268468224;
      14441: inst = 32'd201345832;
      14442: inst = 32'd203442793;
      14443: inst = 32'd471859200;
      14444: inst = 32'd136314880;
      14445: inst = 32'd268468224;
      14446: inst = 32'd201345833;
      14447: inst = 32'd203442793;
      14448: inst = 32'd471859200;
      14449: inst = 32'd136314880;
      14450: inst = 32'd268468224;
      14451: inst = 32'd201345834;
      14452: inst = 32'd203480827;
      14453: inst = 32'd471859200;
      14454: inst = 32'd136314880;
      14455: inst = 32'd268468224;
      14456: inst = 32'd201345835;
      14457: inst = 32'd203442793;
      14458: inst = 32'd471859200;
      14459: inst = 32'd136314880;
      14460: inst = 32'd268468224;
      14461: inst = 32'd201345836;
      14462: inst = 32'd203442793;
      14463: inst = 32'd471859200;
      14464: inst = 32'd136314880;
      14465: inst = 32'd268468224;
      14466: inst = 32'd201345837;
      14467: inst = 32'd203480827;
      14468: inst = 32'd471859200;
      14469: inst = 32'd136314880;
      14470: inst = 32'd268468224;
      14471: inst = 32'd201345838;
      14472: inst = 32'd203480827;
      14473: inst = 32'd471859200;
      14474: inst = 32'd136314880;
      14475: inst = 32'd268468224;
      14476: inst = 32'd201345839;
      14477: inst = 32'd203480827;
      14478: inst = 32'd471859200;
      14479: inst = 32'd136314880;
      14480: inst = 32'd268468224;
      14481: inst = 32'd201345840;
      14482: inst = 32'd203484854;
      14483: inst = 32'd471859200;
      14484: inst = 32'd136314880;
      14485: inst = 32'd268468224;
      14486: inst = 32'd201345841;
      14487: inst = 32'd203484854;
      14488: inst = 32'd471859200;
      14489: inst = 32'd136314880;
      14490: inst = 32'd268468224;
      14491: inst = 32'd201345842;
      14492: inst = 32'd203484854;
      14493: inst = 32'd471859200;
      14494: inst = 32'd136314880;
      14495: inst = 32'd268468224;
      14496: inst = 32'd201345843;
      14497: inst = 32'd203484854;
      14498: inst = 32'd471859200;
      14499: inst = 32'd136314880;
      14500: inst = 32'd268468224;
      14501: inst = 32'd201345844;
      14502: inst = 32'd203484854;
      14503: inst = 32'd471859200;
      14504: inst = 32'd136314880;
      14505: inst = 32'd268468224;
      14506: inst = 32'd201345845;
      14507: inst = 32'd203484854;
      14508: inst = 32'd471859200;
      14509: inst = 32'd136314880;
      14510: inst = 32'd268468224;
      14511: inst = 32'd201345846;
      14512: inst = 32'd203484854;
      14513: inst = 32'd471859200;
      14514: inst = 32'd136314880;
      14515: inst = 32'd268468224;
      14516: inst = 32'd201345847;
      14517: inst = 32'd203484854;
      14518: inst = 32'd471859200;
      14519: inst = 32'd136314880;
      14520: inst = 32'd268468224;
      14521: inst = 32'd201345848;
      14522: inst = 32'd203484854;
      14523: inst = 32'd471859200;
      14524: inst = 32'd136314880;
      14525: inst = 32'd268468224;
      14526: inst = 32'd201345849;
      14527: inst = 32'd203484854;
      14528: inst = 32'd471859200;
      14529: inst = 32'd136314880;
      14530: inst = 32'd268468224;
      14531: inst = 32'd201345850;
      14532: inst = 32'd203484854;
      14533: inst = 32'd471859200;
      14534: inst = 32'd136314880;
      14535: inst = 32'd268468224;
      14536: inst = 32'd201345851;
      14537: inst = 32'd203484854;
      14538: inst = 32'd471859200;
      14539: inst = 32'd136314880;
      14540: inst = 32'd268468224;
      14541: inst = 32'd201345852;
      14542: inst = 32'd203489279;
      14543: inst = 32'd471859200;
      14544: inst = 32'd136314880;
      14545: inst = 32'd268468224;
      14546: inst = 32'd201345853;
      14547: inst = 32'd203489279;
      14548: inst = 32'd471859200;
      14549: inst = 32'd136314880;
      14550: inst = 32'd268468224;
      14551: inst = 32'd201345854;
      14552: inst = 32'd203489279;
      14553: inst = 32'd471859200;
      14554: inst = 32'd136314880;
      14555: inst = 32'd268468224;
      14556: inst = 32'd201345855;
      14557: inst = 32'd203489279;
      14558: inst = 32'd471859200;
      14559: inst = 32'd136314880;
      14560: inst = 32'd268468224;
      14561: inst = 32'd201345856;
      14562: inst = 32'd203489279;
      14563: inst = 32'd471859200;
      14564: inst = 32'd136314880;
      14565: inst = 32'd268468224;
      14566: inst = 32'd201345857;
      14567: inst = 32'd203489279;
      14568: inst = 32'd471859200;
      14569: inst = 32'd136314880;
      14570: inst = 32'd268468224;
      14571: inst = 32'd201345858;
      14572: inst = 32'd203489279;
      14573: inst = 32'd471859200;
      14574: inst = 32'd136314880;
      14575: inst = 32'd268468224;
      14576: inst = 32'd201345859;
      14577: inst = 32'd203489279;
      14578: inst = 32'd471859200;
      14579: inst = 32'd136314880;
      14580: inst = 32'd268468224;
      14581: inst = 32'd201345860;
      14582: inst = 32'd203489279;
      14583: inst = 32'd471859200;
      14584: inst = 32'd136314880;
      14585: inst = 32'd268468224;
      14586: inst = 32'd201345861;
      14587: inst = 32'd203489279;
      14588: inst = 32'd471859200;
      14589: inst = 32'd136314880;
      14590: inst = 32'd268468224;
      14591: inst = 32'd201345862;
      14592: inst = 32'd203489279;
      14593: inst = 32'd471859200;
      14594: inst = 32'd136314880;
      14595: inst = 32'd268468224;
      14596: inst = 32'd201345863;
      14597: inst = 32'd203489279;
      14598: inst = 32'd471859200;
      14599: inst = 32'd136314880;
      14600: inst = 32'd268468224;
      14601: inst = 32'd201345864;
      14602: inst = 32'd203489279;
      14603: inst = 32'd471859200;
      14604: inst = 32'd136314880;
      14605: inst = 32'd268468224;
      14606: inst = 32'd201345865;
      14607: inst = 32'd203489279;
      14608: inst = 32'd471859200;
      14609: inst = 32'd136314880;
      14610: inst = 32'd268468224;
      14611: inst = 32'd201345866;
      14612: inst = 32'd203489279;
      14613: inst = 32'd471859200;
      14614: inst = 32'd136314880;
      14615: inst = 32'd268468224;
      14616: inst = 32'd201345867;
      14617: inst = 32'd203489279;
      14618: inst = 32'd471859200;
      14619: inst = 32'd136314880;
      14620: inst = 32'd268468224;
      14621: inst = 32'd201345868;
      14622: inst = 32'd203489279;
      14623: inst = 32'd471859200;
      14624: inst = 32'd136314880;
      14625: inst = 32'd268468224;
      14626: inst = 32'd201345869;
      14627: inst = 32'd203489279;
      14628: inst = 32'd471859200;
      14629: inst = 32'd136314880;
      14630: inst = 32'd268468224;
      14631: inst = 32'd201345870;
      14632: inst = 32'd203489279;
      14633: inst = 32'd471859200;
      14634: inst = 32'd136314880;
      14635: inst = 32'd268468224;
      14636: inst = 32'd201345871;
      14637: inst = 32'd203489279;
      14638: inst = 32'd471859200;
      14639: inst = 32'd136314880;
      14640: inst = 32'd268468224;
      14641: inst = 32'd201345872;
      14642: inst = 32'd203489279;
      14643: inst = 32'd471859200;
      14644: inst = 32'd136314880;
      14645: inst = 32'd268468224;
      14646: inst = 32'd201345873;
      14647: inst = 32'd203489279;
      14648: inst = 32'd471859200;
      14649: inst = 32'd136314880;
      14650: inst = 32'd268468224;
      14651: inst = 32'd201345874;
      14652: inst = 32'd203489279;
      14653: inst = 32'd471859200;
      14654: inst = 32'd136314880;
      14655: inst = 32'd268468224;
      14656: inst = 32'd201345875;
      14657: inst = 32'd203489279;
      14658: inst = 32'd471859200;
      14659: inst = 32'd136314880;
      14660: inst = 32'd268468224;
      14661: inst = 32'd201345876;
      14662: inst = 32'd203489279;
      14663: inst = 32'd471859200;
      14664: inst = 32'd136314880;
      14665: inst = 32'd268468224;
      14666: inst = 32'd201345877;
      14667: inst = 32'd203489279;
      14668: inst = 32'd471859200;
      14669: inst = 32'd136314880;
      14670: inst = 32'd268468224;
      14671: inst = 32'd201345878;
      14672: inst = 32'd203489279;
      14673: inst = 32'd471859200;
      14674: inst = 32'd136314880;
      14675: inst = 32'd268468224;
      14676: inst = 32'd201345879;
      14677: inst = 32'd203489279;
      14678: inst = 32'd471859200;
      14679: inst = 32'd136314880;
      14680: inst = 32'd268468224;
      14681: inst = 32'd201345880;
      14682: inst = 32'd203489279;
      14683: inst = 32'd471859200;
      14684: inst = 32'd136314880;
      14685: inst = 32'd268468224;
      14686: inst = 32'd201345881;
      14687: inst = 32'd203489279;
      14688: inst = 32'd471859200;
      14689: inst = 32'd136314880;
      14690: inst = 32'd268468224;
      14691: inst = 32'd201345882;
      14692: inst = 32'd203489279;
      14693: inst = 32'd471859200;
      14694: inst = 32'd136314880;
      14695: inst = 32'd268468224;
      14696: inst = 32'd201345883;
      14697: inst = 32'd203489279;
      14698: inst = 32'd471859200;
      14699: inst = 32'd136314880;
      14700: inst = 32'd268468224;
      14701: inst = 32'd201345884;
      14702: inst = 32'd203489279;
      14703: inst = 32'd471859200;
      14704: inst = 32'd136314880;
      14705: inst = 32'd268468224;
      14706: inst = 32'd201345885;
      14707: inst = 32'd203489279;
      14708: inst = 32'd471859200;
      14709: inst = 32'd136314880;
      14710: inst = 32'd268468224;
      14711: inst = 32'd201345886;
      14712: inst = 32'd203489279;
      14713: inst = 32'd471859200;
      14714: inst = 32'd136314880;
      14715: inst = 32'd268468224;
      14716: inst = 32'd201345887;
      14717: inst = 32'd203489279;
      14718: inst = 32'd471859200;
      14719: inst = 32'd136314880;
      14720: inst = 32'd268468224;
      14721: inst = 32'd201345888;
      14722: inst = 32'd203489279;
      14723: inst = 32'd471859200;
      14724: inst = 32'd136314880;
      14725: inst = 32'd268468224;
      14726: inst = 32'd201345889;
      14727: inst = 32'd203489279;
      14728: inst = 32'd471859200;
      14729: inst = 32'd136314880;
      14730: inst = 32'd268468224;
      14731: inst = 32'd201345890;
      14732: inst = 32'd203489279;
      14733: inst = 32'd471859200;
      14734: inst = 32'd136314880;
      14735: inst = 32'd268468224;
      14736: inst = 32'd201345891;
      14737: inst = 32'd203489279;
      14738: inst = 32'd471859200;
      14739: inst = 32'd136314880;
      14740: inst = 32'd268468224;
      14741: inst = 32'd201345892;
      14742: inst = 32'd203484854;
      14743: inst = 32'd471859200;
      14744: inst = 32'd136314880;
      14745: inst = 32'd268468224;
      14746: inst = 32'd201345893;
      14747: inst = 32'd203484854;
      14748: inst = 32'd471859200;
      14749: inst = 32'd136314880;
      14750: inst = 32'd268468224;
      14751: inst = 32'd201345894;
      14752: inst = 32'd203484854;
      14753: inst = 32'd471859200;
      14754: inst = 32'd136314880;
      14755: inst = 32'd268468224;
      14756: inst = 32'd201345895;
      14757: inst = 32'd203484854;
      14758: inst = 32'd471859200;
      14759: inst = 32'd136314880;
      14760: inst = 32'd268468224;
      14761: inst = 32'd201345896;
      14762: inst = 32'd203484854;
      14763: inst = 32'd471859200;
      14764: inst = 32'd136314880;
      14765: inst = 32'd268468224;
      14766: inst = 32'd201345897;
      14767: inst = 32'd203484854;
      14768: inst = 32'd471859200;
      14769: inst = 32'd136314880;
      14770: inst = 32'd268468224;
      14771: inst = 32'd201345898;
      14772: inst = 32'd203484854;
      14773: inst = 32'd471859200;
      14774: inst = 32'd136314880;
      14775: inst = 32'd268468224;
      14776: inst = 32'd201345899;
      14777: inst = 32'd203484854;
      14778: inst = 32'd471859200;
      14779: inst = 32'd136314880;
      14780: inst = 32'd268468224;
      14781: inst = 32'd201345900;
      14782: inst = 32'd203484854;
      14783: inst = 32'd471859200;
      14784: inst = 32'd136314880;
      14785: inst = 32'd268468224;
      14786: inst = 32'd201345901;
      14787: inst = 32'd203484854;
      14788: inst = 32'd471859200;
      14789: inst = 32'd136314880;
      14790: inst = 32'd268468224;
      14791: inst = 32'd201345902;
      14792: inst = 32'd203484854;
      14793: inst = 32'd471859200;
      14794: inst = 32'd136314880;
      14795: inst = 32'd268468224;
      14796: inst = 32'd201345903;
      14797: inst = 32'd203473634;
      14798: inst = 32'd471859200;
      14799: inst = 32'd136314880;
      14800: inst = 32'd268468224;
      14801: inst = 32'd201345904;
      14802: inst = 32'd203480005;
      14803: inst = 32'd471859200;
      14804: inst = 32'd136314880;
      14805: inst = 32'd268468224;
      14806: inst = 32'd201345905;
      14807: inst = 32'd203480005;
      14808: inst = 32'd471859200;
      14809: inst = 32'd136314880;
      14810: inst = 32'd268468224;
      14811: inst = 32'd201345906;
      14812: inst = 32'd203485052;
      14813: inst = 32'd471859200;
      14814: inst = 32'd136314880;
      14815: inst = 32'd268468224;
      14816: inst = 32'd201345907;
      14817: inst = 32'd203485052;
      14818: inst = 32'd471859200;
      14819: inst = 32'd136314880;
      14820: inst = 32'd268468224;
      14821: inst = 32'd201345908;
      14822: inst = 32'd203485052;
      14823: inst = 32'd471859200;
      14824: inst = 32'd136314880;
      14825: inst = 32'd268468224;
      14826: inst = 32'd201345909;
      14827: inst = 32'd203485052;
      14828: inst = 32'd471859200;
      14829: inst = 32'd136314880;
      14830: inst = 32'd268468224;
      14831: inst = 32'd201345910;
      14832: inst = 32'd203480005;
      14833: inst = 32'd471859200;
      14834: inst = 32'd136314880;
      14835: inst = 32'd268468224;
      14836: inst = 32'd201345911;
      14837: inst = 32'd203480005;
      14838: inst = 32'd471859200;
      14839: inst = 32'd136314880;
      14840: inst = 32'd268468224;
      14841: inst = 32'd201345912;
      14842: inst = 32'd203480005;
      14843: inst = 32'd471859200;
      14844: inst = 32'd136314880;
      14845: inst = 32'd268468224;
      14846: inst = 32'd201345913;
      14847: inst = 32'd203480005;
      14848: inst = 32'd471859200;
      14849: inst = 32'd136314880;
      14850: inst = 32'd268468224;
      14851: inst = 32'd201345914;
      14852: inst = 32'd203480005;
      14853: inst = 32'd471859200;
      14854: inst = 32'd136314880;
      14855: inst = 32'd268468224;
      14856: inst = 32'd201345915;
      14857: inst = 32'd203480005;
      14858: inst = 32'd471859200;
      14859: inst = 32'd136314880;
      14860: inst = 32'd268468224;
      14861: inst = 32'd201345916;
      14862: inst = 32'd203480005;
      14863: inst = 32'd471859200;
      14864: inst = 32'd136314880;
      14865: inst = 32'd268468224;
      14866: inst = 32'd201345917;
      14867: inst = 32'd203480005;
      14868: inst = 32'd471859200;
      14869: inst = 32'd136314880;
      14870: inst = 32'd268468224;
      14871: inst = 32'd201345918;
      14872: inst = 32'd203480005;
      14873: inst = 32'd471859200;
      14874: inst = 32'd136314880;
      14875: inst = 32'd268468224;
      14876: inst = 32'd201345919;
      14877: inst = 32'd203473634;
      14878: inst = 32'd471859200;
      14879: inst = 32'd136314880;
      14880: inst = 32'd268468224;
      14881: inst = 32'd201345920;
      14882: inst = 32'd203484854;
      14883: inst = 32'd471859200;
      14884: inst = 32'd136314880;
      14885: inst = 32'd268468224;
      14886: inst = 32'd201345921;
      14887: inst = 32'd203484854;
      14888: inst = 32'd471859200;
      14889: inst = 32'd136314880;
      14890: inst = 32'd268468224;
      14891: inst = 32'd201345922;
      14892: inst = 32'd203484854;
      14893: inst = 32'd471859200;
      14894: inst = 32'd136314880;
      14895: inst = 32'd268468224;
      14896: inst = 32'd201345923;
      14897: inst = 32'd203484854;
      14898: inst = 32'd471859200;
      14899: inst = 32'd136314880;
      14900: inst = 32'd268468224;
      14901: inst = 32'd201345924;
      14902: inst = 32'd203484854;
      14903: inst = 32'd471859200;
      14904: inst = 32'd136314880;
      14905: inst = 32'd268468224;
      14906: inst = 32'd201345925;
      14907: inst = 32'd203484854;
      14908: inst = 32'd471859200;
      14909: inst = 32'd136314880;
      14910: inst = 32'd268468224;
      14911: inst = 32'd201345926;
      14912: inst = 32'd203484854;
      14913: inst = 32'd471859200;
      14914: inst = 32'd136314880;
      14915: inst = 32'd268468224;
      14916: inst = 32'd201345927;
      14917: inst = 32'd203482875;
      14918: inst = 32'd471859200;
      14919: inst = 32'd136314880;
      14920: inst = 32'd268468224;
      14921: inst = 32'd201345928;
      14922: inst = 32'd203442793;
      14923: inst = 32'd471859200;
      14924: inst = 32'd136314880;
      14925: inst = 32'd268468224;
      14926: inst = 32'd201345929;
      14927: inst = 32'd203442793;
      14928: inst = 32'd471859200;
      14929: inst = 32'd136314880;
      14930: inst = 32'd268468224;
      14931: inst = 32'd201345930;
      14932: inst = 32'd203480827;
      14933: inst = 32'd471859200;
      14934: inst = 32'd136314880;
      14935: inst = 32'd268468224;
      14936: inst = 32'd201345931;
      14937: inst = 32'd203442793;
      14938: inst = 32'd471859200;
      14939: inst = 32'd136314880;
      14940: inst = 32'd268468224;
      14941: inst = 32'd201345932;
      14942: inst = 32'd203442793;
      14943: inst = 32'd471859200;
      14944: inst = 32'd136314880;
      14945: inst = 32'd268468224;
      14946: inst = 32'd201345933;
      14947: inst = 32'd203480827;
      14948: inst = 32'd471859200;
      14949: inst = 32'd136314880;
      14950: inst = 32'd268468224;
      14951: inst = 32'd201345934;
      14952: inst = 32'd203480827;
      14953: inst = 32'd471859200;
      14954: inst = 32'd136314880;
      14955: inst = 32'd268468224;
      14956: inst = 32'd201345935;
      14957: inst = 32'd203482875;
      14958: inst = 32'd471859200;
      14959: inst = 32'd136314880;
      14960: inst = 32'd268468224;
      14961: inst = 32'd201345936;
      14962: inst = 32'd203484854;
      14963: inst = 32'd471859200;
      14964: inst = 32'd136314880;
      14965: inst = 32'd268468224;
      14966: inst = 32'd201345937;
      14967: inst = 32'd203484854;
      14968: inst = 32'd471859200;
      14969: inst = 32'd136314880;
      14970: inst = 32'd268468224;
      14971: inst = 32'd201345938;
      14972: inst = 32'd203484854;
      14973: inst = 32'd471859200;
      14974: inst = 32'd136314880;
      14975: inst = 32'd268468224;
      14976: inst = 32'd201345939;
      14977: inst = 32'd203484854;
      14978: inst = 32'd471859200;
      14979: inst = 32'd136314880;
      14980: inst = 32'd268468224;
      14981: inst = 32'd201345940;
      14982: inst = 32'd203484854;
      14983: inst = 32'd471859200;
      14984: inst = 32'd136314880;
      14985: inst = 32'd268468224;
      14986: inst = 32'd201345941;
      14987: inst = 32'd203484854;
      14988: inst = 32'd471859200;
      14989: inst = 32'd136314880;
      14990: inst = 32'd268468224;
      14991: inst = 32'd201345942;
      14992: inst = 32'd203484854;
      14993: inst = 32'd471859200;
      14994: inst = 32'd136314880;
      14995: inst = 32'd268468224;
      14996: inst = 32'd201345943;
      14997: inst = 32'd203484854;
      14998: inst = 32'd471859200;
      14999: inst = 32'd136314880;
      15000: inst = 32'd268468224;
      15001: inst = 32'd201345944;
      15002: inst = 32'd203484854;
      15003: inst = 32'd471859200;
      15004: inst = 32'd136314880;
      15005: inst = 32'd268468224;
      15006: inst = 32'd201345945;
      15007: inst = 32'd203484854;
      15008: inst = 32'd471859200;
      15009: inst = 32'd136314880;
      15010: inst = 32'd268468224;
      15011: inst = 32'd201345946;
      15012: inst = 32'd203484854;
      15013: inst = 32'd471859200;
      15014: inst = 32'd136314880;
      15015: inst = 32'd268468224;
      15016: inst = 32'd201345947;
      15017: inst = 32'd203484854;
      15018: inst = 32'd471859200;
      15019: inst = 32'd136314880;
      15020: inst = 32'd268468224;
      15021: inst = 32'd201345948;
      15022: inst = 32'd203489279;
      15023: inst = 32'd471859200;
      15024: inst = 32'd136314880;
      15025: inst = 32'd268468224;
      15026: inst = 32'd201345949;
      15027: inst = 32'd203489279;
      15028: inst = 32'd471859200;
      15029: inst = 32'd136314880;
      15030: inst = 32'd268468224;
      15031: inst = 32'd201345950;
      15032: inst = 32'd203489279;
      15033: inst = 32'd471859200;
      15034: inst = 32'd136314880;
      15035: inst = 32'd268468224;
      15036: inst = 32'd201345951;
      15037: inst = 32'd203489279;
      15038: inst = 32'd471859200;
      15039: inst = 32'd136314880;
      15040: inst = 32'd268468224;
      15041: inst = 32'd201345952;
      15042: inst = 32'd203489279;
      15043: inst = 32'd471859200;
      15044: inst = 32'd136314880;
      15045: inst = 32'd268468224;
      15046: inst = 32'd201345953;
      15047: inst = 32'd203489279;
      15048: inst = 32'd471859200;
      15049: inst = 32'd136314880;
      15050: inst = 32'd268468224;
      15051: inst = 32'd201345954;
      15052: inst = 32'd203489279;
      15053: inst = 32'd471859200;
      15054: inst = 32'd136314880;
      15055: inst = 32'd268468224;
      15056: inst = 32'd201345955;
      15057: inst = 32'd203489279;
      15058: inst = 32'd471859200;
      15059: inst = 32'd136314880;
      15060: inst = 32'd268468224;
      15061: inst = 32'd201345956;
      15062: inst = 32'd203489279;
      15063: inst = 32'd471859200;
      15064: inst = 32'd136314880;
      15065: inst = 32'd268468224;
      15066: inst = 32'd201345957;
      15067: inst = 32'd203489279;
      15068: inst = 32'd471859200;
      15069: inst = 32'd136314880;
      15070: inst = 32'd268468224;
      15071: inst = 32'd201345958;
      15072: inst = 32'd203489279;
      15073: inst = 32'd471859200;
      15074: inst = 32'd136314880;
      15075: inst = 32'd268468224;
      15076: inst = 32'd201345959;
      15077: inst = 32'd203489279;
      15078: inst = 32'd471859200;
      15079: inst = 32'd136314880;
      15080: inst = 32'd268468224;
      15081: inst = 32'd201345960;
      15082: inst = 32'd203489279;
      15083: inst = 32'd471859200;
      15084: inst = 32'd136314880;
      15085: inst = 32'd268468224;
      15086: inst = 32'd201345961;
      15087: inst = 32'd203489279;
      15088: inst = 32'd471859200;
      15089: inst = 32'd136314880;
      15090: inst = 32'd268468224;
      15091: inst = 32'd201345962;
      15092: inst = 32'd203489279;
      15093: inst = 32'd471859200;
      15094: inst = 32'd136314880;
      15095: inst = 32'd268468224;
      15096: inst = 32'd201345963;
      15097: inst = 32'd203489279;
      15098: inst = 32'd471859200;
      15099: inst = 32'd136314880;
      15100: inst = 32'd268468224;
      15101: inst = 32'd201345964;
      15102: inst = 32'd203489279;
      15103: inst = 32'd471859200;
      15104: inst = 32'd136314880;
      15105: inst = 32'd268468224;
      15106: inst = 32'd201345965;
      15107: inst = 32'd203489279;
      15108: inst = 32'd471859200;
      15109: inst = 32'd136314880;
      15110: inst = 32'd268468224;
      15111: inst = 32'd201345966;
      15112: inst = 32'd203489279;
      15113: inst = 32'd471859200;
      15114: inst = 32'd136314880;
      15115: inst = 32'd268468224;
      15116: inst = 32'd201345967;
      15117: inst = 32'd203489279;
      15118: inst = 32'd471859200;
      15119: inst = 32'd136314880;
      15120: inst = 32'd268468224;
      15121: inst = 32'd201345968;
      15122: inst = 32'd203489279;
      15123: inst = 32'd471859200;
      15124: inst = 32'd136314880;
      15125: inst = 32'd268468224;
      15126: inst = 32'd201345969;
      15127: inst = 32'd203489279;
      15128: inst = 32'd471859200;
      15129: inst = 32'd136314880;
      15130: inst = 32'd268468224;
      15131: inst = 32'd201345970;
      15132: inst = 32'd203489279;
      15133: inst = 32'd471859200;
      15134: inst = 32'd136314880;
      15135: inst = 32'd268468224;
      15136: inst = 32'd201345971;
      15137: inst = 32'd203489279;
      15138: inst = 32'd471859200;
      15139: inst = 32'd136314880;
      15140: inst = 32'd268468224;
      15141: inst = 32'd201345972;
      15142: inst = 32'd203489279;
      15143: inst = 32'd471859200;
      15144: inst = 32'd136314880;
      15145: inst = 32'd268468224;
      15146: inst = 32'd201345973;
      15147: inst = 32'd203489279;
      15148: inst = 32'd471859200;
      15149: inst = 32'd136314880;
      15150: inst = 32'd268468224;
      15151: inst = 32'd201345974;
      15152: inst = 32'd203489279;
      15153: inst = 32'd471859200;
      15154: inst = 32'd136314880;
      15155: inst = 32'd268468224;
      15156: inst = 32'd201345975;
      15157: inst = 32'd203489279;
      15158: inst = 32'd471859200;
      15159: inst = 32'd136314880;
      15160: inst = 32'd268468224;
      15161: inst = 32'd201345976;
      15162: inst = 32'd203489279;
      15163: inst = 32'd471859200;
      15164: inst = 32'd136314880;
      15165: inst = 32'd268468224;
      15166: inst = 32'd201345977;
      15167: inst = 32'd203489279;
      15168: inst = 32'd471859200;
      15169: inst = 32'd136314880;
      15170: inst = 32'd268468224;
      15171: inst = 32'd201345978;
      15172: inst = 32'd203489279;
      15173: inst = 32'd471859200;
      15174: inst = 32'd136314880;
      15175: inst = 32'd268468224;
      15176: inst = 32'd201345979;
      15177: inst = 32'd203489279;
      15178: inst = 32'd471859200;
      15179: inst = 32'd136314880;
      15180: inst = 32'd268468224;
      15181: inst = 32'd201345980;
      15182: inst = 32'd203489279;
      15183: inst = 32'd471859200;
      15184: inst = 32'd136314880;
      15185: inst = 32'd268468224;
      15186: inst = 32'd201345981;
      15187: inst = 32'd203489279;
      15188: inst = 32'd471859200;
      15189: inst = 32'd136314880;
      15190: inst = 32'd268468224;
      15191: inst = 32'd201345982;
      15192: inst = 32'd203489279;
      15193: inst = 32'd471859200;
      15194: inst = 32'd136314880;
      15195: inst = 32'd268468224;
      15196: inst = 32'd201345983;
      15197: inst = 32'd203489279;
      15198: inst = 32'd471859200;
      15199: inst = 32'd136314880;
      15200: inst = 32'd268468224;
      15201: inst = 32'd201345984;
      15202: inst = 32'd203489279;
      15203: inst = 32'd471859200;
      15204: inst = 32'd136314880;
      15205: inst = 32'd268468224;
      15206: inst = 32'd201345985;
      15207: inst = 32'd203489279;
      15208: inst = 32'd471859200;
      15209: inst = 32'd136314880;
      15210: inst = 32'd268468224;
      15211: inst = 32'd201345986;
      15212: inst = 32'd203489279;
      15213: inst = 32'd471859200;
      15214: inst = 32'd136314880;
      15215: inst = 32'd268468224;
      15216: inst = 32'd201345987;
      15217: inst = 32'd203489279;
      15218: inst = 32'd471859200;
      15219: inst = 32'd136314880;
      15220: inst = 32'd268468224;
      15221: inst = 32'd201345988;
      15222: inst = 32'd203484854;
      15223: inst = 32'd471859200;
      15224: inst = 32'd136314880;
      15225: inst = 32'd268468224;
      15226: inst = 32'd201345989;
      15227: inst = 32'd203484854;
      15228: inst = 32'd471859200;
      15229: inst = 32'd136314880;
      15230: inst = 32'd268468224;
      15231: inst = 32'd201345990;
      15232: inst = 32'd203484854;
      15233: inst = 32'd471859200;
      15234: inst = 32'd136314880;
      15235: inst = 32'd268468224;
      15236: inst = 32'd201345991;
      15237: inst = 32'd203484854;
      15238: inst = 32'd471859200;
      15239: inst = 32'd136314880;
      15240: inst = 32'd268468224;
      15241: inst = 32'd201345992;
      15242: inst = 32'd203484854;
      15243: inst = 32'd471859200;
      15244: inst = 32'd136314880;
      15245: inst = 32'd268468224;
      15246: inst = 32'd201345993;
      15247: inst = 32'd203484854;
      15248: inst = 32'd471859200;
      15249: inst = 32'd136314880;
      15250: inst = 32'd268468224;
      15251: inst = 32'd201345994;
      15252: inst = 32'd203484854;
      15253: inst = 32'd471859200;
      15254: inst = 32'd136314880;
      15255: inst = 32'd268468224;
      15256: inst = 32'd201345995;
      15257: inst = 32'd203484854;
      15258: inst = 32'd471859200;
      15259: inst = 32'd136314880;
      15260: inst = 32'd268468224;
      15261: inst = 32'd201345996;
      15262: inst = 32'd203484854;
      15263: inst = 32'd471859200;
      15264: inst = 32'd136314880;
      15265: inst = 32'd268468224;
      15266: inst = 32'd201345997;
      15267: inst = 32'd203484854;
      15268: inst = 32'd471859200;
      15269: inst = 32'd136314880;
      15270: inst = 32'd268468224;
      15271: inst = 32'd201345998;
      15272: inst = 32'd203484854;
      15273: inst = 32'd471859200;
      15274: inst = 32'd136314880;
      15275: inst = 32'd268468224;
      15276: inst = 32'd201345999;
      15277: inst = 32'd203473634;
      15278: inst = 32'd471859200;
      15279: inst = 32'd136314880;
      15280: inst = 32'd268468224;
      15281: inst = 32'd201346000;
      15282: inst = 32'd203480005;
      15283: inst = 32'd471859200;
      15284: inst = 32'd136314880;
      15285: inst = 32'd268468224;
      15286: inst = 32'd201346001;
      15287: inst = 32'd203480005;
      15288: inst = 32'd471859200;
      15289: inst = 32'd136314880;
      15290: inst = 32'd268468224;
      15291: inst = 32'd201346002;
      15292: inst = 32'd203480005;
      15293: inst = 32'd471859200;
      15294: inst = 32'd136314880;
      15295: inst = 32'd268468224;
      15296: inst = 32'd201346003;
      15297: inst = 32'd203480005;
      15298: inst = 32'd471859200;
      15299: inst = 32'd136314880;
      15300: inst = 32'd268468224;
      15301: inst = 32'd201346004;
      15302: inst = 32'd203480005;
      15303: inst = 32'd471859200;
      15304: inst = 32'd136314880;
      15305: inst = 32'd268468224;
      15306: inst = 32'd201346005;
      15307: inst = 32'd203480005;
      15308: inst = 32'd471859200;
      15309: inst = 32'd136314880;
      15310: inst = 32'd268468224;
      15311: inst = 32'd201346006;
      15312: inst = 32'd203480005;
      15313: inst = 32'd471859200;
      15314: inst = 32'd136314880;
      15315: inst = 32'd268468224;
      15316: inst = 32'd201346007;
      15317: inst = 32'd203480005;
      15318: inst = 32'd471859200;
      15319: inst = 32'd136314880;
      15320: inst = 32'd268468224;
      15321: inst = 32'd201346008;
      15322: inst = 32'd203480005;
      15323: inst = 32'd471859200;
      15324: inst = 32'd136314880;
      15325: inst = 32'd268468224;
      15326: inst = 32'd201346009;
      15327: inst = 32'd203480005;
      15328: inst = 32'd471859200;
      15329: inst = 32'd136314880;
      15330: inst = 32'd268468224;
      15331: inst = 32'd201346010;
      15332: inst = 32'd203480005;
      15333: inst = 32'd471859200;
      15334: inst = 32'd136314880;
      15335: inst = 32'd268468224;
      15336: inst = 32'd201346011;
      15337: inst = 32'd203480005;
      15338: inst = 32'd471859200;
      15339: inst = 32'd136314880;
      15340: inst = 32'd268468224;
      15341: inst = 32'd201346012;
      15342: inst = 32'd203480005;
      15343: inst = 32'd471859200;
      15344: inst = 32'd136314880;
      15345: inst = 32'd268468224;
      15346: inst = 32'd201346013;
      15347: inst = 32'd203480005;
      15348: inst = 32'd471859200;
      15349: inst = 32'd136314880;
      15350: inst = 32'd268468224;
      15351: inst = 32'd201346014;
      15352: inst = 32'd203480005;
      15353: inst = 32'd471859200;
      15354: inst = 32'd136314880;
      15355: inst = 32'd268468224;
      15356: inst = 32'd201346015;
      15357: inst = 32'd203473634;
      15358: inst = 32'd471859200;
      15359: inst = 32'd136314880;
      15360: inst = 32'd268468224;
      15361: inst = 32'd201346016;
      15362: inst = 32'd203484854;
      15363: inst = 32'd471859200;
      15364: inst = 32'd136314880;
      15365: inst = 32'd268468224;
      15366: inst = 32'd201346017;
      15367: inst = 32'd203484854;
      15368: inst = 32'd471859200;
      15369: inst = 32'd136314880;
      15370: inst = 32'd268468224;
      15371: inst = 32'd201346018;
      15372: inst = 32'd203484854;
      15373: inst = 32'd471859200;
      15374: inst = 32'd136314880;
      15375: inst = 32'd268468224;
      15376: inst = 32'd201346019;
      15377: inst = 32'd203484854;
      15378: inst = 32'd471859200;
      15379: inst = 32'd136314880;
      15380: inst = 32'd268468224;
      15381: inst = 32'd201346020;
      15382: inst = 32'd203484854;
      15383: inst = 32'd471859200;
      15384: inst = 32'd136314880;
      15385: inst = 32'd268468224;
      15386: inst = 32'd201346021;
      15387: inst = 32'd203484854;
      15388: inst = 32'd471859200;
      15389: inst = 32'd136314880;
      15390: inst = 32'd268468224;
      15391: inst = 32'd201346022;
      15392: inst = 32'd203484854;
      15393: inst = 32'd471859200;
      15394: inst = 32'd136314880;
      15395: inst = 32'd268468224;
      15396: inst = 32'd201346023;
      15397: inst = 32'd203482874;
      15398: inst = 32'd471859200;
      15399: inst = 32'd136314880;
      15400: inst = 32'd268468224;
      15401: inst = 32'd201346024;
      15402: inst = 32'd203480827;
      15403: inst = 32'd471859200;
      15404: inst = 32'd136314880;
      15405: inst = 32'd268468224;
      15406: inst = 32'd201346025;
      15407: inst = 32'd203480827;
      15408: inst = 32'd471859200;
      15409: inst = 32'd136314880;
      15410: inst = 32'd268468224;
      15411: inst = 32'd201346026;
      15412: inst = 32'd203480827;
      15413: inst = 32'd471859200;
      15414: inst = 32'd136314880;
      15415: inst = 32'd268468224;
      15416: inst = 32'd201346027;
      15417: inst = 32'd203480827;
      15418: inst = 32'd471859200;
      15419: inst = 32'd136314880;
      15420: inst = 32'd268468224;
      15421: inst = 32'd201346028;
      15422: inst = 32'd203480827;
      15423: inst = 32'd471859200;
      15424: inst = 32'd136314880;
      15425: inst = 32'd268468224;
      15426: inst = 32'd201346029;
      15427: inst = 32'd203480827;
      15428: inst = 32'd471859200;
      15429: inst = 32'd136314880;
      15430: inst = 32'd268468224;
      15431: inst = 32'd201346030;
      15432: inst = 32'd203480827;
      15433: inst = 32'd471859200;
      15434: inst = 32'd136314880;
      15435: inst = 32'd268468224;
      15436: inst = 32'd201346031;
      15437: inst = 32'd203482841;
      15438: inst = 32'd471859200;
      15439: inst = 32'd136314880;
      15440: inst = 32'd268468224;
      15441: inst = 32'd201346032;
      15442: inst = 32'd203484854;
      15443: inst = 32'd471859200;
      15444: inst = 32'd136314880;
      15445: inst = 32'd268468224;
      15446: inst = 32'd201346033;
      15447: inst = 32'd203484854;
      15448: inst = 32'd471859200;
      15449: inst = 32'd136314880;
      15450: inst = 32'd268468224;
      15451: inst = 32'd201346034;
      15452: inst = 32'd203484854;
      15453: inst = 32'd471859200;
      15454: inst = 32'd136314880;
      15455: inst = 32'd268468224;
      15456: inst = 32'd201346035;
      15457: inst = 32'd203484854;
      15458: inst = 32'd471859200;
      15459: inst = 32'd136314880;
      15460: inst = 32'd268468224;
      15461: inst = 32'd201346036;
      15462: inst = 32'd203484854;
      15463: inst = 32'd471859200;
      15464: inst = 32'd136314880;
      15465: inst = 32'd268468224;
      15466: inst = 32'd201346037;
      15467: inst = 32'd203484854;
      15468: inst = 32'd471859200;
      15469: inst = 32'd136314880;
      15470: inst = 32'd268468224;
      15471: inst = 32'd201346038;
      15472: inst = 32'd203484854;
      15473: inst = 32'd471859200;
      15474: inst = 32'd136314880;
      15475: inst = 32'd268468224;
      15476: inst = 32'd201346039;
      15477: inst = 32'd203484854;
      15478: inst = 32'd471859200;
      15479: inst = 32'd136314880;
      15480: inst = 32'd268468224;
      15481: inst = 32'd201346040;
      15482: inst = 32'd203484854;
      15483: inst = 32'd471859200;
      15484: inst = 32'd136314880;
      15485: inst = 32'd268468224;
      15486: inst = 32'd201346041;
      15487: inst = 32'd203484854;
      15488: inst = 32'd471859200;
      15489: inst = 32'd136314880;
      15490: inst = 32'd268468224;
      15491: inst = 32'd201346042;
      15492: inst = 32'd203470230;
      15493: inst = 32'd471859200;
      15494: inst = 32'd136314880;
      15495: inst = 32'd268468224;
      15496: inst = 32'd201346043;
      15497: inst = 32'd203470230;
      15498: inst = 32'd471859200;
      15499: inst = 32'd136314880;
      15500: inst = 32'd268468224;
      15501: inst = 32'd201346044;
      15502: inst = 32'd203470230;
      15503: inst = 32'd471859200;
      15504: inst = 32'd136314880;
      15505: inst = 32'd268468224;
      15506: inst = 32'd201346045;
      15507: inst = 32'd203470230;
      15508: inst = 32'd471859200;
      15509: inst = 32'd136314880;
      15510: inst = 32'd268468224;
      15511: inst = 32'd201346046;
      15512: inst = 32'd203470230;
      15513: inst = 32'd471859200;
      15514: inst = 32'd136314880;
      15515: inst = 32'd268468224;
      15516: inst = 32'd201346047;
      15517: inst = 32'd203470230;
      15518: inst = 32'd471859200;
      15519: inst = 32'd136314880;
      15520: inst = 32'd268468224;
      15521: inst = 32'd201346048;
      15522: inst = 32'd203470230;
      15523: inst = 32'd471859200;
      15524: inst = 32'd136314880;
      15525: inst = 32'd268468224;
      15526: inst = 32'd201346049;
      15527: inst = 32'd203470230;
      15528: inst = 32'd471859200;
      15529: inst = 32'd136314880;
      15530: inst = 32'd268468224;
      15531: inst = 32'd201346050;
      15532: inst = 32'd203470230;
      15533: inst = 32'd471859200;
      15534: inst = 32'd136314880;
      15535: inst = 32'd268468224;
      15536: inst = 32'd201346051;
      15537: inst = 32'd203470230;
      15538: inst = 32'd471859200;
      15539: inst = 32'd136314880;
      15540: inst = 32'd268468224;
      15541: inst = 32'd201346052;
      15542: inst = 32'd203470230;
      15543: inst = 32'd471859200;
      15544: inst = 32'd136314880;
      15545: inst = 32'd268468224;
      15546: inst = 32'd201346053;
      15547: inst = 32'd203470230;
      15548: inst = 32'd471859200;
      15549: inst = 32'd136314880;
      15550: inst = 32'd268468224;
      15551: inst = 32'd201346054;
      15552: inst = 32'd203470230;
      15553: inst = 32'd471859200;
      15554: inst = 32'd136314880;
      15555: inst = 32'd268468224;
      15556: inst = 32'd201346055;
      15557: inst = 32'd203470230;
      15558: inst = 32'd471859200;
      15559: inst = 32'd136314880;
      15560: inst = 32'd268468224;
      15561: inst = 32'd201346056;
      15562: inst = 32'd203470230;
      15563: inst = 32'd471859200;
      15564: inst = 32'd136314880;
      15565: inst = 32'd268468224;
      15566: inst = 32'd201346057;
      15567: inst = 32'd203470230;
      15568: inst = 32'd471859200;
      15569: inst = 32'd136314880;
      15570: inst = 32'd268468224;
      15571: inst = 32'd201346058;
      15572: inst = 32'd203470230;
      15573: inst = 32'd471859200;
      15574: inst = 32'd136314880;
      15575: inst = 32'd268468224;
      15576: inst = 32'd201346059;
      15577: inst = 32'd203470230;
      15578: inst = 32'd471859200;
      15579: inst = 32'd136314880;
      15580: inst = 32'd268468224;
      15581: inst = 32'd201346060;
      15582: inst = 32'd203470230;
      15583: inst = 32'd471859200;
      15584: inst = 32'd136314880;
      15585: inst = 32'd268468224;
      15586: inst = 32'd201346061;
      15587: inst = 32'd203470230;
      15588: inst = 32'd471859200;
      15589: inst = 32'd136314880;
      15590: inst = 32'd268468224;
      15591: inst = 32'd201346062;
      15592: inst = 32'd203470230;
      15593: inst = 32'd471859200;
      15594: inst = 32'd136314880;
      15595: inst = 32'd268468224;
      15596: inst = 32'd201346063;
      15597: inst = 32'd203470230;
      15598: inst = 32'd471859200;
      15599: inst = 32'd136314880;
      15600: inst = 32'd268468224;
      15601: inst = 32'd201346064;
      15602: inst = 32'd203470230;
      15603: inst = 32'd471859200;
      15604: inst = 32'd136314880;
      15605: inst = 32'd268468224;
      15606: inst = 32'd201346065;
      15607: inst = 32'd203470230;
      15608: inst = 32'd471859200;
      15609: inst = 32'd136314880;
      15610: inst = 32'd268468224;
      15611: inst = 32'd201346066;
      15612: inst = 32'd203470230;
      15613: inst = 32'd471859200;
      15614: inst = 32'd136314880;
      15615: inst = 32'd268468224;
      15616: inst = 32'd201346067;
      15617: inst = 32'd203470230;
      15618: inst = 32'd471859200;
      15619: inst = 32'd136314880;
      15620: inst = 32'd268468224;
      15621: inst = 32'd201346068;
      15622: inst = 32'd203470230;
      15623: inst = 32'd471859200;
      15624: inst = 32'd136314880;
      15625: inst = 32'd268468224;
      15626: inst = 32'd201346069;
      15627: inst = 32'd203470230;
      15628: inst = 32'd471859200;
      15629: inst = 32'd136314880;
      15630: inst = 32'd268468224;
      15631: inst = 32'd201346070;
      15632: inst = 32'd203470230;
      15633: inst = 32'd471859200;
      15634: inst = 32'd136314880;
      15635: inst = 32'd268468224;
      15636: inst = 32'd201346071;
      15637: inst = 32'd203470230;
      15638: inst = 32'd471859200;
      15639: inst = 32'd136314880;
      15640: inst = 32'd268468224;
      15641: inst = 32'd201346072;
      15642: inst = 32'd203470230;
      15643: inst = 32'd471859200;
      15644: inst = 32'd136314880;
      15645: inst = 32'd268468224;
      15646: inst = 32'd201346073;
      15647: inst = 32'd203470230;
      15648: inst = 32'd471859200;
      15649: inst = 32'd136314880;
      15650: inst = 32'd268468224;
      15651: inst = 32'd201346074;
      15652: inst = 32'd203470230;
      15653: inst = 32'd471859200;
      15654: inst = 32'd136314880;
      15655: inst = 32'd268468224;
      15656: inst = 32'd201346075;
      15657: inst = 32'd203470230;
      15658: inst = 32'd471859200;
      15659: inst = 32'd136314880;
      15660: inst = 32'd268468224;
      15661: inst = 32'd201346076;
      15662: inst = 32'd203470230;
      15663: inst = 32'd471859200;
      15664: inst = 32'd136314880;
      15665: inst = 32'd268468224;
      15666: inst = 32'd201346077;
      15667: inst = 32'd203470230;
      15668: inst = 32'd471859200;
      15669: inst = 32'd136314880;
      15670: inst = 32'd268468224;
      15671: inst = 32'd201346078;
      15672: inst = 32'd203470230;
      15673: inst = 32'd471859200;
      15674: inst = 32'd136314880;
      15675: inst = 32'd268468224;
      15676: inst = 32'd201346079;
      15677: inst = 32'd203470230;
      15678: inst = 32'd471859200;
      15679: inst = 32'd136314880;
      15680: inst = 32'd268468224;
      15681: inst = 32'd201346080;
      15682: inst = 32'd203470230;
      15683: inst = 32'd471859200;
      15684: inst = 32'd136314880;
      15685: inst = 32'd268468224;
      15686: inst = 32'd201346081;
      15687: inst = 32'd203470230;
      15688: inst = 32'd471859200;
      15689: inst = 32'd136314880;
      15690: inst = 32'd268468224;
      15691: inst = 32'd201346082;
      15692: inst = 32'd203470230;
      15693: inst = 32'd471859200;
      15694: inst = 32'd136314880;
      15695: inst = 32'd268468224;
      15696: inst = 32'd201346083;
      15697: inst = 32'd203470230;
      15698: inst = 32'd471859200;
      15699: inst = 32'd136314880;
      15700: inst = 32'd268468224;
      15701: inst = 32'd201346084;
      15702: inst = 32'd203470230;
      15703: inst = 32'd471859200;
      15704: inst = 32'd136314880;
      15705: inst = 32'd268468224;
      15706: inst = 32'd201346085;
      15707: inst = 32'd203470230;
      15708: inst = 32'd471859200;
      15709: inst = 32'd136314880;
      15710: inst = 32'd268468224;
      15711: inst = 32'd201346086;
      15712: inst = 32'd203484854;
      15713: inst = 32'd471859200;
      15714: inst = 32'd136314880;
      15715: inst = 32'd268468224;
      15716: inst = 32'd201346087;
      15717: inst = 32'd203484854;
      15718: inst = 32'd471859200;
      15719: inst = 32'd136314880;
      15720: inst = 32'd268468224;
      15721: inst = 32'd201346088;
      15722: inst = 32'd203484854;
      15723: inst = 32'd471859200;
      15724: inst = 32'd136314880;
      15725: inst = 32'd268468224;
      15726: inst = 32'd201346089;
      15727: inst = 32'd203484854;
      15728: inst = 32'd471859200;
      15729: inst = 32'd136314880;
      15730: inst = 32'd268468224;
      15731: inst = 32'd201346090;
      15732: inst = 32'd203484854;
      15733: inst = 32'd471859200;
      15734: inst = 32'd136314880;
      15735: inst = 32'd268468224;
      15736: inst = 32'd201346091;
      15737: inst = 32'd203484854;
      15738: inst = 32'd471859200;
      15739: inst = 32'd136314880;
      15740: inst = 32'd268468224;
      15741: inst = 32'd201346092;
      15742: inst = 32'd203484854;
      15743: inst = 32'd471859200;
      15744: inst = 32'd136314880;
      15745: inst = 32'd268468224;
      15746: inst = 32'd201346093;
      15747: inst = 32'd203484854;
      15748: inst = 32'd471859200;
      15749: inst = 32'd136314880;
      15750: inst = 32'd268468224;
      15751: inst = 32'd201346094;
      15752: inst = 32'd203484854;
      15753: inst = 32'd471859200;
      15754: inst = 32'd136314880;
      15755: inst = 32'd268468224;
      15756: inst = 32'd201346095;
      15757: inst = 32'd203473634;
      15758: inst = 32'd471859200;
      15759: inst = 32'd136314880;
      15760: inst = 32'd268468224;
      15761: inst = 32'd201346096;
      15762: inst = 32'd203480005;
      15763: inst = 32'd471859200;
      15764: inst = 32'd136314880;
      15765: inst = 32'd268468224;
      15766: inst = 32'd201346097;
      15767: inst = 32'd203480005;
      15768: inst = 32'd471859200;
      15769: inst = 32'd136314880;
      15770: inst = 32'd268468224;
      15771: inst = 32'd201346098;
      15772: inst = 32'd203480005;
      15773: inst = 32'd471859200;
      15774: inst = 32'd136314880;
      15775: inst = 32'd268468224;
      15776: inst = 32'd201346099;
      15777: inst = 32'd203480005;
      15778: inst = 32'd471859200;
      15779: inst = 32'd136314880;
      15780: inst = 32'd268468224;
      15781: inst = 32'd201346100;
      15782: inst = 32'd203480005;
      15783: inst = 32'd471859200;
      15784: inst = 32'd136314880;
      15785: inst = 32'd268468224;
      15786: inst = 32'd201346101;
      15787: inst = 32'd203480005;
      15788: inst = 32'd471859200;
      15789: inst = 32'd136314880;
      15790: inst = 32'd268468224;
      15791: inst = 32'd201346102;
      15792: inst = 32'd203480005;
      15793: inst = 32'd471859200;
      15794: inst = 32'd136314880;
      15795: inst = 32'd268468224;
      15796: inst = 32'd201346103;
      15797: inst = 32'd203480005;
      15798: inst = 32'd471859200;
      15799: inst = 32'd136314880;
      15800: inst = 32'd268468224;
      15801: inst = 32'd201346104;
      15802: inst = 32'd203480005;
      15803: inst = 32'd471859200;
      15804: inst = 32'd136314880;
      15805: inst = 32'd268468224;
      15806: inst = 32'd201346105;
      15807: inst = 32'd203480005;
      15808: inst = 32'd471859200;
      15809: inst = 32'd136314880;
      15810: inst = 32'd268468224;
      15811: inst = 32'd201346106;
      15812: inst = 32'd203480005;
      15813: inst = 32'd471859200;
      15814: inst = 32'd136314880;
      15815: inst = 32'd268468224;
      15816: inst = 32'd201346107;
      15817: inst = 32'd203480005;
      15818: inst = 32'd471859200;
      15819: inst = 32'd136314880;
      15820: inst = 32'd268468224;
      15821: inst = 32'd201346108;
      15822: inst = 32'd203480005;
      15823: inst = 32'd471859200;
      15824: inst = 32'd136314880;
      15825: inst = 32'd268468224;
      15826: inst = 32'd201346109;
      15827: inst = 32'd203480005;
      15828: inst = 32'd471859200;
      15829: inst = 32'd136314880;
      15830: inst = 32'd268468224;
      15831: inst = 32'd201346110;
      15832: inst = 32'd203480005;
      15833: inst = 32'd471859200;
      15834: inst = 32'd136314880;
      15835: inst = 32'd268468224;
      15836: inst = 32'd201346111;
      15837: inst = 32'd203473634;
      15838: inst = 32'd471859200;
      15839: inst = 32'd136314880;
      15840: inst = 32'd268468224;
      15841: inst = 32'd201346112;
      15842: inst = 32'd203484854;
      15843: inst = 32'd471859200;
      15844: inst = 32'd136314880;
      15845: inst = 32'd268468224;
      15846: inst = 32'd201346113;
      15847: inst = 32'd203484854;
      15848: inst = 32'd471859200;
      15849: inst = 32'd136314880;
      15850: inst = 32'd268468224;
      15851: inst = 32'd201346114;
      15852: inst = 32'd203484854;
      15853: inst = 32'd471859200;
      15854: inst = 32'd136314880;
      15855: inst = 32'd268468224;
      15856: inst = 32'd201346115;
      15857: inst = 32'd203484854;
      15858: inst = 32'd471859200;
      15859: inst = 32'd136314880;
      15860: inst = 32'd268468224;
      15861: inst = 32'd201346116;
      15862: inst = 32'd203484854;
      15863: inst = 32'd471859200;
      15864: inst = 32'd136314880;
      15865: inst = 32'd268468224;
      15866: inst = 32'd201346117;
      15867: inst = 32'd203484854;
      15868: inst = 32'd471859200;
      15869: inst = 32'd136314880;
      15870: inst = 32'd268468224;
      15871: inst = 32'd201346118;
      15872: inst = 32'd203484854;
      15873: inst = 32'd471859200;
      15874: inst = 32'd136314880;
      15875: inst = 32'd268468224;
      15876: inst = 32'd201346119;
      15877: inst = 32'd203484855;
      15878: inst = 32'd471859200;
      15879: inst = 32'd136314880;
      15880: inst = 32'd268468224;
      15881: inst = 32'd201346120;
      15882: inst = 32'd203442793;
      15883: inst = 32'd471859200;
      15884: inst = 32'd136314880;
      15885: inst = 32'd268468224;
      15886: inst = 32'd201346121;
      15887: inst = 32'd203480827;
      15888: inst = 32'd471859200;
      15889: inst = 32'd136314880;
      15890: inst = 32'd268468224;
      15891: inst = 32'd201346122;
      15892: inst = 32'd203442793;
      15893: inst = 32'd471859200;
      15894: inst = 32'd136314880;
      15895: inst = 32'd268468224;
      15896: inst = 32'd201346123;
      15897: inst = 32'd203480827;
      15898: inst = 32'd471859200;
      15899: inst = 32'd136314880;
      15900: inst = 32'd268468224;
      15901: inst = 32'd201346124;
      15902: inst = 32'd203442793;
      15903: inst = 32'd471859200;
      15904: inst = 32'd136314880;
      15905: inst = 32'd268468224;
      15906: inst = 32'd201346125;
      15907: inst = 32'd203482875;
      15908: inst = 32'd471859200;
      15909: inst = 32'd136314880;
      15910: inst = 32'd268468224;
      15911: inst = 32'd201346126;
      15912: inst = 32'd203482841;
      15913: inst = 32'd471859200;
      15914: inst = 32'd136314880;
      15915: inst = 32'd268468224;
      15916: inst = 32'd201346127;
      15917: inst = 32'd203484854;
      15918: inst = 32'd471859200;
      15919: inst = 32'd136314880;
      15920: inst = 32'd268468224;
      15921: inst = 32'd201346128;
      15922: inst = 32'd203484854;
      15923: inst = 32'd471859200;
      15924: inst = 32'd136314880;
      15925: inst = 32'd268468224;
      15926: inst = 32'd201346129;
      15927: inst = 32'd203484854;
      15928: inst = 32'd471859200;
      15929: inst = 32'd136314880;
      15930: inst = 32'd268468224;
      15931: inst = 32'd201346130;
      15932: inst = 32'd203484854;
      15933: inst = 32'd471859200;
      15934: inst = 32'd136314880;
      15935: inst = 32'd268468224;
      15936: inst = 32'd201346131;
      15937: inst = 32'd203484854;
      15938: inst = 32'd471859200;
      15939: inst = 32'd136314880;
      15940: inst = 32'd268468224;
      15941: inst = 32'd201346132;
      15942: inst = 32'd203484854;
      15943: inst = 32'd471859200;
      15944: inst = 32'd136314880;
      15945: inst = 32'd268468224;
      15946: inst = 32'd201346133;
      15947: inst = 32'd203484854;
      15948: inst = 32'd471859200;
      15949: inst = 32'd136314880;
      15950: inst = 32'd268468224;
      15951: inst = 32'd201346134;
      15952: inst = 32'd203484854;
      15953: inst = 32'd471859200;
      15954: inst = 32'd136314880;
      15955: inst = 32'd268468224;
      15956: inst = 32'd201346135;
      15957: inst = 32'd203484854;
      15958: inst = 32'd471859200;
      15959: inst = 32'd136314880;
      15960: inst = 32'd268468224;
      15961: inst = 32'd201346136;
      15962: inst = 32'd203484854;
      15963: inst = 32'd471859200;
      15964: inst = 32'd136314880;
      15965: inst = 32'd268468224;
      15966: inst = 32'd201346137;
      15967: inst = 32'd203484854;
      15968: inst = 32'd471859200;
      15969: inst = 32'd136314880;
      15970: inst = 32'd268468224;
      15971: inst = 32'd201346138;
      15972: inst = 32'd203484854;
      15973: inst = 32'd471859200;
      15974: inst = 32'd136314880;
      15975: inst = 32'd268468224;
      15976: inst = 32'd201346139;
      15977: inst = 32'd203484854;
      15978: inst = 32'd471859200;
      15979: inst = 32'd136314880;
      15980: inst = 32'd268468224;
      15981: inst = 32'd201346140;
      15982: inst = 32'd203484854;
      15983: inst = 32'd471859200;
      15984: inst = 32'd136314880;
      15985: inst = 32'd268468224;
      15986: inst = 32'd201346141;
      15987: inst = 32'd203484854;
      15988: inst = 32'd471859200;
      15989: inst = 32'd136314880;
      15990: inst = 32'd268468224;
      15991: inst = 32'd201346142;
      15992: inst = 32'd203484854;
      15993: inst = 32'd471859200;
      15994: inst = 32'd136314880;
      15995: inst = 32'd268468224;
      15996: inst = 32'd201346143;
      15997: inst = 32'd203484854;
      15998: inst = 32'd471859200;
      15999: inst = 32'd136314880;
      16000: inst = 32'd268468224;
      16001: inst = 32'd201346144;
      16002: inst = 32'd203484854;
      16003: inst = 32'd471859200;
      16004: inst = 32'd136314880;
      16005: inst = 32'd268468224;
      16006: inst = 32'd201346145;
      16007: inst = 32'd203484854;
      16008: inst = 32'd471859200;
      16009: inst = 32'd136314880;
      16010: inst = 32'd268468224;
      16011: inst = 32'd201346146;
      16012: inst = 32'd203484854;
      16013: inst = 32'd471859200;
      16014: inst = 32'd136314880;
      16015: inst = 32'd268468224;
      16016: inst = 32'd201346147;
      16017: inst = 32'd203484854;
      16018: inst = 32'd471859200;
      16019: inst = 32'd136314880;
      16020: inst = 32'd268468224;
      16021: inst = 32'd201346148;
      16022: inst = 32'd203484854;
      16023: inst = 32'd471859200;
      16024: inst = 32'd136314880;
      16025: inst = 32'd268468224;
      16026: inst = 32'd201346149;
      16027: inst = 32'd203484854;
      16028: inst = 32'd471859200;
      16029: inst = 32'd136314880;
      16030: inst = 32'd268468224;
      16031: inst = 32'd201346150;
      16032: inst = 32'd203484854;
      16033: inst = 32'd471859200;
      16034: inst = 32'd136314880;
      16035: inst = 32'd268468224;
      16036: inst = 32'd201346151;
      16037: inst = 32'd203484854;
      16038: inst = 32'd471859200;
      16039: inst = 32'd136314880;
      16040: inst = 32'd268468224;
      16041: inst = 32'd201346152;
      16042: inst = 32'd203484854;
      16043: inst = 32'd471859200;
      16044: inst = 32'd136314880;
      16045: inst = 32'd268468224;
      16046: inst = 32'd201346153;
      16047: inst = 32'd203484854;
      16048: inst = 32'd471859200;
      16049: inst = 32'd136314880;
      16050: inst = 32'd268468224;
      16051: inst = 32'd201346154;
      16052: inst = 32'd203484854;
      16053: inst = 32'd471859200;
      16054: inst = 32'd136314880;
      16055: inst = 32'd268468224;
      16056: inst = 32'd201346155;
      16057: inst = 32'd203484854;
      16058: inst = 32'd471859200;
      16059: inst = 32'd136314880;
      16060: inst = 32'd268468224;
      16061: inst = 32'd201346156;
      16062: inst = 32'd203484854;
      16063: inst = 32'd471859200;
      16064: inst = 32'd136314880;
      16065: inst = 32'd268468224;
      16066: inst = 32'd201346157;
      16067: inst = 32'd203484854;
      16068: inst = 32'd471859200;
      16069: inst = 32'd136314880;
      16070: inst = 32'd268468224;
      16071: inst = 32'd201346158;
      16072: inst = 32'd203484854;
      16073: inst = 32'd471859200;
      16074: inst = 32'd136314880;
      16075: inst = 32'd268468224;
      16076: inst = 32'd201346159;
      16077: inst = 32'd203484854;
      16078: inst = 32'd471859200;
      16079: inst = 32'd136314880;
      16080: inst = 32'd268468224;
      16081: inst = 32'd201346160;
      16082: inst = 32'd203484854;
      16083: inst = 32'd471859200;
      16084: inst = 32'd136314880;
      16085: inst = 32'd268468224;
      16086: inst = 32'd201346161;
      16087: inst = 32'd203484854;
      16088: inst = 32'd471859200;
      16089: inst = 32'd136314880;
      16090: inst = 32'd268468224;
      16091: inst = 32'd201346162;
      16092: inst = 32'd203484854;
      16093: inst = 32'd471859200;
      16094: inst = 32'd136314880;
      16095: inst = 32'd268468224;
      16096: inst = 32'd201346163;
      16097: inst = 32'd203484854;
      16098: inst = 32'd471859200;
      16099: inst = 32'd136314880;
      16100: inst = 32'd268468224;
      16101: inst = 32'd201346164;
      16102: inst = 32'd203484854;
      16103: inst = 32'd471859200;
      16104: inst = 32'd136314880;
      16105: inst = 32'd268468224;
      16106: inst = 32'd201346165;
      16107: inst = 32'd203484854;
      16108: inst = 32'd471859200;
      16109: inst = 32'd136314880;
      16110: inst = 32'd268468224;
      16111: inst = 32'd201346166;
      16112: inst = 32'd203484854;
      16113: inst = 32'd471859200;
      16114: inst = 32'd136314880;
      16115: inst = 32'd268468224;
      16116: inst = 32'd201346167;
      16117: inst = 32'd203484854;
      16118: inst = 32'd471859200;
      16119: inst = 32'd136314880;
      16120: inst = 32'd268468224;
      16121: inst = 32'd201346168;
      16122: inst = 32'd203484854;
      16123: inst = 32'd471859200;
      16124: inst = 32'd136314880;
      16125: inst = 32'd268468224;
      16126: inst = 32'd201346169;
      16127: inst = 32'd203484854;
      16128: inst = 32'd471859200;
      16129: inst = 32'd136314880;
      16130: inst = 32'd268468224;
      16131: inst = 32'd201346170;
      16132: inst = 32'd203484854;
      16133: inst = 32'd471859200;
      16134: inst = 32'd136314880;
      16135: inst = 32'd268468224;
      16136: inst = 32'd201346171;
      16137: inst = 32'd203484854;
      16138: inst = 32'd471859200;
      16139: inst = 32'd136314880;
      16140: inst = 32'd268468224;
      16141: inst = 32'd201346172;
      16142: inst = 32'd203484854;
      16143: inst = 32'd471859200;
      16144: inst = 32'd136314880;
      16145: inst = 32'd268468224;
      16146: inst = 32'd201346173;
      16147: inst = 32'd203484854;
      16148: inst = 32'd471859200;
      16149: inst = 32'd136314880;
      16150: inst = 32'd268468224;
      16151: inst = 32'd201346174;
      16152: inst = 32'd203484854;
      16153: inst = 32'd471859200;
      16154: inst = 32'd136314880;
      16155: inst = 32'd268468224;
      16156: inst = 32'd201346175;
      16157: inst = 32'd203484854;
      16158: inst = 32'd471859200;
      16159: inst = 32'd136314880;
      16160: inst = 32'd268468224;
      16161: inst = 32'd201346176;
      16162: inst = 32'd203484854;
      16163: inst = 32'd471859200;
      16164: inst = 32'd136314880;
      16165: inst = 32'd268468224;
      16166: inst = 32'd201346177;
      16167: inst = 32'd203484854;
      16168: inst = 32'd471859200;
      16169: inst = 32'd136314880;
      16170: inst = 32'd268468224;
      16171: inst = 32'd201346178;
      16172: inst = 32'd203484854;
      16173: inst = 32'd471859200;
      16174: inst = 32'd136314880;
      16175: inst = 32'd268468224;
      16176: inst = 32'd201346179;
      16177: inst = 32'd203484854;
      16178: inst = 32'd471859200;
      16179: inst = 32'd136314880;
      16180: inst = 32'd268468224;
      16181: inst = 32'd201346180;
      16182: inst = 32'd203484854;
      16183: inst = 32'd471859200;
      16184: inst = 32'd136314880;
      16185: inst = 32'd268468224;
      16186: inst = 32'd201346181;
      16187: inst = 32'd203484854;
      16188: inst = 32'd471859200;
      16189: inst = 32'd136314880;
      16190: inst = 32'd268468224;
      16191: inst = 32'd201346182;
      16192: inst = 32'd203484854;
      16193: inst = 32'd471859200;
      16194: inst = 32'd136314880;
      16195: inst = 32'd268468224;
      16196: inst = 32'd201346183;
      16197: inst = 32'd203484854;
      16198: inst = 32'd471859200;
      16199: inst = 32'd136314880;
      16200: inst = 32'd268468224;
      16201: inst = 32'd201346184;
      16202: inst = 32'd203484854;
      16203: inst = 32'd471859200;
      16204: inst = 32'd136314880;
      16205: inst = 32'd268468224;
      16206: inst = 32'd201346185;
      16207: inst = 32'd203484854;
      16208: inst = 32'd471859200;
      16209: inst = 32'd136314880;
      16210: inst = 32'd268468224;
      16211: inst = 32'd201346186;
      16212: inst = 32'd203484854;
      16213: inst = 32'd471859200;
      16214: inst = 32'd136314880;
      16215: inst = 32'd268468224;
      16216: inst = 32'd201346187;
      16217: inst = 32'd203484854;
      16218: inst = 32'd471859200;
      16219: inst = 32'd136314880;
      16220: inst = 32'd268468224;
      16221: inst = 32'd201346188;
      16222: inst = 32'd203484854;
      16223: inst = 32'd471859200;
      16224: inst = 32'd136314880;
      16225: inst = 32'd268468224;
      16226: inst = 32'd201346189;
      16227: inst = 32'd203484854;
      16228: inst = 32'd471859200;
      16229: inst = 32'd136314880;
      16230: inst = 32'd268468224;
      16231: inst = 32'd201346190;
      16232: inst = 32'd203484854;
      16233: inst = 32'd471859200;
      16234: inst = 32'd136314880;
      16235: inst = 32'd268468224;
      16236: inst = 32'd201346191;
      16237: inst = 32'd203473634;
      16238: inst = 32'd471859200;
      16239: inst = 32'd136314880;
      16240: inst = 32'd268468224;
      16241: inst = 32'd201346192;
      16242: inst = 32'd203480005;
      16243: inst = 32'd471859200;
      16244: inst = 32'd136314880;
      16245: inst = 32'd268468224;
      16246: inst = 32'd201346193;
      16247: inst = 32'd203480005;
      16248: inst = 32'd471859200;
      16249: inst = 32'd136314880;
      16250: inst = 32'd268468224;
      16251: inst = 32'd201346194;
      16252: inst = 32'd203480005;
      16253: inst = 32'd471859200;
      16254: inst = 32'd136314880;
      16255: inst = 32'd268468224;
      16256: inst = 32'd201346195;
      16257: inst = 32'd203480005;
      16258: inst = 32'd471859200;
      16259: inst = 32'd136314880;
      16260: inst = 32'd268468224;
      16261: inst = 32'd201346196;
      16262: inst = 32'd203480005;
      16263: inst = 32'd471859200;
      16264: inst = 32'd136314880;
      16265: inst = 32'd268468224;
      16266: inst = 32'd201346197;
      16267: inst = 32'd203480005;
      16268: inst = 32'd471859200;
      16269: inst = 32'd136314880;
      16270: inst = 32'd268468224;
      16271: inst = 32'd201346198;
      16272: inst = 32'd203480005;
      16273: inst = 32'd471859200;
      16274: inst = 32'd136314880;
      16275: inst = 32'd268468224;
      16276: inst = 32'd201346199;
      16277: inst = 32'd203480005;
      16278: inst = 32'd471859200;
      16279: inst = 32'd136314880;
      16280: inst = 32'd268468224;
      16281: inst = 32'd201346200;
      16282: inst = 32'd203480005;
      16283: inst = 32'd471859200;
      16284: inst = 32'd136314880;
      16285: inst = 32'd268468224;
      16286: inst = 32'd201346201;
      16287: inst = 32'd203480005;
      16288: inst = 32'd471859200;
      16289: inst = 32'd136314880;
      16290: inst = 32'd268468224;
      16291: inst = 32'd201346202;
      16292: inst = 32'd203480005;
      16293: inst = 32'd471859200;
      16294: inst = 32'd136314880;
      16295: inst = 32'd268468224;
      16296: inst = 32'd201346203;
      16297: inst = 32'd203480005;
      16298: inst = 32'd471859200;
      16299: inst = 32'd136314880;
      16300: inst = 32'd268468224;
      16301: inst = 32'd201346204;
      16302: inst = 32'd203480005;
      16303: inst = 32'd471859200;
      16304: inst = 32'd136314880;
      16305: inst = 32'd268468224;
      16306: inst = 32'd201346205;
      16307: inst = 32'd203480005;
      16308: inst = 32'd471859200;
      16309: inst = 32'd136314880;
      16310: inst = 32'd268468224;
      16311: inst = 32'd201346206;
      16312: inst = 32'd203480005;
      16313: inst = 32'd471859200;
      16314: inst = 32'd136314880;
      16315: inst = 32'd268468224;
      16316: inst = 32'd201346207;
      16317: inst = 32'd203473634;
      16318: inst = 32'd471859200;
      16319: inst = 32'd136314880;
      16320: inst = 32'd268468224;
      16321: inst = 32'd201346208;
      16322: inst = 32'd203484854;
      16323: inst = 32'd471859200;
      16324: inst = 32'd136314880;
      16325: inst = 32'd268468224;
      16326: inst = 32'd201346209;
      16327: inst = 32'd203484854;
      16328: inst = 32'd471859200;
      16329: inst = 32'd136314880;
      16330: inst = 32'd268468224;
      16331: inst = 32'd201346210;
      16332: inst = 32'd203478549;
      16333: inst = 32'd471859200;
      16334: inst = 32'd136314880;
      16335: inst = 32'd268468224;
      16336: inst = 32'd201346211;
      16337: inst = 32'd203463825;
      16338: inst = 32'd471859200;
      16339: inst = 32'd136314880;
      16340: inst = 32'd268468224;
      16341: inst = 32'd201346212;
      16342: inst = 32'd203455472;
      16343: inst = 32'd471859200;
      16344: inst = 32'd136314880;
      16345: inst = 32'd268468224;
      16346: inst = 32'd201346213;
      16347: inst = 32'd203455472;
      16348: inst = 32'd471859200;
      16349: inst = 32'd136314880;
      16350: inst = 32'd268468224;
      16351: inst = 32'd201346214;
      16352: inst = 32'd203455472;
      16353: inst = 32'd471859200;
      16354: inst = 32'd136314880;
      16355: inst = 32'd268468224;
      16356: inst = 32'd201346215;
      16357: inst = 32'd203455472;
      16358: inst = 32'd471859200;
      16359: inst = 32'd136314880;
      16360: inst = 32'd268468224;
      16361: inst = 32'd201346216;
      16362: inst = 32'd203442793;
      16363: inst = 32'd471859200;
      16364: inst = 32'd136314880;
      16365: inst = 32'd268468224;
      16366: inst = 32'd201346217;
      16367: inst = 32'd203480827;
      16368: inst = 32'd471859200;
      16369: inst = 32'd136314880;
      16370: inst = 32'd268468224;
      16371: inst = 32'd201346218;
      16372: inst = 32'd203442793;
      16373: inst = 32'd471859200;
      16374: inst = 32'd136314880;
      16375: inst = 32'd268468224;
      16376: inst = 32'd201346219;
      16377: inst = 32'd203480827;
      16378: inst = 32'd471859200;
      16379: inst = 32'd136314880;
      16380: inst = 32'd268468224;
      16381: inst = 32'd201346220;
      16382: inst = 32'd203442793;
      16383: inst = 32'd471859200;
      16384: inst = 32'd136314880;
      16385: inst = 32'd268468224;
      16386: inst = 32'd201346221;
      16387: inst = 32'd203468117;
      16388: inst = 32'd471859200;
      16389: inst = 32'd136314880;
      16390: inst = 32'd268468224;
      16391: inst = 32'd201346222;
      16392: inst = 32'd203457552;
      16393: inst = 32'd471859200;
      16394: inst = 32'd136314880;
      16395: inst = 32'd268468224;
      16396: inst = 32'd201346223;
      16397: inst = 32'd203457552;
      16398: inst = 32'd471859200;
      16399: inst = 32'd136314880;
      16400: inst = 32'd268468224;
      16401: inst = 32'd201346224;
      16402: inst = 32'd203457552;
      16403: inst = 32'd471859200;
      16404: inst = 32'd136314880;
      16405: inst = 32'd268468224;
      16406: inst = 32'd201346225;
      16407: inst = 32'd203457552;
      16408: inst = 32'd471859200;
      16409: inst = 32'd136314880;
      16410: inst = 32'd268468224;
      16411: inst = 32'd201346226;
      16412: inst = 32'd203457552;
      16413: inst = 32'd471859200;
      16414: inst = 32'd136314880;
      16415: inst = 32'd268468224;
      16416: inst = 32'd201346227;
      16417: inst = 32'd203457552;
      16418: inst = 32'd471859200;
      16419: inst = 32'd136314880;
      16420: inst = 32'd268468224;
      16421: inst = 32'd201346228;
      16422: inst = 32'd203457552;
      16423: inst = 32'd471859200;
      16424: inst = 32'd136314880;
      16425: inst = 32'd268468224;
      16426: inst = 32'd201346229;
      16427: inst = 32'd203457552;
      16428: inst = 32'd471859200;
      16429: inst = 32'd136314880;
      16430: inst = 32'd268468224;
      16431: inst = 32'd201346230;
      16432: inst = 32'd203461744;
      16433: inst = 32'd471859200;
      16434: inst = 32'd136314880;
      16435: inst = 32'd268468224;
      16436: inst = 32'd201346231;
      16437: inst = 32'd203484854;
      16438: inst = 32'd471859200;
      16439: inst = 32'd136314880;
      16440: inst = 32'd268468224;
      16441: inst = 32'd201346232;
      16442: inst = 32'd203484854;
      16443: inst = 32'd471859200;
      16444: inst = 32'd136314880;
      16445: inst = 32'd268468224;
      16446: inst = 32'd201346233;
      16447: inst = 32'd203484854;
      16448: inst = 32'd471859200;
      16449: inst = 32'd136314880;
      16450: inst = 32'd268468224;
      16451: inst = 32'd201346234;
      16452: inst = 32'd203484854;
      16453: inst = 32'd471859200;
      16454: inst = 32'd136314880;
      16455: inst = 32'd268468224;
      16456: inst = 32'd201346235;
      16457: inst = 32'd203484854;
      16458: inst = 32'd471859200;
      16459: inst = 32'd136314880;
      16460: inst = 32'd268468224;
      16461: inst = 32'd201346236;
      16462: inst = 32'd203484854;
      16463: inst = 32'd471859200;
      16464: inst = 32'd136314880;
      16465: inst = 32'd268468224;
      16466: inst = 32'd201346237;
      16467: inst = 32'd203484854;
      16468: inst = 32'd471859200;
      16469: inst = 32'd136314880;
      16470: inst = 32'd268468224;
      16471: inst = 32'd201346238;
      16472: inst = 32'd203484854;
      16473: inst = 32'd471859200;
      16474: inst = 32'd136314880;
      16475: inst = 32'd268468224;
      16476: inst = 32'd201346239;
      16477: inst = 32'd203484854;
      16478: inst = 32'd471859200;
      16479: inst = 32'd136314880;
      16480: inst = 32'd268468224;
      16481: inst = 32'd201346240;
      16482: inst = 32'd203484854;
      16483: inst = 32'd471859200;
      16484: inst = 32'd136314880;
      16485: inst = 32'd268468224;
      16486: inst = 32'd201346241;
      16487: inst = 32'd203484854;
      16488: inst = 32'd471859200;
      16489: inst = 32'd136314880;
      16490: inst = 32'd268468224;
      16491: inst = 32'd201346242;
      16492: inst = 32'd203484854;
      16493: inst = 32'd471859200;
      16494: inst = 32'd136314880;
      16495: inst = 32'd268468224;
      16496: inst = 32'd201346243;
      16497: inst = 32'd203484854;
      16498: inst = 32'd471859200;
      16499: inst = 32'd136314880;
      16500: inst = 32'd268468224;
      16501: inst = 32'd201346244;
      16502: inst = 32'd203484854;
      16503: inst = 32'd471859200;
      16504: inst = 32'd136314880;
      16505: inst = 32'd268468224;
      16506: inst = 32'd201346245;
      16507: inst = 32'd203484854;
      16508: inst = 32'd471859200;
      16509: inst = 32'd136314880;
      16510: inst = 32'd268468224;
      16511: inst = 32'd201346246;
      16512: inst = 32'd203484854;
      16513: inst = 32'd471859200;
      16514: inst = 32'd136314880;
      16515: inst = 32'd268468224;
      16516: inst = 32'd201346247;
      16517: inst = 32'd203484854;
      16518: inst = 32'd471859200;
      16519: inst = 32'd136314880;
      16520: inst = 32'd268468224;
      16521: inst = 32'd201346248;
      16522: inst = 32'd203484854;
      16523: inst = 32'd471859200;
      16524: inst = 32'd136314880;
      16525: inst = 32'd268468224;
      16526: inst = 32'd201346249;
      16527: inst = 32'd203484854;
      16528: inst = 32'd471859200;
      16529: inst = 32'd136314880;
      16530: inst = 32'd268468224;
      16531: inst = 32'd201346250;
      16532: inst = 32'd203484854;
      16533: inst = 32'd471859200;
      16534: inst = 32'd136314880;
      16535: inst = 32'd268468224;
      16536: inst = 32'd201346251;
      16537: inst = 32'd203484854;
      16538: inst = 32'd471859200;
      16539: inst = 32'd136314880;
      16540: inst = 32'd268468224;
      16541: inst = 32'd201346252;
      16542: inst = 32'd203484854;
      16543: inst = 32'd471859200;
      16544: inst = 32'd136314880;
      16545: inst = 32'd268468224;
      16546: inst = 32'd201346253;
      16547: inst = 32'd203484854;
      16548: inst = 32'd471859200;
      16549: inst = 32'd136314880;
      16550: inst = 32'd268468224;
      16551: inst = 32'd201346254;
      16552: inst = 32'd203484854;
      16553: inst = 32'd471859200;
      16554: inst = 32'd136314880;
      16555: inst = 32'd268468224;
      16556: inst = 32'd201346255;
      16557: inst = 32'd203484854;
      16558: inst = 32'd471859200;
      16559: inst = 32'd136314880;
      16560: inst = 32'd268468224;
      16561: inst = 32'd201346256;
      16562: inst = 32'd203484854;
      16563: inst = 32'd471859200;
      16564: inst = 32'd136314880;
      16565: inst = 32'd268468224;
      16566: inst = 32'd201346257;
      16567: inst = 32'd203484854;
      16568: inst = 32'd471859200;
      16569: inst = 32'd136314880;
      16570: inst = 32'd268468224;
      16571: inst = 32'd201346258;
      16572: inst = 32'd203484854;
      16573: inst = 32'd471859200;
      16574: inst = 32'd136314880;
      16575: inst = 32'd268468224;
      16576: inst = 32'd201346259;
      16577: inst = 32'd203484854;
      16578: inst = 32'd471859200;
      16579: inst = 32'd136314880;
      16580: inst = 32'd268468224;
      16581: inst = 32'd201346260;
      16582: inst = 32'd203484854;
      16583: inst = 32'd471859200;
      16584: inst = 32'd136314880;
      16585: inst = 32'd268468224;
      16586: inst = 32'd201346261;
      16587: inst = 32'd203484854;
      16588: inst = 32'd471859200;
      16589: inst = 32'd136314880;
      16590: inst = 32'd268468224;
      16591: inst = 32'd201346262;
      16592: inst = 32'd203484854;
      16593: inst = 32'd471859200;
      16594: inst = 32'd136314880;
      16595: inst = 32'd268468224;
      16596: inst = 32'd201346263;
      16597: inst = 32'd203484854;
      16598: inst = 32'd471859200;
      16599: inst = 32'd136314880;
      16600: inst = 32'd268468224;
      16601: inst = 32'd201346264;
      16602: inst = 32'd203484854;
      16603: inst = 32'd471859200;
      16604: inst = 32'd136314880;
      16605: inst = 32'd268468224;
      16606: inst = 32'd201346265;
      16607: inst = 32'd203484854;
      16608: inst = 32'd471859200;
      16609: inst = 32'd136314880;
      16610: inst = 32'd268468224;
      16611: inst = 32'd201346266;
      16612: inst = 32'd203484854;
      16613: inst = 32'd471859200;
      16614: inst = 32'd136314880;
      16615: inst = 32'd268468224;
      16616: inst = 32'd201346267;
      16617: inst = 32'd203484854;
      16618: inst = 32'd471859200;
      16619: inst = 32'd136314880;
      16620: inst = 32'd268468224;
      16621: inst = 32'd201346268;
      16622: inst = 32'd203484854;
      16623: inst = 32'd471859200;
      16624: inst = 32'd136314880;
      16625: inst = 32'd268468224;
      16626: inst = 32'd201346269;
      16627: inst = 32'd203484854;
      16628: inst = 32'd471859200;
      16629: inst = 32'd136314880;
      16630: inst = 32'd268468224;
      16631: inst = 32'd201346270;
      16632: inst = 32'd203484854;
      16633: inst = 32'd471859200;
      16634: inst = 32'd136314880;
      16635: inst = 32'd268468224;
      16636: inst = 32'd201346271;
      16637: inst = 32'd203484854;
      16638: inst = 32'd471859200;
      16639: inst = 32'd136314880;
      16640: inst = 32'd268468224;
      16641: inst = 32'd201346272;
      16642: inst = 32'd203484854;
      16643: inst = 32'd471859200;
      16644: inst = 32'd136314880;
      16645: inst = 32'd268468224;
      16646: inst = 32'd201346273;
      16647: inst = 32'd203484854;
      16648: inst = 32'd471859200;
      16649: inst = 32'd136314880;
      16650: inst = 32'd268468224;
      16651: inst = 32'd201346274;
      16652: inst = 32'd203484854;
      16653: inst = 32'd471859200;
      16654: inst = 32'd136314880;
      16655: inst = 32'd268468224;
      16656: inst = 32'd201346275;
      16657: inst = 32'd203484854;
      16658: inst = 32'd471859200;
      16659: inst = 32'd136314880;
      16660: inst = 32'd268468224;
      16661: inst = 32'd201346276;
      16662: inst = 32'd203484854;
      16663: inst = 32'd471859200;
      16664: inst = 32'd136314880;
      16665: inst = 32'd268468224;
      16666: inst = 32'd201346277;
      16667: inst = 32'd203484854;
      16668: inst = 32'd471859200;
      16669: inst = 32'd136314880;
      16670: inst = 32'd268468224;
      16671: inst = 32'd201346278;
      16672: inst = 32'd203484854;
      16673: inst = 32'd471859200;
      16674: inst = 32'd136314880;
      16675: inst = 32'd268468224;
      16676: inst = 32'd201346279;
      16677: inst = 32'd203484854;
      16678: inst = 32'd471859200;
      16679: inst = 32'd136314880;
      16680: inst = 32'd268468224;
      16681: inst = 32'd201346280;
      16682: inst = 32'd203484854;
      16683: inst = 32'd471859200;
      16684: inst = 32'd136314880;
      16685: inst = 32'd268468224;
      16686: inst = 32'd201346281;
      16687: inst = 32'd203484854;
      16688: inst = 32'd471859200;
      16689: inst = 32'd136314880;
      16690: inst = 32'd268468224;
      16691: inst = 32'd201346282;
      16692: inst = 32'd203484854;
      16693: inst = 32'd471859200;
      16694: inst = 32'd136314880;
      16695: inst = 32'd268468224;
      16696: inst = 32'd201346283;
      16697: inst = 32'd203484854;
      16698: inst = 32'd471859200;
      16699: inst = 32'd136314880;
      16700: inst = 32'd268468224;
      16701: inst = 32'd201346284;
      16702: inst = 32'd203484854;
      16703: inst = 32'd471859200;
      16704: inst = 32'd136314880;
      16705: inst = 32'd268468224;
      16706: inst = 32'd201346285;
      16707: inst = 32'd203484854;
      16708: inst = 32'd471859200;
      16709: inst = 32'd136314880;
      16710: inst = 32'd268468224;
      16711: inst = 32'd201346286;
      16712: inst = 32'd203484854;
      16713: inst = 32'd471859200;
      16714: inst = 32'd136314880;
      16715: inst = 32'd268468224;
      16716: inst = 32'd201346287;
      16717: inst = 32'd203473634;
      16718: inst = 32'd471859200;
      16719: inst = 32'd136314880;
      16720: inst = 32'd268468224;
      16721: inst = 32'd201346288;
      16722: inst = 32'd203480005;
      16723: inst = 32'd471859200;
      16724: inst = 32'd136314880;
      16725: inst = 32'd268468224;
      16726: inst = 32'd201346289;
      16727: inst = 32'd203480005;
      16728: inst = 32'd471859200;
      16729: inst = 32'd136314880;
      16730: inst = 32'd268468224;
      16731: inst = 32'd201346290;
      16732: inst = 32'd203480005;
      16733: inst = 32'd471859200;
      16734: inst = 32'd136314880;
      16735: inst = 32'd268468224;
      16736: inst = 32'd201346291;
      16737: inst = 32'd203480005;
      16738: inst = 32'd471859200;
      16739: inst = 32'd136314880;
      16740: inst = 32'd268468224;
      16741: inst = 32'd201346292;
      16742: inst = 32'd203480005;
      16743: inst = 32'd471859200;
      16744: inst = 32'd136314880;
      16745: inst = 32'd268468224;
      16746: inst = 32'd201346293;
      16747: inst = 32'd203480005;
      16748: inst = 32'd471859200;
      16749: inst = 32'd136314880;
      16750: inst = 32'd268468224;
      16751: inst = 32'd201346294;
      16752: inst = 32'd203480005;
      16753: inst = 32'd471859200;
      16754: inst = 32'd136314880;
      16755: inst = 32'd268468224;
      16756: inst = 32'd201346295;
      16757: inst = 32'd203480005;
      16758: inst = 32'd471859200;
      16759: inst = 32'd136314880;
      16760: inst = 32'd268468224;
      16761: inst = 32'd201346296;
      16762: inst = 32'd203480005;
      16763: inst = 32'd471859200;
      16764: inst = 32'd136314880;
      16765: inst = 32'd268468224;
      16766: inst = 32'd201346297;
      16767: inst = 32'd203480005;
      16768: inst = 32'd471859200;
      16769: inst = 32'd136314880;
      16770: inst = 32'd268468224;
      16771: inst = 32'd201346298;
      16772: inst = 32'd203480005;
      16773: inst = 32'd471859200;
      16774: inst = 32'd136314880;
      16775: inst = 32'd268468224;
      16776: inst = 32'd201346299;
      16777: inst = 32'd203466036;
      16778: inst = 32'd471859200;
      16779: inst = 32'd136314880;
      16780: inst = 32'd268468224;
      16781: inst = 32'd201346300;
      16782: inst = 32'd203459665;
      16783: inst = 32'd471859200;
      16784: inst = 32'd136314880;
      16785: inst = 32'd268468224;
      16786: inst = 32'd201346301;
      16787: inst = 32'd203459665;
      16788: inst = 32'd471859200;
      16789: inst = 32'd136314880;
      16790: inst = 32'd268468224;
      16791: inst = 32'd201346302;
      16792: inst = 32'd203480005;
      16793: inst = 32'd471859200;
      16794: inst = 32'd136314880;
      16795: inst = 32'd268468224;
      16796: inst = 32'd201346303;
      16797: inst = 32'd203473634;
      16798: inst = 32'd471859200;
      16799: inst = 32'd136314880;
      16800: inst = 32'd268468224;
      16801: inst = 32'd201346304;
      16802: inst = 32'd203478549;
      16803: inst = 32'd471859200;
      16804: inst = 32'd136314880;
      16805: inst = 32'd268468224;
      16806: inst = 32'd201346305;
      16807: inst = 32'd203463825;
      16808: inst = 32'd471859200;
      16809: inst = 32'd136314880;
      16810: inst = 32'd268468224;
      16811: inst = 32'd201346306;
      16812: inst = 32'd203455472;
      16813: inst = 32'd471859200;
      16814: inst = 32'd136314880;
      16815: inst = 32'd268468224;
      16816: inst = 32'd201346307;
      16817: inst = 32'd203455472;
      16818: inst = 32'd471859200;
      16819: inst = 32'd136314880;
      16820: inst = 32'd268468224;
      16821: inst = 32'd201346308;
      16822: inst = 32'd203455472;
      16823: inst = 32'd471859200;
      16824: inst = 32'd136314880;
      16825: inst = 32'd268468224;
      16826: inst = 32'd201346309;
      16827: inst = 32'd203455472;
      16828: inst = 32'd471859200;
      16829: inst = 32'd136314880;
      16830: inst = 32'd268468224;
      16831: inst = 32'd201346310;
      16832: inst = 32'd203455472;
      16833: inst = 32'd471859200;
      16834: inst = 32'd136314880;
      16835: inst = 32'd268468224;
      16836: inst = 32'd201346311;
      16837: inst = 32'd203455472;
      16838: inst = 32'd471859200;
      16839: inst = 32'd136314880;
      16840: inst = 32'd268468224;
      16841: inst = 32'd201346312;
      16842: inst = 32'd203455472;
      16843: inst = 32'd471859200;
      16844: inst = 32'd136314880;
      16845: inst = 32'd268468224;
      16846: inst = 32'd201346313;
      16847: inst = 32'd203455472;
      16848: inst = 32'd471859200;
      16849: inst = 32'd136314880;
      16850: inst = 32'd268468224;
      16851: inst = 32'd201346314;
      16852: inst = 32'd203455472;
      16853: inst = 32'd471859200;
      16854: inst = 32'd136314880;
      16855: inst = 32'd268468224;
      16856: inst = 32'd201346315;
      16857: inst = 32'd203455472;
      16858: inst = 32'd471859200;
      16859: inst = 32'd136314880;
      16860: inst = 32'd268468224;
      16861: inst = 32'd201346316;
      16862: inst = 32'd203455472;
      16863: inst = 32'd471859200;
      16864: inst = 32'd136314880;
      16865: inst = 32'd268468224;
      16866: inst = 32'd201346317;
      16867: inst = 32'd203455472;
      16868: inst = 32'd471859200;
      16869: inst = 32'd136314880;
      16870: inst = 32'd268468224;
      16871: inst = 32'd201346318;
      16872: inst = 32'd203455472;
      16873: inst = 32'd471859200;
      16874: inst = 32'd136314880;
      16875: inst = 32'd268468224;
      16876: inst = 32'd201346319;
      16877: inst = 32'd203455472;
      16878: inst = 32'd471859200;
      16879: inst = 32'd136314880;
      16880: inst = 32'd268468224;
      16881: inst = 32'd201346320;
      16882: inst = 32'd203455472;
      16883: inst = 32'd471859200;
      16884: inst = 32'd136314880;
      16885: inst = 32'd268468224;
      16886: inst = 32'd201346321;
      16887: inst = 32'd203455472;
      16888: inst = 32'd471859200;
      16889: inst = 32'd136314880;
      16890: inst = 32'd268468224;
      16891: inst = 32'd201346322;
      16892: inst = 32'd203455472;
      16893: inst = 32'd471859200;
      16894: inst = 32'd136314880;
      16895: inst = 32'd268468224;
      16896: inst = 32'd201346323;
      16897: inst = 32'd203455472;
      16898: inst = 32'd471859200;
      16899: inst = 32'd136314880;
      16900: inst = 32'd268468224;
      16901: inst = 32'd201346324;
      16902: inst = 32'd203455472;
      16903: inst = 32'd471859200;
      16904: inst = 32'd136314880;
      16905: inst = 32'd268468224;
      16906: inst = 32'd201346325;
      16907: inst = 32'd203461744;
      16908: inst = 32'd471859200;
      16909: inst = 32'd136314880;
      16910: inst = 32'd268468224;
      16911: inst = 32'd201346326;
      16912: inst = 32'd203451245;
      16913: inst = 32'd471859200;
      16914: inst = 32'd136314880;
      16915: inst = 32'd268468224;
      16916: inst = 32'd201346327;
      16917: inst = 32'd203484854;
      16918: inst = 32'd471859200;
      16919: inst = 32'd136314880;
      16920: inst = 32'd268468224;
      16921: inst = 32'd201346328;
      16922: inst = 32'd203484854;
      16923: inst = 32'd471859200;
      16924: inst = 32'd136314880;
      16925: inst = 32'd268468224;
      16926: inst = 32'd201346329;
      16927: inst = 32'd203484854;
      16928: inst = 32'd471859200;
      16929: inst = 32'd136314880;
      16930: inst = 32'd268468224;
      16931: inst = 32'd201346330;
      16932: inst = 32'd203484854;
      16933: inst = 32'd471859200;
      16934: inst = 32'd136314880;
      16935: inst = 32'd268468224;
      16936: inst = 32'd201346331;
      16937: inst = 32'd203484854;
      16938: inst = 32'd471859200;
      16939: inst = 32'd136314880;
      16940: inst = 32'd268468224;
      16941: inst = 32'd201346332;
      16942: inst = 32'd203484854;
      16943: inst = 32'd471859200;
      16944: inst = 32'd136314880;
      16945: inst = 32'd268468224;
      16946: inst = 32'd201346333;
      16947: inst = 32'd203484854;
      16948: inst = 32'd471859200;
      16949: inst = 32'd136314880;
      16950: inst = 32'd268468224;
      16951: inst = 32'd201346334;
      16952: inst = 32'd203484854;
      16953: inst = 32'd471859200;
      16954: inst = 32'd136314880;
      16955: inst = 32'd268468224;
      16956: inst = 32'd201346335;
      16957: inst = 32'd203484854;
      16958: inst = 32'd471859200;
      16959: inst = 32'd136314880;
      16960: inst = 32'd268468224;
      16961: inst = 32'd201346336;
      16962: inst = 32'd203484854;
      16963: inst = 32'd471859200;
      16964: inst = 32'd136314880;
      16965: inst = 32'd268468224;
      16966: inst = 32'd201346337;
      16967: inst = 32'd203484854;
      16968: inst = 32'd471859200;
      16969: inst = 32'd136314880;
      16970: inst = 32'd268468224;
      16971: inst = 32'd201346338;
      16972: inst = 32'd203484854;
      16973: inst = 32'd471859200;
      16974: inst = 32'd136314880;
      16975: inst = 32'd268468224;
      16976: inst = 32'd201346339;
      16977: inst = 32'd203484854;
      16978: inst = 32'd471859200;
      16979: inst = 32'd136314880;
      16980: inst = 32'd268468224;
      16981: inst = 32'd201346340;
      16982: inst = 32'd203484854;
      16983: inst = 32'd471859200;
      16984: inst = 32'd136314880;
      16985: inst = 32'd268468224;
      16986: inst = 32'd201346341;
      16987: inst = 32'd203484854;
      16988: inst = 32'd471859200;
      16989: inst = 32'd136314880;
      16990: inst = 32'd268468224;
      16991: inst = 32'd201346342;
      16992: inst = 32'd203484854;
      16993: inst = 32'd471859200;
      16994: inst = 32'd136314880;
      16995: inst = 32'd268468224;
      16996: inst = 32'd201346343;
      16997: inst = 32'd203484854;
      16998: inst = 32'd471859200;
      16999: inst = 32'd136314880;
      17000: inst = 32'd268468224;
      17001: inst = 32'd201346344;
      17002: inst = 32'd203484854;
      17003: inst = 32'd471859200;
      17004: inst = 32'd136314880;
      17005: inst = 32'd268468224;
      17006: inst = 32'd201346345;
      17007: inst = 32'd203484854;
      17008: inst = 32'd471859200;
      17009: inst = 32'd136314880;
      17010: inst = 32'd268468224;
      17011: inst = 32'd201346346;
      17012: inst = 32'd203484854;
      17013: inst = 32'd471859200;
      17014: inst = 32'd136314880;
      17015: inst = 32'd268468224;
      17016: inst = 32'd201346347;
      17017: inst = 32'd203484854;
      17018: inst = 32'd471859200;
      17019: inst = 32'd136314880;
      17020: inst = 32'd268468224;
      17021: inst = 32'd201346348;
      17022: inst = 32'd203484854;
      17023: inst = 32'd471859200;
      17024: inst = 32'd136314880;
      17025: inst = 32'd268468224;
      17026: inst = 32'd201346349;
      17027: inst = 32'd203484854;
      17028: inst = 32'd471859200;
      17029: inst = 32'd136314880;
      17030: inst = 32'd268468224;
      17031: inst = 32'd201346350;
      17032: inst = 32'd203484854;
      17033: inst = 32'd471859200;
      17034: inst = 32'd136314880;
      17035: inst = 32'd268468224;
      17036: inst = 32'd201346351;
      17037: inst = 32'd203484854;
      17038: inst = 32'd471859200;
      17039: inst = 32'd136314880;
      17040: inst = 32'd268468224;
      17041: inst = 32'd201346352;
      17042: inst = 32'd203484854;
      17043: inst = 32'd471859200;
      17044: inst = 32'd136314880;
      17045: inst = 32'd268468224;
      17046: inst = 32'd201346353;
      17047: inst = 32'd203484854;
      17048: inst = 32'd471859200;
      17049: inst = 32'd136314880;
      17050: inst = 32'd268468224;
      17051: inst = 32'd201346354;
      17052: inst = 32'd203484854;
      17053: inst = 32'd471859200;
      17054: inst = 32'd136314880;
      17055: inst = 32'd268468224;
      17056: inst = 32'd201346355;
      17057: inst = 32'd203484854;
      17058: inst = 32'd471859200;
      17059: inst = 32'd136314880;
      17060: inst = 32'd268468224;
      17061: inst = 32'd201346356;
      17062: inst = 32'd203484854;
      17063: inst = 32'd471859200;
      17064: inst = 32'd136314880;
      17065: inst = 32'd268468224;
      17066: inst = 32'd201346357;
      17067: inst = 32'd203484854;
      17068: inst = 32'd471859200;
      17069: inst = 32'd136314880;
      17070: inst = 32'd268468224;
      17071: inst = 32'd201346358;
      17072: inst = 32'd203484854;
      17073: inst = 32'd471859200;
      17074: inst = 32'd136314880;
      17075: inst = 32'd268468224;
      17076: inst = 32'd201346359;
      17077: inst = 32'd203484854;
      17078: inst = 32'd471859200;
      17079: inst = 32'd136314880;
      17080: inst = 32'd268468224;
      17081: inst = 32'd201346360;
      17082: inst = 32'd203484854;
      17083: inst = 32'd471859200;
      17084: inst = 32'd136314880;
      17085: inst = 32'd268468224;
      17086: inst = 32'd201346361;
      17087: inst = 32'd203484854;
      17088: inst = 32'd471859200;
      17089: inst = 32'd136314880;
      17090: inst = 32'd268468224;
      17091: inst = 32'd201346362;
      17092: inst = 32'd203484854;
      17093: inst = 32'd471859200;
      17094: inst = 32'd136314880;
      17095: inst = 32'd268468224;
      17096: inst = 32'd201346363;
      17097: inst = 32'd203484854;
      17098: inst = 32'd471859200;
      17099: inst = 32'd136314880;
      17100: inst = 32'd268468224;
      17101: inst = 32'd201346364;
      17102: inst = 32'd203484854;
      17103: inst = 32'd471859200;
      17104: inst = 32'd136314880;
      17105: inst = 32'd268468224;
      17106: inst = 32'd201346365;
      17107: inst = 32'd203484854;
      17108: inst = 32'd471859200;
      17109: inst = 32'd136314880;
      17110: inst = 32'd268468224;
      17111: inst = 32'd201346366;
      17112: inst = 32'd203484854;
      17113: inst = 32'd471859200;
      17114: inst = 32'd136314880;
      17115: inst = 32'd268468224;
      17116: inst = 32'd201346367;
      17117: inst = 32'd203484854;
      17118: inst = 32'd471859200;
      17119: inst = 32'd136314880;
      17120: inst = 32'd268468224;
      17121: inst = 32'd201346368;
      17122: inst = 32'd203484854;
      17123: inst = 32'd471859200;
      17124: inst = 32'd136314880;
      17125: inst = 32'd268468224;
      17126: inst = 32'd201346369;
      17127: inst = 32'd203484854;
      17128: inst = 32'd471859200;
      17129: inst = 32'd136314880;
      17130: inst = 32'd268468224;
      17131: inst = 32'd201346370;
      17132: inst = 32'd203484854;
      17133: inst = 32'd471859200;
      17134: inst = 32'd136314880;
      17135: inst = 32'd268468224;
      17136: inst = 32'd201346371;
      17137: inst = 32'd203484854;
      17138: inst = 32'd471859200;
      17139: inst = 32'd136314880;
      17140: inst = 32'd268468224;
      17141: inst = 32'd201346372;
      17142: inst = 32'd203484854;
      17143: inst = 32'd471859200;
      17144: inst = 32'd136314880;
      17145: inst = 32'd268468224;
      17146: inst = 32'd201346373;
      17147: inst = 32'd203484854;
      17148: inst = 32'd471859200;
      17149: inst = 32'd136314880;
      17150: inst = 32'd268468224;
      17151: inst = 32'd201346374;
      17152: inst = 32'd203484854;
      17153: inst = 32'd471859200;
      17154: inst = 32'd136314880;
      17155: inst = 32'd268468224;
      17156: inst = 32'd201346375;
      17157: inst = 32'd203484854;
      17158: inst = 32'd471859200;
      17159: inst = 32'd136314880;
      17160: inst = 32'd268468224;
      17161: inst = 32'd201346376;
      17162: inst = 32'd203484854;
      17163: inst = 32'd471859200;
      17164: inst = 32'd136314880;
      17165: inst = 32'd268468224;
      17166: inst = 32'd201346377;
      17167: inst = 32'd203484854;
      17168: inst = 32'd471859200;
      17169: inst = 32'd136314880;
      17170: inst = 32'd268468224;
      17171: inst = 32'd201346378;
      17172: inst = 32'd203484854;
      17173: inst = 32'd471859200;
      17174: inst = 32'd136314880;
      17175: inst = 32'd268468224;
      17176: inst = 32'd201346379;
      17177: inst = 32'd203484854;
      17178: inst = 32'd471859200;
      17179: inst = 32'd136314880;
      17180: inst = 32'd268468224;
      17181: inst = 32'd201346380;
      17182: inst = 32'd203484854;
      17183: inst = 32'd471859200;
      17184: inst = 32'd136314880;
      17185: inst = 32'd268468224;
      17186: inst = 32'd201346381;
      17187: inst = 32'd203484854;
      17188: inst = 32'd471859200;
      17189: inst = 32'd136314880;
      17190: inst = 32'd268468224;
      17191: inst = 32'd201346382;
      17192: inst = 32'd203484854;
      17193: inst = 32'd471859200;
      17194: inst = 32'd136314880;
      17195: inst = 32'd268468224;
      17196: inst = 32'd201346383;
      17197: inst = 32'd203473634;
      17198: inst = 32'd471859200;
      17199: inst = 32'd136314880;
      17200: inst = 32'd268468224;
      17201: inst = 32'd201346384;
      17202: inst = 32'd203480005;
      17203: inst = 32'd471859200;
      17204: inst = 32'd136314880;
      17205: inst = 32'd268468224;
      17206: inst = 32'd201346385;
      17207: inst = 32'd203480005;
      17208: inst = 32'd471859200;
      17209: inst = 32'd136314880;
      17210: inst = 32'd268468224;
      17211: inst = 32'd201346386;
      17212: inst = 32'd203480005;
      17213: inst = 32'd471859200;
      17214: inst = 32'd136314880;
      17215: inst = 32'd268468224;
      17216: inst = 32'd201346387;
      17217: inst = 32'd203480005;
      17218: inst = 32'd471859200;
      17219: inst = 32'd136314880;
      17220: inst = 32'd268468224;
      17221: inst = 32'd201346388;
      17222: inst = 32'd203480005;
      17223: inst = 32'd471859200;
      17224: inst = 32'd136314880;
      17225: inst = 32'd268468224;
      17226: inst = 32'd201346389;
      17227: inst = 32'd203480005;
      17228: inst = 32'd471859200;
      17229: inst = 32'd136314880;
      17230: inst = 32'd268468224;
      17231: inst = 32'd201346390;
      17232: inst = 32'd203480005;
      17233: inst = 32'd471859200;
      17234: inst = 32'd136314880;
      17235: inst = 32'd268468224;
      17236: inst = 32'd201346391;
      17237: inst = 32'd203480005;
      17238: inst = 32'd471859200;
      17239: inst = 32'd136314880;
      17240: inst = 32'd268468224;
      17241: inst = 32'd201346392;
      17242: inst = 32'd203480005;
      17243: inst = 32'd471859200;
      17244: inst = 32'd136314880;
      17245: inst = 32'd268468224;
      17246: inst = 32'd201346393;
      17247: inst = 32'd203480005;
      17248: inst = 32'd471859200;
      17249: inst = 32'd136314880;
      17250: inst = 32'd268468224;
      17251: inst = 32'd201346394;
      17252: inst = 32'd203480005;
      17253: inst = 32'd471859200;
      17254: inst = 32'd136314880;
      17255: inst = 32'd268468224;
      17256: inst = 32'd201346395;
      17257: inst = 32'd203474488;
      17258: inst = 32'd471859200;
      17259: inst = 32'd136314880;
      17260: inst = 32'd268468224;
      17261: inst = 32'd201346396;
      17262: inst = 32'd203480005;
      17263: inst = 32'd471859200;
      17264: inst = 32'd136314880;
      17265: inst = 32'd268468224;
      17266: inst = 32'd201346397;
      17267: inst = 32'd203480005;
      17268: inst = 32'd471859200;
      17269: inst = 32'd136314880;
      17270: inst = 32'd268468224;
      17271: inst = 32'd201346398;
      17272: inst = 32'd203480005;
      17273: inst = 32'd471859200;
      17274: inst = 32'd136314880;
      17275: inst = 32'd268468224;
      17276: inst = 32'd201346399;
      17277: inst = 32'd203473634;
      17278: inst = 32'd471859200;
      17279: inst = 32'd136314880;
      17280: inst = 32'd268468224;
      17281: inst = 32'd201346400;
      17282: inst = 32'd203459697;
      17283: inst = 32'd471859200;
      17284: inst = 32'd136314880;
      17285: inst = 32'd268468224;
      17286: inst = 32'd201346401;
      17287: inst = 32'd203459697;
      17288: inst = 32'd471859200;
      17289: inst = 32'd136314880;
      17290: inst = 32'd268468224;
      17291: inst = 32'd201346402;
      17292: inst = 32'd203459697;
      17293: inst = 32'd471859200;
      17294: inst = 32'd136314880;
      17295: inst = 32'd268468224;
      17296: inst = 32'd201346403;
      17297: inst = 32'd203459697;
      17298: inst = 32'd471859200;
      17299: inst = 32'd136314880;
      17300: inst = 32'd268468224;
      17301: inst = 32'd201346404;
      17302: inst = 32'd203459697;
      17303: inst = 32'd471859200;
      17304: inst = 32'd136314880;
      17305: inst = 32'd268468224;
      17306: inst = 32'd201346405;
      17307: inst = 32'd203459697;
      17308: inst = 32'd471859200;
      17309: inst = 32'd136314880;
      17310: inst = 32'd268468224;
      17311: inst = 32'd201346406;
      17312: inst = 32'd203459697;
      17313: inst = 32'd471859200;
      17314: inst = 32'd136314880;
      17315: inst = 32'd268468224;
      17316: inst = 32'd201346407;
      17317: inst = 32'd203459697;
      17318: inst = 32'd471859200;
      17319: inst = 32'd136314880;
      17320: inst = 32'd268468224;
      17321: inst = 32'd201346408;
      17322: inst = 32'd203459697;
      17323: inst = 32'd471859200;
      17324: inst = 32'd136314880;
      17325: inst = 32'd268468224;
      17326: inst = 32'd201346409;
      17327: inst = 32'd203459697;
      17328: inst = 32'd471859200;
      17329: inst = 32'd136314880;
      17330: inst = 32'd268468224;
      17331: inst = 32'd201346410;
      17332: inst = 32'd203459697;
      17333: inst = 32'd471859200;
      17334: inst = 32'd136314880;
      17335: inst = 32'd268468224;
      17336: inst = 32'd201346411;
      17337: inst = 32'd203459697;
      17338: inst = 32'd471859200;
      17339: inst = 32'd136314880;
      17340: inst = 32'd268468224;
      17341: inst = 32'd201346412;
      17342: inst = 32'd203459697;
      17343: inst = 32'd471859200;
      17344: inst = 32'd136314880;
      17345: inst = 32'd268468224;
      17346: inst = 32'd201346413;
      17347: inst = 32'd203459697;
      17348: inst = 32'd471859200;
      17349: inst = 32'd136314880;
      17350: inst = 32'd268468224;
      17351: inst = 32'd201346414;
      17352: inst = 32'd203459697;
      17353: inst = 32'd471859200;
      17354: inst = 32'd136314880;
      17355: inst = 32'd268468224;
      17356: inst = 32'd201346415;
      17357: inst = 32'd203459697;
      17358: inst = 32'd471859200;
      17359: inst = 32'd136314880;
      17360: inst = 32'd268468224;
      17361: inst = 32'd201346416;
      17362: inst = 32'd203459697;
      17363: inst = 32'd471859200;
      17364: inst = 32'd136314880;
      17365: inst = 32'd268468224;
      17366: inst = 32'd201346417;
      17367: inst = 32'd203459697;
      17368: inst = 32'd471859200;
      17369: inst = 32'd136314880;
      17370: inst = 32'd268468224;
      17371: inst = 32'd201346418;
      17372: inst = 32'd203459697;
      17373: inst = 32'd471859200;
      17374: inst = 32'd136314880;
      17375: inst = 32'd268468224;
      17376: inst = 32'd201346419;
      17377: inst = 32'd203459697;
      17378: inst = 32'd471859200;
      17379: inst = 32'd136314880;
      17380: inst = 32'd268468224;
      17381: inst = 32'd201346420;
      17382: inst = 32'd203459697;
      17383: inst = 32'd471859200;
      17384: inst = 32'd136314880;
      17385: inst = 32'd268468224;
      17386: inst = 32'd201346421;
      17387: inst = 32'd203451245;
      17388: inst = 32'd471859200;
      17389: inst = 32'd136314880;
      17390: inst = 32'd268468224;
      17391: inst = 32'd201346422;
      17392: inst = 32'd203451245;
      17393: inst = 32'd471859200;
      17394: inst = 32'd136314880;
      17395: inst = 32'd268468224;
      17396: inst = 32'd201346423;
      17397: inst = 32'd203484854;
      17398: inst = 32'd471859200;
      17399: inst = 32'd136314880;
      17400: inst = 32'd268468224;
      17401: inst = 32'd201346424;
      17402: inst = 32'd203484854;
      17403: inst = 32'd471859200;
      17404: inst = 32'd136314880;
      17405: inst = 32'd268468224;
      17406: inst = 32'd201346425;
      17407: inst = 32'd203484854;
      17408: inst = 32'd471859200;
      17409: inst = 32'd136314880;
      17410: inst = 32'd268468224;
      17411: inst = 32'd201346426;
      17412: inst = 32'd203484854;
      17413: inst = 32'd471859200;
      17414: inst = 32'd136314880;
      17415: inst = 32'd268468224;
      17416: inst = 32'd201346427;
      17417: inst = 32'd203484854;
      17418: inst = 32'd471859200;
      17419: inst = 32'd136314880;
      17420: inst = 32'd268468224;
      17421: inst = 32'd201346428;
      17422: inst = 32'd203484854;
      17423: inst = 32'd471859200;
      17424: inst = 32'd136314880;
      17425: inst = 32'd268468224;
      17426: inst = 32'd201346429;
      17427: inst = 32'd203484854;
      17428: inst = 32'd471859200;
      17429: inst = 32'd136314880;
      17430: inst = 32'd268468224;
      17431: inst = 32'd201346430;
      17432: inst = 32'd203484854;
      17433: inst = 32'd471859200;
      17434: inst = 32'd136314880;
      17435: inst = 32'd268468224;
      17436: inst = 32'd201346431;
      17437: inst = 32'd203484854;
      17438: inst = 32'd471859200;
      17439: inst = 32'd136314880;
      17440: inst = 32'd268468224;
      17441: inst = 32'd201346432;
      17442: inst = 32'd203484854;
      17443: inst = 32'd471859200;
      17444: inst = 32'd136314880;
      17445: inst = 32'd268468224;
      17446: inst = 32'd201346433;
      17447: inst = 32'd203484854;
      17448: inst = 32'd471859200;
      17449: inst = 32'd136314880;
      17450: inst = 32'd268468224;
      17451: inst = 32'd201346434;
      17452: inst = 32'd203484854;
      17453: inst = 32'd471859200;
      17454: inst = 32'd136314880;
      17455: inst = 32'd268468224;
      17456: inst = 32'd201346435;
      17457: inst = 32'd203484854;
      17458: inst = 32'd471859200;
      17459: inst = 32'd136314880;
      17460: inst = 32'd268468224;
      17461: inst = 32'd201346436;
      17462: inst = 32'd203484854;
      17463: inst = 32'd471859200;
      17464: inst = 32'd136314880;
      17465: inst = 32'd268468224;
      17466: inst = 32'd201346437;
      17467: inst = 32'd203484854;
      17468: inst = 32'd471859200;
      17469: inst = 32'd136314880;
      17470: inst = 32'd268468224;
      17471: inst = 32'd201346438;
      17472: inst = 32'd203484854;
      17473: inst = 32'd471859200;
      17474: inst = 32'd136314880;
      17475: inst = 32'd268468224;
      17476: inst = 32'd201346439;
      17477: inst = 32'd203484854;
      17478: inst = 32'd471859200;
      17479: inst = 32'd136314880;
      17480: inst = 32'd268468224;
      17481: inst = 32'd201346440;
      17482: inst = 32'd203484854;
      17483: inst = 32'd471859200;
      17484: inst = 32'd136314880;
      17485: inst = 32'd268468224;
      17486: inst = 32'd201346441;
      17487: inst = 32'd203484854;
      17488: inst = 32'd471859200;
      17489: inst = 32'd136314880;
      17490: inst = 32'd268468224;
      17491: inst = 32'd201346442;
      17492: inst = 32'd203484854;
      17493: inst = 32'd471859200;
      17494: inst = 32'd136314880;
      17495: inst = 32'd268468224;
      17496: inst = 32'd201346443;
      17497: inst = 32'd203484854;
      17498: inst = 32'd471859200;
      17499: inst = 32'd136314880;
      17500: inst = 32'd268468224;
      17501: inst = 32'd201346444;
      17502: inst = 32'd203484854;
      17503: inst = 32'd471859200;
      17504: inst = 32'd136314880;
      17505: inst = 32'd268468224;
      17506: inst = 32'd201346445;
      17507: inst = 32'd203484854;
      17508: inst = 32'd471859200;
      17509: inst = 32'd136314880;
      17510: inst = 32'd268468224;
      17511: inst = 32'd201346446;
      17512: inst = 32'd203484854;
      17513: inst = 32'd471859200;
      17514: inst = 32'd136314880;
      17515: inst = 32'd268468224;
      17516: inst = 32'd201346447;
      17517: inst = 32'd203484854;
      17518: inst = 32'd471859200;
      17519: inst = 32'd136314880;
      17520: inst = 32'd268468224;
      17521: inst = 32'd201346448;
      17522: inst = 32'd203484854;
      17523: inst = 32'd471859200;
      17524: inst = 32'd136314880;
      17525: inst = 32'd268468224;
      17526: inst = 32'd201346449;
      17527: inst = 32'd203484854;
      17528: inst = 32'd471859200;
      17529: inst = 32'd136314880;
      17530: inst = 32'd268468224;
      17531: inst = 32'd201346450;
      17532: inst = 32'd203484854;
      17533: inst = 32'd471859200;
      17534: inst = 32'd136314880;
      17535: inst = 32'd268468224;
      17536: inst = 32'd201346451;
      17537: inst = 32'd203484854;
      17538: inst = 32'd471859200;
      17539: inst = 32'd136314880;
      17540: inst = 32'd268468224;
      17541: inst = 32'd201346452;
      17542: inst = 32'd203484854;
      17543: inst = 32'd471859200;
      17544: inst = 32'd136314880;
      17545: inst = 32'd268468224;
      17546: inst = 32'd201346453;
      17547: inst = 32'd203484854;
      17548: inst = 32'd471859200;
      17549: inst = 32'd136314880;
      17550: inst = 32'd268468224;
      17551: inst = 32'd201346454;
      17552: inst = 32'd203484854;
      17553: inst = 32'd471859200;
      17554: inst = 32'd136314880;
      17555: inst = 32'd268468224;
      17556: inst = 32'd201346455;
      17557: inst = 32'd203484854;
      17558: inst = 32'd471859200;
      17559: inst = 32'd136314880;
      17560: inst = 32'd268468224;
      17561: inst = 32'd201346456;
      17562: inst = 32'd203484854;
      17563: inst = 32'd471859200;
      17564: inst = 32'd136314880;
      17565: inst = 32'd268468224;
      17566: inst = 32'd201346457;
      17567: inst = 32'd203484854;
      17568: inst = 32'd471859200;
      17569: inst = 32'd136314880;
      17570: inst = 32'd268468224;
      17571: inst = 32'd201346458;
      17572: inst = 32'd203484854;
      17573: inst = 32'd471859200;
      17574: inst = 32'd136314880;
      17575: inst = 32'd268468224;
      17576: inst = 32'd201346459;
      17577: inst = 32'd203484854;
      17578: inst = 32'd471859200;
      17579: inst = 32'd136314880;
      17580: inst = 32'd268468224;
      17581: inst = 32'd201346460;
      17582: inst = 32'd203484854;
      17583: inst = 32'd471859200;
      17584: inst = 32'd136314880;
      17585: inst = 32'd268468224;
      17586: inst = 32'd201346461;
      17587: inst = 32'd203484854;
      17588: inst = 32'd471859200;
      17589: inst = 32'd136314880;
      17590: inst = 32'd268468224;
      17591: inst = 32'd201346462;
      17592: inst = 32'd203484854;
      17593: inst = 32'd471859200;
      17594: inst = 32'd136314880;
      17595: inst = 32'd268468224;
      17596: inst = 32'd201346463;
      17597: inst = 32'd203484854;
      17598: inst = 32'd471859200;
      17599: inst = 32'd136314880;
      17600: inst = 32'd268468224;
      17601: inst = 32'd201346464;
      17602: inst = 32'd203484854;
      17603: inst = 32'd471859200;
      17604: inst = 32'd136314880;
      17605: inst = 32'd268468224;
      17606: inst = 32'd201346465;
      17607: inst = 32'd203484854;
      17608: inst = 32'd471859200;
      17609: inst = 32'd136314880;
      17610: inst = 32'd268468224;
      17611: inst = 32'd201346466;
      17612: inst = 32'd203484854;
      17613: inst = 32'd471859200;
      17614: inst = 32'd136314880;
      17615: inst = 32'd268468224;
      17616: inst = 32'd201346467;
      17617: inst = 32'd203484854;
      17618: inst = 32'd471859200;
      17619: inst = 32'd136314880;
      17620: inst = 32'd268468224;
      17621: inst = 32'd201346468;
      17622: inst = 32'd203484854;
      17623: inst = 32'd471859200;
      17624: inst = 32'd136314880;
      17625: inst = 32'd268468224;
      17626: inst = 32'd201346469;
      17627: inst = 32'd203484854;
      17628: inst = 32'd471859200;
      17629: inst = 32'd136314880;
      17630: inst = 32'd268468224;
      17631: inst = 32'd201346470;
      17632: inst = 32'd203484854;
      17633: inst = 32'd471859200;
      17634: inst = 32'd136314880;
      17635: inst = 32'd268468224;
      17636: inst = 32'd201346471;
      17637: inst = 32'd203484854;
      17638: inst = 32'd471859200;
      17639: inst = 32'd136314880;
      17640: inst = 32'd268468224;
      17641: inst = 32'd201346472;
      17642: inst = 32'd203484854;
      17643: inst = 32'd471859200;
      17644: inst = 32'd136314880;
      17645: inst = 32'd268468224;
      17646: inst = 32'd201346473;
      17647: inst = 32'd203484854;
      17648: inst = 32'd471859200;
      17649: inst = 32'd136314880;
      17650: inst = 32'd268468224;
      17651: inst = 32'd201346474;
      17652: inst = 32'd203484854;
      17653: inst = 32'd471859200;
      17654: inst = 32'd136314880;
      17655: inst = 32'd268468224;
      17656: inst = 32'd201346475;
      17657: inst = 32'd203484854;
      17658: inst = 32'd471859200;
      17659: inst = 32'd136314880;
      17660: inst = 32'd268468224;
      17661: inst = 32'd201346476;
      17662: inst = 32'd203484854;
      17663: inst = 32'd471859200;
      17664: inst = 32'd136314880;
      17665: inst = 32'd268468224;
      17666: inst = 32'd201346477;
      17667: inst = 32'd203484854;
      17668: inst = 32'd471859200;
      17669: inst = 32'd136314880;
      17670: inst = 32'd268468224;
      17671: inst = 32'd201346478;
      17672: inst = 32'd203484854;
      17673: inst = 32'd471859200;
      17674: inst = 32'd136314880;
      17675: inst = 32'd268468224;
      17676: inst = 32'd201346479;
      17677: inst = 32'd203473634;
      17678: inst = 32'd471859200;
      17679: inst = 32'd136314880;
      17680: inst = 32'd268468224;
      17681: inst = 32'd201346480;
      17682: inst = 32'd203480005;
      17683: inst = 32'd471859200;
      17684: inst = 32'd136314880;
      17685: inst = 32'd268468224;
      17686: inst = 32'd201346481;
      17687: inst = 32'd203480005;
      17688: inst = 32'd471859200;
      17689: inst = 32'd136314880;
      17690: inst = 32'd268468224;
      17691: inst = 32'd201346482;
      17692: inst = 32'd203480005;
      17693: inst = 32'd471859200;
      17694: inst = 32'd136314880;
      17695: inst = 32'd268468224;
      17696: inst = 32'd201346483;
      17697: inst = 32'd203480005;
      17698: inst = 32'd471859200;
      17699: inst = 32'd136314880;
      17700: inst = 32'd268468224;
      17701: inst = 32'd201346484;
      17702: inst = 32'd203480005;
      17703: inst = 32'd471859200;
      17704: inst = 32'd136314880;
      17705: inst = 32'd268468224;
      17706: inst = 32'd201346485;
      17707: inst = 32'd203480005;
      17708: inst = 32'd471859200;
      17709: inst = 32'd136314880;
      17710: inst = 32'd268468224;
      17711: inst = 32'd201346486;
      17712: inst = 32'd203480005;
      17713: inst = 32'd471859200;
      17714: inst = 32'd136314880;
      17715: inst = 32'd268468224;
      17716: inst = 32'd201346487;
      17717: inst = 32'd203480005;
      17718: inst = 32'd471859200;
      17719: inst = 32'd136314880;
      17720: inst = 32'd268468224;
      17721: inst = 32'd201346488;
      17722: inst = 32'd203480005;
      17723: inst = 32'd471859200;
      17724: inst = 32'd136314880;
      17725: inst = 32'd268468224;
      17726: inst = 32'd201346489;
      17727: inst = 32'd203480005;
      17728: inst = 32'd471859200;
      17729: inst = 32'd136314880;
      17730: inst = 32'd268468224;
      17731: inst = 32'd201346490;
      17732: inst = 32'd203480005;
      17733: inst = 32'd471859200;
      17734: inst = 32'd136314880;
      17735: inst = 32'd268468224;
      17736: inst = 32'd201346491;
      17737: inst = 32'd203480005;
      17738: inst = 32'd471859200;
      17739: inst = 32'd136314880;
      17740: inst = 32'd268468224;
      17741: inst = 32'd201346492;
      17742: inst = 32'd203480005;
      17743: inst = 32'd471859200;
      17744: inst = 32'd136314880;
      17745: inst = 32'd268468224;
      17746: inst = 32'd201346493;
      17747: inst = 32'd203480005;
      17748: inst = 32'd471859200;
      17749: inst = 32'd136314880;
      17750: inst = 32'd268468224;
      17751: inst = 32'd201346494;
      17752: inst = 32'd203480005;
      17753: inst = 32'd471859200;
      17754: inst = 32'd136314880;
      17755: inst = 32'd268468224;
      17756: inst = 32'd201346495;
      17757: inst = 32'd203473634;
      17758: inst = 32'd471859200;
      17759: inst = 32'd136314880;
      17760: inst = 32'd268468224;
      17761: inst = 32'd201346496;
      17762: inst = 32'd203459697;
      17763: inst = 32'd471859200;
      17764: inst = 32'd136314880;
      17765: inst = 32'd268468224;
      17766: inst = 32'd201346497;
      17767: inst = 32'd203472343;
      17768: inst = 32'd471859200;
      17769: inst = 32'd136314880;
      17770: inst = 32'd268468224;
      17771: inst = 32'd201346498;
      17772: inst = 32'd203472343;
      17773: inst = 32'd471859200;
      17774: inst = 32'd136314880;
      17775: inst = 32'd268468224;
      17776: inst = 32'd201346499;
      17777: inst = 32'd203472343;
      17778: inst = 32'd471859200;
      17779: inst = 32'd136314880;
      17780: inst = 32'd268468224;
      17781: inst = 32'd201346500;
      17782: inst = 32'd203472343;
      17783: inst = 32'd471859200;
      17784: inst = 32'd136314880;
      17785: inst = 32'd268468224;
      17786: inst = 32'd201346501;
      17787: inst = 32'd203472343;
      17788: inst = 32'd471859200;
      17789: inst = 32'd136314880;
      17790: inst = 32'd268468224;
      17791: inst = 32'd201346502;
      17792: inst = 32'd203472343;
      17793: inst = 32'd471859200;
      17794: inst = 32'd136314880;
      17795: inst = 32'd268468224;
      17796: inst = 32'd201346503;
      17797: inst = 32'd203472343;
      17798: inst = 32'd471859200;
      17799: inst = 32'd136314880;
      17800: inst = 32'd268468224;
      17801: inst = 32'd201346504;
      17802: inst = 32'd203472343;
      17803: inst = 32'd471859200;
      17804: inst = 32'd136314880;
      17805: inst = 32'd268468224;
      17806: inst = 32'd201346505;
      17807: inst = 32'd203472343;
      17808: inst = 32'd471859200;
      17809: inst = 32'd136314880;
      17810: inst = 32'd268468224;
      17811: inst = 32'd201346506;
      17812: inst = 32'd203459697;
      17813: inst = 32'd471859200;
      17814: inst = 32'd136314880;
      17815: inst = 32'd268468224;
      17816: inst = 32'd201346507;
      17817: inst = 32'd203472343;
      17818: inst = 32'd471859200;
      17819: inst = 32'd136314880;
      17820: inst = 32'd268468224;
      17821: inst = 32'd201346508;
      17822: inst = 32'd203472343;
      17823: inst = 32'd471859200;
      17824: inst = 32'd136314880;
      17825: inst = 32'd268468224;
      17826: inst = 32'd201346509;
      17827: inst = 32'd203472343;
      17828: inst = 32'd471859200;
      17829: inst = 32'd136314880;
      17830: inst = 32'd268468224;
      17831: inst = 32'd201346510;
      17832: inst = 32'd203472343;
      17833: inst = 32'd471859200;
      17834: inst = 32'd136314880;
      17835: inst = 32'd268468224;
      17836: inst = 32'd201346511;
      17837: inst = 32'd203472343;
      17838: inst = 32'd471859200;
      17839: inst = 32'd136314880;
      17840: inst = 32'd268468224;
      17841: inst = 32'd201346512;
      17842: inst = 32'd203472343;
      17843: inst = 32'd471859200;
      17844: inst = 32'd136314880;
      17845: inst = 32'd268468224;
      17846: inst = 32'd201346513;
      17847: inst = 32'd203472343;
      17848: inst = 32'd471859200;
      17849: inst = 32'd136314880;
      17850: inst = 32'd268468224;
      17851: inst = 32'd201346514;
      17852: inst = 32'd203472343;
      17853: inst = 32'd471859200;
      17854: inst = 32'd136314880;
      17855: inst = 32'd268468224;
      17856: inst = 32'd201346515;
      17857: inst = 32'd203472343;
      17858: inst = 32'd471859200;
      17859: inst = 32'd136314880;
      17860: inst = 32'd268468224;
      17861: inst = 32'd201346516;
      17862: inst = 32'd203459697;
      17863: inst = 32'd471859200;
      17864: inst = 32'd136314880;
      17865: inst = 32'd268468224;
      17866: inst = 32'd201346517;
      17867: inst = 32'd203451245;
      17868: inst = 32'd471859200;
      17869: inst = 32'd136314880;
      17870: inst = 32'd268468224;
      17871: inst = 32'd201346518;
      17872: inst = 32'd203451245;
      17873: inst = 32'd471859200;
      17874: inst = 32'd136314880;
      17875: inst = 32'd268468224;
      17876: inst = 32'd201346519;
      17877: inst = 32'd203484854;
      17878: inst = 32'd471859200;
      17879: inst = 32'd136314880;
      17880: inst = 32'd268468224;
      17881: inst = 32'd201346520;
      17882: inst = 32'd203484854;
      17883: inst = 32'd471859200;
      17884: inst = 32'd136314880;
      17885: inst = 32'd268468224;
      17886: inst = 32'd201346521;
      17887: inst = 32'd203484854;
      17888: inst = 32'd471859200;
      17889: inst = 32'd136314880;
      17890: inst = 32'd268468224;
      17891: inst = 32'd201346522;
      17892: inst = 32'd203484854;
      17893: inst = 32'd471859200;
      17894: inst = 32'd136314880;
      17895: inst = 32'd268468224;
      17896: inst = 32'd201346523;
      17897: inst = 32'd203484854;
      17898: inst = 32'd471859200;
      17899: inst = 32'd136314880;
      17900: inst = 32'd268468224;
      17901: inst = 32'd201346524;
      17902: inst = 32'd203484854;
      17903: inst = 32'd471859200;
      17904: inst = 32'd136314880;
      17905: inst = 32'd268468224;
      17906: inst = 32'd201346525;
      17907: inst = 32'd203484854;
      17908: inst = 32'd471859200;
      17909: inst = 32'd136314880;
      17910: inst = 32'd268468224;
      17911: inst = 32'd201346526;
      17912: inst = 32'd203484854;
      17913: inst = 32'd471859200;
      17914: inst = 32'd136314880;
      17915: inst = 32'd268468224;
      17916: inst = 32'd201346527;
      17917: inst = 32'd203484854;
      17918: inst = 32'd471859200;
      17919: inst = 32'd136314880;
      17920: inst = 32'd268468224;
      17921: inst = 32'd201346528;
      17922: inst = 32'd203484854;
      17923: inst = 32'd471859200;
      17924: inst = 32'd136314880;
      17925: inst = 32'd268468224;
      17926: inst = 32'd201346529;
      17927: inst = 32'd203484854;
      17928: inst = 32'd471859200;
      17929: inst = 32'd136314880;
      17930: inst = 32'd268468224;
      17931: inst = 32'd201346530;
      17932: inst = 32'd203484854;
      17933: inst = 32'd471859200;
      17934: inst = 32'd136314880;
      17935: inst = 32'd268468224;
      17936: inst = 32'd201346531;
      17937: inst = 32'd203484854;
      17938: inst = 32'd471859200;
      17939: inst = 32'd136314880;
      17940: inst = 32'd268468224;
      17941: inst = 32'd201346532;
      17942: inst = 32'd203484854;
      17943: inst = 32'd471859200;
      17944: inst = 32'd136314880;
      17945: inst = 32'd268468224;
      17946: inst = 32'd201346533;
      17947: inst = 32'd203484854;
      17948: inst = 32'd471859200;
      17949: inst = 32'd136314880;
      17950: inst = 32'd268468224;
      17951: inst = 32'd201346534;
      17952: inst = 32'd203484854;
      17953: inst = 32'd471859200;
      17954: inst = 32'd136314880;
      17955: inst = 32'd268468224;
      17956: inst = 32'd201346535;
      17957: inst = 32'd203484854;
      17958: inst = 32'd471859200;
      17959: inst = 32'd136314880;
      17960: inst = 32'd268468224;
      17961: inst = 32'd201346536;
      17962: inst = 32'd203484854;
      17963: inst = 32'd471859200;
      17964: inst = 32'd136314880;
      17965: inst = 32'd268468224;
      17966: inst = 32'd201346537;
      17967: inst = 32'd203484854;
      17968: inst = 32'd471859200;
      17969: inst = 32'd136314880;
      17970: inst = 32'd268468224;
      17971: inst = 32'd201346538;
      17972: inst = 32'd203484854;
      17973: inst = 32'd471859200;
      17974: inst = 32'd136314880;
      17975: inst = 32'd268468224;
      17976: inst = 32'd201346539;
      17977: inst = 32'd203484854;
      17978: inst = 32'd471859200;
      17979: inst = 32'd136314880;
      17980: inst = 32'd268468224;
      17981: inst = 32'd201346540;
      17982: inst = 32'd203484854;
      17983: inst = 32'd471859200;
      17984: inst = 32'd136314880;
      17985: inst = 32'd268468224;
      17986: inst = 32'd201346541;
      17987: inst = 32'd203484854;
      17988: inst = 32'd471859200;
      17989: inst = 32'd136314880;
      17990: inst = 32'd268468224;
      17991: inst = 32'd201346542;
      17992: inst = 32'd203484854;
      17993: inst = 32'd471859200;
      17994: inst = 32'd136314880;
      17995: inst = 32'd268468224;
      17996: inst = 32'd201346543;
      17997: inst = 32'd203484854;
      17998: inst = 32'd471859200;
      17999: inst = 32'd136314880;
      18000: inst = 32'd268468224;
      18001: inst = 32'd201346544;
      18002: inst = 32'd203484854;
      18003: inst = 32'd471859200;
      18004: inst = 32'd136314880;
      18005: inst = 32'd268468224;
      18006: inst = 32'd201346545;
      18007: inst = 32'd203484854;
      18008: inst = 32'd471859200;
      18009: inst = 32'd136314880;
      18010: inst = 32'd268468224;
      18011: inst = 32'd201346546;
      18012: inst = 32'd203484854;
      18013: inst = 32'd471859200;
      18014: inst = 32'd136314880;
      18015: inst = 32'd268468224;
      18016: inst = 32'd201346547;
      18017: inst = 32'd203484854;
      18018: inst = 32'd471859200;
      18019: inst = 32'd136314880;
      18020: inst = 32'd268468224;
      18021: inst = 32'd201346548;
      18022: inst = 32'd203484854;
      18023: inst = 32'd471859200;
      18024: inst = 32'd136314880;
      18025: inst = 32'd268468224;
      18026: inst = 32'd201346549;
      18027: inst = 32'd203484854;
      18028: inst = 32'd471859200;
      18029: inst = 32'd136314880;
      18030: inst = 32'd268468224;
      18031: inst = 32'd201346550;
      18032: inst = 32'd203484854;
      18033: inst = 32'd471859200;
      18034: inst = 32'd136314880;
      18035: inst = 32'd268468224;
      18036: inst = 32'd201346551;
      18037: inst = 32'd203484854;
      18038: inst = 32'd471859200;
      18039: inst = 32'd136314880;
      18040: inst = 32'd268468224;
      18041: inst = 32'd201346552;
      18042: inst = 32'd203484854;
      18043: inst = 32'd471859200;
      18044: inst = 32'd136314880;
      18045: inst = 32'd268468224;
      18046: inst = 32'd201346553;
      18047: inst = 32'd203484854;
      18048: inst = 32'd471859200;
      18049: inst = 32'd136314880;
      18050: inst = 32'd268468224;
      18051: inst = 32'd201346554;
      18052: inst = 32'd203484854;
      18053: inst = 32'd471859200;
      18054: inst = 32'd136314880;
      18055: inst = 32'd268468224;
      18056: inst = 32'd201346555;
      18057: inst = 32'd203484854;
      18058: inst = 32'd471859200;
      18059: inst = 32'd136314880;
      18060: inst = 32'd268468224;
      18061: inst = 32'd201346556;
      18062: inst = 32'd203484854;
      18063: inst = 32'd471859200;
      18064: inst = 32'd136314880;
      18065: inst = 32'd268468224;
      18066: inst = 32'd201346557;
      18067: inst = 32'd203484854;
      18068: inst = 32'd471859200;
      18069: inst = 32'd136314880;
      18070: inst = 32'd268468224;
      18071: inst = 32'd201346558;
      18072: inst = 32'd203484854;
      18073: inst = 32'd471859200;
      18074: inst = 32'd136314880;
      18075: inst = 32'd268468224;
      18076: inst = 32'd201346559;
      18077: inst = 32'd203484854;
      18078: inst = 32'd471859200;
      18079: inst = 32'd136314880;
      18080: inst = 32'd268468224;
      18081: inst = 32'd201346560;
      18082: inst = 32'd203484854;
      18083: inst = 32'd471859200;
      18084: inst = 32'd136314880;
      18085: inst = 32'd268468224;
      18086: inst = 32'd201346561;
      18087: inst = 32'd203484854;
      18088: inst = 32'd471859200;
      18089: inst = 32'd136314880;
      18090: inst = 32'd268468224;
      18091: inst = 32'd201346562;
      18092: inst = 32'd203484854;
      18093: inst = 32'd471859200;
      18094: inst = 32'd136314880;
      18095: inst = 32'd268468224;
      18096: inst = 32'd201346563;
      18097: inst = 32'd203484854;
      18098: inst = 32'd471859200;
      18099: inst = 32'd136314880;
      18100: inst = 32'd268468224;
      18101: inst = 32'd201346564;
      18102: inst = 32'd203484854;
      18103: inst = 32'd471859200;
      18104: inst = 32'd136314880;
      18105: inst = 32'd268468224;
      18106: inst = 32'd201346565;
      18107: inst = 32'd203484854;
      18108: inst = 32'd471859200;
      18109: inst = 32'd136314880;
      18110: inst = 32'd268468224;
      18111: inst = 32'd201346566;
      18112: inst = 32'd203484854;
      18113: inst = 32'd471859200;
      18114: inst = 32'd136314880;
      18115: inst = 32'd268468224;
      18116: inst = 32'd201346567;
      18117: inst = 32'd203484854;
      18118: inst = 32'd471859200;
      18119: inst = 32'd136314880;
      18120: inst = 32'd268468224;
      18121: inst = 32'd201346568;
      18122: inst = 32'd203484854;
      18123: inst = 32'd471859200;
      18124: inst = 32'd136314880;
      18125: inst = 32'd268468224;
      18126: inst = 32'd201346569;
      18127: inst = 32'd203484854;
      18128: inst = 32'd471859200;
      18129: inst = 32'd136314880;
      18130: inst = 32'd268468224;
      18131: inst = 32'd201346570;
      18132: inst = 32'd203484854;
      18133: inst = 32'd471859200;
      18134: inst = 32'd136314880;
      18135: inst = 32'd268468224;
      18136: inst = 32'd201346571;
      18137: inst = 32'd203484854;
      18138: inst = 32'd471859200;
      18139: inst = 32'd136314880;
      18140: inst = 32'd268468224;
      18141: inst = 32'd201346572;
      18142: inst = 32'd203484854;
      18143: inst = 32'd471859200;
      18144: inst = 32'd136314880;
      18145: inst = 32'd268468224;
      18146: inst = 32'd201346573;
      18147: inst = 32'd203484854;
      18148: inst = 32'd471859200;
      18149: inst = 32'd136314880;
      18150: inst = 32'd268468224;
      18151: inst = 32'd201346574;
      18152: inst = 32'd203484854;
      18153: inst = 32'd471859200;
      18154: inst = 32'd136314880;
      18155: inst = 32'd268468224;
      18156: inst = 32'd201346575;
      18157: inst = 32'd203473634;
      18158: inst = 32'd471859200;
      18159: inst = 32'd136314880;
      18160: inst = 32'd268468224;
      18161: inst = 32'd201346576;
      18162: inst = 32'd203480005;
      18163: inst = 32'd471859200;
      18164: inst = 32'd136314880;
      18165: inst = 32'd268468224;
      18166: inst = 32'd201346577;
      18167: inst = 32'd203480005;
      18168: inst = 32'd471859200;
      18169: inst = 32'd136314880;
      18170: inst = 32'd268468224;
      18171: inst = 32'd201346578;
      18172: inst = 32'd203480005;
      18173: inst = 32'd471859200;
      18174: inst = 32'd136314880;
      18175: inst = 32'd268468224;
      18176: inst = 32'd201346579;
      18177: inst = 32'd203480005;
      18178: inst = 32'd471859200;
      18179: inst = 32'd136314880;
      18180: inst = 32'd268468224;
      18181: inst = 32'd201346580;
      18182: inst = 32'd203480005;
      18183: inst = 32'd471859200;
      18184: inst = 32'd136314880;
      18185: inst = 32'd268468224;
      18186: inst = 32'd201346581;
      18187: inst = 32'd203480005;
      18188: inst = 32'd471859200;
      18189: inst = 32'd136314880;
      18190: inst = 32'd268468224;
      18191: inst = 32'd201346582;
      18192: inst = 32'd203480005;
      18193: inst = 32'd471859200;
      18194: inst = 32'd136314880;
      18195: inst = 32'd268468224;
      18196: inst = 32'd201346583;
      18197: inst = 32'd203480005;
      18198: inst = 32'd471859200;
      18199: inst = 32'd136314880;
      18200: inst = 32'd268468224;
      18201: inst = 32'd201346584;
      18202: inst = 32'd203480005;
      18203: inst = 32'd471859200;
      18204: inst = 32'd136314880;
      18205: inst = 32'd268468224;
      18206: inst = 32'd201346585;
      18207: inst = 32'd203480005;
      18208: inst = 32'd471859200;
      18209: inst = 32'd136314880;
      18210: inst = 32'd268468224;
      18211: inst = 32'd201346586;
      18212: inst = 32'd203480005;
      18213: inst = 32'd471859200;
      18214: inst = 32'd136314880;
      18215: inst = 32'd268468224;
      18216: inst = 32'd201346587;
      18217: inst = 32'd203480005;
      18218: inst = 32'd471859200;
      18219: inst = 32'd136314880;
      18220: inst = 32'd268468224;
      18221: inst = 32'd201346588;
      18222: inst = 32'd203480005;
      18223: inst = 32'd471859200;
      18224: inst = 32'd136314880;
      18225: inst = 32'd268468224;
      18226: inst = 32'd201346589;
      18227: inst = 32'd203480005;
      18228: inst = 32'd471859200;
      18229: inst = 32'd136314880;
      18230: inst = 32'd268468224;
      18231: inst = 32'd201346590;
      18232: inst = 32'd203480005;
      18233: inst = 32'd471859200;
      18234: inst = 32'd136314880;
      18235: inst = 32'd268468224;
      18236: inst = 32'd201346591;
      18237: inst = 32'd203473634;
      18238: inst = 32'd471859200;
      18239: inst = 32'd136314880;
      18240: inst = 32'd268468224;
      18241: inst = 32'd201346592;
      18242: inst = 32'd203459697;
      18243: inst = 32'd471859200;
      18244: inst = 32'd136314880;
      18245: inst = 32'd268468224;
      18246: inst = 32'd201346593;
      18247: inst = 32'd203472343;
      18248: inst = 32'd471859200;
      18249: inst = 32'd136314880;
      18250: inst = 32'd268468224;
      18251: inst = 32'd201346594;
      18252: inst = 32'd203472343;
      18253: inst = 32'd471859200;
      18254: inst = 32'd136314880;
      18255: inst = 32'd268468224;
      18256: inst = 32'd201346595;
      18257: inst = 32'd203472343;
      18258: inst = 32'd471859200;
      18259: inst = 32'd136314880;
      18260: inst = 32'd268468224;
      18261: inst = 32'd201346596;
      18262: inst = 32'd203472343;
      18263: inst = 32'd471859200;
      18264: inst = 32'd136314880;
      18265: inst = 32'd268468224;
      18266: inst = 32'd201346597;
      18267: inst = 32'd203472343;
      18268: inst = 32'd471859200;
      18269: inst = 32'd136314880;
      18270: inst = 32'd268468224;
      18271: inst = 32'd201346598;
      18272: inst = 32'd203472343;
      18273: inst = 32'd471859200;
      18274: inst = 32'd136314880;
      18275: inst = 32'd268468224;
      18276: inst = 32'd201346599;
      18277: inst = 32'd203472343;
      18278: inst = 32'd471859200;
      18279: inst = 32'd136314880;
      18280: inst = 32'd268468224;
      18281: inst = 32'd201346600;
      18282: inst = 32'd203472343;
      18283: inst = 32'd471859200;
      18284: inst = 32'd136314880;
      18285: inst = 32'd268468224;
      18286: inst = 32'd201346601;
      18287: inst = 32'd203472343;
      18288: inst = 32'd471859200;
      18289: inst = 32'd136314880;
      18290: inst = 32'd268468224;
      18291: inst = 32'd201346602;
      18292: inst = 32'd203459697;
      18293: inst = 32'd471859200;
      18294: inst = 32'd136314880;
      18295: inst = 32'd268468224;
      18296: inst = 32'd201346603;
      18297: inst = 32'd203472343;
      18298: inst = 32'd471859200;
      18299: inst = 32'd136314880;
      18300: inst = 32'd268468224;
      18301: inst = 32'd201346604;
      18302: inst = 32'd203472343;
      18303: inst = 32'd471859200;
      18304: inst = 32'd136314880;
      18305: inst = 32'd268468224;
      18306: inst = 32'd201346605;
      18307: inst = 32'd203472343;
      18308: inst = 32'd471859200;
      18309: inst = 32'd136314880;
      18310: inst = 32'd268468224;
      18311: inst = 32'd201346606;
      18312: inst = 32'd203472343;
      18313: inst = 32'd471859200;
      18314: inst = 32'd136314880;
      18315: inst = 32'd268468224;
      18316: inst = 32'd201346607;
      18317: inst = 32'd203472343;
      18318: inst = 32'd471859200;
      18319: inst = 32'd136314880;
      18320: inst = 32'd268468224;
      18321: inst = 32'd201346608;
      18322: inst = 32'd203472343;
      18323: inst = 32'd471859200;
      18324: inst = 32'd136314880;
      18325: inst = 32'd268468224;
      18326: inst = 32'd201346609;
      18327: inst = 32'd203472343;
      18328: inst = 32'd471859200;
      18329: inst = 32'd136314880;
      18330: inst = 32'd268468224;
      18331: inst = 32'd201346610;
      18332: inst = 32'd203472343;
      18333: inst = 32'd471859200;
      18334: inst = 32'd136314880;
      18335: inst = 32'd268468224;
      18336: inst = 32'd201346611;
      18337: inst = 32'd203472343;
      18338: inst = 32'd471859200;
      18339: inst = 32'd136314880;
      18340: inst = 32'd268468224;
      18341: inst = 32'd201346612;
      18342: inst = 32'd203459697;
      18343: inst = 32'd471859200;
      18344: inst = 32'd136314880;
      18345: inst = 32'd268468224;
      18346: inst = 32'd201346613;
      18347: inst = 32'd203451245;
      18348: inst = 32'd471859200;
      18349: inst = 32'd136314880;
      18350: inst = 32'd268468224;
      18351: inst = 32'd201346614;
      18352: inst = 32'd203451245;
      18353: inst = 32'd471859200;
      18354: inst = 32'd136314880;
      18355: inst = 32'd268468224;
      18356: inst = 32'd201346615;
      18357: inst = 32'd203484854;
      18358: inst = 32'd471859200;
      18359: inst = 32'd136314880;
      18360: inst = 32'd268468224;
      18361: inst = 32'd201346616;
      18362: inst = 32'd203484854;
      18363: inst = 32'd471859200;
      18364: inst = 32'd136314880;
      18365: inst = 32'd268468224;
      18366: inst = 32'd201346617;
      18367: inst = 32'd203484854;
      18368: inst = 32'd471859200;
      18369: inst = 32'd136314880;
      18370: inst = 32'd268468224;
      18371: inst = 32'd201346618;
      18372: inst = 32'd203484854;
      18373: inst = 32'd471859200;
      18374: inst = 32'd136314880;
      18375: inst = 32'd268468224;
      18376: inst = 32'd201346619;
      18377: inst = 32'd203484854;
      18378: inst = 32'd471859200;
      18379: inst = 32'd136314880;
      18380: inst = 32'd268468224;
      18381: inst = 32'd201346620;
      18382: inst = 32'd203484854;
      18383: inst = 32'd471859200;
      18384: inst = 32'd136314880;
      18385: inst = 32'd268468224;
      18386: inst = 32'd201346621;
      18387: inst = 32'd203484854;
      18388: inst = 32'd471859200;
      18389: inst = 32'd136314880;
      18390: inst = 32'd268468224;
      18391: inst = 32'd201346622;
      18392: inst = 32'd203484854;
      18393: inst = 32'd471859200;
      18394: inst = 32'd136314880;
      18395: inst = 32'd268468224;
      18396: inst = 32'd201346623;
      18397: inst = 32'd203484854;
      18398: inst = 32'd471859200;
      18399: inst = 32'd136314880;
      18400: inst = 32'd268468224;
      18401: inst = 32'd201346624;
      18402: inst = 32'd203484854;
      18403: inst = 32'd471859200;
      18404: inst = 32'd136314880;
      18405: inst = 32'd268468224;
      18406: inst = 32'd201346625;
      18407: inst = 32'd203484854;
      18408: inst = 32'd471859200;
      18409: inst = 32'd136314880;
      18410: inst = 32'd268468224;
      18411: inst = 32'd201346626;
      18412: inst = 32'd203484854;
      18413: inst = 32'd471859200;
      18414: inst = 32'd136314880;
      18415: inst = 32'd268468224;
      18416: inst = 32'd201346627;
      18417: inst = 32'd203484854;
      18418: inst = 32'd471859200;
      18419: inst = 32'd136314880;
      18420: inst = 32'd268468224;
      18421: inst = 32'd201346628;
      18422: inst = 32'd203484854;
      18423: inst = 32'd471859200;
      18424: inst = 32'd136314880;
      18425: inst = 32'd268468224;
      18426: inst = 32'd201346629;
      18427: inst = 32'd203484854;
      18428: inst = 32'd471859200;
      18429: inst = 32'd136314880;
      18430: inst = 32'd268468224;
      18431: inst = 32'd201346630;
      18432: inst = 32'd203484854;
      18433: inst = 32'd471859200;
      18434: inst = 32'd136314880;
      18435: inst = 32'd268468224;
      18436: inst = 32'd201346631;
      18437: inst = 32'd203484854;
      18438: inst = 32'd471859200;
      18439: inst = 32'd136314880;
      18440: inst = 32'd268468224;
      18441: inst = 32'd201346632;
      18442: inst = 32'd203484854;
      18443: inst = 32'd471859200;
      18444: inst = 32'd136314880;
      18445: inst = 32'd268468224;
      18446: inst = 32'd201346633;
      18447: inst = 32'd203484854;
      18448: inst = 32'd471859200;
      18449: inst = 32'd136314880;
      18450: inst = 32'd268468224;
      18451: inst = 32'd201346634;
      18452: inst = 32'd203484854;
      18453: inst = 32'd471859200;
      18454: inst = 32'd136314880;
      18455: inst = 32'd268468224;
      18456: inst = 32'd201346635;
      18457: inst = 32'd203484854;
      18458: inst = 32'd471859200;
      18459: inst = 32'd136314880;
      18460: inst = 32'd268468224;
      18461: inst = 32'd201346636;
      18462: inst = 32'd203484854;
      18463: inst = 32'd471859200;
      18464: inst = 32'd136314880;
      18465: inst = 32'd268468224;
      18466: inst = 32'd201346637;
      18467: inst = 32'd203484854;
      18468: inst = 32'd471859200;
      18469: inst = 32'd136314880;
      18470: inst = 32'd268468224;
      18471: inst = 32'd201346638;
      18472: inst = 32'd203484854;
      18473: inst = 32'd471859200;
      18474: inst = 32'd136314880;
      18475: inst = 32'd268468224;
      18476: inst = 32'd201346639;
      18477: inst = 32'd203484854;
      18478: inst = 32'd471859200;
      18479: inst = 32'd136314880;
      18480: inst = 32'd268468224;
      18481: inst = 32'd201346640;
      18482: inst = 32'd203484854;
      18483: inst = 32'd471859200;
      18484: inst = 32'd136314880;
      18485: inst = 32'd268468224;
      18486: inst = 32'd201346641;
      18487: inst = 32'd203484854;
      18488: inst = 32'd471859200;
      18489: inst = 32'd136314880;
      18490: inst = 32'd268468224;
      18491: inst = 32'd201346642;
      18492: inst = 32'd203484854;
      18493: inst = 32'd471859200;
      18494: inst = 32'd136314880;
      18495: inst = 32'd268468224;
      18496: inst = 32'd201346643;
      18497: inst = 32'd203484854;
      18498: inst = 32'd471859200;
      18499: inst = 32'd136314880;
      18500: inst = 32'd268468224;
      18501: inst = 32'd201346644;
      18502: inst = 32'd203484854;
      18503: inst = 32'd471859200;
      18504: inst = 32'd136314880;
      18505: inst = 32'd268468224;
      18506: inst = 32'd201346645;
      18507: inst = 32'd203484854;
      18508: inst = 32'd471859200;
      18509: inst = 32'd136314880;
      18510: inst = 32'd268468224;
      18511: inst = 32'd201346646;
      18512: inst = 32'd203484854;
      18513: inst = 32'd471859200;
      18514: inst = 32'd136314880;
      18515: inst = 32'd268468224;
      18516: inst = 32'd201346647;
      18517: inst = 32'd203484854;
      18518: inst = 32'd471859200;
      18519: inst = 32'd136314880;
      18520: inst = 32'd268468224;
      18521: inst = 32'd201346648;
      18522: inst = 32'd203484854;
      18523: inst = 32'd471859200;
      18524: inst = 32'd136314880;
      18525: inst = 32'd268468224;
      18526: inst = 32'd201346649;
      18527: inst = 32'd203484854;
      18528: inst = 32'd471859200;
      18529: inst = 32'd136314880;
      18530: inst = 32'd268468224;
      18531: inst = 32'd201346650;
      18532: inst = 32'd203484854;
      18533: inst = 32'd471859200;
      18534: inst = 32'd136314880;
      18535: inst = 32'd268468224;
      18536: inst = 32'd201346651;
      18537: inst = 32'd203484854;
      18538: inst = 32'd471859200;
      18539: inst = 32'd136314880;
      18540: inst = 32'd268468224;
      18541: inst = 32'd201346652;
      18542: inst = 32'd203484854;
      18543: inst = 32'd471859200;
      18544: inst = 32'd136314880;
      18545: inst = 32'd268468224;
      18546: inst = 32'd201346653;
      18547: inst = 32'd203484854;
      18548: inst = 32'd471859200;
      18549: inst = 32'd136314880;
      18550: inst = 32'd268468224;
      18551: inst = 32'd201346654;
      18552: inst = 32'd203484854;
      18553: inst = 32'd471859200;
      18554: inst = 32'd136314880;
      18555: inst = 32'd268468224;
      18556: inst = 32'd201346655;
      18557: inst = 32'd203484854;
      18558: inst = 32'd471859200;
      18559: inst = 32'd136314880;
      18560: inst = 32'd268468224;
      18561: inst = 32'd201346656;
      18562: inst = 32'd203484854;
      18563: inst = 32'd471859200;
      18564: inst = 32'd136314880;
      18565: inst = 32'd268468224;
      18566: inst = 32'd201346657;
      18567: inst = 32'd203484854;
      18568: inst = 32'd471859200;
      18569: inst = 32'd136314880;
      18570: inst = 32'd268468224;
      18571: inst = 32'd201346658;
      18572: inst = 32'd203484854;
      18573: inst = 32'd471859200;
      18574: inst = 32'd136314880;
      18575: inst = 32'd268468224;
      18576: inst = 32'd201346659;
      18577: inst = 32'd203484854;
      18578: inst = 32'd471859200;
      18579: inst = 32'd136314880;
      18580: inst = 32'd268468224;
      18581: inst = 32'd201346660;
      18582: inst = 32'd203484854;
      18583: inst = 32'd471859200;
      18584: inst = 32'd136314880;
      18585: inst = 32'd268468224;
      18586: inst = 32'd201346661;
      18587: inst = 32'd203484854;
      18588: inst = 32'd471859200;
      18589: inst = 32'd136314880;
      18590: inst = 32'd268468224;
      18591: inst = 32'd201346662;
      18592: inst = 32'd203484854;
      18593: inst = 32'd471859200;
      18594: inst = 32'd136314880;
      18595: inst = 32'd268468224;
      18596: inst = 32'd201346663;
      18597: inst = 32'd203484854;
      18598: inst = 32'd471859200;
      18599: inst = 32'd136314880;
      18600: inst = 32'd268468224;
      18601: inst = 32'd201346664;
      18602: inst = 32'd203484854;
      18603: inst = 32'd471859200;
      18604: inst = 32'd136314880;
      18605: inst = 32'd268468224;
      18606: inst = 32'd201346665;
      18607: inst = 32'd203484854;
      18608: inst = 32'd471859200;
      18609: inst = 32'd136314880;
      18610: inst = 32'd268468224;
      18611: inst = 32'd201346666;
      18612: inst = 32'd203484854;
      18613: inst = 32'd471859200;
      18614: inst = 32'd136314880;
      18615: inst = 32'd268468224;
      18616: inst = 32'd201346667;
      18617: inst = 32'd203484854;
      18618: inst = 32'd471859200;
      18619: inst = 32'd136314880;
      18620: inst = 32'd268468224;
      18621: inst = 32'd201346668;
      18622: inst = 32'd203484854;
      18623: inst = 32'd471859200;
      18624: inst = 32'd136314880;
      18625: inst = 32'd268468224;
      18626: inst = 32'd201346669;
      18627: inst = 32'd203484854;
      18628: inst = 32'd471859200;
      18629: inst = 32'd136314880;
      18630: inst = 32'd268468224;
      18631: inst = 32'd201346670;
      18632: inst = 32'd203484854;
      18633: inst = 32'd471859200;
      18634: inst = 32'd136314880;
      18635: inst = 32'd268468224;
      18636: inst = 32'd201346671;
      18637: inst = 32'd203473634;
      18638: inst = 32'd471859200;
      18639: inst = 32'd136314880;
      18640: inst = 32'd268468224;
      18641: inst = 32'd201346672;
      18642: inst = 32'd203480005;
      18643: inst = 32'd471859200;
      18644: inst = 32'd136314880;
      18645: inst = 32'd268468224;
      18646: inst = 32'd201346673;
      18647: inst = 32'd203480005;
      18648: inst = 32'd471859200;
      18649: inst = 32'd136314880;
      18650: inst = 32'd268468224;
      18651: inst = 32'd201346674;
      18652: inst = 32'd203480005;
      18653: inst = 32'd471859200;
      18654: inst = 32'd136314880;
      18655: inst = 32'd268468224;
      18656: inst = 32'd201346675;
      18657: inst = 32'd203480005;
      18658: inst = 32'd471859200;
      18659: inst = 32'd136314880;
      18660: inst = 32'd268468224;
      18661: inst = 32'd201346676;
      18662: inst = 32'd203480005;
      18663: inst = 32'd471859200;
      18664: inst = 32'd136314880;
      18665: inst = 32'd268468224;
      18666: inst = 32'd201346677;
      18667: inst = 32'd203480005;
      18668: inst = 32'd471859200;
      18669: inst = 32'd136314880;
      18670: inst = 32'd268468224;
      18671: inst = 32'd201346678;
      18672: inst = 32'd203480005;
      18673: inst = 32'd471859200;
      18674: inst = 32'd136314880;
      18675: inst = 32'd268468224;
      18676: inst = 32'd201346679;
      18677: inst = 32'd203480005;
      18678: inst = 32'd471859200;
      18679: inst = 32'd136314880;
      18680: inst = 32'd268468224;
      18681: inst = 32'd201346680;
      18682: inst = 32'd203480005;
      18683: inst = 32'd471859200;
      18684: inst = 32'd136314880;
      18685: inst = 32'd268468224;
      18686: inst = 32'd201346681;
      18687: inst = 32'd203480005;
      18688: inst = 32'd471859200;
      18689: inst = 32'd136314880;
      18690: inst = 32'd268468224;
      18691: inst = 32'd201346682;
      18692: inst = 32'd203480005;
      18693: inst = 32'd471859200;
      18694: inst = 32'd136314880;
      18695: inst = 32'd268468224;
      18696: inst = 32'd201346683;
      18697: inst = 32'd203480005;
      18698: inst = 32'd471859200;
      18699: inst = 32'd136314880;
      18700: inst = 32'd268468224;
      18701: inst = 32'd201346684;
      18702: inst = 32'd203480005;
      18703: inst = 32'd471859200;
      18704: inst = 32'd136314880;
      18705: inst = 32'd268468224;
      18706: inst = 32'd201346685;
      18707: inst = 32'd203480005;
      18708: inst = 32'd471859200;
      18709: inst = 32'd136314880;
      18710: inst = 32'd268468224;
      18711: inst = 32'd201346686;
      18712: inst = 32'd203480005;
      18713: inst = 32'd471859200;
      18714: inst = 32'd136314880;
      18715: inst = 32'd268468224;
      18716: inst = 32'd201346687;
      18717: inst = 32'd203473634;
      18718: inst = 32'd471859200;
      18719: inst = 32'd136314880;
      18720: inst = 32'd268468224;
      18721: inst = 32'd201346688;
      18722: inst = 32'd203459697;
      18723: inst = 32'd471859200;
      18724: inst = 32'd136314880;
      18725: inst = 32'd268468224;
      18726: inst = 32'd201346689;
      18727: inst = 32'd203472343;
      18728: inst = 32'd471859200;
      18729: inst = 32'd136314880;
      18730: inst = 32'd268468224;
      18731: inst = 32'd201346690;
      18732: inst = 32'd203472343;
      18733: inst = 32'd471859200;
      18734: inst = 32'd136314880;
      18735: inst = 32'd268468224;
      18736: inst = 32'd201346691;
      18737: inst = 32'd203472343;
      18738: inst = 32'd471859200;
      18739: inst = 32'd136314880;
      18740: inst = 32'd268468224;
      18741: inst = 32'd201346692;
      18742: inst = 32'd203472343;
      18743: inst = 32'd471859200;
      18744: inst = 32'd136314880;
      18745: inst = 32'd268468224;
      18746: inst = 32'd201346693;
      18747: inst = 32'd203472343;
      18748: inst = 32'd471859200;
      18749: inst = 32'd136314880;
      18750: inst = 32'd268468224;
      18751: inst = 32'd201346694;
      18752: inst = 32'd203472343;
      18753: inst = 32'd471859200;
      18754: inst = 32'd136314880;
      18755: inst = 32'd268468224;
      18756: inst = 32'd201346695;
      18757: inst = 32'd203472343;
      18758: inst = 32'd471859200;
      18759: inst = 32'd136314880;
      18760: inst = 32'd268468224;
      18761: inst = 32'd201346696;
      18762: inst = 32'd203472343;
      18763: inst = 32'd471859200;
      18764: inst = 32'd136314880;
      18765: inst = 32'd268468224;
      18766: inst = 32'd201346697;
      18767: inst = 32'd203472343;
      18768: inst = 32'd471859200;
      18769: inst = 32'd136314880;
      18770: inst = 32'd268468224;
      18771: inst = 32'd201346698;
      18772: inst = 32'd203459697;
      18773: inst = 32'd471859200;
      18774: inst = 32'd136314880;
      18775: inst = 32'd268468224;
      18776: inst = 32'd201346699;
      18777: inst = 32'd203472343;
      18778: inst = 32'd471859200;
      18779: inst = 32'd136314880;
      18780: inst = 32'd268468224;
      18781: inst = 32'd201346700;
      18782: inst = 32'd203472343;
      18783: inst = 32'd471859200;
      18784: inst = 32'd136314880;
      18785: inst = 32'd268468224;
      18786: inst = 32'd201346701;
      18787: inst = 32'd203472343;
      18788: inst = 32'd471859200;
      18789: inst = 32'd136314880;
      18790: inst = 32'd268468224;
      18791: inst = 32'd201346702;
      18792: inst = 32'd203472343;
      18793: inst = 32'd471859200;
      18794: inst = 32'd136314880;
      18795: inst = 32'd268468224;
      18796: inst = 32'd201346703;
      18797: inst = 32'd203472343;
      18798: inst = 32'd471859200;
      18799: inst = 32'd136314880;
      18800: inst = 32'd268468224;
      18801: inst = 32'd201346704;
      18802: inst = 32'd203472343;
      18803: inst = 32'd471859200;
      18804: inst = 32'd136314880;
      18805: inst = 32'd268468224;
      18806: inst = 32'd201346705;
      18807: inst = 32'd203472343;
      18808: inst = 32'd471859200;
      18809: inst = 32'd136314880;
      18810: inst = 32'd268468224;
      18811: inst = 32'd201346706;
      18812: inst = 32'd203472343;
      18813: inst = 32'd471859200;
      18814: inst = 32'd136314880;
      18815: inst = 32'd268468224;
      18816: inst = 32'd201346707;
      18817: inst = 32'd203472343;
      18818: inst = 32'd471859200;
      18819: inst = 32'd136314880;
      18820: inst = 32'd268468224;
      18821: inst = 32'd201346708;
      18822: inst = 32'd203459697;
      18823: inst = 32'd471859200;
      18824: inst = 32'd136314880;
      18825: inst = 32'd268468224;
      18826: inst = 32'd201346709;
      18827: inst = 32'd203451245;
      18828: inst = 32'd471859200;
      18829: inst = 32'd136314880;
      18830: inst = 32'd268468224;
      18831: inst = 32'd201346710;
      18832: inst = 32'd203451245;
      18833: inst = 32'd471859200;
      18834: inst = 32'd136314880;
      18835: inst = 32'd268468224;
      18836: inst = 32'd201346711;
      18837: inst = 32'd203484854;
      18838: inst = 32'd471859200;
      18839: inst = 32'd136314880;
      18840: inst = 32'd268468224;
      18841: inst = 32'd201346712;
      18842: inst = 32'd203484854;
      18843: inst = 32'd471859200;
      18844: inst = 32'd136314880;
      18845: inst = 32'd268468224;
      18846: inst = 32'd201346713;
      18847: inst = 32'd203484854;
      18848: inst = 32'd471859200;
      18849: inst = 32'd136314880;
      18850: inst = 32'd268468224;
      18851: inst = 32'd201346714;
      18852: inst = 32'd203484854;
      18853: inst = 32'd471859200;
      18854: inst = 32'd136314880;
      18855: inst = 32'd268468224;
      18856: inst = 32'd201346715;
      18857: inst = 32'd203484854;
      18858: inst = 32'd471859200;
      18859: inst = 32'd136314880;
      18860: inst = 32'd268468224;
      18861: inst = 32'd201346716;
      18862: inst = 32'd203484854;
      18863: inst = 32'd471859200;
      18864: inst = 32'd136314880;
      18865: inst = 32'd268468224;
      18866: inst = 32'd201346717;
      18867: inst = 32'd203484854;
      18868: inst = 32'd471859200;
      18869: inst = 32'd136314880;
      18870: inst = 32'd268468224;
      18871: inst = 32'd201346718;
      18872: inst = 32'd203484854;
      18873: inst = 32'd471859200;
      18874: inst = 32'd136314880;
      18875: inst = 32'd268468224;
      18876: inst = 32'd201346719;
      18877: inst = 32'd203472243;
      18878: inst = 32'd471859200;
      18879: inst = 32'd136314880;
      18880: inst = 32'd268468224;
      18881: inst = 32'd201346720;
      18882: inst = 32'd203447021;
      18883: inst = 32'd471859200;
      18884: inst = 32'd136314880;
      18885: inst = 32'd268468224;
      18886: inst = 32'd201346721;
      18887: inst = 32'd203447021;
      18888: inst = 32'd471859200;
      18889: inst = 32'd136314880;
      18890: inst = 32'd268468224;
      18891: inst = 32'd201346722;
      18892: inst = 32'd203447021;
      18893: inst = 32'd471859200;
      18894: inst = 32'd136314880;
      18895: inst = 32'd268468224;
      18896: inst = 32'd201346723;
      18897: inst = 32'd203447021;
      18898: inst = 32'd471859200;
      18899: inst = 32'd136314880;
      18900: inst = 32'd268468224;
      18901: inst = 32'd201346724;
      18902: inst = 32'd203447021;
      18903: inst = 32'd471859200;
      18904: inst = 32'd136314880;
      18905: inst = 32'd268468224;
      18906: inst = 32'd201346725;
      18907: inst = 32'd203455406;
      18908: inst = 32'd471859200;
      18909: inst = 32'd136314880;
      18910: inst = 32'd268468224;
      18911: inst = 32'd201346726;
      18912: inst = 32'd203474356;
      18913: inst = 32'd471859200;
      18914: inst = 32'd136314880;
      18915: inst = 32'd268468224;
      18916: inst = 32'd201346727;
      18917: inst = 32'd203478516;
      18918: inst = 32'd471859200;
      18919: inst = 32'd136314880;
      18920: inst = 32'd268468224;
      18921: inst = 32'd201346728;
      18922: inst = 32'd203484854;
      18923: inst = 32'd471859200;
      18924: inst = 32'd136314880;
      18925: inst = 32'd268468224;
      18926: inst = 32'd201346729;
      18927: inst = 32'd203484854;
      18928: inst = 32'd471859200;
      18929: inst = 32'd136314880;
      18930: inst = 32'd268468224;
      18931: inst = 32'd201346730;
      18932: inst = 32'd203484854;
      18933: inst = 32'd471859200;
      18934: inst = 32'd136314880;
      18935: inst = 32'd268468224;
      18936: inst = 32'd201346731;
      18937: inst = 32'd203484854;
      18938: inst = 32'd471859200;
      18939: inst = 32'd136314880;
      18940: inst = 32'd268468224;
      18941: inst = 32'd201346732;
      18942: inst = 32'd203484854;
      18943: inst = 32'd471859200;
      18944: inst = 32'd136314880;
      18945: inst = 32'd268468224;
      18946: inst = 32'd201346733;
      18947: inst = 32'd203484854;
      18948: inst = 32'd471859200;
      18949: inst = 32'd136314880;
      18950: inst = 32'd268468224;
      18951: inst = 32'd201346734;
      18952: inst = 32'd203484854;
      18953: inst = 32'd471859200;
      18954: inst = 32'd136314880;
      18955: inst = 32'd268468224;
      18956: inst = 32'd201346735;
      18957: inst = 32'd203484854;
      18958: inst = 32'd471859200;
      18959: inst = 32'd136314880;
      18960: inst = 32'd268468224;
      18961: inst = 32'd201346736;
      18962: inst = 32'd203484854;
      18963: inst = 32'd471859200;
      18964: inst = 32'd136314880;
      18965: inst = 32'd268468224;
      18966: inst = 32'd201346737;
      18967: inst = 32'd203484854;
      18968: inst = 32'd471859200;
      18969: inst = 32'd136314880;
      18970: inst = 32'd268468224;
      18971: inst = 32'd201346738;
      18972: inst = 32'd203484854;
      18973: inst = 32'd471859200;
      18974: inst = 32'd136314880;
      18975: inst = 32'd268468224;
      18976: inst = 32'd201346739;
      18977: inst = 32'd203484854;
      18978: inst = 32'd471859200;
      18979: inst = 32'd136314880;
      18980: inst = 32'd268468224;
      18981: inst = 32'd201346740;
      18982: inst = 32'd203484854;
      18983: inst = 32'd471859200;
      18984: inst = 32'd136314880;
      18985: inst = 32'd268468224;
      18986: inst = 32'd201346741;
      18987: inst = 32'd203484854;
      18988: inst = 32'd471859200;
      18989: inst = 32'd136314880;
      18990: inst = 32'd268468224;
      18991: inst = 32'd201346742;
      18992: inst = 32'd203484854;
      18993: inst = 32'd471859200;
      18994: inst = 32'd136314880;
      18995: inst = 32'd268468224;
      18996: inst = 32'd201346743;
      18997: inst = 32'd203484854;
      18998: inst = 32'd471859200;
      18999: inst = 32'd136314880;
      19000: inst = 32'd268468224;
      19001: inst = 32'd201346744;
      19002: inst = 32'd203478516;
      19003: inst = 32'd471859200;
      19004: inst = 32'd136314880;
      19005: inst = 32'd268468224;
      19006: inst = 32'd201346745;
      19007: inst = 32'd203474356;
      19008: inst = 32'd471859200;
      19009: inst = 32'd136314880;
      19010: inst = 32'd268468224;
      19011: inst = 32'd201346746;
      19012: inst = 32'd203455406;
      19013: inst = 32'd471859200;
      19014: inst = 32'd136314880;
      19015: inst = 32'd268468224;
      19016: inst = 32'd201346747;
      19017: inst = 32'd203447021;
      19018: inst = 32'd471859200;
      19019: inst = 32'd136314880;
      19020: inst = 32'd268468224;
      19021: inst = 32'd201346748;
      19022: inst = 32'd203447021;
      19023: inst = 32'd471859200;
      19024: inst = 32'd136314880;
      19025: inst = 32'd268468224;
      19026: inst = 32'd201346749;
      19027: inst = 32'd203447021;
      19028: inst = 32'd471859200;
      19029: inst = 32'd136314880;
      19030: inst = 32'd268468224;
      19031: inst = 32'd201346750;
      19032: inst = 32'd203447021;
      19033: inst = 32'd471859200;
      19034: inst = 32'd136314880;
      19035: inst = 32'd268468224;
      19036: inst = 32'd201346751;
      19037: inst = 32'd203447021;
      19038: inst = 32'd471859200;
      19039: inst = 32'd136314880;
      19040: inst = 32'd268468224;
      19041: inst = 32'd201346752;
      19042: inst = 32'd203472243;
      19043: inst = 32'd471859200;
      19044: inst = 32'd136314880;
      19045: inst = 32'd268468224;
      19046: inst = 32'd201346753;
      19047: inst = 32'd203484854;
      19048: inst = 32'd471859200;
      19049: inst = 32'd136314880;
      19050: inst = 32'd268468224;
      19051: inst = 32'd201346754;
      19052: inst = 32'd203484854;
      19053: inst = 32'd471859200;
      19054: inst = 32'd136314880;
      19055: inst = 32'd268468224;
      19056: inst = 32'd201346755;
      19057: inst = 32'd203484854;
      19058: inst = 32'd471859200;
      19059: inst = 32'd136314880;
      19060: inst = 32'd268468224;
      19061: inst = 32'd201346756;
      19062: inst = 32'd203484854;
      19063: inst = 32'd471859200;
      19064: inst = 32'd136314880;
      19065: inst = 32'd268468224;
      19066: inst = 32'd201346757;
      19067: inst = 32'd203484854;
      19068: inst = 32'd471859200;
      19069: inst = 32'd136314880;
      19070: inst = 32'd268468224;
      19071: inst = 32'd201346758;
      19072: inst = 32'd203484854;
      19073: inst = 32'd471859200;
      19074: inst = 32'd136314880;
      19075: inst = 32'd268468224;
      19076: inst = 32'd201346759;
      19077: inst = 32'd203484854;
      19078: inst = 32'd471859200;
      19079: inst = 32'd136314880;
      19080: inst = 32'd268468224;
      19081: inst = 32'd201346760;
      19082: inst = 32'd203484854;
      19083: inst = 32'd471859200;
      19084: inst = 32'd136314880;
      19085: inst = 32'd268468224;
      19086: inst = 32'd201346761;
      19087: inst = 32'd203484854;
      19088: inst = 32'd471859200;
      19089: inst = 32'd136314880;
      19090: inst = 32'd268468224;
      19091: inst = 32'd201346762;
      19092: inst = 32'd203484854;
      19093: inst = 32'd471859200;
      19094: inst = 32'd136314880;
      19095: inst = 32'd268468224;
      19096: inst = 32'd201346763;
      19097: inst = 32'd203484854;
      19098: inst = 32'd471859200;
      19099: inst = 32'd136314880;
      19100: inst = 32'd268468224;
      19101: inst = 32'd201346764;
      19102: inst = 32'd203484854;
      19103: inst = 32'd471859200;
      19104: inst = 32'd136314880;
      19105: inst = 32'd268468224;
      19106: inst = 32'd201346765;
      19107: inst = 32'd203484854;
      19108: inst = 32'd471859200;
      19109: inst = 32'd136314880;
      19110: inst = 32'd268468224;
      19111: inst = 32'd201346766;
      19112: inst = 32'd203484854;
      19113: inst = 32'd471859200;
      19114: inst = 32'd136314880;
      19115: inst = 32'd268468224;
      19116: inst = 32'd201346767;
      19117: inst = 32'd203473634;
      19118: inst = 32'd471859200;
      19119: inst = 32'd136314880;
      19120: inst = 32'd268468224;
      19121: inst = 32'd201346768;
      19122: inst = 32'd203480005;
      19123: inst = 32'd471859200;
      19124: inst = 32'd136314880;
      19125: inst = 32'd268468224;
      19126: inst = 32'd201346769;
      19127: inst = 32'd203480005;
      19128: inst = 32'd471859200;
      19129: inst = 32'd136314880;
      19130: inst = 32'd268468224;
      19131: inst = 32'd201346770;
      19132: inst = 32'd203480005;
      19133: inst = 32'd471859200;
      19134: inst = 32'd136314880;
      19135: inst = 32'd268468224;
      19136: inst = 32'd201346771;
      19137: inst = 32'd203480005;
      19138: inst = 32'd471859200;
      19139: inst = 32'd136314880;
      19140: inst = 32'd268468224;
      19141: inst = 32'd201346772;
      19142: inst = 32'd203480005;
      19143: inst = 32'd471859200;
      19144: inst = 32'd136314880;
      19145: inst = 32'd268468224;
      19146: inst = 32'd201346773;
      19147: inst = 32'd203480005;
      19148: inst = 32'd471859200;
      19149: inst = 32'd136314880;
      19150: inst = 32'd268468224;
      19151: inst = 32'd201346774;
      19152: inst = 32'd203480005;
      19153: inst = 32'd471859200;
      19154: inst = 32'd136314880;
      19155: inst = 32'd268468224;
      19156: inst = 32'd201346775;
      19157: inst = 32'd203480005;
      19158: inst = 32'd471859200;
      19159: inst = 32'd136314880;
      19160: inst = 32'd268468224;
      19161: inst = 32'd201346776;
      19162: inst = 32'd203480005;
      19163: inst = 32'd471859200;
      19164: inst = 32'd136314880;
      19165: inst = 32'd268468224;
      19166: inst = 32'd201346777;
      19167: inst = 32'd203480005;
      19168: inst = 32'd471859200;
      19169: inst = 32'd136314880;
      19170: inst = 32'd268468224;
      19171: inst = 32'd201346778;
      19172: inst = 32'd203480005;
      19173: inst = 32'd471859200;
      19174: inst = 32'd136314880;
      19175: inst = 32'd268468224;
      19176: inst = 32'd201346779;
      19177: inst = 32'd203480005;
      19178: inst = 32'd471859200;
      19179: inst = 32'd136314880;
      19180: inst = 32'd268468224;
      19181: inst = 32'd201346780;
      19182: inst = 32'd203480005;
      19183: inst = 32'd471859200;
      19184: inst = 32'd136314880;
      19185: inst = 32'd268468224;
      19186: inst = 32'd201346781;
      19187: inst = 32'd203480005;
      19188: inst = 32'd471859200;
      19189: inst = 32'd136314880;
      19190: inst = 32'd268468224;
      19191: inst = 32'd201346782;
      19192: inst = 32'd203480005;
      19193: inst = 32'd471859200;
      19194: inst = 32'd136314880;
      19195: inst = 32'd268468224;
      19196: inst = 32'd201346783;
      19197: inst = 32'd203473634;
      19198: inst = 32'd471859200;
      19199: inst = 32'd136314880;
      19200: inst = 32'd268468224;
      19201: inst = 32'd201346784;
      19202: inst = 32'd203459697;
      19203: inst = 32'd471859200;
      19204: inst = 32'd136314880;
      19205: inst = 32'd268468224;
      19206: inst = 32'd201346785;
      19207: inst = 32'd203472343;
      19208: inst = 32'd471859200;
      19209: inst = 32'd136314880;
      19210: inst = 32'd268468224;
      19211: inst = 32'd201346786;
      19212: inst = 32'd203472343;
      19213: inst = 32'd471859200;
      19214: inst = 32'd136314880;
      19215: inst = 32'd268468224;
      19216: inst = 32'd201346787;
      19217: inst = 32'd203472343;
      19218: inst = 32'd471859200;
      19219: inst = 32'd136314880;
      19220: inst = 32'd268468224;
      19221: inst = 32'd201346788;
      19222: inst = 32'd203472343;
      19223: inst = 32'd471859200;
      19224: inst = 32'd136314880;
      19225: inst = 32'd268468224;
      19226: inst = 32'd201346789;
      19227: inst = 32'd203472343;
      19228: inst = 32'd471859200;
      19229: inst = 32'd136314880;
      19230: inst = 32'd268468224;
      19231: inst = 32'd201346790;
      19232: inst = 32'd203472343;
      19233: inst = 32'd471859200;
      19234: inst = 32'd136314880;
      19235: inst = 32'd268468224;
      19236: inst = 32'd201346791;
      19237: inst = 32'd203472343;
      19238: inst = 32'd471859200;
      19239: inst = 32'd136314880;
      19240: inst = 32'd268468224;
      19241: inst = 32'd201346792;
      19242: inst = 32'd203472343;
      19243: inst = 32'd471859200;
      19244: inst = 32'd136314880;
      19245: inst = 32'd268468224;
      19246: inst = 32'd201346793;
      19247: inst = 32'd203472343;
      19248: inst = 32'd471859200;
      19249: inst = 32'd136314880;
      19250: inst = 32'd268468224;
      19251: inst = 32'd201346794;
      19252: inst = 32'd203459697;
      19253: inst = 32'd471859200;
      19254: inst = 32'd136314880;
      19255: inst = 32'd268468224;
      19256: inst = 32'd201346795;
      19257: inst = 32'd203472343;
      19258: inst = 32'd471859200;
      19259: inst = 32'd136314880;
      19260: inst = 32'd268468224;
      19261: inst = 32'd201346796;
      19262: inst = 32'd203472343;
      19263: inst = 32'd471859200;
      19264: inst = 32'd136314880;
      19265: inst = 32'd268468224;
      19266: inst = 32'd201346797;
      19267: inst = 32'd203472343;
      19268: inst = 32'd471859200;
      19269: inst = 32'd136314880;
      19270: inst = 32'd268468224;
      19271: inst = 32'd201346798;
      19272: inst = 32'd203472343;
      19273: inst = 32'd471859200;
      19274: inst = 32'd136314880;
      19275: inst = 32'd268468224;
      19276: inst = 32'd201346799;
      19277: inst = 32'd203472343;
      19278: inst = 32'd471859200;
      19279: inst = 32'd136314880;
      19280: inst = 32'd268468224;
      19281: inst = 32'd201346800;
      19282: inst = 32'd203472343;
      19283: inst = 32'd471859200;
      19284: inst = 32'd136314880;
      19285: inst = 32'd268468224;
      19286: inst = 32'd201346801;
      19287: inst = 32'd203472343;
      19288: inst = 32'd471859200;
      19289: inst = 32'd136314880;
      19290: inst = 32'd268468224;
      19291: inst = 32'd201346802;
      19292: inst = 32'd203472343;
      19293: inst = 32'd471859200;
      19294: inst = 32'd136314880;
      19295: inst = 32'd268468224;
      19296: inst = 32'd201346803;
      19297: inst = 32'd203472343;
      19298: inst = 32'd471859200;
      19299: inst = 32'd136314880;
      19300: inst = 32'd268468224;
      19301: inst = 32'd201346804;
      19302: inst = 32'd203459697;
      19303: inst = 32'd471859200;
      19304: inst = 32'd136314880;
      19305: inst = 32'd268468224;
      19306: inst = 32'd201346805;
      19307: inst = 32'd203451245;
      19308: inst = 32'd471859200;
      19309: inst = 32'd136314880;
      19310: inst = 32'd268468224;
      19311: inst = 32'd201346806;
      19312: inst = 32'd203451245;
      19313: inst = 32'd471859200;
      19314: inst = 32'd136314880;
      19315: inst = 32'd268468224;
      19316: inst = 32'd201346807;
      19317: inst = 32'd203484854;
      19318: inst = 32'd471859200;
      19319: inst = 32'd136314880;
      19320: inst = 32'd268468224;
      19321: inst = 32'd201346808;
      19322: inst = 32'd203484854;
      19323: inst = 32'd471859200;
      19324: inst = 32'd136314880;
      19325: inst = 32'd268468224;
      19326: inst = 32'd201346809;
      19327: inst = 32'd203484854;
      19328: inst = 32'd471859200;
      19329: inst = 32'd136314880;
      19330: inst = 32'd268468224;
      19331: inst = 32'd201346810;
      19332: inst = 32'd203484854;
      19333: inst = 32'd471859200;
      19334: inst = 32'd136314880;
      19335: inst = 32'd268468224;
      19336: inst = 32'd201346811;
      19337: inst = 32'd203484854;
      19338: inst = 32'd471859200;
      19339: inst = 32'd136314880;
      19340: inst = 32'd268468224;
      19341: inst = 32'd201346812;
      19342: inst = 32'd203484854;
      19343: inst = 32'd471859200;
      19344: inst = 32'd136314880;
      19345: inst = 32'd268468224;
      19346: inst = 32'd201346813;
      19347: inst = 32'd203484854;
      19348: inst = 32'd471859200;
      19349: inst = 32'd136314880;
      19350: inst = 32'd268468224;
      19351: inst = 32'd201346814;
      19352: inst = 32'd203484854;
      19353: inst = 32'd471859200;
      19354: inst = 32'd136314880;
      19355: inst = 32'd268468224;
      19356: inst = 32'd201346815;
      19357: inst = 32'd203465905;
      19358: inst = 32'd471859200;
      19359: inst = 32'd136314880;
      19360: inst = 32'd268468224;
      19361: inst = 32'd201346816;
      19362: inst = 32'd203447021;
      19363: inst = 32'd471859200;
      19364: inst = 32'd136314880;
      19365: inst = 32'd268468224;
      19366: inst = 32'd201346817;
      19367: inst = 32'd203447021;
      19368: inst = 32'd471859200;
      19369: inst = 32'd136314880;
      19370: inst = 32'd268468224;
      19371: inst = 32'd201346818;
      19372: inst = 32'd203447021;
      19373: inst = 32'd471859200;
      19374: inst = 32'd136314880;
      19375: inst = 32'd268468224;
      19376: inst = 32'd201346819;
      19377: inst = 32'd203447021;
      19378: inst = 32'd471859200;
      19379: inst = 32'd136314880;
      19380: inst = 32'd268468224;
      19381: inst = 32'd201346820;
      19382: inst = 32'd203447021;
      19383: inst = 32'd471859200;
      19384: inst = 32'd136314880;
      19385: inst = 32'd268468224;
      19386: inst = 32'd201346821;
      19387: inst = 32'd203447021;
      19388: inst = 32'd471859200;
      19389: inst = 32'd136314880;
      19390: inst = 32'd268468224;
      19391: inst = 32'd201346822;
      19392: inst = 32'd203449069;
      19393: inst = 32'd471859200;
      19394: inst = 32'd136314880;
      19395: inst = 32'd268468224;
      19396: inst = 32'd201346823;
      19397: inst = 32'd203461712;
      19398: inst = 32'd471859200;
      19399: inst = 32'd136314880;
      19400: inst = 32'd268468224;
      19401: inst = 32'd201346824;
      19402: inst = 32'd203484854;
      19403: inst = 32'd471859200;
      19404: inst = 32'd136314880;
      19405: inst = 32'd268468224;
      19406: inst = 32'd201346825;
      19407: inst = 32'd203484854;
      19408: inst = 32'd471859200;
      19409: inst = 32'd136314880;
      19410: inst = 32'd268468224;
      19411: inst = 32'd201346826;
      19412: inst = 32'd203484854;
      19413: inst = 32'd471859200;
      19414: inst = 32'd136314880;
      19415: inst = 32'd268468224;
      19416: inst = 32'd201346827;
      19417: inst = 32'd203484854;
      19418: inst = 32'd471859200;
      19419: inst = 32'd136314880;
      19420: inst = 32'd268468224;
      19421: inst = 32'd201346828;
      19422: inst = 32'd203484854;
      19423: inst = 32'd471859200;
      19424: inst = 32'd136314880;
      19425: inst = 32'd268468224;
      19426: inst = 32'd201346829;
      19427: inst = 32'd203484854;
      19428: inst = 32'd471859200;
      19429: inst = 32'd136314880;
      19430: inst = 32'd268468224;
      19431: inst = 32'd201346830;
      19432: inst = 32'd203484854;
      19433: inst = 32'd471859200;
      19434: inst = 32'd136314880;
      19435: inst = 32'd268468224;
      19436: inst = 32'd201346831;
      19437: inst = 32'd203484854;
      19438: inst = 32'd471859200;
      19439: inst = 32'd136314880;
      19440: inst = 32'd268468224;
      19441: inst = 32'd201346832;
      19442: inst = 32'd203484854;
      19443: inst = 32'd471859200;
      19444: inst = 32'd136314880;
      19445: inst = 32'd268468224;
      19446: inst = 32'd201346833;
      19447: inst = 32'd203484854;
      19448: inst = 32'd471859200;
      19449: inst = 32'd136314880;
      19450: inst = 32'd268468224;
      19451: inst = 32'd201346834;
      19452: inst = 32'd203484854;
      19453: inst = 32'd471859200;
      19454: inst = 32'd136314880;
      19455: inst = 32'd268468224;
      19456: inst = 32'd201346835;
      19457: inst = 32'd203484854;
      19458: inst = 32'd471859200;
      19459: inst = 32'd136314880;
      19460: inst = 32'd268468224;
      19461: inst = 32'd201346836;
      19462: inst = 32'd203484854;
      19463: inst = 32'd471859200;
      19464: inst = 32'd136314880;
      19465: inst = 32'd268468224;
      19466: inst = 32'd201346837;
      19467: inst = 32'd203484854;
      19468: inst = 32'd471859200;
      19469: inst = 32'd136314880;
      19470: inst = 32'd268468224;
      19471: inst = 32'd201346838;
      19472: inst = 32'd203484854;
      19473: inst = 32'd471859200;
      19474: inst = 32'd136314880;
      19475: inst = 32'd268468224;
      19476: inst = 32'd201346839;
      19477: inst = 32'd203484854;
      19478: inst = 32'd471859200;
      19479: inst = 32'd136314880;
      19480: inst = 32'd268468224;
      19481: inst = 32'd201346840;
      19482: inst = 32'd203461712;
      19483: inst = 32'd471859200;
      19484: inst = 32'd136314880;
      19485: inst = 32'd268468224;
      19486: inst = 32'd201346841;
      19487: inst = 32'd203449069;
      19488: inst = 32'd471859200;
      19489: inst = 32'd136314880;
      19490: inst = 32'd268468224;
      19491: inst = 32'd201346842;
      19492: inst = 32'd203447021;
      19493: inst = 32'd471859200;
      19494: inst = 32'd136314880;
      19495: inst = 32'd268468224;
      19496: inst = 32'd201346843;
      19497: inst = 32'd203447021;
      19498: inst = 32'd471859200;
      19499: inst = 32'd136314880;
      19500: inst = 32'd268468224;
      19501: inst = 32'd201346844;
      19502: inst = 32'd203447021;
      19503: inst = 32'd471859200;
      19504: inst = 32'd136314880;
      19505: inst = 32'd268468224;
      19506: inst = 32'd201346845;
      19507: inst = 32'd203447021;
      19508: inst = 32'd471859200;
      19509: inst = 32'd136314880;
      19510: inst = 32'd268468224;
      19511: inst = 32'd201346846;
      19512: inst = 32'd203447021;
      19513: inst = 32'd471859200;
      19514: inst = 32'd136314880;
      19515: inst = 32'd268468224;
      19516: inst = 32'd201346847;
      19517: inst = 32'd203447021;
      19518: inst = 32'd471859200;
      19519: inst = 32'd136314880;
      19520: inst = 32'd268468224;
      19521: inst = 32'd201346848;
      19522: inst = 32'd203465905;
      19523: inst = 32'd471859200;
      19524: inst = 32'd136314880;
      19525: inst = 32'd268468224;
      19526: inst = 32'd201346849;
      19527: inst = 32'd203484854;
      19528: inst = 32'd471859200;
      19529: inst = 32'd136314880;
      19530: inst = 32'd268468224;
      19531: inst = 32'd201346850;
      19532: inst = 32'd203484854;
      19533: inst = 32'd471859200;
      19534: inst = 32'd136314880;
      19535: inst = 32'd268468224;
      19536: inst = 32'd201346851;
      19537: inst = 32'd203484854;
      19538: inst = 32'd471859200;
      19539: inst = 32'd136314880;
      19540: inst = 32'd268468224;
      19541: inst = 32'd201346852;
      19542: inst = 32'd203484854;
      19543: inst = 32'd471859200;
      19544: inst = 32'd136314880;
      19545: inst = 32'd268468224;
      19546: inst = 32'd201346853;
      19547: inst = 32'd203484854;
      19548: inst = 32'd471859200;
      19549: inst = 32'd136314880;
      19550: inst = 32'd268468224;
      19551: inst = 32'd201346854;
      19552: inst = 32'd203484854;
      19553: inst = 32'd471859200;
      19554: inst = 32'd136314880;
      19555: inst = 32'd268468224;
      19556: inst = 32'd201346855;
      19557: inst = 32'd203484854;
      19558: inst = 32'd471859200;
      19559: inst = 32'd136314880;
      19560: inst = 32'd268468224;
      19561: inst = 32'd201346856;
      19562: inst = 32'd203484854;
      19563: inst = 32'd471859200;
      19564: inst = 32'd136314880;
      19565: inst = 32'd268468224;
      19566: inst = 32'd201346857;
      19567: inst = 32'd203484854;
      19568: inst = 32'd471859200;
      19569: inst = 32'd136314880;
      19570: inst = 32'd268468224;
      19571: inst = 32'd201346858;
      19572: inst = 32'd203484854;
      19573: inst = 32'd471859200;
      19574: inst = 32'd136314880;
      19575: inst = 32'd268468224;
      19576: inst = 32'd201346859;
      19577: inst = 32'd203484854;
      19578: inst = 32'd471859200;
      19579: inst = 32'd136314880;
      19580: inst = 32'd268468224;
      19581: inst = 32'd201346860;
      19582: inst = 32'd203484854;
      19583: inst = 32'd471859200;
      19584: inst = 32'd136314880;
      19585: inst = 32'd268468224;
      19586: inst = 32'd201346861;
      19587: inst = 32'd203484854;
      19588: inst = 32'd471859200;
      19589: inst = 32'd136314880;
      19590: inst = 32'd268468224;
      19591: inst = 32'd201346862;
      19592: inst = 32'd203484854;
      19593: inst = 32'd471859200;
      19594: inst = 32'd136314880;
      19595: inst = 32'd268468224;
      19596: inst = 32'd201346863;
      19597: inst = 32'd203473634;
      19598: inst = 32'd471859200;
      19599: inst = 32'd136314880;
      19600: inst = 32'd268468224;
      19601: inst = 32'd201346864;
      19602: inst = 32'd203480005;
      19603: inst = 32'd471859200;
      19604: inst = 32'd136314880;
      19605: inst = 32'd268468224;
      19606: inst = 32'd201346865;
      19607: inst = 32'd203480005;
      19608: inst = 32'd471859200;
      19609: inst = 32'd136314880;
      19610: inst = 32'd268468224;
      19611: inst = 32'd201346866;
      19612: inst = 32'd203480005;
      19613: inst = 32'd471859200;
      19614: inst = 32'd136314880;
      19615: inst = 32'd268468224;
      19616: inst = 32'd201346867;
      19617: inst = 32'd203480005;
      19618: inst = 32'd471859200;
      19619: inst = 32'd136314880;
      19620: inst = 32'd268468224;
      19621: inst = 32'd201346868;
      19622: inst = 32'd203480005;
      19623: inst = 32'd471859200;
      19624: inst = 32'd136314880;
      19625: inst = 32'd268468224;
      19626: inst = 32'd201346869;
      19627: inst = 32'd203480005;
      19628: inst = 32'd471859200;
      19629: inst = 32'd136314880;
      19630: inst = 32'd268468224;
      19631: inst = 32'd201346870;
      19632: inst = 32'd203480005;
      19633: inst = 32'd471859200;
      19634: inst = 32'd136314880;
      19635: inst = 32'd268468224;
      19636: inst = 32'd201346871;
      19637: inst = 32'd203480005;
      19638: inst = 32'd471859200;
      19639: inst = 32'd136314880;
      19640: inst = 32'd268468224;
      19641: inst = 32'd201346872;
      19642: inst = 32'd203480005;
      19643: inst = 32'd471859200;
      19644: inst = 32'd136314880;
      19645: inst = 32'd268468224;
      19646: inst = 32'd201346873;
      19647: inst = 32'd203480005;
      19648: inst = 32'd471859200;
      19649: inst = 32'd136314880;
      19650: inst = 32'd268468224;
      19651: inst = 32'd201346874;
      19652: inst = 32'd203480005;
      19653: inst = 32'd471859200;
      19654: inst = 32'd136314880;
      19655: inst = 32'd268468224;
      19656: inst = 32'd201346875;
      19657: inst = 32'd203480005;
      19658: inst = 32'd471859200;
      19659: inst = 32'd136314880;
      19660: inst = 32'd268468224;
      19661: inst = 32'd201346876;
      19662: inst = 32'd203480005;
      19663: inst = 32'd471859200;
      19664: inst = 32'd136314880;
      19665: inst = 32'd268468224;
      19666: inst = 32'd201346877;
      19667: inst = 32'd203480005;
      19668: inst = 32'd471859200;
      19669: inst = 32'd136314880;
      19670: inst = 32'd268468224;
      19671: inst = 32'd201346878;
      19672: inst = 32'd203480005;
      19673: inst = 32'd471859200;
      19674: inst = 32'd136314880;
      19675: inst = 32'd268468224;
      19676: inst = 32'd201346879;
      19677: inst = 32'd203473634;
      19678: inst = 32'd471859200;
      19679: inst = 32'd136314880;
      19680: inst = 32'd268468224;
      19681: inst = 32'd201346880;
      19682: inst = 32'd203459697;
      19683: inst = 32'd471859200;
      19684: inst = 32'd136314880;
      19685: inst = 32'd268468224;
      19686: inst = 32'd201346881;
      19687: inst = 32'd203472343;
      19688: inst = 32'd471859200;
      19689: inst = 32'd136314880;
      19690: inst = 32'd268468224;
      19691: inst = 32'd201346882;
      19692: inst = 32'd203472343;
      19693: inst = 32'd471859200;
      19694: inst = 32'd136314880;
      19695: inst = 32'd268468224;
      19696: inst = 32'd201346883;
      19697: inst = 32'd203472343;
      19698: inst = 32'd471859200;
      19699: inst = 32'd136314880;
      19700: inst = 32'd268468224;
      19701: inst = 32'd201346884;
      19702: inst = 32'd203472343;
      19703: inst = 32'd471859200;
      19704: inst = 32'd136314880;
      19705: inst = 32'd268468224;
      19706: inst = 32'd201346885;
      19707: inst = 32'd203472343;
      19708: inst = 32'd471859200;
      19709: inst = 32'd136314880;
      19710: inst = 32'd268468224;
      19711: inst = 32'd201346886;
      19712: inst = 32'd203472343;
      19713: inst = 32'd471859200;
      19714: inst = 32'd136314880;
      19715: inst = 32'd268468224;
      19716: inst = 32'd201346887;
      19717: inst = 32'd203472343;
      19718: inst = 32'd471859200;
      19719: inst = 32'd136314880;
      19720: inst = 32'd268468224;
      19721: inst = 32'd201346888;
      19722: inst = 32'd203472343;
      19723: inst = 32'd471859200;
      19724: inst = 32'd136314880;
      19725: inst = 32'd268468224;
      19726: inst = 32'd201346889;
      19727: inst = 32'd203472343;
      19728: inst = 32'd471859200;
      19729: inst = 32'd136314880;
      19730: inst = 32'd268468224;
      19731: inst = 32'd201346890;
      19732: inst = 32'd203459697;
      19733: inst = 32'd471859200;
      19734: inst = 32'd136314880;
      19735: inst = 32'd268468224;
      19736: inst = 32'd201346891;
      19737: inst = 32'd203472343;
      19738: inst = 32'd471859200;
      19739: inst = 32'd136314880;
      19740: inst = 32'd268468224;
      19741: inst = 32'd201346892;
      19742: inst = 32'd203472343;
      19743: inst = 32'd471859200;
      19744: inst = 32'd136314880;
      19745: inst = 32'd268468224;
      19746: inst = 32'd201346893;
      19747: inst = 32'd203472343;
      19748: inst = 32'd471859200;
      19749: inst = 32'd136314880;
      19750: inst = 32'd268468224;
      19751: inst = 32'd201346894;
      19752: inst = 32'd203472343;
      19753: inst = 32'd471859200;
      19754: inst = 32'd136314880;
      19755: inst = 32'd268468224;
      19756: inst = 32'd201346895;
      19757: inst = 32'd203472343;
      19758: inst = 32'd471859200;
      19759: inst = 32'd136314880;
      19760: inst = 32'd268468224;
      19761: inst = 32'd201346896;
      19762: inst = 32'd203472343;
      19763: inst = 32'd471859200;
      19764: inst = 32'd136314880;
      19765: inst = 32'd268468224;
      19766: inst = 32'd201346897;
      19767: inst = 32'd203472343;
      19768: inst = 32'd471859200;
      19769: inst = 32'd136314880;
      19770: inst = 32'd268468224;
      19771: inst = 32'd201346898;
      19772: inst = 32'd203472343;
      19773: inst = 32'd471859200;
      19774: inst = 32'd136314880;
      19775: inst = 32'd268468224;
      19776: inst = 32'd201346899;
      19777: inst = 32'd203472343;
      19778: inst = 32'd471859200;
      19779: inst = 32'd136314880;
      19780: inst = 32'd268468224;
      19781: inst = 32'd201346900;
      19782: inst = 32'd203459697;
      19783: inst = 32'd471859200;
      19784: inst = 32'd136314880;
      19785: inst = 32'd268468224;
      19786: inst = 32'd201346901;
      19787: inst = 32'd203451245;
      19788: inst = 32'd471859200;
      19789: inst = 32'd136314880;
      19790: inst = 32'd268468224;
      19791: inst = 32'd201346902;
      19792: inst = 32'd203451245;
      19793: inst = 32'd471859200;
      19794: inst = 32'd136314880;
      19795: inst = 32'd268468224;
      19796: inst = 32'd201346903;
      19797: inst = 32'd203484854;
      19798: inst = 32'd471859200;
      19799: inst = 32'd136314880;
      19800: inst = 32'd268468224;
      19801: inst = 32'd201346904;
      19802: inst = 32'd203484854;
      19803: inst = 32'd471859200;
      19804: inst = 32'd136314880;
      19805: inst = 32'd268468224;
      19806: inst = 32'd201346905;
      19807: inst = 32'd203484854;
      19808: inst = 32'd471859200;
      19809: inst = 32'd136314880;
      19810: inst = 32'd268468224;
      19811: inst = 32'd201346906;
      19812: inst = 32'd203484854;
      19813: inst = 32'd471859200;
      19814: inst = 32'd136314880;
      19815: inst = 32'd268468224;
      19816: inst = 32'd201346907;
      19817: inst = 32'd203484854;
      19818: inst = 32'd471859200;
      19819: inst = 32'd136314880;
      19820: inst = 32'd268468224;
      19821: inst = 32'd201346908;
      19822: inst = 32'd203484854;
      19823: inst = 32'd471859200;
      19824: inst = 32'd136314880;
      19825: inst = 32'd268468224;
      19826: inst = 32'd201346909;
      19827: inst = 32'd203484854;
      19828: inst = 32'd471859200;
      19829: inst = 32'd136314880;
      19830: inst = 32'd268468224;
      19831: inst = 32'd201346910;
      19832: inst = 32'd203484854;
      19833: inst = 32'd471859200;
      19834: inst = 32'd136314880;
      19835: inst = 32'd268468224;
      19836: inst = 32'd201346911;
      19837: inst = 32'd203465937;
      19838: inst = 32'd471859200;
      19839: inst = 32'd136314880;
      19840: inst = 32'd268468224;
      19841: inst = 32'd201346912;
      19842: inst = 32'd203447021;
      19843: inst = 32'd471859200;
      19844: inst = 32'd136314880;
      19845: inst = 32'd268468224;
      19846: inst = 32'd201346913;
      19847: inst = 32'd203447021;
      19848: inst = 32'd471859200;
      19849: inst = 32'd136314880;
      19850: inst = 32'd268468224;
      19851: inst = 32'd201346914;
      19852: inst = 32'd203447021;
      19853: inst = 32'd471859200;
      19854: inst = 32'd136314880;
      19855: inst = 32'd268468224;
      19856: inst = 32'd201346915;
      19857: inst = 32'd203447021;
      19858: inst = 32'd471859200;
      19859: inst = 32'd136314880;
      19860: inst = 32'd268468224;
      19861: inst = 32'd201346916;
      19862: inst = 32'd203447021;
      19863: inst = 32'd471859200;
      19864: inst = 32'd136314880;
      19865: inst = 32'd268468224;
      19866: inst = 32'd201346917;
      19867: inst = 32'd203447021;
      19868: inst = 32'd471859200;
      19869: inst = 32'd136314880;
      19870: inst = 32'd268468224;
      19871: inst = 32'd201346918;
      19872: inst = 32'd203447021;
      19873: inst = 32'd471859200;
      19874: inst = 32'd136314880;
      19875: inst = 32'd268468224;
      19876: inst = 32'd201346919;
      19877: inst = 32'd203447021;
      19878: inst = 32'd471859200;
      19879: inst = 32'd136314880;
      19880: inst = 32'd268468224;
      19881: inst = 32'd201346920;
      19882: inst = 32'd203484854;
      19883: inst = 32'd471859200;
      19884: inst = 32'd136314880;
      19885: inst = 32'd268468224;
      19886: inst = 32'd201346921;
      19887: inst = 32'd203484854;
      19888: inst = 32'd471859200;
      19889: inst = 32'd136314880;
      19890: inst = 32'd268468224;
      19891: inst = 32'd201346922;
      19892: inst = 32'd203484854;
      19893: inst = 32'd471859200;
      19894: inst = 32'd136314880;
      19895: inst = 32'd268468224;
      19896: inst = 32'd201346923;
      19897: inst = 32'd203484854;
      19898: inst = 32'd471859200;
      19899: inst = 32'd136314880;
      19900: inst = 32'd268468224;
      19901: inst = 32'd201346924;
      19902: inst = 32'd203484854;
      19903: inst = 32'd471859200;
      19904: inst = 32'd136314880;
      19905: inst = 32'd268468224;
      19906: inst = 32'd201346925;
      19907: inst = 32'd203484854;
      19908: inst = 32'd471859200;
      19909: inst = 32'd136314880;
      19910: inst = 32'd268468224;
      19911: inst = 32'd201346926;
      19912: inst = 32'd203484854;
      19913: inst = 32'd471859200;
      19914: inst = 32'd136314880;
      19915: inst = 32'd268468224;
      19916: inst = 32'd201346927;
      19917: inst = 32'd203484854;
      19918: inst = 32'd471859200;
      19919: inst = 32'd136314880;
      19920: inst = 32'd268468224;
      19921: inst = 32'd201346928;
      19922: inst = 32'd203484854;
      19923: inst = 32'd471859200;
      19924: inst = 32'd136314880;
      19925: inst = 32'd268468224;
      19926: inst = 32'd201346929;
      19927: inst = 32'd203484854;
      19928: inst = 32'd471859200;
      19929: inst = 32'd136314880;
      19930: inst = 32'd268468224;
      19931: inst = 32'd201346930;
      19932: inst = 32'd203484854;
      19933: inst = 32'd471859200;
      19934: inst = 32'd136314880;
      19935: inst = 32'd268468224;
      19936: inst = 32'd201346931;
      19937: inst = 32'd203484854;
      19938: inst = 32'd471859200;
      19939: inst = 32'd136314880;
      19940: inst = 32'd268468224;
      19941: inst = 32'd201346932;
      19942: inst = 32'd203484854;
      19943: inst = 32'd471859200;
      19944: inst = 32'd136314880;
      19945: inst = 32'd268468224;
      19946: inst = 32'd201346933;
      19947: inst = 32'd203484854;
      19948: inst = 32'd471859200;
      19949: inst = 32'd136314880;
      19950: inst = 32'd268468224;
      19951: inst = 32'd201346934;
      19952: inst = 32'd203484854;
      19953: inst = 32'd471859200;
      19954: inst = 32'd136314880;
      19955: inst = 32'd268468224;
      19956: inst = 32'd201346935;
      19957: inst = 32'd203484854;
      19958: inst = 32'd471859200;
      19959: inst = 32'd136314880;
      19960: inst = 32'd268468224;
      19961: inst = 32'd201346936;
      19962: inst = 32'd203447021;
      19963: inst = 32'd471859200;
      19964: inst = 32'd136314880;
      19965: inst = 32'd268468224;
      19966: inst = 32'd201346937;
      19967: inst = 32'd203447021;
      19968: inst = 32'd471859200;
      19969: inst = 32'd136314880;
      19970: inst = 32'd268468224;
      19971: inst = 32'd201346938;
      19972: inst = 32'd203447021;
      19973: inst = 32'd471859200;
      19974: inst = 32'd136314880;
      19975: inst = 32'd268468224;
      19976: inst = 32'd201346939;
      19977: inst = 32'd203447021;
      19978: inst = 32'd471859200;
      19979: inst = 32'd136314880;
      19980: inst = 32'd268468224;
      19981: inst = 32'd201346940;
      19982: inst = 32'd203447021;
      19983: inst = 32'd471859200;
      19984: inst = 32'd136314880;
      19985: inst = 32'd268468224;
      19986: inst = 32'd201346941;
      19987: inst = 32'd203447021;
      19988: inst = 32'd471859200;
      19989: inst = 32'd136314880;
      19990: inst = 32'd268468224;
      19991: inst = 32'd201346942;
      19992: inst = 32'd203447021;
      19993: inst = 32'd471859200;
      19994: inst = 32'd136314880;
      19995: inst = 32'd268468224;
      19996: inst = 32'd201346943;
      19997: inst = 32'd203447021;
      19998: inst = 32'd471859200;
      19999: inst = 32'd136314880;
      20000: inst = 32'd268468224;
      20001: inst = 32'd201346944;
      20002: inst = 32'd203465937;
      20003: inst = 32'd471859200;
      20004: inst = 32'd136314880;
      20005: inst = 32'd268468224;
      20006: inst = 32'd201346945;
      20007: inst = 32'd203484854;
      20008: inst = 32'd471859200;
      20009: inst = 32'd136314880;
      20010: inst = 32'd268468224;
      20011: inst = 32'd201346946;
      20012: inst = 32'd203484854;
      20013: inst = 32'd471859200;
      20014: inst = 32'd136314880;
      20015: inst = 32'd268468224;
      20016: inst = 32'd201346947;
      20017: inst = 32'd203484854;
      20018: inst = 32'd471859200;
      20019: inst = 32'd136314880;
      20020: inst = 32'd268468224;
      20021: inst = 32'd201346948;
      20022: inst = 32'd203484854;
      20023: inst = 32'd471859200;
      20024: inst = 32'd136314880;
      20025: inst = 32'd268468224;
      20026: inst = 32'd201346949;
      20027: inst = 32'd203484854;
      20028: inst = 32'd471859200;
      20029: inst = 32'd136314880;
      20030: inst = 32'd268468224;
      20031: inst = 32'd201346950;
      20032: inst = 32'd203484854;
      20033: inst = 32'd471859200;
      20034: inst = 32'd136314880;
      20035: inst = 32'd268468224;
      20036: inst = 32'd201346951;
      20037: inst = 32'd203484854;
      20038: inst = 32'd471859200;
      20039: inst = 32'd136314880;
      20040: inst = 32'd268468224;
      20041: inst = 32'd201346952;
      20042: inst = 32'd203484854;
      20043: inst = 32'd471859200;
      20044: inst = 32'd136314880;
      20045: inst = 32'd268468224;
      20046: inst = 32'd201346953;
      20047: inst = 32'd203484854;
      20048: inst = 32'd471859200;
      20049: inst = 32'd136314880;
      20050: inst = 32'd268468224;
      20051: inst = 32'd201346954;
      20052: inst = 32'd203484854;
      20053: inst = 32'd471859200;
      20054: inst = 32'd136314880;
      20055: inst = 32'd268468224;
      20056: inst = 32'd201346955;
      20057: inst = 32'd203484854;
      20058: inst = 32'd471859200;
      20059: inst = 32'd136314880;
      20060: inst = 32'd268468224;
      20061: inst = 32'd201346956;
      20062: inst = 32'd203484854;
      20063: inst = 32'd471859200;
      20064: inst = 32'd136314880;
      20065: inst = 32'd268468224;
      20066: inst = 32'd201346957;
      20067: inst = 32'd203484854;
      20068: inst = 32'd471859200;
      20069: inst = 32'd136314880;
      20070: inst = 32'd268468224;
      20071: inst = 32'd201346958;
      20072: inst = 32'd203484854;
      20073: inst = 32'd471859200;
      20074: inst = 32'd136314880;
      20075: inst = 32'd268468224;
      20076: inst = 32'd201346959;
      20077: inst = 32'd203473634;
      20078: inst = 32'd471859200;
      20079: inst = 32'd136314880;
      20080: inst = 32'd268468224;
      20081: inst = 32'd201346960;
      20082: inst = 32'd203480005;
      20083: inst = 32'd471859200;
      20084: inst = 32'd136314880;
      20085: inst = 32'd268468224;
      20086: inst = 32'd201346961;
      20087: inst = 32'd203480005;
      20088: inst = 32'd471859200;
      20089: inst = 32'd136314880;
      20090: inst = 32'd268468224;
      20091: inst = 32'd201346962;
      20092: inst = 32'd203480005;
      20093: inst = 32'd471859200;
      20094: inst = 32'd136314880;
      20095: inst = 32'd268468224;
      20096: inst = 32'd201346963;
      20097: inst = 32'd203480005;
      20098: inst = 32'd471859200;
      20099: inst = 32'd136314880;
      20100: inst = 32'd268468224;
      20101: inst = 32'd201346964;
      20102: inst = 32'd203480005;
      20103: inst = 32'd471859200;
      20104: inst = 32'd136314880;
      20105: inst = 32'd268468224;
      20106: inst = 32'd201346965;
      20107: inst = 32'd203480005;
      20108: inst = 32'd471859200;
      20109: inst = 32'd136314880;
      20110: inst = 32'd268468224;
      20111: inst = 32'd201346966;
      20112: inst = 32'd203480005;
      20113: inst = 32'd471859200;
      20114: inst = 32'd136314880;
      20115: inst = 32'd268468224;
      20116: inst = 32'd201346967;
      20117: inst = 32'd203480005;
      20118: inst = 32'd471859200;
      20119: inst = 32'd136314880;
      20120: inst = 32'd268468224;
      20121: inst = 32'd201346968;
      20122: inst = 32'd203480005;
      20123: inst = 32'd471859200;
      20124: inst = 32'd136314880;
      20125: inst = 32'd268468224;
      20126: inst = 32'd201346969;
      20127: inst = 32'd203480005;
      20128: inst = 32'd471859200;
      20129: inst = 32'd136314880;
      20130: inst = 32'd268468224;
      20131: inst = 32'd201346970;
      20132: inst = 32'd203480005;
      20133: inst = 32'd471859200;
      20134: inst = 32'd136314880;
      20135: inst = 32'd268468224;
      20136: inst = 32'd201346971;
      20137: inst = 32'd203480005;
      20138: inst = 32'd471859200;
      20139: inst = 32'd136314880;
      20140: inst = 32'd268468224;
      20141: inst = 32'd201346972;
      20142: inst = 32'd203480005;
      20143: inst = 32'd471859200;
      20144: inst = 32'd136314880;
      20145: inst = 32'd268468224;
      20146: inst = 32'd201346973;
      20147: inst = 32'd203480005;
      20148: inst = 32'd471859200;
      20149: inst = 32'd136314880;
      20150: inst = 32'd268468224;
      20151: inst = 32'd201346974;
      20152: inst = 32'd203480005;
      20153: inst = 32'd471859200;
      20154: inst = 32'd136314880;
      20155: inst = 32'd268468224;
      20156: inst = 32'd201346975;
      20157: inst = 32'd203473634;
      20158: inst = 32'd471859200;
      20159: inst = 32'd136314880;
      20160: inst = 32'd268468224;
      20161: inst = 32'd201346976;
      20162: inst = 32'd203459697;
      20163: inst = 32'd471859200;
      20164: inst = 32'd136314880;
      20165: inst = 32'd268468224;
      20166: inst = 32'd201346977;
      20167: inst = 32'd203472343;
      20168: inst = 32'd471859200;
      20169: inst = 32'd136314880;
      20170: inst = 32'd268468224;
      20171: inst = 32'd201346978;
      20172: inst = 32'd203472343;
      20173: inst = 32'd471859200;
      20174: inst = 32'd136314880;
      20175: inst = 32'd268468224;
      20176: inst = 32'd201346979;
      20177: inst = 32'd203472343;
      20178: inst = 32'd471859200;
      20179: inst = 32'd136314880;
      20180: inst = 32'd268468224;
      20181: inst = 32'd201346980;
      20182: inst = 32'd203472343;
      20183: inst = 32'd471859200;
      20184: inst = 32'd136314880;
      20185: inst = 32'd268468224;
      20186: inst = 32'd201346981;
      20187: inst = 32'd203472343;
      20188: inst = 32'd471859200;
      20189: inst = 32'd136314880;
      20190: inst = 32'd268468224;
      20191: inst = 32'd201346982;
      20192: inst = 32'd203472343;
      20193: inst = 32'd471859200;
      20194: inst = 32'd136314880;
      20195: inst = 32'd268468224;
      20196: inst = 32'd201346983;
      20197: inst = 32'd203472343;
      20198: inst = 32'd471859200;
      20199: inst = 32'd136314880;
      20200: inst = 32'd268468224;
      20201: inst = 32'd201346984;
      20202: inst = 32'd203442761;
      20203: inst = 32'd471859200;
      20204: inst = 32'd136314880;
      20205: inst = 32'd268468224;
      20206: inst = 32'd201346985;
      20207: inst = 32'd203472343;
      20208: inst = 32'd471859200;
      20209: inst = 32'd136314880;
      20210: inst = 32'd268468224;
      20211: inst = 32'd201346986;
      20212: inst = 32'd203459697;
      20213: inst = 32'd471859200;
      20214: inst = 32'd136314880;
      20215: inst = 32'd268468224;
      20216: inst = 32'd201346987;
      20217: inst = 32'd203472343;
      20218: inst = 32'd471859200;
      20219: inst = 32'd136314880;
      20220: inst = 32'd268468224;
      20221: inst = 32'd201346988;
      20222: inst = 32'd203442761;
      20223: inst = 32'd471859200;
      20224: inst = 32'd136314880;
      20225: inst = 32'd268468224;
      20226: inst = 32'd201346989;
      20227: inst = 32'd203472343;
      20228: inst = 32'd471859200;
      20229: inst = 32'd136314880;
      20230: inst = 32'd268468224;
      20231: inst = 32'd201346990;
      20232: inst = 32'd203472343;
      20233: inst = 32'd471859200;
      20234: inst = 32'd136314880;
      20235: inst = 32'd268468224;
      20236: inst = 32'd201346991;
      20237: inst = 32'd203472343;
      20238: inst = 32'd471859200;
      20239: inst = 32'd136314880;
      20240: inst = 32'd268468224;
      20241: inst = 32'd201346992;
      20242: inst = 32'd203472343;
      20243: inst = 32'd471859200;
      20244: inst = 32'd136314880;
      20245: inst = 32'd268468224;
      20246: inst = 32'd201346993;
      20247: inst = 32'd203472343;
      20248: inst = 32'd471859200;
      20249: inst = 32'd136314880;
      20250: inst = 32'd268468224;
      20251: inst = 32'd201346994;
      20252: inst = 32'd203472343;
      20253: inst = 32'd471859200;
      20254: inst = 32'd136314880;
      20255: inst = 32'd268468224;
      20256: inst = 32'd201346995;
      20257: inst = 32'd203472343;
      20258: inst = 32'd471859200;
      20259: inst = 32'd136314880;
      20260: inst = 32'd268468224;
      20261: inst = 32'd201346996;
      20262: inst = 32'd203459697;
      20263: inst = 32'd471859200;
      20264: inst = 32'd136314880;
      20265: inst = 32'd268468224;
      20266: inst = 32'd201346997;
      20267: inst = 32'd203451245;
      20268: inst = 32'd471859200;
      20269: inst = 32'd136314880;
      20270: inst = 32'd268468224;
      20271: inst = 32'd201346998;
      20272: inst = 32'd203451245;
      20273: inst = 32'd471859200;
      20274: inst = 32'd136314880;
      20275: inst = 32'd268468224;
      20276: inst = 32'd201346999;
      20277: inst = 32'd203484854;
      20278: inst = 32'd471859200;
      20279: inst = 32'd136314880;
      20280: inst = 32'd268468224;
      20281: inst = 32'd201347000;
      20282: inst = 32'd203484854;
      20283: inst = 32'd471859200;
      20284: inst = 32'd136314880;
      20285: inst = 32'd268468224;
      20286: inst = 32'd201347001;
      20287: inst = 32'd203484854;
      20288: inst = 32'd471859200;
      20289: inst = 32'd136314880;
      20290: inst = 32'd268468224;
      20291: inst = 32'd201347002;
      20292: inst = 32'd203484854;
      20293: inst = 32'd471859200;
      20294: inst = 32'd136314880;
      20295: inst = 32'd268468224;
      20296: inst = 32'd201347003;
      20297: inst = 32'd203484854;
      20298: inst = 32'd471859200;
      20299: inst = 32'd136314880;
      20300: inst = 32'd268468224;
      20301: inst = 32'd201347004;
      20302: inst = 32'd203484854;
      20303: inst = 32'd471859200;
      20304: inst = 32'd136314880;
      20305: inst = 32'd268468224;
      20306: inst = 32'd201347005;
      20307: inst = 32'd203484854;
      20308: inst = 32'd471859200;
      20309: inst = 32'd136314880;
      20310: inst = 32'd268468224;
      20311: inst = 32'd201347006;
      20312: inst = 32'd203484854;
      20313: inst = 32'd471859200;
      20314: inst = 32'd136314880;
      20315: inst = 32'd268468224;
      20316: inst = 32'd201347007;
      20317: inst = 32'd203465905;
      20318: inst = 32'd471859200;
      20319: inst = 32'd136314880;
      20320: inst = 32'd268468224;
      20321: inst = 32'd201347008;
      20322: inst = 32'd203447021;
      20323: inst = 32'd471859200;
      20324: inst = 32'd136314880;
      20325: inst = 32'd268468224;
      20326: inst = 32'd201347009;
      20327: inst = 32'd203447021;
      20328: inst = 32'd471859200;
      20329: inst = 32'd136314880;
      20330: inst = 32'd268468224;
      20331: inst = 32'd201347010;
      20332: inst = 32'd203447021;
      20333: inst = 32'd471859200;
      20334: inst = 32'd136314880;
      20335: inst = 32'd268468224;
      20336: inst = 32'd201347011;
      20337: inst = 32'd203447021;
      20338: inst = 32'd471859200;
      20339: inst = 32'd136314880;
      20340: inst = 32'd268468224;
      20341: inst = 32'd201347012;
      20342: inst = 32'd203447021;
      20343: inst = 32'd471859200;
      20344: inst = 32'd136314880;
      20345: inst = 32'd268468224;
      20346: inst = 32'd201347013;
      20347: inst = 32'd203446987;
      20348: inst = 32'd471859200;
      20349: inst = 32'd136314880;
      20350: inst = 32'd268468224;
      20351: inst = 32'd201347014;
      20352: inst = 32'd203447021;
      20353: inst = 32'd471859200;
      20354: inst = 32'd136314880;
      20355: inst = 32'd268468224;
      20356: inst = 32'd201347015;
      20357: inst = 32'd203447021;
      20358: inst = 32'd471859200;
      20359: inst = 32'd136314880;
      20360: inst = 32'd268468224;
      20361: inst = 32'd201347016;
      20362: inst = 32'd203484854;
      20363: inst = 32'd471859200;
      20364: inst = 32'd136314880;
      20365: inst = 32'd268468224;
      20366: inst = 32'd201347017;
      20367: inst = 32'd203484854;
      20368: inst = 32'd471859200;
      20369: inst = 32'd136314880;
      20370: inst = 32'd268468224;
      20371: inst = 32'd201347018;
      20372: inst = 32'd203484854;
      20373: inst = 32'd471859200;
      20374: inst = 32'd136314880;
      20375: inst = 32'd268468224;
      20376: inst = 32'd201347019;
      20377: inst = 32'd203484854;
      20378: inst = 32'd471859200;
      20379: inst = 32'd136314880;
      20380: inst = 32'd268468224;
      20381: inst = 32'd201347020;
      20382: inst = 32'd203484854;
      20383: inst = 32'd471859200;
      20384: inst = 32'd136314880;
      20385: inst = 32'd268468224;
      20386: inst = 32'd201347021;
      20387: inst = 32'd203484854;
      20388: inst = 32'd471859200;
      20389: inst = 32'd136314880;
      20390: inst = 32'd268468224;
      20391: inst = 32'd201347022;
      20392: inst = 32'd203484854;
      20393: inst = 32'd471859200;
      20394: inst = 32'd136314880;
      20395: inst = 32'd268468224;
      20396: inst = 32'd201347023;
      20397: inst = 32'd203484854;
      20398: inst = 32'd471859200;
      20399: inst = 32'd136314880;
      20400: inst = 32'd268468224;
      20401: inst = 32'd201347024;
      20402: inst = 32'd203484854;
      20403: inst = 32'd471859200;
      20404: inst = 32'd136314880;
      20405: inst = 32'd268468224;
      20406: inst = 32'd201347025;
      20407: inst = 32'd203484854;
      20408: inst = 32'd471859200;
      20409: inst = 32'd136314880;
      20410: inst = 32'd268468224;
      20411: inst = 32'd201347026;
      20412: inst = 32'd203484854;
      20413: inst = 32'd471859200;
      20414: inst = 32'd136314880;
      20415: inst = 32'd268468224;
      20416: inst = 32'd201347027;
      20417: inst = 32'd203484854;
      20418: inst = 32'd471859200;
      20419: inst = 32'd136314880;
      20420: inst = 32'd268468224;
      20421: inst = 32'd201347028;
      20422: inst = 32'd203484854;
      20423: inst = 32'd471859200;
      20424: inst = 32'd136314880;
      20425: inst = 32'd268468224;
      20426: inst = 32'd201347029;
      20427: inst = 32'd203484854;
      20428: inst = 32'd471859200;
      20429: inst = 32'd136314880;
      20430: inst = 32'd268468224;
      20431: inst = 32'd201347030;
      20432: inst = 32'd203484854;
      20433: inst = 32'd471859200;
      20434: inst = 32'd136314880;
      20435: inst = 32'd268468224;
      20436: inst = 32'd201347031;
      20437: inst = 32'd203484854;
      20438: inst = 32'd471859200;
      20439: inst = 32'd136314880;
      20440: inst = 32'd268468224;
      20441: inst = 32'd201347032;
      20442: inst = 32'd203447021;
      20443: inst = 32'd471859200;
      20444: inst = 32'd136314880;
      20445: inst = 32'd268468224;
      20446: inst = 32'd201347033;
      20447: inst = 32'd203447021;
      20448: inst = 32'd471859200;
      20449: inst = 32'd136314880;
      20450: inst = 32'd268468224;
      20451: inst = 32'd201347034;
      20452: inst = 32'd203446987;
      20453: inst = 32'd471859200;
      20454: inst = 32'd136314880;
      20455: inst = 32'd268468224;
      20456: inst = 32'd201347035;
      20457: inst = 32'd203447021;
      20458: inst = 32'd471859200;
      20459: inst = 32'd136314880;
      20460: inst = 32'd268468224;
      20461: inst = 32'd201347036;
      20462: inst = 32'd203447021;
      20463: inst = 32'd471859200;
      20464: inst = 32'd136314880;
      20465: inst = 32'd268468224;
      20466: inst = 32'd201347037;
      20467: inst = 32'd203447021;
      20468: inst = 32'd471859200;
      20469: inst = 32'd136314880;
      20470: inst = 32'd268468224;
      20471: inst = 32'd201347038;
      20472: inst = 32'd203447021;
      20473: inst = 32'd471859200;
      20474: inst = 32'd136314880;
      20475: inst = 32'd268468224;
      20476: inst = 32'd201347039;
      20477: inst = 32'd203447021;
      20478: inst = 32'd471859200;
      20479: inst = 32'd136314880;
      20480: inst = 32'd268468224;
      20481: inst = 32'd201347040;
      20482: inst = 32'd203465905;
      20483: inst = 32'd471859200;
      20484: inst = 32'd136314880;
      20485: inst = 32'd268468224;
      20486: inst = 32'd201347041;
      20487: inst = 32'd203484854;
      20488: inst = 32'd471859200;
      20489: inst = 32'd136314880;
      20490: inst = 32'd268468224;
      20491: inst = 32'd201347042;
      20492: inst = 32'd203484854;
      20493: inst = 32'd471859200;
      20494: inst = 32'd136314880;
      20495: inst = 32'd268468224;
      20496: inst = 32'd201347043;
      20497: inst = 32'd203484854;
      20498: inst = 32'd471859200;
      20499: inst = 32'd136314880;
      20500: inst = 32'd268468224;
      20501: inst = 32'd201347044;
      20502: inst = 32'd203484854;
      20503: inst = 32'd471859200;
      20504: inst = 32'd136314880;
      20505: inst = 32'd268468224;
      20506: inst = 32'd201347045;
      20507: inst = 32'd203484854;
      20508: inst = 32'd471859200;
      20509: inst = 32'd136314880;
      20510: inst = 32'd268468224;
      20511: inst = 32'd201347046;
      20512: inst = 32'd203484854;
      20513: inst = 32'd471859200;
      20514: inst = 32'd136314880;
      20515: inst = 32'd268468224;
      20516: inst = 32'd201347047;
      20517: inst = 32'd203484854;
      20518: inst = 32'd471859200;
      20519: inst = 32'd136314880;
      20520: inst = 32'd268468224;
      20521: inst = 32'd201347048;
      20522: inst = 32'd203484854;
      20523: inst = 32'd471859200;
      20524: inst = 32'd136314880;
      20525: inst = 32'd268468224;
      20526: inst = 32'd201347049;
      20527: inst = 32'd203484854;
      20528: inst = 32'd471859200;
      20529: inst = 32'd136314880;
      20530: inst = 32'd268468224;
      20531: inst = 32'd201347050;
      20532: inst = 32'd203484854;
      20533: inst = 32'd471859200;
      20534: inst = 32'd136314880;
      20535: inst = 32'd268468224;
      20536: inst = 32'd201347051;
      20537: inst = 32'd203484854;
      20538: inst = 32'd471859200;
      20539: inst = 32'd136314880;
      20540: inst = 32'd268468224;
      20541: inst = 32'd201347052;
      20542: inst = 32'd203484854;
      20543: inst = 32'd471859200;
      20544: inst = 32'd136314880;
      20545: inst = 32'd268468224;
      20546: inst = 32'd201347053;
      20547: inst = 32'd203484854;
      20548: inst = 32'd471859200;
      20549: inst = 32'd136314880;
      20550: inst = 32'd268468224;
      20551: inst = 32'd201347054;
      20552: inst = 32'd203484854;
      20553: inst = 32'd471859200;
      20554: inst = 32'd136314880;
      20555: inst = 32'd268468224;
      20556: inst = 32'd201347055;
      20557: inst = 32'd203473634;
      20558: inst = 32'd471859200;
      20559: inst = 32'd136314880;
      20560: inst = 32'd268468224;
      20561: inst = 32'd201347056;
      20562: inst = 32'd203480005;
      20563: inst = 32'd471859200;
      20564: inst = 32'd136314880;
      20565: inst = 32'd268468224;
      20566: inst = 32'd201347057;
      20567: inst = 32'd203480005;
      20568: inst = 32'd471859200;
      20569: inst = 32'd136314880;
      20570: inst = 32'd268468224;
      20571: inst = 32'd201347058;
      20572: inst = 32'd203480005;
      20573: inst = 32'd471859200;
      20574: inst = 32'd136314880;
      20575: inst = 32'd268468224;
      20576: inst = 32'd201347059;
      20577: inst = 32'd203480005;
      20578: inst = 32'd471859200;
      20579: inst = 32'd136314880;
      20580: inst = 32'd268468224;
      20581: inst = 32'd201347060;
      20582: inst = 32'd203480005;
      20583: inst = 32'd471859200;
      20584: inst = 32'd136314880;
      20585: inst = 32'd268468224;
      20586: inst = 32'd201347061;
      20587: inst = 32'd203480005;
      20588: inst = 32'd471859200;
      20589: inst = 32'd136314880;
      20590: inst = 32'd268468224;
      20591: inst = 32'd201347062;
      20592: inst = 32'd203480005;
      20593: inst = 32'd471859200;
      20594: inst = 32'd136314880;
      20595: inst = 32'd268468224;
      20596: inst = 32'd201347063;
      20597: inst = 32'd203480005;
      20598: inst = 32'd471859200;
      20599: inst = 32'd136314880;
      20600: inst = 32'd268468224;
      20601: inst = 32'd201347064;
      20602: inst = 32'd203480005;
      20603: inst = 32'd471859200;
      20604: inst = 32'd136314880;
      20605: inst = 32'd268468224;
      20606: inst = 32'd201347065;
      20607: inst = 32'd203480005;
      20608: inst = 32'd471859200;
      20609: inst = 32'd136314880;
      20610: inst = 32'd268468224;
      20611: inst = 32'd201347066;
      20612: inst = 32'd203480005;
      20613: inst = 32'd471859200;
      20614: inst = 32'd136314880;
      20615: inst = 32'd268468224;
      20616: inst = 32'd201347067;
      20617: inst = 32'd203480005;
      20618: inst = 32'd471859200;
      20619: inst = 32'd136314880;
      20620: inst = 32'd268468224;
      20621: inst = 32'd201347068;
      20622: inst = 32'd203480005;
      20623: inst = 32'd471859200;
      20624: inst = 32'd136314880;
      20625: inst = 32'd268468224;
      20626: inst = 32'd201347069;
      20627: inst = 32'd203480005;
      20628: inst = 32'd471859200;
      20629: inst = 32'd136314880;
      20630: inst = 32'd268468224;
      20631: inst = 32'd201347070;
      20632: inst = 32'd203480005;
      20633: inst = 32'd471859200;
      20634: inst = 32'd136314880;
      20635: inst = 32'd268468224;
      20636: inst = 32'd201347071;
      20637: inst = 32'd203473634;
      20638: inst = 32'd471859200;
      20639: inst = 32'd136314880;
      20640: inst = 32'd268468224;
      20641: inst = 32'd201347072;
      20642: inst = 32'd203459697;
      20643: inst = 32'd471859200;
      20644: inst = 32'd136314880;
      20645: inst = 32'd268468224;
      20646: inst = 32'd201347073;
      20647: inst = 32'd203472343;
      20648: inst = 32'd471859200;
      20649: inst = 32'd136314880;
      20650: inst = 32'd268468224;
      20651: inst = 32'd201347074;
      20652: inst = 32'd203472343;
      20653: inst = 32'd471859200;
      20654: inst = 32'd136314880;
      20655: inst = 32'd268468224;
      20656: inst = 32'd201347075;
      20657: inst = 32'd203472343;
      20658: inst = 32'd471859200;
      20659: inst = 32'd136314880;
      20660: inst = 32'd268468224;
      20661: inst = 32'd201347076;
      20662: inst = 32'd203472343;
      20663: inst = 32'd471859200;
      20664: inst = 32'd136314880;
      20665: inst = 32'd268468224;
      20666: inst = 32'd201347077;
      20667: inst = 32'd203472343;
      20668: inst = 32'd471859200;
      20669: inst = 32'd136314880;
      20670: inst = 32'd268468224;
      20671: inst = 32'd201347078;
      20672: inst = 32'd203472343;
      20673: inst = 32'd471859200;
      20674: inst = 32'd136314880;
      20675: inst = 32'd268468224;
      20676: inst = 32'd201347079;
      20677: inst = 32'd203472343;
      20678: inst = 32'd471859200;
      20679: inst = 32'd136314880;
      20680: inst = 32'd268468224;
      20681: inst = 32'd201347080;
      20682: inst = 32'd203442761;
      20683: inst = 32'd471859200;
      20684: inst = 32'd136314880;
      20685: inst = 32'd268468224;
      20686: inst = 32'd201347081;
      20687: inst = 32'd203472343;
      20688: inst = 32'd471859200;
      20689: inst = 32'd136314880;
      20690: inst = 32'd268468224;
      20691: inst = 32'd201347082;
      20692: inst = 32'd203459697;
      20693: inst = 32'd471859200;
      20694: inst = 32'd136314880;
      20695: inst = 32'd268468224;
      20696: inst = 32'd201347083;
      20697: inst = 32'd203472343;
      20698: inst = 32'd471859200;
      20699: inst = 32'd136314880;
      20700: inst = 32'd268468224;
      20701: inst = 32'd201347084;
      20702: inst = 32'd203442761;
      20703: inst = 32'd471859200;
      20704: inst = 32'd136314880;
      20705: inst = 32'd268468224;
      20706: inst = 32'd201347085;
      20707: inst = 32'd203472343;
      20708: inst = 32'd471859200;
      20709: inst = 32'd136314880;
      20710: inst = 32'd268468224;
      20711: inst = 32'd201347086;
      20712: inst = 32'd203472343;
      20713: inst = 32'd471859200;
      20714: inst = 32'd136314880;
      20715: inst = 32'd268468224;
      20716: inst = 32'd201347087;
      20717: inst = 32'd203472343;
      20718: inst = 32'd471859200;
      20719: inst = 32'd136314880;
      20720: inst = 32'd268468224;
      20721: inst = 32'd201347088;
      20722: inst = 32'd203472343;
      20723: inst = 32'd471859200;
      20724: inst = 32'd136314880;
      20725: inst = 32'd268468224;
      20726: inst = 32'd201347089;
      20727: inst = 32'd203472343;
      20728: inst = 32'd471859200;
      20729: inst = 32'd136314880;
      20730: inst = 32'd268468224;
      20731: inst = 32'd201347090;
      20732: inst = 32'd203472343;
      20733: inst = 32'd471859200;
      20734: inst = 32'd136314880;
      20735: inst = 32'd268468224;
      20736: inst = 32'd201347091;
      20737: inst = 32'd203472343;
      20738: inst = 32'd471859200;
      20739: inst = 32'd136314880;
      20740: inst = 32'd268468224;
      20741: inst = 32'd201347092;
      20742: inst = 32'd203459697;
      20743: inst = 32'd471859200;
      20744: inst = 32'd136314880;
      20745: inst = 32'd268468224;
      20746: inst = 32'd201347093;
      20747: inst = 32'd203451245;
      20748: inst = 32'd471859200;
      20749: inst = 32'd136314880;
      20750: inst = 32'd268468224;
      20751: inst = 32'd201347094;
      20752: inst = 32'd203451245;
      20753: inst = 32'd471859200;
      20754: inst = 32'd136314880;
      20755: inst = 32'd268468224;
      20756: inst = 32'd201347095;
      20757: inst = 32'd203484854;
      20758: inst = 32'd471859200;
      20759: inst = 32'd136314880;
      20760: inst = 32'd268468224;
      20761: inst = 32'd201347096;
      20762: inst = 32'd203484854;
      20763: inst = 32'd471859200;
      20764: inst = 32'd136314880;
      20765: inst = 32'd268468224;
      20766: inst = 32'd201347097;
      20767: inst = 32'd203484854;
      20768: inst = 32'd471859200;
      20769: inst = 32'd136314880;
      20770: inst = 32'd268468224;
      20771: inst = 32'd201347098;
      20772: inst = 32'd203484854;
      20773: inst = 32'd471859200;
      20774: inst = 32'd136314880;
      20775: inst = 32'd268468224;
      20776: inst = 32'd201347099;
      20777: inst = 32'd203484854;
      20778: inst = 32'd471859200;
      20779: inst = 32'd136314880;
      20780: inst = 32'd268468224;
      20781: inst = 32'd201347100;
      20782: inst = 32'd203484854;
      20783: inst = 32'd471859200;
      20784: inst = 32'd136314880;
      20785: inst = 32'd268468224;
      20786: inst = 32'd201347101;
      20787: inst = 32'd203484854;
      20788: inst = 32'd471859200;
      20789: inst = 32'd136314880;
      20790: inst = 32'd268468224;
      20791: inst = 32'd201347102;
      20792: inst = 32'd203484854;
      20793: inst = 32'd471859200;
      20794: inst = 32'd136314880;
      20795: inst = 32'd268468224;
      20796: inst = 32'd201347103;
      20797: inst = 32'd203449101;
      20798: inst = 32'd471859200;
      20799: inst = 32'd136314880;
      20800: inst = 32'd268468224;
      20801: inst = 32'd201347104;
      20802: inst = 32'd203447021;
      20803: inst = 32'd471859200;
      20804: inst = 32'd136314880;
      20805: inst = 32'd268468224;
      20806: inst = 32'd201347105;
      20807: inst = 32'd203447021;
      20808: inst = 32'd471859200;
      20809: inst = 32'd136314880;
      20810: inst = 32'd268468224;
      20811: inst = 32'd201347106;
      20812: inst = 32'd203447021;
      20813: inst = 32'd471859200;
      20814: inst = 32'd136314880;
      20815: inst = 32'd268468224;
      20816: inst = 32'd201347107;
      20817: inst = 32'd203447021;
      20818: inst = 32'd471859200;
      20819: inst = 32'd136314880;
      20820: inst = 32'd268468224;
      20821: inst = 32'd201347108;
      20822: inst = 32'd203447020;
      20823: inst = 32'd471859200;
      20824: inst = 32'd136314880;
      20825: inst = 32'd268468224;
      20826: inst = 32'd201347109;
      20827: inst = 32'd203444841;
      20828: inst = 32'd471859200;
      20829: inst = 32'd136314880;
      20830: inst = 32'd268468224;
      20831: inst = 32'd201347110;
      20832: inst = 32'd203447021;
      20833: inst = 32'd471859200;
      20834: inst = 32'd136314880;
      20835: inst = 32'd268468224;
      20836: inst = 32'd201347111;
      20837: inst = 32'd203447021;
      20838: inst = 32'd471859200;
      20839: inst = 32'd136314880;
      20840: inst = 32'd268468224;
      20841: inst = 32'd201347112;
      20842: inst = 32'd203484854;
      20843: inst = 32'd471859200;
      20844: inst = 32'd136314880;
      20845: inst = 32'd268468224;
      20846: inst = 32'd201347113;
      20847: inst = 32'd203484854;
      20848: inst = 32'd471859200;
      20849: inst = 32'd136314880;
      20850: inst = 32'd268468224;
      20851: inst = 32'd201347114;
      20852: inst = 32'd203484854;
      20853: inst = 32'd471859200;
      20854: inst = 32'd136314880;
      20855: inst = 32'd268468224;
      20856: inst = 32'd201347115;
      20857: inst = 32'd203484854;
      20858: inst = 32'd471859200;
      20859: inst = 32'd136314880;
      20860: inst = 32'd268468224;
      20861: inst = 32'd201347116;
      20862: inst = 32'd203484854;
      20863: inst = 32'd471859200;
      20864: inst = 32'd136314880;
      20865: inst = 32'd268468224;
      20866: inst = 32'd201347117;
      20867: inst = 32'd203484854;
      20868: inst = 32'd471859200;
      20869: inst = 32'd136314880;
      20870: inst = 32'd268468224;
      20871: inst = 32'd201347118;
      20872: inst = 32'd203484854;
      20873: inst = 32'd471859200;
      20874: inst = 32'd136314880;
      20875: inst = 32'd268468224;
      20876: inst = 32'd201347119;
      20877: inst = 32'd203484854;
      20878: inst = 32'd471859200;
      20879: inst = 32'd136314880;
      20880: inst = 32'd268468224;
      20881: inst = 32'd201347120;
      20882: inst = 32'd203484854;
      20883: inst = 32'd471859200;
      20884: inst = 32'd136314880;
      20885: inst = 32'd268468224;
      20886: inst = 32'd201347121;
      20887: inst = 32'd203484854;
      20888: inst = 32'd471859200;
      20889: inst = 32'd136314880;
      20890: inst = 32'd268468224;
      20891: inst = 32'd201347122;
      20892: inst = 32'd203484854;
      20893: inst = 32'd471859200;
      20894: inst = 32'd136314880;
      20895: inst = 32'd268468224;
      20896: inst = 32'd201347123;
      20897: inst = 32'd203484854;
      20898: inst = 32'd471859200;
      20899: inst = 32'd136314880;
      20900: inst = 32'd268468224;
      20901: inst = 32'd201347124;
      20902: inst = 32'd203484854;
      20903: inst = 32'd471859200;
      20904: inst = 32'd136314880;
      20905: inst = 32'd268468224;
      20906: inst = 32'd201347125;
      20907: inst = 32'd203484854;
      20908: inst = 32'd471859200;
      20909: inst = 32'd136314880;
      20910: inst = 32'd268468224;
      20911: inst = 32'd201347126;
      20912: inst = 32'd203484854;
      20913: inst = 32'd471859200;
      20914: inst = 32'd136314880;
      20915: inst = 32'd268468224;
      20916: inst = 32'd201347127;
      20917: inst = 32'd203484854;
      20918: inst = 32'd471859200;
      20919: inst = 32'd136314880;
      20920: inst = 32'd268468224;
      20921: inst = 32'd201347128;
      20922: inst = 32'd203447021;
      20923: inst = 32'd471859200;
      20924: inst = 32'd136314880;
      20925: inst = 32'd268468224;
      20926: inst = 32'd201347129;
      20927: inst = 32'd203447021;
      20928: inst = 32'd471859200;
      20929: inst = 32'd136314880;
      20930: inst = 32'd268468224;
      20931: inst = 32'd201347130;
      20932: inst = 32'd203444841;
      20933: inst = 32'd471859200;
      20934: inst = 32'd136314880;
      20935: inst = 32'd268468224;
      20936: inst = 32'd201347131;
      20937: inst = 32'd203447020;
      20938: inst = 32'd471859200;
      20939: inst = 32'd136314880;
      20940: inst = 32'd268468224;
      20941: inst = 32'd201347132;
      20942: inst = 32'd203447021;
      20943: inst = 32'd471859200;
      20944: inst = 32'd136314880;
      20945: inst = 32'd268468224;
      20946: inst = 32'd201347133;
      20947: inst = 32'd203447021;
      20948: inst = 32'd471859200;
      20949: inst = 32'd136314880;
      20950: inst = 32'd268468224;
      20951: inst = 32'd201347134;
      20952: inst = 32'd203447021;
      20953: inst = 32'd471859200;
      20954: inst = 32'd136314880;
      20955: inst = 32'd268468224;
      20956: inst = 32'd201347135;
      20957: inst = 32'd203447021;
      20958: inst = 32'd471859200;
      20959: inst = 32'd136314880;
      20960: inst = 32'd268468224;
      20961: inst = 32'd201347136;
      20962: inst = 32'd203449101;
      20963: inst = 32'd471859200;
      20964: inst = 32'd136314880;
      20965: inst = 32'd268468224;
      20966: inst = 32'd201347137;
      20967: inst = 32'd203484854;
      20968: inst = 32'd471859200;
      20969: inst = 32'd136314880;
      20970: inst = 32'd268468224;
      20971: inst = 32'd201347138;
      20972: inst = 32'd203484854;
      20973: inst = 32'd471859200;
      20974: inst = 32'd136314880;
      20975: inst = 32'd268468224;
      20976: inst = 32'd201347139;
      20977: inst = 32'd203484854;
      20978: inst = 32'd471859200;
      20979: inst = 32'd136314880;
      20980: inst = 32'd268468224;
      20981: inst = 32'd201347140;
      20982: inst = 32'd203484854;
      20983: inst = 32'd471859200;
      20984: inst = 32'd136314880;
      20985: inst = 32'd268468224;
      20986: inst = 32'd201347141;
      20987: inst = 32'd203484854;
      20988: inst = 32'd471859200;
      20989: inst = 32'd136314880;
      20990: inst = 32'd268468224;
      20991: inst = 32'd201347142;
      20992: inst = 32'd203484854;
      20993: inst = 32'd471859200;
      20994: inst = 32'd136314880;
      20995: inst = 32'd268468224;
      20996: inst = 32'd201347143;
      20997: inst = 32'd203484854;
      20998: inst = 32'd471859200;
      20999: inst = 32'd136314880;
      21000: inst = 32'd268468224;
      21001: inst = 32'd201347144;
      21002: inst = 32'd203484854;
      21003: inst = 32'd471859200;
      21004: inst = 32'd136314880;
      21005: inst = 32'd268468224;
      21006: inst = 32'd201347145;
      21007: inst = 32'd203484854;
      21008: inst = 32'd471859200;
      21009: inst = 32'd136314880;
      21010: inst = 32'd268468224;
      21011: inst = 32'd201347146;
      21012: inst = 32'd203484854;
      21013: inst = 32'd471859200;
      21014: inst = 32'd136314880;
      21015: inst = 32'd268468224;
      21016: inst = 32'd201347147;
      21017: inst = 32'd203484854;
      21018: inst = 32'd471859200;
      21019: inst = 32'd136314880;
      21020: inst = 32'd268468224;
      21021: inst = 32'd201347148;
      21022: inst = 32'd203484854;
      21023: inst = 32'd471859200;
      21024: inst = 32'd136314880;
      21025: inst = 32'd268468224;
      21026: inst = 32'd201347149;
      21027: inst = 32'd203484854;
      21028: inst = 32'd471859200;
      21029: inst = 32'd136314880;
      21030: inst = 32'd268468224;
      21031: inst = 32'd201347150;
      21032: inst = 32'd203484854;
      21033: inst = 32'd471859200;
      21034: inst = 32'd136314880;
      21035: inst = 32'd268468224;
      21036: inst = 32'd201347151;
      21037: inst = 32'd203473634;
      21038: inst = 32'd471859200;
      21039: inst = 32'd136314880;
      21040: inst = 32'd268468224;
      21041: inst = 32'd201347152;
      21042: inst = 32'd203480005;
      21043: inst = 32'd471859200;
      21044: inst = 32'd136314880;
      21045: inst = 32'd268468224;
      21046: inst = 32'd201347153;
      21047: inst = 32'd203480005;
      21048: inst = 32'd471859200;
      21049: inst = 32'd136314880;
      21050: inst = 32'd268468224;
      21051: inst = 32'd201347154;
      21052: inst = 32'd203480005;
      21053: inst = 32'd471859200;
      21054: inst = 32'd136314880;
      21055: inst = 32'd268468224;
      21056: inst = 32'd201347155;
      21057: inst = 32'd203480005;
      21058: inst = 32'd471859200;
      21059: inst = 32'd136314880;
      21060: inst = 32'd268468224;
      21061: inst = 32'd201347156;
      21062: inst = 32'd203480005;
      21063: inst = 32'd471859200;
      21064: inst = 32'd136314880;
      21065: inst = 32'd268468224;
      21066: inst = 32'd201347157;
      21067: inst = 32'd203480005;
      21068: inst = 32'd471859200;
      21069: inst = 32'd136314880;
      21070: inst = 32'd268468224;
      21071: inst = 32'd201347158;
      21072: inst = 32'd203480005;
      21073: inst = 32'd471859200;
      21074: inst = 32'd136314880;
      21075: inst = 32'd268468224;
      21076: inst = 32'd201347159;
      21077: inst = 32'd203480005;
      21078: inst = 32'd471859200;
      21079: inst = 32'd136314880;
      21080: inst = 32'd268468224;
      21081: inst = 32'd201347160;
      21082: inst = 32'd203480005;
      21083: inst = 32'd471859200;
      21084: inst = 32'd136314880;
      21085: inst = 32'd268468224;
      21086: inst = 32'd201347161;
      21087: inst = 32'd203480005;
      21088: inst = 32'd471859200;
      21089: inst = 32'd136314880;
      21090: inst = 32'd268468224;
      21091: inst = 32'd201347162;
      21092: inst = 32'd203480005;
      21093: inst = 32'd471859200;
      21094: inst = 32'd136314880;
      21095: inst = 32'd268468224;
      21096: inst = 32'd201347163;
      21097: inst = 32'd203480005;
      21098: inst = 32'd471859200;
      21099: inst = 32'd136314880;
      21100: inst = 32'd268468224;
      21101: inst = 32'd201347164;
      21102: inst = 32'd203480005;
      21103: inst = 32'd471859200;
      21104: inst = 32'd136314880;
      21105: inst = 32'd268468224;
      21106: inst = 32'd201347165;
      21107: inst = 32'd203480005;
      21108: inst = 32'd471859200;
      21109: inst = 32'd136314880;
      21110: inst = 32'd268468224;
      21111: inst = 32'd201347166;
      21112: inst = 32'd203480005;
      21113: inst = 32'd471859200;
      21114: inst = 32'd136314880;
      21115: inst = 32'd268468224;
      21116: inst = 32'd201347167;
      21117: inst = 32'd203473634;
      21118: inst = 32'd471859200;
      21119: inst = 32'd136314880;
      21120: inst = 32'd268468224;
      21121: inst = 32'd201347168;
      21122: inst = 32'd203459697;
      21123: inst = 32'd471859200;
      21124: inst = 32'd136314880;
      21125: inst = 32'd268468224;
      21126: inst = 32'd201347169;
      21127: inst = 32'd203472343;
      21128: inst = 32'd471859200;
      21129: inst = 32'd136314880;
      21130: inst = 32'd268468224;
      21131: inst = 32'd201347170;
      21132: inst = 32'd203472343;
      21133: inst = 32'd471859200;
      21134: inst = 32'd136314880;
      21135: inst = 32'd268468224;
      21136: inst = 32'd201347171;
      21137: inst = 32'd203472343;
      21138: inst = 32'd471859200;
      21139: inst = 32'd136314880;
      21140: inst = 32'd268468224;
      21141: inst = 32'd201347172;
      21142: inst = 32'd203472343;
      21143: inst = 32'd471859200;
      21144: inst = 32'd136314880;
      21145: inst = 32'd268468224;
      21146: inst = 32'd201347173;
      21147: inst = 32'd203472343;
      21148: inst = 32'd471859200;
      21149: inst = 32'd136314880;
      21150: inst = 32'd268468224;
      21151: inst = 32'd201347174;
      21152: inst = 32'd203472343;
      21153: inst = 32'd471859200;
      21154: inst = 32'd136314880;
      21155: inst = 32'd268468224;
      21156: inst = 32'd201347175;
      21157: inst = 32'd203472343;
      21158: inst = 32'd471859200;
      21159: inst = 32'd136314880;
      21160: inst = 32'd268468224;
      21161: inst = 32'd201347176;
      21162: inst = 32'd203472343;
      21163: inst = 32'd471859200;
      21164: inst = 32'd136314880;
      21165: inst = 32'd268468224;
      21166: inst = 32'd201347177;
      21167: inst = 32'd203472343;
      21168: inst = 32'd471859200;
      21169: inst = 32'd136314880;
      21170: inst = 32'd268468224;
      21171: inst = 32'd201347178;
      21172: inst = 32'd203459697;
      21173: inst = 32'd471859200;
      21174: inst = 32'd136314880;
      21175: inst = 32'd268468224;
      21176: inst = 32'd201347179;
      21177: inst = 32'd203472343;
      21178: inst = 32'd471859200;
      21179: inst = 32'd136314880;
      21180: inst = 32'd268468224;
      21181: inst = 32'd201347180;
      21182: inst = 32'd203472343;
      21183: inst = 32'd471859200;
      21184: inst = 32'd136314880;
      21185: inst = 32'd268468224;
      21186: inst = 32'd201347181;
      21187: inst = 32'd203472343;
      21188: inst = 32'd471859200;
      21189: inst = 32'd136314880;
      21190: inst = 32'd268468224;
      21191: inst = 32'd201347182;
      21192: inst = 32'd203472343;
      21193: inst = 32'd471859200;
      21194: inst = 32'd136314880;
      21195: inst = 32'd268468224;
      21196: inst = 32'd201347183;
      21197: inst = 32'd203472343;
      21198: inst = 32'd471859200;
      21199: inst = 32'd136314880;
      21200: inst = 32'd268468224;
      21201: inst = 32'd201347184;
      21202: inst = 32'd203472343;
      21203: inst = 32'd471859200;
      21204: inst = 32'd136314880;
      21205: inst = 32'd268468224;
      21206: inst = 32'd201347185;
      21207: inst = 32'd203472343;
      21208: inst = 32'd471859200;
      21209: inst = 32'd136314880;
      21210: inst = 32'd268468224;
      21211: inst = 32'd201347186;
      21212: inst = 32'd203472343;
      21213: inst = 32'd471859200;
      21214: inst = 32'd136314880;
      21215: inst = 32'd268468224;
      21216: inst = 32'd201347187;
      21217: inst = 32'd203472343;
      21218: inst = 32'd471859200;
      21219: inst = 32'd136314880;
      21220: inst = 32'd268468224;
      21221: inst = 32'd201347188;
      21222: inst = 32'd203459697;
      21223: inst = 32'd471859200;
      21224: inst = 32'd136314880;
      21225: inst = 32'd268468224;
      21226: inst = 32'd201347189;
      21227: inst = 32'd203451245;
      21228: inst = 32'd471859200;
      21229: inst = 32'd136314880;
      21230: inst = 32'd268468224;
      21231: inst = 32'd201347190;
      21232: inst = 32'd203451245;
      21233: inst = 32'd471859200;
      21234: inst = 32'd136314880;
      21235: inst = 32'd268468224;
      21236: inst = 32'd201347191;
      21237: inst = 32'd203484854;
      21238: inst = 32'd471859200;
      21239: inst = 32'd136314880;
      21240: inst = 32'd268468224;
      21241: inst = 32'd201347192;
      21242: inst = 32'd203484854;
      21243: inst = 32'd471859200;
      21244: inst = 32'd136314880;
      21245: inst = 32'd268468224;
      21246: inst = 32'd201347193;
      21247: inst = 32'd203484854;
      21248: inst = 32'd471859200;
      21249: inst = 32'd136314880;
      21250: inst = 32'd268468224;
      21251: inst = 32'd201347194;
      21252: inst = 32'd203484854;
      21253: inst = 32'd471859200;
      21254: inst = 32'd136314880;
      21255: inst = 32'd268468224;
      21256: inst = 32'd201347195;
      21257: inst = 32'd203484854;
      21258: inst = 32'd471859200;
      21259: inst = 32'd136314880;
      21260: inst = 32'd268468224;
      21261: inst = 32'd201347196;
      21262: inst = 32'd203484854;
      21263: inst = 32'd471859200;
      21264: inst = 32'd136314880;
      21265: inst = 32'd268468224;
      21266: inst = 32'd201347197;
      21267: inst = 32'd203484854;
      21268: inst = 32'd471859200;
      21269: inst = 32'd136314880;
      21270: inst = 32'd268468224;
      21271: inst = 32'd201347198;
      21272: inst = 32'd203484854;
      21273: inst = 32'd471859200;
      21274: inst = 32'd136314880;
      21275: inst = 32'd268468224;
      21276: inst = 32'd201347199;
      21277: inst = 32'd203447021;
      21278: inst = 32'd471859200;
      21279: inst = 32'd136314880;
      21280: inst = 32'd268468224;
      21281: inst = 32'd201347200;
      21282: inst = 32'd203447021;
      21283: inst = 32'd471859200;
      21284: inst = 32'd136314880;
      21285: inst = 32'd268468224;
      21286: inst = 32'd201347201;
      21287: inst = 32'd203447021;
      21288: inst = 32'd471859200;
      21289: inst = 32'd136314880;
      21290: inst = 32'd268468224;
      21291: inst = 32'd201347202;
      21292: inst = 32'd203447021;
      21293: inst = 32'd471859200;
      21294: inst = 32'd136314880;
      21295: inst = 32'd268468224;
      21296: inst = 32'd201347203;
      21297: inst = 32'd203447020;
      21298: inst = 32'd471859200;
      21299: inst = 32'd136314880;
      21300: inst = 32'd268468224;
      21301: inst = 32'd201347204;
      21302: inst = 32'd203444874;
      21303: inst = 32'd471859200;
      21304: inst = 32'd136314880;
      21305: inst = 32'd268468224;
      21306: inst = 32'd201347205;
      21307: inst = 32'd203442793;
      21308: inst = 32'd471859200;
      21309: inst = 32'd136314880;
      21310: inst = 32'd268468224;
      21311: inst = 32'd201347206;
      21312: inst = 32'd203447021;
      21313: inst = 32'd471859200;
      21314: inst = 32'd136314880;
      21315: inst = 32'd268468224;
      21316: inst = 32'd201347207;
      21317: inst = 32'd203447021;
      21318: inst = 32'd471859200;
      21319: inst = 32'd136314880;
      21320: inst = 32'd268468224;
      21321: inst = 32'd201347208;
      21322: inst = 32'd203484854;
      21323: inst = 32'd471859200;
      21324: inst = 32'd136314880;
      21325: inst = 32'd268468224;
      21326: inst = 32'd201347209;
      21327: inst = 32'd203484854;
      21328: inst = 32'd471859200;
      21329: inst = 32'd136314880;
      21330: inst = 32'd268468224;
      21331: inst = 32'd201347210;
      21332: inst = 32'd203484854;
      21333: inst = 32'd471859200;
      21334: inst = 32'd136314880;
      21335: inst = 32'd268468224;
      21336: inst = 32'd201347211;
      21337: inst = 32'd203484854;
      21338: inst = 32'd471859200;
      21339: inst = 32'd136314880;
      21340: inst = 32'd268468224;
      21341: inst = 32'd201347212;
      21342: inst = 32'd203484854;
      21343: inst = 32'd471859200;
      21344: inst = 32'd136314880;
      21345: inst = 32'd268468224;
      21346: inst = 32'd201347213;
      21347: inst = 32'd203484854;
      21348: inst = 32'd471859200;
      21349: inst = 32'd136314880;
      21350: inst = 32'd268468224;
      21351: inst = 32'd201347214;
      21352: inst = 32'd203484854;
      21353: inst = 32'd471859200;
      21354: inst = 32'd136314880;
      21355: inst = 32'd268468224;
      21356: inst = 32'd201347215;
      21357: inst = 32'd203484854;
      21358: inst = 32'd471859200;
      21359: inst = 32'd136314880;
      21360: inst = 32'd268468224;
      21361: inst = 32'd201347216;
      21362: inst = 32'd203484854;
      21363: inst = 32'd471859200;
      21364: inst = 32'd136314880;
      21365: inst = 32'd268468224;
      21366: inst = 32'd201347217;
      21367: inst = 32'd203484854;
      21368: inst = 32'd471859200;
      21369: inst = 32'd136314880;
      21370: inst = 32'd268468224;
      21371: inst = 32'd201347218;
      21372: inst = 32'd203484854;
      21373: inst = 32'd471859200;
      21374: inst = 32'd136314880;
      21375: inst = 32'd268468224;
      21376: inst = 32'd201347219;
      21377: inst = 32'd203484854;
      21378: inst = 32'd471859200;
      21379: inst = 32'd136314880;
      21380: inst = 32'd268468224;
      21381: inst = 32'd201347220;
      21382: inst = 32'd203484854;
      21383: inst = 32'd471859200;
      21384: inst = 32'd136314880;
      21385: inst = 32'd268468224;
      21386: inst = 32'd201347221;
      21387: inst = 32'd203484854;
      21388: inst = 32'd471859200;
      21389: inst = 32'd136314880;
      21390: inst = 32'd268468224;
      21391: inst = 32'd201347222;
      21392: inst = 32'd203484854;
      21393: inst = 32'd471859200;
      21394: inst = 32'd136314880;
      21395: inst = 32'd268468224;
      21396: inst = 32'd201347223;
      21397: inst = 32'd203484854;
      21398: inst = 32'd471859200;
      21399: inst = 32'd136314880;
      21400: inst = 32'd268468224;
      21401: inst = 32'd201347224;
      21402: inst = 32'd203447021;
      21403: inst = 32'd471859200;
      21404: inst = 32'd136314880;
      21405: inst = 32'd268468224;
      21406: inst = 32'd201347225;
      21407: inst = 32'd203447021;
      21408: inst = 32'd471859200;
      21409: inst = 32'd136314880;
      21410: inst = 32'd268468224;
      21411: inst = 32'd201347226;
      21412: inst = 32'd203442793;
      21413: inst = 32'd471859200;
      21414: inst = 32'd136314880;
      21415: inst = 32'd268468224;
      21416: inst = 32'd201347227;
      21417: inst = 32'd203444874;
      21418: inst = 32'd471859200;
      21419: inst = 32'd136314880;
      21420: inst = 32'd268468224;
      21421: inst = 32'd201347228;
      21422: inst = 32'd203447020;
      21423: inst = 32'd471859200;
      21424: inst = 32'd136314880;
      21425: inst = 32'd268468224;
      21426: inst = 32'd201347229;
      21427: inst = 32'd203447021;
      21428: inst = 32'd471859200;
      21429: inst = 32'd136314880;
      21430: inst = 32'd268468224;
      21431: inst = 32'd201347230;
      21432: inst = 32'd203447021;
      21433: inst = 32'd471859200;
      21434: inst = 32'd136314880;
      21435: inst = 32'd268468224;
      21436: inst = 32'd201347231;
      21437: inst = 32'd203447021;
      21438: inst = 32'd471859200;
      21439: inst = 32'd136314880;
      21440: inst = 32'd268468224;
      21441: inst = 32'd201347232;
      21442: inst = 32'd203447021;
      21443: inst = 32'd471859200;
      21444: inst = 32'd136314880;
      21445: inst = 32'd268468224;
      21446: inst = 32'd201347233;
      21447: inst = 32'd203484854;
      21448: inst = 32'd471859200;
      21449: inst = 32'd136314880;
      21450: inst = 32'd268468224;
      21451: inst = 32'd201347234;
      21452: inst = 32'd203484854;
      21453: inst = 32'd471859200;
      21454: inst = 32'd136314880;
      21455: inst = 32'd268468224;
      21456: inst = 32'd201347235;
      21457: inst = 32'd203484854;
      21458: inst = 32'd471859200;
      21459: inst = 32'd136314880;
      21460: inst = 32'd268468224;
      21461: inst = 32'd201347236;
      21462: inst = 32'd203484854;
      21463: inst = 32'd471859200;
      21464: inst = 32'd136314880;
      21465: inst = 32'd268468224;
      21466: inst = 32'd201347237;
      21467: inst = 32'd203484854;
      21468: inst = 32'd471859200;
      21469: inst = 32'd136314880;
      21470: inst = 32'd268468224;
      21471: inst = 32'd201347238;
      21472: inst = 32'd203484854;
      21473: inst = 32'd471859200;
      21474: inst = 32'd136314880;
      21475: inst = 32'd268468224;
      21476: inst = 32'd201347239;
      21477: inst = 32'd203484854;
      21478: inst = 32'd471859200;
      21479: inst = 32'd136314880;
      21480: inst = 32'd268468224;
      21481: inst = 32'd201347240;
      21482: inst = 32'd203484854;
      21483: inst = 32'd471859200;
      21484: inst = 32'd136314880;
      21485: inst = 32'd268468224;
      21486: inst = 32'd201347241;
      21487: inst = 32'd203484854;
      21488: inst = 32'd471859200;
      21489: inst = 32'd136314880;
      21490: inst = 32'd268468224;
      21491: inst = 32'd201347242;
      21492: inst = 32'd203484854;
      21493: inst = 32'd471859200;
      21494: inst = 32'd136314880;
      21495: inst = 32'd268468224;
      21496: inst = 32'd201347243;
      21497: inst = 32'd203484854;
      21498: inst = 32'd471859200;
      21499: inst = 32'd136314880;
      21500: inst = 32'd268468224;
      21501: inst = 32'd201347244;
      21502: inst = 32'd203484854;
      21503: inst = 32'd471859200;
      21504: inst = 32'd136314880;
      21505: inst = 32'd268468224;
      21506: inst = 32'd201347245;
      21507: inst = 32'd203484854;
      21508: inst = 32'd471859200;
      21509: inst = 32'd136314880;
      21510: inst = 32'd268468224;
      21511: inst = 32'd201347246;
      21512: inst = 32'd203484854;
      21513: inst = 32'd471859200;
      21514: inst = 32'd136314880;
      21515: inst = 32'd268468224;
      21516: inst = 32'd201347247;
      21517: inst = 32'd203473634;
      21518: inst = 32'd471859200;
      21519: inst = 32'd136314880;
      21520: inst = 32'd268468224;
      21521: inst = 32'd201347248;
      21522: inst = 32'd203480005;
      21523: inst = 32'd471859200;
      21524: inst = 32'd136314880;
      21525: inst = 32'd268468224;
      21526: inst = 32'd201347249;
      21527: inst = 32'd203480005;
      21528: inst = 32'd471859200;
      21529: inst = 32'd136314880;
      21530: inst = 32'd268468224;
      21531: inst = 32'd201347250;
      21532: inst = 32'd203480005;
      21533: inst = 32'd471859200;
      21534: inst = 32'd136314880;
      21535: inst = 32'd268468224;
      21536: inst = 32'd201347251;
      21537: inst = 32'd203480005;
      21538: inst = 32'd471859200;
      21539: inst = 32'd136314880;
      21540: inst = 32'd268468224;
      21541: inst = 32'd201347252;
      21542: inst = 32'd203480005;
      21543: inst = 32'd471859200;
      21544: inst = 32'd136314880;
      21545: inst = 32'd268468224;
      21546: inst = 32'd201347253;
      21547: inst = 32'd203480005;
      21548: inst = 32'd471859200;
      21549: inst = 32'd136314880;
      21550: inst = 32'd268468224;
      21551: inst = 32'd201347254;
      21552: inst = 32'd203480005;
      21553: inst = 32'd471859200;
      21554: inst = 32'd136314880;
      21555: inst = 32'd268468224;
      21556: inst = 32'd201347255;
      21557: inst = 32'd203480005;
      21558: inst = 32'd471859200;
      21559: inst = 32'd136314880;
      21560: inst = 32'd268468224;
      21561: inst = 32'd201347256;
      21562: inst = 32'd203480005;
      21563: inst = 32'd471859200;
      21564: inst = 32'd136314880;
      21565: inst = 32'd268468224;
      21566: inst = 32'd201347257;
      21567: inst = 32'd203480005;
      21568: inst = 32'd471859200;
      21569: inst = 32'd136314880;
      21570: inst = 32'd268468224;
      21571: inst = 32'd201347258;
      21572: inst = 32'd203480005;
      21573: inst = 32'd471859200;
      21574: inst = 32'd136314880;
      21575: inst = 32'd268468224;
      21576: inst = 32'd201347259;
      21577: inst = 32'd203480005;
      21578: inst = 32'd471859200;
      21579: inst = 32'd136314880;
      21580: inst = 32'd268468224;
      21581: inst = 32'd201347260;
      21582: inst = 32'd203480005;
      21583: inst = 32'd471859200;
      21584: inst = 32'd136314880;
      21585: inst = 32'd268468224;
      21586: inst = 32'd201347261;
      21587: inst = 32'd203480005;
      21588: inst = 32'd471859200;
      21589: inst = 32'd136314880;
      21590: inst = 32'd268468224;
      21591: inst = 32'd201347262;
      21592: inst = 32'd203480005;
      21593: inst = 32'd471859200;
      21594: inst = 32'd136314880;
      21595: inst = 32'd268468224;
      21596: inst = 32'd201347263;
      21597: inst = 32'd203473634;
      21598: inst = 32'd471859200;
      21599: inst = 32'd136314880;
      21600: inst = 32'd268468224;
      21601: inst = 32'd201347264;
      21602: inst = 32'd203459697;
      21603: inst = 32'd471859200;
      21604: inst = 32'd136314880;
      21605: inst = 32'd268468224;
      21606: inst = 32'd201347265;
      21607: inst = 32'd203472343;
      21608: inst = 32'd471859200;
      21609: inst = 32'd136314880;
      21610: inst = 32'd268468224;
      21611: inst = 32'd201347266;
      21612: inst = 32'd203472343;
      21613: inst = 32'd471859200;
      21614: inst = 32'd136314880;
      21615: inst = 32'd268468224;
      21616: inst = 32'd201347267;
      21617: inst = 32'd203472343;
      21618: inst = 32'd471859200;
      21619: inst = 32'd136314880;
      21620: inst = 32'd268468224;
      21621: inst = 32'd201347268;
      21622: inst = 32'd203472343;
      21623: inst = 32'd471859200;
      21624: inst = 32'd136314880;
      21625: inst = 32'd268468224;
      21626: inst = 32'd201347269;
      21627: inst = 32'd203472343;
      21628: inst = 32'd471859200;
      21629: inst = 32'd136314880;
      21630: inst = 32'd268468224;
      21631: inst = 32'd201347270;
      21632: inst = 32'd203472343;
      21633: inst = 32'd471859200;
      21634: inst = 32'd136314880;
      21635: inst = 32'd268468224;
      21636: inst = 32'd201347271;
      21637: inst = 32'd203472343;
      21638: inst = 32'd471859200;
      21639: inst = 32'd136314880;
      21640: inst = 32'd268468224;
      21641: inst = 32'd201347272;
      21642: inst = 32'd203472343;
      21643: inst = 32'd471859200;
      21644: inst = 32'd136314880;
      21645: inst = 32'd268468224;
      21646: inst = 32'd201347273;
      21647: inst = 32'd203472343;
      21648: inst = 32'd471859200;
      21649: inst = 32'd136314880;
      21650: inst = 32'd268468224;
      21651: inst = 32'd201347274;
      21652: inst = 32'd203459697;
      21653: inst = 32'd471859200;
      21654: inst = 32'd136314880;
      21655: inst = 32'd268468224;
      21656: inst = 32'd201347275;
      21657: inst = 32'd203472343;
      21658: inst = 32'd471859200;
      21659: inst = 32'd136314880;
      21660: inst = 32'd268468224;
      21661: inst = 32'd201347276;
      21662: inst = 32'd203472343;
      21663: inst = 32'd471859200;
      21664: inst = 32'd136314880;
      21665: inst = 32'd268468224;
      21666: inst = 32'd201347277;
      21667: inst = 32'd203472343;
      21668: inst = 32'd471859200;
      21669: inst = 32'd136314880;
      21670: inst = 32'd268468224;
      21671: inst = 32'd201347278;
      21672: inst = 32'd203472343;
      21673: inst = 32'd471859200;
      21674: inst = 32'd136314880;
      21675: inst = 32'd268468224;
      21676: inst = 32'd201347279;
      21677: inst = 32'd203472343;
      21678: inst = 32'd471859200;
      21679: inst = 32'd136314880;
      21680: inst = 32'd268468224;
      21681: inst = 32'd201347280;
      21682: inst = 32'd203472343;
      21683: inst = 32'd471859200;
      21684: inst = 32'd136314880;
      21685: inst = 32'd268468224;
      21686: inst = 32'd201347281;
      21687: inst = 32'd203472343;
      21688: inst = 32'd471859200;
      21689: inst = 32'd136314880;
      21690: inst = 32'd268468224;
      21691: inst = 32'd201347282;
      21692: inst = 32'd203472343;
      21693: inst = 32'd471859200;
      21694: inst = 32'd136314880;
      21695: inst = 32'd268468224;
      21696: inst = 32'd201347283;
      21697: inst = 32'd203472343;
      21698: inst = 32'd471859200;
      21699: inst = 32'd136314880;
      21700: inst = 32'd268468224;
      21701: inst = 32'd201347284;
      21702: inst = 32'd203459697;
      21703: inst = 32'd471859200;
      21704: inst = 32'd136314880;
      21705: inst = 32'd268468224;
      21706: inst = 32'd201347285;
      21707: inst = 32'd203451245;
      21708: inst = 32'd471859200;
      21709: inst = 32'd136314880;
      21710: inst = 32'd268468224;
      21711: inst = 32'd201347286;
      21712: inst = 32'd203451245;
      21713: inst = 32'd471859200;
      21714: inst = 32'd136314880;
      21715: inst = 32'd268468224;
      21716: inst = 32'd201347287;
      21717: inst = 32'd203484854;
      21718: inst = 32'd471859200;
      21719: inst = 32'd136314880;
      21720: inst = 32'd268468224;
      21721: inst = 32'd201347288;
      21722: inst = 32'd203484854;
      21723: inst = 32'd471859200;
      21724: inst = 32'd136314880;
      21725: inst = 32'd268468224;
      21726: inst = 32'd201347289;
      21727: inst = 32'd203484854;
      21728: inst = 32'd471859200;
      21729: inst = 32'd136314880;
      21730: inst = 32'd268468224;
      21731: inst = 32'd201347290;
      21732: inst = 32'd203484854;
      21733: inst = 32'd471859200;
      21734: inst = 32'd136314880;
      21735: inst = 32'd268468224;
      21736: inst = 32'd201347291;
      21737: inst = 32'd203484854;
      21738: inst = 32'd471859200;
      21739: inst = 32'd136314880;
      21740: inst = 32'd268468224;
      21741: inst = 32'd201347292;
      21742: inst = 32'd203484854;
      21743: inst = 32'd471859200;
      21744: inst = 32'd136314880;
      21745: inst = 32'd268468224;
      21746: inst = 32'd201347293;
      21747: inst = 32'd203484854;
      21748: inst = 32'd471859200;
      21749: inst = 32'd136314880;
      21750: inst = 32'd268468224;
      21751: inst = 32'd201347294;
      21752: inst = 32'd203484854;
      21753: inst = 32'd471859200;
      21754: inst = 32'd136314880;
      21755: inst = 32'd268468224;
      21756: inst = 32'd201347295;
      21757: inst = 32'd203447021;
      21758: inst = 32'd471859200;
      21759: inst = 32'd136314880;
      21760: inst = 32'd268468224;
      21761: inst = 32'd201347296;
      21762: inst = 32'd203447021;
      21763: inst = 32'd471859200;
      21764: inst = 32'd136314880;
      21765: inst = 32'd268468224;
      21766: inst = 32'd201347297;
      21767: inst = 32'd203447021;
      21768: inst = 32'd471859200;
      21769: inst = 32'd136314880;
      21770: inst = 32'd268468224;
      21771: inst = 32'd201347298;
      21772: inst = 32'd203447021;
      21773: inst = 32'd471859200;
      21774: inst = 32'd136314880;
      21775: inst = 32'd268468224;
      21776: inst = 32'd201347299;
      21777: inst = 32'd203444874;
      21778: inst = 32'd471859200;
      21779: inst = 32'd136314880;
      21780: inst = 32'd268468224;
      21781: inst = 32'd201347300;
      21782: inst = 32'd203442793;
      21783: inst = 32'd471859200;
      21784: inst = 32'd136314880;
      21785: inst = 32'd268468224;
      21786: inst = 32'd201347301;
      21787: inst = 32'd203442793;
      21788: inst = 32'd471859200;
      21789: inst = 32'd136314880;
      21790: inst = 32'd268468224;
      21791: inst = 32'd201347302;
      21792: inst = 32'd203447021;
      21793: inst = 32'd471859200;
      21794: inst = 32'd136314880;
      21795: inst = 32'd268468224;
      21796: inst = 32'd201347303;
      21797: inst = 32'd203447021;
      21798: inst = 32'd471859200;
      21799: inst = 32'd136314880;
      21800: inst = 32'd268468224;
      21801: inst = 32'd201347304;
      21802: inst = 32'd203484854;
      21803: inst = 32'd471859200;
      21804: inst = 32'd136314880;
      21805: inst = 32'd268468224;
      21806: inst = 32'd201347305;
      21807: inst = 32'd203484854;
      21808: inst = 32'd471859200;
      21809: inst = 32'd136314880;
      21810: inst = 32'd268468224;
      21811: inst = 32'd201347306;
      21812: inst = 32'd203484854;
      21813: inst = 32'd471859200;
      21814: inst = 32'd136314880;
      21815: inst = 32'd268468224;
      21816: inst = 32'd201347307;
      21817: inst = 32'd203484854;
      21818: inst = 32'd471859200;
      21819: inst = 32'd136314880;
      21820: inst = 32'd268468224;
      21821: inst = 32'd201347308;
      21822: inst = 32'd203484854;
      21823: inst = 32'd471859200;
      21824: inst = 32'd136314880;
      21825: inst = 32'd268468224;
      21826: inst = 32'd201347309;
      21827: inst = 32'd203484854;
      21828: inst = 32'd471859200;
      21829: inst = 32'd136314880;
      21830: inst = 32'd268468224;
      21831: inst = 32'd201347310;
      21832: inst = 32'd203484854;
      21833: inst = 32'd471859200;
      21834: inst = 32'd136314880;
      21835: inst = 32'd268468224;
      21836: inst = 32'd201347311;
      21837: inst = 32'd203484854;
      21838: inst = 32'd471859200;
      21839: inst = 32'd136314880;
      21840: inst = 32'd268468224;
      21841: inst = 32'd201347312;
      21842: inst = 32'd203484854;
      21843: inst = 32'd471859200;
      21844: inst = 32'd136314880;
      21845: inst = 32'd268468224;
      21846: inst = 32'd201347313;
      21847: inst = 32'd203484854;
      21848: inst = 32'd471859200;
      21849: inst = 32'd136314880;
      21850: inst = 32'd268468224;
      21851: inst = 32'd201347314;
      21852: inst = 32'd203484854;
      21853: inst = 32'd471859200;
      21854: inst = 32'd136314880;
      21855: inst = 32'd268468224;
      21856: inst = 32'd201347315;
      21857: inst = 32'd203484854;
      21858: inst = 32'd471859200;
      21859: inst = 32'd136314880;
      21860: inst = 32'd268468224;
      21861: inst = 32'd201347316;
      21862: inst = 32'd203484854;
      21863: inst = 32'd471859200;
      21864: inst = 32'd136314880;
      21865: inst = 32'd268468224;
      21866: inst = 32'd201347317;
      21867: inst = 32'd203484854;
      21868: inst = 32'd471859200;
      21869: inst = 32'd136314880;
      21870: inst = 32'd268468224;
      21871: inst = 32'd201347318;
      21872: inst = 32'd203484854;
      21873: inst = 32'd471859200;
      21874: inst = 32'd136314880;
      21875: inst = 32'd268468224;
      21876: inst = 32'd201347319;
      21877: inst = 32'd203484854;
      21878: inst = 32'd471859200;
      21879: inst = 32'd136314880;
      21880: inst = 32'd268468224;
      21881: inst = 32'd201347320;
      21882: inst = 32'd203447021;
      21883: inst = 32'd471859200;
      21884: inst = 32'd136314880;
      21885: inst = 32'd268468224;
      21886: inst = 32'd201347321;
      21887: inst = 32'd203447021;
      21888: inst = 32'd471859200;
      21889: inst = 32'd136314880;
      21890: inst = 32'd268468224;
      21891: inst = 32'd201347322;
      21892: inst = 32'd203442793;
      21893: inst = 32'd471859200;
      21894: inst = 32'd136314880;
      21895: inst = 32'd268468224;
      21896: inst = 32'd201347323;
      21897: inst = 32'd203442793;
      21898: inst = 32'd471859200;
      21899: inst = 32'd136314880;
      21900: inst = 32'd268468224;
      21901: inst = 32'd201347324;
      21902: inst = 32'd203444874;
      21903: inst = 32'd471859200;
      21904: inst = 32'd136314880;
      21905: inst = 32'd268468224;
      21906: inst = 32'd201347325;
      21907: inst = 32'd203447021;
      21908: inst = 32'd471859200;
      21909: inst = 32'd136314880;
      21910: inst = 32'd268468224;
      21911: inst = 32'd201347326;
      21912: inst = 32'd203447021;
      21913: inst = 32'd471859200;
      21914: inst = 32'd136314880;
      21915: inst = 32'd268468224;
      21916: inst = 32'd201347327;
      21917: inst = 32'd203447021;
      21918: inst = 32'd471859200;
      21919: inst = 32'd136314880;
      21920: inst = 32'd268468224;
      21921: inst = 32'd201347328;
      21922: inst = 32'd203447021;
      21923: inst = 32'd471859200;
      21924: inst = 32'd136314880;
      21925: inst = 32'd268468224;
      21926: inst = 32'd201347329;
      21927: inst = 32'd203484854;
      21928: inst = 32'd471859200;
      21929: inst = 32'd136314880;
      21930: inst = 32'd268468224;
      21931: inst = 32'd201347330;
      21932: inst = 32'd203484854;
      21933: inst = 32'd471859200;
      21934: inst = 32'd136314880;
      21935: inst = 32'd268468224;
      21936: inst = 32'd201347331;
      21937: inst = 32'd203484854;
      21938: inst = 32'd471859200;
      21939: inst = 32'd136314880;
      21940: inst = 32'd268468224;
      21941: inst = 32'd201347332;
      21942: inst = 32'd203484854;
      21943: inst = 32'd471859200;
      21944: inst = 32'd136314880;
      21945: inst = 32'd268468224;
      21946: inst = 32'd201347333;
      21947: inst = 32'd203484854;
      21948: inst = 32'd471859200;
      21949: inst = 32'd136314880;
      21950: inst = 32'd268468224;
      21951: inst = 32'd201347334;
      21952: inst = 32'd203484854;
      21953: inst = 32'd471859200;
      21954: inst = 32'd136314880;
      21955: inst = 32'd268468224;
      21956: inst = 32'd201347335;
      21957: inst = 32'd203484854;
      21958: inst = 32'd471859200;
      21959: inst = 32'd136314880;
      21960: inst = 32'd268468224;
      21961: inst = 32'd201347336;
      21962: inst = 32'd203484854;
      21963: inst = 32'd471859200;
      21964: inst = 32'd136314880;
      21965: inst = 32'd268468224;
      21966: inst = 32'd201347337;
      21967: inst = 32'd203484854;
      21968: inst = 32'd471859200;
      21969: inst = 32'd136314880;
      21970: inst = 32'd268468224;
      21971: inst = 32'd201347338;
      21972: inst = 32'd203484854;
      21973: inst = 32'd471859200;
      21974: inst = 32'd136314880;
      21975: inst = 32'd268468224;
      21976: inst = 32'd201347339;
      21977: inst = 32'd203484854;
      21978: inst = 32'd471859200;
      21979: inst = 32'd136314880;
      21980: inst = 32'd268468224;
      21981: inst = 32'd201347340;
      21982: inst = 32'd203484854;
      21983: inst = 32'd471859200;
      21984: inst = 32'd136314880;
      21985: inst = 32'd268468224;
      21986: inst = 32'd201347341;
      21987: inst = 32'd203484854;
      21988: inst = 32'd471859200;
      21989: inst = 32'd136314880;
      21990: inst = 32'd268468224;
      21991: inst = 32'd201347342;
      21992: inst = 32'd203484854;
      21993: inst = 32'd471859200;
      21994: inst = 32'd136314880;
      21995: inst = 32'd268468224;
      21996: inst = 32'd201347343;
      21997: inst = 32'd203473634;
      21998: inst = 32'd471859200;
      21999: inst = 32'd136314880;
      22000: inst = 32'd268468224;
      22001: inst = 32'd201347344;
      22002: inst = 32'd203480005;
      22003: inst = 32'd471859200;
      22004: inst = 32'd136314880;
      22005: inst = 32'd268468224;
      22006: inst = 32'd201347345;
      22007: inst = 32'd203480005;
      22008: inst = 32'd471859200;
      22009: inst = 32'd136314880;
      22010: inst = 32'd268468224;
      22011: inst = 32'd201347346;
      22012: inst = 32'd203480005;
      22013: inst = 32'd471859200;
      22014: inst = 32'd136314880;
      22015: inst = 32'd268468224;
      22016: inst = 32'd201347347;
      22017: inst = 32'd203480005;
      22018: inst = 32'd471859200;
      22019: inst = 32'd136314880;
      22020: inst = 32'd268468224;
      22021: inst = 32'd201347348;
      22022: inst = 32'd203480005;
      22023: inst = 32'd471859200;
      22024: inst = 32'd136314880;
      22025: inst = 32'd268468224;
      22026: inst = 32'd201347349;
      22027: inst = 32'd203480005;
      22028: inst = 32'd471859200;
      22029: inst = 32'd136314880;
      22030: inst = 32'd268468224;
      22031: inst = 32'd201347350;
      22032: inst = 32'd203480005;
      22033: inst = 32'd471859200;
      22034: inst = 32'd136314880;
      22035: inst = 32'd268468224;
      22036: inst = 32'd201347351;
      22037: inst = 32'd203480005;
      22038: inst = 32'd471859200;
      22039: inst = 32'd136314880;
      22040: inst = 32'd268468224;
      22041: inst = 32'd201347352;
      22042: inst = 32'd203480005;
      22043: inst = 32'd471859200;
      22044: inst = 32'd136314880;
      22045: inst = 32'd268468224;
      22046: inst = 32'd201347353;
      22047: inst = 32'd203480005;
      22048: inst = 32'd471859200;
      22049: inst = 32'd136314880;
      22050: inst = 32'd268468224;
      22051: inst = 32'd201347354;
      22052: inst = 32'd203480005;
      22053: inst = 32'd471859200;
      22054: inst = 32'd136314880;
      22055: inst = 32'd268468224;
      22056: inst = 32'd201347355;
      22057: inst = 32'd203480005;
      22058: inst = 32'd471859200;
      22059: inst = 32'd136314880;
      22060: inst = 32'd268468224;
      22061: inst = 32'd201347356;
      22062: inst = 32'd203480005;
      22063: inst = 32'd471859200;
      22064: inst = 32'd136314880;
      22065: inst = 32'd268468224;
      22066: inst = 32'd201347357;
      22067: inst = 32'd203480005;
      22068: inst = 32'd471859200;
      22069: inst = 32'd136314880;
      22070: inst = 32'd268468224;
      22071: inst = 32'd201347358;
      22072: inst = 32'd203480005;
      22073: inst = 32'd471859200;
      22074: inst = 32'd136314880;
      22075: inst = 32'd268468224;
      22076: inst = 32'd201347359;
      22077: inst = 32'd203473634;
      22078: inst = 32'd471859200;
      22079: inst = 32'd136314880;
      22080: inst = 32'd268468224;
      22081: inst = 32'd201347360;
      22082: inst = 32'd203459697;
      22083: inst = 32'd471859200;
      22084: inst = 32'd136314880;
      22085: inst = 32'd268468224;
      22086: inst = 32'd201347361;
      22087: inst = 32'd203472343;
      22088: inst = 32'd471859200;
      22089: inst = 32'd136314880;
      22090: inst = 32'd268468224;
      22091: inst = 32'd201347362;
      22092: inst = 32'd203472343;
      22093: inst = 32'd471859200;
      22094: inst = 32'd136314880;
      22095: inst = 32'd268468224;
      22096: inst = 32'd201347363;
      22097: inst = 32'd203472343;
      22098: inst = 32'd471859200;
      22099: inst = 32'd136314880;
      22100: inst = 32'd268468224;
      22101: inst = 32'd201347364;
      22102: inst = 32'd203472343;
      22103: inst = 32'd471859200;
      22104: inst = 32'd136314880;
      22105: inst = 32'd268468224;
      22106: inst = 32'd201347365;
      22107: inst = 32'd203472343;
      22108: inst = 32'd471859200;
      22109: inst = 32'd136314880;
      22110: inst = 32'd268468224;
      22111: inst = 32'd201347366;
      22112: inst = 32'd203472343;
      22113: inst = 32'd471859200;
      22114: inst = 32'd136314880;
      22115: inst = 32'd268468224;
      22116: inst = 32'd201347367;
      22117: inst = 32'd203472343;
      22118: inst = 32'd471859200;
      22119: inst = 32'd136314880;
      22120: inst = 32'd268468224;
      22121: inst = 32'd201347368;
      22122: inst = 32'd203472343;
      22123: inst = 32'd471859200;
      22124: inst = 32'd136314880;
      22125: inst = 32'd268468224;
      22126: inst = 32'd201347369;
      22127: inst = 32'd203472343;
      22128: inst = 32'd471859200;
      22129: inst = 32'd136314880;
      22130: inst = 32'd268468224;
      22131: inst = 32'd201347370;
      22132: inst = 32'd203459697;
      22133: inst = 32'd471859200;
      22134: inst = 32'd136314880;
      22135: inst = 32'd268468224;
      22136: inst = 32'd201347371;
      22137: inst = 32'd203472343;
      22138: inst = 32'd471859200;
      22139: inst = 32'd136314880;
      22140: inst = 32'd268468224;
      22141: inst = 32'd201347372;
      22142: inst = 32'd203472343;
      22143: inst = 32'd471859200;
      22144: inst = 32'd136314880;
      22145: inst = 32'd268468224;
      22146: inst = 32'd201347373;
      22147: inst = 32'd203472343;
      22148: inst = 32'd471859200;
      22149: inst = 32'd136314880;
      22150: inst = 32'd268468224;
      22151: inst = 32'd201347374;
      22152: inst = 32'd203472343;
      22153: inst = 32'd471859200;
      22154: inst = 32'd136314880;
      22155: inst = 32'd268468224;
      22156: inst = 32'd201347375;
      22157: inst = 32'd203472343;
      22158: inst = 32'd471859200;
      22159: inst = 32'd136314880;
      22160: inst = 32'd268468224;
      22161: inst = 32'd201347376;
      22162: inst = 32'd203472343;
      22163: inst = 32'd471859200;
      22164: inst = 32'd136314880;
      22165: inst = 32'd268468224;
      22166: inst = 32'd201347377;
      22167: inst = 32'd203472343;
      22168: inst = 32'd471859200;
      22169: inst = 32'd136314880;
      22170: inst = 32'd268468224;
      22171: inst = 32'd201347378;
      22172: inst = 32'd203472343;
      22173: inst = 32'd471859200;
      22174: inst = 32'd136314880;
      22175: inst = 32'd268468224;
      22176: inst = 32'd201347379;
      22177: inst = 32'd203472343;
      22178: inst = 32'd471859200;
      22179: inst = 32'd136314880;
      22180: inst = 32'd268468224;
      22181: inst = 32'd201347380;
      22182: inst = 32'd203459697;
      22183: inst = 32'd471859200;
      22184: inst = 32'd136314880;
      22185: inst = 32'd268468224;
      22186: inst = 32'd201347381;
      22187: inst = 32'd203451245;
      22188: inst = 32'd471859200;
      22189: inst = 32'd136314880;
      22190: inst = 32'd268468224;
      22191: inst = 32'd201347382;
      22192: inst = 32'd203451245;
      22193: inst = 32'd471859200;
      22194: inst = 32'd136314880;
      22195: inst = 32'd268468224;
      22196: inst = 32'd201347383;
      22197: inst = 32'd203484854;
      22198: inst = 32'd471859200;
      22199: inst = 32'd136314880;
      22200: inst = 32'd268468224;
      22201: inst = 32'd201347384;
      22202: inst = 32'd203484854;
      22203: inst = 32'd471859200;
      22204: inst = 32'd136314880;
      22205: inst = 32'd268468224;
      22206: inst = 32'd201347385;
      22207: inst = 32'd203484854;
      22208: inst = 32'd471859200;
      22209: inst = 32'd136314880;
      22210: inst = 32'd268468224;
      22211: inst = 32'd201347386;
      22212: inst = 32'd203484854;
      22213: inst = 32'd471859200;
      22214: inst = 32'd136314880;
      22215: inst = 32'd268468224;
      22216: inst = 32'd201347387;
      22217: inst = 32'd203484854;
      22218: inst = 32'd471859200;
      22219: inst = 32'd136314880;
      22220: inst = 32'd268468224;
      22221: inst = 32'd201347388;
      22222: inst = 32'd203484854;
      22223: inst = 32'd471859200;
      22224: inst = 32'd136314880;
      22225: inst = 32'd268468224;
      22226: inst = 32'd201347389;
      22227: inst = 32'd203484854;
      22228: inst = 32'd471859200;
      22229: inst = 32'd136314880;
      22230: inst = 32'd268468224;
      22231: inst = 32'd201347390;
      22232: inst = 32'd203484854;
      22233: inst = 32'd471859200;
      22234: inst = 32'd136314880;
      22235: inst = 32'd268468224;
      22236: inst = 32'd201347391;
      22237: inst = 32'd203447021;
      22238: inst = 32'd471859200;
      22239: inst = 32'd136314880;
      22240: inst = 32'd268468224;
      22241: inst = 32'd201347392;
      22242: inst = 32'd203447021;
      22243: inst = 32'd471859200;
      22244: inst = 32'd136314880;
      22245: inst = 32'd268468224;
      22246: inst = 32'd201347393;
      22247: inst = 32'd203447021;
      22248: inst = 32'd471859200;
      22249: inst = 32'd136314880;
      22250: inst = 32'd268468224;
      22251: inst = 32'd201347394;
      22252: inst = 32'd203446955;
      22253: inst = 32'd471859200;
      22254: inst = 32'd136314880;
      22255: inst = 32'd268468224;
      22256: inst = 32'd201347395;
      22257: inst = 32'd203442793;
      22258: inst = 32'd471859200;
      22259: inst = 32'd136314880;
      22260: inst = 32'd268468224;
      22261: inst = 32'd201347396;
      22262: inst = 32'd203442793;
      22263: inst = 32'd471859200;
      22264: inst = 32'd136314880;
      22265: inst = 32'd268468224;
      22266: inst = 32'd201347397;
      22267: inst = 32'd203442793;
      22268: inst = 32'd471859200;
      22269: inst = 32'd136314880;
      22270: inst = 32'd268468224;
      22271: inst = 32'd201347398;
      22272: inst = 32'd203447021;
      22273: inst = 32'd471859200;
      22274: inst = 32'd136314880;
      22275: inst = 32'd268468224;
      22276: inst = 32'd201347399;
      22277: inst = 32'd203447021;
      22278: inst = 32'd471859200;
      22279: inst = 32'd136314880;
      22280: inst = 32'd268468224;
      22281: inst = 32'd201347400;
      22282: inst = 32'd203484854;
      22283: inst = 32'd471859200;
      22284: inst = 32'd136314880;
      22285: inst = 32'd268468224;
      22286: inst = 32'd201347401;
      22287: inst = 32'd203484854;
      22288: inst = 32'd471859200;
      22289: inst = 32'd136314880;
      22290: inst = 32'd268468224;
      22291: inst = 32'd201347402;
      22292: inst = 32'd203484854;
      22293: inst = 32'd471859200;
      22294: inst = 32'd136314880;
      22295: inst = 32'd268468224;
      22296: inst = 32'd201347403;
      22297: inst = 32'd203484854;
      22298: inst = 32'd471859200;
      22299: inst = 32'd136314880;
      22300: inst = 32'd268468224;
      22301: inst = 32'd201347404;
      22302: inst = 32'd203484854;
      22303: inst = 32'd471859200;
      22304: inst = 32'd136314880;
      22305: inst = 32'd268468224;
      22306: inst = 32'd201347405;
      22307: inst = 32'd203484854;
      22308: inst = 32'd471859200;
      22309: inst = 32'd136314880;
      22310: inst = 32'd268468224;
      22311: inst = 32'd201347406;
      22312: inst = 32'd203484854;
      22313: inst = 32'd471859200;
      22314: inst = 32'd136314880;
      22315: inst = 32'd268468224;
      22316: inst = 32'd201347407;
      22317: inst = 32'd203484854;
      22318: inst = 32'd471859200;
      22319: inst = 32'd136314880;
      22320: inst = 32'd268468224;
      22321: inst = 32'd201347408;
      22322: inst = 32'd203484854;
      22323: inst = 32'd471859200;
      22324: inst = 32'd136314880;
      22325: inst = 32'd268468224;
      22326: inst = 32'd201347409;
      22327: inst = 32'd203484854;
      22328: inst = 32'd471859200;
      22329: inst = 32'd136314880;
      22330: inst = 32'd268468224;
      22331: inst = 32'd201347410;
      22332: inst = 32'd203484854;
      22333: inst = 32'd471859200;
      22334: inst = 32'd136314880;
      22335: inst = 32'd268468224;
      22336: inst = 32'd201347411;
      22337: inst = 32'd203484854;
      22338: inst = 32'd471859200;
      22339: inst = 32'd136314880;
      22340: inst = 32'd268468224;
      22341: inst = 32'd201347412;
      22342: inst = 32'd203484854;
      22343: inst = 32'd471859200;
      22344: inst = 32'd136314880;
      22345: inst = 32'd268468224;
      22346: inst = 32'd201347413;
      22347: inst = 32'd203484854;
      22348: inst = 32'd471859200;
      22349: inst = 32'd136314880;
      22350: inst = 32'd268468224;
      22351: inst = 32'd201347414;
      22352: inst = 32'd203484854;
      22353: inst = 32'd471859200;
      22354: inst = 32'd136314880;
      22355: inst = 32'd268468224;
      22356: inst = 32'd201347415;
      22357: inst = 32'd203484854;
      22358: inst = 32'd471859200;
      22359: inst = 32'd136314880;
      22360: inst = 32'd268468224;
      22361: inst = 32'd201347416;
      22362: inst = 32'd203447021;
      22363: inst = 32'd471859200;
      22364: inst = 32'd136314880;
      22365: inst = 32'd268468224;
      22366: inst = 32'd201347417;
      22367: inst = 32'd203447021;
      22368: inst = 32'd471859200;
      22369: inst = 32'd136314880;
      22370: inst = 32'd268468224;
      22371: inst = 32'd201347418;
      22372: inst = 32'd203442793;
      22373: inst = 32'd471859200;
      22374: inst = 32'd136314880;
      22375: inst = 32'd268468224;
      22376: inst = 32'd201347419;
      22377: inst = 32'd203442793;
      22378: inst = 32'd471859200;
      22379: inst = 32'd136314880;
      22380: inst = 32'd268468224;
      22381: inst = 32'd201347420;
      22382: inst = 32'd203442793;
      22383: inst = 32'd471859200;
      22384: inst = 32'd136314880;
      22385: inst = 32'd268468224;
      22386: inst = 32'd201347421;
      22387: inst = 32'd203446955;
      22388: inst = 32'd471859200;
      22389: inst = 32'd136314880;
      22390: inst = 32'd268468224;
      22391: inst = 32'd201347422;
      22392: inst = 32'd203447021;
      22393: inst = 32'd471859200;
      22394: inst = 32'd136314880;
      22395: inst = 32'd268468224;
      22396: inst = 32'd201347423;
      22397: inst = 32'd203447021;
      22398: inst = 32'd471859200;
      22399: inst = 32'd136314880;
      22400: inst = 32'd268468224;
      22401: inst = 32'd201347424;
      22402: inst = 32'd203447021;
      22403: inst = 32'd471859200;
      22404: inst = 32'd136314880;
      22405: inst = 32'd268468224;
      22406: inst = 32'd201347425;
      22407: inst = 32'd203484854;
      22408: inst = 32'd471859200;
      22409: inst = 32'd136314880;
      22410: inst = 32'd268468224;
      22411: inst = 32'd201347426;
      22412: inst = 32'd203484854;
      22413: inst = 32'd471859200;
      22414: inst = 32'd136314880;
      22415: inst = 32'd268468224;
      22416: inst = 32'd201347427;
      22417: inst = 32'd203484854;
      22418: inst = 32'd471859200;
      22419: inst = 32'd136314880;
      22420: inst = 32'd268468224;
      22421: inst = 32'd201347428;
      22422: inst = 32'd203484854;
      22423: inst = 32'd471859200;
      22424: inst = 32'd136314880;
      22425: inst = 32'd268468224;
      22426: inst = 32'd201347429;
      22427: inst = 32'd203484854;
      22428: inst = 32'd471859200;
      22429: inst = 32'd136314880;
      22430: inst = 32'd268468224;
      22431: inst = 32'd201347430;
      22432: inst = 32'd203484854;
      22433: inst = 32'd471859200;
      22434: inst = 32'd136314880;
      22435: inst = 32'd268468224;
      22436: inst = 32'd201347431;
      22437: inst = 32'd203484854;
      22438: inst = 32'd471859200;
      22439: inst = 32'd136314880;
      22440: inst = 32'd268468224;
      22441: inst = 32'd201347432;
      22442: inst = 32'd203484854;
      22443: inst = 32'd471859200;
      22444: inst = 32'd136314880;
      22445: inst = 32'd268468224;
      22446: inst = 32'd201347433;
      22447: inst = 32'd203484854;
      22448: inst = 32'd471859200;
      22449: inst = 32'd136314880;
      22450: inst = 32'd268468224;
      22451: inst = 32'd201347434;
      22452: inst = 32'd203484854;
      22453: inst = 32'd471859200;
      22454: inst = 32'd136314880;
      22455: inst = 32'd268468224;
      22456: inst = 32'd201347435;
      22457: inst = 32'd203484854;
      22458: inst = 32'd471859200;
      22459: inst = 32'd136314880;
      22460: inst = 32'd268468224;
      22461: inst = 32'd201347436;
      22462: inst = 32'd203484854;
      22463: inst = 32'd471859200;
      22464: inst = 32'd136314880;
      22465: inst = 32'd268468224;
      22466: inst = 32'd201347437;
      22467: inst = 32'd203484854;
      22468: inst = 32'd471859200;
      22469: inst = 32'd136314880;
      22470: inst = 32'd268468224;
      22471: inst = 32'd201347438;
      22472: inst = 32'd203484854;
      22473: inst = 32'd471859200;
      22474: inst = 32'd136314880;
      22475: inst = 32'd268468224;
      22476: inst = 32'd201347439;
      22477: inst = 32'd203473634;
      22478: inst = 32'd471859200;
      22479: inst = 32'd136314880;
      22480: inst = 32'd268468224;
      22481: inst = 32'd201347440;
      22482: inst = 32'd203480005;
      22483: inst = 32'd471859200;
      22484: inst = 32'd136314880;
      22485: inst = 32'd268468224;
      22486: inst = 32'd201347441;
      22487: inst = 32'd203480005;
      22488: inst = 32'd471859200;
      22489: inst = 32'd136314880;
      22490: inst = 32'd268468224;
      22491: inst = 32'd201347442;
      22492: inst = 32'd203480005;
      22493: inst = 32'd471859200;
      22494: inst = 32'd136314880;
      22495: inst = 32'd268468224;
      22496: inst = 32'd201347443;
      22497: inst = 32'd203480005;
      22498: inst = 32'd471859200;
      22499: inst = 32'd136314880;
      22500: inst = 32'd268468224;
      22501: inst = 32'd201347444;
      22502: inst = 32'd203480005;
      22503: inst = 32'd471859200;
      22504: inst = 32'd136314880;
      22505: inst = 32'd268468224;
      22506: inst = 32'd201347445;
      22507: inst = 32'd203480005;
      22508: inst = 32'd471859200;
      22509: inst = 32'd136314880;
      22510: inst = 32'd268468224;
      22511: inst = 32'd201347446;
      22512: inst = 32'd203480005;
      22513: inst = 32'd471859200;
      22514: inst = 32'd136314880;
      22515: inst = 32'd268468224;
      22516: inst = 32'd201347447;
      22517: inst = 32'd203480005;
      22518: inst = 32'd471859200;
      22519: inst = 32'd136314880;
      22520: inst = 32'd268468224;
      22521: inst = 32'd201347448;
      22522: inst = 32'd203480005;
      22523: inst = 32'd471859200;
      22524: inst = 32'd136314880;
      22525: inst = 32'd268468224;
      22526: inst = 32'd201347449;
      22527: inst = 32'd203480005;
      22528: inst = 32'd471859200;
      22529: inst = 32'd136314880;
      22530: inst = 32'd268468224;
      22531: inst = 32'd201347450;
      22532: inst = 32'd203480005;
      22533: inst = 32'd471859200;
      22534: inst = 32'd136314880;
      22535: inst = 32'd268468224;
      22536: inst = 32'd201347451;
      22537: inst = 32'd203480005;
      22538: inst = 32'd471859200;
      22539: inst = 32'd136314880;
      22540: inst = 32'd268468224;
      22541: inst = 32'd201347452;
      22542: inst = 32'd203480005;
      22543: inst = 32'd471859200;
      22544: inst = 32'd136314880;
      22545: inst = 32'd268468224;
      22546: inst = 32'd201347453;
      22547: inst = 32'd203480005;
      22548: inst = 32'd471859200;
      22549: inst = 32'd136314880;
      22550: inst = 32'd268468224;
      22551: inst = 32'd201347454;
      22552: inst = 32'd203480005;
      22553: inst = 32'd471859200;
      22554: inst = 32'd136314880;
      22555: inst = 32'd268468224;
      22556: inst = 32'd201347455;
      22557: inst = 32'd203473634;
      22558: inst = 32'd471859200;
      22559: inst = 32'd136314880;
      22560: inst = 32'd268468224;
      22561: inst = 32'd201347456;
      22562: inst = 32'd203459697;
      22563: inst = 32'd471859200;
      22564: inst = 32'd136314880;
      22565: inst = 32'd268468224;
      22566: inst = 32'd201347457;
      22567: inst = 32'd203472343;
      22568: inst = 32'd471859200;
      22569: inst = 32'd136314880;
      22570: inst = 32'd268468224;
      22571: inst = 32'd201347458;
      22572: inst = 32'd203472343;
      22573: inst = 32'd471859200;
      22574: inst = 32'd136314880;
      22575: inst = 32'd268468224;
      22576: inst = 32'd201347459;
      22577: inst = 32'd203472343;
      22578: inst = 32'd471859200;
      22579: inst = 32'd136314880;
      22580: inst = 32'd268468224;
      22581: inst = 32'd201347460;
      22582: inst = 32'd203472343;
      22583: inst = 32'd471859200;
      22584: inst = 32'd136314880;
      22585: inst = 32'd268468224;
      22586: inst = 32'd201347461;
      22587: inst = 32'd203472343;
      22588: inst = 32'd471859200;
      22589: inst = 32'd136314880;
      22590: inst = 32'd268468224;
      22591: inst = 32'd201347462;
      22592: inst = 32'd203472343;
      22593: inst = 32'd471859200;
      22594: inst = 32'd136314880;
      22595: inst = 32'd268468224;
      22596: inst = 32'd201347463;
      22597: inst = 32'd203472343;
      22598: inst = 32'd471859200;
      22599: inst = 32'd136314880;
      22600: inst = 32'd268468224;
      22601: inst = 32'd201347464;
      22602: inst = 32'd203472343;
      22603: inst = 32'd471859200;
      22604: inst = 32'd136314880;
      22605: inst = 32'd268468224;
      22606: inst = 32'd201347465;
      22607: inst = 32'd203472343;
      22608: inst = 32'd471859200;
      22609: inst = 32'd136314880;
      22610: inst = 32'd268468224;
      22611: inst = 32'd201347466;
      22612: inst = 32'd203459697;
      22613: inst = 32'd471859200;
      22614: inst = 32'd136314880;
      22615: inst = 32'd268468224;
      22616: inst = 32'd201347467;
      22617: inst = 32'd203472343;
      22618: inst = 32'd471859200;
      22619: inst = 32'd136314880;
      22620: inst = 32'd268468224;
      22621: inst = 32'd201347468;
      22622: inst = 32'd203472343;
      22623: inst = 32'd471859200;
      22624: inst = 32'd136314880;
      22625: inst = 32'd268468224;
      22626: inst = 32'd201347469;
      22627: inst = 32'd203472343;
      22628: inst = 32'd471859200;
      22629: inst = 32'd136314880;
      22630: inst = 32'd268468224;
      22631: inst = 32'd201347470;
      22632: inst = 32'd203472343;
      22633: inst = 32'd471859200;
      22634: inst = 32'd136314880;
      22635: inst = 32'd268468224;
      22636: inst = 32'd201347471;
      22637: inst = 32'd203472343;
      22638: inst = 32'd471859200;
      22639: inst = 32'd136314880;
      22640: inst = 32'd268468224;
      22641: inst = 32'd201347472;
      22642: inst = 32'd203472343;
      22643: inst = 32'd471859200;
      22644: inst = 32'd136314880;
      22645: inst = 32'd268468224;
      22646: inst = 32'd201347473;
      22647: inst = 32'd203472343;
      22648: inst = 32'd471859200;
      22649: inst = 32'd136314880;
      22650: inst = 32'd268468224;
      22651: inst = 32'd201347474;
      22652: inst = 32'd203472343;
      22653: inst = 32'd471859200;
      22654: inst = 32'd136314880;
      22655: inst = 32'd268468224;
      22656: inst = 32'd201347475;
      22657: inst = 32'd203472343;
      22658: inst = 32'd471859200;
      22659: inst = 32'd136314880;
      22660: inst = 32'd268468224;
      22661: inst = 32'd201347476;
      22662: inst = 32'd203459697;
      22663: inst = 32'd471859200;
      22664: inst = 32'd136314880;
      22665: inst = 32'd268468224;
      22666: inst = 32'd201347477;
      22667: inst = 32'd203451245;
      22668: inst = 32'd471859200;
      22669: inst = 32'd136314880;
      22670: inst = 32'd268468224;
      22671: inst = 32'd201347478;
      22672: inst = 32'd203451245;
      22673: inst = 32'd471859200;
      22674: inst = 32'd136314880;
      22675: inst = 32'd268468224;
      22676: inst = 32'd201347479;
      22677: inst = 32'd203484854;
      22678: inst = 32'd471859200;
      22679: inst = 32'd136314880;
      22680: inst = 32'd268468224;
      22681: inst = 32'd201347480;
      22682: inst = 32'd203484854;
      22683: inst = 32'd471859200;
      22684: inst = 32'd136314880;
      22685: inst = 32'd268468224;
      22686: inst = 32'd201347481;
      22687: inst = 32'd203484854;
      22688: inst = 32'd471859200;
      22689: inst = 32'd136314880;
      22690: inst = 32'd268468224;
      22691: inst = 32'd201347482;
      22692: inst = 32'd203484854;
      22693: inst = 32'd471859200;
      22694: inst = 32'd136314880;
      22695: inst = 32'd268468224;
      22696: inst = 32'd201347483;
      22697: inst = 32'd203484854;
      22698: inst = 32'd471859200;
      22699: inst = 32'd136314880;
      22700: inst = 32'd268468224;
      22701: inst = 32'd201347484;
      22702: inst = 32'd203484854;
      22703: inst = 32'd471859200;
      22704: inst = 32'd136314880;
      22705: inst = 32'd268468224;
      22706: inst = 32'd201347485;
      22707: inst = 32'd203484854;
      22708: inst = 32'd471859200;
      22709: inst = 32'd136314880;
      22710: inst = 32'd268468224;
      22711: inst = 32'd201347486;
      22712: inst = 32'd203476436;
      22713: inst = 32'd471859200;
      22714: inst = 32'd136314880;
      22715: inst = 32'd268468224;
      22716: inst = 32'd201347487;
      22717: inst = 32'd203447021;
      22718: inst = 32'd471859200;
      22719: inst = 32'd136314880;
      22720: inst = 32'd268468224;
      22721: inst = 32'd201347488;
      22722: inst = 32'd203447021;
      22723: inst = 32'd471859200;
      22724: inst = 32'd136314880;
      22725: inst = 32'd268468224;
      22726: inst = 32'd201347489;
      22727: inst = 32'd203447020;
      22728: inst = 32'd471859200;
      22729: inst = 32'd136314880;
      22730: inst = 32'd268468224;
      22731: inst = 32'd201347490;
      22732: inst = 32'd203442793;
      22733: inst = 32'd471859200;
      22734: inst = 32'd136314880;
      22735: inst = 32'd268468224;
      22736: inst = 32'd201347491;
      22737: inst = 32'd203442793;
      22738: inst = 32'd471859200;
      22739: inst = 32'd136314880;
      22740: inst = 32'd268468224;
      22741: inst = 32'd201347492;
      22742: inst = 32'd203442793;
      22743: inst = 32'd471859200;
      22744: inst = 32'd136314880;
      22745: inst = 32'd268468224;
      22746: inst = 32'd201347493;
      22747: inst = 32'd203442793;
      22748: inst = 32'd471859200;
      22749: inst = 32'd136314880;
      22750: inst = 32'd268468224;
      22751: inst = 32'd201347494;
      22752: inst = 32'd203447021;
      22753: inst = 32'd471859200;
      22754: inst = 32'd136314880;
      22755: inst = 32'd268468224;
      22756: inst = 32'd201347495;
      22757: inst = 32'd203447021;
      22758: inst = 32'd471859200;
      22759: inst = 32'd136314880;
      22760: inst = 32'd268468224;
      22761: inst = 32'd201347496;
      22762: inst = 32'd203459697;
      22763: inst = 32'd471859200;
      22764: inst = 32'd136314880;
      22765: inst = 32'd268468224;
      22766: inst = 32'd201347497;
      22767: inst = 32'd203459697;
      22768: inst = 32'd471859200;
      22769: inst = 32'd136314880;
      22770: inst = 32'd268468224;
      22771: inst = 32'd201347498;
      22772: inst = 32'd203484854;
      22773: inst = 32'd471859200;
      22774: inst = 32'd136314880;
      22775: inst = 32'd268468224;
      22776: inst = 32'd201347499;
      22777: inst = 32'd203484854;
      22778: inst = 32'd471859200;
      22779: inst = 32'd136314880;
      22780: inst = 32'd268468224;
      22781: inst = 32'd201347500;
      22782: inst = 32'd203484854;
      22783: inst = 32'd471859200;
      22784: inst = 32'd136314880;
      22785: inst = 32'd268468224;
      22786: inst = 32'd201347501;
      22787: inst = 32'd203484854;
      22788: inst = 32'd471859200;
      22789: inst = 32'd136314880;
      22790: inst = 32'd268468224;
      22791: inst = 32'd201347502;
      22792: inst = 32'd203484854;
      22793: inst = 32'd471859200;
      22794: inst = 32'd136314880;
      22795: inst = 32'd268468224;
      22796: inst = 32'd201347503;
      22797: inst = 32'd203484854;
      22798: inst = 32'd471859200;
      22799: inst = 32'd136314880;
      22800: inst = 32'd268468224;
      22801: inst = 32'd201347504;
      22802: inst = 32'd203484854;
      22803: inst = 32'd471859200;
      22804: inst = 32'd136314880;
      22805: inst = 32'd268468224;
      22806: inst = 32'd201347505;
      22807: inst = 32'd203484854;
      22808: inst = 32'd471859200;
      22809: inst = 32'd136314880;
      22810: inst = 32'd268468224;
      22811: inst = 32'd201347506;
      22812: inst = 32'd203484854;
      22813: inst = 32'd471859200;
      22814: inst = 32'd136314880;
      22815: inst = 32'd268468224;
      22816: inst = 32'd201347507;
      22817: inst = 32'd203484854;
      22818: inst = 32'd471859200;
      22819: inst = 32'd136314880;
      22820: inst = 32'd268468224;
      22821: inst = 32'd201347508;
      22822: inst = 32'd203484854;
      22823: inst = 32'd471859200;
      22824: inst = 32'd136314880;
      22825: inst = 32'd268468224;
      22826: inst = 32'd201347509;
      22827: inst = 32'd203484854;
      22828: inst = 32'd471859200;
      22829: inst = 32'd136314880;
      22830: inst = 32'd268468224;
      22831: inst = 32'd201347510;
      22832: inst = 32'd203461745;
      22833: inst = 32'd471859200;
      22834: inst = 32'd136314880;
      22835: inst = 32'd268468224;
      22836: inst = 32'd201347511;
      22837: inst = 32'd203459697;
      22838: inst = 32'd471859200;
      22839: inst = 32'd136314880;
      22840: inst = 32'd268468224;
      22841: inst = 32'd201347512;
      22842: inst = 32'd203447021;
      22843: inst = 32'd471859200;
      22844: inst = 32'd136314880;
      22845: inst = 32'd268468224;
      22846: inst = 32'd201347513;
      22847: inst = 32'd203447021;
      22848: inst = 32'd471859200;
      22849: inst = 32'd136314880;
      22850: inst = 32'd268468224;
      22851: inst = 32'd201347514;
      22852: inst = 32'd203442793;
      22853: inst = 32'd471859200;
      22854: inst = 32'd136314880;
      22855: inst = 32'd268468224;
      22856: inst = 32'd201347515;
      22857: inst = 32'd203442793;
      22858: inst = 32'd471859200;
      22859: inst = 32'd136314880;
      22860: inst = 32'd268468224;
      22861: inst = 32'd201347516;
      22862: inst = 32'd203442793;
      22863: inst = 32'd471859200;
      22864: inst = 32'd136314880;
      22865: inst = 32'd268468224;
      22866: inst = 32'd201347517;
      22867: inst = 32'd203442793;
      22868: inst = 32'd471859200;
      22869: inst = 32'd136314880;
      22870: inst = 32'd268468224;
      22871: inst = 32'd201347518;
      22872: inst = 32'd203447020;
      22873: inst = 32'd471859200;
      22874: inst = 32'd136314880;
      22875: inst = 32'd268468224;
      22876: inst = 32'd201347519;
      22877: inst = 32'd203447021;
      22878: inst = 32'd471859200;
      22879: inst = 32'd136314880;
      22880: inst = 32'd268468224;
      22881: inst = 32'd201347520;
      22882: inst = 32'd203447021;
      22883: inst = 32'd471859200;
      22884: inst = 32'd136314880;
      22885: inst = 32'd268468224;
      22886: inst = 32'd201347521;
      22887: inst = 32'd203476436;
      22888: inst = 32'd471859200;
      22889: inst = 32'd136314880;
      22890: inst = 32'd268468224;
      22891: inst = 32'd201347522;
      22892: inst = 32'd203484854;
      22893: inst = 32'd471859200;
      22894: inst = 32'd136314880;
      22895: inst = 32'd268468224;
      22896: inst = 32'd201347523;
      22897: inst = 32'd203484854;
      22898: inst = 32'd471859200;
      22899: inst = 32'd136314880;
      22900: inst = 32'd268468224;
      22901: inst = 32'd201347524;
      22902: inst = 32'd203484854;
      22903: inst = 32'd471859200;
      22904: inst = 32'd136314880;
      22905: inst = 32'd268468224;
      22906: inst = 32'd201347525;
      22907: inst = 32'd203484854;
      22908: inst = 32'd471859200;
      22909: inst = 32'd136314880;
      22910: inst = 32'd268468224;
      22911: inst = 32'd201347526;
      22912: inst = 32'd203484854;
      22913: inst = 32'd471859200;
      22914: inst = 32'd136314880;
      22915: inst = 32'd268468224;
      22916: inst = 32'd201347527;
      22917: inst = 32'd203484854;
      22918: inst = 32'd471859200;
      22919: inst = 32'd136314880;
      22920: inst = 32'd268468224;
      22921: inst = 32'd201347528;
      22922: inst = 32'd203484854;
      22923: inst = 32'd471859200;
      22924: inst = 32'd136314880;
      22925: inst = 32'd268468224;
      22926: inst = 32'd201347529;
      22927: inst = 32'd203484854;
      22928: inst = 32'd471859200;
      22929: inst = 32'd136314880;
      22930: inst = 32'd268468224;
      22931: inst = 32'd201347530;
      22932: inst = 32'd203484854;
      22933: inst = 32'd471859200;
      22934: inst = 32'd136314880;
      22935: inst = 32'd268468224;
      22936: inst = 32'd201347531;
      22937: inst = 32'd203484854;
      22938: inst = 32'd471859200;
      22939: inst = 32'd136314880;
      22940: inst = 32'd268468224;
      22941: inst = 32'd201347532;
      22942: inst = 32'd203484854;
      22943: inst = 32'd471859200;
      22944: inst = 32'd136314880;
      22945: inst = 32'd268468224;
      22946: inst = 32'd201347533;
      22947: inst = 32'd203484854;
      22948: inst = 32'd471859200;
      22949: inst = 32'd136314880;
      22950: inst = 32'd268468224;
      22951: inst = 32'd201347534;
      22952: inst = 32'd203484854;
      22953: inst = 32'd471859200;
      22954: inst = 32'd136314880;
      22955: inst = 32'd268468224;
      22956: inst = 32'd201347535;
      22957: inst = 32'd203473634;
      22958: inst = 32'd471859200;
      22959: inst = 32'd136314880;
      22960: inst = 32'd268468224;
      22961: inst = 32'd201347536;
      22962: inst = 32'd203480005;
      22963: inst = 32'd471859200;
      22964: inst = 32'd136314880;
      22965: inst = 32'd268468224;
      22966: inst = 32'd201347537;
      22967: inst = 32'd203480005;
      22968: inst = 32'd471859200;
      22969: inst = 32'd136314880;
      22970: inst = 32'd268468224;
      22971: inst = 32'd201347538;
      22972: inst = 32'd203480005;
      22973: inst = 32'd471859200;
      22974: inst = 32'd136314880;
      22975: inst = 32'd268468224;
      22976: inst = 32'd201347539;
      22977: inst = 32'd203480005;
      22978: inst = 32'd471859200;
      22979: inst = 32'd136314880;
      22980: inst = 32'd268468224;
      22981: inst = 32'd201347540;
      22982: inst = 32'd203480005;
      22983: inst = 32'd471859200;
      22984: inst = 32'd136314880;
      22985: inst = 32'd268468224;
      22986: inst = 32'd201347541;
      22987: inst = 32'd203480005;
      22988: inst = 32'd471859200;
      22989: inst = 32'd136314880;
      22990: inst = 32'd268468224;
      22991: inst = 32'd201347542;
      22992: inst = 32'd203480005;
      22993: inst = 32'd471859200;
      22994: inst = 32'd136314880;
      22995: inst = 32'd268468224;
      22996: inst = 32'd201347543;
      22997: inst = 32'd203480005;
      22998: inst = 32'd471859200;
      22999: inst = 32'd136314880;
      23000: inst = 32'd268468224;
      23001: inst = 32'd201347544;
      23002: inst = 32'd203480005;
      23003: inst = 32'd471859200;
      23004: inst = 32'd136314880;
      23005: inst = 32'd268468224;
      23006: inst = 32'd201347545;
      23007: inst = 32'd203480005;
      23008: inst = 32'd471859200;
      23009: inst = 32'd136314880;
      23010: inst = 32'd268468224;
      23011: inst = 32'd201347546;
      23012: inst = 32'd203480005;
      23013: inst = 32'd471859200;
      23014: inst = 32'd136314880;
      23015: inst = 32'd268468224;
      23016: inst = 32'd201347547;
      23017: inst = 32'd203480005;
      23018: inst = 32'd471859200;
      23019: inst = 32'd136314880;
      23020: inst = 32'd268468224;
      23021: inst = 32'd201347548;
      23022: inst = 32'd203480005;
      23023: inst = 32'd471859200;
      23024: inst = 32'd136314880;
      23025: inst = 32'd268468224;
      23026: inst = 32'd201347549;
      23027: inst = 32'd203480005;
      23028: inst = 32'd471859200;
      23029: inst = 32'd136314880;
      23030: inst = 32'd268468224;
      23031: inst = 32'd201347550;
      23032: inst = 32'd203480005;
      23033: inst = 32'd471859200;
      23034: inst = 32'd136314880;
      23035: inst = 32'd268468224;
      23036: inst = 32'd201347551;
      23037: inst = 32'd203473634;
      23038: inst = 32'd471859200;
      23039: inst = 32'd136314880;
      23040: inst = 32'd268468224;
      23041: inst = 32'd201347552;
      23042: inst = 32'd203459697;
      23043: inst = 32'd471859200;
      23044: inst = 32'd136314880;
      23045: inst = 32'd268468224;
      23046: inst = 32'd201347553;
      23047: inst = 32'd203472343;
      23048: inst = 32'd471859200;
      23049: inst = 32'd136314880;
      23050: inst = 32'd268468224;
      23051: inst = 32'd201347554;
      23052: inst = 32'd203472343;
      23053: inst = 32'd471859200;
      23054: inst = 32'd136314880;
      23055: inst = 32'd268468224;
      23056: inst = 32'd201347555;
      23057: inst = 32'd203472343;
      23058: inst = 32'd471859200;
      23059: inst = 32'd136314880;
      23060: inst = 32'd268468224;
      23061: inst = 32'd201347556;
      23062: inst = 32'd203472343;
      23063: inst = 32'd471859200;
      23064: inst = 32'd136314880;
      23065: inst = 32'd268468224;
      23066: inst = 32'd201347557;
      23067: inst = 32'd203472343;
      23068: inst = 32'd471859200;
      23069: inst = 32'd136314880;
      23070: inst = 32'd268468224;
      23071: inst = 32'd201347558;
      23072: inst = 32'd203472343;
      23073: inst = 32'd471859200;
      23074: inst = 32'd136314880;
      23075: inst = 32'd268468224;
      23076: inst = 32'd201347559;
      23077: inst = 32'd203472343;
      23078: inst = 32'd471859200;
      23079: inst = 32'd136314880;
      23080: inst = 32'd268468224;
      23081: inst = 32'd201347560;
      23082: inst = 32'd203472343;
      23083: inst = 32'd471859200;
      23084: inst = 32'd136314880;
      23085: inst = 32'd268468224;
      23086: inst = 32'd201347561;
      23087: inst = 32'd203472343;
      23088: inst = 32'd471859200;
      23089: inst = 32'd136314880;
      23090: inst = 32'd268468224;
      23091: inst = 32'd201347562;
      23092: inst = 32'd203459697;
      23093: inst = 32'd471859200;
      23094: inst = 32'd136314880;
      23095: inst = 32'd268468224;
      23096: inst = 32'd201347563;
      23097: inst = 32'd203472343;
      23098: inst = 32'd471859200;
      23099: inst = 32'd136314880;
      23100: inst = 32'd268468224;
      23101: inst = 32'd201347564;
      23102: inst = 32'd203472343;
      23103: inst = 32'd471859200;
      23104: inst = 32'd136314880;
      23105: inst = 32'd268468224;
      23106: inst = 32'd201347565;
      23107: inst = 32'd203472343;
      23108: inst = 32'd471859200;
      23109: inst = 32'd136314880;
      23110: inst = 32'd268468224;
      23111: inst = 32'd201347566;
      23112: inst = 32'd203472343;
      23113: inst = 32'd471859200;
      23114: inst = 32'd136314880;
      23115: inst = 32'd268468224;
      23116: inst = 32'd201347567;
      23117: inst = 32'd203472343;
      23118: inst = 32'd471859200;
      23119: inst = 32'd136314880;
      23120: inst = 32'd268468224;
      23121: inst = 32'd201347568;
      23122: inst = 32'd203472343;
      23123: inst = 32'd471859200;
      23124: inst = 32'd136314880;
      23125: inst = 32'd268468224;
      23126: inst = 32'd201347569;
      23127: inst = 32'd203472343;
      23128: inst = 32'd471859200;
      23129: inst = 32'd136314880;
      23130: inst = 32'd268468224;
      23131: inst = 32'd201347570;
      23132: inst = 32'd203472343;
      23133: inst = 32'd471859200;
      23134: inst = 32'd136314880;
      23135: inst = 32'd268468224;
      23136: inst = 32'd201347571;
      23137: inst = 32'd203472343;
      23138: inst = 32'd471859200;
      23139: inst = 32'd136314880;
      23140: inst = 32'd268468224;
      23141: inst = 32'd201347572;
      23142: inst = 32'd203459697;
      23143: inst = 32'd471859200;
      23144: inst = 32'd136314880;
      23145: inst = 32'd268468224;
      23146: inst = 32'd201347573;
      23147: inst = 32'd203451245;
      23148: inst = 32'd471859200;
      23149: inst = 32'd136314880;
      23150: inst = 32'd268468224;
      23151: inst = 32'd201347574;
      23152: inst = 32'd203451245;
      23153: inst = 32'd471859200;
      23154: inst = 32'd136314880;
      23155: inst = 32'd268468224;
      23156: inst = 32'd201347575;
      23157: inst = 32'd203484854;
      23158: inst = 32'd471859200;
      23159: inst = 32'd136314880;
      23160: inst = 32'd268468224;
      23161: inst = 32'd201347576;
      23162: inst = 32'd203484854;
      23163: inst = 32'd471859200;
      23164: inst = 32'd136314880;
      23165: inst = 32'd268468224;
      23166: inst = 32'd201347577;
      23167: inst = 32'd203484854;
      23168: inst = 32'd471859200;
      23169: inst = 32'd136314880;
      23170: inst = 32'd268468224;
      23171: inst = 32'd201347578;
      23172: inst = 32'd203484854;
      23173: inst = 32'd471859200;
      23174: inst = 32'd136314880;
      23175: inst = 32'd268468224;
      23176: inst = 32'd201347579;
      23177: inst = 32'd203484854;
      23178: inst = 32'd471859200;
      23179: inst = 32'd136314880;
      23180: inst = 32'd268468224;
      23181: inst = 32'd201347580;
      23182: inst = 32'd203484854;
      23183: inst = 32'd471859200;
      23184: inst = 32'd136314880;
      23185: inst = 32'd268468224;
      23186: inst = 32'd201347581;
      23187: inst = 32'd203480661;
      23188: inst = 32'd471859200;
      23189: inst = 32'd136314880;
      23190: inst = 32'd268468224;
      23191: inst = 32'd201347582;
      23192: inst = 32'd203461778;
      23193: inst = 32'd471859200;
      23194: inst = 32'd136314880;
      23195: inst = 32'd268468224;
      23196: inst = 32'd201347583;
      23197: inst = 32'd203447021;
      23198: inst = 32'd471859200;
      23199: inst = 32'd136314880;
      23200: inst = 32'd268468224;
      23201: inst = 32'd201347584;
      23202: inst = 32'd203447021;
      23203: inst = 32'd471859200;
      23204: inst = 32'd136314880;
      23205: inst = 32'd268468224;
      23206: inst = 32'd201347585;
      23207: inst = 32'd203446988;
      23208: inst = 32'd471859200;
      23209: inst = 32'd136314880;
      23210: inst = 32'd268468224;
      23211: inst = 32'd201347586;
      23212: inst = 32'd203442793;
      23213: inst = 32'd471859200;
      23214: inst = 32'd136314880;
      23215: inst = 32'd268468224;
      23216: inst = 32'd201347587;
      23217: inst = 32'd203442793;
      23218: inst = 32'd471859200;
      23219: inst = 32'd136314880;
      23220: inst = 32'd268468224;
      23221: inst = 32'd201347588;
      23222: inst = 32'd203442793;
      23223: inst = 32'd471859200;
      23224: inst = 32'd136314880;
      23225: inst = 32'd268468224;
      23226: inst = 32'd201347589;
      23227: inst = 32'd203442793;
      23228: inst = 32'd471859200;
      23229: inst = 32'd136314880;
      23230: inst = 32'd268468224;
      23231: inst = 32'd201347590;
      23232: inst = 32'd203447021;
      23233: inst = 32'd471859200;
      23234: inst = 32'd136314880;
      23235: inst = 32'd268468224;
      23236: inst = 32'd201347591;
      23237: inst = 32'd203447021;
      23238: inst = 32'd471859200;
      23239: inst = 32'd136314880;
      23240: inst = 32'd268468224;
      23241: inst = 32'd201347592;
      23242: inst = 32'd203459697;
      23243: inst = 32'd471859200;
      23244: inst = 32'd136314880;
      23245: inst = 32'd268468224;
      23246: inst = 32'd201347593;
      23247: inst = 32'd203461712;
      23248: inst = 32'd471859200;
      23249: inst = 32'd136314880;
      23250: inst = 32'd268468224;
      23251: inst = 32'd201347594;
      23252: inst = 32'd203484854;
      23253: inst = 32'd471859200;
      23254: inst = 32'd136314880;
      23255: inst = 32'd268468224;
      23256: inst = 32'd201347595;
      23257: inst = 32'd203484854;
      23258: inst = 32'd471859200;
      23259: inst = 32'd136314880;
      23260: inst = 32'd268468224;
      23261: inst = 32'd201347596;
      23262: inst = 32'd203484854;
      23263: inst = 32'd471859200;
      23264: inst = 32'd136314880;
      23265: inst = 32'd268468224;
      23266: inst = 32'd201347597;
      23267: inst = 32'd203484854;
      23268: inst = 32'd471859200;
      23269: inst = 32'd136314880;
      23270: inst = 32'd268468224;
      23271: inst = 32'd201347598;
      23272: inst = 32'd203484854;
      23273: inst = 32'd471859200;
      23274: inst = 32'd136314880;
      23275: inst = 32'd268468224;
      23276: inst = 32'd201347599;
      23277: inst = 32'd203484854;
      23278: inst = 32'd471859200;
      23279: inst = 32'd136314880;
      23280: inst = 32'd268468224;
      23281: inst = 32'd201347600;
      23282: inst = 32'd203484854;
      23283: inst = 32'd471859200;
      23284: inst = 32'd136314880;
      23285: inst = 32'd268468224;
      23286: inst = 32'd201347601;
      23287: inst = 32'd203484854;
      23288: inst = 32'd471859200;
      23289: inst = 32'd136314880;
      23290: inst = 32'd268468224;
      23291: inst = 32'd201347602;
      23292: inst = 32'd203484854;
      23293: inst = 32'd471859200;
      23294: inst = 32'd136314880;
      23295: inst = 32'd268468224;
      23296: inst = 32'd201347603;
      23297: inst = 32'd203484854;
      23298: inst = 32'd471859200;
      23299: inst = 32'd136314880;
      23300: inst = 32'd268468224;
      23301: inst = 32'd201347604;
      23302: inst = 32'd203484854;
      23303: inst = 32'd471859200;
      23304: inst = 32'd136314880;
      23305: inst = 32'd268468224;
      23306: inst = 32'd201347605;
      23307: inst = 32'd203484854;
      23308: inst = 32'd471859200;
      23309: inst = 32'd136314880;
      23310: inst = 32'd268468224;
      23311: inst = 32'd201347606;
      23312: inst = 32'd203461712;
      23313: inst = 32'd471859200;
      23314: inst = 32'd136314880;
      23315: inst = 32'd268468224;
      23316: inst = 32'd201347607;
      23317: inst = 32'd203459697;
      23318: inst = 32'd471859200;
      23319: inst = 32'd136314880;
      23320: inst = 32'd268468224;
      23321: inst = 32'd201347608;
      23322: inst = 32'd203447021;
      23323: inst = 32'd471859200;
      23324: inst = 32'd136314880;
      23325: inst = 32'd268468224;
      23326: inst = 32'd201347609;
      23327: inst = 32'd203447021;
      23328: inst = 32'd471859200;
      23329: inst = 32'd136314880;
      23330: inst = 32'd268468224;
      23331: inst = 32'd201347610;
      23332: inst = 32'd203442793;
      23333: inst = 32'd471859200;
      23334: inst = 32'd136314880;
      23335: inst = 32'd268468224;
      23336: inst = 32'd201347611;
      23337: inst = 32'd203442793;
      23338: inst = 32'd471859200;
      23339: inst = 32'd136314880;
      23340: inst = 32'd268468224;
      23341: inst = 32'd201347612;
      23342: inst = 32'd203442793;
      23343: inst = 32'd471859200;
      23344: inst = 32'd136314880;
      23345: inst = 32'd268468224;
      23346: inst = 32'd201347613;
      23347: inst = 32'd203442793;
      23348: inst = 32'd471859200;
      23349: inst = 32'd136314880;
      23350: inst = 32'd268468224;
      23351: inst = 32'd201347614;
      23352: inst = 32'd203446988;
      23353: inst = 32'd471859200;
      23354: inst = 32'd136314880;
      23355: inst = 32'd268468224;
      23356: inst = 32'd201347615;
      23357: inst = 32'd203447021;
      23358: inst = 32'd471859200;
      23359: inst = 32'd136314880;
      23360: inst = 32'd268468224;
      23361: inst = 32'd201347616;
      23362: inst = 32'd203447021;
      23363: inst = 32'd471859200;
      23364: inst = 32'd136314880;
      23365: inst = 32'd268468224;
      23366: inst = 32'd201347617;
      23367: inst = 32'd203461778;
      23368: inst = 32'd471859200;
      23369: inst = 32'd136314880;
      23370: inst = 32'd268468224;
      23371: inst = 32'd201347618;
      23372: inst = 32'd203480661;
      23373: inst = 32'd471859200;
      23374: inst = 32'd136314880;
      23375: inst = 32'd268468224;
      23376: inst = 32'd201347619;
      23377: inst = 32'd203484854;
      23378: inst = 32'd471859200;
      23379: inst = 32'd136314880;
      23380: inst = 32'd268468224;
      23381: inst = 32'd201347620;
      23382: inst = 32'd203484854;
      23383: inst = 32'd471859200;
      23384: inst = 32'd136314880;
      23385: inst = 32'd268468224;
      23386: inst = 32'd201347621;
      23387: inst = 32'd203484854;
      23388: inst = 32'd471859200;
      23389: inst = 32'd136314880;
      23390: inst = 32'd268468224;
      23391: inst = 32'd201347622;
      23392: inst = 32'd203484854;
      23393: inst = 32'd471859200;
      23394: inst = 32'd136314880;
      23395: inst = 32'd268468224;
      23396: inst = 32'd201347623;
      23397: inst = 32'd203484854;
      23398: inst = 32'd471859200;
      23399: inst = 32'd136314880;
      23400: inst = 32'd268468224;
      23401: inst = 32'd201347624;
      23402: inst = 32'd203484854;
      23403: inst = 32'd471859200;
      23404: inst = 32'd136314880;
      23405: inst = 32'd268468224;
      23406: inst = 32'd201347625;
      23407: inst = 32'd203484854;
      23408: inst = 32'd471859200;
      23409: inst = 32'd136314880;
      23410: inst = 32'd268468224;
      23411: inst = 32'd201347626;
      23412: inst = 32'd203484854;
      23413: inst = 32'd471859200;
      23414: inst = 32'd136314880;
      23415: inst = 32'd268468224;
      23416: inst = 32'd201347627;
      23417: inst = 32'd203484854;
      23418: inst = 32'd471859200;
      23419: inst = 32'd136314880;
      23420: inst = 32'd268468224;
      23421: inst = 32'd201347628;
      23422: inst = 32'd203484854;
      23423: inst = 32'd471859200;
      23424: inst = 32'd136314880;
      23425: inst = 32'd268468224;
      23426: inst = 32'd201347629;
      23427: inst = 32'd203484854;
      23428: inst = 32'd471859200;
      23429: inst = 32'd136314880;
      23430: inst = 32'd268468224;
      23431: inst = 32'd201347630;
      23432: inst = 32'd203484854;
      23433: inst = 32'd471859200;
      23434: inst = 32'd136314880;
      23435: inst = 32'd268468224;
      23436: inst = 32'd201347631;
      23437: inst = 32'd203473634;
      23438: inst = 32'd471859200;
      23439: inst = 32'd136314880;
      23440: inst = 32'd268468224;
      23441: inst = 32'd201347632;
      23442: inst = 32'd203480005;
      23443: inst = 32'd471859200;
      23444: inst = 32'd136314880;
      23445: inst = 32'd268468224;
      23446: inst = 32'd201347633;
      23447: inst = 32'd203480005;
      23448: inst = 32'd471859200;
      23449: inst = 32'd136314880;
      23450: inst = 32'd268468224;
      23451: inst = 32'd201347634;
      23452: inst = 32'd203480005;
      23453: inst = 32'd471859200;
      23454: inst = 32'd136314880;
      23455: inst = 32'd268468224;
      23456: inst = 32'd201347635;
      23457: inst = 32'd203480005;
      23458: inst = 32'd471859200;
      23459: inst = 32'd136314880;
      23460: inst = 32'd268468224;
      23461: inst = 32'd201347636;
      23462: inst = 32'd203480005;
      23463: inst = 32'd471859200;
      23464: inst = 32'd136314880;
      23465: inst = 32'd268468224;
      23466: inst = 32'd201347637;
      23467: inst = 32'd203480005;
      23468: inst = 32'd471859200;
      23469: inst = 32'd136314880;
      23470: inst = 32'd268468224;
      23471: inst = 32'd201347638;
      23472: inst = 32'd203480005;
      23473: inst = 32'd471859200;
      23474: inst = 32'd136314880;
      23475: inst = 32'd268468224;
      23476: inst = 32'd201347639;
      23477: inst = 32'd203480005;
      23478: inst = 32'd471859200;
      23479: inst = 32'd136314880;
      23480: inst = 32'd268468224;
      23481: inst = 32'd201347640;
      23482: inst = 32'd203480005;
      23483: inst = 32'd471859200;
      23484: inst = 32'd136314880;
      23485: inst = 32'd268468224;
      23486: inst = 32'd201347641;
      23487: inst = 32'd203480005;
      23488: inst = 32'd471859200;
      23489: inst = 32'd136314880;
      23490: inst = 32'd268468224;
      23491: inst = 32'd201347642;
      23492: inst = 32'd203480005;
      23493: inst = 32'd471859200;
      23494: inst = 32'd136314880;
      23495: inst = 32'd268468224;
      23496: inst = 32'd201347643;
      23497: inst = 32'd203480005;
      23498: inst = 32'd471859200;
      23499: inst = 32'd136314880;
      23500: inst = 32'd268468224;
      23501: inst = 32'd201347644;
      23502: inst = 32'd203480005;
      23503: inst = 32'd471859200;
      23504: inst = 32'd136314880;
      23505: inst = 32'd268468224;
      23506: inst = 32'd201347645;
      23507: inst = 32'd203480005;
      23508: inst = 32'd471859200;
      23509: inst = 32'd136314880;
      23510: inst = 32'd268468224;
      23511: inst = 32'd201347646;
      23512: inst = 32'd203480005;
      23513: inst = 32'd471859200;
      23514: inst = 32'd136314880;
      23515: inst = 32'd268468224;
      23516: inst = 32'd201347647;
      23517: inst = 32'd203473634;
      23518: inst = 32'd471859200;
      23519: inst = 32'd136314880;
      23520: inst = 32'd268468224;
      23521: inst = 32'd201347648;
      23522: inst = 32'd203459697;
      23523: inst = 32'd471859200;
      23524: inst = 32'd136314880;
      23525: inst = 32'd268468224;
      23526: inst = 32'd201347649;
      23527: inst = 32'd203472343;
      23528: inst = 32'd471859200;
      23529: inst = 32'd136314880;
      23530: inst = 32'd268468224;
      23531: inst = 32'd201347650;
      23532: inst = 32'd203472343;
      23533: inst = 32'd471859200;
      23534: inst = 32'd136314880;
      23535: inst = 32'd268468224;
      23536: inst = 32'd201347651;
      23537: inst = 32'd203472343;
      23538: inst = 32'd471859200;
      23539: inst = 32'd136314880;
      23540: inst = 32'd268468224;
      23541: inst = 32'd201347652;
      23542: inst = 32'd203472343;
      23543: inst = 32'd471859200;
      23544: inst = 32'd136314880;
      23545: inst = 32'd268468224;
      23546: inst = 32'd201347653;
      23547: inst = 32'd203472343;
      23548: inst = 32'd471859200;
      23549: inst = 32'd136314880;
      23550: inst = 32'd268468224;
      23551: inst = 32'd201347654;
      23552: inst = 32'd203472343;
      23553: inst = 32'd471859200;
      23554: inst = 32'd136314880;
      23555: inst = 32'd268468224;
      23556: inst = 32'd201347655;
      23557: inst = 32'd203472343;
      23558: inst = 32'd471859200;
      23559: inst = 32'd136314880;
      23560: inst = 32'd268468224;
      23561: inst = 32'd201347656;
      23562: inst = 32'd203472343;
      23563: inst = 32'd471859200;
      23564: inst = 32'd136314880;
      23565: inst = 32'd268468224;
      23566: inst = 32'd201347657;
      23567: inst = 32'd203472343;
      23568: inst = 32'd471859200;
      23569: inst = 32'd136314880;
      23570: inst = 32'd268468224;
      23571: inst = 32'd201347658;
      23572: inst = 32'd203459697;
      23573: inst = 32'd471859200;
      23574: inst = 32'd136314880;
      23575: inst = 32'd268468224;
      23576: inst = 32'd201347659;
      23577: inst = 32'd203472343;
      23578: inst = 32'd471859200;
      23579: inst = 32'd136314880;
      23580: inst = 32'd268468224;
      23581: inst = 32'd201347660;
      23582: inst = 32'd203472343;
      23583: inst = 32'd471859200;
      23584: inst = 32'd136314880;
      23585: inst = 32'd268468224;
      23586: inst = 32'd201347661;
      23587: inst = 32'd203472343;
      23588: inst = 32'd471859200;
      23589: inst = 32'd136314880;
      23590: inst = 32'd268468224;
      23591: inst = 32'd201347662;
      23592: inst = 32'd203472343;
      23593: inst = 32'd471859200;
      23594: inst = 32'd136314880;
      23595: inst = 32'd268468224;
      23596: inst = 32'd201347663;
      23597: inst = 32'd203472343;
      23598: inst = 32'd471859200;
      23599: inst = 32'd136314880;
      23600: inst = 32'd268468224;
      23601: inst = 32'd201347664;
      23602: inst = 32'd203472343;
      23603: inst = 32'd471859200;
      23604: inst = 32'd136314880;
      23605: inst = 32'd268468224;
      23606: inst = 32'd201347665;
      23607: inst = 32'd203472343;
      23608: inst = 32'd471859200;
      23609: inst = 32'd136314880;
      23610: inst = 32'd268468224;
      23611: inst = 32'd201347666;
      23612: inst = 32'd203472343;
      23613: inst = 32'd471859200;
      23614: inst = 32'd136314880;
      23615: inst = 32'd268468224;
      23616: inst = 32'd201347667;
      23617: inst = 32'd203472343;
      23618: inst = 32'd471859200;
      23619: inst = 32'd136314880;
      23620: inst = 32'd268468224;
      23621: inst = 32'd201347668;
      23622: inst = 32'd203459697;
      23623: inst = 32'd471859200;
      23624: inst = 32'd136314880;
      23625: inst = 32'd268468224;
      23626: inst = 32'd201347669;
      23627: inst = 32'd203451245;
      23628: inst = 32'd471859200;
      23629: inst = 32'd136314880;
      23630: inst = 32'd268468224;
      23631: inst = 32'd201347670;
      23632: inst = 32'd203451245;
      23633: inst = 32'd471859200;
      23634: inst = 32'd136314880;
      23635: inst = 32'd268468224;
      23636: inst = 32'd201347671;
      23637: inst = 32'd203484854;
      23638: inst = 32'd471859200;
      23639: inst = 32'd136314880;
      23640: inst = 32'd268468224;
      23641: inst = 32'd201347672;
      23642: inst = 32'd203484854;
      23643: inst = 32'd471859200;
      23644: inst = 32'd136314880;
      23645: inst = 32'd268468224;
      23646: inst = 32'd201347673;
      23647: inst = 32'd203484854;
      23648: inst = 32'd471859200;
      23649: inst = 32'd136314880;
      23650: inst = 32'd268468224;
      23651: inst = 32'd201347674;
      23652: inst = 32'd203484854;
      23653: inst = 32'd471859200;
      23654: inst = 32'd136314880;
      23655: inst = 32'd268468224;
      23656: inst = 32'd201347675;
      23657: inst = 32'd203484854;
      23658: inst = 32'd471859200;
      23659: inst = 32'd136314880;
      23660: inst = 32'd268468224;
      23661: inst = 32'd201347676;
      23662: inst = 32'd203482774;
      23663: inst = 32'd471859200;
      23664: inst = 32'd136314880;
      23665: inst = 32'd268468224;
      23666: inst = 32'd201347677;
      23667: inst = 32'd203463858;
      23668: inst = 32'd471859200;
      23669: inst = 32'd136314880;
      23670: inst = 32'd268468224;
      23671: inst = 32'd201347678;
      23672: inst = 32'd203459697;
      23673: inst = 32'd471859200;
      23674: inst = 32'd136314880;
      23675: inst = 32'd268468224;
      23676: inst = 32'd201347679;
      23677: inst = 32'd203447021;
      23678: inst = 32'd471859200;
      23679: inst = 32'd136314880;
      23680: inst = 32'd268468224;
      23681: inst = 32'd201347680;
      23682: inst = 32'd203447021;
      23683: inst = 32'd471859200;
      23684: inst = 32'd136314880;
      23685: inst = 32'd268468224;
      23686: inst = 32'd201347681;
      23687: inst = 32'd203446988;
      23688: inst = 32'd471859200;
      23689: inst = 32'd136314880;
      23690: inst = 32'd268468224;
      23691: inst = 32'd201347682;
      23692: inst = 32'd203442793;
      23693: inst = 32'd471859200;
      23694: inst = 32'd136314880;
      23695: inst = 32'd268468224;
      23696: inst = 32'd201347683;
      23697: inst = 32'd203442793;
      23698: inst = 32'd471859200;
      23699: inst = 32'd136314880;
      23700: inst = 32'd268468224;
      23701: inst = 32'd201347684;
      23702: inst = 32'd203442793;
      23703: inst = 32'd471859200;
      23704: inst = 32'd136314880;
      23705: inst = 32'd268468224;
      23706: inst = 32'd201347685;
      23707: inst = 32'd203442793;
      23708: inst = 32'd471859200;
      23709: inst = 32'd136314880;
      23710: inst = 32'd268468224;
      23711: inst = 32'd201347686;
      23712: inst = 32'd203447021;
      23713: inst = 32'd471859200;
      23714: inst = 32'd136314880;
      23715: inst = 32'd268468224;
      23716: inst = 32'd201347687;
      23717: inst = 32'd203447021;
      23718: inst = 32'd471859200;
      23719: inst = 32'd136314880;
      23720: inst = 32'd268468224;
      23721: inst = 32'd201347688;
      23722: inst = 32'd203459697;
      23723: inst = 32'd471859200;
      23724: inst = 32'd136314880;
      23725: inst = 32'd268468224;
      23726: inst = 32'd201347689;
      23727: inst = 32'd203459631;
      23728: inst = 32'd471859200;
      23729: inst = 32'd136314880;
      23730: inst = 32'd268468224;
      23731: inst = 32'd201347690;
      23732: inst = 32'd203484854;
      23733: inst = 32'd471859200;
      23734: inst = 32'd136314880;
      23735: inst = 32'd268468224;
      23736: inst = 32'd201347691;
      23737: inst = 32'd203484854;
      23738: inst = 32'd471859200;
      23739: inst = 32'd136314880;
      23740: inst = 32'd268468224;
      23741: inst = 32'd201347692;
      23742: inst = 32'd203484854;
      23743: inst = 32'd471859200;
      23744: inst = 32'd136314880;
      23745: inst = 32'd268468224;
      23746: inst = 32'd201347693;
      23747: inst = 32'd203484854;
      23748: inst = 32'd471859200;
      23749: inst = 32'd136314880;
      23750: inst = 32'd268468224;
      23751: inst = 32'd201347694;
      23752: inst = 32'd203484854;
      23753: inst = 32'd471859200;
      23754: inst = 32'd136314880;
      23755: inst = 32'd268468224;
      23756: inst = 32'd201347695;
      23757: inst = 32'd203484854;
      23758: inst = 32'd471859200;
      23759: inst = 32'd136314880;
      23760: inst = 32'd268468224;
      23761: inst = 32'd201347696;
      23762: inst = 32'd203484854;
      23763: inst = 32'd471859200;
      23764: inst = 32'd136314880;
      23765: inst = 32'd268468224;
      23766: inst = 32'd201347697;
      23767: inst = 32'd203484854;
      23768: inst = 32'd471859200;
      23769: inst = 32'd136314880;
      23770: inst = 32'd268468224;
      23771: inst = 32'd201347698;
      23772: inst = 32'd203484854;
      23773: inst = 32'd471859200;
      23774: inst = 32'd136314880;
      23775: inst = 32'd268468224;
      23776: inst = 32'd201347699;
      23777: inst = 32'd203484854;
      23778: inst = 32'd471859200;
      23779: inst = 32'd136314880;
      23780: inst = 32'd268468224;
      23781: inst = 32'd201347700;
      23782: inst = 32'd203484854;
      23783: inst = 32'd471859200;
      23784: inst = 32'd136314880;
      23785: inst = 32'd268468224;
      23786: inst = 32'd201347701;
      23787: inst = 32'd203484854;
      23788: inst = 32'd471859200;
      23789: inst = 32'd136314880;
      23790: inst = 32'd268468224;
      23791: inst = 32'd201347702;
      23792: inst = 32'd203459631;
      23793: inst = 32'd471859200;
      23794: inst = 32'd136314880;
      23795: inst = 32'd268468224;
      23796: inst = 32'd201347703;
      23797: inst = 32'd203459697;
      23798: inst = 32'd471859200;
      23799: inst = 32'd136314880;
      23800: inst = 32'd268468224;
      23801: inst = 32'd201347704;
      23802: inst = 32'd203447021;
      23803: inst = 32'd471859200;
      23804: inst = 32'd136314880;
      23805: inst = 32'd268468224;
      23806: inst = 32'd201347705;
      23807: inst = 32'd203447021;
      23808: inst = 32'd471859200;
      23809: inst = 32'd136314880;
      23810: inst = 32'd268468224;
      23811: inst = 32'd201347706;
      23812: inst = 32'd203442793;
      23813: inst = 32'd471859200;
      23814: inst = 32'd136314880;
      23815: inst = 32'd268468224;
      23816: inst = 32'd201347707;
      23817: inst = 32'd203442793;
      23818: inst = 32'd471859200;
      23819: inst = 32'd136314880;
      23820: inst = 32'd268468224;
      23821: inst = 32'd201347708;
      23822: inst = 32'd203442793;
      23823: inst = 32'd471859200;
      23824: inst = 32'd136314880;
      23825: inst = 32'd268468224;
      23826: inst = 32'd201347709;
      23827: inst = 32'd203442793;
      23828: inst = 32'd471859200;
      23829: inst = 32'd136314880;
      23830: inst = 32'd268468224;
      23831: inst = 32'd201347710;
      23832: inst = 32'd203446988;
      23833: inst = 32'd471859200;
      23834: inst = 32'd136314880;
      23835: inst = 32'd268468224;
      23836: inst = 32'd201347711;
      23837: inst = 32'd203447021;
      23838: inst = 32'd471859200;
      23839: inst = 32'd136314880;
      23840: inst = 32'd268468224;
      23841: inst = 32'd201347712;
      23842: inst = 32'd203447021;
      23843: inst = 32'd471859200;
      23844: inst = 32'd136314880;
      23845: inst = 32'd268468224;
      23846: inst = 32'd201347713;
      23847: inst = 32'd203459697;
      23848: inst = 32'd471859200;
      23849: inst = 32'd136314880;
      23850: inst = 32'd268468224;
      23851: inst = 32'd201347714;
      23852: inst = 32'd203463858;
      23853: inst = 32'd471859200;
      23854: inst = 32'd136314880;
      23855: inst = 32'd268468224;
      23856: inst = 32'd201347715;
      23857: inst = 32'd203482774;
      23858: inst = 32'd471859200;
      23859: inst = 32'd136314880;
      23860: inst = 32'd268468224;
      23861: inst = 32'd201347716;
      23862: inst = 32'd203484854;
      23863: inst = 32'd471859200;
      23864: inst = 32'd136314880;
      23865: inst = 32'd268468224;
      23866: inst = 32'd201347717;
      23867: inst = 32'd203484854;
      23868: inst = 32'd471859200;
      23869: inst = 32'd136314880;
      23870: inst = 32'd268468224;
      23871: inst = 32'd201347718;
      23872: inst = 32'd203484854;
      23873: inst = 32'd471859200;
      23874: inst = 32'd136314880;
      23875: inst = 32'd268468224;
      23876: inst = 32'd201347719;
      23877: inst = 32'd203484854;
      23878: inst = 32'd471859200;
      23879: inst = 32'd136314880;
      23880: inst = 32'd268468224;
      23881: inst = 32'd201347720;
      23882: inst = 32'd203484854;
      23883: inst = 32'd471859200;
      23884: inst = 32'd136314880;
      23885: inst = 32'd268468224;
      23886: inst = 32'd201347721;
      23887: inst = 32'd203484854;
      23888: inst = 32'd471859200;
      23889: inst = 32'd136314880;
      23890: inst = 32'd268468224;
      23891: inst = 32'd201347722;
      23892: inst = 32'd203484854;
      23893: inst = 32'd471859200;
      23894: inst = 32'd136314880;
      23895: inst = 32'd268468224;
      23896: inst = 32'd201347723;
      23897: inst = 32'd203484854;
      23898: inst = 32'd471859200;
      23899: inst = 32'd136314880;
      23900: inst = 32'd268468224;
      23901: inst = 32'd201347724;
      23902: inst = 32'd203484854;
      23903: inst = 32'd471859200;
      23904: inst = 32'd136314880;
      23905: inst = 32'd268468224;
      23906: inst = 32'd201347725;
      23907: inst = 32'd203484854;
      23908: inst = 32'd471859200;
      23909: inst = 32'd136314880;
      23910: inst = 32'd268468224;
      23911: inst = 32'd201347726;
      23912: inst = 32'd203484854;
      23913: inst = 32'd471859200;
      23914: inst = 32'd136314880;
      23915: inst = 32'd268468224;
      23916: inst = 32'd201347727;
      23917: inst = 32'd203473634;
      23918: inst = 32'd471859200;
      23919: inst = 32'd136314880;
      23920: inst = 32'd268468224;
      23921: inst = 32'd201347728;
      23922: inst = 32'd203480005;
      23923: inst = 32'd471859200;
      23924: inst = 32'd136314880;
      23925: inst = 32'd268468224;
      23926: inst = 32'd201347729;
      23927: inst = 32'd203480005;
      23928: inst = 32'd471859200;
      23929: inst = 32'd136314880;
      23930: inst = 32'd268468224;
      23931: inst = 32'd201347730;
      23932: inst = 32'd203480005;
      23933: inst = 32'd471859200;
      23934: inst = 32'd136314880;
      23935: inst = 32'd268468224;
      23936: inst = 32'd201347731;
      23937: inst = 32'd203480005;
      23938: inst = 32'd471859200;
      23939: inst = 32'd136314880;
      23940: inst = 32'd268468224;
      23941: inst = 32'd201347732;
      23942: inst = 32'd203480005;
      23943: inst = 32'd471859200;
      23944: inst = 32'd136314880;
      23945: inst = 32'd268468224;
      23946: inst = 32'd201347733;
      23947: inst = 32'd203480005;
      23948: inst = 32'd471859200;
      23949: inst = 32'd136314880;
      23950: inst = 32'd268468224;
      23951: inst = 32'd201347734;
      23952: inst = 32'd203480005;
      23953: inst = 32'd471859200;
      23954: inst = 32'd136314880;
      23955: inst = 32'd268468224;
      23956: inst = 32'd201347735;
      23957: inst = 32'd203480005;
      23958: inst = 32'd471859200;
      23959: inst = 32'd136314880;
      23960: inst = 32'd268468224;
      23961: inst = 32'd201347736;
      23962: inst = 32'd203480005;
      23963: inst = 32'd471859200;
      23964: inst = 32'd136314880;
      23965: inst = 32'd268468224;
      23966: inst = 32'd201347737;
      23967: inst = 32'd203480005;
      23968: inst = 32'd471859200;
      23969: inst = 32'd136314880;
      23970: inst = 32'd268468224;
      23971: inst = 32'd201347738;
      23972: inst = 32'd203480005;
      23973: inst = 32'd471859200;
      23974: inst = 32'd136314880;
      23975: inst = 32'd268468224;
      23976: inst = 32'd201347739;
      23977: inst = 32'd203480005;
      23978: inst = 32'd471859200;
      23979: inst = 32'd136314880;
      23980: inst = 32'd268468224;
      23981: inst = 32'd201347740;
      23982: inst = 32'd203480005;
      23983: inst = 32'd471859200;
      23984: inst = 32'd136314880;
      23985: inst = 32'd268468224;
      23986: inst = 32'd201347741;
      23987: inst = 32'd203480005;
      23988: inst = 32'd471859200;
      23989: inst = 32'd136314880;
      23990: inst = 32'd268468224;
      23991: inst = 32'd201347742;
      23992: inst = 32'd203480005;
      23993: inst = 32'd471859200;
      23994: inst = 32'd136314880;
      23995: inst = 32'd268468224;
      23996: inst = 32'd201347743;
      23997: inst = 32'd203473634;
      23998: inst = 32'd471859200;
      23999: inst = 32'd136314880;
      24000: inst = 32'd268468224;
      24001: inst = 32'd201347744;
      24002: inst = 32'd203459697;
      24003: inst = 32'd471859200;
      24004: inst = 32'd136314880;
      24005: inst = 32'd268468224;
      24006: inst = 32'd201347745;
      24007: inst = 32'd203459697;
      24008: inst = 32'd471859200;
      24009: inst = 32'd136314880;
      24010: inst = 32'd268468224;
      24011: inst = 32'd201347746;
      24012: inst = 32'd203459697;
      24013: inst = 32'd471859200;
      24014: inst = 32'd136314880;
      24015: inst = 32'd268468224;
      24016: inst = 32'd201347747;
      24017: inst = 32'd203459697;
      24018: inst = 32'd471859200;
      24019: inst = 32'd136314880;
      24020: inst = 32'd268468224;
      24021: inst = 32'd201347748;
      24022: inst = 32'd203459697;
      24023: inst = 32'd471859200;
      24024: inst = 32'd136314880;
      24025: inst = 32'd268468224;
      24026: inst = 32'd201347749;
      24027: inst = 32'd203459697;
      24028: inst = 32'd471859200;
      24029: inst = 32'd136314880;
      24030: inst = 32'd268468224;
      24031: inst = 32'd201347750;
      24032: inst = 32'd203459697;
      24033: inst = 32'd471859200;
      24034: inst = 32'd136314880;
      24035: inst = 32'd268468224;
      24036: inst = 32'd201347751;
      24037: inst = 32'd203459697;
      24038: inst = 32'd471859200;
      24039: inst = 32'd136314880;
      24040: inst = 32'd268468224;
      24041: inst = 32'd201347752;
      24042: inst = 32'd203459697;
      24043: inst = 32'd471859200;
      24044: inst = 32'd136314880;
      24045: inst = 32'd268468224;
      24046: inst = 32'd201347753;
      24047: inst = 32'd203459697;
      24048: inst = 32'd471859200;
      24049: inst = 32'd136314880;
      24050: inst = 32'd268468224;
      24051: inst = 32'd201347754;
      24052: inst = 32'd203459697;
      24053: inst = 32'd471859200;
      24054: inst = 32'd136314880;
      24055: inst = 32'd268468224;
      24056: inst = 32'd201347755;
      24057: inst = 32'd203459697;
      24058: inst = 32'd471859200;
      24059: inst = 32'd136314880;
      24060: inst = 32'd268468224;
      24061: inst = 32'd201347756;
      24062: inst = 32'd203459697;
      24063: inst = 32'd471859200;
      24064: inst = 32'd136314880;
      24065: inst = 32'd268468224;
      24066: inst = 32'd201347757;
      24067: inst = 32'd203459697;
      24068: inst = 32'd471859200;
      24069: inst = 32'd136314880;
      24070: inst = 32'd268468224;
      24071: inst = 32'd201347758;
      24072: inst = 32'd203459697;
      24073: inst = 32'd471859200;
      24074: inst = 32'd136314880;
      24075: inst = 32'd268468224;
      24076: inst = 32'd201347759;
      24077: inst = 32'd203459697;
      24078: inst = 32'd471859200;
      24079: inst = 32'd136314880;
      24080: inst = 32'd268468224;
      24081: inst = 32'd201347760;
      24082: inst = 32'd203459697;
      24083: inst = 32'd471859200;
      24084: inst = 32'd136314880;
      24085: inst = 32'd268468224;
      24086: inst = 32'd201347761;
      24087: inst = 32'd203459697;
      24088: inst = 32'd471859200;
      24089: inst = 32'd136314880;
      24090: inst = 32'd268468224;
      24091: inst = 32'd201347762;
      24092: inst = 32'd203459697;
      24093: inst = 32'd471859200;
      24094: inst = 32'd136314880;
      24095: inst = 32'd268468224;
      24096: inst = 32'd201347763;
      24097: inst = 32'd203459697;
      24098: inst = 32'd471859200;
      24099: inst = 32'd136314880;
      24100: inst = 32'd268468224;
      24101: inst = 32'd201347764;
      24102: inst = 32'd203459697;
      24103: inst = 32'd471859200;
      24104: inst = 32'd136314880;
      24105: inst = 32'd268468224;
      24106: inst = 32'd201347765;
      24107: inst = 32'd203451245;
      24108: inst = 32'd471859200;
      24109: inst = 32'd136314880;
      24110: inst = 32'd268468224;
      24111: inst = 32'd201347766;
      24112: inst = 32'd203451245;
      24113: inst = 32'd471859200;
      24114: inst = 32'd136314880;
      24115: inst = 32'd268468224;
      24116: inst = 32'd201347767;
      24117: inst = 32'd203484854;
      24118: inst = 32'd471859200;
      24119: inst = 32'd136314880;
      24120: inst = 32'd268468224;
      24121: inst = 32'd201347768;
      24122: inst = 32'd203484854;
      24123: inst = 32'd471859200;
      24124: inst = 32'd136314880;
      24125: inst = 32'd268468224;
      24126: inst = 32'd201347769;
      24127: inst = 32'd203484854;
      24128: inst = 32'd471859200;
      24129: inst = 32'd136314880;
      24130: inst = 32'd268468224;
      24131: inst = 32'd201347770;
      24132: inst = 32'd203484854;
      24133: inst = 32'd471859200;
      24134: inst = 32'd136314880;
      24135: inst = 32'd268468224;
      24136: inst = 32'd201347771;
      24137: inst = 32'd203484854;
      24138: inst = 32'd471859200;
      24139: inst = 32'd136314880;
      24140: inst = 32'd268468224;
      24141: inst = 32'd201347772;
      24142: inst = 32'd203468083;
      24143: inst = 32'd471859200;
      24144: inst = 32'd136314880;
      24145: inst = 32'd268468224;
      24146: inst = 32'd201347773;
      24147: inst = 32'd203459697;
      24148: inst = 32'd471859200;
      24149: inst = 32'd136314880;
      24150: inst = 32'd268468224;
      24151: inst = 32'd201347774;
      24152: inst = 32'd203459697;
      24153: inst = 32'd471859200;
      24154: inst = 32'd136314880;
      24155: inst = 32'd268468224;
      24156: inst = 32'd201347775;
      24157: inst = 32'd203447021;
      24158: inst = 32'd471859200;
      24159: inst = 32'd136314880;
      24160: inst = 32'd268468224;
      24161: inst = 32'd201347776;
      24162: inst = 32'd203447021;
      24163: inst = 32'd471859200;
      24164: inst = 32'd136314880;
      24165: inst = 32'd268468224;
      24166: inst = 32'd201347777;
      24167: inst = 32'd203446988;
      24168: inst = 32'd471859200;
      24169: inst = 32'd136314880;
      24170: inst = 32'd268468224;
      24171: inst = 32'd201347778;
      24172: inst = 32'd203442793;
      24173: inst = 32'd471859200;
      24174: inst = 32'd136314880;
      24175: inst = 32'd268468224;
      24176: inst = 32'd201347779;
      24177: inst = 32'd203442793;
      24178: inst = 32'd471859200;
      24179: inst = 32'd136314880;
      24180: inst = 32'd268468224;
      24181: inst = 32'd201347780;
      24182: inst = 32'd203442793;
      24183: inst = 32'd471859200;
      24184: inst = 32'd136314880;
      24185: inst = 32'd268468224;
      24186: inst = 32'd201347781;
      24187: inst = 32'd203444874;
      24188: inst = 32'd471859200;
      24189: inst = 32'd136314880;
      24190: inst = 32'd268468224;
      24191: inst = 32'd201347782;
      24192: inst = 32'd203447021;
      24193: inst = 32'd471859200;
      24194: inst = 32'd136314880;
      24195: inst = 32'd268468224;
      24196: inst = 32'd201347783;
      24197: inst = 32'd203447021;
      24198: inst = 32'd471859200;
      24199: inst = 32'd136314880;
      24200: inst = 32'd268468224;
      24201: inst = 32'd201347784;
      24202: inst = 32'd203459697;
      24203: inst = 32'd471859200;
      24204: inst = 32'd136314880;
      24205: inst = 32'd268468224;
      24206: inst = 32'd201347785;
      24207: inst = 32'd203457518;
      24208: inst = 32'd471859200;
      24209: inst = 32'd136314880;
      24210: inst = 32'd268468224;
      24211: inst = 32'd201347786;
      24212: inst = 32'd203484854;
      24213: inst = 32'd471859200;
      24214: inst = 32'd136314880;
      24215: inst = 32'd268468224;
      24216: inst = 32'd201347787;
      24217: inst = 32'd203484854;
      24218: inst = 32'd471859200;
      24219: inst = 32'd136314880;
      24220: inst = 32'd268468224;
      24221: inst = 32'd201347788;
      24222: inst = 32'd203484854;
      24223: inst = 32'd471859200;
      24224: inst = 32'd136314880;
      24225: inst = 32'd268468224;
      24226: inst = 32'd201347789;
      24227: inst = 32'd203484854;
      24228: inst = 32'd471859200;
      24229: inst = 32'd136314880;
      24230: inst = 32'd268468224;
      24231: inst = 32'd201347790;
      24232: inst = 32'd203484854;
      24233: inst = 32'd471859200;
      24234: inst = 32'd136314880;
      24235: inst = 32'd268468224;
      24236: inst = 32'd201347791;
      24237: inst = 32'd203484854;
      24238: inst = 32'd471859200;
      24239: inst = 32'd136314880;
      24240: inst = 32'd268468224;
      24241: inst = 32'd201347792;
      24242: inst = 32'd203484854;
      24243: inst = 32'd471859200;
      24244: inst = 32'd136314880;
      24245: inst = 32'd268468224;
      24246: inst = 32'd201347793;
      24247: inst = 32'd203484854;
      24248: inst = 32'd471859200;
      24249: inst = 32'd136314880;
      24250: inst = 32'd268468224;
      24251: inst = 32'd201347794;
      24252: inst = 32'd203484854;
      24253: inst = 32'd471859200;
      24254: inst = 32'd136314880;
      24255: inst = 32'd268468224;
      24256: inst = 32'd201347795;
      24257: inst = 32'd203484854;
      24258: inst = 32'd471859200;
      24259: inst = 32'd136314880;
      24260: inst = 32'd268468224;
      24261: inst = 32'd201347796;
      24262: inst = 32'd203484854;
      24263: inst = 32'd471859200;
      24264: inst = 32'd136314880;
      24265: inst = 32'd268468224;
      24266: inst = 32'd201347797;
      24267: inst = 32'd203484854;
      24268: inst = 32'd471859200;
      24269: inst = 32'd136314880;
      24270: inst = 32'd268468224;
      24271: inst = 32'd201347798;
      24272: inst = 32'd203457518;
      24273: inst = 32'd471859200;
      24274: inst = 32'd136314880;
      24275: inst = 32'd268468224;
      24276: inst = 32'd201347799;
      24277: inst = 32'd203459697;
      24278: inst = 32'd471859200;
      24279: inst = 32'd136314880;
      24280: inst = 32'd268468224;
      24281: inst = 32'd201347800;
      24282: inst = 32'd203447021;
      24283: inst = 32'd471859200;
      24284: inst = 32'd136314880;
      24285: inst = 32'd268468224;
      24286: inst = 32'd201347801;
      24287: inst = 32'd203447021;
      24288: inst = 32'd471859200;
      24289: inst = 32'd136314880;
      24290: inst = 32'd268468224;
      24291: inst = 32'd201347802;
      24292: inst = 32'd203444874;
      24293: inst = 32'd471859200;
      24294: inst = 32'd136314880;
      24295: inst = 32'd268468224;
      24296: inst = 32'd201347803;
      24297: inst = 32'd203442793;
      24298: inst = 32'd471859200;
      24299: inst = 32'd136314880;
      24300: inst = 32'd268468224;
      24301: inst = 32'd201347804;
      24302: inst = 32'd203442793;
      24303: inst = 32'd471859200;
      24304: inst = 32'd136314880;
      24305: inst = 32'd268468224;
      24306: inst = 32'd201347805;
      24307: inst = 32'd203442793;
      24308: inst = 32'd471859200;
      24309: inst = 32'd136314880;
      24310: inst = 32'd268468224;
      24311: inst = 32'd201347806;
      24312: inst = 32'd203446988;
      24313: inst = 32'd471859200;
      24314: inst = 32'd136314880;
      24315: inst = 32'd268468224;
      24316: inst = 32'd201347807;
      24317: inst = 32'd203447021;
      24318: inst = 32'd471859200;
      24319: inst = 32'd136314880;
      24320: inst = 32'd268468224;
      24321: inst = 32'd201347808;
      24322: inst = 32'd203447021;
      24323: inst = 32'd471859200;
      24324: inst = 32'd136314880;
      24325: inst = 32'd268468224;
      24326: inst = 32'd201347809;
      24327: inst = 32'd203459697;
      24328: inst = 32'd471859200;
      24329: inst = 32'd136314880;
      24330: inst = 32'd268468224;
      24331: inst = 32'd201347810;
      24332: inst = 32'd203459697;
      24333: inst = 32'd471859200;
      24334: inst = 32'd136314880;
      24335: inst = 32'd268468224;
      24336: inst = 32'd201347811;
      24337: inst = 32'd203468083;
      24338: inst = 32'd471859200;
      24339: inst = 32'd136314880;
      24340: inst = 32'd268468224;
      24341: inst = 32'd201347812;
      24342: inst = 32'd203484854;
      24343: inst = 32'd471859200;
      24344: inst = 32'd136314880;
      24345: inst = 32'd268468224;
      24346: inst = 32'd201347813;
      24347: inst = 32'd203484854;
      24348: inst = 32'd471859200;
      24349: inst = 32'd136314880;
      24350: inst = 32'd268468224;
      24351: inst = 32'd201347814;
      24352: inst = 32'd203484854;
      24353: inst = 32'd471859200;
      24354: inst = 32'd136314880;
      24355: inst = 32'd268468224;
      24356: inst = 32'd201347815;
      24357: inst = 32'd203484854;
      24358: inst = 32'd471859200;
      24359: inst = 32'd136314880;
      24360: inst = 32'd268468224;
      24361: inst = 32'd201347816;
      24362: inst = 32'd203484854;
      24363: inst = 32'd471859200;
      24364: inst = 32'd136314880;
      24365: inst = 32'd268468224;
      24366: inst = 32'd201347817;
      24367: inst = 32'd203484854;
      24368: inst = 32'd471859200;
      24369: inst = 32'd136314880;
      24370: inst = 32'd268468224;
      24371: inst = 32'd201347818;
      24372: inst = 32'd203484854;
      24373: inst = 32'd471859200;
      24374: inst = 32'd136314880;
      24375: inst = 32'd268468224;
      24376: inst = 32'd201347819;
      24377: inst = 32'd203484854;
      24378: inst = 32'd471859200;
      24379: inst = 32'd136314880;
      24380: inst = 32'd268468224;
      24381: inst = 32'd201347820;
      24382: inst = 32'd203484854;
      24383: inst = 32'd471859200;
      24384: inst = 32'd136314880;
      24385: inst = 32'd268468224;
      24386: inst = 32'd201347821;
      24387: inst = 32'd203484854;
      24388: inst = 32'd471859200;
      24389: inst = 32'd136314880;
      24390: inst = 32'd268468224;
      24391: inst = 32'd201347822;
      24392: inst = 32'd203484854;
      24393: inst = 32'd471859200;
      24394: inst = 32'd136314880;
      24395: inst = 32'd268468224;
      24396: inst = 32'd201347823;
      24397: inst = 32'd203473634;
      24398: inst = 32'd471859200;
      24399: inst = 32'd136314880;
      24400: inst = 32'd268468224;
      24401: inst = 32'd201347824;
      24402: inst = 32'd203473634;
      24403: inst = 32'd471859200;
      24404: inst = 32'd136314880;
      24405: inst = 32'd268468224;
      24406: inst = 32'd201347825;
      24407: inst = 32'd203473634;
      24408: inst = 32'd471859200;
      24409: inst = 32'd136314880;
      24410: inst = 32'd268468224;
      24411: inst = 32'd201347826;
      24412: inst = 32'd203473634;
      24413: inst = 32'd471859200;
      24414: inst = 32'd136314880;
      24415: inst = 32'd268468224;
      24416: inst = 32'd201347827;
      24417: inst = 32'd203473634;
      24418: inst = 32'd471859200;
      24419: inst = 32'd136314880;
      24420: inst = 32'd268468224;
      24421: inst = 32'd201347828;
      24422: inst = 32'd203473634;
      24423: inst = 32'd471859200;
      24424: inst = 32'd136314880;
      24425: inst = 32'd268468224;
      24426: inst = 32'd201347829;
      24427: inst = 32'd203473634;
      24428: inst = 32'd471859200;
      24429: inst = 32'd136314880;
      24430: inst = 32'd268468224;
      24431: inst = 32'd201347830;
      24432: inst = 32'd203473634;
      24433: inst = 32'd471859200;
      24434: inst = 32'd136314880;
      24435: inst = 32'd268468224;
      24436: inst = 32'd201347831;
      24437: inst = 32'd203473634;
      24438: inst = 32'd471859200;
      24439: inst = 32'd136314880;
      24440: inst = 32'd268468224;
      24441: inst = 32'd201347832;
      24442: inst = 32'd203473634;
      24443: inst = 32'd471859200;
      24444: inst = 32'd136314880;
      24445: inst = 32'd268468224;
      24446: inst = 32'd201347833;
      24447: inst = 32'd203473634;
      24448: inst = 32'd471859200;
      24449: inst = 32'd136314880;
      24450: inst = 32'd268468224;
      24451: inst = 32'd201347834;
      24452: inst = 32'd203473634;
      24453: inst = 32'd471859200;
      24454: inst = 32'd136314880;
      24455: inst = 32'd268468224;
      24456: inst = 32'd201347835;
      24457: inst = 32'd203473634;
      24458: inst = 32'd471859200;
      24459: inst = 32'd136314880;
      24460: inst = 32'd268468224;
      24461: inst = 32'd201347836;
      24462: inst = 32'd203473634;
      24463: inst = 32'd471859200;
      24464: inst = 32'd136314880;
      24465: inst = 32'd268468224;
      24466: inst = 32'd201347837;
      24467: inst = 32'd203473634;
      24468: inst = 32'd471859200;
      24469: inst = 32'd136314880;
      24470: inst = 32'd268468224;
      24471: inst = 32'd201347838;
      24472: inst = 32'd203473634;
      24473: inst = 32'd471859200;
      24474: inst = 32'd136314880;
      24475: inst = 32'd268468224;
      24476: inst = 32'd201347839;
      24477: inst = 32'd203473634;
      24478: inst = 32'd471859200;
      24479: inst = 32'd136314880;
      24480: inst = 32'd268468224;
      24481: inst = 32'd201347840;
      24482: inst = 32'd203451216;
      24483: inst = 32'd471859200;
      24484: inst = 32'd136314880;
      24485: inst = 32'd268468224;
      24486: inst = 32'd201347841;
      24487: inst = 32'd203451216;
      24488: inst = 32'd471859200;
      24489: inst = 32'd136314880;
      24490: inst = 32'd268468224;
      24491: inst = 32'd201347842;
      24492: inst = 32'd203451216;
      24493: inst = 32'd471859200;
      24494: inst = 32'd136314880;
      24495: inst = 32'd268468224;
      24496: inst = 32'd201347843;
      24497: inst = 32'd203451216;
      24498: inst = 32'd471859200;
      24499: inst = 32'd136314880;
      24500: inst = 32'd268468224;
      24501: inst = 32'd201347844;
      24502: inst = 32'd203451216;
      24503: inst = 32'd471859200;
      24504: inst = 32'd136314880;
      24505: inst = 32'd268468224;
      24506: inst = 32'd201347845;
      24507: inst = 32'd203451216;
      24508: inst = 32'd471859200;
      24509: inst = 32'd136314880;
      24510: inst = 32'd268468224;
      24511: inst = 32'd201347846;
      24512: inst = 32'd203451216;
      24513: inst = 32'd471859200;
      24514: inst = 32'd136314880;
      24515: inst = 32'd268468224;
      24516: inst = 32'd201347847;
      24517: inst = 32'd203451216;
      24518: inst = 32'd471859200;
      24519: inst = 32'd136314880;
      24520: inst = 32'd268468224;
      24521: inst = 32'd201347848;
      24522: inst = 32'd203451216;
      24523: inst = 32'd471859200;
      24524: inst = 32'd136314880;
      24525: inst = 32'd268468224;
      24526: inst = 32'd201347849;
      24527: inst = 32'd203451216;
      24528: inst = 32'd471859200;
      24529: inst = 32'd136314880;
      24530: inst = 32'd268468224;
      24531: inst = 32'd201347850;
      24532: inst = 32'd203451216;
      24533: inst = 32'd471859200;
      24534: inst = 32'd136314880;
      24535: inst = 32'd268468224;
      24536: inst = 32'd201347851;
      24537: inst = 32'd203451216;
      24538: inst = 32'd471859200;
      24539: inst = 32'd136314880;
      24540: inst = 32'd268468224;
      24541: inst = 32'd201347852;
      24542: inst = 32'd203451216;
      24543: inst = 32'd471859200;
      24544: inst = 32'd136314880;
      24545: inst = 32'd268468224;
      24546: inst = 32'd201347853;
      24547: inst = 32'd203451216;
      24548: inst = 32'd471859200;
      24549: inst = 32'd136314880;
      24550: inst = 32'd268468224;
      24551: inst = 32'd201347854;
      24552: inst = 32'd203451216;
      24553: inst = 32'd471859200;
      24554: inst = 32'd136314880;
      24555: inst = 32'd268468224;
      24556: inst = 32'd201347855;
      24557: inst = 32'd203451216;
      24558: inst = 32'd471859200;
      24559: inst = 32'd136314880;
      24560: inst = 32'd268468224;
      24561: inst = 32'd201347856;
      24562: inst = 32'd203451216;
      24563: inst = 32'd471859200;
      24564: inst = 32'd136314880;
      24565: inst = 32'd268468224;
      24566: inst = 32'd201347857;
      24567: inst = 32'd203451216;
      24568: inst = 32'd471859200;
      24569: inst = 32'd136314880;
      24570: inst = 32'd268468224;
      24571: inst = 32'd201347858;
      24572: inst = 32'd203451216;
      24573: inst = 32'd471859200;
      24574: inst = 32'd136314880;
      24575: inst = 32'd268468224;
      24576: inst = 32'd201347859;
      24577: inst = 32'd203451216;
      24578: inst = 32'd471859200;
      24579: inst = 32'd136314880;
      24580: inst = 32'd268468224;
      24581: inst = 32'd201347860;
      24582: inst = 32'd203451216;
      24583: inst = 32'd471859200;
      24584: inst = 32'd136314880;
      24585: inst = 32'd268468224;
      24586: inst = 32'd201347861;
      24587: inst = 32'd203451216;
      24588: inst = 32'd471859200;
      24589: inst = 32'd136314880;
      24590: inst = 32'd268468224;
      24591: inst = 32'd201347862;
      24592: inst = 32'd203451216;
      24593: inst = 32'd471859200;
      24594: inst = 32'd136314880;
      24595: inst = 32'd268468224;
      24596: inst = 32'd201347863;
      24597: inst = 32'd203451216;
      24598: inst = 32'd471859200;
      24599: inst = 32'd136314880;
      24600: inst = 32'd268468224;
      24601: inst = 32'd201347864;
      24602: inst = 32'd203451216;
      24603: inst = 32'd471859200;
      24604: inst = 32'd136314880;
      24605: inst = 32'd268468224;
      24606: inst = 32'd201347865;
      24607: inst = 32'd203451216;
      24608: inst = 32'd471859200;
      24609: inst = 32'd136314880;
      24610: inst = 32'd268468224;
      24611: inst = 32'd201347866;
      24612: inst = 32'd203451216;
      24613: inst = 32'd471859200;
      24614: inst = 32'd136314880;
      24615: inst = 32'd268468224;
      24616: inst = 32'd201347867;
      24617: inst = 32'd203455440;
      24618: inst = 32'd471859200;
      24619: inst = 32'd136314880;
      24620: inst = 32'd268468224;
      24621: inst = 32'd201347868;
      24622: inst = 32'd203459697;
      24623: inst = 32'd471859200;
      24624: inst = 32'd136314880;
      24625: inst = 32'd268468224;
      24626: inst = 32'd201347869;
      24627: inst = 32'd203459697;
      24628: inst = 32'd471859200;
      24629: inst = 32'd136314880;
      24630: inst = 32'd268468224;
      24631: inst = 32'd201347870;
      24632: inst = 32'd203459697;
      24633: inst = 32'd471859200;
      24634: inst = 32'd136314880;
      24635: inst = 32'd268468224;
      24636: inst = 32'd201347871;
      24637: inst = 32'd203459697;
      24638: inst = 32'd471859200;
      24639: inst = 32'd136314880;
      24640: inst = 32'd268468224;
      24641: inst = 32'd201347872;
      24642: inst = 32'd203459697;
      24643: inst = 32'd471859200;
      24644: inst = 32'd136314880;
      24645: inst = 32'd268468224;
      24646: inst = 32'd201347873;
      24647: inst = 32'd203455439;
      24648: inst = 32'd471859200;
      24649: inst = 32'd136314880;
      24650: inst = 32'd268468224;
      24651: inst = 32'd201347874;
      24652: inst = 32'd203442793;
      24653: inst = 32'd471859200;
      24654: inst = 32'd136314880;
      24655: inst = 32'd268468224;
      24656: inst = 32'd201347875;
      24657: inst = 32'd203442793;
      24658: inst = 32'd471859200;
      24659: inst = 32'd136314880;
      24660: inst = 32'd268468224;
      24661: inst = 32'd201347876;
      24662: inst = 32'd203442793;
      24663: inst = 32'd471859200;
      24664: inst = 32'd136314880;
      24665: inst = 32'd268468224;
      24666: inst = 32'd201347877;
      24667: inst = 32'd203451245;
      24668: inst = 32'd471859200;
      24669: inst = 32'd136314880;
      24670: inst = 32'd268468224;
      24671: inst = 32'd201347878;
      24672: inst = 32'd203459697;
      24673: inst = 32'd471859200;
      24674: inst = 32'd136314880;
      24675: inst = 32'd268468224;
      24676: inst = 32'd201347879;
      24677: inst = 32'd203459697;
      24678: inst = 32'd471859200;
      24679: inst = 32'd136314880;
      24680: inst = 32'd268468224;
      24681: inst = 32'd201347880;
      24682: inst = 32'd203459697;
      24683: inst = 32'd471859200;
      24684: inst = 32'd136314880;
      24685: inst = 32'd268468224;
      24686: inst = 32'd201347881;
      24687: inst = 32'd203447020;
      24688: inst = 32'd471859200;
      24689: inst = 32'd136314880;
      24690: inst = 32'd268468224;
      24691: inst = 32'd201347882;
      24692: inst = 32'd203451216;
      24693: inst = 32'd471859200;
      24694: inst = 32'd136314880;
      24695: inst = 32'd268468224;
      24696: inst = 32'd201347883;
      24697: inst = 32'd203451216;
      24698: inst = 32'd471859200;
      24699: inst = 32'd136314880;
      24700: inst = 32'd268468224;
      24701: inst = 32'd201347884;
      24702: inst = 32'd203451216;
      24703: inst = 32'd471859200;
      24704: inst = 32'd136314880;
      24705: inst = 32'd268468224;
      24706: inst = 32'd201347885;
      24707: inst = 32'd203451216;
      24708: inst = 32'd471859200;
      24709: inst = 32'd136314880;
      24710: inst = 32'd268468224;
      24711: inst = 32'd201347886;
      24712: inst = 32'd203451216;
      24713: inst = 32'd471859200;
      24714: inst = 32'd136314880;
      24715: inst = 32'd268468224;
      24716: inst = 32'd201347887;
      24717: inst = 32'd203451216;
      24718: inst = 32'd471859200;
      24719: inst = 32'd136314880;
      24720: inst = 32'd268468224;
      24721: inst = 32'd201347888;
      24722: inst = 32'd203451216;
      24723: inst = 32'd471859200;
      24724: inst = 32'd136314880;
      24725: inst = 32'd268468224;
      24726: inst = 32'd201347889;
      24727: inst = 32'd203451216;
      24728: inst = 32'd471859200;
      24729: inst = 32'd136314880;
      24730: inst = 32'd268468224;
      24731: inst = 32'd201347890;
      24732: inst = 32'd203451216;
      24733: inst = 32'd471859200;
      24734: inst = 32'd136314880;
      24735: inst = 32'd268468224;
      24736: inst = 32'd201347891;
      24737: inst = 32'd203451216;
      24738: inst = 32'd471859200;
      24739: inst = 32'd136314880;
      24740: inst = 32'd268468224;
      24741: inst = 32'd201347892;
      24742: inst = 32'd203451216;
      24743: inst = 32'd471859200;
      24744: inst = 32'd136314880;
      24745: inst = 32'd268468224;
      24746: inst = 32'd201347893;
      24747: inst = 32'd203451216;
      24748: inst = 32'd471859200;
      24749: inst = 32'd136314880;
      24750: inst = 32'd268468224;
      24751: inst = 32'd201347894;
      24752: inst = 32'd203446987;
      24753: inst = 32'd471859200;
      24754: inst = 32'd136314880;
      24755: inst = 32'd268468224;
      24756: inst = 32'd201347895;
      24757: inst = 32'd203459697;
      24758: inst = 32'd471859200;
      24759: inst = 32'd136314880;
      24760: inst = 32'd268468224;
      24761: inst = 32'd201347896;
      24762: inst = 32'd203459697;
      24763: inst = 32'd471859200;
      24764: inst = 32'd136314880;
      24765: inst = 32'd268468224;
      24766: inst = 32'd201347897;
      24767: inst = 32'd203459697;
      24768: inst = 32'd471859200;
      24769: inst = 32'd136314880;
      24770: inst = 32'd268468224;
      24771: inst = 32'd201347898;
      24772: inst = 32'd203451245;
      24773: inst = 32'd471859200;
      24774: inst = 32'd136314880;
      24775: inst = 32'd268468224;
      24776: inst = 32'd201347899;
      24777: inst = 32'd203442793;
      24778: inst = 32'd471859200;
      24779: inst = 32'd136314880;
      24780: inst = 32'd268468224;
      24781: inst = 32'd201347900;
      24782: inst = 32'd203442793;
      24783: inst = 32'd471859200;
      24784: inst = 32'd136314880;
      24785: inst = 32'd268468224;
      24786: inst = 32'd201347901;
      24787: inst = 32'd203442793;
      24788: inst = 32'd471859200;
      24789: inst = 32'd136314880;
      24790: inst = 32'd268468224;
      24791: inst = 32'd201347902;
      24792: inst = 32'd203455439;
      24793: inst = 32'd471859200;
      24794: inst = 32'd136314880;
      24795: inst = 32'd268468224;
      24796: inst = 32'd201347903;
      24797: inst = 32'd203459697;
      24798: inst = 32'd471859200;
      24799: inst = 32'd136314880;
      24800: inst = 32'd268468224;
      24801: inst = 32'd201347904;
      24802: inst = 32'd203459697;
      24803: inst = 32'd471859200;
      24804: inst = 32'd136314880;
      24805: inst = 32'd268468224;
      24806: inst = 32'd201347905;
      24807: inst = 32'd203459697;
      24808: inst = 32'd471859200;
      24809: inst = 32'd136314880;
      24810: inst = 32'd268468224;
      24811: inst = 32'd201347906;
      24812: inst = 32'd203459697;
      24813: inst = 32'd471859200;
      24814: inst = 32'd136314880;
      24815: inst = 32'd268468224;
      24816: inst = 32'd201347907;
      24817: inst = 32'd203459697;
      24818: inst = 32'd471859200;
      24819: inst = 32'd136314880;
      24820: inst = 32'd268468224;
      24821: inst = 32'd201347908;
      24822: inst = 32'd203455440;
      24823: inst = 32'd471859200;
      24824: inst = 32'd136314880;
      24825: inst = 32'd268468224;
      24826: inst = 32'd201347909;
      24827: inst = 32'd203451216;
      24828: inst = 32'd471859200;
      24829: inst = 32'd136314880;
      24830: inst = 32'd268468224;
      24831: inst = 32'd201347910;
      24832: inst = 32'd203451216;
      24833: inst = 32'd471859200;
      24834: inst = 32'd136314880;
      24835: inst = 32'd268468224;
      24836: inst = 32'd201347911;
      24837: inst = 32'd203451216;
      24838: inst = 32'd471859200;
      24839: inst = 32'd136314880;
      24840: inst = 32'd268468224;
      24841: inst = 32'd201347912;
      24842: inst = 32'd203451216;
      24843: inst = 32'd471859200;
      24844: inst = 32'd136314880;
      24845: inst = 32'd268468224;
      24846: inst = 32'd201347913;
      24847: inst = 32'd203451216;
      24848: inst = 32'd471859200;
      24849: inst = 32'd136314880;
      24850: inst = 32'd268468224;
      24851: inst = 32'd201347914;
      24852: inst = 32'd203451216;
      24853: inst = 32'd471859200;
      24854: inst = 32'd136314880;
      24855: inst = 32'd268468224;
      24856: inst = 32'd201347915;
      24857: inst = 32'd203451216;
      24858: inst = 32'd471859200;
      24859: inst = 32'd136314880;
      24860: inst = 32'd268468224;
      24861: inst = 32'd201347916;
      24862: inst = 32'd203451216;
      24863: inst = 32'd471859200;
      24864: inst = 32'd136314880;
      24865: inst = 32'd268468224;
      24866: inst = 32'd201347917;
      24867: inst = 32'd203451216;
      24868: inst = 32'd471859200;
      24869: inst = 32'd136314880;
      24870: inst = 32'd268468224;
      24871: inst = 32'd201347918;
      24872: inst = 32'd203451216;
      24873: inst = 32'd471859200;
      24874: inst = 32'd136314880;
      24875: inst = 32'd268468224;
      24876: inst = 32'd201347919;
      24877: inst = 32'd203451216;
      24878: inst = 32'd471859200;
      24879: inst = 32'd136314880;
      24880: inst = 32'd268468224;
      24881: inst = 32'd201347920;
      24882: inst = 32'd203451216;
      24883: inst = 32'd471859200;
      24884: inst = 32'd136314880;
      24885: inst = 32'd268468224;
      24886: inst = 32'd201347921;
      24887: inst = 32'd203451216;
      24888: inst = 32'd471859200;
      24889: inst = 32'd136314880;
      24890: inst = 32'd268468224;
      24891: inst = 32'd201347922;
      24892: inst = 32'd203451216;
      24893: inst = 32'd471859200;
      24894: inst = 32'd136314880;
      24895: inst = 32'd268468224;
      24896: inst = 32'd201347923;
      24897: inst = 32'd203451216;
      24898: inst = 32'd471859200;
      24899: inst = 32'd136314880;
      24900: inst = 32'd268468224;
      24901: inst = 32'd201347924;
      24902: inst = 32'd203451216;
      24903: inst = 32'd471859200;
      24904: inst = 32'd136314880;
      24905: inst = 32'd268468224;
      24906: inst = 32'd201347925;
      24907: inst = 32'd203451216;
      24908: inst = 32'd471859200;
      24909: inst = 32'd136314880;
      24910: inst = 32'd268468224;
      24911: inst = 32'd201347926;
      24912: inst = 32'd203451216;
      24913: inst = 32'd471859200;
      24914: inst = 32'd136314880;
      24915: inst = 32'd268468224;
      24916: inst = 32'd201347927;
      24917: inst = 32'd203451216;
      24918: inst = 32'd471859200;
      24919: inst = 32'd136314880;
      24920: inst = 32'd268468224;
      24921: inst = 32'd201347928;
      24922: inst = 32'd203451216;
      24923: inst = 32'd471859200;
      24924: inst = 32'd136314880;
      24925: inst = 32'd268468224;
      24926: inst = 32'd201347929;
      24927: inst = 32'd203451216;
      24928: inst = 32'd471859200;
      24929: inst = 32'd136314880;
      24930: inst = 32'd268468224;
      24931: inst = 32'd201347930;
      24932: inst = 32'd203451216;
      24933: inst = 32'd471859200;
      24934: inst = 32'd136314880;
      24935: inst = 32'd268468224;
      24936: inst = 32'd201347931;
      24937: inst = 32'd203451216;
      24938: inst = 32'd471859200;
      24939: inst = 32'd136314880;
      24940: inst = 32'd268468224;
      24941: inst = 32'd201347932;
      24942: inst = 32'd203451216;
      24943: inst = 32'd471859200;
      24944: inst = 32'd136314880;
      24945: inst = 32'd268468224;
      24946: inst = 32'd201347933;
      24947: inst = 32'd203451216;
      24948: inst = 32'd471859200;
      24949: inst = 32'd136314880;
      24950: inst = 32'd268468224;
      24951: inst = 32'd201347934;
      24952: inst = 32'd203451216;
      24953: inst = 32'd471859200;
      24954: inst = 32'd136314880;
      24955: inst = 32'd268468224;
      24956: inst = 32'd201347935;
      24957: inst = 32'd203451216;
      24958: inst = 32'd471859200;
      24959: inst = 32'd136314880;
      24960: inst = 32'd268468224;
      24961: inst = 32'd201347936;
      24962: inst = 32'd203451216;
      24963: inst = 32'd471859200;
      24964: inst = 32'd136314880;
      24965: inst = 32'd268468224;
      24966: inst = 32'd201347937;
      24967: inst = 32'd203451216;
      24968: inst = 32'd471859200;
      24969: inst = 32'd136314880;
      24970: inst = 32'd268468224;
      24971: inst = 32'd201347938;
      24972: inst = 32'd203451216;
      24973: inst = 32'd471859200;
      24974: inst = 32'd136314880;
      24975: inst = 32'd268468224;
      24976: inst = 32'd201347939;
      24977: inst = 32'd203451216;
      24978: inst = 32'd471859200;
      24979: inst = 32'd136314880;
      24980: inst = 32'd268468224;
      24981: inst = 32'd201347940;
      24982: inst = 32'd203451216;
      24983: inst = 32'd471859200;
      24984: inst = 32'd136314880;
      24985: inst = 32'd268468224;
      24986: inst = 32'd201347941;
      24987: inst = 32'd203451216;
      24988: inst = 32'd471859200;
      24989: inst = 32'd136314880;
      24990: inst = 32'd268468224;
      24991: inst = 32'd201347942;
      24992: inst = 32'd203451216;
      24993: inst = 32'd471859200;
      24994: inst = 32'd136314880;
      24995: inst = 32'd268468224;
      24996: inst = 32'd201347943;
      24997: inst = 32'd203451216;
      24998: inst = 32'd471859200;
      24999: inst = 32'd136314880;
      25000: inst = 32'd268468224;
      25001: inst = 32'd201347944;
      25002: inst = 32'd203451216;
      25003: inst = 32'd471859200;
      25004: inst = 32'd136314880;
      25005: inst = 32'd268468224;
      25006: inst = 32'd201347945;
      25007: inst = 32'd203451216;
      25008: inst = 32'd471859200;
      25009: inst = 32'd136314880;
      25010: inst = 32'd268468224;
      25011: inst = 32'd201347946;
      25012: inst = 32'd203451216;
      25013: inst = 32'd471859200;
      25014: inst = 32'd136314880;
      25015: inst = 32'd268468224;
      25016: inst = 32'd201347947;
      25017: inst = 32'd203451216;
      25018: inst = 32'd471859200;
      25019: inst = 32'd136314880;
      25020: inst = 32'd268468224;
      25021: inst = 32'd201347948;
      25022: inst = 32'd203451216;
      25023: inst = 32'd471859200;
      25024: inst = 32'd136314880;
      25025: inst = 32'd268468224;
      25026: inst = 32'd201347949;
      25027: inst = 32'd203451216;
      25028: inst = 32'd471859200;
      25029: inst = 32'd136314880;
      25030: inst = 32'd268468224;
      25031: inst = 32'd201347950;
      25032: inst = 32'd203451216;
      25033: inst = 32'd471859200;
      25034: inst = 32'd136314880;
      25035: inst = 32'd268468224;
      25036: inst = 32'd201347951;
      25037: inst = 32'd203451216;
      25038: inst = 32'd471859200;
      25039: inst = 32'd136314880;
      25040: inst = 32'd268468224;
      25041: inst = 32'd201347952;
      25042: inst = 32'd203451216;
      25043: inst = 32'd471859200;
      25044: inst = 32'd136314880;
      25045: inst = 32'd268468224;
      25046: inst = 32'd201347953;
      25047: inst = 32'd203451216;
      25048: inst = 32'd471859200;
      25049: inst = 32'd136314880;
      25050: inst = 32'd268468224;
      25051: inst = 32'd201347954;
      25052: inst = 32'd203451216;
      25053: inst = 32'd471859200;
      25054: inst = 32'd136314880;
      25055: inst = 32'd268468224;
      25056: inst = 32'd201347955;
      25057: inst = 32'd203451216;
      25058: inst = 32'd471859200;
      25059: inst = 32'd136314880;
      25060: inst = 32'd268468224;
      25061: inst = 32'd201347956;
      25062: inst = 32'd203451216;
      25063: inst = 32'd471859200;
      25064: inst = 32'd136314880;
      25065: inst = 32'd268468224;
      25066: inst = 32'd201347957;
      25067: inst = 32'd203451216;
      25068: inst = 32'd471859200;
      25069: inst = 32'd136314880;
      25070: inst = 32'd268468224;
      25071: inst = 32'd201347958;
      25072: inst = 32'd203451216;
      25073: inst = 32'd471859200;
      25074: inst = 32'd136314880;
      25075: inst = 32'd268468224;
      25076: inst = 32'd201347959;
      25077: inst = 32'd203451216;
      25078: inst = 32'd471859200;
      25079: inst = 32'd136314880;
      25080: inst = 32'd268468224;
      25081: inst = 32'd201347960;
      25082: inst = 32'd203451216;
      25083: inst = 32'd471859200;
      25084: inst = 32'd136314880;
      25085: inst = 32'd268468224;
      25086: inst = 32'd201347961;
      25087: inst = 32'd203451216;
      25088: inst = 32'd471859200;
      25089: inst = 32'd136314880;
      25090: inst = 32'd268468224;
      25091: inst = 32'd201347962;
      25092: inst = 32'd203453328;
      25093: inst = 32'd471859200;
      25094: inst = 32'd136314880;
      25095: inst = 32'd268468224;
      25096: inst = 32'd201347963;
      25097: inst = 32'd203459697;
      25098: inst = 32'd471859200;
      25099: inst = 32'd136314880;
      25100: inst = 32'd268468224;
      25101: inst = 32'd201347964;
      25102: inst = 32'd203459697;
      25103: inst = 32'd471859200;
      25104: inst = 32'd136314880;
      25105: inst = 32'd268468224;
      25106: inst = 32'd201347965;
      25107: inst = 32'd203457552;
      25108: inst = 32'd471859200;
      25109: inst = 32'd136314880;
      25110: inst = 32'd268468224;
      25111: inst = 32'd201347966;
      25112: inst = 32'd203444841;
      25113: inst = 32'd471859200;
      25114: inst = 32'd136314880;
      25115: inst = 32'd268468224;
      25116: inst = 32'd201347967;
      25117: inst = 32'd203442793;
      25118: inst = 32'd471859200;
      25119: inst = 32'd136314880;
      25120: inst = 32'd268468224;
      25121: inst = 32'd201347968;
      25122: inst = 32'd203446987;
      25123: inst = 32'd471859200;
      25124: inst = 32'd136314880;
      25125: inst = 32'd268468224;
      25126: inst = 32'd201347969;
      25127: inst = 32'd203455439;
      25128: inst = 32'd471859200;
      25129: inst = 32'd136314880;
      25130: inst = 32'd268468224;
      25131: inst = 32'd201347970;
      25132: inst = 32'd203442793;
      25133: inst = 32'd471859200;
      25134: inst = 32'd136314880;
      25135: inst = 32'd268468224;
      25136: inst = 32'd201347971;
      25137: inst = 32'd203442793;
      25138: inst = 32'd471859200;
      25139: inst = 32'd136314880;
      25140: inst = 32'd268468224;
      25141: inst = 32'd201347972;
      25142: inst = 32'd203442793;
      25143: inst = 32'd471859200;
      25144: inst = 32'd136314880;
      25145: inst = 32'd268468224;
      25146: inst = 32'd201347973;
      25147: inst = 32'd203457552;
      25148: inst = 32'd471859200;
      25149: inst = 32'd136314880;
      25150: inst = 32'd268468224;
      25151: inst = 32'd201347974;
      25152: inst = 32'd203459697;
      25153: inst = 32'd471859200;
      25154: inst = 32'd136314880;
      25155: inst = 32'd268468224;
      25156: inst = 32'd201347975;
      25157: inst = 32'd203459697;
      25158: inst = 32'd471859200;
      25159: inst = 32'd136314880;
      25160: inst = 32'd268468224;
      25161: inst = 32'd201347976;
      25162: inst = 32'd203459697;
      25163: inst = 32'd471859200;
      25164: inst = 32'd136314880;
      25165: inst = 32'd268468224;
      25166: inst = 32'd201347977;
      25167: inst = 32'd203444906;
      25168: inst = 32'd471859200;
      25169: inst = 32'd136314880;
      25170: inst = 32'd268468224;
      25171: inst = 32'd201347978;
      25172: inst = 32'd203451216;
      25173: inst = 32'd471859200;
      25174: inst = 32'd136314880;
      25175: inst = 32'd268468224;
      25176: inst = 32'd201347979;
      25177: inst = 32'd203451216;
      25178: inst = 32'd471859200;
      25179: inst = 32'd136314880;
      25180: inst = 32'd268468224;
      25181: inst = 32'd201347980;
      25182: inst = 32'd203451216;
      25183: inst = 32'd471859200;
      25184: inst = 32'd136314880;
      25185: inst = 32'd268468224;
      25186: inst = 32'd201347981;
      25187: inst = 32'd203451216;
      25188: inst = 32'd471859200;
      25189: inst = 32'd136314880;
      25190: inst = 32'd268468224;
      25191: inst = 32'd201347982;
      25192: inst = 32'd203451216;
      25193: inst = 32'd471859200;
      25194: inst = 32'd136314880;
      25195: inst = 32'd268468224;
      25196: inst = 32'd201347983;
      25197: inst = 32'd203451216;
      25198: inst = 32'd471859200;
      25199: inst = 32'd136314880;
      25200: inst = 32'd268468224;
      25201: inst = 32'd201347984;
      25202: inst = 32'd203451216;
      25203: inst = 32'd471859200;
      25204: inst = 32'd136314880;
      25205: inst = 32'd268468224;
      25206: inst = 32'd201347985;
      25207: inst = 32'd203451216;
      25208: inst = 32'd471859200;
      25209: inst = 32'd136314880;
      25210: inst = 32'd268468224;
      25211: inst = 32'd201347986;
      25212: inst = 32'd203451216;
      25213: inst = 32'd471859200;
      25214: inst = 32'd136314880;
      25215: inst = 32'd268468224;
      25216: inst = 32'd201347987;
      25217: inst = 32'd203451216;
      25218: inst = 32'd471859200;
      25219: inst = 32'd136314880;
      25220: inst = 32'd268468224;
      25221: inst = 32'd201347988;
      25222: inst = 32'd203451216;
      25223: inst = 32'd471859200;
      25224: inst = 32'd136314880;
      25225: inst = 32'd268468224;
      25226: inst = 32'd201347989;
      25227: inst = 32'd203451216;
      25228: inst = 32'd471859200;
      25229: inst = 32'd136314880;
      25230: inst = 32'd268468224;
      25231: inst = 32'd201347990;
      25232: inst = 32'd203444906;
      25233: inst = 32'd471859200;
      25234: inst = 32'd136314880;
      25235: inst = 32'd268468224;
      25236: inst = 32'd201347991;
      25237: inst = 32'd203459697;
      25238: inst = 32'd471859200;
      25239: inst = 32'd136314880;
      25240: inst = 32'd268468224;
      25241: inst = 32'd201347992;
      25242: inst = 32'd203459697;
      25243: inst = 32'd471859200;
      25244: inst = 32'd136314880;
      25245: inst = 32'd268468224;
      25246: inst = 32'd201347993;
      25247: inst = 32'd203459697;
      25248: inst = 32'd471859200;
      25249: inst = 32'd136314880;
      25250: inst = 32'd268468224;
      25251: inst = 32'd201347994;
      25252: inst = 32'd203457552;
      25253: inst = 32'd471859200;
      25254: inst = 32'd136314880;
      25255: inst = 32'd268468224;
      25256: inst = 32'd201347995;
      25257: inst = 32'd203442793;
      25258: inst = 32'd471859200;
      25259: inst = 32'd136314880;
      25260: inst = 32'd268468224;
      25261: inst = 32'd201347996;
      25262: inst = 32'd203442793;
      25263: inst = 32'd471859200;
      25264: inst = 32'd136314880;
      25265: inst = 32'd268468224;
      25266: inst = 32'd201347997;
      25267: inst = 32'd203442793;
      25268: inst = 32'd471859200;
      25269: inst = 32'd136314880;
      25270: inst = 32'd268468224;
      25271: inst = 32'd201347998;
      25272: inst = 32'd203455439;
      25273: inst = 32'd471859200;
      25274: inst = 32'd136314880;
      25275: inst = 32'd268468224;
      25276: inst = 32'd201347999;
      25277: inst = 32'd203446987;
      25278: inst = 32'd471859200;
      25279: inst = 32'd136314880;
      25280: inst = 32'd268468224;
      25281: inst = 32'd201348000;
      25282: inst = 32'd203442793;
      25283: inst = 32'd471859200;
      25284: inst = 32'd136314880;
      25285: inst = 32'd268468224;
      25286: inst = 32'd201348001;
      25287: inst = 32'd203444841;
      25288: inst = 32'd471859200;
      25289: inst = 32'd136314880;
      25290: inst = 32'd268468224;
      25291: inst = 32'd201348002;
      25292: inst = 32'd203457552;
      25293: inst = 32'd471859200;
      25294: inst = 32'd136314880;
      25295: inst = 32'd268468224;
      25296: inst = 32'd201348003;
      25297: inst = 32'd203459697;
      25298: inst = 32'd471859200;
      25299: inst = 32'd136314880;
      25300: inst = 32'd268468224;
      25301: inst = 32'd201348004;
      25302: inst = 32'd203459697;
      25303: inst = 32'd471859200;
      25304: inst = 32'd136314880;
      25305: inst = 32'd268468224;
      25306: inst = 32'd201348005;
      25307: inst = 32'd203453328;
      25308: inst = 32'd471859200;
      25309: inst = 32'd136314880;
      25310: inst = 32'd268468224;
      25311: inst = 32'd201348006;
      25312: inst = 32'd203451216;
      25313: inst = 32'd471859200;
      25314: inst = 32'd136314880;
      25315: inst = 32'd268468224;
      25316: inst = 32'd201348007;
      25317: inst = 32'd203451216;
      25318: inst = 32'd471859200;
      25319: inst = 32'd136314880;
      25320: inst = 32'd268468224;
      25321: inst = 32'd201348008;
      25322: inst = 32'd203451216;
      25323: inst = 32'd471859200;
      25324: inst = 32'd136314880;
      25325: inst = 32'd268468224;
      25326: inst = 32'd201348009;
      25327: inst = 32'd203451216;
      25328: inst = 32'd471859200;
      25329: inst = 32'd136314880;
      25330: inst = 32'd268468224;
      25331: inst = 32'd201348010;
      25332: inst = 32'd203451216;
      25333: inst = 32'd471859200;
      25334: inst = 32'd136314880;
      25335: inst = 32'd268468224;
      25336: inst = 32'd201348011;
      25337: inst = 32'd203451216;
      25338: inst = 32'd471859200;
      25339: inst = 32'd136314880;
      25340: inst = 32'd268468224;
      25341: inst = 32'd201348012;
      25342: inst = 32'd203451216;
      25343: inst = 32'd471859200;
      25344: inst = 32'd136314880;
      25345: inst = 32'd268468224;
      25346: inst = 32'd201348013;
      25347: inst = 32'd203451216;
      25348: inst = 32'd471859200;
      25349: inst = 32'd136314880;
      25350: inst = 32'd268468224;
      25351: inst = 32'd201348014;
      25352: inst = 32'd203451216;
      25353: inst = 32'd471859200;
      25354: inst = 32'd136314880;
      25355: inst = 32'd268468224;
      25356: inst = 32'd201348015;
      25357: inst = 32'd203451216;
      25358: inst = 32'd471859200;
      25359: inst = 32'd136314880;
      25360: inst = 32'd268468224;
      25361: inst = 32'd201348016;
      25362: inst = 32'd203451216;
      25363: inst = 32'd471859200;
      25364: inst = 32'd136314880;
      25365: inst = 32'd268468224;
      25366: inst = 32'd201348017;
      25367: inst = 32'd203451216;
      25368: inst = 32'd471859200;
      25369: inst = 32'd136314880;
      25370: inst = 32'd268468224;
      25371: inst = 32'd201348018;
      25372: inst = 32'd203451216;
      25373: inst = 32'd471859200;
      25374: inst = 32'd136314880;
      25375: inst = 32'd268468224;
      25376: inst = 32'd201348019;
      25377: inst = 32'd203451216;
      25378: inst = 32'd471859200;
      25379: inst = 32'd136314880;
      25380: inst = 32'd268468224;
      25381: inst = 32'd201348020;
      25382: inst = 32'd203451216;
      25383: inst = 32'd471859200;
      25384: inst = 32'd136314880;
      25385: inst = 32'd268468224;
      25386: inst = 32'd201348021;
      25387: inst = 32'd203451216;
      25388: inst = 32'd471859200;
      25389: inst = 32'd136314880;
      25390: inst = 32'd268468224;
      25391: inst = 32'd201348022;
      25392: inst = 32'd203451216;
      25393: inst = 32'd471859200;
      25394: inst = 32'd136314880;
      25395: inst = 32'd268468224;
      25396: inst = 32'd201348023;
      25397: inst = 32'd203451216;
      25398: inst = 32'd471859200;
      25399: inst = 32'd136314880;
      25400: inst = 32'd268468224;
      25401: inst = 32'd201348024;
      25402: inst = 32'd203451216;
      25403: inst = 32'd471859200;
      25404: inst = 32'd136314880;
      25405: inst = 32'd268468224;
      25406: inst = 32'd201348025;
      25407: inst = 32'd203451216;
      25408: inst = 32'd471859200;
      25409: inst = 32'd136314880;
      25410: inst = 32'd268468224;
      25411: inst = 32'd201348026;
      25412: inst = 32'd203451216;
      25413: inst = 32'd471859200;
      25414: inst = 32'd136314880;
      25415: inst = 32'd268468224;
      25416: inst = 32'd201348027;
      25417: inst = 32'd203451216;
      25418: inst = 32'd471859200;
      25419: inst = 32'd136314880;
      25420: inst = 32'd268468224;
      25421: inst = 32'd201348028;
      25422: inst = 32'd203451216;
      25423: inst = 32'd471859200;
      25424: inst = 32'd136314880;
      25425: inst = 32'd268468224;
      25426: inst = 32'd201348029;
      25427: inst = 32'd203451216;
      25428: inst = 32'd471859200;
      25429: inst = 32'd136314880;
      25430: inst = 32'd268468224;
      25431: inst = 32'd201348030;
      25432: inst = 32'd203451216;
      25433: inst = 32'd471859200;
      25434: inst = 32'd136314880;
      25435: inst = 32'd268468224;
      25436: inst = 32'd201348031;
      25437: inst = 32'd203451216;
      25438: inst = 32'd471859200;
      25439: inst = 32'd136314880;
      25440: inst = 32'd268468224;
      25441: inst = 32'd201348032;
      25442: inst = 32'd203451216;
      25443: inst = 32'd471859200;
      25444: inst = 32'd136314880;
      25445: inst = 32'd268468224;
      25446: inst = 32'd201348033;
      25447: inst = 32'd203451216;
      25448: inst = 32'd471859200;
      25449: inst = 32'd136314880;
      25450: inst = 32'd268468224;
      25451: inst = 32'd201348034;
      25452: inst = 32'd203451216;
      25453: inst = 32'd471859200;
      25454: inst = 32'd136314880;
      25455: inst = 32'd268468224;
      25456: inst = 32'd201348035;
      25457: inst = 32'd203451216;
      25458: inst = 32'd471859200;
      25459: inst = 32'd136314880;
      25460: inst = 32'd268468224;
      25461: inst = 32'd201348036;
      25462: inst = 32'd203451216;
      25463: inst = 32'd471859200;
      25464: inst = 32'd136314880;
      25465: inst = 32'd268468224;
      25466: inst = 32'd201348037;
      25467: inst = 32'd203451216;
      25468: inst = 32'd471859200;
      25469: inst = 32'd136314880;
      25470: inst = 32'd268468224;
      25471: inst = 32'd201348038;
      25472: inst = 32'd203451216;
      25473: inst = 32'd471859200;
      25474: inst = 32'd136314880;
      25475: inst = 32'd268468224;
      25476: inst = 32'd201348039;
      25477: inst = 32'd203451216;
      25478: inst = 32'd471859200;
      25479: inst = 32'd136314880;
      25480: inst = 32'd268468224;
      25481: inst = 32'd201348040;
      25482: inst = 32'd203451216;
      25483: inst = 32'd471859200;
      25484: inst = 32'd136314880;
      25485: inst = 32'd268468224;
      25486: inst = 32'd201348041;
      25487: inst = 32'd203451216;
      25488: inst = 32'd471859200;
      25489: inst = 32'd136314880;
      25490: inst = 32'd268468224;
      25491: inst = 32'd201348042;
      25492: inst = 32'd203451216;
      25493: inst = 32'd471859200;
      25494: inst = 32'd136314880;
      25495: inst = 32'd268468224;
      25496: inst = 32'd201348043;
      25497: inst = 32'd203451216;
      25498: inst = 32'd471859200;
      25499: inst = 32'd136314880;
      25500: inst = 32'd268468224;
      25501: inst = 32'd201348044;
      25502: inst = 32'd203451216;
      25503: inst = 32'd471859200;
      25504: inst = 32'd136314880;
      25505: inst = 32'd268468224;
      25506: inst = 32'd201348045;
      25507: inst = 32'd203451216;
      25508: inst = 32'd471859200;
      25509: inst = 32'd136314880;
      25510: inst = 32'd268468224;
      25511: inst = 32'd201348046;
      25512: inst = 32'd203451216;
      25513: inst = 32'd471859200;
      25514: inst = 32'd136314880;
      25515: inst = 32'd268468224;
      25516: inst = 32'd201348047;
      25517: inst = 32'd203451216;
      25518: inst = 32'd471859200;
      25519: inst = 32'd136314880;
      25520: inst = 32'd268468224;
      25521: inst = 32'd201348048;
      25522: inst = 32'd203451216;
      25523: inst = 32'd471859200;
      25524: inst = 32'd136314880;
      25525: inst = 32'd268468224;
      25526: inst = 32'd201348049;
      25527: inst = 32'd203451216;
      25528: inst = 32'd471859200;
      25529: inst = 32'd136314880;
      25530: inst = 32'd268468224;
      25531: inst = 32'd201348050;
      25532: inst = 32'd203451216;
      25533: inst = 32'd471859200;
      25534: inst = 32'd136314880;
      25535: inst = 32'd268468224;
      25536: inst = 32'd201348051;
      25537: inst = 32'd203451216;
      25538: inst = 32'd471859200;
      25539: inst = 32'd136314880;
      25540: inst = 32'd268468224;
      25541: inst = 32'd201348052;
      25542: inst = 32'd203451216;
      25543: inst = 32'd471859200;
      25544: inst = 32'd136314880;
      25545: inst = 32'd268468224;
      25546: inst = 32'd201348053;
      25547: inst = 32'd203451216;
      25548: inst = 32'd471859200;
      25549: inst = 32'd136314880;
      25550: inst = 32'd268468224;
      25551: inst = 32'd201348054;
      25552: inst = 32'd203451216;
      25553: inst = 32'd471859200;
      25554: inst = 32'd136314880;
      25555: inst = 32'd268468224;
      25556: inst = 32'd201348055;
      25557: inst = 32'd203451216;
      25558: inst = 32'd471859200;
      25559: inst = 32'd136314880;
      25560: inst = 32'd268468224;
      25561: inst = 32'd201348056;
      25562: inst = 32'd203451216;
      25563: inst = 32'd471859200;
      25564: inst = 32'd136314880;
      25565: inst = 32'd268468224;
      25566: inst = 32'd201348057;
      25567: inst = 32'd203451248;
      25568: inst = 32'd471859200;
      25569: inst = 32'd136314880;
      25570: inst = 32'd268468224;
      25571: inst = 32'd201348058;
      25572: inst = 32'd203459665;
      25573: inst = 32'd471859200;
      25574: inst = 32'd136314880;
      25575: inst = 32'd268468224;
      25576: inst = 32'd201348059;
      25577: inst = 32'd203459697;
      25578: inst = 32'd471859200;
      25579: inst = 32'd136314880;
      25580: inst = 32'd268468224;
      25581: inst = 32'd201348060;
      25582: inst = 32'd203459665;
      25583: inst = 32'd471859200;
      25584: inst = 32'd136314880;
      25585: inst = 32'd268468224;
      25586: inst = 32'd201348061;
      25587: inst = 32'd203446987;
      25588: inst = 32'd471859200;
      25589: inst = 32'd136314880;
      25590: inst = 32'd268468224;
      25591: inst = 32'd201348062;
      25592: inst = 32'd203442793;
      25593: inst = 32'd471859200;
      25594: inst = 32'd136314880;
      25595: inst = 32'd268468224;
      25596: inst = 32'd201348063;
      25597: inst = 32'd203442793;
      25598: inst = 32'd471859200;
      25599: inst = 32'd136314880;
      25600: inst = 32'd268468224;
      25601: inst = 32'd201348064;
      25602: inst = 32'd203453294;
      25603: inst = 32'd471859200;
      25604: inst = 32'd136314880;
      25605: inst = 32'd268468224;
      25606: inst = 32'd201348065;
      25607: inst = 32'd203455439;
      25608: inst = 32'd471859200;
      25609: inst = 32'd136314880;
      25610: inst = 32'd268468224;
      25611: inst = 32'd201348066;
      25612: inst = 32'd203442793;
      25613: inst = 32'd471859200;
      25614: inst = 32'd136314880;
      25615: inst = 32'd268468224;
      25616: inst = 32'd201348067;
      25617: inst = 32'd203442793;
      25618: inst = 32'd471859200;
      25619: inst = 32'd136314880;
      25620: inst = 32'd268468224;
      25621: inst = 32'd201348068;
      25622: inst = 32'd203446954;
      25623: inst = 32'd471859200;
      25624: inst = 32'd136314880;
      25625: inst = 32'd268468224;
      25626: inst = 32'd201348069;
      25627: inst = 32'd203459697;
      25628: inst = 32'd471859200;
      25629: inst = 32'd136314880;
      25630: inst = 32'd268468224;
      25631: inst = 32'd201348070;
      25632: inst = 32'd203459697;
      25633: inst = 32'd471859200;
      25634: inst = 32'd136314880;
      25635: inst = 32'd268468224;
      25636: inst = 32'd201348071;
      25637: inst = 32'd203459697;
      25638: inst = 32'd471859200;
      25639: inst = 32'd136314880;
      25640: inst = 32'd268468224;
      25641: inst = 32'd201348072;
      25642: inst = 32'd203457585;
      25643: inst = 32'd471859200;
      25644: inst = 32'd136314880;
      25645: inst = 32'd268468224;
      25646: inst = 32'd201348073;
      25647: inst = 32'd203444874;
      25648: inst = 32'd471859200;
      25649: inst = 32'd136314880;
      25650: inst = 32'd268468224;
      25651: inst = 32'd201348074;
      25652: inst = 32'd203451216;
      25653: inst = 32'd471859200;
      25654: inst = 32'd136314880;
      25655: inst = 32'd268468224;
      25656: inst = 32'd201348075;
      25657: inst = 32'd203451216;
      25658: inst = 32'd471859200;
      25659: inst = 32'd136314880;
      25660: inst = 32'd268468224;
      25661: inst = 32'd201348076;
      25662: inst = 32'd203451216;
      25663: inst = 32'd471859200;
      25664: inst = 32'd136314880;
      25665: inst = 32'd268468224;
      25666: inst = 32'd201348077;
      25667: inst = 32'd203451216;
      25668: inst = 32'd471859200;
      25669: inst = 32'd136314880;
      25670: inst = 32'd268468224;
      25671: inst = 32'd201348078;
      25672: inst = 32'd203451216;
      25673: inst = 32'd471859200;
      25674: inst = 32'd136314880;
      25675: inst = 32'd268468224;
      25676: inst = 32'd201348079;
      25677: inst = 32'd203451216;
      25678: inst = 32'd471859200;
      25679: inst = 32'd136314880;
      25680: inst = 32'd268468224;
      25681: inst = 32'd201348080;
      25682: inst = 32'd203451216;
      25683: inst = 32'd471859200;
      25684: inst = 32'd136314880;
      25685: inst = 32'd268468224;
      25686: inst = 32'd201348081;
      25687: inst = 32'd203451216;
      25688: inst = 32'd471859200;
      25689: inst = 32'd136314880;
      25690: inst = 32'd268468224;
      25691: inst = 32'd201348082;
      25692: inst = 32'd203451216;
      25693: inst = 32'd471859200;
      25694: inst = 32'd136314880;
      25695: inst = 32'd268468224;
      25696: inst = 32'd201348083;
      25697: inst = 32'd203451216;
      25698: inst = 32'd471859200;
      25699: inst = 32'd136314880;
      25700: inst = 32'd268468224;
      25701: inst = 32'd201348084;
      25702: inst = 32'd203451216;
      25703: inst = 32'd471859200;
      25704: inst = 32'd136314880;
      25705: inst = 32'd268468224;
      25706: inst = 32'd201348085;
      25707: inst = 32'd203451216;
      25708: inst = 32'd471859200;
      25709: inst = 32'd136314880;
      25710: inst = 32'd268468224;
      25711: inst = 32'd201348086;
      25712: inst = 32'd203444874;
      25713: inst = 32'd471859200;
      25714: inst = 32'd136314880;
      25715: inst = 32'd268468224;
      25716: inst = 32'd201348087;
      25717: inst = 32'd203457585;
      25718: inst = 32'd471859200;
      25719: inst = 32'd136314880;
      25720: inst = 32'd268468224;
      25721: inst = 32'd201348088;
      25722: inst = 32'd203459697;
      25723: inst = 32'd471859200;
      25724: inst = 32'd136314880;
      25725: inst = 32'd268468224;
      25726: inst = 32'd201348089;
      25727: inst = 32'd203459697;
      25728: inst = 32'd471859200;
      25729: inst = 32'd136314880;
      25730: inst = 32'd268468224;
      25731: inst = 32'd201348090;
      25732: inst = 32'd203459697;
      25733: inst = 32'd471859200;
      25734: inst = 32'd136314880;
      25735: inst = 32'd268468224;
      25736: inst = 32'd201348091;
      25737: inst = 32'd203446954;
      25738: inst = 32'd471859200;
      25739: inst = 32'd136314880;
      25740: inst = 32'd268468224;
      25741: inst = 32'd201348092;
      25742: inst = 32'd203442793;
      25743: inst = 32'd471859200;
      25744: inst = 32'd136314880;
      25745: inst = 32'd268468224;
      25746: inst = 32'd201348093;
      25747: inst = 32'd203442793;
      25748: inst = 32'd471859200;
      25749: inst = 32'd136314880;
      25750: inst = 32'd268468224;
      25751: inst = 32'd201348094;
      25752: inst = 32'd203455439;
      25753: inst = 32'd471859200;
      25754: inst = 32'd136314880;
      25755: inst = 32'd268468224;
      25756: inst = 32'd201348095;
      25757: inst = 32'd203453294;
      25758: inst = 32'd471859200;
      25759: inst = 32'd136314880;
      25760: inst = 32'd268468224;
      25761: inst = 32'd201348096;
      25762: inst = 32'd203442793;
      25763: inst = 32'd471859200;
      25764: inst = 32'd136314880;
      25765: inst = 32'd268468224;
      25766: inst = 32'd201348097;
      25767: inst = 32'd203442793;
      25768: inst = 32'd471859200;
      25769: inst = 32'd136314880;
      25770: inst = 32'd268468224;
      25771: inst = 32'd201348098;
      25772: inst = 32'd203446987;
      25773: inst = 32'd471859200;
      25774: inst = 32'd136314880;
      25775: inst = 32'd268468224;
      25776: inst = 32'd201348099;
      25777: inst = 32'd203459665;
      25778: inst = 32'd471859200;
      25779: inst = 32'd136314880;
      25780: inst = 32'd268468224;
      25781: inst = 32'd201348100;
      25782: inst = 32'd203459697;
      25783: inst = 32'd471859200;
      25784: inst = 32'd136314880;
      25785: inst = 32'd268468224;
      25786: inst = 32'd201348101;
      25787: inst = 32'd203459665;
      25788: inst = 32'd471859200;
      25789: inst = 32'd136314880;
      25790: inst = 32'd268468224;
      25791: inst = 32'd201348102;
      25792: inst = 32'd203451248;
      25793: inst = 32'd471859200;
      25794: inst = 32'd136314880;
      25795: inst = 32'd268468224;
      25796: inst = 32'd201348103;
      25797: inst = 32'd203451216;
      25798: inst = 32'd471859200;
      25799: inst = 32'd136314880;
      25800: inst = 32'd268468224;
      25801: inst = 32'd201348104;
      25802: inst = 32'd203451216;
      25803: inst = 32'd471859200;
      25804: inst = 32'd136314880;
      25805: inst = 32'd268468224;
      25806: inst = 32'd201348105;
      25807: inst = 32'd203451216;
      25808: inst = 32'd471859200;
      25809: inst = 32'd136314880;
      25810: inst = 32'd268468224;
      25811: inst = 32'd201348106;
      25812: inst = 32'd203451216;
      25813: inst = 32'd471859200;
      25814: inst = 32'd136314880;
      25815: inst = 32'd268468224;
      25816: inst = 32'd201348107;
      25817: inst = 32'd203451216;
      25818: inst = 32'd471859200;
      25819: inst = 32'd136314880;
      25820: inst = 32'd268468224;
      25821: inst = 32'd201348108;
      25822: inst = 32'd203451216;
      25823: inst = 32'd471859200;
      25824: inst = 32'd136314880;
      25825: inst = 32'd268468224;
      25826: inst = 32'd201348109;
      25827: inst = 32'd203451216;
      25828: inst = 32'd471859200;
      25829: inst = 32'd136314880;
      25830: inst = 32'd268468224;
      25831: inst = 32'd201348110;
      25832: inst = 32'd203451216;
      25833: inst = 32'd471859200;
      25834: inst = 32'd136314880;
      25835: inst = 32'd268468224;
      25836: inst = 32'd201348111;
      25837: inst = 32'd203451216;
      25838: inst = 32'd471859200;
      25839: inst = 32'd136314880;
      25840: inst = 32'd268468224;
      25841: inst = 32'd201348112;
      25842: inst = 32'd203451216;
      25843: inst = 32'd471859200;
      25844: inst = 32'd136314880;
      25845: inst = 32'd268468224;
      25846: inst = 32'd201348113;
      25847: inst = 32'd203451216;
      25848: inst = 32'd471859200;
      25849: inst = 32'd136314880;
      25850: inst = 32'd268468224;
      25851: inst = 32'd201348114;
      25852: inst = 32'd203451216;
      25853: inst = 32'd471859200;
      25854: inst = 32'd136314880;
      25855: inst = 32'd268468224;
      25856: inst = 32'd201348115;
      25857: inst = 32'd203451216;
      25858: inst = 32'd471859200;
      25859: inst = 32'd136314880;
      25860: inst = 32'd268468224;
      25861: inst = 32'd201348116;
      25862: inst = 32'd203451216;
      25863: inst = 32'd471859200;
      25864: inst = 32'd136314880;
      25865: inst = 32'd268468224;
      25866: inst = 32'd201348117;
      25867: inst = 32'd203451216;
      25868: inst = 32'd471859200;
      25869: inst = 32'd136314880;
      25870: inst = 32'd268468224;
      25871: inst = 32'd201348118;
      25872: inst = 32'd203451216;
      25873: inst = 32'd471859200;
      25874: inst = 32'd136314880;
      25875: inst = 32'd268468224;
      25876: inst = 32'd201348119;
      25877: inst = 32'd203451216;
      25878: inst = 32'd471859200;
      25879: inst = 32'd136314880;
      25880: inst = 32'd268468224;
      25881: inst = 32'd201348120;
      25882: inst = 32'd203451216;
      25883: inst = 32'd471859200;
      25884: inst = 32'd136314880;
      25885: inst = 32'd268468224;
      25886: inst = 32'd201348121;
      25887: inst = 32'd203451216;
      25888: inst = 32'd471859200;
      25889: inst = 32'd136314880;
      25890: inst = 32'd268468224;
      25891: inst = 32'd201348122;
      25892: inst = 32'd203451216;
      25893: inst = 32'd471859200;
      25894: inst = 32'd136314880;
      25895: inst = 32'd268468224;
      25896: inst = 32'd201348123;
      25897: inst = 32'd203451216;
      25898: inst = 32'd471859200;
      25899: inst = 32'd136314880;
      25900: inst = 32'd268468224;
      25901: inst = 32'd201348124;
      25902: inst = 32'd203451216;
      25903: inst = 32'd471859200;
      25904: inst = 32'd136314880;
      25905: inst = 32'd268468224;
      25906: inst = 32'd201348125;
      25907: inst = 32'd203451216;
      25908: inst = 32'd471859200;
      25909: inst = 32'd136314880;
      25910: inst = 32'd268468224;
      25911: inst = 32'd201348126;
      25912: inst = 32'd203451216;
      25913: inst = 32'd471859200;
      25914: inst = 32'd136314880;
      25915: inst = 32'd268468224;
      25916: inst = 32'd201348127;
      25917: inst = 32'd203451216;
      25918: inst = 32'd471859200;
      25919: inst = 32'd136314880;
      25920: inst = 32'd268468224;
      25921: inst = 32'd201348128;
      25922: inst = 32'd203451216;
      25923: inst = 32'd471859200;
      25924: inst = 32'd136314880;
      25925: inst = 32'd268468224;
      25926: inst = 32'd201348129;
      25927: inst = 32'd203451216;
      25928: inst = 32'd471859200;
      25929: inst = 32'd136314880;
      25930: inst = 32'd268468224;
      25931: inst = 32'd201348130;
      25932: inst = 32'd203451216;
      25933: inst = 32'd471859200;
      25934: inst = 32'd136314880;
      25935: inst = 32'd268468224;
      25936: inst = 32'd201348131;
      25937: inst = 32'd203451216;
      25938: inst = 32'd471859200;
      25939: inst = 32'd136314880;
      25940: inst = 32'd268468224;
      25941: inst = 32'd201348132;
      25942: inst = 32'd203451216;
      25943: inst = 32'd471859200;
      25944: inst = 32'd136314880;
      25945: inst = 32'd268468224;
      25946: inst = 32'd201348133;
      25947: inst = 32'd203451216;
      25948: inst = 32'd471859200;
      25949: inst = 32'd136314880;
      25950: inst = 32'd268468224;
      25951: inst = 32'd201348134;
      25952: inst = 32'd203451216;
      25953: inst = 32'd471859200;
      25954: inst = 32'd136314880;
      25955: inst = 32'd268468224;
      25956: inst = 32'd201348135;
      25957: inst = 32'd203451216;
      25958: inst = 32'd471859200;
      25959: inst = 32'd136314880;
      25960: inst = 32'd268468224;
      25961: inst = 32'd201348136;
      25962: inst = 32'd203451216;
      25963: inst = 32'd471859200;
      25964: inst = 32'd136314880;
      25965: inst = 32'd268468224;
      25966: inst = 32'd201348137;
      25967: inst = 32'd203451216;
      25968: inst = 32'd471859200;
      25969: inst = 32'd136314880;
      25970: inst = 32'd268468224;
      25971: inst = 32'd201348138;
      25972: inst = 32'd203451216;
      25973: inst = 32'd471859200;
      25974: inst = 32'd136314880;
      25975: inst = 32'd268468224;
      25976: inst = 32'd201348139;
      25977: inst = 32'd203451216;
      25978: inst = 32'd471859200;
      25979: inst = 32'd136314880;
      25980: inst = 32'd268468224;
      25981: inst = 32'd201348140;
      25982: inst = 32'd203451216;
      25983: inst = 32'd471859200;
      25984: inst = 32'd136314880;
      25985: inst = 32'd268468224;
      25986: inst = 32'd201348141;
      25987: inst = 32'd203451216;
      25988: inst = 32'd471859200;
      25989: inst = 32'd136314880;
      25990: inst = 32'd268468224;
      25991: inst = 32'd201348142;
      25992: inst = 32'd203451216;
      25993: inst = 32'd471859200;
      25994: inst = 32'd136314880;
      25995: inst = 32'd268468224;
      25996: inst = 32'd201348143;
      25997: inst = 32'd203451216;
      25998: inst = 32'd471859200;
      25999: inst = 32'd136314880;
      26000: inst = 32'd268468224;
      26001: inst = 32'd201348144;
      26002: inst = 32'd203451216;
      26003: inst = 32'd471859200;
      26004: inst = 32'd136314880;
      26005: inst = 32'd268468224;
      26006: inst = 32'd201348145;
      26007: inst = 32'd203451216;
      26008: inst = 32'd471859200;
      26009: inst = 32'd136314880;
      26010: inst = 32'd268468224;
      26011: inst = 32'd201348146;
      26012: inst = 32'd203451216;
      26013: inst = 32'd471859200;
      26014: inst = 32'd136314880;
      26015: inst = 32'd268468224;
      26016: inst = 32'd201348147;
      26017: inst = 32'd203451216;
      26018: inst = 32'd471859200;
      26019: inst = 32'd136314880;
      26020: inst = 32'd268468224;
      26021: inst = 32'd201348148;
      26022: inst = 32'd203451216;
      26023: inst = 32'd471859200;
      26024: inst = 32'd136314880;
      26025: inst = 32'd268468224;
      26026: inst = 32'd201348149;
      26027: inst = 32'd203451216;
      26028: inst = 32'd471859200;
      26029: inst = 32'd136314880;
      26030: inst = 32'd268468224;
      26031: inst = 32'd201348150;
      26032: inst = 32'd203451216;
      26033: inst = 32'd471859200;
      26034: inst = 32'd136314880;
      26035: inst = 32'd268468224;
      26036: inst = 32'd201348151;
      26037: inst = 32'd203451216;
      26038: inst = 32'd471859200;
      26039: inst = 32'd136314880;
      26040: inst = 32'd268468224;
      26041: inst = 32'd201348152;
      26042: inst = 32'd203451216;
      26043: inst = 32'd471859200;
      26044: inst = 32'd136314880;
      26045: inst = 32'd268468224;
      26046: inst = 32'd201348153;
      26047: inst = 32'd203457585;
      26048: inst = 32'd471859200;
      26049: inst = 32'd136314880;
      26050: inst = 32'd268468224;
      26051: inst = 32'd201348154;
      26052: inst = 32'd203459697;
      26053: inst = 32'd471859200;
      26054: inst = 32'd136314880;
      26055: inst = 32'd268468224;
      26056: inst = 32'd201348155;
      26057: inst = 32'd203459697;
      26058: inst = 32'd471859200;
      26059: inst = 32'd136314880;
      26060: inst = 32'd268468224;
      26061: inst = 32'd201348156;
      26062: inst = 32'd203451213;
      26063: inst = 32'd471859200;
      26064: inst = 32'd136314880;
      26065: inst = 32'd268468224;
      26066: inst = 32'd201348157;
      26067: inst = 32'd203442793;
      26068: inst = 32'd471859200;
      26069: inst = 32'd136314880;
      26070: inst = 32'd268468224;
      26071: inst = 32'd201348158;
      26072: inst = 32'd203442793;
      26073: inst = 32'd471859200;
      26074: inst = 32'd136314880;
      26075: inst = 32'd268468224;
      26076: inst = 32'd201348159;
      26077: inst = 32'd203442793;
      26078: inst = 32'd471859200;
      26079: inst = 32'd136314880;
      26080: inst = 32'd268468224;
      26081: inst = 32'd201348160;
      26082: inst = 32'd203457584;
      26083: inst = 32'd471859200;
      26084: inst = 32'd136314880;
      26085: inst = 32'd268468224;
      26086: inst = 32'd201348161;
      26087: inst = 32'd203455439;
      26088: inst = 32'd471859200;
      26089: inst = 32'd136314880;
      26090: inst = 32'd268468224;
      26091: inst = 32'd201348162;
      26092: inst = 32'd203442793;
      26093: inst = 32'd471859200;
      26094: inst = 32'd136314880;
      26095: inst = 32'd268468224;
      26096: inst = 32'd201348163;
      26097: inst = 32'd203442793;
      26098: inst = 32'd471859200;
      26099: inst = 32'd136314880;
      26100: inst = 32'd268468224;
      26101: inst = 32'd201348164;
      26102: inst = 32'd203451213;
      26103: inst = 32'd471859200;
      26104: inst = 32'd136314880;
      26105: inst = 32'd268468224;
      26106: inst = 32'd201348165;
      26107: inst = 32'd203459697;
      26108: inst = 32'd471859200;
      26109: inst = 32'd136314880;
      26110: inst = 32'd268468224;
      26111: inst = 32'd201348166;
      26112: inst = 32'd203459697;
      26113: inst = 32'd471859200;
      26114: inst = 32'd136314880;
      26115: inst = 32'd268468224;
      26116: inst = 32'd201348167;
      26117: inst = 32'd203459697;
      26118: inst = 32'd471859200;
      26119: inst = 32'd136314880;
      26120: inst = 32'd268468224;
      26121: inst = 32'd201348168;
      26122: inst = 32'd203455439;
      26123: inst = 32'd471859200;
      26124: inst = 32'd136314880;
      26125: inst = 32'd268468224;
      26126: inst = 32'd201348169;
      26127: inst = 32'd203444874;
      26128: inst = 32'd471859200;
      26129: inst = 32'd136314880;
      26130: inst = 32'd268468224;
      26131: inst = 32'd201348170;
      26132: inst = 32'd203451216;
      26133: inst = 32'd471859200;
      26134: inst = 32'd136314880;
      26135: inst = 32'd268468224;
      26136: inst = 32'd201348171;
      26137: inst = 32'd203451216;
      26138: inst = 32'd471859200;
      26139: inst = 32'd136314880;
      26140: inst = 32'd268468224;
      26141: inst = 32'd201348172;
      26142: inst = 32'd203451216;
      26143: inst = 32'd471859200;
      26144: inst = 32'd136314880;
      26145: inst = 32'd268468224;
      26146: inst = 32'd201348173;
      26147: inst = 32'd203451216;
      26148: inst = 32'd471859200;
      26149: inst = 32'd136314880;
      26150: inst = 32'd268468224;
      26151: inst = 32'd201348174;
      26152: inst = 32'd203451216;
      26153: inst = 32'd471859200;
      26154: inst = 32'd136314880;
      26155: inst = 32'd268468224;
      26156: inst = 32'd201348175;
      26157: inst = 32'd203451216;
      26158: inst = 32'd471859200;
      26159: inst = 32'd136314880;
      26160: inst = 32'd268468224;
      26161: inst = 32'd201348176;
      26162: inst = 32'd203451216;
      26163: inst = 32'd471859200;
      26164: inst = 32'd136314880;
      26165: inst = 32'd268468224;
      26166: inst = 32'd201348177;
      26167: inst = 32'd203451216;
      26168: inst = 32'd471859200;
      26169: inst = 32'd136314880;
      26170: inst = 32'd268468224;
      26171: inst = 32'd201348178;
      26172: inst = 32'd203451216;
      26173: inst = 32'd471859200;
      26174: inst = 32'd136314880;
      26175: inst = 32'd268468224;
      26176: inst = 32'd201348179;
      26177: inst = 32'd203451216;
      26178: inst = 32'd471859200;
      26179: inst = 32'd136314880;
      26180: inst = 32'd268468224;
      26181: inst = 32'd201348180;
      26182: inst = 32'd203451216;
      26183: inst = 32'd471859200;
      26184: inst = 32'd136314880;
      26185: inst = 32'd268468224;
      26186: inst = 32'd201348181;
      26187: inst = 32'd203451216;
      26188: inst = 32'd471859200;
      26189: inst = 32'd136314880;
      26190: inst = 32'd268468224;
      26191: inst = 32'd201348182;
      26192: inst = 32'd203444874;
      26193: inst = 32'd471859200;
      26194: inst = 32'd136314880;
      26195: inst = 32'd268468224;
      26196: inst = 32'd201348183;
      26197: inst = 32'd203455439;
      26198: inst = 32'd471859200;
      26199: inst = 32'd136314880;
      26200: inst = 32'd268468224;
      26201: inst = 32'd201348184;
      26202: inst = 32'd203459697;
      26203: inst = 32'd471859200;
      26204: inst = 32'd136314880;
      26205: inst = 32'd268468224;
      26206: inst = 32'd201348185;
      26207: inst = 32'd203459697;
      26208: inst = 32'd471859200;
      26209: inst = 32'd136314880;
      26210: inst = 32'd268468224;
      26211: inst = 32'd201348186;
      26212: inst = 32'd203459697;
      26213: inst = 32'd471859200;
      26214: inst = 32'd136314880;
      26215: inst = 32'd268468224;
      26216: inst = 32'd201348187;
      26217: inst = 32'd203451213;
      26218: inst = 32'd471859200;
      26219: inst = 32'd136314880;
      26220: inst = 32'd268468224;
      26221: inst = 32'd201348188;
      26222: inst = 32'd203442793;
      26223: inst = 32'd471859200;
      26224: inst = 32'd136314880;
      26225: inst = 32'd268468224;
      26226: inst = 32'd201348189;
      26227: inst = 32'd203442793;
      26228: inst = 32'd471859200;
      26229: inst = 32'd136314880;
      26230: inst = 32'd268468224;
      26231: inst = 32'd201348190;
      26232: inst = 32'd203455439;
      26233: inst = 32'd471859200;
      26234: inst = 32'd136314880;
      26235: inst = 32'd268468224;
      26236: inst = 32'd201348191;
      26237: inst = 32'd203457584;
      26238: inst = 32'd471859200;
      26239: inst = 32'd136314880;
      26240: inst = 32'd268468224;
      26241: inst = 32'd201348192;
      26242: inst = 32'd203442793;
      26243: inst = 32'd471859200;
      26244: inst = 32'd136314880;
      26245: inst = 32'd268468224;
      26246: inst = 32'd201348193;
      26247: inst = 32'd203442793;
      26248: inst = 32'd471859200;
      26249: inst = 32'd136314880;
      26250: inst = 32'd268468224;
      26251: inst = 32'd201348194;
      26252: inst = 32'd203442793;
      26253: inst = 32'd471859200;
      26254: inst = 32'd136314880;
      26255: inst = 32'd268468224;
      26256: inst = 32'd201348195;
      26257: inst = 32'd203451213;
      26258: inst = 32'd471859200;
      26259: inst = 32'd136314880;
      26260: inst = 32'd268468224;
      26261: inst = 32'd201348196;
      26262: inst = 32'd203459697;
      26263: inst = 32'd471859200;
      26264: inst = 32'd136314880;
      26265: inst = 32'd268468224;
      26266: inst = 32'd201348197;
      26267: inst = 32'd203459697;
      26268: inst = 32'd471859200;
      26269: inst = 32'd136314880;
      26270: inst = 32'd268468224;
      26271: inst = 32'd201348198;
      26272: inst = 32'd203457585;
      26273: inst = 32'd471859200;
      26274: inst = 32'd136314880;
      26275: inst = 32'd268468224;
      26276: inst = 32'd201348199;
      26277: inst = 32'd203451216;
      26278: inst = 32'd471859200;
      26279: inst = 32'd136314880;
      26280: inst = 32'd268468224;
      26281: inst = 32'd201348200;
      26282: inst = 32'd203451216;
      26283: inst = 32'd471859200;
      26284: inst = 32'd136314880;
      26285: inst = 32'd268468224;
      26286: inst = 32'd201348201;
      26287: inst = 32'd203451216;
      26288: inst = 32'd471859200;
      26289: inst = 32'd136314880;
      26290: inst = 32'd268468224;
      26291: inst = 32'd201348202;
      26292: inst = 32'd203451216;
      26293: inst = 32'd471859200;
      26294: inst = 32'd136314880;
      26295: inst = 32'd268468224;
      26296: inst = 32'd201348203;
      26297: inst = 32'd203451216;
      26298: inst = 32'd471859200;
      26299: inst = 32'd136314880;
      26300: inst = 32'd268468224;
      26301: inst = 32'd201348204;
      26302: inst = 32'd203451216;
      26303: inst = 32'd471859200;
      26304: inst = 32'd136314880;
      26305: inst = 32'd268468224;
      26306: inst = 32'd201348205;
      26307: inst = 32'd203451216;
      26308: inst = 32'd471859200;
      26309: inst = 32'd136314880;
      26310: inst = 32'd268468224;
      26311: inst = 32'd201348206;
      26312: inst = 32'd203451216;
      26313: inst = 32'd471859200;
      26314: inst = 32'd136314880;
      26315: inst = 32'd268468224;
      26316: inst = 32'd201348207;
      26317: inst = 32'd203451216;
      26318: inst = 32'd471859200;
      26319: inst = 32'd136314880;
      26320: inst = 32'd268468224;
      26321: inst = 32'd201348208;
      26322: inst = 32'd203451216;
      26323: inst = 32'd471859200;
      26324: inst = 32'd136314880;
      26325: inst = 32'd268468224;
      26326: inst = 32'd201348209;
      26327: inst = 32'd203451216;
      26328: inst = 32'd471859200;
      26329: inst = 32'd136314880;
      26330: inst = 32'd268468224;
      26331: inst = 32'd201348210;
      26332: inst = 32'd203451216;
      26333: inst = 32'd471859200;
      26334: inst = 32'd136314880;
      26335: inst = 32'd268468224;
      26336: inst = 32'd201348211;
      26337: inst = 32'd203451216;
      26338: inst = 32'd471859200;
      26339: inst = 32'd136314880;
      26340: inst = 32'd268468224;
      26341: inst = 32'd201348212;
      26342: inst = 32'd203451216;
      26343: inst = 32'd471859200;
      26344: inst = 32'd136314880;
      26345: inst = 32'd268468224;
      26346: inst = 32'd201348213;
      26347: inst = 32'd203451216;
      26348: inst = 32'd471859200;
      26349: inst = 32'd136314880;
      26350: inst = 32'd268468224;
      26351: inst = 32'd201348214;
      26352: inst = 32'd203451216;
      26353: inst = 32'd471859200;
      26354: inst = 32'd136314880;
      26355: inst = 32'd268468224;
      26356: inst = 32'd201348215;
      26357: inst = 32'd203451216;
      26358: inst = 32'd471859200;
      26359: inst = 32'd136314880;
      26360: inst = 32'd268468224;
      26361: inst = 32'd201348216;
      26362: inst = 32'd203451216;
      26363: inst = 32'd471859200;
      26364: inst = 32'd136314880;
      26365: inst = 32'd268468224;
      26366: inst = 32'd201348217;
      26367: inst = 32'd203451216;
      26368: inst = 32'd471859200;
      26369: inst = 32'd136314880;
      26370: inst = 32'd268468224;
      26371: inst = 32'd201348218;
      26372: inst = 32'd203451216;
      26373: inst = 32'd471859200;
      26374: inst = 32'd136314880;
      26375: inst = 32'd268468224;
      26376: inst = 32'd201348219;
      26377: inst = 32'd203451216;
      26378: inst = 32'd471859200;
      26379: inst = 32'd136314880;
      26380: inst = 32'd268468224;
      26381: inst = 32'd201348220;
      26382: inst = 32'd203451216;
      26383: inst = 32'd471859200;
      26384: inst = 32'd136314880;
      26385: inst = 32'd268468224;
      26386: inst = 32'd201348221;
      26387: inst = 32'd203451216;
      26388: inst = 32'd471859200;
      26389: inst = 32'd136314880;
      26390: inst = 32'd268468224;
      26391: inst = 32'd201348222;
      26392: inst = 32'd203451216;
      26393: inst = 32'd471859200;
      26394: inst = 32'd136314880;
      26395: inst = 32'd268468224;
      26396: inst = 32'd201348223;
      26397: inst = 32'd203451216;
      26398: inst = 32'd471859200;
      26399: inst = 32'd136314880;
      26400: inst = 32'd268468224;
      26401: inst = 32'd201348224;
      26402: inst = 32'd203451216;
      26403: inst = 32'd471859200;
      26404: inst = 32'd136314880;
      26405: inst = 32'd268468224;
      26406: inst = 32'd201348225;
      26407: inst = 32'd203451216;
      26408: inst = 32'd471859200;
      26409: inst = 32'd136314880;
      26410: inst = 32'd268468224;
      26411: inst = 32'd201348226;
      26412: inst = 32'd203451216;
      26413: inst = 32'd471859200;
      26414: inst = 32'd136314880;
      26415: inst = 32'd268468224;
      26416: inst = 32'd201348227;
      26417: inst = 32'd203451216;
      26418: inst = 32'd471859200;
      26419: inst = 32'd136314880;
      26420: inst = 32'd268468224;
      26421: inst = 32'd201348228;
      26422: inst = 32'd203451216;
      26423: inst = 32'd471859200;
      26424: inst = 32'd136314880;
      26425: inst = 32'd268468224;
      26426: inst = 32'd201348229;
      26427: inst = 32'd203451216;
      26428: inst = 32'd471859200;
      26429: inst = 32'd136314880;
      26430: inst = 32'd268468224;
      26431: inst = 32'd201348230;
      26432: inst = 32'd203451216;
      26433: inst = 32'd471859200;
      26434: inst = 32'd136314880;
      26435: inst = 32'd268468224;
      26436: inst = 32'd201348231;
      26437: inst = 32'd203451216;
      26438: inst = 32'd471859200;
      26439: inst = 32'd136314880;
      26440: inst = 32'd268468224;
      26441: inst = 32'd201348232;
      26442: inst = 32'd203451216;
      26443: inst = 32'd471859200;
      26444: inst = 32'd136314880;
      26445: inst = 32'd268468224;
      26446: inst = 32'd201348233;
      26447: inst = 32'd203451216;
      26448: inst = 32'd471859200;
      26449: inst = 32'd136314880;
      26450: inst = 32'd268468224;
      26451: inst = 32'd201348234;
      26452: inst = 32'd203451216;
      26453: inst = 32'd471859200;
      26454: inst = 32'd136314880;
      26455: inst = 32'd268468224;
      26456: inst = 32'd201348235;
      26457: inst = 32'd203451216;
      26458: inst = 32'd471859200;
      26459: inst = 32'd136314880;
      26460: inst = 32'd268468224;
      26461: inst = 32'd201348236;
      26462: inst = 32'd203451216;
      26463: inst = 32'd471859200;
      26464: inst = 32'd136314880;
      26465: inst = 32'd268468224;
      26466: inst = 32'd201348237;
      26467: inst = 32'd203451216;
      26468: inst = 32'd471859200;
      26469: inst = 32'd136314880;
      26470: inst = 32'd268468224;
      26471: inst = 32'd201348238;
      26472: inst = 32'd203451216;
      26473: inst = 32'd471859200;
      26474: inst = 32'd136314880;
      26475: inst = 32'd268468224;
      26476: inst = 32'd201348239;
      26477: inst = 32'd203451216;
      26478: inst = 32'd471859200;
      26479: inst = 32'd136314880;
      26480: inst = 32'd268468224;
      26481: inst = 32'd201348240;
      26482: inst = 32'd203451216;
      26483: inst = 32'd471859200;
      26484: inst = 32'd136314880;
      26485: inst = 32'd268468224;
      26486: inst = 32'd201348241;
      26487: inst = 32'd203451216;
      26488: inst = 32'd471859200;
      26489: inst = 32'd136314880;
      26490: inst = 32'd268468224;
      26491: inst = 32'd201348242;
      26492: inst = 32'd203451216;
      26493: inst = 32'd471859200;
      26494: inst = 32'd136314880;
      26495: inst = 32'd268468224;
      26496: inst = 32'd201348243;
      26497: inst = 32'd203451216;
      26498: inst = 32'd471859200;
      26499: inst = 32'd136314880;
      26500: inst = 32'd268468224;
      26501: inst = 32'd201348244;
      26502: inst = 32'd203451216;
      26503: inst = 32'd471859200;
      26504: inst = 32'd136314880;
      26505: inst = 32'd268468224;
      26506: inst = 32'd201348245;
      26507: inst = 32'd203451216;
      26508: inst = 32'd471859200;
      26509: inst = 32'd136314880;
      26510: inst = 32'd268468224;
      26511: inst = 32'd201348246;
      26512: inst = 32'd203451216;
      26513: inst = 32'd471859200;
      26514: inst = 32'd136314880;
      26515: inst = 32'd268468224;
      26516: inst = 32'd201348247;
      26517: inst = 32'd203451216;
      26518: inst = 32'd471859200;
      26519: inst = 32'd136314880;
      26520: inst = 32'd268468224;
      26521: inst = 32'd201348248;
      26522: inst = 32'd203455473;
      26523: inst = 32'd471859200;
      26524: inst = 32'd136314880;
      26525: inst = 32'd268468224;
      26526: inst = 32'd201348249;
      26527: inst = 32'd203459697;
      26528: inst = 32'd471859200;
      26529: inst = 32'd136314880;
      26530: inst = 32'd268468224;
      26531: inst = 32'd201348250;
      26532: inst = 32'd203459697;
      26533: inst = 32'd471859200;
      26534: inst = 32'd136314880;
      26535: inst = 32'd268468224;
      26536: inst = 32'd201348251;
      26537: inst = 32'd203455471;
      26538: inst = 32'd471859200;
      26539: inst = 32'd136314880;
      26540: inst = 32'd268468224;
      26541: inst = 32'd201348252;
      26542: inst = 32'd203444841;
      26543: inst = 32'd471859200;
      26544: inst = 32'd136314880;
      26545: inst = 32'd268468224;
      26546: inst = 32'd201348253;
      26547: inst = 32'd203442793;
      26548: inst = 32'd471859200;
      26549: inst = 32'd136314880;
      26550: inst = 32'd268468224;
      26551: inst = 32'd201348254;
      26552: inst = 32'd203442793;
      26553: inst = 32'd471859200;
      26554: inst = 32'd136314880;
      26555: inst = 32'd268468224;
      26556: inst = 32'd201348255;
      26557: inst = 32'd203447019;
      26558: inst = 32'd471859200;
      26559: inst = 32'd136314880;
      26560: inst = 32'd268468224;
      26561: inst = 32'd201348256;
      26562: inst = 32'd203442793;
      26563: inst = 32'd471859200;
      26564: inst = 32'd136314880;
      26565: inst = 32'd268468224;
      26566: inst = 32'd201348257;
      26567: inst = 32'd203442793;
      26568: inst = 32'd471859200;
      26569: inst = 32'd136314880;
      26570: inst = 32'd268468224;
      26571: inst = 32'd201348258;
      26572: inst = 32'd203442793;
      26573: inst = 32'd471859200;
      26574: inst = 32'd136314880;
      26575: inst = 32'd268468224;
      26576: inst = 32'd201348259;
      26577: inst = 32'd203442793;
      26578: inst = 32'd471859200;
      26579: inst = 32'd136314880;
      26580: inst = 32'd268468224;
      26581: inst = 32'd201348260;
      26582: inst = 32'd203457552;
      26583: inst = 32'd471859200;
      26584: inst = 32'd136314880;
      26585: inst = 32'd268468224;
      26586: inst = 32'd201348261;
      26587: inst = 32'd203459697;
      26588: inst = 32'd471859200;
      26589: inst = 32'd136314880;
      26590: inst = 32'd268468224;
      26591: inst = 32'd201348262;
      26592: inst = 32'd203459697;
      26593: inst = 32'd471859200;
      26594: inst = 32'd136314880;
      26595: inst = 32'd268468224;
      26596: inst = 32'd201348263;
      26597: inst = 32'd203459697;
      26598: inst = 32'd471859200;
      26599: inst = 32'd136314880;
      26600: inst = 32'd268468224;
      26601: inst = 32'd201348264;
      26602: inst = 32'd203451246;
      26603: inst = 32'd471859200;
      26604: inst = 32'd136314880;
      26605: inst = 32'd268468224;
      26606: inst = 32'd201348265;
      26607: inst = 32'd203444874;
      26608: inst = 32'd471859200;
      26609: inst = 32'd136314880;
      26610: inst = 32'd268468224;
      26611: inst = 32'd201348266;
      26612: inst = 32'd203451216;
      26613: inst = 32'd471859200;
      26614: inst = 32'd136314880;
      26615: inst = 32'd268468224;
      26616: inst = 32'd201348267;
      26617: inst = 32'd203451216;
      26618: inst = 32'd471859200;
      26619: inst = 32'd136314880;
      26620: inst = 32'd268468224;
      26621: inst = 32'd201348268;
      26622: inst = 32'd203451216;
      26623: inst = 32'd471859200;
      26624: inst = 32'd136314880;
      26625: inst = 32'd268468224;
      26626: inst = 32'd201348269;
      26627: inst = 32'd203451216;
      26628: inst = 32'd471859200;
      26629: inst = 32'd136314880;
      26630: inst = 32'd268468224;
      26631: inst = 32'd201348270;
      26632: inst = 32'd203451216;
      26633: inst = 32'd471859200;
      26634: inst = 32'd136314880;
      26635: inst = 32'd268468224;
      26636: inst = 32'd201348271;
      26637: inst = 32'd203451216;
      26638: inst = 32'd471859200;
      26639: inst = 32'd136314880;
      26640: inst = 32'd268468224;
      26641: inst = 32'd201348272;
      26642: inst = 32'd203451216;
      26643: inst = 32'd471859200;
      26644: inst = 32'd136314880;
      26645: inst = 32'd268468224;
      26646: inst = 32'd201348273;
      26647: inst = 32'd203451216;
      26648: inst = 32'd471859200;
      26649: inst = 32'd136314880;
      26650: inst = 32'd268468224;
      26651: inst = 32'd201348274;
      26652: inst = 32'd203451216;
      26653: inst = 32'd471859200;
      26654: inst = 32'd136314880;
      26655: inst = 32'd268468224;
      26656: inst = 32'd201348275;
      26657: inst = 32'd203451216;
      26658: inst = 32'd471859200;
      26659: inst = 32'd136314880;
      26660: inst = 32'd268468224;
      26661: inst = 32'd201348276;
      26662: inst = 32'd203451216;
      26663: inst = 32'd471859200;
      26664: inst = 32'd136314880;
      26665: inst = 32'd268468224;
      26666: inst = 32'd201348277;
      26667: inst = 32'd203451216;
      26668: inst = 32'd471859200;
      26669: inst = 32'd136314880;
      26670: inst = 32'd268468224;
      26671: inst = 32'd201348278;
      26672: inst = 32'd203444874;
      26673: inst = 32'd471859200;
      26674: inst = 32'd136314880;
      26675: inst = 32'd268468224;
      26676: inst = 32'd201348279;
      26677: inst = 32'd203451246;
      26678: inst = 32'd471859200;
      26679: inst = 32'd136314880;
      26680: inst = 32'd268468224;
      26681: inst = 32'd201348280;
      26682: inst = 32'd203459697;
      26683: inst = 32'd471859200;
      26684: inst = 32'd136314880;
      26685: inst = 32'd268468224;
      26686: inst = 32'd201348281;
      26687: inst = 32'd203459697;
      26688: inst = 32'd471859200;
      26689: inst = 32'd136314880;
      26690: inst = 32'd268468224;
      26691: inst = 32'd201348282;
      26692: inst = 32'd203459697;
      26693: inst = 32'd471859200;
      26694: inst = 32'd136314880;
      26695: inst = 32'd268468224;
      26696: inst = 32'd201348283;
      26697: inst = 32'd203457552;
      26698: inst = 32'd471859200;
      26699: inst = 32'd136314880;
      26700: inst = 32'd268468224;
      26701: inst = 32'd201348284;
      26702: inst = 32'd203442793;
      26703: inst = 32'd471859200;
      26704: inst = 32'd136314880;
      26705: inst = 32'd268468224;
      26706: inst = 32'd201348285;
      26707: inst = 32'd203442793;
      26708: inst = 32'd471859200;
      26709: inst = 32'd136314880;
      26710: inst = 32'd268468224;
      26711: inst = 32'd201348286;
      26712: inst = 32'd203442793;
      26713: inst = 32'd471859200;
      26714: inst = 32'd136314880;
      26715: inst = 32'd268468224;
      26716: inst = 32'd201348287;
      26717: inst = 32'd203442793;
      26718: inst = 32'd471859200;
      26719: inst = 32'd136314880;
      26720: inst = 32'd268468224;
      26721: inst = 32'd201348288;
      26722: inst = 32'd203447019;
      26723: inst = 32'd471859200;
      26724: inst = 32'd136314880;
      26725: inst = 32'd268468224;
      26726: inst = 32'd201348289;
      26727: inst = 32'd203442793;
      26728: inst = 32'd471859200;
      26729: inst = 32'd136314880;
      26730: inst = 32'd268468224;
      26731: inst = 32'd201348290;
      26732: inst = 32'd203442793;
      26733: inst = 32'd471859200;
      26734: inst = 32'd136314880;
      26735: inst = 32'd268468224;
      26736: inst = 32'd201348291;
      26737: inst = 32'd203444841;
      26738: inst = 32'd471859200;
      26739: inst = 32'd136314880;
      26740: inst = 32'd268468224;
      26741: inst = 32'd201348292;
      26742: inst = 32'd203455471;
      26743: inst = 32'd471859200;
      26744: inst = 32'd136314880;
      26745: inst = 32'd268468224;
      26746: inst = 32'd201348293;
      26747: inst = 32'd203459697;
      26748: inst = 32'd471859200;
      26749: inst = 32'd136314880;
      26750: inst = 32'd268468224;
      26751: inst = 32'd201348294;
      26752: inst = 32'd203459697;
      26753: inst = 32'd471859200;
      26754: inst = 32'd136314880;
      26755: inst = 32'd268468224;
      26756: inst = 32'd201348295;
      26757: inst = 32'd203455473;
      26758: inst = 32'd471859200;
      26759: inst = 32'd136314880;
      26760: inst = 32'd268468224;
      26761: inst = 32'd201348296;
      26762: inst = 32'd203451216;
      26763: inst = 32'd471859200;
      26764: inst = 32'd136314880;
      26765: inst = 32'd268468224;
      26766: inst = 32'd201348297;
      26767: inst = 32'd203451216;
      26768: inst = 32'd471859200;
      26769: inst = 32'd136314880;
      26770: inst = 32'd268468224;
      26771: inst = 32'd201348298;
      26772: inst = 32'd203451216;
      26773: inst = 32'd471859200;
      26774: inst = 32'd136314880;
      26775: inst = 32'd268468224;
      26776: inst = 32'd201348299;
      26777: inst = 32'd203451216;
      26778: inst = 32'd471859200;
      26779: inst = 32'd136314880;
      26780: inst = 32'd268468224;
      26781: inst = 32'd201348300;
      26782: inst = 32'd203451216;
      26783: inst = 32'd471859200;
      26784: inst = 32'd136314880;
      26785: inst = 32'd268468224;
      26786: inst = 32'd201348301;
      26787: inst = 32'd203451216;
      26788: inst = 32'd471859200;
      26789: inst = 32'd136314880;
      26790: inst = 32'd268468224;
      26791: inst = 32'd201348302;
      26792: inst = 32'd203451216;
      26793: inst = 32'd471859200;
      26794: inst = 32'd136314880;
      26795: inst = 32'd268468224;
      26796: inst = 32'd201348303;
      26797: inst = 32'd203451216;
      26798: inst = 32'd471859200;
      26799: inst = 32'd136314880;
      26800: inst = 32'd268468224;
      26801: inst = 32'd201348304;
      26802: inst = 32'd203451216;
      26803: inst = 32'd471859200;
      26804: inst = 32'd136314880;
      26805: inst = 32'd268468224;
      26806: inst = 32'd201348305;
      26807: inst = 32'd203451216;
      26808: inst = 32'd471859200;
      26809: inst = 32'd136314880;
      26810: inst = 32'd268468224;
      26811: inst = 32'd201348306;
      26812: inst = 32'd203451216;
      26813: inst = 32'd471859200;
      26814: inst = 32'd136314880;
      26815: inst = 32'd268468224;
      26816: inst = 32'd201348307;
      26817: inst = 32'd203451216;
      26818: inst = 32'd471859200;
      26819: inst = 32'd136314880;
      26820: inst = 32'd268468224;
      26821: inst = 32'd201348308;
      26822: inst = 32'd203451216;
      26823: inst = 32'd471859200;
      26824: inst = 32'd136314880;
      26825: inst = 32'd268468224;
      26826: inst = 32'd201348309;
      26827: inst = 32'd203451216;
      26828: inst = 32'd471859200;
      26829: inst = 32'd136314880;
      26830: inst = 32'd268468224;
      26831: inst = 32'd201348310;
      26832: inst = 32'd203451216;
      26833: inst = 32'd471859200;
      26834: inst = 32'd136314880;
      26835: inst = 32'd268468224;
      26836: inst = 32'd201348311;
      26837: inst = 32'd203451216;
      26838: inst = 32'd471859200;
      26839: inst = 32'd136314880;
      26840: inst = 32'd268468224;
      26841: inst = 32'd201348312;
      26842: inst = 32'd203451216;
      26843: inst = 32'd471859200;
      26844: inst = 32'd136314880;
      26845: inst = 32'd268468224;
      26846: inst = 32'd201348313;
      26847: inst = 32'd203451216;
      26848: inst = 32'd471859200;
      26849: inst = 32'd136314880;
      26850: inst = 32'd268468224;
      26851: inst = 32'd201348314;
      26852: inst = 32'd203451216;
      26853: inst = 32'd471859200;
      26854: inst = 32'd136314880;
      26855: inst = 32'd268468224;
      26856: inst = 32'd201348315;
      26857: inst = 32'd203451216;
      26858: inst = 32'd471859200;
      26859: inst = 32'd136314880;
      26860: inst = 32'd268468224;
      26861: inst = 32'd201348316;
      26862: inst = 32'd203451216;
      26863: inst = 32'd471859200;
      26864: inst = 32'd136314880;
      26865: inst = 32'd268468224;
      26866: inst = 32'd201348317;
      26867: inst = 32'd203451216;
      26868: inst = 32'd471859200;
      26869: inst = 32'd136314880;
      26870: inst = 32'd268468224;
      26871: inst = 32'd201348318;
      26872: inst = 32'd203451216;
      26873: inst = 32'd471859200;
      26874: inst = 32'd136314880;
      26875: inst = 32'd268468224;
      26876: inst = 32'd201348319;
      26877: inst = 32'd203451216;
      26878: inst = 32'd471859200;
      26879: inst = 32'd136314880;
      26880: inst = 32'd268468224;
      26881: inst = 32'd201348320;
      26882: inst = 32'd203451216;
      26883: inst = 32'd471859200;
      26884: inst = 32'd136314880;
      26885: inst = 32'd268468224;
      26886: inst = 32'd201348321;
      26887: inst = 32'd203451216;
      26888: inst = 32'd471859200;
      26889: inst = 32'd136314880;
      26890: inst = 32'd268468224;
      26891: inst = 32'd201348322;
      26892: inst = 32'd203451216;
      26893: inst = 32'd471859200;
      26894: inst = 32'd136314880;
      26895: inst = 32'd268468224;
      26896: inst = 32'd201348323;
      26897: inst = 32'd203451216;
      26898: inst = 32'd471859200;
      26899: inst = 32'd136314880;
      26900: inst = 32'd268468224;
      26901: inst = 32'd201348324;
      26902: inst = 32'd203451216;
      26903: inst = 32'd471859200;
      26904: inst = 32'd136314880;
      26905: inst = 32'd268468224;
      26906: inst = 32'd201348325;
      26907: inst = 32'd203451216;
      26908: inst = 32'd471859200;
      26909: inst = 32'd136314880;
      26910: inst = 32'd268468224;
      26911: inst = 32'd201348326;
      26912: inst = 32'd203451216;
      26913: inst = 32'd471859200;
      26914: inst = 32'd136314880;
      26915: inst = 32'd268468224;
      26916: inst = 32'd201348327;
      26917: inst = 32'd203451216;
      26918: inst = 32'd471859200;
      26919: inst = 32'd136314880;
      26920: inst = 32'd268468224;
      26921: inst = 32'd201348328;
      26922: inst = 32'd203451216;
      26923: inst = 32'd471859200;
      26924: inst = 32'd136314880;
      26925: inst = 32'd268468224;
      26926: inst = 32'd201348329;
      26927: inst = 32'd203451216;
      26928: inst = 32'd471859200;
      26929: inst = 32'd136314880;
      26930: inst = 32'd268468224;
      26931: inst = 32'd201348330;
      26932: inst = 32'd203451216;
      26933: inst = 32'd471859200;
      26934: inst = 32'd136314880;
      26935: inst = 32'd268468224;
      26936: inst = 32'd201348331;
      26937: inst = 32'd203451216;
      26938: inst = 32'd471859200;
      26939: inst = 32'd136314880;
      26940: inst = 32'd268468224;
      26941: inst = 32'd201348332;
      26942: inst = 32'd203451216;
      26943: inst = 32'd471859200;
      26944: inst = 32'd136314880;
      26945: inst = 32'd268468224;
      26946: inst = 32'd201348333;
      26947: inst = 32'd203451216;
      26948: inst = 32'd471859200;
      26949: inst = 32'd136314880;
      26950: inst = 32'd268468224;
      26951: inst = 32'd201348334;
      26952: inst = 32'd203451216;
      26953: inst = 32'd471859200;
      26954: inst = 32'd136314880;
      26955: inst = 32'd268468224;
      26956: inst = 32'd201348335;
      26957: inst = 32'd203451216;
      26958: inst = 32'd471859200;
      26959: inst = 32'd136314880;
      26960: inst = 32'd268468224;
      26961: inst = 32'd201348336;
      26962: inst = 32'd203451216;
      26963: inst = 32'd471859200;
      26964: inst = 32'd136314880;
      26965: inst = 32'd268468224;
      26966: inst = 32'd201348337;
      26967: inst = 32'd203451216;
      26968: inst = 32'd471859200;
      26969: inst = 32'd136314880;
      26970: inst = 32'd268468224;
      26971: inst = 32'd201348338;
      26972: inst = 32'd203451216;
      26973: inst = 32'd471859200;
      26974: inst = 32'd136314880;
      26975: inst = 32'd268468224;
      26976: inst = 32'd201348339;
      26977: inst = 32'd203451216;
      26978: inst = 32'd471859200;
      26979: inst = 32'd136314880;
      26980: inst = 32'd268468224;
      26981: inst = 32'd201348340;
      26982: inst = 32'd203451216;
      26983: inst = 32'd471859200;
      26984: inst = 32'd136314880;
      26985: inst = 32'd268468224;
      26986: inst = 32'd201348341;
      26987: inst = 32'd203451216;
      26988: inst = 32'd471859200;
      26989: inst = 32'd136314880;
      26990: inst = 32'd268468224;
      26991: inst = 32'd201348342;
      26992: inst = 32'd203451216;
      26993: inst = 32'd471859200;
      26994: inst = 32'd136314880;
      26995: inst = 32'd268468224;
      26996: inst = 32'd201348343;
      26997: inst = 32'd203453360;
      26998: inst = 32'd471859200;
      26999: inst = 32'd136314880;
      27000: inst = 32'd268468224;
      27001: inst = 32'd201348344;
      27002: inst = 32'd203459697;
      27003: inst = 32'd471859200;
      27004: inst = 32'd136314880;
      27005: inst = 32'd268468224;
      27006: inst = 32'd201348345;
      27007: inst = 32'd203459697;
      27008: inst = 32'd471859200;
      27009: inst = 32'd136314880;
      27010: inst = 32'd268468224;
      27011: inst = 32'd201348346;
      27012: inst = 32'd203459665;
      27013: inst = 32'd471859200;
      27014: inst = 32'd136314880;
      27015: inst = 32'd268468224;
      27016: inst = 32'd201348347;
      27017: inst = 32'd203444906;
      27018: inst = 32'd471859200;
      27019: inst = 32'd136314880;
      27020: inst = 32'd268468224;
      27021: inst = 32'd201348348;
      27022: inst = 32'd203442793;
      27023: inst = 32'd471859200;
      27024: inst = 32'd136314880;
      27025: inst = 32'd268468224;
      27026: inst = 32'd201348349;
      27027: inst = 32'd203442793;
      27028: inst = 32'd471859200;
      27029: inst = 32'd136314880;
      27030: inst = 32'd268468224;
      27031: inst = 32'd201348350;
      27032: inst = 32'd203442793;
      27033: inst = 32'd471859200;
      27034: inst = 32'd136314880;
      27035: inst = 32'd268468224;
      27036: inst = 32'd201348351;
      27037: inst = 32'd203453358;
      27038: inst = 32'd471859200;
      27039: inst = 32'd136314880;
      27040: inst = 32'd268468224;
      27041: inst = 32'd201348352;
      27042: inst = 32'd203459697;
      27043: inst = 32'd471859200;
      27044: inst = 32'd136314880;
      27045: inst = 32'd268468224;
      27046: inst = 32'd201348353;
      27047: inst = 32'd203455439;
      27048: inst = 32'd471859200;
      27049: inst = 32'd136314880;
      27050: inst = 32'd268468224;
      27051: inst = 32'd201348354;
      27052: inst = 32'd203442793;
      27053: inst = 32'd471859200;
      27054: inst = 32'd136314880;
      27055: inst = 32'd268468224;
      27056: inst = 32'd201348355;
      27057: inst = 32'd203444906;
      27058: inst = 32'd471859200;
      27059: inst = 32'd136314880;
      27060: inst = 32'd268468224;
      27061: inst = 32'd201348356;
      27062: inst = 32'd203459697;
      27063: inst = 32'd471859200;
      27064: inst = 32'd136314880;
      27065: inst = 32'd268468224;
      27066: inst = 32'd201348357;
      27067: inst = 32'd203459697;
      27068: inst = 32'd471859200;
      27069: inst = 32'd136314880;
      27070: inst = 32'd268468224;
      27071: inst = 32'd201348358;
      27072: inst = 32'd203459697;
      27073: inst = 32'd471859200;
      27074: inst = 32'd136314880;
      27075: inst = 32'd268468224;
      27076: inst = 32'd201348359;
      27077: inst = 32'd203459697;
      27078: inst = 32'd471859200;
      27079: inst = 32'd136314880;
      27080: inst = 32'd268468224;
      27081: inst = 32'd201348360;
      27082: inst = 32'd203449133;
      27083: inst = 32'd471859200;
      27084: inst = 32'd136314880;
      27085: inst = 32'd268468224;
      27086: inst = 32'd201348361;
      27087: inst = 32'd203444874;
      27088: inst = 32'd471859200;
      27089: inst = 32'd136314880;
      27090: inst = 32'd268468224;
      27091: inst = 32'd201348362;
      27092: inst = 32'd203451216;
      27093: inst = 32'd471859200;
      27094: inst = 32'd136314880;
      27095: inst = 32'd268468224;
      27096: inst = 32'd201348363;
      27097: inst = 32'd203451216;
      27098: inst = 32'd471859200;
      27099: inst = 32'd136314880;
      27100: inst = 32'd268468224;
      27101: inst = 32'd201348364;
      27102: inst = 32'd203451216;
      27103: inst = 32'd471859200;
      27104: inst = 32'd136314880;
      27105: inst = 32'd268468224;
      27106: inst = 32'd201348365;
      27107: inst = 32'd203451216;
      27108: inst = 32'd471859200;
      27109: inst = 32'd136314880;
      27110: inst = 32'd268468224;
      27111: inst = 32'd201348366;
      27112: inst = 32'd203451216;
      27113: inst = 32'd471859200;
      27114: inst = 32'd136314880;
      27115: inst = 32'd268468224;
      27116: inst = 32'd201348367;
      27117: inst = 32'd203451216;
      27118: inst = 32'd471859200;
      27119: inst = 32'd136314880;
      27120: inst = 32'd268468224;
      27121: inst = 32'd201348368;
      27122: inst = 32'd203451216;
      27123: inst = 32'd471859200;
      27124: inst = 32'd136314880;
      27125: inst = 32'd268468224;
      27126: inst = 32'd201348369;
      27127: inst = 32'd203451216;
      27128: inst = 32'd471859200;
      27129: inst = 32'd136314880;
      27130: inst = 32'd268468224;
      27131: inst = 32'd201348370;
      27132: inst = 32'd203451216;
      27133: inst = 32'd471859200;
      27134: inst = 32'd136314880;
      27135: inst = 32'd268468224;
      27136: inst = 32'd201348371;
      27137: inst = 32'd203451216;
      27138: inst = 32'd471859200;
      27139: inst = 32'd136314880;
      27140: inst = 32'd268468224;
      27141: inst = 32'd201348372;
      27142: inst = 32'd203451216;
      27143: inst = 32'd471859200;
      27144: inst = 32'd136314880;
      27145: inst = 32'd268468224;
      27146: inst = 32'd201348373;
      27147: inst = 32'd203451216;
      27148: inst = 32'd471859200;
      27149: inst = 32'd136314880;
      27150: inst = 32'd268468224;
      27151: inst = 32'd201348374;
      27152: inst = 32'd203444874;
      27153: inst = 32'd471859200;
      27154: inst = 32'd136314880;
      27155: inst = 32'd268468224;
      27156: inst = 32'd201348375;
      27157: inst = 32'd203449133;
      27158: inst = 32'd471859200;
      27159: inst = 32'd136314880;
      27160: inst = 32'd268468224;
      27161: inst = 32'd201348376;
      27162: inst = 32'd203459697;
      27163: inst = 32'd471859200;
      27164: inst = 32'd136314880;
      27165: inst = 32'd268468224;
      27166: inst = 32'd201348377;
      27167: inst = 32'd203459697;
      27168: inst = 32'd471859200;
      27169: inst = 32'd136314880;
      27170: inst = 32'd268468224;
      27171: inst = 32'd201348378;
      27172: inst = 32'd203459697;
      27173: inst = 32'd471859200;
      27174: inst = 32'd136314880;
      27175: inst = 32'd268468224;
      27176: inst = 32'd201348379;
      27177: inst = 32'd203459697;
      27178: inst = 32'd471859200;
      27179: inst = 32'd136314880;
      27180: inst = 32'd268468224;
      27181: inst = 32'd201348380;
      27182: inst = 32'd203444906;
      27183: inst = 32'd471859200;
      27184: inst = 32'd136314880;
      27185: inst = 32'd268468224;
      27186: inst = 32'd201348381;
      27187: inst = 32'd203442793;
      27188: inst = 32'd471859200;
      27189: inst = 32'd136314880;
      27190: inst = 32'd268468224;
      27191: inst = 32'd201348382;
      27192: inst = 32'd203455439;
      27193: inst = 32'd471859200;
      27194: inst = 32'd136314880;
      27195: inst = 32'd268468224;
      27196: inst = 32'd201348383;
      27197: inst = 32'd203459697;
      27198: inst = 32'd471859200;
      27199: inst = 32'd136314880;
      27200: inst = 32'd268468224;
      27201: inst = 32'd201348384;
      27202: inst = 32'd203453358;
      27203: inst = 32'd471859200;
      27204: inst = 32'd136314880;
      27205: inst = 32'd268468224;
      27206: inst = 32'd201348385;
      27207: inst = 32'd203442793;
      27208: inst = 32'd471859200;
      27209: inst = 32'd136314880;
      27210: inst = 32'd268468224;
      27211: inst = 32'd201348386;
      27212: inst = 32'd203442793;
      27213: inst = 32'd471859200;
      27214: inst = 32'd136314880;
      27215: inst = 32'd268468224;
      27216: inst = 32'd201348387;
      27217: inst = 32'd203442793;
      27218: inst = 32'd471859200;
      27219: inst = 32'd136314880;
      27220: inst = 32'd268468224;
      27221: inst = 32'd201348388;
      27222: inst = 32'd203444906;
      27223: inst = 32'd471859200;
      27224: inst = 32'd136314880;
      27225: inst = 32'd268468224;
      27226: inst = 32'd201348389;
      27227: inst = 32'd203459665;
      27228: inst = 32'd471859200;
      27229: inst = 32'd136314880;
      27230: inst = 32'd268468224;
      27231: inst = 32'd201348390;
      27232: inst = 32'd203459697;
      27233: inst = 32'd471859200;
      27234: inst = 32'd136314880;
      27235: inst = 32'd268468224;
      27236: inst = 32'd201348391;
      27237: inst = 32'd203459697;
      27238: inst = 32'd471859200;
      27239: inst = 32'd136314880;
      27240: inst = 32'd268468224;
      27241: inst = 32'd201348392;
      27242: inst = 32'd203453360;
      27243: inst = 32'd471859200;
      27244: inst = 32'd136314880;
      27245: inst = 32'd268468224;
      27246: inst = 32'd201348393;
      27247: inst = 32'd203451216;
      27248: inst = 32'd471859200;
      27249: inst = 32'd136314880;
      27250: inst = 32'd268468224;
      27251: inst = 32'd201348394;
      27252: inst = 32'd203451216;
      27253: inst = 32'd471859200;
      27254: inst = 32'd136314880;
      27255: inst = 32'd268468224;
      27256: inst = 32'd201348395;
      27257: inst = 32'd203451216;
      27258: inst = 32'd471859200;
      27259: inst = 32'd136314880;
      27260: inst = 32'd268468224;
      27261: inst = 32'd201348396;
      27262: inst = 32'd203451216;
      27263: inst = 32'd471859200;
      27264: inst = 32'd136314880;
      27265: inst = 32'd268468224;
      27266: inst = 32'd201348397;
      27267: inst = 32'd203451216;
      27268: inst = 32'd471859200;
      27269: inst = 32'd136314880;
      27270: inst = 32'd268468224;
      27271: inst = 32'd201348398;
      27272: inst = 32'd203451216;
      27273: inst = 32'd471859200;
      27274: inst = 32'd136314880;
      27275: inst = 32'd268468224;
      27276: inst = 32'd201348399;
      27277: inst = 32'd203451216;
      27278: inst = 32'd471859200;
      27279: inst = 32'd136314880;
      27280: inst = 32'd268468224;
      27281: inst = 32'd201348400;
      27282: inst = 32'd203451216;
      27283: inst = 32'd471859200;
      27284: inst = 32'd136314880;
      27285: inst = 32'd268468224;
      27286: inst = 32'd201348401;
      27287: inst = 32'd203451216;
      27288: inst = 32'd471859200;
      27289: inst = 32'd136314880;
      27290: inst = 32'd268468224;
      27291: inst = 32'd201348402;
      27292: inst = 32'd203451216;
      27293: inst = 32'd471859200;
      27294: inst = 32'd136314880;
      27295: inst = 32'd268468224;
      27296: inst = 32'd201348403;
      27297: inst = 32'd203451216;
      27298: inst = 32'd471859200;
      27299: inst = 32'd136314880;
      27300: inst = 32'd268468224;
      27301: inst = 32'd201348404;
      27302: inst = 32'd203451216;
      27303: inst = 32'd471859200;
      27304: inst = 32'd136314880;
      27305: inst = 32'd268468224;
      27306: inst = 32'd201348405;
      27307: inst = 32'd203451216;
      27308: inst = 32'd471859200;
      27309: inst = 32'd136314880;
      27310: inst = 32'd268468224;
      27311: inst = 32'd201348406;
      27312: inst = 32'd203451216;
      27313: inst = 32'd471859200;
      27314: inst = 32'd136314880;
      27315: inst = 32'd268468224;
      27316: inst = 32'd201348407;
      27317: inst = 32'd203451216;
      27318: inst = 32'd471859200;
      27319: inst = 32'd136314880;
      27320: inst = 32'd268468224;
      27321: inst = 32'd201348408;
      27322: inst = 32'd203451216;
      27323: inst = 32'd471859200;
      27324: inst = 32'd136314880;
      27325: inst = 32'd268468224;
      27326: inst = 32'd201348409;
      27327: inst = 32'd203451216;
      27328: inst = 32'd471859200;
      27329: inst = 32'd136314880;
      27330: inst = 32'd268468224;
      27331: inst = 32'd201348410;
      27332: inst = 32'd203451216;
      27333: inst = 32'd471859200;
      27334: inst = 32'd136314880;
      27335: inst = 32'd268468224;
      27336: inst = 32'd201348411;
      27337: inst = 32'd203451216;
      27338: inst = 32'd471859200;
      27339: inst = 32'd136314880;
      27340: inst = 32'd268468224;
      27341: inst = 32'd201348412;
      27342: inst = 32'd203451216;
      27343: inst = 32'd471859200;
      27344: inst = 32'd136314880;
      27345: inst = 32'd268468224;
      27346: inst = 32'd201348413;
      27347: inst = 32'd203451216;
      27348: inst = 32'd471859200;
      27349: inst = 32'd136314880;
      27350: inst = 32'd268468224;
      27351: inst = 32'd201348414;
      27352: inst = 32'd203451216;
      27353: inst = 32'd471859200;
      27354: inst = 32'd136314880;
      27355: inst = 32'd268468224;
      27356: inst = 32'd201348415;
      27357: inst = 32'd203451216;
      27358: inst = 32'd471859200;
      27359: inst = 32'd136314880;
      27360: inst = 32'd268468224;
      27361: inst = 32'd201348416;
      27362: inst = 32'd203451216;
      27363: inst = 32'd471859200;
      27364: inst = 32'd136314880;
      27365: inst = 32'd268468224;
      27366: inst = 32'd201348417;
      27367: inst = 32'd203451216;
      27368: inst = 32'd471859200;
      27369: inst = 32'd136314880;
      27370: inst = 32'd268468224;
      27371: inst = 32'd201348418;
      27372: inst = 32'd203451216;
      27373: inst = 32'd471859200;
      27374: inst = 32'd136314880;
      27375: inst = 32'd268468224;
      27376: inst = 32'd201348419;
      27377: inst = 32'd203451216;
      27378: inst = 32'd471859200;
      27379: inst = 32'd136314880;
      27380: inst = 32'd268468224;
      27381: inst = 32'd201348420;
      27382: inst = 32'd203451216;
      27383: inst = 32'd471859200;
      27384: inst = 32'd136314880;
      27385: inst = 32'd268468224;
      27386: inst = 32'd201348421;
      27387: inst = 32'd203451216;
      27388: inst = 32'd471859200;
      27389: inst = 32'd136314880;
      27390: inst = 32'd268468224;
      27391: inst = 32'd201348422;
      27392: inst = 32'd203451216;
      27393: inst = 32'd471859200;
      27394: inst = 32'd136314880;
      27395: inst = 32'd268468224;
      27396: inst = 32'd201348423;
      27397: inst = 32'd203451216;
      27398: inst = 32'd471859200;
      27399: inst = 32'd136314880;
      27400: inst = 32'd268468224;
      27401: inst = 32'd201348424;
      27402: inst = 32'd203451216;
      27403: inst = 32'd471859200;
      27404: inst = 32'd136314880;
      27405: inst = 32'd268468224;
      27406: inst = 32'd201348425;
      27407: inst = 32'd203451216;
      27408: inst = 32'd471859200;
      27409: inst = 32'd136314880;
      27410: inst = 32'd268468224;
      27411: inst = 32'd201348426;
      27412: inst = 32'd203451216;
      27413: inst = 32'd471859200;
      27414: inst = 32'd136314880;
      27415: inst = 32'd268468224;
      27416: inst = 32'd201348427;
      27417: inst = 32'd203451216;
      27418: inst = 32'd471859200;
      27419: inst = 32'd136314880;
      27420: inst = 32'd268468224;
      27421: inst = 32'd201348428;
      27422: inst = 32'd203451216;
      27423: inst = 32'd471859200;
      27424: inst = 32'd136314880;
      27425: inst = 32'd268468224;
      27426: inst = 32'd201348429;
      27427: inst = 32'd203451216;
      27428: inst = 32'd471859200;
      27429: inst = 32'd136314880;
      27430: inst = 32'd268468224;
      27431: inst = 32'd201348430;
      27432: inst = 32'd203451216;
      27433: inst = 32'd471859200;
      27434: inst = 32'd136314880;
      27435: inst = 32'd268468224;
      27436: inst = 32'd201348431;
      27437: inst = 32'd203451216;
      27438: inst = 32'd471859200;
      27439: inst = 32'd136314880;
      27440: inst = 32'd268468224;
      27441: inst = 32'd201348432;
      27442: inst = 32'd203451216;
      27443: inst = 32'd471859200;
      27444: inst = 32'd136314880;
      27445: inst = 32'd268468224;
      27446: inst = 32'd201348433;
      27447: inst = 32'd203451216;
      27448: inst = 32'd471859200;
      27449: inst = 32'd136314880;
      27450: inst = 32'd268468224;
      27451: inst = 32'd201348434;
      27452: inst = 32'd203451216;
      27453: inst = 32'd471859200;
      27454: inst = 32'd136314880;
      27455: inst = 32'd268468224;
      27456: inst = 32'd201348435;
      27457: inst = 32'd203451216;
      27458: inst = 32'd471859200;
      27459: inst = 32'd136314880;
      27460: inst = 32'd268468224;
      27461: inst = 32'd201348436;
      27462: inst = 32'd203451216;
      27463: inst = 32'd471859200;
      27464: inst = 32'd136314880;
      27465: inst = 32'd268468224;
      27466: inst = 32'd201348437;
      27467: inst = 32'd203451216;
      27468: inst = 32'd471859200;
      27469: inst = 32'd136314880;
      27470: inst = 32'd268468224;
      27471: inst = 32'd201348438;
      27472: inst = 32'd203451248;
      27473: inst = 32'd471859200;
      27474: inst = 32'd136314880;
      27475: inst = 32'd268468224;
      27476: inst = 32'd201348439;
      27477: inst = 32'd203459665;
      27478: inst = 32'd471859200;
      27479: inst = 32'd136314880;
      27480: inst = 32'd268468224;
      27481: inst = 32'd201348440;
      27482: inst = 32'd203459697;
      27483: inst = 32'd471859200;
      27484: inst = 32'd136314880;
      27485: inst = 32'd268468224;
      27486: inst = 32'd201348441;
      27487: inst = 32'd203459697;
      27488: inst = 32'd471859200;
      27489: inst = 32'd136314880;
      27490: inst = 32'd268468224;
      27491: inst = 32'd201348442;
      27492: inst = 32'd203451181;
      27493: inst = 32'd471859200;
      27494: inst = 32'd136314880;
      27495: inst = 32'd268468224;
      27496: inst = 32'd201348443;
      27497: inst = 32'd203442793;
      27498: inst = 32'd471859200;
      27499: inst = 32'd136314880;
      27500: inst = 32'd268468224;
      27501: inst = 32'd201348444;
      27502: inst = 32'd203442793;
      27503: inst = 32'd471859200;
      27504: inst = 32'd136314880;
      27505: inst = 32'd268468224;
      27506: inst = 32'd201348445;
      27507: inst = 32'd203442793;
      27508: inst = 32'd471859200;
      27509: inst = 32'd136314880;
      27510: inst = 32'd268468224;
      27511: inst = 32'd201348446;
      27512: inst = 32'd203444874;
      27513: inst = 32'd471859200;
      27514: inst = 32'd136314880;
      27515: inst = 32'd268468224;
      27516: inst = 32'd201348447;
      27517: inst = 32'd203459665;
      27518: inst = 32'd471859200;
      27519: inst = 32'd136314880;
      27520: inst = 32'd268468224;
      27521: inst = 32'd201348448;
      27522: inst = 32'd203459697;
      27523: inst = 32'd471859200;
      27524: inst = 32'd136314880;
      27525: inst = 32'd268468224;
      27526: inst = 32'd201348449;
      27527: inst = 32'd203455439;
      27528: inst = 32'd471859200;
      27529: inst = 32'd136314880;
      27530: inst = 32'd268468224;
      27531: inst = 32'd201348450;
      27532: inst = 32'd203442793;
      27533: inst = 32'd471859200;
      27534: inst = 32'd136314880;
      27535: inst = 32'd268468224;
      27536: inst = 32'd201348451;
      27537: inst = 32'd203451213;
      27538: inst = 32'd471859200;
      27539: inst = 32'd136314880;
      27540: inst = 32'd268468224;
      27541: inst = 32'd201348452;
      27542: inst = 32'd203459697;
      27543: inst = 32'd471859200;
      27544: inst = 32'd136314880;
      27545: inst = 32'd268468224;
      27546: inst = 32'd201348453;
      27547: inst = 32'd203459697;
      27548: inst = 32'd471859200;
      27549: inst = 32'd136314880;
      27550: inst = 32'd268468224;
      27551: inst = 32'd201348454;
      27552: inst = 32'd203459697;
      27553: inst = 32'd471859200;
      27554: inst = 32'd136314880;
      27555: inst = 32'd268468224;
      27556: inst = 32'd201348455;
      27557: inst = 32'd203459697;
      27558: inst = 32'd471859200;
      27559: inst = 32'd136314880;
      27560: inst = 32'd268468224;
      27561: inst = 32'd201348456;
      27562: inst = 32'd203447020;
      27563: inst = 32'd471859200;
      27564: inst = 32'd136314880;
      27565: inst = 32'd268468224;
      27566: inst = 32'd201348457;
      27567: inst = 32'd203444874;
      27568: inst = 32'd471859200;
      27569: inst = 32'd136314880;
      27570: inst = 32'd268468224;
      27571: inst = 32'd201348458;
      27572: inst = 32'd203451216;
      27573: inst = 32'd471859200;
      27574: inst = 32'd136314880;
      27575: inst = 32'd268468224;
      27576: inst = 32'd201348459;
      27577: inst = 32'd203451216;
      27578: inst = 32'd471859200;
      27579: inst = 32'd136314880;
      27580: inst = 32'd268468224;
      27581: inst = 32'd201348460;
      27582: inst = 32'd203451216;
      27583: inst = 32'd471859200;
      27584: inst = 32'd136314880;
      27585: inst = 32'd268468224;
      27586: inst = 32'd201348461;
      27587: inst = 32'd203451216;
      27588: inst = 32'd471859200;
      27589: inst = 32'd136314880;
      27590: inst = 32'd268468224;
      27591: inst = 32'd201348462;
      27592: inst = 32'd203451216;
      27593: inst = 32'd471859200;
      27594: inst = 32'd136314880;
      27595: inst = 32'd268468224;
      27596: inst = 32'd201348463;
      27597: inst = 32'd203451216;
      27598: inst = 32'd471859200;
      27599: inst = 32'd136314880;
      27600: inst = 32'd268468224;
      27601: inst = 32'd201348464;
      27602: inst = 32'd203451216;
      27603: inst = 32'd471859200;
      27604: inst = 32'd136314880;
      27605: inst = 32'd268468224;
      27606: inst = 32'd201348465;
      27607: inst = 32'd203451216;
      27608: inst = 32'd471859200;
      27609: inst = 32'd136314880;
      27610: inst = 32'd268468224;
      27611: inst = 32'd201348466;
      27612: inst = 32'd203451216;
      27613: inst = 32'd471859200;
      27614: inst = 32'd136314880;
      27615: inst = 32'd268468224;
      27616: inst = 32'd201348467;
      27617: inst = 32'd203451216;
      27618: inst = 32'd471859200;
      27619: inst = 32'd136314880;
      27620: inst = 32'd268468224;
      27621: inst = 32'd201348468;
      27622: inst = 32'd203451216;
      27623: inst = 32'd471859200;
      27624: inst = 32'd136314880;
      27625: inst = 32'd268468224;
      27626: inst = 32'd201348469;
      27627: inst = 32'd203451216;
      27628: inst = 32'd471859200;
      27629: inst = 32'd136314880;
      27630: inst = 32'd268468224;
      27631: inst = 32'd201348470;
      27632: inst = 32'd203444874;
      27633: inst = 32'd471859200;
      27634: inst = 32'd136314880;
      27635: inst = 32'd268468224;
      27636: inst = 32'd201348471;
      27637: inst = 32'd203447020;
      27638: inst = 32'd471859200;
      27639: inst = 32'd136314880;
      27640: inst = 32'd268468224;
      27641: inst = 32'd201348472;
      27642: inst = 32'd203459697;
      27643: inst = 32'd471859200;
      27644: inst = 32'd136314880;
      27645: inst = 32'd268468224;
      27646: inst = 32'd201348473;
      27647: inst = 32'd203459697;
      27648: inst = 32'd471859200;
      27649: inst = 32'd136314880;
      27650: inst = 32'd268468224;
      27651: inst = 32'd201348474;
      27652: inst = 32'd203459697;
      27653: inst = 32'd471859200;
      27654: inst = 32'd136314880;
      27655: inst = 32'd268468224;
      27656: inst = 32'd201348475;
      27657: inst = 32'd203459697;
      27658: inst = 32'd471859200;
      27659: inst = 32'd136314880;
      27660: inst = 32'd268468224;
      27661: inst = 32'd201348476;
      27662: inst = 32'd203451213;
      27663: inst = 32'd471859200;
      27664: inst = 32'd136314880;
      27665: inst = 32'd268468224;
      27666: inst = 32'd201348477;
      27667: inst = 32'd203442793;
      27668: inst = 32'd471859200;
      27669: inst = 32'd136314880;
      27670: inst = 32'd268468224;
      27671: inst = 32'd201348478;
      27672: inst = 32'd203455439;
      27673: inst = 32'd471859200;
      27674: inst = 32'd136314880;
      27675: inst = 32'd268468224;
      27676: inst = 32'd201348479;
      27677: inst = 32'd203459697;
      27678: inst = 32'd471859200;
      27679: inst = 32'd136314880;
      27680: inst = 32'd268468224;
      27681: inst = 32'd201348480;
      27682: inst = 32'd203459665;
      27683: inst = 32'd471859200;
      27684: inst = 32'd136314880;
      27685: inst = 32'd268468224;
      27686: inst = 32'd201348481;
      27687: inst = 32'd203444874;
      27688: inst = 32'd471859200;
      27689: inst = 32'd136314880;
      27690: inst = 32'd268468224;
      27691: inst = 32'd201348482;
      27692: inst = 32'd203442793;
      27693: inst = 32'd471859200;
      27694: inst = 32'd136314880;
      27695: inst = 32'd268468224;
      27696: inst = 32'd201348483;
      27697: inst = 32'd203442793;
      27698: inst = 32'd471859200;
      27699: inst = 32'd136314880;
      27700: inst = 32'd268468224;
      27701: inst = 32'd201348484;
      27702: inst = 32'd203442793;
      27703: inst = 32'd471859200;
      27704: inst = 32'd136314880;
      27705: inst = 32'd268468224;
      27706: inst = 32'd201348485;
      27707: inst = 32'd203451181;
      27708: inst = 32'd471859200;
      27709: inst = 32'd136314880;
      27710: inst = 32'd268468224;
      27711: inst = 32'd201348486;
      27712: inst = 32'd203459697;
      27713: inst = 32'd471859200;
      27714: inst = 32'd136314880;
      27715: inst = 32'd268468224;
      27716: inst = 32'd201348487;
      27717: inst = 32'd203459697;
      27718: inst = 32'd471859200;
      27719: inst = 32'd136314880;
      27720: inst = 32'd268468224;
      27721: inst = 32'd201348488;
      27722: inst = 32'd203459665;
      27723: inst = 32'd471859200;
      27724: inst = 32'd136314880;
      27725: inst = 32'd268468224;
      27726: inst = 32'd201348489;
      27727: inst = 32'd203451248;
      27728: inst = 32'd471859200;
      27729: inst = 32'd136314880;
      27730: inst = 32'd268468224;
      27731: inst = 32'd201348490;
      27732: inst = 32'd203451216;
      27733: inst = 32'd471859200;
      27734: inst = 32'd136314880;
      27735: inst = 32'd268468224;
      27736: inst = 32'd201348491;
      27737: inst = 32'd203451216;
      27738: inst = 32'd471859200;
      27739: inst = 32'd136314880;
      27740: inst = 32'd268468224;
      27741: inst = 32'd201348492;
      27742: inst = 32'd203451216;
      27743: inst = 32'd471859200;
      27744: inst = 32'd136314880;
      27745: inst = 32'd268468224;
      27746: inst = 32'd201348493;
      27747: inst = 32'd203451216;
      27748: inst = 32'd471859200;
      27749: inst = 32'd136314880;
      27750: inst = 32'd268468224;
      27751: inst = 32'd201348494;
      27752: inst = 32'd203451216;
      27753: inst = 32'd471859200;
      27754: inst = 32'd136314880;
      27755: inst = 32'd268468224;
      27756: inst = 32'd201348495;
      27757: inst = 32'd203451216;
      27758: inst = 32'd471859200;
      27759: inst = 32'd136314880;
      27760: inst = 32'd268468224;
      27761: inst = 32'd201348496;
      27762: inst = 32'd203451216;
      27763: inst = 32'd471859200;
      27764: inst = 32'd136314880;
      27765: inst = 32'd268468224;
      27766: inst = 32'd201348497;
      27767: inst = 32'd203451216;
      27768: inst = 32'd471859200;
      27769: inst = 32'd136314880;
      27770: inst = 32'd268468224;
      27771: inst = 32'd201348498;
      27772: inst = 32'd203451216;
      27773: inst = 32'd471859200;
      27774: inst = 32'd136314880;
      27775: inst = 32'd268468224;
      27776: inst = 32'd201348499;
      27777: inst = 32'd203451216;
      27778: inst = 32'd471859200;
      27779: inst = 32'd136314880;
      27780: inst = 32'd268468224;
      27781: inst = 32'd201348500;
      27782: inst = 32'd203451216;
      27783: inst = 32'd471859200;
      27784: inst = 32'd136314880;
      27785: inst = 32'd268468224;
      27786: inst = 32'd201348501;
      27787: inst = 32'd203451216;
      27788: inst = 32'd471859200;
      27789: inst = 32'd136314880;
      27790: inst = 32'd268468224;
      27791: inst = 32'd201348502;
      27792: inst = 32'd203451216;
      27793: inst = 32'd471859200;
      27794: inst = 32'd136314880;
      27795: inst = 32'd268468224;
      27796: inst = 32'd201348503;
      27797: inst = 32'd203451216;
      27798: inst = 32'd471859200;
      27799: inst = 32'd136314880;
      27800: inst = 32'd268468224;
      27801: inst = 32'd201348504;
      27802: inst = 32'd203451216;
      27803: inst = 32'd471859200;
      27804: inst = 32'd136314880;
      27805: inst = 32'd268468224;
      27806: inst = 32'd201348505;
      27807: inst = 32'd203451216;
      27808: inst = 32'd471859200;
      27809: inst = 32'd136314880;
      27810: inst = 32'd268468224;
      27811: inst = 32'd201348506;
      27812: inst = 32'd203451216;
      27813: inst = 32'd471859200;
      27814: inst = 32'd136314880;
      27815: inst = 32'd268468224;
      27816: inst = 32'd201348507;
      27817: inst = 32'd203451216;
      27818: inst = 32'd471859200;
      27819: inst = 32'd136314880;
      27820: inst = 32'd268468224;
      27821: inst = 32'd201348508;
      27822: inst = 32'd203451216;
      27823: inst = 32'd471859200;
      27824: inst = 32'd136314880;
      27825: inst = 32'd268468224;
      27826: inst = 32'd201348509;
      27827: inst = 32'd203451216;
      27828: inst = 32'd471859200;
      27829: inst = 32'd136314880;
      27830: inst = 32'd268468224;
      27831: inst = 32'd201348510;
      27832: inst = 32'd203451216;
      27833: inst = 32'd471859200;
      27834: inst = 32'd136314880;
      27835: inst = 32'd268468224;
      27836: inst = 32'd201348511;
      27837: inst = 32'd203451216;
      27838: inst = 32'd471859200;
      27839: inst = 32'd136314880;
      27840: inst = 32'd268468224;
      27841: inst = 32'd201348512;
      27842: inst = 32'd203451216;
      27843: inst = 32'd471859200;
      27844: inst = 32'd136314880;
      27845: inst = 32'd268468224;
      27846: inst = 32'd201348513;
      27847: inst = 32'd203451216;
      27848: inst = 32'd471859200;
      27849: inst = 32'd136314880;
      27850: inst = 32'd268468224;
      27851: inst = 32'd201348514;
      27852: inst = 32'd203451216;
      27853: inst = 32'd471859200;
      27854: inst = 32'd136314880;
      27855: inst = 32'd268468224;
      27856: inst = 32'd201348515;
      27857: inst = 32'd203451216;
      27858: inst = 32'd471859200;
      27859: inst = 32'd136314880;
      27860: inst = 32'd268468224;
      27861: inst = 32'd201348516;
      27862: inst = 32'd203451216;
      27863: inst = 32'd471859200;
      27864: inst = 32'd136314880;
      27865: inst = 32'd268468224;
      27866: inst = 32'd201348517;
      27867: inst = 32'd203451216;
      27868: inst = 32'd471859200;
      27869: inst = 32'd136314880;
      27870: inst = 32'd268468224;
      27871: inst = 32'd201348518;
      27872: inst = 32'd203451216;
      27873: inst = 32'd471859200;
      27874: inst = 32'd136314880;
      27875: inst = 32'd268468224;
      27876: inst = 32'd201348519;
      27877: inst = 32'd203451216;
      27878: inst = 32'd471859200;
      27879: inst = 32'd136314880;
      27880: inst = 32'd268468224;
      27881: inst = 32'd201348520;
      27882: inst = 32'd203451216;
      27883: inst = 32'd471859200;
      27884: inst = 32'd136314880;
      27885: inst = 32'd268468224;
      27886: inst = 32'd201348521;
      27887: inst = 32'd203451216;
      27888: inst = 32'd471859200;
      27889: inst = 32'd136314880;
      27890: inst = 32'd268468224;
      27891: inst = 32'd201348522;
      27892: inst = 32'd203451216;
      27893: inst = 32'd471859200;
      27894: inst = 32'd136314880;
      27895: inst = 32'd268468224;
      27896: inst = 32'd201348523;
      27897: inst = 32'd203451216;
      27898: inst = 32'd471859200;
      27899: inst = 32'd136314880;
      27900: inst = 32'd268468224;
      27901: inst = 32'd201348524;
      27902: inst = 32'd203451216;
      27903: inst = 32'd471859200;
      27904: inst = 32'd136314880;
      27905: inst = 32'd268468224;
      27906: inst = 32'd201348525;
      27907: inst = 32'd203451216;
      27908: inst = 32'd471859200;
      27909: inst = 32'd136314880;
      27910: inst = 32'd268468224;
      27911: inst = 32'd201348526;
      27912: inst = 32'd203451216;
      27913: inst = 32'd471859200;
      27914: inst = 32'd136314880;
      27915: inst = 32'd268468224;
      27916: inst = 32'd201348527;
      27917: inst = 32'd203451216;
      27918: inst = 32'd471859200;
      27919: inst = 32'd136314880;
      27920: inst = 32'd268468224;
      27921: inst = 32'd201348528;
      27922: inst = 32'd203451216;
      27923: inst = 32'd471859200;
      27924: inst = 32'd136314880;
      27925: inst = 32'd268468224;
      27926: inst = 32'd201348529;
      27927: inst = 32'd203451216;
      27928: inst = 32'd471859200;
      27929: inst = 32'd136314880;
      27930: inst = 32'd268468224;
      27931: inst = 32'd201348530;
      27932: inst = 32'd203451216;
      27933: inst = 32'd471859200;
      27934: inst = 32'd136314880;
      27935: inst = 32'd268468224;
      27936: inst = 32'd201348531;
      27937: inst = 32'd203451216;
      27938: inst = 32'd471859200;
      27939: inst = 32'd136314880;
      27940: inst = 32'd268468224;
      27941: inst = 32'd201348532;
      27942: inst = 32'd203451216;
      27943: inst = 32'd471859200;
      27944: inst = 32'd136314880;
      27945: inst = 32'd268468224;
      27946: inst = 32'd201348533;
      27947: inst = 32'd203451248;
      27948: inst = 32'd471859200;
      27949: inst = 32'd136314880;
      27950: inst = 32'd268468224;
      27951: inst = 32'd201348534;
      27952: inst = 32'd203457585;
      27953: inst = 32'd471859200;
      27954: inst = 32'd136314880;
      27955: inst = 32'd268468224;
      27956: inst = 32'd201348535;
      27957: inst = 32'd203459697;
      27958: inst = 32'd471859200;
      27959: inst = 32'd136314880;
      27960: inst = 32'd268468224;
      27961: inst = 32'd201348536;
      27962: inst = 32'd203459697;
      27963: inst = 32'd471859200;
      27964: inst = 32'd136314880;
      27965: inst = 32'd268468224;
      27966: inst = 32'd201348537;
      27967: inst = 32'd203455439;
      27968: inst = 32'd471859200;
      27969: inst = 32'd136314880;
      27970: inst = 32'd268468224;
      27971: inst = 32'd201348538;
      27972: inst = 32'd203442793;
      27973: inst = 32'd471859200;
      27974: inst = 32'd136314880;
      27975: inst = 32'd268468224;
      27976: inst = 32'd201348539;
      27977: inst = 32'd203442793;
      27978: inst = 32'd471859200;
      27979: inst = 32'd136314880;
      27980: inst = 32'd268468224;
      27981: inst = 32'd201348540;
      27982: inst = 32'd203442793;
      27983: inst = 32'd471859200;
      27984: inst = 32'd136314880;
      27985: inst = 32'd268468224;
      27986: inst = 32'd201348541;
      27987: inst = 32'd203442793;
      27988: inst = 32'd471859200;
      27989: inst = 32'd136314880;
      27990: inst = 32'd268468224;
      27991: inst = 32'd201348542;
      27992: inst = 32'd203449100;
      27993: inst = 32'd471859200;
      27994: inst = 32'd136314880;
      27995: inst = 32'd268468224;
      27996: inst = 32'd201348543;
      27997: inst = 32'd203459697;
      27998: inst = 32'd471859200;
      27999: inst = 32'd136314880;
      28000: inst = 32'd268468224;
      28001: inst = 32'd201348544;
      28002: inst = 32'd203459697;
      28003: inst = 32'd471859200;
      28004: inst = 32'd136314880;
      28005: inst = 32'd268468224;
      28006: inst = 32'd201348545;
      28007: inst = 32'd203455439;
      28008: inst = 32'd471859200;
      28009: inst = 32'd136314880;
      28010: inst = 32'd268468224;
      28011: inst = 32'd201348546;
      28012: inst = 32'd203442793;
      28013: inst = 32'd471859200;
      28014: inst = 32'd136314880;
      28015: inst = 32'd268468224;
      28016: inst = 32'd201348547;
      28017: inst = 32'd203455472;
      28018: inst = 32'd471859200;
      28019: inst = 32'd136314880;
      28020: inst = 32'd268468224;
      28021: inst = 32'd201348548;
      28022: inst = 32'd203459697;
      28023: inst = 32'd471859200;
      28024: inst = 32'd136314880;
      28025: inst = 32'd268468224;
      28026: inst = 32'd201348549;
      28027: inst = 32'd203459697;
      28028: inst = 32'd471859200;
      28029: inst = 32'd136314880;
      28030: inst = 32'd268468224;
      28031: inst = 32'd201348550;
      28032: inst = 32'd203459697;
      28033: inst = 32'd471859200;
      28034: inst = 32'd136314880;
      28035: inst = 32'd268468224;
      28036: inst = 32'd201348551;
      28037: inst = 32'd203459697;
      28038: inst = 32'd471859200;
      28039: inst = 32'd136314880;
      28040: inst = 32'd268468224;
      28041: inst = 32'd201348552;
      28042: inst = 32'd203444906;
      28043: inst = 32'd471859200;
      28044: inst = 32'd136314880;
      28045: inst = 32'd268468224;
      28046: inst = 32'd201348553;
      28047: inst = 32'd203444874;
      28048: inst = 32'd471859200;
      28049: inst = 32'd136314880;
      28050: inst = 32'd268468224;
      28051: inst = 32'd201348554;
      28052: inst = 32'd203451216;
      28053: inst = 32'd471859200;
      28054: inst = 32'd136314880;
      28055: inst = 32'd268468224;
      28056: inst = 32'd201348555;
      28057: inst = 32'd203451216;
      28058: inst = 32'd471859200;
      28059: inst = 32'd136314880;
      28060: inst = 32'd268468224;
      28061: inst = 32'd201348556;
      28062: inst = 32'd203451216;
      28063: inst = 32'd471859200;
      28064: inst = 32'd136314880;
      28065: inst = 32'd268468224;
      28066: inst = 32'd201348557;
      28067: inst = 32'd203451216;
      28068: inst = 32'd471859200;
      28069: inst = 32'd136314880;
      28070: inst = 32'd268468224;
      28071: inst = 32'd201348558;
      28072: inst = 32'd203451216;
      28073: inst = 32'd471859200;
      28074: inst = 32'd136314880;
      28075: inst = 32'd268468224;
      28076: inst = 32'd201348559;
      28077: inst = 32'd203451216;
      28078: inst = 32'd471859200;
      28079: inst = 32'd136314880;
      28080: inst = 32'd268468224;
      28081: inst = 32'd201348560;
      28082: inst = 32'd203451216;
      28083: inst = 32'd471859200;
      28084: inst = 32'd136314880;
      28085: inst = 32'd268468224;
      28086: inst = 32'd201348561;
      28087: inst = 32'd203451216;
      28088: inst = 32'd471859200;
      28089: inst = 32'd136314880;
      28090: inst = 32'd268468224;
      28091: inst = 32'd201348562;
      28092: inst = 32'd203451216;
      28093: inst = 32'd471859200;
      28094: inst = 32'd136314880;
      28095: inst = 32'd268468224;
      28096: inst = 32'd201348563;
      28097: inst = 32'd203451216;
      28098: inst = 32'd471859200;
      28099: inst = 32'd136314880;
      28100: inst = 32'd268468224;
      28101: inst = 32'd201348564;
      28102: inst = 32'd203451216;
      28103: inst = 32'd471859200;
      28104: inst = 32'd136314880;
      28105: inst = 32'd268468224;
      28106: inst = 32'd201348565;
      28107: inst = 32'd203451216;
      28108: inst = 32'd471859200;
      28109: inst = 32'd136314880;
      28110: inst = 32'd268468224;
      28111: inst = 32'd201348566;
      28112: inst = 32'd203444874;
      28113: inst = 32'd471859200;
      28114: inst = 32'd136314880;
      28115: inst = 32'd268468224;
      28116: inst = 32'd201348567;
      28117: inst = 32'd203444906;
      28118: inst = 32'd471859200;
      28119: inst = 32'd136314880;
      28120: inst = 32'd268468224;
      28121: inst = 32'd201348568;
      28122: inst = 32'd203459697;
      28123: inst = 32'd471859200;
      28124: inst = 32'd136314880;
      28125: inst = 32'd268468224;
      28126: inst = 32'd201348569;
      28127: inst = 32'd203459697;
      28128: inst = 32'd471859200;
      28129: inst = 32'd136314880;
      28130: inst = 32'd268468224;
      28131: inst = 32'd201348570;
      28132: inst = 32'd203459697;
      28133: inst = 32'd471859200;
      28134: inst = 32'd136314880;
      28135: inst = 32'd268468224;
      28136: inst = 32'd201348571;
      28137: inst = 32'd203459697;
      28138: inst = 32'd471859200;
      28139: inst = 32'd136314880;
      28140: inst = 32'd268468224;
      28141: inst = 32'd201348572;
      28142: inst = 32'd203455472;
      28143: inst = 32'd471859200;
      28144: inst = 32'd136314880;
      28145: inst = 32'd268468224;
      28146: inst = 32'd201348573;
      28147: inst = 32'd203442793;
      28148: inst = 32'd471859200;
      28149: inst = 32'd136314880;
      28150: inst = 32'd268468224;
      28151: inst = 32'd201348574;
      28152: inst = 32'd203455439;
      28153: inst = 32'd471859200;
      28154: inst = 32'd136314880;
      28155: inst = 32'd268468224;
      28156: inst = 32'd201348575;
      28157: inst = 32'd203459697;
      28158: inst = 32'd471859200;
      28159: inst = 32'd136314880;
      28160: inst = 32'd268468224;
      28161: inst = 32'd201348576;
      28162: inst = 32'd203459697;
      28163: inst = 32'd471859200;
      28164: inst = 32'd136314880;
      28165: inst = 32'd268468224;
      28166: inst = 32'd201348577;
      28167: inst = 32'd203449100;
      28168: inst = 32'd471859200;
      28169: inst = 32'd136314880;
      28170: inst = 32'd268468224;
      28171: inst = 32'd201348578;
      28172: inst = 32'd203442793;
      28173: inst = 32'd471859200;
      28174: inst = 32'd136314880;
      28175: inst = 32'd268468224;
      28176: inst = 32'd201348579;
      28177: inst = 32'd203442793;
      28178: inst = 32'd471859200;
      28179: inst = 32'd136314880;
      28180: inst = 32'd268468224;
      28181: inst = 32'd201348580;
      28182: inst = 32'd203442793;
      28183: inst = 32'd471859200;
      28184: inst = 32'd136314880;
      28185: inst = 32'd268468224;
      28186: inst = 32'd201348581;
      28187: inst = 32'd203442793;
      28188: inst = 32'd471859200;
      28189: inst = 32'd136314880;
      28190: inst = 32'd268468224;
      28191: inst = 32'd201348582;
      28192: inst = 32'd203455439;
      28193: inst = 32'd471859200;
      28194: inst = 32'd136314880;
      28195: inst = 32'd268468224;
      28196: inst = 32'd201348583;
      28197: inst = 32'd203459697;
      28198: inst = 32'd471859200;
      28199: inst = 32'd136314880;
      28200: inst = 32'd268468224;
      28201: inst = 32'd201348584;
      28202: inst = 32'd203459697;
      28203: inst = 32'd471859200;
      28204: inst = 32'd136314880;
      28205: inst = 32'd268468224;
      28206: inst = 32'd201348585;
      28207: inst = 32'd203457585;
      28208: inst = 32'd471859200;
      28209: inst = 32'd136314880;
      28210: inst = 32'd268468224;
      28211: inst = 32'd201348586;
      28212: inst = 32'd203451248;
      28213: inst = 32'd471859200;
      28214: inst = 32'd136314880;
      28215: inst = 32'd268468224;
      28216: inst = 32'd201348587;
      28217: inst = 32'd203451216;
      28218: inst = 32'd471859200;
      28219: inst = 32'd136314880;
      28220: inst = 32'd268468224;
      28221: inst = 32'd201348588;
      28222: inst = 32'd203451216;
      28223: inst = 32'd471859200;
      28224: inst = 32'd136314880;
      28225: inst = 32'd268468224;
      28226: inst = 32'd201348589;
      28227: inst = 32'd203451216;
      28228: inst = 32'd471859200;
      28229: inst = 32'd136314880;
      28230: inst = 32'd268468224;
      28231: inst = 32'd201348590;
      28232: inst = 32'd203451216;
      28233: inst = 32'd471859200;
      28234: inst = 32'd136314880;
      28235: inst = 32'd268468224;
      28236: inst = 32'd201348591;
      28237: inst = 32'd203451216;
      28238: inst = 32'd471859200;
      28239: inst = 32'd136314880;
      28240: inst = 32'd268468224;
      28241: inst = 32'd201348592;
      28242: inst = 32'd203451216;
      28243: inst = 32'd471859200;
      28244: inst = 32'd136314880;
      28245: inst = 32'd268468224;
      28246: inst = 32'd201348593;
      28247: inst = 32'd203451216;
      28248: inst = 32'd471859200;
      28249: inst = 32'd136314880;
      28250: inst = 32'd268468224;
      28251: inst = 32'd201348594;
      28252: inst = 32'd203451216;
      28253: inst = 32'd471859200;
      28254: inst = 32'd136314880;
      28255: inst = 32'd268468224;
      28256: inst = 32'd201348595;
      28257: inst = 32'd203451216;
      28258: inst = 32'd471859200;
      28259: inst = 32'd136314880;
      28260: inst = 32'd268468224;
      28261: inst = 32'd201348596;
      28262: inst = 32'd203451216;
      28263: inst = 32'd471859200;
      28264: inst = 32'd136314880;
      28265: inst = 32'd268468224;
      28266: inst = 32'd201348597;
      28267: inst = 32'd203451216;
      28268: inst = 32'd471859200;
      28269: inst = 32'd136314880;
      28270: inst = 32'd268468224;
      28271: inst = 32'd201348598;
      28272: inst = 32'd203451216;
      28273: inst = 32'd471859200;
      28274: inst = 32'd136314880;
      28275: inst = 32'd268468224;
      28276: inst = 32'd201348599;
      28277: inst = 32'd203451216;
      28278: inst = 32'd471859200;
      28279: inst = 32'd136314880;
      28280: inst = 32'd268468224;
      28281: inst = 32'd201348600;
      28282: inst = 32'd203451216;
      28283: inst = 32'd471859200;
      28284: inst = 32'd136314880;
      28285: inst = 32'd268468224;
      28286: inst = 32'd201348601;
      28287: inst = 32'd203451216;
      28288: inst = 32'd471859200;
      28289: inst = 32'd136314880;
      28290: inst = 32'd268468224;
      28291: inst = 32'd201348602;
      28292: inst = 32'd203451216;
      28293: inst = 32'd471859200;
      28294: inst = 32'd136314880;
      28295: inst = 32'd268468224;
      28296: inst = 32'd201348603;
      28297: inst = 32'd203451216;
      28298: inst = 32'd471859200;
      28299: inst = 32'd136314880;
      28300: inst = 32'd268468224;
      28301: inst = 32'd201348604;
      28302: inst = 32'd203451216;
      28303: inst = 32'd471859200;
      28304: inst = 32'd136314880;
      28305: inst = 32'd268468224;
      28306: inst = 32'd201348605;
      28307: inst = 32'd203451216;
      28308: inst = 32'd471859200;
      28309: inst = 32'd136314880;
      28310: inst = 32'd268468224;
      28311: inst = 32'd201348606;
      28312: inst = 32'd203451216;
      28313: inst = 32'd471859200;
      28314: inst = 32'd136314880;
      28315: inst = 32'd268468224;
      28316: inst = 32'd201348607;
      28317: inst = 32'd203451216;
      28318: inst = 32'd471859200;
      28319: inst = 32'd136314880;
      28320: inst = 32'd268468224;
      28321: inst = 32'd201348608;
      28322: inst = 32'd203451216;
      28323: inst = 32'd471859200;
      28324: inst = 32'd136314880;
      28325: inst = 32'd268468224;
      28326: inst = 32'd201348609;
      28327: inst = 32'd203451216;
      28328: inst = 32'd471859200;
      28329: inst = 32'd136314880;
      28330: inst = 32'd268468224;
      28331: inst = 32'd201348610;
      28332: inst = 32'd203451216;
      28333: inst = 32'd471859200;
      28334: inst = 32'd136314880;
      28335: inst = 32'd268468224;
      28336: inst = 32'd201348611;
      28337: inst = 32'd203451216;
      28338: inst = 32'd471859200;
      28339: inst = 32'd136314880;
      28340: inst = 32'd268468224;
      28341: inst = 32'd201348612;
      28342: inst = 32'd203451216;
      28343: inst = 32'd471859200;
      28344: inst = 32'd136314880;
      28345: inst = 32'd268468224;
      28346: inst = 32'd201348613;
      28347: inst = 32'd203451216;
      28348: inst = 32'd471859200;
      28349: inst = 32'd136314880;
      28350: inst = 32'd268468224;
      28351: inst = 32'd201348614;
      28352: inst = 32'd203451216;
      28353: inst = 32'd471859200;
      28354: inst = 32'd136314880;
      28355: inst = 32'd268468224;
      28356: inst = 32'd201348615;
      28357: inst = 32'd203451216;
      28358: inst = 32'd471859200;
      28359: inst = 32'd136314880;
      28360: inst = 32'd268468224;
      28361: inst = 32'd201348616;
      28362: inst = 32'd203451216;
      28363: inst = 32'd471859200;
      28364: inst = 32'd136314880;
      28365: inst = 32'd268468224;
      28366: inst = 32'd201348617;
      28367: inst = 32'd203451216;
      28368: inst = 32'd471859200;
      28369: inst = 32'd136314880;
      28370: inst = 32'd268468224;
      28371: inst = 32'd201348618;
      28372: inst = 32'd203451216;
      28373: inst = 32'd471859200;
      28374: inst = 32'd136314880;
      28375: inst = 32'd268468224;
      28376: inst = 32'd201348619;
      28377: inst = 32'd203451216;
      28378: inst = 32'd471859200;
      28379: inst = 32'd136314880;
      28380: inst = 32'd268468224;
      28381: inst = 32'd201348620;
      28382: inst = 32'd203451216;
      28383: inst = 32'd471859200;
      28384: inst = 32'd136314880;
      28385: inst = 32'd268468224;
      28386: inst = 32'd201348621;
      28387: inst = 32'd203451216;
      28388: inst = 32'd471859200;
      28389: inst = 32'd136314880;
      28390: inst = 32'd268468224;
      28391: inst = 32'd201348622;
      28392: inst = 32'd203451216;
      28393: inst = 32'd471859200;
      28394: inst = 32'd136314880;
      28395: inst = 32'd268468224;
      28396: inst = 32'd201348623;
      28397: inst = 32'd203451216;
      28398: inst = 32'd471859200;
      28399: inst = 32'd136314880;
      28400: inst = 32'd268468224;
      28401: inst = 32'd201348624;
      28402: inst = 32'd203451216;
      28403: inst = 32'd471859200;
      28404: inst = 32'd136314880;
      28405: inst = 32'd268468224;
      28406: inst = 32'd201348625;
      28407: inst = 32'd203451216;
      28408: inst = 32'd471859200;
      28409: inst = 32'd136314880;
      28410: inst = 32'd268468224;
      28411: inst = 32'd201348626;
      28412: inst = 32'd203451216;
      28413: inst = 32'd471859200;
      28414: inst = 32'd136314880;
      28415: inst = 32'd268468224;
      28416: inst = 32'd201348627;
      28417: inst = 32'd203451216;
      28418: inst = 32'd471859200;
      28419: inst = 32'd136314880;
      28420: inst = 32'd268468224;
      28421: inst = 32'd201348628;
      28422: inst = 32'd203451216;
      28423: inst = 32'd471859200;
      28424: inst = 32'd136314880;
      28425: inst = 32'd268468224;
      28426: inst = 32'd201348629;
      28427: inst = 32'd203455473;
      28428: inst = 32'd471859200;
      28429: inst = 32'd136314880;
      28430: inst = 32'd268468224;
      28431: inst = 32'd201348630;
      28432: inst = 32'd203459697;
      28433: inst = 32'd471859200;
      28434: inst = 32'd136314880;
      28435: inst = 32'd268468224;
      28436: inst = 32'd201348631;
      28437: inst = 32'd203459697;
      28438: inst = 32'd471859200;
      28439: inst = 32'd136314880;
      28440: inst = 32'd268468224;
      28441: inst = 32'd201348632;
      28442: inst = 32'd203459665;
      28443: inst = 32'd471859200;
      28444: inst = 32'd136314880;
      28445: inst = 32'd268468224;
      28446: inst = 32'd201348633;
      28447: inst = 32'd203444906;
      28448: inst = 32'd471859200;
      28449: inst = 32'd136314880;
      28450: inst = 32'd268468224;
      28451: inst = 32'd201348634;
      28452: inst = 32'd203442793;
      28453: inst = 32'd471859200;
      28454: inst = 32'd136314880;
      28455: inst = 32'd268468224;
      28456: inst = 32'd201348635;
      28457: inst = 32'd203442793;
      28458: inst = 32'd471859200;
      28459: inst = 32'd136314880;
      28460: inst = 32'd268468224;
      28461: inst = 32'd201348636;
      28462: inst = 32'd203442793;
      28463: inst = 32'd471859200;
      28464: inst = 32'd136314880;
      28465: inst = 32'd268468224;
      28466: inst = 32'd201348637;
      28467: inst = 32'd203442793;
      28468: inst = 32'd471859200;
      28469: inst = 32'd136314880;
      28470: inst = 32'd268468224;
      28471: inst = 32'd201348638;
      28472: inst = 32'd203455439;
      28473: inst = 32'd471859200;
      28474: inst = 32'd136314880;
      28475: inst = 32'd268468224;
      28476: inst = 32'd201348639;
      28477: inst = 32'd203459697;
      28478: inst = 32'd471859200;
      28479: inst = 32'd136314880;
      28480: inst = 32'd268468224;
      28481: inst = 32'd201348640;
      28482: inst = 32'd203459697;
      28483: inst = 32'd471859200;
      28484: inst = 32'd136314880;
      28485: inst = 32'd268468224;
      28486: inst = 32'd201348641;
      28487: inst = 32'd203455439;
      28488: inst = 32'd471859200;
      28489: inst = 32'd136314880;
      28490: inst = 32'd268468224;
      28491: inst = 32'd201348642;
      28492: inst = 32'd203444906;
      28493: inst = 32'd471859200;
      28494: inst = 32'd136314880;
      28495: inst = 32'd268468224;
      28496: inst = 32'd201348643;
      28497: inst = 32'd203459697;
      28498: inst = 32'd471859200;
      28499: inst = 32'd136314880;
      28500: inst = 32'd268468224;
      28501: inst = 32'd201348644;
      28502: inst = 32'd203459697;
      28503: inst = 32'd471859200;
      28504: inst = 32'd136314880;
      28505: inst = 32'd268468224;
      28506: inst = 32'd201348645;
      28507: inst = 32'd203459697;
      28508: inst = 32'd471859200;
      28509: inst = 32'd136314880;
      28510: inst = 32'd268468224;
      28511: inst = 32'd201348646;
      28512: inst = 32'd203459697;
      28513: inst = 32'd471859200;
      28514: inst = 32'd136314880;
      28515: inst = 32'd268468224;
      28516: inst = 32'd201348647;
      28517: inst = 32'd203459665;
      28518: inst = 32'd471859200;
      28519: inst = 32'd136314880;
      28520: inst = 32'd268468224;
      28521: inst = 32'd201348648;
      28522: inst = 32'd203444874;
      28523: inst = 32'd471859200;
      28524: inst = 32'd136314880;
      28525: inst = 32'd268468224;
      28526: inst = 32'd201348649;
      28527: inst = 32'd203444874;
      28528: inst = 32'd471859200;
      28529: inst = 32'd136314880;
      28530: inst = 32'd268468224;
      28531: inst = 32'd201348650;
      28532: inst = 32'd203451216;
      28533: inst = 32'd471859200;
      28534: inst = 32'd136314880;
      28535: inst = 32'd268468224;
      28536: inst = 32'd201348651;
      28537: inst = 32'd203451216;
      28538: inst = 32'd471859200;
      28539: inst = 32'd136314880;
      28540: inst = 32'd268468224;
      28541: inst = 32'd201348652;
      28542: inst = 32'd203451216;
      28543: inst = 32'd471859200;
      28544: inst = 32'd136314880;
      28545: inst = 32'd268468224;
      28546: inst = 32'd201348653;
      28547: inst = 32'd203451216;
      28548: inst = 32'd471859200;
      28549: inst = 32'd136314880;
      28550: inst = 32'd268468224;
      28551: inst = 32'd201348654;
      28552: inst = 32'd203451216;
      28553: inst = 32'd471859200;
      28554: inst = 32'd136314880;
      28555: inst = 32'd268468224;
      28556: inst = 32'd201348655;
      28557: inst = 32'd203451216;
      28558: inst = 32'd471859200;
      28559: inst = 32'd136314880;
      28560: inst = 32'd268468224;
      28561: inst = 32'd201348656;
      28562: inst = 32'd203451216;
      28563: inst = 32'd471859200;
      28564: inst = 32'd136314880;
      28565: inst = 32'd268468224;
      28566: inst = 32'd201348657;
      28567: inst = 32'd203451216;
      28568: inst = 32'd471859200;
      28569: inst = 32'd136314880;
      28570: inst = 32'd268468224;
      28571: inst = 32'd201348658;
      28572: inst = 32'd203451216;
      28573: inst = 32'd471859200;
      28574: inst = 32'd136314880;
      28575: inst = 32'd268468224;
      28576: inst = 32'd201348659;
      28577: inst = 32'd203451216;
      28578: inst = 32'd471859200;
      28579: inst = 32'd136314880;
      28580: inst = 32'd268468224;
      28581: inst = 32'd201348660;
      28582: inst = 32'd203451216;
      28583: inst = 32'd471859200;
      28584: inst = 32'd136314880;
      28585: inst = 32'd268468224;
      28586: inst = 32'd201348661;
      28587: inst = 32'd203451216;
      28588: inst = 32'd471859200;
      28589: inst = 32'd136314880;
      28590: inst = 32'd268468224;
      28591: inst = 32'd201348662;
      28592: inst = 32'd203444874;
      28593: inst = 32'd471859200;
      28594: inst = 32'd136314880;
      28595: inst = 32'd268468224;
      28596: inst = 32'd201348663;
      28597: inst = 32'd203444874;
      28598: inst = 32'd471859200;
      28599: inst = 32'd136314880;
      28600: inst = 32'd268468224;
      28601: inst = 32'd201348664;
      28602: inst = 32'd203459665;
      28603: inst = 32'd471859200;
      28604: inst = 32'd136314880;
      28605: inst = 32'd268468224;
      28606: inst = 32'd201348665;
      28607: inst = 32'd203459697;
      28608: inst = 32'd471859200;
      28609: inst = 32'd136314880;
      28610: inst = 32'd268468224;
      28611: inst = 32'd201348666;
      28612: inst = 32'd203459697;
      28613: inst = 32'd471859200;
      28614: inst = 32'd136314880;
      28615: inst = 32'd268468224;
      28616: inst = 32'd201348667;
      28617: inst = 32'd203459697;
      28618: inst = 32'd471859200;
      28619: inst = 32'd136314880;
      28620: inst = 32'd268468224;
      28621: inst = 32'd201348668;
      28622: inst = 32'd203459697;
      28623: inst = 32'd471859200;
      28624: inst = 32'd136314880;
      28625: inst = 32'd268468224;
      28626: inst = 32'd201348669;
      28627: inst = 32'd203444906;
      28628: inst = 32'd471859200;
      28629: inst = 32'd136314880;
      28630: inst = 32'd268468224;
      28631: inst = 32'd201348670;
      28632: inst = 32'd203455439;
      28633: inst = 32'd471859200;
      28634: inst = 32'd136314880;
      28635: inst = 32'd268468224;
      28636: inst = 32'd201348671;
      28637: inst = 32'd203459697;
      28638: inst = 32'd471859200;
      28639: inst = 32'd136314880;
      28640: inst = 32'd268468224;
      28641: inst = 32'd201348672;
      28642: inst = 32'd203459697;
      28643: inst = 32'd471859200;
      28644: inst = 32'd136314880;
      28645: inst = 32'd268468224;
      28646: inst = 32'd201348673;
      28647: inst = 32'd203455439;
      28648: inst = 32'd471859200;
      28649: inst = 32'd136314880;
      28650: inst = 32'd268468224;
      28651: inst = 32'd201348674;
      28652: inst = 32'd203442793;
      28653: inst = 32'd471859200;
      28654: inst = 32'd136314880;
      28655: inst = 32'd268468224;
      28656: inst = 32'd201348675;
      28657: inst = 32'd203442793;
      28658: inst = 32'd471859200;
      28659: inst = 32'd136314880;
      28660: inst = 32'd268468224;
      28661: inst = 32'd201348676;
      28662: inst = 32'd203442793;
      28663: inst = 32'd471859200;
      28664: inst = 32'd136314880;
      28665: inst = 32'd268468224;
      28666: inst = 32'd201348677;
      28667: inst = 32'd203442793;
      28668: inst = 32'd471859200;
      28669: inst = 32'd136314880;
      28670: inst = 32'd268468224;
      28671: inst = 32'd201348678;
      28672: inst = 32'd203444906;
      28673: inst = 32'd471859200;
      28674: inst = 32'd136314880;
      28675: inst = 32'd268468224;
      28676: inst = 32'd201348679;
      28677: inst = 32'd203459665;
      28678: inst = 32'd471859200;
      28679: inst = 32'd136314880;
      28680: inst = 32'd268468224;
      28681: inst = 32'd201348680;
      28682: inst = 32'd203459697;
      28683: inst = 32'd471859200;
      28684: inst = 32'd136314880;
      28685: inst = 32'd268468224;
      28686: inst = 32'd201348681;
      28687: inst = 32'd203459697;
      28688: inst = 32'd471859200;
      28689: inst = 32'd136314880;
      28690: inst = 32'd268468224;
      28691: inst = 32'd201348682;
      28692: inst = 32'd203455473;
      28693: inst = 32'd471859200;
      28694: inst = 32'd136314880;
      28695: inst = 32'd268468224;
      28696: inst = 32'd201348683;
      28697: inst = 32'd203451216;
      28698: inst = 32'd471859200;
      28699: inst = 32'd136314880;
      28700: inst = 32'd268468224;
      28701: inst = 32'd201348684;
      28702: inst = 32'd203451216;
      28703: inst = 32'd471859200;
      28704: inst = 32'd136314880;
      28705: inst = 32'd268468224;
      28706: inst = 32'd201348685;
      28707: inst = 32'd203451216;
      28708: inst = 32'd471859200;
      28709: inst = 32'd136314880;
      28710: inst = 32'd268468224;
      28711: inst = 32'd201348686;
      28712: inst = 32'd203451216;
      28713: inst = 32'd471859200;
      28714: inst = 32'd136314880;
      28715: inst = 32'd268468224;
      28716: inst = 32'd201348687;
      28717: inst = 32'd203451216;
      28718: inst = 32'd471859200;
      28719: inst = 32'd136314880;
      28720: inst = 32'd268468224;
      28721: inst = 32'd201348688;
      28722: inst = 32'd203451216;
      28723: inst = 32'd471859200;
      28724: inst = 32'd136314880;
      28725: inst = 32'd268468224;
      28726: inst = 32'd201348689;
      28727: inst = 32'd203451216;
      28728: inst = 32'd471859200;
      28729: inst = 32'd136314880;
      28730: inst = 32'd268468224;
      28731: inst = 32'd201348690;
      28732: inst = 32'd203451216;
      28733: inst = 32'd471859200;
      28734: inst = 32'd136314880;
      28735: inst = 32'd268468224;
      28736: inst = 32'd201348691;
      28737: inst = 32'd203451216;
      28738: inst = 32'd471859200;
      28739: inst = 32'd136314880;
      28740: inst = 32'd268468224;
      28741: inst = 32'd201348692;
      28742: inst = 32'd203451216;
      28743: inst = 32'd471859200;
      28744: inst = 32'd136314880;
      28745: inst = 32'd268468224;
      28746: inst = 32'd201348693;
      28747: inst = 32'd203451216;
      28748: inst = 32'd471859200;
      28749: inst = 32'd136314880;
      28750: inst = 32'd268468224;
      28751: inst = 32'd201348694;
      28752: inst = 32'd203451216;
      28753: inst = 32'd471859200;
      28754: inst = 32'd136314880;
      28755: inst = 32'd268468224;
      28756: inst = 32'd201348695;
      28757: inst = 32'd203451216;
      28758: inst = 32'd471859200;
      28759: inst = 32'd136314880;
      28760: inst = 32'd268468224;
      28761: inst = 32'd201348696;
      28762: inst = 32'd203451216;
      28763: inst = 32'd471859200;
      28764: inst = 32'd136314880;
      28765: inst = 32'd268468224;
      28766: inst = 32'd201348697;
      28767: inst = 32'd203451216;
      28768: inst = 32'd471859200;
      28769: inst = 32'd136314880;
      28770: inst = 32'd268468224;
      28771: inst = 32'd201348698;
      28772: inst = 32'd203451216;
      28773: inst = 32'd471859200;
      28774: inst = 32'd136314880;
      28775: inst = 32'd268468224;
      28776: inst = 32'd201348699;
      28777: inst = 32'd203451216;
      28778: inst = 32'd471859200;
      28779: inst = 32'd136314880;
      28780: inst = 32'd268468224;
      28781: inst = 32'd201348700;
      28782: inst = 32'd203451216;
      28783: inst = 32'd471859200;
      28784: inst = 32'd136314880;
      28785: inst = 32'd268468224;
      28786: inst = 32'd201348701;
      28787: inst = 32'd203451216;
      28788: inst = 32'd471859200;
      28789: inst = 32'd136314880;
      28790: inst = 32'd268468224;
      28791: inst = 32'd201348702;
      28792: inst = 32'd203451216;
      28793: inst = 32'd471859200;
      28794: inst = 32'd136314880;
      28795: inst = 32'd268468224;
      28796: inst = 32'd201348703;
      28797: inst = 32'd203451216;
      28798: inst = 32'd471859200;
      28799: inst = 32'd136314880;
      28800: inst = 32'd268468224;
      28801: inst = 32'd201348704;
      28802: inst = 32'd203451216;
      28803: inst = 32'd471859200;
      28804: inst = 32'd136314880;
      28805: inst = 32'd268468224;
      28806: inst = 32'd201348705;
      28807: inst = 32'd203451216;
      28808: inst = 32'd471859200;
      28809: inst = 32'd136314880;
      28810: inst = 32'd268468224;
      28811: inst = 32'd201348706;
      28812: inst = 32'd203451216;
      28813: inst = 32'd471859200;
      28814: inst = 32'd136314880;
      28815: inst = 32'd268468224;
      28816: inst = 32'd201348707;
      28817: inst = 32'd203451216;
      28818: inst = 32'd471859200;
      28819: inst = 32'd136314880;
      28820: inst = 32'd268468224;
      28821: inst = 32'd201348708;
      28822: inst = 32'd203451216;
      28823: inst = 32'd471859200;
      28824: inst = 32'd136314880;
      28825: inst = 32'd268468224;
      28826: inst = 32'd201348709;
      28827: inst = 32'd203451216;
      28828: inst = 32'd471859200;
      28829: inst = 32'd136314880;
      28830: inst = 32'd268468224;
      28831: inst = 32'd201348710;
      28832: inst = 32'd203451216;
      28833: inst = 32'd471859200;
      28834: inst = 32'd136314880;
      28835: inst = 32'd268468224;
      28836: inst = 32'd201348711;
      28837: inst = 32'd203451216;
      28838: inst = 32'd471859200;
      28839: inst = 32'd136314880;
      28840: inst = 32'd268468224;
      28841: inst = 32'd201348712;
      28842: inst = 32'd203451216;
      28843: inst = 32'd471859200;
      28844: inst = 32'd136314880;
      28845: inst = 32'd268468224;
      28846: inst = 32'd201348713;
      28847: inst = 32'd203451216;
      28848: inst = 32'd471859200;
      28849: inst = 32'd136314880;
      28850: inst = 32'd268468224;
      28851: inst = 32'd201348714;
      28852: inst = 32'd203451216;
      28853: inst = 32'd471859200;
      28854: inst = 32'd136314880;
      28855: inst = 32'd268468224;
      28856: inst = 32'd201348715;
      28857: inst = 32'd203451216;
      28858: inst = 32'd471859200;
      28859: inst = 32'd136314880;
      28860: inst = 32'd268468224;
      28861: inst = 32'd201348716;
      28862: inst = 32'd203451216;
      28863: inst = 32'd471859200;
      28864: inst = 32'd136314880;
      28865: inst = 32'd268468224;
      28866: inst = 32'd201348717;
      28867: inst = 32'd203451216;
      28868: inst = 32'd471859200;
      28869: inst = 32'd136314880;
      28870: inst = 32'd268468224;
      28871: inst = 32'd201348718;
      28872: inst = 32'd203451216;
      28873: inst = 32'd471859200;
      28874: inst = 32'd136314880;
      28875: inst = 32'd268468224;
      28876: inst = 32'd201348719;
      28877: inst = 32'd203451216;
      28878: inst = 32'd471859200;
      28879: inst = 32'd136314880;
      28880: inst = 32'd268468224;
      28881: inst = 32'd201348720;
      28882: inst = 32'd203451216;
      28883: inst = 32'd471859200;
      28884: inst = 32'd136314880;
      28885: inst = 32'd268468224;
      28886: inst = 32'd201348721;
      28887: inst = 32'd203451216;
      28888: inst = 32'd471859200;
      28889: inst = 32'd136314880;
      28890: inst = 32'd268468224;
      28891: inst = 32'd201348722;
      28892: inst = 32'd203451216;
      28893: inst = 32'd471859200;
      28894: inst = 32'd136314880;
      28895: inst = 32'd268468224;
      28896: inst = 32'd201348723;
      28897: inst = 32'd203451216;
      28898: inst = 32'd471859200;
      28899: inst = 32'd136314880;
      28900: inst = 32'd268468224;
      28901: inst = 32'd201348724;
      28902: inst = 32'd203453360;
      28903: inst = 32'd471859200;
      28904: inst = 32'd136314880;
      28905: inst = 32'd268468224;
      28906: inst = 32'd201348725;
      28907: inst = 32'd203459697;
      28908: inst = 32'd471859200;
      28909: inst = 32'd136314880;
      28910: inst = 32'd268468224;
      28911: inst = 32'd201348726;
      28912: inst = 32'd203459697;
      28913: inst = 32'd471859200;
      28914: inst = 32'd136314880;
      28915: inst = 32'd268468224;
      28916: inst = 32'd201348727;
      28917: inst = 32'd203459697;
      28918: inst = 32'd471859200;
      28919: inst = 32'd136314880;
      28920: inst = 32'd268468224;
      28921: inst = 32'd201348728;
      28922: inst = 32'd203449100;
      28923: inst = 32'd471859200;
      28924: inst = 32'd136314880;
      28925: inst = 32'd268468224;
      28926: inst = 32'd201348729;
      28927: inst = 32'd203442793;
      28928: inst = 32'd471859200;
      28929: inst = 32'd136314880;
      28930: inst = 32'd268468224;
      28931: inst = 32'd201348730;
      28932: inst = 32'd203442793;
      28933: inst = 32'd471859200;
      28934: inst = 32'd136314880;
      28935: inst = 32'd268468224;
      28936: inst = 32'd201348731;
      28937: inst = 32'd203442793;
      28938: inst = 32'd471859200;
      28939: inst = 32'd136314880;
      28940: inst = 32'd268468224;
      28941: inst = 32'd201348732;
      28942: inst = 32'd203442793;
      28943: inst = 32'd471859200;
      28944: inst = 32'd136314880;
      28945: inst = 32'd268468224;
      28946: inst = 32'd201348733;
      28947: inst = 32'd203444874;
      28948: inst = 32'd471859200;
      28949: inst = 32'd136314880;
      28950: inst = 32'd268468224;
      28951: inst = 32'd201348734;
      28952: inst = 32'd203459697;
      28953: inst = 32'd471859200;
      28954: inst = 32'd136314880;
      28955: inst = 32'd268468224;
      28956: inst = 32'd201348735;
      28957: inst = 32'd203459697;
      28958: inst = 32'd471859200;
      28959: inst = 32'd136314880;
      28960: inst = 32'd268468224;
      28961: inst = 32'd201348736;
      28962: inst = 32'd203459697;
      28963: inst = 32'd471859200;
      28964: inst = 32'd136314880;
      28965: inst = 32'd268468224;
      28966: inst = 32'd201348737;
      28967: inst = 32'd203455439;
      28968: inst = 32'd471859200;
      28969: inst = 32'd136314880;
      28970: inst = 32'd268468224;
      28971: inst = 32'd201348738;
      28972: inst = 32'd203451213;
      28973: inst = 32'd471859200;
      28974: inst = 32'd136314880;
      28975: inst = 32'd268468224;
      28976: inst = 32'd201348739;
      28977: inst = 32'd203459697;
      28978: inst = 32'd471859200;
      28979: inst = 32'd136314880;
      28980: inst = 32'd268468224;
      28981: inst = 32'd201348740;
      28982: inst = 32'd203459697;
      28983: inst = 32'd471859200;
      28984: inst = 32'd136314880;
      28985: inst = 32'd268468224;
      28986: inst = 32'd201348741;
      28987: inst = 32'd203459697;
      28988: inst = 32'd471859200;
      28989: inst = 32'd136314880;
      28990: inst = 32'd268468224;
      28991: inst = 32'd201348742;
      28992: inst = 32'd203459697;
      28993: inst = 32'd471859200;
      28994: inst = 32'd136314880;
      28995: inst = 32'd268468224;
      28996: inst = 32'd201348743;
      28997: inst = 32'd203455471;
      28998: inst = 32'd471859200;
      28999: inst = 32'd136314880;
      29000: inst = 32'd268468224;
      29001: inst = 32'd201348744;
      29002: inst = 32'd203444874;
      29003: inst = 32'd471859200;
      29004: inst = 32'd136314880;
      29005: inst = 32'd268468224;
      29006: inst = 32'd201348745;
      29007: inst = 32'd203444874;
      29008: inst = 32'd471859200;
      29009: inst = 32'd136314880;
      29010: inst = 32'd268468224;
      29011: inst = 32'd201348746;
      29012: inst = 32'd203451216;
      29013: inst = 32'd471859200;
      29014: inst = 32'd136314880;
      29015: inst = 32'd268468224;
      29016: inst = 32'd201348747;
      29017: inst = 32'd203451216;
      29018: inst = 32'd471859200;
      29019: inst = 32'd136314880;
      29020: inst = 32'd268468224;
      29021: inst = 32'd201348748;
      29022: inst = 32'd203451216;
      29023: inst = 32'd471859200;
      29024: inst = 32'd136314880;
      29025: inst = 32'd268468224;
      29026: inst = 32'd201348749;
      29027: inst = 32'd203451216;
      29028: inst = 32'd471859200;
      29029: inst = 32'd136314880;
      29030: inst = 32'd268468224;
      29031: inst = 32'd201348750;
      29032: inst = 32'd203451216;
      29033: inst = 32'd471859200;
      29034: inst = 32'd136314880;
      29035: inst = 32'd268468224;
      29036: inst = 32'd201348751;
      29037: inst = 32'd203451216;
      29038: inst = 32'd471859200;
      29039: inst = 32'd136314880;
      29040: inst = 32'd268468224;
      29041: inst = 32'd201348752;
      29042: inst = 32'd203451216;
      29043: inst = 32'd471859200;
      29044: inst = 32'd136314880;
      29045: inst = 32'd268468224;
      29046: inst = 32'd201348753;
      29047: inst = 32'd203451216;
      29048: inst = 32'd471859200;
      29049: inst = 32'd136314880;
      29050: inst = 32'd268468224;
      29051: inst = 32'd201348754;
      29052: inst = 32'd203451216;
      29053: inst = 32'd471859200;
      29054: inst = 32'd136314880;
      29055: inst = 32'd268468224;
      29056: inst = 32'd201348755;
      29057: inst = 32'd203451216;
      29058: inst = 32'd471859200;
      29059: inst = 32'd136314880;
      29060: inst = 32'd268468224;
      29061: inst = 32'd201348756;
      29062: inst = 32'd203451216;
      29063: inst = 32'd471859200;
      29064: inst = 32'd136314880;
      29065: inst = 32'd268468224;
      29066: inst = 32'd201348757;
      29067: inst = 32'd203451216;
      29068: inst = 32'd471859200;
      29069: inst = 32'd136314880;
      29070: inst = 32'd268468224;
      29071: inst = 32'd201348758;
      29072: inst = 32'd203444874;
      29073: inst = 32'd471859200;
      29074: inst = 32'd136314880;
      29075: inst = 32'd268468224;
      29076: inst = 32'd201348759;
      29077: inst = 32'd203444874;
      29078: inst = 32'd471859200;
      29079: inst = 32'd136314880;
      29080: inst = 32'd268468224;
      29081: inst = 32'd201348760;
      29082: inst = 32'd203455439;
      29083: inst = 32'd471859200;
      29084: inst = 32'd136314880;
      29085: inst = 32'd268468224;
      29086: inst = 32'd201348761;
      29087: inst = 32'd203459697;
      29088: inst = 32'd471859200;
      29089: inst = 32'd136314880;
      29090: inst = 32'd268468224;
      29091: inst = 32'd201348762;
      29092: inst = 32'd203459697;
      29093: inst = 32'd471859200;
      29094: inst = 32'd136314880;
      29095: inst = 32'd268468224;
      29096: inst = 32'd201348763;
      29097: inst = 32'd203459697;
      29098: inst = 32'd471859200;
      29099: inst = 32'd136314880;
      29100: inst = 32'd268468224;
      29101: inst = 32'd201348764;
      29102: inst = 32'd203459697;
      29103: inst = 32'd471859200;
      29104: inst = 32'd136314880;
      29105: inst = 32'd268468224;
      29106: inst = 32'd201348765;
      29107: inst = 32'd203451213;
      29108: inst = 32'd471859200;
      29109: inst = 32'd136314880;
      29110: inst = 32'd268468224;
      29111: inst = 32'd201348766;
      29112: inst = 32'd203455439;
      29113: inst = 32'd471859200;
      29114: inst = 32'd136314880;
      29115: inst = 32'd268468224;
      29116: inst = 32'd201348767;
      29117: inst = 32'd203459697;
      29118: inst = 32'd471859200;
      29119: inst = 32'd136314880;
      29120: inst = 32'd268468224;
      29121: inst = 32'd201348768;
      29122: inst = 32'd203459697;
      29123: inst = 32'd471859200;
      29124: inst = 32'd136314880;
      29125: inst = 32'd268468224;
      29126: inst = 32'd201348769;
      29127: inst = 32'd203459697;
      29128: inst = 32'd471859200;
      29129: inst = 32'd136314880;
      29130: inst = 32'd268468224;
      29131: inst = 32'd201348770;
      29132: inst = 32'd203444874;
      29133: inst = 32'd471859200;
      29134: inst = 32'd136314880;
      29135: inst = 32'd268468224;
      29136: inst = 32'd201348771;
      29137: inst = 32'd203442793;
      29138: inst = 32'd471859200;
      29139: inst = 32'd136314880;
      29140: inst = 32'd268468224;
      29141: inst = 32'd201348772;
      29142: inst = 32'd203442793;
      29143: inst = 32'd471859200;
      29144: inst = 32'd136314880;
      29145: inst = 32'd268468224;
      29146: inst = 32'd201348773;
      29147: inst = 32'd203442793;
      29148: inst = 32'd471859200;
      29149: inst = 32'd136314880;
      29150: inst = 32'd268468224;
      29151: inst = 32'd201348774;
      29152: inst = 32'd203442793;
      29153: inst = 32'd471859200;
      29154: inst = 32'd136314880;
      29155: inst = 32'd268468224;
      29156: inst = 32'd201348775;
      29157: inst = 32'd203449132;
      29158: inst = 32'd471859200;
      29159: inst = 32'd136314880;
      29160: inst = 32'd268468224;
      29161: inst = 32'd201348776;
      29162: inst = 32'd203459697;
      29163: inst = 32'd471859200;
      29164: inst = 32'd136314880;
      29165: inst = 32'd268468224;
      29166: inst = 32'd201348777;
      29167: inst = 32'd203459697;
      29168: inst = 32'd471859200;
      29169: inst = 32'd136314880;
      29170: inst = 32'd268468224;
      29171: inst = 32'd201348778;
      29172: inst = 32'd203459697;
      29173: inst = 32'd471859200;
      29174: inst = 32'd136314880;
      29175: inst = 32'd268468224;
      29176: inst = 32'd201348779;
      29177: inst = 32'd203453360;
      29178: inst = 32'd471859200;
      29179: inst = 32'd136314880;
      29180: inst = 32'd268468224;
      29181: inst = 32'd201348780;
      29182: inst = 32'd203451216;
      29183: inst = 32'd471859200;
      29184: inst = 32'd136314880;
      29185: inst = 32'd268468224;
      29186: inst = 32'd201348781;
      29187: inst = 32'd203451216;
      29188: inst = 32'd471859200;
      29189: inst = 32'd136314880;
      29190: inst = 32'd268468224;
      29191: inst = 32'd201348782;
      29192: inst = 32'd203451216;
      29193: inst = 32'd471859200;
      29194: inst = 32'd136314880;
      29195: inst = 32'd268468224;
      29196: inst = 32'd201348783;
      29197: inst = 32'd203451216;
      29198: inst = 32'd471859200;
      29199: inst = 32'd136314880;
      29200: inst = 32'd268468224;
      29201: inst = 32'd201348784;
      29202: inst = 32'd203451216;
      29203: inst = 32'd471859200;
      29204: inst = 32'd136314880;
      29205: inst = 32'd268468224;
      29206: inst = 32'd201348785;
      29207: inst = 32'd203451216;
      29208: inst = 32'd471859200;
      29209: inst = 32'd136314880;
      29210: inst = 32'd268468224;
      29211: inst = 32'd201348786;
      29212: inst = 32'd203451216;
      29213: inst = 32'd471859200;
      29214: inst = 32'd136314880;
      29215: inst = 32'd268468224;
      29216: inst = 32'd201348787;
      29217: inst = 32'd203451216;
      29218: inst = 32'd471859200;
      29219: inst = 32'd136314880;
      29220: inst = 32'd268468224;
      29221: inst = 32'd201348788;
      29222: inst = 32'd203451216;
      29223: inst = 32'd471859200;
      29224: inst = 32'd136314880;
      29225: inst = 32'd268468224;
      29226: inst = 32'd201348789;
      29227: inst = 32'd203451216;
      29228: inst = 32'd471859200;
      29229: inst = 32'd136314880;
      29230: inst = 32'd268468224;
      29231: inst = 32'd201348790;
      29232: inst = 32'd203451216;
      29233: inst = 32'd471859200;
      29234: inst = 32'd136314880;
      29235: inst = 32'd268468224;
      29236: inst = 32'd201348791;
      29237: inst = 32'd203451216;
      29238: inst = 32'd471859200;
      29239: inst = 32'd136314880;
      29240: inst = 32'd268468224;
      29241: inst = 32'd201348792;
      29242: inst = 32'd203451216;
      29243: inst = 32'd471859200;
      29244: inst = 32'd136314880;
      29245: inst = 32'd268468224;
      29246: inst = 32'd201348793;
      29247: inst = 32'd203451216;
      29248: inst = 32'd471859200;
      29249: inst = 32'd136314880;
      29250: inst = 32'd268468224;
      29251: inst = 32'd201348794;
      29252: inst = 32'd203451216;
      29253: inst = 32'd471859200;
      29254: inst = 32'd136314880;
      29255: inst = 32'd268468224;
      29256: inst = 32'd201348795;
      29257: inst = 32'd203451216;
      29258: inst = 32'd471859200;
      29259: inst = 32'd136314880;
      29260: inst = 32'd268468224;
      29261: inst = 32'd201348796;
      29262: inst = 32'd203451216;
      29263: inst = 32'd471859200;
      29264: inst = 32'd136314880;
      29265: inst = 32'd268468224;
      29266: inst = 32'd201348797;
      29267: inst = 32'd203451216;
      29268: inst = 32'd471859200;
      29269: inst = 32'd136314880;
      29270: inst = 32'd268468224;
      29271: inst = 32'd201348798;
      29272: inst = 32'd203451216;
      29273: inst = 32'd471859200;
      29274: inst = 32'd136314880;
      29275: inst = 32'd268468224;
      29276: inst = 32'd201348799;
      29277: inst = 32'd203451216;
      29278: inst = 32'd471859200;
      29279: inst = 32'd136314880;
      29280: inst = 32'd268468224;
      29281: inst = 32'd201348800;
      29282: inst = 32'd203451216;
      29283: inst = 32'd471859200;
      29284: inst = 32'd136314880;
      29285: inst = 32'd268468224;
      29286: inst = 32'd201348801;
      29287: inst = 32'd203451216;
      29288: inst = 32'd471859200;
      29289: inst = 32'd136314880;
      29290: inst = 32'd268468224;
      29291: inst = 32'd201348802;
      29292: inst = 32'd203451216;
      29293: inst = 32'd471859200;
      29294: inst = 32'd136314880;
      29295: inst = 32'd268468224;
      29296: inst = 32'd201348803;
      29297: inst = 32'd203451216;
      29298: inst = 32'd471859200;
      29299: inst = 32'd136314880;
      29300: inst = 32'd268468224;
      29301: inst = 32'd201348804;
      29302: inst = 32'd203451216;
      29303: inst = 32'd471859200;
      29304: inst = 32'd136314880;
      29305: inst = 32'd268468224;
      29306: inst = 32'd201348805;
      29307: inst = 32'd203451216;
      29308: inst = 32'd471859200;
      29309: inst = 32'd136314880;
      29310: inst = 32'd268468224;
      29311: inst = 32'd201348806;
      29312: inst = 32'd203451216;
      29313: inst = 32'd471859200;
      29314: inst = 32'd136314880;
      29315: inst = 32'd268468224;
      29316: inst = 32'd201348807;
      29317: inst = 32'd203451216;
      29318: inst = 32'd471859200;
      29319: inst = 32'd136314880;
      29320: inst = 32'd268468224;
      29321: inst = 32'd201348808;
      29322: inst = 32'd203451216;
      29323: inst = 32'd471859200;
      29324: inst = 32'd136314880;
      29325: inst = 32'd268468224;
      29326: inst = 32'd201348809;
      29327: inst = 32'd203451216;
      29328: inst = 32'd471859200;
      29329: inst = 32'd136314880;
      29330: inst = 32'd268468224;
      29331: inst = 32'd201348810;
      29332: inst = 32'd203451216;
      29333: inst = 32'd471859200;
      29334: inst = 32'd136314880;
      29335: inst = 32'd268468224;
      29336: inst = 32'd201348811;
      29337: inst = 32'd203451216;
      29338: inst = 32'd471859200;
      29339: inst = 32'd136314880;
      29340: inst = 32'd268468224;
      29341: inst = 32'd201348812;
      29342: inst = 32'd203451216;
      29343: inst = 32'd471859200;
      29344: inst = 32'd136314880;
      29345: inst = 32'd268468224;
      29346: inst = 32'd201348813;
      29347: inst = 32'd203451216;
      29348: inst = 32'd471859200;
      29349: inst = 32'd136314880;
      29350: inst = 32'd268468224;
      29351: inst = 32'd201348814;
      29352: inst = 32'd203451216;
      29353: inst = 32'd471859200;
      29354: inst = 32'd136314880;
      29355: inst = 32'd268468224;
      29356: inst = 32'd201348815;
      29357: inst = 32'd203451216;
      29358: inst = 32'd471859200;
      29359: inst = 32'd136314880;
      29360: inst = 32'd268468224;
      29361: inst = 32'd201348816;
      29362: inst = 32'd203451216;
      29363: inst = 32'd471859200;
      29364: inst = 32'd136314880;
      29365: inst = 32'd268468224;
      29366: inst = 32'd201348817;
      29367: inst = 32'd203451216;
      29368: inst = 32'd471859200;
      29369: inst = 32'd136314880;
      29370: inst = 32'd268468224;
      29371: inst = 32'd201348818;
      29372: inst = 32'd203451216;
      29373: inst = 32'd471859200;
      29374: inst = 32'd136314880;
      29375: inst = 32'd268468224;
      29376: inst = 32'd201348819;
      29377: inst = 32'd203451280;
      29378: inst = 32'd471859200;
      29379: inst = 32'd136314880;
      29380: inst = 32'd268468224;
      29381: inst = 32'd201348820;
      29382: inst = 32'd203459697;
      29383: inst = 32'd471859200;
      29384: inst = 32'd136314880;
      29385: inst = 32'd268468224;
      29386: inst = 32'd201348821;
      29387: inst = 32'd203459697;
      29388: inst = 32'd471859200;
      29389: inst = 32'd136314880;
      29390: inst = 32'd268468224;
      29391: inst = 32'd201348822;
      29392: inst = 32'd203459697;
      29393: inst = 32'd471859200;
      29394: inst = 32'd136314880;
      29395: inst = 32'd268468224;
      29396: inst = 32'd201348823;
      29397: inst = 32'd203459697;
      29398: inst = 32'd471859200;
      29399: inst = 32'd136314880;
      29400: inst = 32'd268468224;
      29401: inst = 32'd201348824;
      29402: inst = 32'd203459697;
      29403: inst = 32'd471859200;
      29404: inst = 32'd136314880;
      29405: inst = 32'd268468224;
      29406: inst = 32'd201348825;
      29407: inst = 32'd203459697;
      29408: inst = 32'd471859200;
      29409: inst = 32'd136314880;
      29410: inst = 32'd268468224;
      29411: inst = 32'd201348826;
      29412: inst = 32'd203459697;
      29413: inst = 32'd471859200;
      29414: inst = 32'd136314880;
      29415: inst = 32'd268468224;
      29416: inst = 32'd201348827;
      29417: inst = 32'd203459697;
      29418: inst = 32'd471859200;
      29419: inst = 32'd136314880;
      29420: inst = 32'd268468224;
      29421: inst = 32'd201348828;
      29422: inst = 32'd203459697;
      29423: inst = 32'd471859200;
      29424: inst = 32'd136314880;
      29425: inst = 32'd268468224;
      29426: inst = 32'd201348829;
      29427: inst = 32'd203459697;
      29428: inst = 32'd471859200;
      29429: inst = 32'd136314880;
      29430: inst = 32'd268468224;
      29431: inst = 32'd201348830;
      29432: inst = 32'd203459697;
      29433: inst = 32'd471859200;
      29434: inst = 32'd136314880;
      29435: inst = 32'd268468224;
      29436: inst = 32'd201348831;
      29437: inst = 32'd203459697;
      29438: inst = 32'd471859200;
      29439: inst = 32'd136314880;
      29440: inst = 32'd268468224;
      29441: inst = 32'd201348832;
      29442: inst = 32'd203459697;
      29443: inst = 32'd471859200;
      29444: inst = 32'd136314880;
      29445: inst = 32'd268468224;
      29446: inst = 32'd201348833;
      29447: inst = 32'd203455439;
      29448: inst = 32'd471859200;
      29449: inst = 32'd136314880;
      29450: inst = 32'd268468224;
      29451: inst = 32'd201348834;
      29452: inst = 32'd203455471;
      29453: inst = 32'd471859200;
      29454: inst = 32'd136314880;
      29455: inst = 32'd268468224;
      29456: inst = 32'd201348835;
      29457: inst = 32'd203459697;
      29458: inst = 32'd471859200;
      29459: inst = 32'd136314880;
      29460: inst = 32'd268468224;
      29461: inst = 32'd201348836;
      29462: inst = 32'd203459697;
      29463: inst = 32'd471859200;
      29464: inst = 32'd136314880;
      29465: inst = 32'd268468224;
      29466: inst = 32'd201348837;
      29467: inst = 32'd203459697;
      29468: inst = 32'd471859200;
      29469: inst = 32'd136314880;
      29470: inst = 32'd268468224;
      29471: inst = 32'd201348838;
      29472: inst = 32'd203459697;
      29473: inst = 32'd471859200;
      29474: inst = 32'd136314880;
      29475: inst = 32'd268468224;
      29476: inst = 32'd201348839;
      29477: inst = 32'd203451246;
      29478: inst = 32'd471859200;
      29479: inst = 32'd136314880;
      29480: inst = 32'd268468224;
      29481: inst = 32'd201348840;
      29482: inst = 32'd203444874;
      29483: inst = 32'd471859200;
      29484: inst = 32'd136314880;
      29485: inst = 32'd268468224;
      29486: inst = 32'd201348841;
      29487: inst = 32'd203444874;
      29488: inst = 32'd471859200;
      29489: inst = 32'd136314880;
      29490: inst = 32'd268468224;
      29491: inst = 32'd201348842;
      29492: inst = 32'd203451216;
      29493: inst = 32'd471859200;
      29494: inst = 32'd136314880;
      29495: inst = 32'd268468224;
      29496: inst = 32'd201348843;
      29497: inst = 32'd203451216;
      29498: inst = 32'd471859200;
      29499: inst = 32'd136314880;
      29500: inst = 32'd268468224;
      29501: inst = 32'd201348844;
      29502: inst = 32'd203451216;
      29503: inst = 32'd471859200;
      29504: inst = 32'd136314880;
      29505: inst = 32'd268468224;
      29506: inst = 32'd201348845;
      29507: inst = 32'd203451216;
      29508: inst = 32'd471859200;
      29509: inst = 32'd136314880;
      29510: inst = 32'd268468224;
      29511: inst = 32'd201348846;
      29512: inst = 32'd203451216;
      29513: inst = 32'd471859200;
      29514: inst = 32'd136314880;
      29515: inst = 32'd268468224;
      29516: inst = 32'd201348847;
      29517: inst = 32'd203451216;
      29518: inst = 32'd471859200;
      29519: inst = 32'd136314880;
      29520: inst = 32'd268468224;
      29521: inst = 32'd201348848;
      29522: inst = 32'd203451216;
      29523: inst = 32'd471859200;
      29524: inst = 32'd136314880;
      29525: inst = 32'd268468224;
      29526: inst = 32'd201348849;
      29527: inst = 32'd203451216;
      29528: inst = 32'd471859200;
      29529: inst = 32'd136314880;
      29530: inst = 32'd268468224;
      29531: inst = 32'd201348850;
      29532: inst = 32'd203451216;
      29533: inst = 32'd471859200;
      29534: inst = 32'd136314880;
      29535: inst = 32'd268468224;
      29536: inst = 32'd201348851;
      29537: inst = 32'd203451216;
      29538: inst = 32'd471859200;
      29539: inst = 32'd136314880;
      29540: inst = 32'd268468224;
      29541: inst = 32'd201348852;
      29542: inst = 32'd203451216;
      29543: inst = 32'd471859200;
      29544: inst = 32'd136314880;
      29545: inst = 32'd268468224;
      29546: inst = 32'd201348853;
      29547: inst = 32'd203451216;
      29548: inst = 32'd471859200;
      29549: inst = 32'd136314880;
      29550: inst = 32'd268468224;
      29551: inst = 32'd201348854;
      29552: inst = 32'd203444874;
      29553: inst = 32'd471859200;
      29554: inst = 32'd136314880;
      29555: inst = 32'd268468224;
      29556: inst = 32'd201348855;
      29557: inst = 32'd203444874;
      29558: inst = 32'd471859200;
      29559: inst = 32'd136314880;
      29560: inst = 32'd268468224;
      29561: inst = 32'd201348856;
      29562: inst = 32'd203451246;
      29563: inst = 32'd471859200;
      29564: inst = 32'd136314880;
      29565: inst = 32'd268468224;
      29566: inst = 32'd201348857;
      29567: inst = 32'd203459697;
      29568: inst = 32'd471859200;
      29569: inst = 32'd136314880;
      29570: inst = 32'd268468224;
      29571: inst = 32'd201348858;
      29572: inst = 32'd203459697;
      29573: inst = 32'd471859200;
      29574: inst = 32'd136314880;
      29575: inst = 32'd268468224;
      29576: inst = 32'd201348859;
      29577: inst = 32'd203459697;
      29578: inst = 32'd471859200;
      29579: inst = 32'd136314880;
      29580: inst = 32'd268468224;
      29581: inst = 32'd201348860;
      29582: inst = 32'd203459697;
      29583: inst = 32'd471859200;
      29584: inst = 32'd136314880;
      29585: inst = 32'd268468224;
      29586: inst = 32'd201348861;
      29587: inst = 32'd203455471;
      29588: inst = 32'd471859200;
      29589: inst = 32'd136314880;
      29590: inst = 32'd268468224;
      29591: inst = 32'd201348862;
      29592: inst = 32'd203455439;
      29593: inst = 32'd471859200;
      29594: inst = 32'd136314880;
      29595: inst = 32'd268468224;
      29596: inst = 32'd201348863;
      29597: inst = 32'd203459697;
      29598: inst = 32'd471859200;
      29599: inst = 32'd136314880;
      29600: inst = 32'd268468224;
      29601: inst = 32'd201348864;
      29602: inst = 32'd203459697;
      29603: inst = 32'd471859200;
      29604: inst = 32'd136314880;
      29605: inst = 32'd268468224;
      29606: inst = 32'd201348865;
      29607: inst = 32'd203459697;
      29608: inst = 32'd471859200;
      29609: inst = 32'd136314880;
      29610: inst = 32'd268468224;
      29611: inst = 32'd201348866;
      29612: inst = 32'd203459697;
      29613: inst = 32'd471859200;
      29614: inst = 32'd136314880;
      29615: inst = 32'd268468224;
      29616: inst = 32'd201348867;
      29617: inst = 32'd203459697;
      29618: inst = 32'd471859200;
      29619: inst = 32'd136314880;
      29620: inst = 32'd268468224;
      29621: inst = 32'd201348868;
      29622: inst = 32'd203459697;
      29623: inst = 32'd471859200;
      29624: inst = 32'd136314880;
      29625: inst = 32'd268468224;
      29626: inst = 32'd201348869;
      29627: inst = 32'd203459697;
      29628: inst = 32'd471859200;
      29629: inst = 32'd136314880;
      29630: inst = 32'd268468224;
      29631: inst = 32'd201348870;
      29632: inst = 32'd203459697;
      29633: inst = 32'd471859200;
      29634: inst = 32'd136314880;
      29635: inst = 32'd268468224;
      29636: inst = 32'd201348871;
      29637: inst = 32'd203459697;
      29638: inst = 32'd471859200;
      29639: inst = 32'd136314880;
      29640: inst = 32'd268468224;
      29641: inst = 32'd201348872;
      29642: inst = 32'd203459697;
      29643: inst = 32'd471859200;
      29644: inst = 32'd136314880;
      29645: inst = 32'd268468224;
      29646: inst = 32'd201348873;
      29647: inst = 32'd203459697;
      29648: inst = 32'd471859200;
      29649: inst = 32'd136314880;
      29650: inst = 32'd268468224;
      29651: inst = 32'd201348874;
      29652: inst = 32'd203459697;
      29653: inst = 32'd471859200;
      29654: inst = 32'd136314880;
      29655: inst = 32'd268468224;
      29656: inst = 32'd201348875;
      29657: inst = 32'd203459665;
      29658: inst = 32'd471859200;
      29659: inst = 32'd136314880;
      29660: inst = 32'd268468224;
      29661: inst = 32'd201348876;
      29662: inst = 32'd203451280;
      29663: inst = 32'd471859200;
      29664: inst = 32'd136314880;
      29665: inst = 32'd268468224;
      29666: inst = 32'd201348877;
      29667: inst = 32'd203451216;
      29668: inst = 32'd471859200;
      29669: inst = 32'd136314880;
      29670: inst = 32'd268468224;
      29671: inst = 32'd201348878;
      29672: inst = 32'd203451216;
      29673: inst = 32'd471859200;
      29674: inst = 32'd136314880;
      29675: inst = 32'd268468224;
      29676: inst = 32'd201348879;
      29677: inst = 32'd203451216;
      29678: inst = 32'd471859200;
      29679: inst = 32'd136314880;
      29680: inst = 32'd268468224;
      29681: inst = 32'd201348880;
      29682: inst = 32'd203451216;
      29683: inst = 32'd471859200;
      29684: inst = 32'd136314880;
      29685: inst = 32'd268468224;
      29686: inst = 32'd201348881;
      29687: inst = 32'd203451216;
      29688: inst = 32'd471859200;
      29689: inst = 32'd136314880;
      29690: inst = 32'd268468224;
      29691: inst = 32'd201348882;
      29692: inst = 32'd203451216;
      29693: inst = 32'd471859200;
      29694: inst = 32'd136314880;
      29695: inst = 32'd268468224;
      29696: inst = 32'd201348883;
      29697: inst = 32'd203451216;
      29698: inst = 32'd471859200;
      29699: inst = 32'd136314880;
      29700: inst = 32'd268468224;
      29701: inst = 32'd201348884;
      29702: inst = 32'd203451216;
      29703: inst = 32'd471859200;
      29704: inst = 32'd136314880;
      29705: inst = 32'd268468224;
      29706: inst = 32'd201348885;
      29707: inst = 32'd203451216;
      29708: inst = 32'd471859200;
      29709: inst = 32'd136314880;
      29710: inst = 32'd268468224;
      29711: inst = 32'd201348886;
      29712: inst = 32'd203451216;
      29713: inst = 32'd471859200;
      29714: inst = 32'd136314880;
      29715: inst = 32'd268468224;
      29716: inst = 32'd201348887;
      29717: inst = 32'd203451216;
      29718: inst = 32'd471859200;
      29719: inst = 32'd136314880;
      29720: inst = 32'd268468224;
      29721: inst = 32'd201348888;
      29722: inst = 32'd203451216;
      29723: inst = 32'd471859200;
      29724: inst = 32'd136314880;
      29725: inst = 32'd268468224;
      29726: inst = 32'd201348889;
      29727: inst = 32'd203451216;
      29728: inst = 32'd471859200;
      29729: inst = 32'd136314880;
      29730: inst = 32'd268468224;
      29731: inst = 32'd201348890;
      29732: inst = 32'd203451216;
      29733: inst = 32'd471859200;
      29734: inst = 32'd136314880;
      29735: inst = 32'd268468224;
      29736: inst = 32'd201348891;
      29737: inst = 32'd203451216;
      29738: inst = 32'd471859200;
      29739: inst = 32'd136314880;
      29740: inst = 32'd268468224;
      29741: inst = 32'd201348892;
      29742: inst = 32'd203451216;
      29743: inst = 32'd471859200;
      29744: inst = 32'd136314880;
      29745: inst = 32'd268468224;
      29746: inst = 32'd201348893;
      29747: inst = 32'd203451216;
      29748: inst = 32'd471859200;
      29749: inst = 32'd136314880;
      29750: inst = 32'd268468224;
      29751: inst = 32'd201348894;
      29752: inst = 32'd203451216;
      29753: inst = 32'd471859200;
      29754: inst = 32'd136314880;
      29755: inst = 32'd268468224;
      29756: inst = 32'd201348895;
      29757: inst = 32'd203451216;
      29758: inst = 32'd471859200;
      29759: inst = 32'd136314880;
      29760: inst = 32'd268468224;
      29761: inst = 32'd201348896;
      29762: inst = 32'd203451216;
      29763: inst = 32'd471859200;
      29764: inst = 32'd136314880;
      29765: inst = 32'd268468224;
      29766: inst = 32'd201348897;
      29767: inst = 32'd203451216;
      29768: inst = 32'd471859200;
      29769: inst = 32'd136314880;
      29770: inst = 32'd268468224;
      29771: inst = 32'd201348898;
      29772: inst = 32'd203451216;
      29773: inst = 32'd471859200;
      29774: inst = 32'd136314880;
      29775: inst = 32'd268468224;
      29776: inst = 32'd201348899;
      29777: inst = 32'd203451216;
      29778: inst = 32'd471859200;
      29779: inst = 32'd136314880;
      29780: inst = 32'd268468224;
      29781: inst = 32'd201348900;
      29782: inst = 32'd203451216;
      29783: inst = 32'd471859200;
      29784: inst = 32'd136314880;
      29785: inst = 32'd268468224;
      29786: inst = 32'd201348901;
      29787: inst = 32'd203451216;
      29788: inst = 32'd471859200;
      29789: inst = 32'd136314880;
      29790: inst = 32'd268468224;
      29791: inst = 32'd201348902;
      29792: inst = 32'd203451216;
      29793: inst = 32'd471859200;
      29794: inst = 32'd136314880;
      29795: inst = 32'd268468224;
      29796: inst = 32'd201348903;
      29797: inst = 32'd203451216;
      29798: inst = 32'd471859200;
      29799: inst = 32'd136314880;
      29800: inst = 32'd268468224;
      29801: inst = 32'd201348904;
      29802: inst = 32'd203451216;
      29803: inst = 32'd471859200;
      29804: inst = 32'd136314880;
      29805: inst = 32'd268468224;
      29806: inst = 32'd201348905;
      29807: inst = 32'd203451216;
      29808: inst = 32'd471859200;
      29809: inst = 32'd136314880;
      29810: inst = 32'd268468224;
      29811: inst = 32'd201348906;
      29812: inst = 32'd203451216;
      29813: inst = 32'd471859200;
      29814: inst = 32'd136314880;
      29815: inst = 32'd268468224;
      29816: inst = 32'd201348907;
      29817: inst = 32'd203451216;
      29818: inst = 32'd471859200;
      29819: inst = 32'd136314880;
      29820: inst = 32'd268468224;
      29821: inst = 32'd201348908;
      29822: inst = 32'd203451216;
      29823: inst = 32'd471859200;
      29824: inst = 32'd136314880;
      29825: inst = 32'd268468224;
      29826: inst = 32'd201348909;
      29827: inst = 32'd203451216;
      29828: inst = 32'd471859200;
      29829: inst = 32'd136314880;
      29830: inst = 32'd268468224;
      29831: inst = 32'd201348910;
      29832: inst = 32'd203451216;
      29833: inst = 32'd471859200;
      29834: inst = 32'd136314880;
      29835: inst = 32'd268468224;
      29836: inst = 32'd201348911;
      29837: inst = 32'd203451216;
      29838: inst = 32'd471859200;
      29839: inst = 32'd136314880;
      29840: inst = 32'd268468224;
      29841: inst = 32'd201348912;
      29842: inst = 32'd203451216;
      29843: inst = 32'd471859200;
      29844: inst = 32'd136314880;
      29845: inst = 32'd268468224;
      29846: inst = 32'd201348913;
      29847: inst = 32'd203451216;
      29848: inst = 32'd471859200;
      29849: inst = 32'd136314880;
      29850: inst = 32'd268468224;
      29851: inst = 32'd201348914;
      29852: inst = 32'd203451248;
      29853: inst = 32'd471859200;
      29854: inst = 32'd136314880;
      29855: inst = 32'd268468224;
      29856: inst = 32'd201348915;
      29857: inst = 32'd203457585;
      29858: inst = 32'd471859200;
      29859: inst = 32'd136314880;
      29860: inst = 32'd268468224;
      29861: inst = 32'd201348916;
      29862: inst = 32'd203459697;
      29863: inst = 32'd471859200;
      29864: inst = 32'd136314880;
      29865: inst = 32'd268468224;
      29866: inst = 32'd201348917;
      29867: inst = 32'd203459697;
      29868: inst = 32'd471859200;
      29869: inst = 32'd136314880;
      29870: inst = 32'd268468224;
      29871: inst = 32'd201348918;
      29872: inst = 32'd203459697;
      29873: inst = 32'd471859200;
      29874: inst = 32'd136314880;
      29875: inst = 32'd268468224;
      29876: inst = 32'd201348919;
      29877: inst = 32'd203459697;
      29878: inst = 32'd471859200;
      29879: inst = 32'd136314880;
      29880: inst = 32'd268468224;
      29881: inst = 32'd201348920;
      29882: inst = 32'd203459697;
      29883: inst = 32'd471859200;
      29884: inst = 32'd136314880;
      29885: inst = 32'd268468224;
      29886: inst = 32'd201348921;
      29887: inst = 32'd203459697;
      29888: inst = 32'd471859200;
      29889: inst = 32'd136314880;
      29890: inst = 32'd268468224;
      29891: inst = 32'd201348922;
      29892: inst = 32'd203459697;
      29893: inst = 32'd471859200;
      29894: inst = 32'd136314880;
      29895: inst = 32'd268468224;
      29896: inst = 32'd201348923;
      29897: inst = 32'd203459697;
      29898: inst = 32'd471859200;
      29899: inst = 32'd136314880;
      29900: inst = 32'd268468224;
      29901: inst = 32'd201348924;
      29902: inst = 32'd203459697;
      29903: inst = 32'd471859200;
      29904: inst = 32'd136314880;
      29905: inst = 32'd268468224;
      29906: inst = 32'd201348925;
      29907: inst = 32'd203459697;
      29908: inst = 32'd471859200;
      29909: inst = 32'd136314880;
      29910: inst = 32'd268468224;
      29911: inst = 32'd201348926;
      29912: inst = 32'd203459697;
      29913: inst = 32'd471859200;
      29914: inst = 32'd136314880;
      29915: inst = 32'd268468224;
      29916: inst = 32'd201348927;
      29917: inst = 32'd203459697;
      29918: inst = 32'd471859200;
      29919: inst = 32'd136314880;
      29920: inst = 32'd268468224;
      29921: inst = 32'd201348928;
      29922: inst = 32'd203459697;
      29923: inst = 32'd471859200;
      29924: inst = 32'd136314880;
      29925: inst = 32'd268468224;
      29926: inst = 32'd201348929;
      29927: inst = 32'd203457552;
      29928: inst = 32'd471859200;
      29929: inst = 32'd136314880;
      29930: inst = 32'd268468224;
      29931: inst = 32'd201348930;
      29932: inst = 32'd203459697;
      29933: inst = 32'd471859200;
      29934: inst = 32'd136314880;
      29935: inst = 32'd268468224;
      29936: inst = 32'd201348931;
      29937: inst = 32'd203459697;
      29938: inst = 32'd471859200;
      29939: inst = 32'd136314880;
      29940: inst = 32'd268468224;
      29941: inst = 32'd201348932;
      29942: inst = 32'd203459697;
      29943: inst = 32'd471859200;
      29944: inst = 32'd136314880;
      29945: inst = 32'd268468224;
      29946: inst = 32'd201348933;
      29947: inst = 32'd203459697;
      29948: inst = 32'd471859200;
      29949: inst = 32'd136314880;
      29950: inst = 32'd268468224;
      29951: inst = 32'd201348934;
      29952: inst = 32'd203459697;
      29953: inst = 32'd471859200;
      29954: inst = 32'd136314880;
      29955: inst = 32'd268468224;
      29956: inst = 32'd201348935;
      29957: inst = 32'd203449133;
      29958: inst = 32'd471859200;
      29959: inst = 32'd136314880;
      29960: inst = 32'd268468224;
      29961: inst = 32'd201348936;
      29962: inst = 32'd203444874;
      29963: inst = 32'd471859200;
      29964: inst = 32'd136314880;
      29965: inst = 32'd268468224;
      29966: inst = 32'd201348937;
      29967: inst = 32'd203444874;
      29968: inst = 32'd471859200;
      29969: inst = 32'd136314880;
      29970: inst = 32'd268468224;
      29971: inst = 32'd201348938;
      29972: inst = 32'd203451216;
      29973: inst = 32'd471859200;
      29974: inst = 32'd136314880;
      29975: inst = 32'd268468224;
      29976: inst = 32'd201348939;
      29977: inst = 32'd203451216;
      29978: inst = 32'd471859200;
      29979: inst = 32'd136314880;
      29980: inst = 32'd268468224;
      29981: inst = 32'd201348940;
      29982: inst = 32'd203451216;
      29983: inst = 32'd471859200;
      29984: inst = 32'd136314880;
      29985: inst = 32'd268468224;
      29986: inst = 32'd201348941;
      29987: inst = 32'd203451216;
      29988: inst = 32'd471859200;
      29989: inst = 32'd136314880;
      29990: inst = 32'd268468224;
      29991: inst = 32'd201348942;
      29992: inst = 32'd203451216;
      29993: inst = 32'd471859200;
      29994: inst = 32'd136314880;
      29995: inst = 32'd268468224;
      29996: inst = 32'd201348943;
      29997: inst = 32'd203451216;
      29998: inst = 32'd471859200;
      29999: inst = 32'd136314880;
      30000: inst = 32'd268468224;
      30001: inst = 32'd201348944;
      30002: inst = 32'd203451216;
      30003: inst = 32'd471859200;
      30004: inst = 32'd136314880;
      30005: inst = 32'd268468224;
      30006: inst = 32'd201348945;
      30007: inst = 32'd203451216;
      30008: inst = 32'd471859200;
      30009: inst = 32'd136314880;
      30010: inst = 32'd268468224;
      30011: inst = 32'd201348946;
      30012: inst = 32'd203451216;
      30013: inst = 32'd471859200;
      30014: inst = 32'd136314880;
      30015: inst = 32'd268468224;
      30016: inst = 32'd201348947;
      30017: inst = 32'd203451216;
      30018: inst = 32'd471859200;
      30019: inst = 32'd136314880;
      30020: inst = 32'd268468224;
      30021: inst = 32'd201348948;
      30022: inst = 32'd203451216;
      30023: inst = 32'd471859200;
      30024: inst = 32'd136314880;
      30025: inst = 32'd268468224;
      30026: inst = 32'd201348949;
      30027: inst = 32'd203451216;
      30028: inst = 32'd471859200;
      30029: inst = 32'd136314880;
      30030: inst = 32'd268468224;
      30031: inst = 32'd201348950;
      30032: inst = 32'd203444874;
      30033: inst = 32'd471859200;
      30034: inst = 32'd136314880;
      30035: inst = 32'd268468224;
      30036: inst = 32'd201348951;
      30037: inst = 32'd203444874;
      30038: inst = 32'd471859200;
      30039: inst = 32'd136314880;
      30040: inst = 32'd268468224;
      30041: inst = 32'd201348952;
      30042: inst = 32'd203449133;
      30043: inst = 32'd471859200;
      30044: inst = 32'd136314880;
      30045: inst = 32'd268468224;
      30046: inst = 32'd201348953;
      30047: inst = 32'd203459697;
      30048: inst = 32'd471859200;
      30049: inst = 32'd136314880;
      30050: inst = 32'd268468224;
      30051: inst = 32'd201348954;
      30052: inst = 32'd203459697;
      30053: inst = 32'd471859200;
      30054: inst = 32'd136314880;
      30055: inst = 32'd268468224;
      30056: inst = 32'd201348955;
      30057: inst = 32'd203459697;
      30058: inst = 32'd471859200;
      30059: inst = 32'd136314880;
      30060: inst = 32'd268468224;
      30061: inst = 32'd201348956;
      30062: inst = 32'd203459697;
      30063: inst = 32'd471859200;
      30064: inst = 32'd136314880;
      30065: inst = 32'd268468224;
      30066: inst = 32'd201348957;
      30067: inst = 32'd203459697;
      30068: inst = 32'd471859200;
      30069: inst = 32'd136314880;
      30070: inst = 32'd268468224;
      30071: inst = 32'd201348958;
      30072: inst = 32'd203457552;
      30073: inst = 32'd471859200;
      30074: inst = 32'd136314880;
      30075: inst = 32'd268468224;
      30076: inst = 32'd201348959;
      30077: inst = 32'd203459697;
      30078: inst = 32'd471859200;
      30079: inst = 32'd136314880;
      30080: inst = 32'd268468224;
      30081: inst = 32'd201348960;
      30082: inst = 32'd203459697;
      30083: inst = 32'd471859200;
      30084: inst = 32'd136314880;
      30085: inst = 32'd268468224;
      30086: inst = 32'd201348961;
      30087: inst = 32'd203459697;
      30088: inst = 32'd471859200;
      30089: inst = 32'd136314880;
      30090: inst = 32'd268468224;
      30091: inst = 32'd201348962;
      30092: inst = 32'd203459697;
      30093: inst = 32'd471859200;
      30094: inst = 32'd136314880;
      30095: inst = 32'd268468224;
      30096: inst = 32'd201348963;
      30097: inst = 32'd203459697;
      30098: inst = 32'd471859200;
      30099: inst = 32'd136314880;
      30100: inst = 32'd268468224;
      30101: inst = 32'd201348964;
      30102: inst = 32'd203459697;
      30103: inst = 32'd471859200;
      30104: inst = 32'd136314880;
      30105: inst = 32'd268468224;
      30106: inst = 32'd201348965;
      30107: inst = 32'd203459697;
      30108: inst = 32'd471859200;
      30109: inst = 32'd136314880;
      30110: inst = 32'd268468224;
      30111: inst = 32'd201348966;
      30112: inst = 32'd203459697;
      30113: inst = 32'd471859200;
      30114: inst = 32'd136314880;
      30115: inst = 32'd268468224;
      30116: inst = 32'd201348967;
      30117: inst = 32'd203459697;
      30118: inst = 32'd471859200;
      30119: inst = 32'd136314880;
      30120: inst = 32'd268468224;
      30121: inst = 32'd201348968;
      30122: inst = 32'd203459697;
      30123: inst = 32'd471859200;
      30124: inst = 32'd136314880;
      30125: inst = 32'd268468224;
      30126: inst = 32'd201348969;
      30127: inst = 32'd203459697;
      30128: inst = 32'd471859200;
      30129: inst = 32'd136314880;
      30130: inst = 32'd268468224;
      30131: inst = 32'd201348970;
      30132: inst = 32'd203459697;
      30133: inst = 32'd471859200;
      30134: inst = 32'd136314880;
      30135: inst = 32'd268468224;
      30136: inst = 32'd201348971;
      30137: inst = 32'd203459697;
      30138: inst = 32'd471859200;
      30139: inst = 32'd136314880;
      30140: inst = 32'd268468224;
      30141: inst = 32'd201348972;
      30142: inst = 32'd203457585;
      30143: inst = 32'd471859200;
      30144: inst = 32'd136314880;
      30145: inst = 32'd268468224;
      30146: inst = 32'd201348973;
      30147: inst = 32'd203451248;
      30148: inst = 32'd471859200;
      30149: inst = 32'd136314880;
      30150: inst = 32'd268468224;
      30151: inst = 32'd201348974;
      30152: inst = 32'd203451216;
      30153: inst = 32'd471859200;
      30154: inst = 32'd136314880;
      30155: inst = 32'd268468224;
      30156: inst = 32'd201348975;
      30157: inst = 32'd203451216;
      30158: inst = 32'd471859200;
      30159: inst = 32'd136314880;
      30160: inst = 32'd268468224;
      30161: inst = 32'd201348976;
      30162: inst = 32'd203451216;
      30163: inst = 32'd471859200;
      30164: inst = 32'd136314880;
      30165: inst = 32'd268468224;
      30166: inst = 32'd201348977;
      30167: inst = 32'd203451216;
      30168: inst = 32'd471859200;
      30169: inst = 32'd136314880;
      30170: inst = 32'd268468224;
      30171: inst = 32'd201348978;
      30172: inst = 32'd203451216;
      30173: inst = 32'd471859200;
      30174: inst = 32'd136314880;
      30175: inst = 32'd268468224;
      30176: inst = 32'd201348979;
      30177: inst = 32'd203451216;
      30178: inst = 32'd471859200;
      30179: inst = 32'd136314880;
      30180: inst = 32'd268468224;
      30181: inst = 32'd201348980;
      30182: inst = 32'd203451216;
      30183: inst = 32'd471859200;
      30184: inst = 32'd136314880;
      30185: inst = 32'd268468224;
      30186: inst = 32'd201348981;
      30187: inst = 32'd203451216;
      30188: inst = 32'd471859200;
      30189: inst = 32'd136314880;
      30190: inst = 32'd268468224;
      30191: inst = 32'd201348982;
      30192: inst = 32'd203451216;
      30193: inst = 32'd471859200;
      30194: inst = 32'd136314880;
      30195: inst = 32'd268468224;
      30196: inst = 32'd201348983;
      30197: inst = 32'd203451216;
      30198: inst = 32'd471859200;
      30199: inst = 32'd136314880;
      30200: inst = 32'd268468224;
      30201: inst = 32'd201348984;
      30202: inst = 32'd203451216;
      30203: inst = 32'd471859200;
      30204: inst = 32'd136314880;
      30205: inst = 32'd268468224;
      30206: inst = 32'd201348985;
      30207: inst = 32'd203451216;
      30208: inst = 32'd471859200;
      30209: inst = 32'd136314880;
      30210: inst = 32'd268468224;
      30211: inst = 32'd201348986;
      30212: inst = 32'd203451216;
      30213: inst = 32'd471859200;
      30214: inst = 32'd136314880;
      30215: inst = 32'd268468224;
      30216: inst = 32'd201348987;
      30217: inst = 32'd203451216;
      30218: inst = 32'd471859200;
      30219: inst = 32'd136314880;
      30220: inst = 32'd268468224;
      30221: inst = 32'd201348988;
      30222: inst = 32'd203451216;
      30223: inst = 32'd471859200;
      30224: inst = 32'd136314880;
      30225: inst = 32'd268468224;
      30226: inst = 32'd201348989;
      30227: inst = 32'd203451216;
      30228: inst = 32'd471859200;
      30229: inst = 32'd136314880;
      30230: inst = 32'd268468224;
      30231: inst = 32'd201348990;
      30232: inst = 32'd203451216;
      30233: inst = 32'd471859200;
      30234: inst = 32'd136314880;
      30235: inst = 32'd268468224;
      30236: inst = 32'd201348991;
      30237: inst = 32'd203451216;
      30238: inst = 32'd471859200;
      30239: inst = 32'd136314880;
      30240: inst = 32'd268468224;
      30241: inst = 32'd201348992;
      30242: inst = 32'd203451216;
      30243: inst = 32'd471859200;
      30244: inst = 32'd136314880;
      30245: inst = 32'd268468224;
      30246: inst = 32'd201348993;
      30247: inst = 32'd203451216;
      30248: inst = 32'd471859200;
      30249: inst = 32'd136314880;
      30250: inst = 32'd268468224;
      30251: inst = 32'd201348994;
      30252: inst = 32'd203451216;
      30253: inst = 32'd471859200;
      30254: inst = 32'd136314880;
      30255: inst = 32'd268468224;
      30256: inst = 32'd201348995;
      30257: inst = 32'd203451216;
      30258: inst = 32'd471859200;
      30259: inst = 32'd136314880;
      30260: inst = 32'd268468224;
      30261: inst = 32'd201348996;
      30262: inst = 32'd203451216;
      30263: inst = 32'd471859200;
      30264: inst = 32'd136314880;
      30265: inst = 32'd268468224;
      30266: inst = 32'd201348997;
      30267: inst = 32'd203451216;
      30268: inst = 32'd471859200;
      30269: inst = 32'd136314880;
      30270: inst = 32'd268468224;
      30271: inst = 32'd201348998;
      30272: inst = 32'd203451216;
      30273: inst = 32'd471859200;
      30274: inst = 32'd136314880;
      30275: inst = 32'd268468224;
      30276: inst = 32'd201348999;
      30277: inst = 32'd203451216;
      30278: inst = 32'd471859200;
      30279: inst = 32'd136314880;
      30280: inst = 32'd268468224;
      30281: inst = 32'd201349000;
      30282: inst = 32'd203451216;
      30283: inst = 32'd471859200;
      30284: inst = 32'd136314880;
      30285: inst = 32'd268468224;
      30286: inst = 32'd201349001;
      30287: inst = 32'd203451216;
      30288: inst = 32'd471859200;
      30289: inst = 32'd136314880;
      30290: inst = 32'd268468224;
      30291: inst = 32'd201349002;
      30292: inst = 32'd203451216;
      30293: inst = 32'd471859200;
      30294: inst = 32'd136314880;
      30295: inst = 32'd268468224;
      30296: inst = 32'd201349003;
      30297: inst = 32'd203451216;
      30298: inst = 32'd471859200;
      30299: inst = 32'd136314880;
      30300: inst = 32'd268468224;
      30301: inst = 32'd201349004;
      30302: inst = 32'd203451216;
      30303: inst = 32'd471859200;
      30304: inst = 32'd136314880;
      30305: inst = 32'd268468224;
      30306: inst = 32'd201349005;
      30307: inst = 32'd203451216;
      30308: inst = 32'd471859200;
      30309: inst = 32'd136314880;
      30310: inst = 32'd268468224;
      30311: inst = 32'd201349006;
      30312: inst = 32'd203451216;
      30313: inst = 32'd471859200;
      30314: inst = 32'd136314880;
      30315: inst = 32'd268468224;
      30316: inst = 32'd201349007;
      30317: inst = 32'd203451216;
      30318: inst = 32'd471859200;
      30319: inst = 32'd136314880;
      30320: inst = 32'd268468224;
      30321: inst = 32'd201349008;
      30322: inst = 32'd203451216;
      30323: inst = 32'd471859200;
      30324: inst = 32'd136314880;
      30325: inst = 32'd268468224;
      30326: inst = 32'd201349009;
      30327: inst = 32'd203451216;
      30328: inst = 32'd471859200;
      30329: inst = 32'd136314880;
      30330: inst = 32'd268468224;
      30331: inst = 32'd201349010;
      30332: inst = 32'd203455505;
      30333: inst = 32'd471859200;
      30334: inst = 32'd136314880;
      30335: inst = 32'd268468224;
      30336: inst = 32'd201349011;
      30337: inst = 32'd203459697;
      30338: inst = 32'd471859200;
      30339: inst = 32'd136314880;
      30340: inst = 32'd268468224;
      30341: inst = 32'd201349012;
      30342: inst = 32'd203459697;
      30343: inst = 32'd471859200;
      30344: inst = 32'd136314880;
      30345: inst = 32'd268468224;
      30346: inst = 32'd201349013;
      30347: inst = 32'd203459697;
      30348: inst = 32'd471859200;
      30349: inst = 32'd136314880;
      30350: inst = 32'd268468224;
      30351: inst = 32'd201349014;
      30352: inst = 32'd203459697;
      30353: inst = 32'd471859200;
      30354: inst = 32'd136314880;
      30355: inst = 32'd268468224;
      30356: inst = 32'd201349015;
      30357: inst = 32'd203459697;
      30358: inst = 32'd471859200;
      30359: inst = 32'd136314880;
      30360: inst = 32'd268468224;
      30361: inst = 32'd201349016;
      30362: inst = 32'd203459697;
      30363: inst = 32'd471859200;
      30364: inst = 32'd136314880;
      30365: inst = 32'd268468224;
      30366: inst = 32'd201349017;
      30367: inst = 32'd203459697;
      30368: inst = 32'd471859200;
      30369: inst = 32'd136314880;
      30370: inst = 32'd268468224;
      30371: inst = 32'd201349018;
      30372: inst = 32'd203459697;
      30373: inst = 32'd471859200;
      30374: inst = 32'd136314880;
      30375: inst = 32'd268468224;
      30376: inst = 32'd201349019;
      30377: inst = 32'd203459697;
      30378: inst = 32'd471859200;
      30379: inst = 32'd136314880;
      30380: inst = 32'd268468224;
      30381: inst = 32'd201349020;
      30382: inst = 32'd203459697;
      30383: inst = 32'd471859200;
      30384: inst = 32'd136314880;
      30385: inst = 32'd268468224;
      30386: inst = 32'd201349021;
      30387: inst = 32'd203459697;
      30388: inst = 32'd471859200;
      30389: inst = 32'd136314880;
      30390: inst = 32'd268468224;
      30391: inst = 32'd201349022;
      30392: inst = 32'd203459697;
      30393: inst = 32'd471859200;
      30394: inst = 32'd136314880;
      30395: inst = 32'd268468224;
      30396: inst = 32'd201349023;
      30397: inst = 32'd203459697;
      30398: inst = 32'd471859200;
      30399: inst = 32'd136314880;
      30400: inst = 32'd268468224;
      30401: inst = 32'd201349024;
      30402: inst = 32'd203459697;
      30403: inst = 32'd471859200;
      30404: inst = 32'd136314880;
      30405: inst = 32'd268468224;
      30406: inst = 32'd201349025;
      30407: inst = 32'd203459697;
      30408: inst = 32'd471859200;
      30409: inst = 32'd136314880;
      30410: inst = 32'd268468224;
      30411: inst = 32'd201349026;
      30412: inst = 32'd203459697;
      30413: inst = 32'd471859200;
      30414: inst = 32'd136314880;
      30415: inst = 32'd268468224;
      30416: inst = 32'd201349027;
      30417: inst = 32'd203459697;
      30418: inst = 32'd471859200;
      30419: inst = 32'd136314880;
      30420: inst = 32'd268468224;
      30421: inst = 32'd201349028;
      30422: inst = 32'd203459697;
      30423: inst = 32'd471859200;
      30424: inst = 32'd136314880;
      30425: inst = 32'd268468224;
      30426: inst = 32'd201349029;
      30427: inst = 32'd203459697;
      30428: inst = 32'd471859200;
      30429: inst = 32'd136314880;
      30430: inst = 32'd268468224;
      30431: inst = 32'd201349030;
      30432: inst = 32'd203459697;
      30433: inst = 32'd471859200;
      30434: inst = 32'd136314880;
      30435: inst = 32'd268468224;
      30436: inst = 32'd201349031;
      30437: inst = 32'd203447020;
      30438: inst = 32'd471859200;
      30439: inst = 32'd136314880;
      30440: inst = 32'd268468224;
      30441: inst = 32'd201349032;
      30442: inst = 32'd203444874;
      30443: inst = 32'd471859200;
      30444: inst = 32'd136314880;
      30445: inst = 32'd268468224;
      30446: inst = 32'd201349033;
      30447: inst = 32'd203444874;
      30448: inst = 32'd471859200;
      30449: inst = 32'd136314880;
      30450: inst = 32'd268468224;
      30451: inst = 32'd201349034;
      30452: inst = 32'd203451216;
      30453: inst = 32'd471859200;
      30454: inst = 32'd136314880;
      30455: inst = 32'd268468224;
      30456: inst = 32'd201349035;
      30457: inst = 32'd203451216;
      30458: inst = 32'd471859200;
      30459: inst = 32'd136314880;
      30460: inst = 32'd268468224;
      30461: inst = 32'd201349036;
      30462: inst = 32'd203451216;
      30463: inst = 32'd471859200;
      30464: inst = 32'd136314880;
      30465: inst = 32'd268468224;
      30466: inst = 32'd201349037;
      30467: inst = 32'd203451216;
      30468: inst = 32'd471859200;
      30469: inst = 32'd136314880;
      30470: inst = 32'd268468224;
      30471: inst = 32'd201349038;
      30472: inst = 32'd203451216;
      30473: inst = 32'd471859200;
      30474: inst = 32'd136314880;
      30475: inst = 32'd268468224;
      30476: inst = 32'd201349039;
      30477: inst = 32'd203451216;
      30478: inst = 32'd471859200;
      30479: inst = 32'd136314880;
      30480: inst = 32'd268468224;
      30481: inst = 32'd201349040;
      30482: inst = 32'd203451216;
      30483: inst = 32'd471859200;
      30484: inst = 32'd136314880;
      30485: inst = 32'd268468224;
      30486: inst = 32'd201349041;
      30487: inst = 32'd203451216;
      30488: inst = 32'd471859200;
      30489: inst = 32'd136314880;
      30490: inst = 32'd268468224;
      30491: inst = 32'd201349042;
      30492: inst = 32'd203451216;
      30493: inst = 32'd471859200;
      30494: inst = 32'd136314880;
      30495: inst = 32'd268468224;
      30496: inst = 32'd201349043;
      30497: inst = 32'd203451216;
      30498: inst = 32'd471859200;
      30499: inst = 32'd136314880;
      30500: inst = 32'd268468224;
      30501: inst = 32'd201349044;
      30502: inst = 32'd203451216;
      30503: inst = 32'd471859200;
      30504: inst = 32'd136314880;
      30505: inst = 32'd268468224;
      30506: inst = 32'd201349045;
      30507: inst = 32'd203451216;
      30508: inst = 32'd471859200;
      30509: inst = 32'd136314880;
      30510: inst = 32'd268468224;
      30511: inst = 32'd201349046;
      30512: inst = 32'd203444874;
      30513: inst = 32'd471859200;
      30514: inst = 32'd136314880;
      30515: inst = 32'd268468224;
      30516: inst = 32'd201349047;
      30517: inst = 32'd203444874;
      30518: inst = 32'd471859200;
      30519: inst = 32'd136314880;
      30520: inst = 32'd268468224;
      30521: inst = 32'd201349048;
      30522: inst = 32'd203447020;
      30523: inst = 32'd471859200;
      30524: inst = 32'd136314880;
      30525: inst = 32'd268468224;
      30526: inst = 32'd201349049;
      30527: inst = 32'd203459697;
      30528: inst = 32'd471859200;
      30529: inst = 32'd136314880;
      30530: inst = 32'd268468224;
      30531: inst = 32'd201349050;
      30532: inst = 32'd203459697;
      30533: inst = 32'd471859200;
      30534: inst = 32'd136314880;
      30535: inst = 32'd268468224;
      30536: inst = 32'd201349051;
      30537: inst = 32'd203459697;
      30538: inst = 32'd471859200;
      30539: inst = 32'd136314880;
      30540: inst = 32'd268468224;
      30541: inst = 32'd201349052;
      30542: inst = 32'd203459697;
      30543: inst = 32'd471859200;
      30544: inst = 32'd136314880;
      30545: inst = 32'd268468224;
      30546: inst = 32'd201349053;
      30547: inst = 32'd203459697;
      30548: inst = 32'd471859200;
      30549: inst = 32'd136314880;
      30550: inst = 32'd268468224;
      30551: inst = 32'd201349054;
      30552: inst = 32'd203459697;
      30553: inst = 32'd471859200;
      30554: inst = 32'd136314880;
      30555: inst = 32'd268468224;
      30556: inst = 32'd201349055;
      30557: inst = 32'd203459697;
      30558: inst = 32'd471859200;
      30559: inst = 32'd136314880;
      30560: inst = 32'd268468224;
      30561: inst = 32'd201349056;
      30562: inst = 32'd203459697;
      30563: inst = 32'd471859200;
      30564: inst = 32'd136314880;
      30565: inst = 32'd268468224;
      30566: inst = 32'd201349057;
      30567: inst = 32'd203459697;
      30568: inst = 32'd471859200;
      30569: inst = 32'd136314880;
      30570: inst = 32'd268468224;
      30571: inst = 32'd201349058;
      30572: inst = 32'd203459697;
      30573: inst = 32'd471859200;
      30574: inst = 32'd136314880;
      30575: inst = 32'd268468224;
      30576: inst = 32'd201349059;
      30577: inst = 32'd203459697;
      30578: inst = 32'd471859200;
      30579: inst = 32'd136314880;
      30580: inst = 32'd268468224;
      30581: inst = 32'd201349060;
      30582: inst = 32'd203459697;
      30583: inst = 32'd471859200;
      30584: inst = 32'd136314880;
      30585: inst = 32'd268468224;
      30586: inst = 32'd201349061;
      30587: inst = 32'd203459697;
      30588: inst = 32'd471859200;
      30589: inst = 32'd136314880;
      30590: inst = 32'd268468224;
      30591: inst = 32'd201349062;
      30592: inst = 32'd203459697;
      30593: inst = 32'd471859200;
      30594: inst = 32'd136314880;
      30595: inst = 32'd268468224;
      30596: inst = 32'd201349063;
      30597: inst = 32'd203459697;
      30598: inst = 32'd471859200;
      30599: inst = 32'd136314880;
      30600: inst = 32'd268468224;
      30601: inst = 32'd201349064;
      30602: inst = 32'd203459697;
      30603: inst = 32'd471859200;
      30604: inst = 32'd136314880;
      30605: inst = 32'd268468224;
      30606: inst = 32'd201349065;
      30607: inst = 32'd203459697;
      30608: inst = 32'd471859200;
      30609: inst = 32'd136314880;
      30610: inst = 32'd268468224;
      30611: inst = 32'd201349066;
      30612: inst = 32'd203459697;
      30613: inst = 32'd471859200;
      30614: inst = 32'd136314880;
      30615: inst = 32'd268468224;
      30616: inst = 32'd201349067;
      30617: inst = 32'd203459697;
      30618: inst = 32'd471859200;
      30619: inst = 32'd136314880;
      30620: inst = 32'd268468224;
      30621: inst = 32'd201349068;
      30622: inst = 32'd203459697;
      30623: inst = 32'd471859200;
      30624: inst = 32'd136314880;
      30625: inst = 32'd268468224;
      30626: inst = 32'd201349069;
      30627: inst = 32'd203455505;
      30628: inst = 32'd471859200;
      30629: inst = 32'd136314880;
      30630: inst = 32'd268468224;
      30631: inst = 32'd201349070;
      30632: inst = 32'd203451216;
      30633: inst = 32'd471859200;
      30634: inst = 32'd136314880;
      30635: inst = 32'd268468224;
      30636: inst = 32'd201349071;
      30637: inst = 32'd203451216;
      30638: inst = 32'd471859200;
      30639: inst = 32'd136314880;
      30640: inst = 32'd268468224;
      30641: inst = 32'd201349072;
      30642: inst = 32'd203451216;
      30643: inst = 32'd471859200;
      30644: inst = 32'd136314880;
      30645: inst = 32'd268468224;
      30646: inst = 32'd201349073;
      30647: inst = 32'd203451216;
      30648: inst = 32'd471859200;
      30649: inst = 32'd136314880;
      30650: inst = 32'd268468224;
      30651: inst = 32'd201349074;
      30652: inst = 32'd203451216;
      30653: inst = 32'd471859200;
      30654: inst = 32'd136314880;
      30655: inst = 32'd268468224;
      30656: inst = 32'd201349075;
      30657: inst = 32'd203451216;
      30658: inst = 32'd471859200;
      30659: inst = 32'd136314880;
      30660: inst = 32'd268468224;
      30661: inst = 32'd201349076;
      30662: inst = 32'd203451216;
      30663: inst = 32'd471859200;
      30664: inst = 32'd136314880;
      30665: inst = 32'd268468224;
      30666: inst = 32'd201349077;
      30667: inst = 32'd203451216;
      30668: inst = 32'd471859200;
      30669: inst = 32'd136314880;
      30670: inst = 32'd268468224;
      30671: inst = 32'd201349078;
      30672: inst = 32'd203451216;
      30673: inst = 32'd471859200;
      30674: inst = 32'd136314880;
      30675: inst = 32'd268468224;
      30676: inst = 32'd201349079;
      30677: inst = 32'd203451216;
      30678: inst = 32'd471859200;
      30679: inst = 32'd136314880;
      30680: inst = 32'd268468224;
      30681: inst = 32'd201349080;
      30682: inst = 32'd203451216;
      30683: inst = 32'd471859200;
      30684: inst = 32'd136314880;
      30685: inst = 32'd268468224;
      30686: inst = 32'd201349081;
      30687: inst = 32'd203451216;
      30688: inst = 32'd471859200;
      30689: inst = 32'd136314880;
      30690: inst = 32'd268468224;
      30691: inst = 32'd201349082;
      30692: inst = 32'd203451216;
      30693: inst = 32'd471859200;
      30694: inst = 32'd136314880;
      30695: inst = 32'd268468224;
      30696: inst = 32'd201349083;
      30697: inst = 32'd203451216;
      30698: inst = 32'd471859200;
      30699: inst = 32'd136314880;
      30700: inst = 32'd268468224;
      30701: inst = 32'd201349084;
      30702: inst = 32'd203451216;
      30703: inst = 32'd471859200;
      30704: inst = 32'd136314880;
      30705: inst = 32'd268468224;
      30706: inst = 32'd201349085;
      30707: inst = 32'd203451216;
      30708: inst = 32'd471859200;
      30709: inst = 32'd136314880;
      30710: inst = 32'd268468224;
      30711: inst = 32'd201349086;
      30712: inst = 32'd203451216;
      30713: inst = 32'd471859200;
      30714: inst = 32'd136314880;
      30715: inst = 32'd268468224;
      30716: inst = 32'd201349087;
      30717: inst = 32'd203451216;
      30718: inst = 32'd471859200;
      30719: inst = 32'd136314880;
      30720: inst = 32'd272629792;
      30721: inst = 32'd205520896;
      30722: inst = 32'd809631745;
      30723: inst = 32'd333447168;
      30724: inst = 32'd266369026;
      30725: inst = 32'd473956352;
      30726: inst = 32'd1541406720;
      30727: inst = 32'd268468224;
      30728: inst = 32'd201342944;
      30729: inst = 32'd203423744;
      30730: inst = 32'd471859200;
      30731: inst = 32'd136314880;
      30732: inst = 32'd268468224;
      30733: inst = 32'd201342945;
      30734: inst = 32'd203423744;
      30735: inst = 32'd471859200;
      30736: inst = 32'd136314880;
      30737: inst = 32'd268468224;
      30738: inst = 32'd201342946;
      30739: inst = 32'd203423744;
      30740: inst = 32'd471859200;
      30741: inst = 32'd136314880;
      30742: inst = 32'd268468224;
      30743: inst = 32'd201342947;
      30744: inst = 32'd203423744;
      30745: inst = 32'd471859200;
      30746: inst = 32'd136314880;
      30747: inst = 32'd268468224;
      30748: inst = 32'd201342948;
      30749: inst = 32'd203423744;
      30750: inst = 32'd471859200;
      30751: inst = 32'd136314880;
      30752: inst = 32'd268468224;
      30753: inst = 32'd201342949;
      30754: inst = 32'd203423744;
      30755: inst = 32'd471859200;
      30756: inst = 32'd136314880;
      30757: inst = 32'd268468224;
      30758: inst = 32'd201342950;
      30759: inst = 32'd203423744;
      30760: inst = 32'd471859200;
      30761: inst = 32'd136314880;
      30762: inst = 32'd268468224;
      30763: inst = 32'd201342951;
      30764: inst = 32'd203423744;
      30765: inst = 32'd471859200;
      30766: inst = 32'd136314880;
      30767: inst = 32'd268468224;
      30768: inst = 32'd201342952;
      30769: inst = 32'd203423744;
      30770: inst = 32'd471859200;
      30771: inst = 32'd136314880;
      30772: inst = 32'd268468224;
      30773: inst = 32'd201342953;
      30774: inst = 32'd203423744;
      30775: inst = 32'd471859200;
      30776: inst = 32'd136314880;
      30777: inst = 32'd268468224;
      30778: inst = 32'd201342954;
      30779: inst = 32'd203423744;
      30780: inst = 32'd471859200;
      30781: inst = 32'd136314880;
      30782: inst = 32'd268468224;
      30783: inst = 32'd201342955;
      30784: inst = 32'd203423744;
      30785: inst = 32'd471859200;
      30786: inst = 32'd136314880;
      30787: inst = 32'd268468224;
      30788: inst = 32'd201342956;
      30789: inst = 32'd203423744;
      30790: inst = 32'd471859200;
      30791: inst = 32'd136314880;
      30792: inst = 32'd268468224;
      30793: inst = 32'd201342957;
      30794: inst = 32'd203423744;
      30795: inst = 32'd471859200;
      30796: inst = 32'd136314880;
      30797: inst = 32'd268468224;
      30798: inst = 32'd201342958;
      30799: inst = 32'd203423744;
      30800: inst = 32'd471859200;
      30801: inst = 32'd136314880;
      30802: inst = 32'd268468224;
      30803: inst = 32'd201342959;
      30804: inst = 32'd203423744;
      30805: inst = 32'd471859200;
      30806: inst = 32'd136314880;
      30807: inst = 32'd268468224;
      30808: inst = 32'd201342960;
      30809: inst = 32'd203423744;
      30810: inst = 32'd471859200;
      30811: inst = 32'd136314880;
      30812: inst = 32'd268468224;
      30813: inst = 32'd201342961;
      30814: inst = 32'd203423744;
      30815: inst = 32'd471859200;
      30816: inst = 32'd136314880;
      30817: inst = 32'd268468224;
      30818: inst = 32'd201342962;
      30819: inst = 32'd203423744;
      30820: inst = 32'd471859200;
      30821: inst = 32'd136314880;
      30822: inst = 32'd268468224;
      30823: inst = 32'd201342963;
      30824: inst = 32'd203423744;
      30825: inst = 32'd471859200;
      30826: inst = 32'd136314880;
      30827: inst = 32'd268468224;
      30828: inst = 32'd201342964;
      30829: inst = 32'd203423744;
      30830: inst = 32'd471859200;
      30831: inst = 32'd136314880;
      30832: inst = 32'd268468224;
      30833: inst = 32'd201342965;
      30834: inst = 32'd203423744;
      30835: inst = 32'd471859200;
      30836: inst = 32'd136314880;
      30837: inst = 32'd268468224;
      30838: inst = 32'd201342966;
      30839: inst = 32'd203423744;
      30840: inst = 32'd471859200;
      30841: inst = 32'd136314880;
      30842: inst = 32'd268468224;
      30843: inst = 32'd201342967;
      30844: inst = 32'd203423744;
      30845: inst = 32'd471859200;
      30846: inst = 32'd136314880;
      30847: inst = 32'd268468224;
      30848: inst = 32'd201342968;
      30849: inst = 32'd203423744;
      30850: inst = 32'd471859200;
      30851: inst = 32'd136314880;
      30852: inst = 32'd268468224;
      30853: inst = 32'd201342969;
      30854: inst = 32'd203423744;
      30855: inst = 32'd471859200;
      30856: inst = 32'd136314880;
      30857: inst = 32'd268468224;
      30858: inst = 32'd201342970;
      30859: inst = 32'd203423744;
      30860: inst = 32'd471859200;
      30861: inst = 32'd136314880;
      30862: inst = 32'd268468224;
      30863: inst = 32'd201342971;
      30864: inst = 32'd203423744;
      30865: inst = 32'd471859200;
      30866: inst = 32'd136314880;
      30867: inst = 32'd268468224;
      30868: inst = 32'd201342972;
      30869: inst = 32'd203423744;
      30870: inst = 32'd471859200;
      30871: inst = 32'd136314880;
      30872: inst = 32'd268468224;
      30873: inst = 32'd201342973;
      30874: inst = 32'd203423744;
      30875: inst = 32'd471859200;
      30876: inst = 32'd136314880;
      30877: inst = 32'd268468224;
      30878: inst = 32'd201342974;
      30879: inst = 32'd203423744;
      30880: inst = 32'd471859200;
      30881: inst = 32'd136314880;
      30882: inst = 32'd268468224;
      30883: inst = 32'd201342975;
      30884: inst = 32'd203423744;
      30885: inst = 32'd471859200;
      30886: inst = 32'd136314880;
      30887: inst = 32'd268468224;
      30888: inst = 32'd201342976;
      30889: inst = 32'd203423744;
      30890: inst = 32'd471859200;
      30891: inst = 32'd136314880;
      30892: inst = 32'd268468224;
      30893: inst = 32'd201342977;
      30894: inst = 32'd203423744;
      30895: inst = 32'd471859200;
      30896: inst = 32'd136314880;
      30897: inst = 32'd268468224;
      30898: inst = 32'd201342978;
      30899: inst = 32'd203423744;
      30900: inst = 32'd471859200;
      30901: inst = 32'd136314880;
      30902: inst = 32'd268468224;
      30903: inst = 32'd201342979;
      30904: inst = 32'd203423744;
      30905: inst = 32'd471859200;
      30906: inst = 32'd136314880;
      30907: inst = 32'd268468224;
      30908: inst = 32'd201342980;
      30909: inst = 32'd203423744;
      30910: inst = 32'd471859200;
      30911: inst = 32'd136314880;
      30912: inst = 32'd268468224;
      30913: inst = 32'd201342981;
      30914: inst = 32'd203423744;
      30915: inst = 32'd471859200;
      30916: inst = 32'd136314880;
      30917: inst = 32'd268468224;
      30918: inst = 32'd201342982;
      30919: inst = 32'd203423744;
      30920: inst = 32'd471859200;
      30921: inst = 32'd136314880;
      30922: inst = 32'd268468224;
      30923: inst = 32'd201342983;
      30924: inst = 32'd203423744;
      30925: inst = 32'd471859200;
      30926: inst = 32'd136314880;
      30927: inst = 32'd268468224;
      30928: inst = 32'd201342984;
      30929: inst = 32'd203423744;
      30930: inst = 32'd471859200;
      30931: inst = 32'd136314880;
      30932: inst = 32'd268468224;
      30933: inst = 32'd201342985;
      30934: inst = 32'd203423744;
      30935: inst = 32'd471859200;
      30936: inst = 32'd136314880;
      30937: inst = 32'd268468224;
      30938: inst = 32'd201342986;
      30939: inst = 32'd203423744;
      30940: inst = 32'd471859200;
      30941: inst = 32'd136314880;
      30942: inst = 32'd268468224;
      30943: inst = 32'd201342987;
      30944: inst = 32'd203423744;
      30945: inst = 32'd471859200;
      30946: inst = 32'd136314880;
      30947: inst = 32'd268468224;
      30948: inst = 32'd201342988;
      30949: inst = 32'd203423744;
      30950: inst = 32'd471859200;
      30951: inst = 32'd136314880;
      30952: inst = 32'd268468224;
      30953: inst = 32'd201342989;
      30954: inst = 32'd203423744;
      30955: inst = 32'd471859200;
      30956: inst = 32'd136314880;
      30957: inst = 32'd268468224;
      30958: inst = 32'd201342990;
      30959: inst = 32'd203423744;
      30960: inst = 32'd471859200;
      30961: inst = 32'd136314880;
      30962: inst = 32'd268468224;
      30963: inst = 32'd201342991;
      30964: inst = 32'd203423744;
      30965: inst = 32'd471859200;
      30966: inst = 32'd136314880;
      30967: inst = 32'd268468224;
      30968: inst = 32'd201342992;
      30969: inst = 32'd203423744;
      30970: inst = 32'd471859200;
      30971: inst = 32'd136314880;
      30972: inst = 32'd268468224;
      30973: inst = 32'd201342993;
      30974: inst = 32'd203423744;
      30975: inst = 32'd471859200;
      30976: inst = 32'd136314880;
      30977: inst = 32'd268468224;
      30978: inst = 32'd201342994;
      30979: inst = 32'd203423744;
      30980: inst = 32'd471859200;
      30981: inst = 32'd136314880;
      30982: inst = 32'd268468224;
      30983: inst = 32'd201342995;
      30984: inst = 32'd203423744;
      30985: inst = 32'd471859200;
      30986: inst = 32'd136314880;
      30987: inst = 32'd268468224;
      30988: inst = 32'd201342996;
      30989: inst = 32'd203423744;
      30990: inst = 32'd471859200;
      30991: inst = 32'd136314880;
      30992: inst = 32'd268468224;
      30993: inst = 32'd201342997;
      30994: inst = 32'd203423744;
      30995: inst = 32'd471859200;
      30996: inst = 32'd136314880;
      30997: inst = 32'd268468224;
      30998: inst = 32'd201342998;
      30999: inst = 32'd203423744;
      31000: inst = 32'd471859200;
      31001: inst = 32'd136314880;
      31002: inst = 32'd268468224;
      31003: inst = 32'd201342999;
      31004: inst = 32'd203423744;
      31005: inst = 32'd471859200;
      31006: inst = 32'd136314880;
      31007: inst = 32'd268468224;
      31008: inst = 32'd201343000;
      31009: inst = 32'd203423744;
      31010: inst = 32'd471859200;
      31011: inst = 32'd136314880;
      31012: inst = 32'd268468224;
      31013: inst = 32'd201343001;
      31014: inst = 32'd203423744;
      31015: inst = 32'd471859200;
      31016: inst = 32'd136314880;
      31017: inst = 32'd268468224;
      31018: inst = 32'd201343002;
      31019: inst = 32'd203423744;
      31020: inst = 32'd471859200;
      31021: inst = 32'd136314880;
      31022: inst = 32'd268468224;
      31023: inst = 32'd201343003;
      31024: inst = 32'd203423744;
      31025: inst = 32'd471859200;
      31026: inst = 32'd136314880;
      31027: inst = 32'd268468224;
      31028: inst = 32'd201343004;
      31029: inst = 32'd203423744;
      31030: inst = 32'd471859200;
      31031: inst = 32'd136314880;
      31032: inst = 32'd268468224;
      31033: inst = 32'd201343005;
      31034: inst = 32'd203423744;
      31035: inst = 32'd471859200;
      31036: inst = 32'd136314880;
      31037: inst = 32'd268468224;
      31038: inst = 32'd201343006;
      31039: inst = 32'd203423744;
      31040: inst = 32'd471859200;
      31041: inst = 32'd136314880;
      31042: inst = 32'd268468224;
      31043: inst = 32'd201343007;
      31044: inst = 32'd203423744;
      31045: inst = 32'd471859200;
      31046: inst = 32'd136314880;
      31047: inst = 32'd268468224;
      31048: inst = 32'd201343008;
      31049: inst = 32'd203423744;
      31050: inst = 32'd471859200;
      31051: inst = 32'd136314880;
      31052: inst = 32'd268468224;
      31053: inst = 32'd201343009;
      31054: inst = 32'd203423744;
      31055: inst = 32'd471859200;
      31056: inst = 32'd136314880;
      31057: inst = 32'd268468224;
      31058: inst = 32'd201343010;
      31059: inst = 32'd203423744;
      31060: inst = 32'd471859200;
      31061: inst = 32'd136314880;
      31062: inst = 32'd268468224;
      31063: inst = 32'd201343011;
      31064: inst = 32'd203423744;
      31065: inst = 32'd471859200;
      31066: inst = 32'd136314880;
      31067: inst = 32'd268468224;
      31068: inst = 32'd201343012;
      31069: inst = 32'd203423744;
      31070: inst = 32'd471859200;
      31071: inst = 32'd136314880;
      31072: inst = 32'd268468224;
      31073: inst = 32'd201343013;
      31074: inst = 32'd203423744;
      31075: inst = 32'd471859200;
      31076: inst = 32'd136314880;
      31077: inst = 32'd268468224;
      31078: inst = 32'd201343014;
      31079: inst = 32'd203423744;
      31080: inst = 32'd471859200;
      31081: inst = 32'd136314880;
      31082: inst = 32'd268468224;
      31083: inst = 32'd201343015;
      31084: inst = 32'd203423744;
      31085: inst = 32'd471859200;
      31086: inst = 32'd136314880;
      31087: inst = 32'd268468224;
      31088: inst = 32'd201343016;
      31089: inst = 32'd203423744;
      31090: inst = 32'd471859200;
      31091: inst = 32'd136314880;
      31092: inst = 32'd268468224;
      31093: inst = 32'd201343017;
      31094: inst = 32'd203423744;
      31095: inst = 32'd471859200;
      31096: inst = 32'd136314880;
      31097: inst = 32'd268468224;
      31098: inst = 32'd201343018;
      31099: inst = 32'd203423744;
      31100: inst = 32'd471859200;
      31101: inst = 32'd136314880;
      31102: inst = 32'd268468224;
      31103: inst = 32'd201343019;
      31104: inst = 32'd203423744;
      31105: inst = 32'd471859200;
      31106: inst = 32'd136314880;
      31107: inst = 32'd268468224;
      31108: inst = 32'd201343020;
      31109: inst = 32'd203423744;
      31110: inst = 32'd471859200;
      31111: inst = 32'd136314880;
      31112: inst = 32'd268468224;
      31113: inst = 32'd201343021;
      31114: inst = 32'd203423744;
      31115: inst = 32'd471859200;
      31116: inst = 32'd136314880;
      31117: inst = 32'd268468224;
      31118: inst = 32'd201343022;
      31119: inst = 32'd203423744;
      31120: inst = 32'd471859200;
      31121: inst = 32'd136314880;
      31122: inst = 32'd268468224;
      31123: inst = 32'd201343023;
      31124: inst = 32'd203423744;
      31125: inst = 32'd471859200;
      31126: inst = 32'd136314880;
      31127: inst = 32'd268468224;
      31128: inst = 32'd201343024;
      31129: inst = 32'd203423744;
      31130: inst = 32'd471859200;
      31131: inst = 32'd136314880;
      31132: inst = 32'd268468224;
      31133: inst = 32'd201343025;
      31134: inst = 32'd203423744;
      31135: inst = 32'd471859200;
      31136: inst = 32'd136314880;
      31137: inst = 32'd268468224;
      31138: inst = 32'd201343026;
      31139: inst = 32'd203423744;
      31140: inst = 32'd471859200;
      31141: inst = 32'd136314880;
      31142: inst = 32'd268468224;
      31143: inst = 32'd201343027;
      31144: inst = 32'd203423744;
      31145: inst = 32'd471859200;
      31146: inst = 32'd136314880;
      31147: inst = 32'd268468224;
      31148: inst = 32'd201343028;
      31149: inst = 32'd203423744;
      31150: inst = 32'd471859200;
      31151: inst = 32'd136314880;
      31152: inst = 32'd268468224;
      31153: inst = 32'd201343029;
      31154: inst = 32'd203423744;
      31155: inst = 32'd471859200;
      31156: inst = 32'd136314880;
      31157: inst = 32'd268468224;
      31158: inst = 32'd201343030;
      31159: inst = 32'd203423744;
      31160: inst = 32'd471859200;
      31161: inst = 32'd136314880;
      31162: inst = 32'd268468224;
      31163: inst = 32'd201343031;
      31164: inst = 32'd203423744;
      31165: inst = 32'd471859200;
      31166: inst = 32'd136314880;
      31167: inst = 32'd268468224;
      31168: inst = 32'd201343032;
      31169: inst = 32'd203423744;
      31170: inst = 32'd471859200;
      31171: inst = 32'd136314880;
      31172: inst = 32'd268468224;
      31173: inst = 32'd201343033;
      31174: inst = 32'd203423744;
      31175: inst = 32'd471859200;
      31176: inst = 32'd136314880;
      31177: inst = 32'd268468224;
      31178: inst = 32'd201343034;
      31179: inst = 32'd203423744;
      31180: inst = 32'd471859200;
      31181: inst = 32'd136314880;
      31182: inst = 32'd268468224;
      31183: inst = 32'd201343035;
      31184: inst = 32'd203423744;
      31185: inst = 32'd471859200;
      31186: inst = 32'd136314880;
      31187: inst = 32'd268468224;
      31188: inst = 32'd201343036;
      31189: inst = 32'd203423744;
      31190: inst = 32'd471859200;
      31191: inst = 32'd136314880;
      31192: inst = 32'd268468224;
      31193: inst = 32'd201343037;
      31194: inst = 32'd203423744;
      31195: inst = 32'd471859200;
      31196: inst = 32'd136314880;
      31197: inst = 32'd268468224;
      31198: inst = 32'd201343038;
      31199: inst = 32'd203423744;
      31200: inst = 32'd471859200;
      31201: inst = 32'd136314880;
      31202: inst = 32'd268468224;
      31203: inst = 32'd201343039;
      31204: inst = 32'd203423744;
      31205: inst = 32'd471859200;
      31206: inst = 32'd136314880;
      31207: inst = 32'd268468224;
      31208: inst = 32'd201343040;
      31209: inst = 32'd203423744;
      31210: inst = 32'd471859200;
      31211: inst = 32'd136314880;
      31212: inst = 32'd268468224;
      31213: inst = 32'd201343041;
      31214: inst = 32'd203423744;
      31215: inst = 32'd471859200;
      31216: inst = 32'd136314880;
      31217: inst = 32'd268468224;
      31218: inst = 32'd201343042;
      31219: inst = 32'd203423744;
      31220: inst = 32'd471859200;
      31221: inst = 32'd136314880;
      31222: inst = 32'd268468224;
      31223: inst = 32'd201343043;
      31224: inst = 32'd203423744;
      31225: inst = 32'd471859200;
      31226: inst = 32'd136314880;
      31227: inst = 32'd268468224;
      31228: inst = 32'd201343044;
      31229: inst = 32'd203423744;
      31230: inst = 32'd471859200;
      31231: inst = 32'd136314880;
      31232: inst = 32'd268468224;
      31233: inst = 32'd201343045;
      31234: inst = 32'd203423744;
      31235: inst = 32'd471859200;
      31236: inst = 32'd136314880;
      31237: inst = 32'd268468224;
      31238: inst = 32'd201343046;
      31239: inst = 32'd203423744;
      31240: inst = 32'd471859200;
      31241: inst = 32'd136314880;
      31242: inst = 32'd268468224;
      31243: inst = 32'd201343047;
      31244: inst = 32'd203423744;
      31245: inst = 32'd471859200;
      31246: inst = 32'd136314880;
      31247: inst = 32'd268468224;
      31248: inst = 32'd201343048;
      31249: inst = 32'd203423744;
      31250: inst = 32'd471859200;
      31251: inst = 32'd136314880;
      31252: inst = 32'd268468224;
      31253: inst = 32'd201343049;
      31254: inst = 32'd203423744;
      31255: inst = 32'd471859200;
      31256: inst = 32'd136314880;
      31257: inst = 32'd268468224;
      31258: inst = 32'd201343050;
      31259: inst = 32'd203423744;
      31260: inst = 32'd471859200;
      31261: inst = 32'd136314880;
      31262: inst = 32'd268468224;
      31263: inst = 32'd201343051;
      31264: inst = 32'd203423744;
      31265: inst = 32'd471859200;
      31266: inst = 32'd136314880;
      31267: inst = 32'd268468224;
      31268: inst = 32'd201343052;
      31269: inst = 32'd203423744;
      31270: inst = 32'd471859200;
      31271: inst = 32'd136314880;
      31272: inst = 32'd268468224;
      31273: inst = 32'd201343053;
      31274: inst = 32'd203423744;
      31275: inst = 32'd471859200;
      31276: inst = 32'd136314880;
      31277: inst = 32'd268468224;
      31278: inst = 32'd201343054;
      31279: inst = 32'd203423744;
      31280: inst = 32'd471859200;
      31281: inst = 32'd136314880;
      31282: inst = 32'd268468224;
      31283: inst = 32'd201343055;
      31284: inst = 32'd203423744;
      31285: inst = 32'd471859200;
      31286: inst = 32'd136314880;
      31287: inst = 32'd268468224;
      31288: inst = 32'd201343056;
      31289: inst = 32'd203423744;
      31290: inst = 32'd471859200;
      31291: inst = 32'd136314880;
      31292: inst = 32'd268468224;
      31293: inst = 32'd201343057;
      31294: inst = 32'd203423744;
      31295: inst = 32'd471859200;
      31296: inst = 32'd136314880;
      31297: inst = 32'd268468224;
      31298: inst = 32'd201343058;
      31299: inst = 32'd203423744;
      31300: inst = 32'd471859200;
      31301: inst = 32'd136314880;
      31302: inst = 32'd268468224;
      31303: inst = 32'd201343059;
      31304: inst = 32'd203423744;
      31305: inst = 32'd471859200;
      31306: inst = 32'd136314880;
      31307: inst = 32'd268468224;
      31308: inst = 32'd201343060;
      31309: inst = 32'd203423744;
      31310: inst = 32'd471859200;
      31311: inst = 32'd136314880;
      31312: inst = 32'd268468224;
      31313: inst = 32'd201343061;
      31314: inst = 32'd203423744;
      31315: inst = 32'd471859200;
      31316: inst = 32'd136314880;
      31317: inst = 32'd268468224;
      31318: inst = 32'd201343062;
      31319: inst = 32'd203423744;
      31320: inst = 32'd471859200;
      31321: inst = 32'd136314880;
      31322: inst = 32'd268468224;
      31323: inst = 32'd201343063;
      31324: inst = 32'd203423744;
      31325: inst = 32'd471859200;
      31326: inst = 32'd136314880;
      31327: inst = 32'd268468224;
      31328: inst = 32'd201343064;
      31329: inst = 32'd203423744;
      31330: inst = 32'd471859200;
      31331: inst = 32'd136314880;
      31332: inst = 32'd268468224;
      31333: inst = 32'd201343065;
      31334: inst = 32'd203423744;
      31335: inst = 32'd471859200;
      31336: inst = 32'd136314880;
      31337: inst = 32'd268468224;
      31338: inst = 32'd201343066;
      31339: inst = 32'd203423744;
      31340: inst = 32'd471859200;
      31341: inst = 32'd136314880;
      31342: inst = 32'd268468224;
      31343: inst = 32'd201343067;
      31344: inst = 32'd203423744;
      31345: inst = 32'd471859200;
      31346: inst = 32'd136314880;
      31347: inst = 32'd268468224;
      31348: inst = 32'd201343068;
      31349: inst = 32'd203423744;
      31350: inst = 32'd471859200;
      31351: inst = 32'd136314880;
      31352: inst = 32'd268468224;
      31353: inst = 32'd201343069;
      31354: inst = 32'd203423744;
      31355: inst = 32'd471859200;
      31356: inst = 32'd136314880;
      31357: inst = 32'd268468224;
      31358: inst = 32'd201343070;
      31359: inst = 32'd203423744;
      31360: inst = 32'd471859200;
      31361: inst = 32'd136314880;
      31362: inst = 32'd268468224;
      31363: inst = 32'd201343071;
      31364: inst = 32'd203423744;
      31365: inst = 32'd471859200;
      31366: inst = 32'd136314880;
      31367: inst = 32'd268468224;
      31368: inst = 32'd201343072;
      31369: inst = 32'd203423744;
      31370: inst = 32'd471859200;
      31371: inst = 32'd136314880;
      31372: inst = 32'd268468224;
      31373: inst = 32'd201343073;
      31374: inst = 32'd203423744;
      31375: inst = 32'd471859200;
      31376: inst = 32'd136314880;
      31377: inst = 32'd268468224;
      31378: inst = 32'd201343074;
      31379: inst = 32'd203423744;
      31380: inst = 32'd471859200;
      31381: inst = 32'd136314880;
      31382: inst = 32'd268468224;
      31383: inst = 32'd201343075;
      31384: inst = 32'd203423744;
      31385: inst = 32'd471859200;
      31386: inst = 32'd136314880;
      31387: inst = 32'd268468224;
      31388: inst = 32'd201343076;
      31389: inst = 32'd203423744;
      31390: inst = 32'd471859200;
      31391: inst = 32'd136314880;
      31392: inst = 32'd268468224;
      31393: inst = 32'd201343077;
      31394: inst = 32'd203423744;
      31395: inst = 32'd471859200;
      31396: inst = 32'd136314880;
      31397: inst = 32'd268468224;
      31398: inst = 32'd201343078;
      31399: inst = 32'd203423744;
      31400: inst = 32'd471859200;
      31401: inst = 32'd136314880;
      31402: inst = 32'd268468224;
      31403: inst = 32'd201343079;
      31404: inst = 32'd203423744;
      31405: inst = 32'd471859200;
      31406: inst = 32'd136314880;
      31407: inst = 32'd268468224;
      31408: inst = 32'd201343080;
      31409: inst = 32'd203423744;
      31410: inst = 32'd471859200;
      31411: inst = 32'd136314880;
      31412: inst = 32'd268468224;
      31413: inst = 32'd201343081;
      31414: inst = 32'd203423744;
      31415: inst = 32'd471859200;
      31416: inst = 32'd136314880;
      31417: inst = 32'd268468224;
      31418: inst = 32'd201343082;
      31419: inst = 32'd203423744;
      31420: inst = 32'd471859200;
      31421: inst = 32'd136314880;
      31422: inst = 32'd268468224;
      31423: inst = 32'd201343083;
      31424: inst = 32'd203423744;
      31425: inst = 32'd471859200;
      31426: inst = 32'd136314880;
      31427: inst = 32'd268468224;
      31428: inst = 32'd201343084;
      31429: inst = 32'd203423744;
      31430: inst = 32'd471859200;
      31431: inst = 32'd136314880;
      31432: inst = 32'd268468224;
      31433: inst = 32'd201343085;
      31434: inst = 32'd203423744;
      31435: inst = 32'd471859200;
      31436: inst = 32'd136314880;
      31437: inst = 32'd268468224;
      31438: inst = 32'd201343086;
      31439: inst = 32'd203423744;
      31440: inst = 32'd471859200;
      31441: inst = 32'd136314880;
      31442: inst = 32'd268468224;
      31443: inst = 32'd201343087;
      31444: inst = 32'd203423744;
      31445: inst = 32'd471859200;
      31446: inst = 32'd136314880;
      31447: inst = 32'd268468224;
      31448: inst = 32'd201343088;
      31449: inst = 32'd203423744;
      31450: inst = 32'd471859200;
      31451: inst = 32'd136314880;
      31452: inst = 32'd268468224;
      31453: inst = 32'd201343089;
      31454: inst = 32'd203423744;
      31455: inst = 32'd471859200;
      31456: inst = 32'd136314880;
      31457: inst = 32'd268468224;
      31458: inst = 32'd201343090;
      31459: inst = 32'd203423744;
      31460: inst = 32'd471859200;
      31461: inst = 32'd136314880;
      31462: inst = 32'd268468224;
      31463: inst = 32'd201343091;
      31464: inst = 32'd203423744;
      31465: inst = 32'd471859200;
      31466: inst = 32'd136314880;
      31467: inst = 32'd268468224;
      31468: inst = 32'd201343092;
      31469: inst = 32'd203423744;
      31470: inst = 32'd471859200;
      31471: inst = 32'd136314880;
      31472: inst = 32'd268468224;
      31473: inst = 32'd201343093;
      31474: inst = 32'd203423744;
      31475: inst = 32'd471859200;
      31476: inst = 32'd136314880;
      31477: inst = 32'd268468224;
      31478: inst = 32'd201343094;
      31479: inst = 32'd203423744;
      31480: inst = 32'd471859200;
      31481: inst = 32'd136314880;
      31482: inst = 32'd268468224;
      31483: inst = 32'd201343095;
      31484: inst = 32'd203423744;
      31485: inst = 32'd471859200;
      31486: inst = 32'd136314880;
      31487: inst = 32'd268468224;
      31488: inst = 32'd201343096;
      31489: inst = 32'd203423744;
      31490: inst = 32'd471859200;
      31491: inst = 32'd136314880;
      31492: inst = 32'd268468224;
      31493: inst = 32'd201343097;
      31494: inst = 32'd203423744;
      31495: inst = 32'd471859200;
      31496: inst = 32'd136314880;
      31497: inst = 32'd268468224;
      31498: inst = 32'd201343098;
      31499: inst = 32'd203423744;
      31500: inst = 32'd471859200;
      31501: inst = 32'd136314880;
      31502: inst = 32'd268468224;
      31503: inst = 32'd201343099;
      31504: inst = 32'd203423744;
      31505: inst = 32'd471859200;
      31506: inst = 32'd136314880;
      31507: inst = 32'd268468224;
      31508: inst = 32'd201343100;
      31509: inst = 32'd203423744;
      31510: inst = 32'd471859200;
      31511: inst = 32'd136314880;
      31512: inst = 32'd268468224;
      31513: inst = 32'd201343101;
      31514: inst = 32'd203423744;
      31515: inst = 32'd471859200;
      31516: inst = 32'd136314880;
      31517: inst = 32'd268468224;
      31518: inst = 32'd201343102;
      31519: inst = 32'd203423744;
      31520: inst = 32'd471859200;
      31521: inst = 32'd136314880;
      31522: inst = 32'd268468224;
      31523: inst = 32'd201343103;
      31524: inst = 32'd203423744;
      31525: inst = 32'd471859200;
      31526: inst = 32'd136314880;
      31527: inst = 32'd268468224;
      31528: inst = 32'd201343104;
      31529: inst = 32'd203423744;
      31530: inst = 32'd471859200;
      31531: inst = 32'd136314880;
      31532: inst = 32'd268468224;
      31533: inst = 32'd201343105;
      31534: inst = 32'd203423744;
      31535: inst = 32'd471859200;
      31536: inst = 32'd136314880;
      31537: inst = 32'd268468224;
      31538: inst = 32'd201343106;
      31539: inst = 32'd203423744;
      31540: inst = 32'd471859200;
      31541: inst = 32'd136314880;
      31542: inst = 32'd268468224;
      31543: inst = 32'd201343107;
      31544: inst = 32'd203423744;
      31545: inst = 32'd471859200;
      31546: inst = 32'd136314880;
      31547: inst = 32'd268468224;
      31548: inst = 32'd201343108;
      31549: inst = 32'd203423744;
      31550: inst = 32'd471859200;
      31551: inst = 32'd136314880;
      31552: inst = 32'd268468224;
      31553: inst = 32'd201343109;
      31554: inst = 32'd203423744;
      31555: inst = 32'd471859200;
      31556: inst = 32'd136314880;
      31557: inst = 32'd268468224;
      31558: inst = 32'd201343110;
      31559: inst = 32'd203423744;
      31560: inst = 32'd471859200;
      31561: inst = 32'd136314880;
      31562: inst = 32'd268468224;
      31563: inst = 32'd201343111;
      31564: inst = 32'd203423744;
      31565: inst = 32'd471859200;
      31566: inst = 32'd136314880;
      31567: inst = 32'd268468224;
      31568: inst = 32'd201343112;
      31569: inst = 32'd203423744;
      31570: inst = 32'd471859200;
      31571: inst = 32'd136314880;
      31572: inst = 32'd268468224;
      31573: inst = 32'd201343113;
      31574: inst = 32'd203423744;
      31575: inst = 32'd471859200;
      31576: inst = 32'd136314880;
      31577: inst = 32'd268468224;
      31578: inst = 32'd201343114;
      31579: inst = 32'd203423744;
      31580: inst = 32'd471859200;
      31581: inst = 32'd136314880;
      31582: inst = 32'd268468224;
      31583: inst = 32'd201343115;
      31584: inst = 32'd203423744;
      31585: inst = 32'd471859200;
      31586: inst = 32'd136314880;
      31587: inst = 32'd268468224;
      31588: inst = 32'd201343116;
      31589: inst = 32'd203423744;
      31590: inst = 32'd471859200;
      31591: inst = 32'd136314880;
      31592: inst = 32'd268468224;
      31593: inst = 32'd201343117;
      31594: inst = 32'd203423744;
      31595: inst = 32'd471859200;
      31596: inst = 32'd136314880;
      31597: inst = 32'd268468224;
      31598: inst = 32'd201343118;
      31599: inst = 32'd203423744;
      31600: inst = 32'd471859200;
      31601: inst = 32'd136314880;
      31602: inst = 32'd268468224;
      31603: inst = 32'd201343119;
      31604: inst = 32'd203423744;
      31605: inst = 32'd471859200;
      31606: inst = 32'd136314880;
      31607: inst = 32'd268468224;
      31608: inst = 32'd201343120;
      31609: inst = 32'd203423744;
      31610: inst = 32'd471859200;
      31611: inst = 32'd136314880;
      31612: inst = 32'd268468224;
      31613: inst = 32'd201343121;
      31614: inst = 32'd203423744;
      31615: inst = 32'd471859200;
      31616: inst = 32'd136314880;
      31617: inst = 32'd268468224;
      31618: inst = 32'd201343122;
      31619: inst = 32'd203423744;
      31620: inst = 32'd471859200;
      31621: inst = 32'd136314880;
      31622: inst = 32'd268468224;
      31623: inst = 32'd201343123;
      31624: inst = 32'd203423744;
      31625: inst = 32'd471859200;
      31626: inst = 32'd136314880;
      31627: inst = 32'd268468224;
      31628: inst = 32'd201343124;
      31629: inst = 32'd203423744;
      31630: inst = 32'd471859200;
      31631: inst = 32'd136314880;
      31632: inst = 32'd268468224;
      31633: inst = 32'd201343125;
      31634: inst = 32'd203423744;
      31635: inst = 32'd471859200;
      31636: inst = 32'd136314880;
      31637: inst = 32'd268468224;
      31638: inst = 32'd201343126;
      31639: inst = 32'd203423744;
      31640: inst = 32'd471859200;
      31641: inst = 32'd136314880;
      31642: inst = 32'd268468224;
      31643: inst = 32'd201343127;
      31644: inst = 32'd203423744;
      31645: inst = 32'd471859200;
      31646: inst = 32'd136314880;
      31647: inst = 32'd268468224;
      31648: inst = 32'd201343128;
      31649: inst = 32'd203423744;
      31650: inst = 32'd471859200;
      31651: inst = 32'd136314880;
      31652: inst = 32'd268468224;
      31653: inst = 32'd201343129;
      31654: inst = 32'd203423744;
      31655: inst = 32'd471859200;
      31656: inst = 32'd136314880;
      31657: inst = 32'd268468224;
      31658: inst = 32'd201343130;
      31659: inst = 32'd203423744;
      31660: inst = 32'd471859200;
      31661: inst = 32'd136314880;
      31662: inst = 32'd268468224;
      31663: inst = 32'd201343131;
      31664: inst = 32'd203423744;
      31665: inst = 32'd471859200;
      31666: inst = 32'd136314880;
      31667: inst = 32'd268468224;
      31668: inst = 32'd201343132;
      31669: inst = 32'd203423744;
      31670: inst = 32'd471859200;
      31671: inst = 32'd136314880;
      31672: inst = 32'd268468224;
      31673: inst = 32'd201343133;
      31674: inst = 32'd203423744;
      31675: inst = 32'd471859200;
      31676: inst = 32'd136314880;
      31677: inst = 32'd268468224;
      31678: inst = 32'd201343134;
      31679: inst = 32'd203423744;
      31680: inst = 32'd471859200;
      31681: inst = 32'd136314880;
      31682: inst = 32'd268468224;
      31683: inst = 32'd201343135;
      31684: inst = 32'd203423744;
      31685: inst = 32'd471859200;
      31686: inst = 32'd136314880;
      31687: inst = 32'd268468224;
      31688: inst = 32'd201343136;
      31689: inst = 32'd203423744;
      31690: inst = 32'd471859200;
      31691: inst = 32'd136314880;
      31692: inst = 32'd268468224;
      31693: inst = 32'd201343137;
      31694: inst = 32'd203423744;
      31695: inst = 32'd471859200;
      31696: inst = 32'd136314880;
      31697: inst = 32'd268468224;
      31698: inst = 32'd201343138;
      31699: inst = 32'd203423744;
      31700: inst = 32'd471859200;
      31701: inst = 32'd136314880;
      31702: inst = 32'd268468224;
      31703: inst = 32'd201343139;
      31704: inst = 32'd203423744;
      31705: inst = 32'd471859200;
      31706: inst = 32'd136314880;
      31707: inst = 32'd268468224;
      31708: inst = 32'd201343140;
      31709: inst = 32'd203423744;
      31710: inst = 32'd471859200;
      31711: inst = 32'd136314880;
      31712: inst = 32'd268468224;
      31713: inst = 32'd201343141;
      31714: inst = 32'd203423744;
      31715: inst = 32'd471859200;
      31716: inst = 32'd136314880;
      31717: inst = 32'd268468224;
      31718: inst = 32'd201343142;
      31719: inst = 32'd203423744;
      31720: inst = 32'd471859200;
      31721: inst = 32'd136314880;
      31722: inst = 32'd268468224;
      31723: inst = 32'd201343143;
      31724: inst = 32'd203423744;
      31725: inst = 32'd471859200;
      31726: inst = 32'd136314880;
      31727: inst = 32'd268468224;
      31728: inst = 32'd201343144;
      31729: inst = 32'd203423744;
      31730: inst = 32'd471859200;
      31731: inst = 32'd136314880;
      31732: inst = 32'd268468224;
      31733: inst = 32'd201343145;
      31734: inst = 32'd203423744;
      31735: inst = 32'd471859200;
      31736: inst = 32'd136314880;
      31737: inst = 32'd268468224;
      31738: inst = 32'd201343146;
      31739: inst = 32'd203423744;
      31740: inst = 32'd471859200;
      31741: inst = 32'd136314880;
      31742: inst = 32'd268468224;
      31743: inst = 32'd201343147;
      31744: inst = 32'd203423744;
      31745: inst = 32'd471859200;
      31746: inst = 32'd136314880;
      31747: inst = 32'd268468224;
      31748: inst = 32'd201343148;
      31749: inst = 32'd203423744;
      31750: inst = 32'd471859200;
      31751: inst = 32'd136314880;
      31752: inst = 32'd268468224;
      31753: inst = 32'd201343149;
      31754: inst = 32'd203423744;
      31755: inst = 32'd471859200;
      31756: inst = 32'd136314880;
      31757: inst = 32'd268468224;
      31758: inst = 32'd201343150;
      31759: inst = 32'd203423744;
      31760: inst = 32'd471859200;
      31761: inst = 32'd136314880;
      31762: inst = 32'd268468224;
      31763: inst = 32'd201343151;
      31764: inst = 32'd203423744;
      31765: inst = 32'd471859200;
      31766: inst = 32'd136314880;
      31767: inst = 32'd268468224;
      31768: inst = 32'd201343152;
      31769: inst = 32'd203423744;
      31770: inst = 32'd471859200;
      31771: inst = 32'd136314880;
      31772: inst = 32'd268468224;
      31773: inst = 32'd201343153;
      31774: inst = 32'd203423744;
      31775: inst = 32'd471859200;
      31776: inst = 32'd136314880;
      31777: inst = 32'd268468224;
      31778: inst = 32'd201343154;
      31779: inst = 32'd203423744;
      31780: inst = 32'd471859200;
      31781: inst = 32'd136314880;
      31782: inst = 32'd268468224;
      31783: inst = 32'd201343155;
      31784: inst = 32'd203423744;
      31785: inst = 32'd471859200;
      31786: inst = 32'd136314880;
      31787: inst = 32'd268468224;
      31788: inst = 32'd201343156;
      31789: inst = 32'd203423744;
      31790: inst = 32'd471859200;
      31791: inst = 32'd136314880;
      31792: inst = 32'd268468224;
      31793: inst = 32'd201343157;
      31794: inst = 32'd203423744;
      31795: inst = 32'd471859200;
      31796: inst = 32'd136314880;
      31797: inst = 32'd268468224;
      31798: inst = 32'd201343158;
      31799: inst = 32'd203423744;
      31800: inst = 32'd471859200;
      31801: inst = 32'd136314880;
      31802: inst = 32'd268468224;
      31803: inst = 32'd201343159;
      31804: inst = 32'd203423744;
      31805: inst = 32'd471859200;
      31806: inst = 32'd136314880;
      31807: inst = 32'd268468224;
      31808: inst = 32'd201343160;
      31809: inst = 32'd203423744;
      31810: inst = 32'd471859200;
      31811: inst = 32'd136314880;
      31812: inst = 32'd268468224;
      31813: inst = 32'd201343161;
      31814: inst = 32'd203423744;
      31815: inst = 32'd471859200;
      31816: inst = 32'd136314880;
      31817: inst = 32'd268468224;
      31818: inst = 32'd201343162;
      31819: inst = 32'd203423744;
      31820: inst = 32'd471859200;
      31821: inst = 32'd136314880;
      31822: inst = 32'd268468224;
      31823: inst = 32'd201343163;
      31824: inst = 32'd203423744;
      31825: inst = 32'd471859200;
      31826: inst = 32'd136314880;
      31827: inst = 32'd268468224;
      31828: inst = 32'd201343164;
      31829: inst = 32'd203423744;
      31830: inst = 32'd471859200;
      31831: inst = 32'd136314880;
      31832: inst = 32'd268468224;
      31833: inst = 32'd201343165;
      31834: inst = 32'd203423744;
      31835: inst = 32'd471859200;
      31836: inst = 32'd136314880;
      31837: inst = 32'd268468224;
      31838: inst = 32'd201343166;
      31839: inst = 32'd203423744;
      31840: inst = 32'd471859200;
      31841: inst = 32'd136314880;
      31842: inst = 32'd268468224;
      31843: inst = 32'd201343167;
      31844: inst = 32'd203423744;
      31845: inst = 32'd471859200;
      31846: inst = 32'd136314880;
      31847: inst = 32'd268468224;
      31848: inst = 32'd201343168;
      31849: inst = 32'd203423744;
      31850: inst = 32'd471859200;
      31851: inst = 32'd136314880;
      31852: inst = 32'd268468224;
      31853: inst = 32'd201343169;
      31854: inst = 32'd203423744;
      31855: inst = 32'd471859200;
      31856: inst = 32'd136314880;
      31857: inst = 32'd268468224;
      31858: inst = 32'd201343170;
      31859: inst = 32'd203423744;
      31860: inst = 32'd471859200;
      31861: inst = 32'd136314880;
      31862: inst = 32'd268468224;
      31863: inst = 32'd201343171;
      31864: inst = 32'd203423744;
      31865: inst = 32'd471859200;
      31866: inst = 32'd136314880;
      31867: inst = 32'd268468224;
      31868: inst = 32'd201343172;
      31869: inst = 32'd203423744;
      31870: inst = 32'd471859200;
      31871: inst = 32'd136314880;
      31872: inst = 32'd268468224;
      31873: inst = 32'd201343173;
      31874: inst = 32'd203423744;
      31875: inst = 32'd471859200;
      31876: inst = 32'd136314880;
      31877: inst = 32'd268468224;
      31878: inst = 32'd201343174;
      31879: inst = 32'd203423744;
      31880: inst = 32'd471859200;
      31881: inst = 32'd136314880;
      31882: inst = 32'd268468224;
      31883: inst = 32'd201343175;
      31884: inst = 32'd203423744;
      31885: inst = 32'd471859200;
      31886: inst = 32'd136314880;
      31887: inst = 32'd268468224;
      31888: inst = 32'd201343176;
      31889: inst = 32'd203423744;
      31890: inst = 32'd471859200;
      31891: inst = 32'd136314880;
      31892: inst = 32'd268468224;
      31893: inst = 32'd201343177;
      31894: inst = 32'd203423744;
      31895: inst = 32'd471859200;
      31896: inst = 32'd136314880;
      31897: inst = 32'd268468224;
      31898: inst = 32'd201343178;
      31899: inst = 32'd203423744;
      31900: inst = 32'd471859200;
      31901: inst = 32'd136314880;
      31902: inst = 32'd268468224;
      31903: inst = 32'd201343179;
      31904: inst = 32'd203423744;
      31905: inst = 32'd471859200;
      31906: inst = 32'd136314880;
      31907: inst = 32'd268468224;
      31908: inst = 32'd201343180;
      31909: inst = 32'd203423744;
      31910: inst = 32'd471859200;
      31911: inst = 32'd136314880;
      31912: inst = 32'd268468224;
      31913: inst = 32'd201343181;
      31914: inst = 32'd203423744;
      31915: inst = 32'd471859200;
      31916: inst = 32'd136314880;
      31917: inst = 32'd268468224;
      31918: inst = 32'd201343182;
      31919: inst = 32'd203423744;
      31920: inst = 32'd471859200;
      31921: inst = 32'd136314880;
      31922: inst = 32'd268468224;
      31923: inst = 32'd201343183;
      31924: inst = 32'd203423744;
      31925: inst = 32'd471859200;
      31926: inst = 32'd136314880;
      31927: inst = 32'd268468224;
      31928: inst = 32'd201343184;
      31929: inst = 32'd203423744;
      31930: inst = 32'd471859200;
      31931: inst = 32'd136314880;
      31932: inst = 32'd268468224;
      31933: inst = 32'd201343185;
      31934: inst = 32'd203423744;
      31935: inst = 32'd471859200;
      31936: inst = 32'd136314880;
      31937: inst = 32'd268468224;
      31938: inst = 32'd201343186;
      31939: inst = 32'd203423744;
      31940: inst = 32'd471859200;
      31941: inst = 32'd136314880;
      31942: inst = 32'd268468224;
      31943: inst = 32'd201343187;
      31944: inst = 32'd203423744;
      31945: inst = 32'd471859200;
      31946: inst = 32'd136314880;
      31947: inst = 32'd268468224;
      31948: inst = 32'd201343188;
      31949: inst = 32'd203423744;
      31950: inst = 32'd471859200;
      31951: inst = 32'd136314880;
      31952: inst = 32'd268468224;
      31953: inst = 32'd201343189;
      31954: inst = 32'd203423744;
      31955: inst = 32'd471859200;
      31956: inst = 32'd136314880;
      31957: inst = 32'd268468224;
      31958: inst = 32'd201343190;
      31959: inst = 32'd203423744;
      31960: inst = 32'd471859200;
      31961: inst = 32'd136314880;
      31962: inst = 32'd268468224;
      31963: inst = 32'd201343191;
      31964: inst = 32'd203423744;
      31965: inst = 32'd471859200;
      31966: inst = 32'd136314880;
      31967: inst = 32'd268468224;
      31968: inst = 32'd201343192;
      31969: inst = 32'd203423744;
      31970: inst = 32'd471859200;
      31971: inst = 32'd136314880;
      31972: inst = 32'd268468224;
      31973: inst = 32'd201343193;
      31974: inst = 32'd203423744;
      31975: inst = 32'd471859200;
      31976: inst = 32'd136314880;
      31977: inst = 32'd268468224;
      31978: inst = 32'd201343194;
      31979: inst = 32'd203423744;
      31980: inst = 32'd471859200;
      31981: inst = 32'd136314880;
      31982: inst = 32'd268468224;
      31983: inst = 32'd201343195;
      31984: inst = 32'd203423744;
      31985: inst = 32'd471859200;
      31986: inst = 32'd136314880;
      31987: inst = 32'd268468224;
      31988: inst = 32'd201343196;
      31989: inst = 32'd203423744;
      31990: inst = 32'd471859200;
      31991: inst = 32'd136314880;
      31992: inst = 32'd268468224;
      31993: inst = 32'd201343197;
      31994: inst = 32'd203423744;
      31995: inst = 32'd471859200;
      31996: inst = 32'd136314880;
      31997: inst = 32'd268468224;
      31998: inst = 32'd201343198;
      31999: inst = 32'd203423744;
      32000: inst = 32'd471859200;
      32001: inst = 32'd136314880;
      32002: inst = 32'd268468224;
      32003: inst = 32'd201343199;
      32004: inst = 32'd203423744;
      32005: inst = 32'd471859200;
      32006: inst = 32'd136314880;
      32007: inst = 32'd268468224;
      32008: inst = 32'd201343200;
      32009: inst = 32'd203423744;
      32010: inst = 32'd471859200;
      32011: inst = 32'd136314880;
      32012: inst = 32'd268468224;
      32013: inst = 32'd201343201;
      32014: inst = 32'd203423744;
      32015: inst = 32'd471859200;
      32016: inst = 32'd136314880;
      32017: inst = 32'd268468224;
      32018: inst = 32'd201343202;
      32019: inst = 32'd203423744;
      32020: inst = 32'd471859200;
      32021: inst = 32'd136314880;
      32022: inst = 32'd268468224;
      32023: inst = 32'd201343203;
      32024: inst = 32'd203423744;
      32025: inst = 32'd471859200;
      32026: inst = 32'd136314880;
      32027: inst = 32'd268468224;
      32028: inst = 32'd201343204;
      32029: inst = 32'd203423744;
      32030: inst = 32'd471859200;
      32031: inst = 32'd136314880;
      32032: inst = 32'd268468224;
      32033: inst = 32'd201343205;
      32034: inst = 32'd203423744;
      32035: inst = 32'd471859200;
      32036: inst = 32'd136314880;
      32037: inst = 32'd268468224;
      32038: inst = 32'd201343206;
      32039: inst = 32'd203423744;
      32040: inst = 32'd471859200;
      32041: inst = 32'd136314880;
      32042: inst = 32'd268468224;
      32043: inst = 32'd201343207;
      32044: inst = 32'd203423744;
      32045: inst = 32'd471859200;
      32046: inst = 32'd136314880;
      32047: inst = 32'd268468224;
      32048: inst = 32'd201343208;
      32049: inst = 32'd203423744;
      32050: inst = 32'd471859200;
      32051: inst = 32'd136314880;
      32052: inst = 32'd268468224;
      32053: inst = 32'd201343209;
      32054: inst = 32'd203423744;
      32055: inst = 32'd471859200;
      32056: inst = 32'd136314880;
      32057: inst = 32'd268468224;
      32058: inst = 32'd201343210;
      32059: inst = 32'd203423744;
      32060: inst = 32'd471859200;
      32061: inst = 32'd136314880;
      32062: inst = 32'd268468224;
      32063: inst = 32'd201343211;
      32064: inst = 32'd203423744;
      32065: inst = 32'd471859200;
      32066: inst = 32'd136314880;
      32067: inst = 32'd268468224;
      32068: inst = 32'd201343212;
      32069: inst = 32'd203423744;
      32070: inst = 32'd471859200;
      32071: inst = 32'd136314880;
      32072: inst = 32'd268468224;
      32073: inst = 32'd201343213;
      32074: inst = 32'd203423744;
      32075: inst = 32'd471859200;
      32076: inst = 32'd136314880;
      32077: inst = 32'd268468224;
      32078: inst = 32'd201343214;
      32079: inst = 32'd203423744;
      32080: inst = 32'd471859200;
      32081: inst = 32'd136314880;
      32082: inst = 32'd268468224;
      32083: inst = 32'd201343215;
      32084: inst = 32'd203423744;
      32085: inst = 32'd471859200;
      32086: inst = 32'd136314880;
      32087: inst = 32'd268468224;
      32088: inst = 32'd201343216;
      32089: inst = 32'd203423744;
      32090: inst = 32'd471859200;
      32091: inst = 32'd136314880;
      32092: inst = 32'd268468224;
      32093: inst = 32'd201343217;
      32094: inst = 32'd203423744;
      32095: inst = 32'd471859200;
      32096: inst = 32'd136314880;
      32097: inst = 32'd268468224;
      32098: inst = 32'd201343218;
      32099: inst = 32'd203423744;
      32100: inst = 32'd471859200;
      32101: inst = 32'd136314880;
      32102: inst = 32'd268468224;
      32103: inst = 32'd201343219;
      32104: inst = 32'd203423744;
      32105: inst = 32'd471859200;
      32106: inst = 32'd136314880;
      32107: inst = 32'd268468224;
      32108: inst = 32'd201343220;
      32109: inst = 32'd203423744;
      32110: inst = 32'd471859200;
      32111: inst = 32'd136314880;
      32112: inst = 32'd268468224;
      32113: inst = 32'd201343221;
      32114: inst = 32'd203423744;
      32115: inst = 32'd471859200;
      32116: inst = 32'd136314880;
      32117: inst = 32'd268468224;
      32118: inst = 32'd201343222;
      32119: inst = 32'd203423744;
      32120: inst = 32'd471859200;
      32121: inst = 32'd136314880;
      32122: inst = 32'd268468224;
      32123: inst = 32'd201343223;
      32124: inst = 32'd203423744;
      32125: inst = 32'd471859200;
      32126: inst = 32'd136314880;
      32127: inst = 32'd268468224;
      32128: inst = 32'd201343224;
      32129: inst = 32'd203423744;
      32130: inst = 32'd471859200;
      32131: inst = 32'd136314880;
      32132: inst = 32'd268468224;
      32133: inst = 32'd201343225;
      32134: inst = 32'd203423744;
      32135: inst = 32'd471859200;
      32136: inst = 32'd136314880;
      32137: inst = 32'd268468224;
      32138: inst = 32'd201343226;
      32139: inst = 32'd203423744;
      32140: inst = 32'd471859200;
      32141: inst = 32'd136314880;
      32142: inst = 32'd268468224;
      32143: inst = 32'd201343227;
      32144: inst = 32'd203423744;
      32145: inst = 32'd471859200;
      32146: inst = 32'd136314880;
      32147: inst = 32'd268468224;
      32148: inst = 32'd201343228;
      32149: inst = 32'd203423744;
      32150: inst = 32'd471859200;
      32151: inst = 32'd136314880;
      32152: inst = 32'd268468224;
      32153: inst = 32'd201343229;
      32154: inst = 32'd203423744;
      32155: inst = 32'd471859200;
      32156: inst = 32'd136314880;
      32157: inst = 32'd268468224;
      32158: inst = 32'd201343230;
      32159: inst = 32'd203423744;
      32160: inst = 32'd471859200;
      32161: inst = 32'd136314880;
      32162: inst = 32'd268468224;
      32163: inst = 32'd201343231;
      32164: inst = 32'd203423744;
      32165: inst = 32'd471859200;
      32166: inst = 32'd136314880;
      32167: inst = 32'd268468224;
      32168: inst = 32'd201343232;
      32169: inst = 32'd203423744;
      32170: inst = 32'd471859200;
      32171: inst = 32'd136314880;
      32172: inst = 32'd268468224;
      32173: inst = 32'd201343233;
      32174: inst = 32'd203423744;
      32175: inst = 32'd471859200;
      32176: inst = 32'd136314880;
      32177: inst = 32'd268468224;
      32178: inst = 32'd201343234;
      32179: inst = 32'd203423744;
      32180: inst = 32'd471859200;
      32181: inst = 32'd136314880;
      32182: inst = 32'd268468224;
      32183: inst = 32'd201343235;
      32184: inst = 32'd203423744;
      32185: inst = 32'd471859200;
      32186: inst = 32'd136314880;
      32187: inst = 32'd268468224;
      32188: inst = 32'd201343236;
      32189: inst = 32'd203423744;
      32190: inst = 32'd471859200;
      32191: inst = 32'd136314880;
      32192: inst = 32'd268468224;
      32193: inst = 32'd201343237;
      32194: inst = 32'd203423744;
      32195: inst = 32'd471859200;
      32196: inst = 32'd136314880;
      32197: inst = 32'd268468224;
      32198: inst = 32'd201343238;
      32199: inst = 32'd203423744;
      32200: inst = 32'd471859200;
      32201: inst = 32'd136314880;
      32202: inst = 32'd268468224;
      32203: inst = 32'd201343239;
      32204: inst = 32'd203423744;
      32205: inst = 32'd471859200;
      32206: inst = 32'd136314880;
      32207: inst = 32'd268468224;
      32208: inst = 32'd201343240;
      32209: inst = 32'd203423744;
      32210: inst = 32'd471859200;
      32211: inst = 32'd136314880;
      32212: inst = 32'd268468224;
      32213: inst = 32'd201343241;
      32214: inst = 32'd203423744;
      32215: inst = 32'd471859200;
      32216: inst = 32'd136314880;
      32217: inst = 32'd268468224;
      32218: inst = 32'd201343242;
      32219: inst = 32'd203423744;
      32220: inst = 32'd471859200;
      32221: inst = 32'd136314880;
      32222: inst = 32'd268468224;
      32223: inst = 32'd201343243;
      32224: inst = 32'd203423744;
      32225: inst = 32'd471859200;
      32226: inst = 32'd136314880;
      32227: inst = 32'd268468224;
      32228: inst = 32'd201343244;
      32229: inst = 32'd203423744;
      32230: inst = 32'd471859200;
      32231: inst = 32'd136314880;
      32232: inst = 32'd268468224;
      32233: inst = 32'd201343245;
      32234: inst = 32'd203423744;
      32235: inst = 32'd471859200;
      32236: inst = 32'd136314880;
      32237: inst = 32'd268468224;
      32238: inst = 32'd201343246;
      32239: inst = 32'd203423744;
      32240: inst = 32'd471859200;
      32241: inst = 32'd136314880;
      32242: inst = 32'd268468224;
      32243: inst = 32'd201343247;
      32244: inst = 32'd203423744;
      32245: inst = 32'd471859200;
      32246: inst = 32'd136314880;
      32247: inst = 32'd268468224;
      32248: inst = 32'd201343248;
      32249: inst = 32'd203423744;
      32250: inst = 32'd471859200;
      32251: inst = 32'd136314880;
      32252: inst = 32'd268468224;
      32253: inst = 32'd201343249;
      32254: inst = 32'd203423744;
      32255: inst = 32'd471859200;
      32256: inst = 32'd136314880;
      32257: inst = 32'd268468224;
      32258: inst = 32'd201343250;
      32259: inst = 32'd203423744;
      32260: inst = 32'd471859200;
      32261: inst = 32'd136314880;
      32262: inst = 32'd268468224;
      32263: inst = 32'd201343251;
      32264: inst = 32'd203423744;
      32265: inst = 32'd471859200;
      32266: inst = 32'd136314880;
      32267: inst = 32'd268468224;
      32268: inst = 32'd201343252;
      32269: inst = 32'd203423744;
      32270: inst = 32'd471859200;
      32271: inst = 32'd136314880;
      32272: inst = 32'd268468224;
      32273: inst = 32'd201343253;
      32274: inst = 32'd203423744;
      32275: inst = 32'd471859200;
      32276: inst = 32'd136314880;
      32277: inst = 32'd268468224;
      32278: inst = 32'd201343254;
      32279: inst = 32'd203423744;
      32280: inst = 32'd471859200;
      32281: inst = 32'd136314880;
      32282: inst = 32'd268468224;
      32283: inst = 32'd201343255;
      32284: inst = 32'd203423744;
      32285: inst = 32'd471859200;
      32286: inst = 32'd136314880;
      32287: inst = 32'd268468224;
      32288: inst = 32'd201343256;
      32289: inst = 32'd203423744;
      32290: inst = 32'd471859200;
      32291: inst = 32'd136314880;
      32292: inst = 32'd268468224;
      32293: inst = 32'd201343257;
      32294: inst = 32'd203423744;
      32295: inst = 32'd471859200;
      32296: inst = 32'd136314880;
      32297: inst = 32'd268468224;
      32298: inst = 32'd201343258;
      32299: inst = 32'd203423744;
      32300: inst = 32'd471859200;
      32301: inst = 32'd136314880;
      32302: inst = 32'd268468224;
      32303: inst = 32'd201343259;
      32304: inst = 32'd203423744;
      32305: inst = 32'd471859200;
      32306: inst = 32'd136314880;
      32307: inst = 32'd268468224;
      32308: inst = 32'd201343260;
      32309: inst = 32'd203423744;
      32310: inst = 32'd471859200;
      32311: inst = 32'd136314880;
      32312: inst = 32'd268468224;
      32313: inst = 32'd201343261;
      32314: inst = 32'd203423744;
      32315: inst = 32'd471859200;
      32316: inst = 32'd136314880;
      32317: inst = 32'd268468224;
      32318: inst = 32'd201343262;
      32319: inst = 32'd203423744;
      32320: inst = 32'd471859200;
      32321: inst = 32'd136314880;
      32322: inst = 32'd268468224;
      32323: inst = 32'd201343263;
      32324: inst = 32'd203423744;
      32325: inst = 32'd471859200;
      32326: inst = 32'd136314880;
      32327: inst = 32'd268468224;
      32328: inst = 32'd201343264;
      32329: inst = 32'd203423744;
      32330: inst = 32'd471859200;
      32331: inst = 32'd136314880;
      32332: inst = 32'd268468224;
      32333: inst = 32'd201343265;
      32334: inst = 32'd203423744;
      32335: inst = 32'd471859200;
      32336: inst = 32'd136314880;
      32337: inst = 32'd268468224;
      32338: inst = 32'd201343266;
      32339: inst = 32'd203423744;
      32340: inst = 32'd471859200;
      32341: inst = 32'd136314880;
      32342: inst = 32'd268468224;
      32343: inst = 32'd201343267;
      32344: inst = 32'd203423744;
      32345: inst = 32'd471859200;
      32346: inst = 32'd136314880;
      32347: inst = 32'd268468224;
      32348: inst = 32'd201343268;
      32349: inst = 32'd203423744;
      32350: inst = 32'd471859200;
      32351: inst = 32'd136314880;
      32352: inst = 32'd268468224;
      32353: inst = 32'd201343269;
      32354: inst = 32'd203423744;
      32355: inst = 32'd471859200;
      32356: inst = 32'd136314880;
      32357: inst = 32'd268468224;
      32358: inst = 32'd201343270;
      32359: inst = 32'd203423744;
      32360: inst = 32'd471859200;
      32361: inst = 32'd136314880;
      32362: inst = 32'd268468224;
      32363: inst = 32'd201343271;
      32364: inst = 32'd203423744;
      32365: inst = 32'd471859200;
      32366: inst = 32'd136314880;
      32367: inst = 32'd268468224;
      32368: inst = 32'd201343272;
      32369: inst = 32'd203423744;
      32370: inst = 32'd471859200;
      32371: inst = 32'd136314880;
      32372: inst = 32'd268468224;
      32373: inst = 32'd201343273;
      32374: inst = 32'd203423744;
      32375: inst = 32'd471859200;
      32376: inst = 32'd136314880;
      32377: inst = 32'd268468224;
      32378: inst = 32'd201343274;
      32379: inst = 32'd203423744;
      32380: inst = 32'd471859200;
      32381: inst = 32'd136314880;
      32382: inst = 32'd268468224;
      32383: inst = 32'd201343275;
      32384: inst = 32'd203423744;
      32385: inst = 32'd471859200;
      32386: inst = 32'd136314880;
      32387: inst = 32'd268468224;
      32388: inst = 32'd201343276;
      32389: inst = 32'd203423744;
      32390: inst = 32'd471859200;
      32391: inst = 32'd136314880;
      32392: inst = 32'd268468224;
      32393: inst = 32'd201343277;
      32394: inst = 32'd203423744;
      32395: inst = 32'd471859200;
      32396: inst = 32'd136314880;
      32397: inst = 32'd268468224;
      32398: inst = 32'd201343278;
      32399: inst = 32'd203423744;
      32400: inst = 32'd471859200;
      32401: inst = 32'd136314880;
      32402: inst = 32'd268468224;
      32403: inst = 32'd201343279;
      32404: inst = 32'd203423744;
      32405: inst = 32'd471859200;
      32406: inst = 32'd136314880;
      32407: inst = 32'd268468224;
      32408: inst = 32'd201343280;
      32409: inst = 32'd203423744;
      32410: inst = 32'd471859200;
      32411: inst = 32'd136314880;
      32412: inst = 32'd268468224;
      32413: inst = 32'd201343281;
      32414: inst = 32'd203423744;
      32415: inst = 32'd471859200;
      32416: inst = 32'd136314880;
      32417: inst = 32'd268468224;
      32418: inst = 32'd201343282;
      32419: inst = 32'd203423744;
      32420: inst = 32'd471859200;
      32421: inst = 32'd136314880;
      32422: inst = 32'd268468224;
      32423: inst = 32'd201343283;
      32424: inst = 32'd203423744;
      32425: inst = 32'd471859200;
      32426: inst = 32'd136314880;
      32427: inst = 32'd268468224;
      32428: inst = 32'd201343284;
      32429: inst = 32'd203423744;
      32430: inst = 32'd471859200;
      32431: inst = 32'd136314880;
      32432: inst = 32'd268468224;
      32433: inst = 32'd201343285;
      32434: inst = 32'd203423744;
      32435: inst = 32'd471859200;
      32436: inst = 32'd136314880;
      32437: inst = 32'd268468224;
      32438: inst = 32'd201343286;
      32439: inst = 32'd203423744;
      32440: inst = 32'd471859200;
      32441: inst = 32'd136314880;
      32442: inst = 32'd268468224;
      32443: inst = 32'd201343287;
      32444: inst = 32'd203423744;
      32445: inst = 32'd471859200;
      32446: inst = 32'd136314880;
      32447: inst = 32'd268468224;
      32448: inst = 32'd201343288;
      32449: inst = 32'd203423744;
      32450: inst = 32'd471859200;
      32451: inst = 32'd136314880;
      32452: inst = 32'd268468224;
      32453: inst = 32'd201343289;
      32454: inst = 32'd203423744;
      32455: inst = 32'd471859200;
      32456: inst = 32'd136314880;
      32457: inst = 32'd268468224;
      32458: inst = 32'd201343290;
      32459: inst = 32'd203423744;
      32460: inst = 32'd471859200;
      32461: inst = 32'd136314880;
      32462: inst = 32'd268468224;
      32463: inst = 32'd201343291;
      32464: inst = 32'd203423744;
      32465: inst = 32'd471859200;
      32466: inst = 32'd136314880;
      32467: inst = 32'd268468224;
      32468: inst = 32'd201343292;
      32469: inst = 32'd203423744;
      32470: inst = 32'd471859200;
      32471: inst = 32'd136314880;
      32472: inst = 32'd268468224;
      32473: inst = 32'd201343293;
      32474: inst = 32'd203423744;
      32475: inst = 32'd471859200;
      32476: inst = 32'd136314880;
      32477: inst = 32'd268468224;
      32478: inst = 32'd201343294;
      32479: inst = 32'd203423744;
      32480: inst = 32'd471859200;
      32481: inst = 32'd136314880;
      32482: inst = 32'd268468224;
      32483: inst = 32'd201343295;
      32484: inst = 32'd203423744;
      32485: inst = 32'd471859200;
      32486: inst = 32'd136314880;
      32487: inst = 32'd268468224;
      32488: inst = 32'd201343296;
      32489: inst = 32'd203423744;
      32490: inst = 32'd471859200;
      32491: inst = 32'd136314880;
      32492: inst = 32'd268468224;
      32493: inst = 32'd201343297;
      32494: inst = 32'd203423744;
      32495: inst = 32'd471859200;
      32496: inst = 32'd136314880;
      32497: inst = 32'd268468224;
      32498: inst = 32'd201343298;
      32499: inst = 32'd203423744;
      32500: inst = 32'd471859200;
      32501: inst = 32'd136314880;
      32502: inst = 32'd268468224;
      32503: inst = 32'd201343299;
      32504: inst = 32'd203423744;
      32505: inst = 32'd471859200;
      32506: inst = 32'd136314880;
      32507: inst = 32'd268468224;
      32508: inst = 32'd201343300;
      32509: inst = 32'd203423744;
      32510: inst = 32'd471859200;
      32511: inst = 32'd136314880;
      32512: inst = 32'd268468224;
      32513: inst = 32'd201343301;
      32514: inst = 32'd203423744;
      32515: inst = 32'd471859200;
      32516: inst = 32'd136314880;
      32517: inst = 32'd268468224;
      32518: inst = 32'd201343302;
      32519: inst = 32'd203423744;
      32520: inst = 32'd471859200;
      32521: inst = 32'd136314880;
      32522: inst = 32'd268468224;
      32523: inst = 32'd201343303;
      32524: inst = 32'd203423744;
      32525: inst = 32'd471859200;
      32526: inst = 32'd136314880;
      32527: inst = 32'd268468224;
      32528: inst = 32'd201343304;
      32529: inst = 32'd203423744;
      32530: inst = 32'd471859200;
      32531: inst = 32'd136314880;
      32532: inst = 32'd268468224;
      32533: inst = 32'd201343305;
      32534: inst = 32'd203423744;
      32535: inst = 32'd471859200;
      32536: inst = 32'd136314880;
      32537: inst = 32'd268468224;
      32538: inst = 32'd201343306;
      32539: inst = 32'd203423744;
      32540: inst = 32'd471859200;
      32541: inst = 32'd136314880;
      32542: inst = 32'd268468224;
      32543: inst = 32'd201343307;
      32544: inst = 32'd203423744;
      32545: inst = 32'd471859200;
      32546: inst = 32'd136314880;
      32547: inst = 32'd268468224;
      32548: inst = 32'd201343308;
      32549: inst = 32'd203423744;
      32550: inst = 32'd471859200;
      32551: inst = 32'd136314880;
      32552: inst = 32'd268468224;
      32553: inst = 32'd201343309;
      32554: inst = 32'd203423744;
      32555: inst = 32'd471859200;
      32556: inst = 32'd136314880;
      32557: inst = 32'd268468224;
      32558: inst = 32'd201343310;
      32559: inst = 32'd203423744;
      32560: inst = 32'd471859200;
      32561: inst = 32'd136314880;
      32562: inst = 32'd268468224;
      32563: inst = 32'd201343311;
      32564: inst = 32'd203423744;
      32565: inst = 32'd471859200;
      32566: inst = 32'd136314880;
      32567: inst = 32'd268468224;
      32568: inst = 32'd201343312;
      32569: inst = 32'd203423744;
      32570: inst = 32'd471859200;
      32571: inst = 32'd136314880;
      32572: inst = 32'd268468224;
      32573: inst = 32'd201343313;
      32574: inst = 32'd203423744;
      32575: inst = 32'd471859200;
      32576: inst = 32'd136314880;
      32577: inst = 32'd268468224;
      32578: inst = 32'd201343314;
      32579: inst = 32'd203423744;
      32580: inst = 32'd471859200;
      32581: inst = 32'd136314880;
      32582: inst = 32'd268468224;
      32583: inst = 32'd201343315;
      32584: inst = 32'd203423744;
      32585: inst = 32'd471859200;
      32586: inst = 32'd136314880;
      32587: inst = 32'd268468224;
      32588: inst = 32'd201343316;
      32589: inst = 32'd203423744;
      32590: inst = 32'd471859200;
      32591: inst = 32'd136314880;
      32592: inst = 32'd268468224;
      32593: inst = 32'd201343317;
      32594: inst = 32'd203423744;
      32595: inst = 32'd471859200;
      32596: inst = 32'd136314880;
      32597: inst = 32'd268468224;
      32598: inst = 32'd201343318;
      32599: inst = 32'd203423744;
      32600: inst = 32'd471859200;
      32601: inst = 32'd136314880;
      32602: inst = 32'd268468224;
      32603: inst = 32'd201343319;
      32604: inst = 32'd203423744;
      32605: inst = 32'd471859200;
      32606: inst = 32'd136314880;
      32607: inst = 32'd268468224;
      32608: inst = 32'd201343320;
      32609: inst = 32'd203423744;
      32610: inst = 32'd471859200;
      32611: inst = 32'd136314880;
      32612: inst = 32'd268468224;
      32613: inst = 32'd201343321;
      32614: inst = 32'd203423744;
      32615: inst = 32'd471859200;
      32616: inst = 32'd136314880;
      32617: inst = 32'd268468224;
      32618: inst = 32'd201343322;
      32619: inst = 32'd203423744;
      32620: inst = 32'd471859200;
      32621: inst = 32'd136314880;
      32622: inst = 32'd268468224;
      32623: inst = 32'd201343323;
      32624: inst = 32'd203423744;
      32625: inst = 32'd471859200;
      32626: inst = 32'd136314880;
      32627: inst = 32'd268468224;
      32628: inst = 32'd201343324;
      32629: inst = 32'd203423744;
      32630: inst = 32'd471859200;
      32631: inst = 32'd136314880;
      32632: inst = 32'd268468224;
      32633: inst = 32'd201343325;
      32634: inst = 32'd203423744;
      32635: inst = 32'd471859200;
      32636: inst = 32'd136314880;
      32637: inst = 32'd268468224;
      32638: inst = 32'd201343326;
      32639: inst = 32'd203423744;
      32640: inst = 32'd471859200;
      32641: inst = 32'd136314880;
      32642: inst = 32'd268468224;
      32643: inst = 32'd201343327;
      32644: inst = 32'd203423744;
      32645: inst = 32'd471859200;
      32646: inst = 32'd136314880;
      32647: inst = 32'd268468224;
      32648: inst = 32'd201343328;
      32649: inst = 32'd203423744;
      32650: inst = 32'd471859200;
      32651: inst = 32'd136314880;
      32652: inst = 32'd268468224;
      32653: inst = 32'd201343329;
      32654: inst = 32'd203423744;
      32655: inst = 32'd471859200;
      32656: inst = 32'd136314880;
      32657: inst = 32'd268468224;
      32658: inst = 32'd201343330;
      32659: inst = 32'd203423744;
      32660: inst = 32'd471859200;
      32661: inst = 32'd136314880;
      32662: inst = 32'd268468224;
      32663: inst = 32'd201343331;
      32664: inst = 32'd203423744;
      32665: inst = 32'd471859200;
      32666: inst = 32'd136314880;
      32667: inst = 32'd268468224;
      32668: inst = 32'd201343332;
      32669: inst = 32'd203423744;
      32670: inst = 32'd471859200;
      32671: inst = 32'd136314880;
      32672: inst = 32'd268468224;
      32673: inst = 32'd201343333;
      32674: inst = 32'd203423744;
      32675: inst = 32'd471859200;
      32676: inst = 32'd136314880;
      32677: inst = 32'd268468224;
      32678: inst = 32'd201343334;
      32679: inst = 32'd203423744;
      32680: inst = 32'd471859200;
      32681: inst = 32'd136314880;
      32682: inst = 32'd268468224;
      32683: inst = 32'd201343335;
      32684: inst = 32'd203423744;
      32685: inst = 32'd471859200;
      32686: inst = 32'd136314880;
      32687: inst = 32'd268468224;
      32688: inst = 32'd201343336;
      32689: inst = 32'd203423744;
      32690: inst = 32'd471859200;
      32691: inst = 32'd136314880;
      32692: inst = 32'd268468224;
      32693: inst = 32'd201343337;
      32694: inst = 32'd203423744;
      32695: inst = 32'd471859200;
      32696: inst = 32'd136314880;
      32697: inst = 32'd268468224;
      32698: inst = 32'd201343338;
      32699: inst = 32'd203423744;
      32700: inst = 32'd471859200;
      32701: inst = 32'd136314880;
      32702: inst = 32'd268468224;
      32703: inst = 32'd201343339;
      32704: inst = 32'd203423744;
      32705: inst = 32'd471859200;
      32706: inst = 32'd136314880;
      32707: inst = 32'd268468224;
      32708: inst = 32'd201343340;
      32709: inst = 32'd203423744;
      32710: inst = 32'd471859200;
      32711: inst = 32'd136314880;
      32712: inst = 32'd268468224;
      32713: inst = 32'd201343341;
      32714: inst = 32'd203423744;
      32715: inst = 32'd471859200;
      32716: inst = 32'd136314880;
      32717: inst = 32'd268468224;
      32718: inst = 32'd201343342;
      32719: inst = 32'd203423744;
      32720: inst = 32'd471859200;
      32721: inst = 32'd136314880;
      32722: inst = 32'd268468224;
      32723: inst = 32'd201343343;
      32724: inst = 32'd203423744;
      32725: inst = 32'd471859200;
      32726: inst = 32'd136314880;
      32727: inst = 32'd268468224;
      32728: inst = 32'd201343344;
      32729: inst = 32'd203423744;
      32730: inst = 32'd471859200;
      32731: inst = 32'd136314880;
      32732: inst = 32'd268468224;
      32733: inst = 32'd201343345;
      32734: inst = 32'd203423744;
      32735: inst = 32'd471859200;
      32736: inst = 32'd136314880;
      32737: inst = 32'd268468224;
      32738: inst = 32'd201343346;
      32739: inst = 32'd203423744;
      32740: inst = 32'd471859200;
      32741: inst = 32'd136314880;
      32742: inst = 32'd268468224;
      32743: inst = 32'd201343347;
      32744: inst = 32'd203423744;
      32745: inst = 32'd471859200;
      32746: inst = 32'd136314880;
      32747: inst = 32'd268468224;
      32748: inst = 32'd201343348;
      32749: inst = 32'd203423744;
      32750: inst = 32'd471859200;
      32751: inst = 32'd136314880;
      32752: inst = 32'd268468224;
      32753: inst = 32'd201343349;
      32754: inst = 32'd203423744;
      32755: inst = 32'd471859200;
      32756: inst = 32'd136314880;
      32757: inst = 32'd268468224;
      32758: inst = 32'd201343350;
      32759: inst = 32'd203423744;
      32760: inst = 32'd471859200;
      32761: inst = 32'd136314880;
      32762: inst = 32'd268468224;
      32763: inst = 32'd201343351;
      32764: inst = 32'd203423744;
      32765: inst = 32'd471859200;
      32766: inst = 32'd136314880;
      32767: inst = 32'd268468224;
      32768: inst = 32'd201343352;
      32769: inst = 32'd203423744;
      32770: inst = 32'd471859200;
      32771: inst = 32'd136314880;
      32772: inst = 32'd268468224;
      32773: inst = 32'd201343353;
      32774: inst = 32'd203423744;
      32775: inst = 32'd471859200;
      32776: inst = 32'd136314880;
      32777: inst = 32'd268468224;
      32778: inst = 32'd201343354;
      32779: inst = 32'd203423744;
      32780: inst = 32'd471859200;
      32781: inst = 32'd136314880;
      32782: inst = 32'd268468224;
      32783: inst = 32'd201343355;
      32784: inst = 32'd203423744;
      32785: inst = 32'd471859200;
      32786: inst = 32'd136314880;
      32787: inst = 32'd268468224;
      32788: inst = 32'd201343356;
      32789: inst = 32'd203423744;
      32790: inst = 32'd471859200;
      32791: inst = 32'd136314880;
      32792: inst = 32'd268468224;
      32793: inst = 32'd201343357;
      32794: inst = 32'd203423744;
      32795: inst = 32'd471859200;
      32796: inst = 32'd136314880;
      32797: inst = 32'd268468224;
      32798: inst = 32'd201343358;
      32799: inst = 32'd203423744;
      32800: inst = 32'd471859200;
      32801: inst = 32'd136314880;
      32802: inst = 32'd268468224;
      32803: inst = 32'd201343359;
      32804: inst = 32'd203423744;
      32805: inst = 32'd471859200;
      32806: inst = 32'd136314880;
      32807: inst = 32'd268468224;
      32808: inst = 32'd201343360;
      32809: inst = 32'd203423744;
      32810: inst = 32'd471859200;
      32811: inst = 32'd136314880;
      32812: inst = 32'd268468224;
      32813: inst = 32'd201343361;
      32814: inst = 32'd203423744;
      32815: inst = 32'd471859200;
      32816: inst = 32'd136314880;
      32817: inst = 32'd268468224;
      32818: inst = 32'd201343362;
      32819: inst = 32'd203423744;
      32820: inst = 32'd471859200;
      32821: inst = 32'd136314880;
      32822: inst = 32'd268468224;
      32823: inst = 32'd201343363;
      32824: inst = 32'd203423744;
      32825: inst = 32'd471859200;
      32826: inst = 32'd136314880;
      32827: inst = 32'd268468224;
      32828: inst = 32'd201343364;
      32829: inst = 32'd203423744;
      32830: inst = 32'd471859200;
      32831: inst = 32'd136314880;
      32832: inst = 32'd268468224;
      32833: inst = 32'd201343365;
      32834: inst = 32'd203423744;
      32835: inst = 32'd471859200;
      32836: inst = 32'd136314880;
      32837: inst = 32'd268468224;
      32838: inst = 32'd201343366;
      32839: inst = 32'd203423744;
      32840: inst = 32'd471859200;
      32841: inst = 32'd136314880;
      32842: inst = 32'd268468224;
      32843: inst = 32'd201343367;
      32844: inst = 32'd203423744;
      32845: inst = 32'd471859200;
      32846: inst = 32'd136314880;
      32847: inst = 32'd268468224;
      32848: inst = 32'd201343368;
      32849: inst = 32'd203423744;
      32850: inst = 32'd471859200;
      32851: inst = 32'd136314880;
      32852: inst = 32'd268468224;
      32853: inst = 32'd201343369;
      32854: inst = 32'd203423744;
      32855: inst = 32'd471859200;
      32856: inst = 32'd136314880;
      32857: inst = 32'd268468224;
      32858: inst = 32'd201343370;
      32859: inst = 32'd203423744;
      32860: inst = 32'd471859200;
      32861: inst = 32'd136314880;
      32862: inst = 32'd268468224;
      32863: inst = 32'd201343371;
      32864: inst = 32'd203423744;
      32865: inst = 32'd471859200;
      32866: inst = 32'd136314880;
      32867: inst = 32'd268468224;
      32868: inst = 32'd201343372;
      32869: inst = 32'd203423744;
      32870: inst = 32'd471859200;
      32871: inst = 32'd136314880;
      32872: inst = 32'd268468224;
      32873: inst = 32'd201343373;
      32874: inst = 32'd203423744;
      32875: inst = 32'd471859200;
      32876: inst = 32'd136314880;
      32877: inst = 32'd268468224;
      32878: inst = 32'd201343374;
      32879: inst = 32'd203423744;
      32880: inst = 32'd471859200;
      32881: inst = 32'd136314880;
      32882: inst = 32'd268468224;
      32883: inst = 32'd201343375;
      32884: inst = 32'd203423744;
      32885: inst = 32'd471859200;
      32886: inst = 32'd136314880;
      32887: inst = 32'd268468224;
      32888: inst = 32'd201343376;
      32889: inst = 32'd203423744;
      32890: inst = 32'd471859200;
      32891: inst = 32'd136314880;
      32892: inst = 32'd268468224;
      32893: inst = 32'd201343377;
      32894: inst = 32'd203423744;
      32895: inst = 32'd471859200;
      32896: inst = 32'd136314880;
      32897: inst = 32'd268468224;
      32898: inst = 32'd201343378;
      32899: inst = 32'd203423744;
      32900: inst = 32'd471859200;
      32901: inst = 32'd136314880;
      32902: inst = 32'd268468224;
      32903: inst = 32'd201343379;
      32904: inst = 32'd203423744;
      32905: inst = 32'd471859200;
      32906: inst = 32'd136314880;
      32907: inst = 32'd268468224;
      32908: inst = 32'd201343380;
      32909: inst = 32'd203423744;
      32910: inst = 32'd471859200;
      32911: inst = 32'd136314880;
      32912: inst = 32'd268468224;
      32913: inst = 32'd201343381;
      32914: inst = 32'd203423744;
      32915: inst = 32'd471859200;
      32916: inst = 32'd136314880;
      32917: inst = 32'd268468224;
      32918: inst = 32'd201343382;
      32919: inst = 32'd203423744;
      32920: inst = 32'd471859200;
      32921: inst = 32'd136314880;
      32922: inst = 32'd268468224;
      32923: inst = 32'd201343383;
      32924: inst = 32'd203423744;
      32925: inst = 32'd471859200;
      32926: inst = 32'd136314880;
      32927: inst = 32'd268468224;
      32928: inst = 32'd201343384;
      32929: inst = 32'd203423744;
      32930: inst = 32'd471859200;
      32931: inst = 32'd136314880;
      32932: inst = 32'd268468224;
      32933: inst = 32'd201343385;
      32934: inst = 32'd203423744;
      32935: inst = 32'd471859200;
      32936: inst = 32'd136314880;
      32937: inst = 32'd268468224;
      32938: inst = 32'd201343386;
      32939: inst = 32'd203423744;
      32940: inst = 32'd471859200;
      32941: inst = 32'd136314880;
      32942: inst = 32'd268468224;
      32943: inst = 32'd201343387;
      32944: inst = 32'd203423744;
      32945: inst = 32'd471859200;
      32946: inst = 32'd136314880;
      32947: inst = 32'd268468224;
      32948: inst = 32'd201343388;
      32949: inst = 32'd203423744;
      32950: inst = 32'd471859200;
      32951: inst = 32'd136314880;
      32952: inst = 32'd268468224;
      32953: inst = 32'd201343389;
      32954: inst = 32'd203423744;
      32955: inst = 32'd471859200;
      32956: inst = 32'd136314880;
      32957: inst = 32'd268468224;
      32958: inst = 32'd201343390;
      32959: inst = 32'd203423744;
      32960: inst = 32'd471859200;
      32961: inst = 32'd136314880;
      32962: inst = 32'd268468224;
      32963: inst = 32'd201343391;
      32964: inst = 32'd203423744;
      32965: inst = 32'd471859200;
      32966: inst = 32'd136314880;
      32967: inst = 32'd268468224;
      32968: inst = 32'd201343392;
      32969: inst = 32'd203423744;
      32970: inst = 32'd471859200;
      32971: inst = 32'd136314880;
      32972: inst = 32'd268468224;
      32973: inst = 32'd201343393;
      32974: inst = 32'd203423744;
      32975: inst = 32'd471859200;
      32976: inst = 32'd136314880;
      32977: inst = 32'd268468224;
      32978: inst = 32'd201343394;
      32979: inst = 32'd203423744;
      32980: inst = 32'd471859200;
      32981: inst = 32'd136314880;
      32982: inst = 32'd268468224;
      32983: inst = 32'd201343395;
      32984: inst = 32'd203423744;
      32985: inst = 32'd471859200;
      32986: inst = 32'd136314880;
      32987: inst = 32'd268468224;
      32988: inst = 32'd201343396;
      32989: inst = 32'd203423744;
      32990: inst = 32'd471859200;
      32991: inst = 32'd136314880;
      32992: inst = 32'd268468224;
      32993: inst = 32'd201343397;
      32994: inst = 32'd203423744;
      32995: inst = 32'd471859200;
      32996: inst = 32'd136314880;
      32997: inst = 32'd268468224;
      32998: inst = 32'd201343398;
      32999: inst = 32'd203423744;
      33000: inst = 32'd471859200;
      33001: inst = 32'd136314880;
      33002: inst = 32'd268468224;
      33003: inst = 32'd201343399;
      33004: inst = 32'd203423744;
      33005: inst = 32'd471859200;
      33006: inst = 32'd136314880;
      33007: inst = 32'd268468224;
      33008: inst = 32'd201343400;
      33009: inst = 32'd203423744;
      33010: inst = 32'd471859200;
      33011: inst = 32'd136314880;
      33012: inst = 32'd268468224;
      33013: inst = 32'd201343401;
      33014: inst = 32'd203423744;
      33015: inst = 32'd471859200;
      33016: inst = 32'd136314880;
      33017: inst = 32'd268468224;
      33018: inst = 32'd201343402;
      33019: inst = 32'd203423744;
      33020: inst = 32'd471859200;
      33021: inst = 32'd136314880;
      33022: inst = 32'd268468224;
      33023: inst = 32'd201343403;
      33024: inst = 32'd203423744;
      33025: inst = 32'd471859200;
      33026: inst = 32'd136314880;
      33027: inst = 32'd268468224;
      33028: inst = 32'd201343404;
      33029: inst = 32'd203423744;
      33030: inst = 32'd471859200;
      33031: inst = 32'd136314880;
      33032: inst = 32'd268468224;
      33033: inst = 32'd201343405;
      33034: inst = 32'd203423744;
      33035: inst = 32'd471859200;
      33036: inst = 32'd136314880;
      33037: inst = 32'd268468224;
      33038: inst = 32'd201343406;
      33039: inst = 32'd203423744;
      33040: inst = 32'd471859200;
      33041: inst = 32'd136314880;
      33042: inst = 32'd268468224;
      33043: inst = 32'd201343407;
      33044: inst = 32'd203423744;
      33045: inst = 32'd471859200;
      33046: inst = 32'd136314880;
      33047: inst = 32'd268468224;
      33048: inst = 32'd201343408;
      33049: inst = 32'd203423744;
      33050: inst = 32'd471859200;
      33051: inst = 32'd136314880;
      33052: inst = 32'd268468224;
      33053: inst = 32'd201343409;
      33054: inst = 32'd203423744;
      33055: inst = 32'd471859200;
      33056: inst = 32'd136314880;
      33057: inst = 32'd268468224;
      33058: inst = 32'd201343410;
      33059: inst = 32'd203423744;
      33060: inst = 32'd471859200;
      33061: inst = 32'd136314880;
      33062: inst = 32'd268468224;
      33063: inst = 32'd201343411;
      33064: inst = 32'd203423744;
      33065: inst = 32'd471859200;
      33066: inst = 32'd136314880;
      33067: inst = 32'd268468224;
      33068: inst = 32'd201343412;
      33069: inst = 32'd203423744;
      33070: inst = 32'd471859200;
      33071: inst = 32'd136314880;
      33072: inst = 32'd268468224;
      33073: inst = 32'd201343413;
      33074: inst = 32'd203423744;
      33075: inst = 32'd471859200;
      33076: inst = 32'd136314880;
      33077: inst = 32'd268468224;
      33078: inst = 32'd201343414;
      33079: inst = 32'd203423744;
      33080: inst = 32'd471859200;
      33081: inst = 32'd136314880;
      33082: inst = 32'd268468224;
      33083: inst = 32'd201343415;
      33084: inst = 32'd203423744;
      33085: inst = 32'd471859200;
      33086: inst = 32'd136314880;
      33087: inst = 32'd268468224;
      33088: inst = 32'd201343416;
      33089: inst = 32'd203423744;
      33090: inst = 32'd471859200;
      33091: inst = 32'd136314880;
      33092: inst = 32'd268468224;
      33093: inst = 32'd201343417;
      33094: inst = 32'd203423744;
      33095: inst = 32'd471859200;
      33096: inst = 32'd136314880;
      33097: inst = 32'd268468224;
      33098: inst = 32'd201343418;
      33099: inst = 32'd203423744;
      33100: inst = 32'd471859200;
      33101: inst = 32'd136314880;
      33102: inst = 32'd268468224;
      33103: inst = 32'd201343419;
      33104: inst = 32'd203423744;
      33105: inst = 32'd471859200;
      33106: inst = 32'd136314880;
      33107: inst = 32'd268468224;
      33108: inst = 32'd201343420;
      33109: inst = 32'd203423744;
      33110: inst = 32'd471859200;
      33111: inst = 32'd136314880;
      33112: inst = 32'd268468224;
      33113: inst = 32'd201343421;
      33114: inst = 32'd203423744;
      33115: inst = 32'd471859200;
      33116: inst = 32'd136314880;
      33117: inst = 32'd268468224;
      33118: inst = 32'd201343422;
      33119: inst = 32'd203423744;
      33120: inst = 32'd471859200;
      33121: inst = 32'd136314880;
      33122: inst = 32'd268468224;
      33123: inst = 32'd201343423;
      33124: inst = 32'd203423744;
      33125: inst = 32'd471859200;
      33126: inst = 32'd136314880;
      33127: inst = 32'd268468224;
      33128: inst = 32'd201343424;
      33129: inst = 32'd203423744;
      33130: inst = 32'd471859200;
      33131: inst = 32'd136314880;
      33132: inst = 32'd268468224;
      33133: inst = 32'd201343425;
      33134: inst = 32'd203423744;
      33135: inst = 32'd471859200;
      33136: inst = 32'd136314880;
      33137: inst = 32'd268468224;
      33138: inst = 32'd201343426;
      33139: inst = 32'd203423744;
      33140: inst = 32'd471859200;
      33141: inst = 32'd136314880;
      33142: inst = 32'd268468224;
      33143: inst = 32'd201343427;
      33144: inst = 32'd203423744;
      33145: inst = 32'd471859200;
      33146: inst = 32'd136314880;
      33147: inst = 32'd268468224;
      33148: inst = 32'd201343428;
      33149: inst = 32'd203423744;
      33150: inst = 32'd471859200;
      33151: inst = 32'd136314880;
      33152: inst = 32'd268468224;
      33153: inst = 32'd201343429;
      33154: inst = 32'd203423744;
      33155: inst = 32'd471859200;
      33156: inst = 32'd136314880;
      33157: inst = 32'd268468224;
      33158: inst = 32'd201343430;
      33159: inst = 32'd203423744;
      33160: inst = 32'd471859200;
      33161: inst = 32'd136314880;
      33162: inst = 32'd268468224;
      33163: inst = 32'd201343431;
      33164: inst = 32'd203423744;
      33165: inst = 32'd471859200;
      33166: inst = 32'd136314880;
      33167: inst = 32'd268468224;
      33168: inst = 32'd201343432;
      33169: inst = 32'd203423744;
      33170: inst = 32'd471859200;
      33171: inst = 32'd136314880;
      33172: inst = 32'd268468224;
      33173: inst = 32'd201343433;
      33174: inst = 32'd203423744;
      33175: inst = 32'd471859200;
      33176: inst = 32'd136314880;
      33177: inst = 32'd268468224;
      33178: inst = 32'd201343434;
      33179: inst = 32'd203423744;
      33180: inst = 32'd471859200;
      33181: inst = 32'd136314880;
      33182: inst = 32'd268468224;
      33183: inst = 32'd201343435;
      33184: inst = 32'd203423744;
      33185: inst = 32'd471859200;
      33186: inst = 32'd136314880;
      33187: inst = 32'd268468224;
      33188: inst = 32'd201343436;
      33189: inst = 32'd203423744;
      33190: inst = 32'd471859200;
      33191: inst = 32'd136314880;
      33192: inst = 32'd268468224;
      33193: inst = 32'd201343437;
      33194: inst = 32'd203423744;
      33195: inst = 32'd471859200;
      33196: inst = 32'd136314880;
      33197: inst = 32'd268468224;
      33198: inst = 32'd201343438;
      33199: inst = 32'd203423744;
      33200: inst = 32'd471859200;
      33201: inst = 32'd136314880;
      33202: inst = 32'd268468224;
      33203: inst = 32'd201343439;
      33204: inst = 32'd203423744;
      33205: inst = 32'd471859200;
      33206: inst = 32'd136314880;
      33207: inst = 32'd268468224;
      33208: inst = 32'd201343440;
      33209: inst = 32'd203423744;
      33210: inst = 32'd471859200;
      33211: inst = 32'd136314880;
      33212: inst = 32'd268468224;
      33213: inst = 32'd201343441;
      33214: inst = 32'd203423744;
      33215: inst = 32'd471859200;
      33216: inst = 32'd136314880;
      33217: inst = 32'd268468224;
      33218: inst = 32'd201343442;
      33219: inst = 32'd203423744;
      33220: inst = 32'd471859200;
      33221: inst = 32'd136314880;
      33222: inst = 32'd268468224;
      33223: inst = 32'd201343443;
      33224: inst = 32'd203423744;
      33225: inst = 32'd471859200;
      33226: inst = 32'd136314880;
      33227: inst = 32'd268468224;
      33228: inst = 32'd201343444;
      33229: inst = 32'd203423744;
      33230: inst = 32'd471859200;
      33231: inst = 32'd136314880;
      33232: inst = 32'd268468224;
      33233: inst = 32'd201343445;
      33234: inst = 32'd203423744;
      33235: inst = 32'd471859200;
      33236: inst = 32'd136314880;
      33237: inst = 32'd268468224;
      33238: inst = 32'd201343446;
      33239: inst = 32'd203423744;
      33240: inst = 32'd471859200;
      33241: inst = 32'd136314880;
      33242: inst = 32'd268468224;
      33243: inst = 32'd201343447;
      33244: inst = 32'd203423744;
      33245: inst = 32'd471859200;
      33246: inst = 32'd136314880;
      33247: inst = 32'd268468224;
      33248: inst = 32'd201343448;
      33249: inst = 32'd203423744;
      33250: inst = 32'd471859200;
      33251: inst = 32'd136314880;
      33252: inst = 32'd268468224;
      33253: inst = 32'd201343449;
      33254: inst = 32'd203423744;
      33255: inst = 32'd471859200;
      33256: inst = 32'd136314880;
      33257: inst = 32'd268468224;
      33258: inst = 32'd201343450;
      33259: inst = 32'd203423744;
      33260: inst = 32'd471859200;
      33261: inst = 32'd136314880;
      33262: inst = 32'd268468224;
      33263: inst = 32'd201343451;
      33264: inst = 32'd203423744;
      33265: inst = 32'd471859200;
      33266: inst = 32'd136314880;
      33267: inst = 32'd268468224;
      33268: inst = 32'd201343452;
      33269: inst = 32'd203423744;
      33270: inst = 32'd471859200;
      33271: inst = 32'd136314880;
      33272: inst = 32'd268468224;
      33273: inst = 32'd201343453;
      33274: inst = 32'd203423744;
      33275: inst = 32'd471859200;
      33276: inst = 32'd136314880;
      33277: inst = 32'd268468224;
      33278: inst = 32'd201343454;
      33279: inst = 32'd203423744;
      33280: inst = 32'd471859200;
      33281: inst = 32'd136314880;
      33282: inst = 32'd268468224;
      33283: inst = 32'd201343455;
      33284: inst = 32'd203423744;
      33285: inst = 32'd471859200;
      33286: inst = 32'd136314880;
      33287: inst = 32'd268468224;
      33288: inst = 32'd201343456;
      33289: inst = 32'd203423744;
      33290: inst = 32'd471859200;
      33291: inst = 32'd136314880;
      33292: inst = 32'd268468224;
      33293: inst = 32'd201343457;
      33294: inst = 32'd203423744;
      33295: inst = 32'd471859200;
      33296: inst = 32'd136314880;
      33297: inst = 32'd268468224;
      33298: inst = 32'd201343458;
      33299: inst = 32'd203423744;
      33300: inst = 32'd471859200;
      33301: inst = 32'd136314880;
      33302: inst = 32'd268468224;
      33303: inst = 32'd201343459;
      33304: inst = 32'd203423744;
      33305: inst = 32'd471859200;
      33306: inst = 32'd136314880;
      33307: inst = 32'd268468224;
      33308: inst = 32'd201343460;
      33309: inst = 32'd203423744;
      33310: inst = 32'd471859200;
      33311: inst = 32'd136314880;
      33312: inst = 32'd268468224;
      33313: inst = 32'd201343461;
      33314: inst = 32'd203423744;
      33315: inst = 32'd471859200;
      33316: inst = 32'd136314880;
      33317: inst = 32'd268468224;
      33318: inst = 32'd201343462;
      33319: inst = 32'd203423744;
      33320: inst = 32'd471859200;
      33321: inst = 32'd136314880;
      33322: inst = 32'd268468224;
      33323: inst = 32'd201343463;
      33324: inst = 32'd203423744;
      33325: inst = 32'd471859200;
      33326: inst = 32'd136314880;
      33327: inst = 32'd268468224;
      33328: inst = 32'd201343464;
      33329: inst = 32'd203423744;
      33330: inst = 32'd471859200;
      33331: inst = 32'd136314880;
      33332: inst = 32'd268468224;
      33333: inst = 32'd201343465;
      33334: inst = 32'd203423744;
      33335: inst = 32'd471859200;
      33336: inst = 32'd136314880;
      33337: inst = 32'd268468224;
      33338: inst = 32'd201343466;
      33339: inst = 32'd203423744;
      33340: inst = 32'd471859200;
      33341: inst = 32'd136314880;
      33342: inst = 32'd268468224;
      33343: inst = 32'd201343467;
      33344: inst = 32'd203423744;
      33345: inst = 32'd471859200;
      33346: inst = 32'd136314880;
      33347: inst = 32'd268468224;
      33348: inst = 32'd201343468;
      33349: inst = 32'd203423744;
      33350: inst = 32'd471859200;
      33351: inst = 32'd136314880;
      33352: inst = 32'd268468224;
      33353: inst = 32'd201343469;
      33354: inst = 32'd203423744;
      33355: inst = 32'd471859200;
      33356: inst = 32'd136314880;
      33357: inst = 32'd268468224;
      33358: inst = 32'd201343470;
      33359: inst = 32'd203423744;
      33360: inst = 32'd471859200;
      33361: inst = 32'd136314880;
      33362: inst = 32'd268468224;
      33363: inst = 32'd201343471;
      33364: inst = 32'd203423744;
      33365: inst = 32'd471859200;
      33366: inst = 32'd136314880;
      33367: inst = 32'd268468224;
      33368: inst = 32'd201343472;
      33369: inst = 32'd203423744;
      33370: inst = 32'd471859200;
      33371: inst = 32'd136314880;
      33372: inst = 32'd268468224;
      33373: inst = 32'd201343473;
      33374: inst = 32'd203423744;
      33375: inst = 32'd471859200;
      33376: inst = 32'd136314880;
      33377: inst = 32'd268468224;
      33378: inst = 32'd201343474;
      33379: inst = 32'd203423744;
      33380: inst = 32'd471859200;
      33381: inst = 32'd136314880;
      33382: inst = 32'd268468224;
      33383: inst = 32'd201343475;
      33384: inst = 32'd203423744;
      33385: inst = 32'd471859200;
      33386: inst = 32'd136314880;
      33387: inst = 32'd268468224;
      33388: inst = 32'd201343476;
      33389: inst = 32'd203423744;
      33390: inst = 32'd471859200;
      33391: inst = 32'd136314880;
      33392: inst = 32'd268468224;
      33393: inst = 32'd201343477;
      33394: inst = 32'd203423744;
      33395: inst = 32'd471859200;
      33396: inst = 32'd136314880;
      33397: inst = 32'd268468224;
      33398: inst = 32'd201343478;
      33399: inst = 32'd203423744;
      33400: inst = 32'd471859200;
      33401: inst = 32'd136314880;
      33402: inst = 32'd268468224;
      33403: inst = 32'd201343479;
      33404: inst = 32'd203423744;
      33405: inst = 32'd471859200;
      33406: inst = 32'd136314880;
      33407: inst = 32'd268468224;
      33408: inst = 32'd201343480;
      33409: inst = 32'd203423744;
      33410: inst = 32'd471859200;
      33411: inst = 32'd136314880;
      33412: inst = 32'd268468224;
      33413: inst = 32'd201343481;
      33414: inst = 32'd203423744;
      33415: inst = 32'd471859200;
      33416: inst = 32'd136314880;
      33417: inst = 32'd268468224;
      33418: inst = 32'd201343482;
      33419: inst = 32'd203423744;
      33420: inst = 32'd471859200;
      33421: inst = 32'd136314880;
      33422: inst = 32'd268468224;
      33423: inst = 32'd201343483;
      33424: inst = 32'd203423744;
      33425: inst = 32'd471859200;
      33426: inst = 32'd136314880;
      33427: inst = 32'd268468224;
      33428: inst = 32'd201343484;
      33429: inst = 32'd203423744;
      33430: inst = 32'd471859200;
      33431: inst = 32'd136314880;
      33432: inst = 32'd268468224;
      33433: inst = 32'd201343485;
      33434: inst = 32'd203423744;
      33435: inst = 32'd471859200;
      33436: inst = 32'd136314880;
      33437: inst = 32'd268468224;
      33438: inst = 32'd201343486;
      33439: inst = 32'd203423744;
      33440: inst = 32'd471859200;
      33441: inst = 32'd136314880;
      33442: inst = 32'd268468224;
      33443: inst = 32'd201343487;
      33444: inst = 32'd203423744;
      33445: inst = 32'd471859200;
      33446: inst = 32'd136314880;
      33447: inst = 32'd268468224;
      33448: inst = 32'd201343488;
      33449: inst = 32'd203423744;
      33450: inst = 32'd471859200;
      33451: inst = 32'd136314880;
      33452: inst = 32'd268468224;
      33453: inst = 32'd201343489;
      33454: inst = 32'd203423744;
      33455: inst = 32'd471859200;
      33456: inst = 32'd136314880;
      33457: inst = 32'd268468224;
      33458: inst = 32'd201343490;
      33459: inst = 32'd203423744;
      33460: inst = 32'd471859200;
      33461: inst = 32'd136314880;
      33462: inst = 32'd268468224;
      33463: inst = 32'd201343491;
      33464: inst = 32'd203423744;
      33465: inst = 32'd471859200;
      33466: inst = 32'd136314880;
      33467: inst = 32'd268468224;
      33468: inst = 32'd201343492;
      33469: inst = 32'd203423744;
      33470: inst = 32'd471859200;
      33471: inst = 32'd136314880;
      33472: inst = 32'd268468224;
      33473: inst = 32'd201343493;
      33474: inst = 32'd203423744;
      33475: inst = 32'd471859200;
      33476: inst = 32'd136314880;
      33477: inst = 32'd268468224;
      33478: inst = 32'd201343494;
      33479: inst = 32'd203423744;
      33480: inst = 32'd471859200;
      33481: inst = 32'd136314880;
      33482: inst = 32'd268468224;
      33483: inst = 32'd201343495;
      33484: inst = 32'd203423744;
      33485: inst = 32'd471859200;
      33486: inst = 32'd136314880;
      33487: inst = 32'd268468224;
      33488: inst = 32'd201343496;
      33489: inst = 32'd203423744;
      33490: inst = 32'd471859200;
      33491: inst = 32'd136314880;
      33492: inst = 32'd268468224;
      33493: inst = 32'd201343497;
      33494: inst = 32'd203423744;
      33495: inst = 32'd471859200;
      33496: inst = 32'd136314880;
      33497: inst = 32'd268468224;
      33498: inst = 32'd201343498;
      33499: inst = 32'd203423744;
      33500: inst = 32'd471859200;
      33501: inst = 32'd136314880;
      33502: inst = 32'd268468224;
      33503: inst = 32'd201343499;
      33504: inst = 32'd203423744;
      33505: inst = 32'd471859200;
      33506: inst = 32'd136314880;
      33507: inst = 32'd268468224;
      33508: inst = 32'd201343500;
      33509: inst = 32'd203423744;
      33510: inst = 32'd471859200;
      33511: inst = 32'd136314880;
      33512: inst = 32'd268468224;
      33513: inst = 32'd201343501;
      33514: inst = 32'd203423744;
      33515: inst = 32'd471859200;
      33516: inst = 32'd136314880;
      33517: inst = 32'd268468224;
      33518: inst = 32'd201343502;
      33519: inst = 32'd203423744;
      33520: inst = 32'd471859200;
      33521: inst = 32'd136314880;
      33522: inst = 32'd268468224;
      33523: inst = 32'd201343503;
      33524: inst = 32'd203423744;
      33525: inst = 32'd471859200;
      33526: inst = 32'd136314880;
      33527: inst = 32'd268468224;
      33528: inst = 32'd201343504;
      33529: inst = 32'd203423744;
      33530: inst = 32'd471859200;
      33531: inst = 32'd136314880;
      33532: inst = 32'd268468224;
      33533: inst = 32'd201343505;
      33534: inst = 32'd203423744;
      33535: inst = 32'd471859200;
      33536: inst = 32'd136314880;
      33537: inst = 32'd268468224;
      33538: inst = 32'd201343506;
      33539: inst = 32'd203423744;
      33540: inst = 32'd471859200;
      33541: inst = 32'd136314880;
      33542: inst = 32'd268468224;
      33543: inst = 32'd201343507;
      33544: inst = 32'd203423744;
      33545: inst = 32'd471859200;
      33546: inst = 32'd136314880;
      33547: inst = 32'd268468224;
      33548: inst = 32'd201343508;
      33549: inst = 32'd203423744;
      33550: inst = 32'd471859200;
      33551: inst = 32'd136314880;
      33552: inst = 32'd268468224;
      33553: inst = 32'd201343509;
      33554: inst = 32'd203423744;
      33555: inst = 32'd471859200;
      33556: inst = 32'd136314880;
      33557: inst = 32'd268468224;
      33558: inst = 32'd201343510;
      33559: inst = 32'd203423744;
      33560: inst = 32'd471859200;
      33561: inst = 32'd136314880;
      33562: inst = 32'd268468224;
      33563: inst = 32'd201343511;
      33564: inst = 32'd203423744;
      33565: inst = 32'd471859200;
      33566: inst = 32'd136314880;
      33567: inst = 32'd268468224;
      33568: inst = 32'd201343512;
      33569: inst = 32'd203423744;
      33570: inst = 32'd471859200;
      33571: inst = 32'd136314880;
      33572: inst = 32'd268468224;
      33573: inst = 32'd201343513;
      33574: inst = 32'd203423744;
      33575: inst = 32'd471859200;
      33576: inst = 32'd136314880;
      33577: inst = 32'd268468224;
      33578: inst = 32'd201343514;
      33579: inst = 32'd203423744;
      33580: inst = 32'd471859200;
      33581: inst = 32'd136314880;
      33582: inst = 32'd268468224;
      33583: inst = 32'd201343515;
      33584: inst = 32'd203423744;
      33585: inst = 32'd471859200;
      33586: inst = 32'd136314880;
      33587: inst = 32'd268468224;
      33588: inst = 32'd201343516;
      33589: inst = 32'd203423744;
      33590: inst = 32'd471859200;
      33591: inst = 32'd136314880;
      33592: inst = 32'd268468224;
      33593: inst = 32'd201343517;
      33594: inst = 32'd203423744;
      33595: inst = 32'd471859200;
      33596: inst = 32'd136314880;
      33597: inst = 32'd268468224;
      33598: inst = 32'd201343518;
      33599: inst = 32'd203423744;
      33600: inst = 32'd471859200;
      33601: inst = 32'd136314880;
      33602: inst = 32'd268468224;
      33603: inst = 32'd201343519;
      33604: inst = 32'd203423744;
      33605: inst = 32'd471859200;
      33606: inst = 32'd136314880;
      33607: inst = 32'd268468224;
      33608: inst = 32'd201343520;
      33609: inst = 32'd203423744;
      33610: inst = 32'd471859200;
      33611: inst = 32'd136314880;
      33612: inst = 32'd268468224;
      33613: inst = 32'd201343521;
      33614: inst = 32'd203423744;
      33615: inst = 32'd471859200;
      33616: inst = 32'd136314880;
      33617: inst = 32'd268468224;
      33618: inst = 32'd201343522;
      33619: inst = 32'd203423744;
      33620: inst = 32'd471859200;
      33621: inst = 32'd136314880;
      33622: inst = 32'd268468224;
      33623: inst = 32'd201343523;
      33624: inst = 32'd203423744;
      33625: inst = 32'd471859200;
      33626: inst = 32'd136314880;
      33627: inst = 32'd268468224;
      33628: inst = 32'd201343524;
      33629: inst = 32'd203423744;
      33630: inst = 32'd471859200;
      33631: inst = 32'd136314880;
      33632: inst = 32'd268468224;
      33633: inst = 32'd201343525;
      33634: inst = 32'd203423744;
      33635: inst = 32'd471859200;
      33636: inst = 32'd136314880;
      33637: inst = 32'd268468224;
      33638: inst = 32'd201343526;
      33639: inst = 32'd203423744;
      33640: inst = 32'd471859200;
      33641: inst = 32'd136314880;
      33642: inst = 32'd268468224;
      33643: inst = 32'd201343527;
      33644: inst = 32'd203423744;
      33645: inst = 32'd471859200;
      33646: inst = 32'd136314880;
      33647: inst = 32'd268468224;
      33648: inst = 32'd201343528;
      33649: inst = 32'd203423744;
      33650: inst = 32'd471859200;
      33651: inst = 32'd136314880;
      33652: inst = 32'd268468224;
      33653: inst = 32'd201343529;
      33654: inst = 32'd203423744;
      33655: inst = 32'd471859200;
      33656: inst = 32'd136314880;
      33657: inst = 32'd268468224;
      33658: inst = 32'd201343530;
      33659: inst = 32'd203423744;
      33660: inst = 32'd471859200;
      33661: inst = 32'd136314880;
      33662: inst = 32'd268468224;
      33663: inst = 32'd201343531;
      33664: inst = 32'd203423744;
      33665: inst = 32'd471859200;
      33666: inst = 32'd136314880;
      33667: inst = 32'd268468224;
      33668: inst = 32'd201343532;
      33669: inst = 32'd203423744;
      33670: inst = 32'd471859200;
      33671: inst = 32'd136314880;
      33672: inst = 32'd268468224;
      33673: inst = 32'd201343533;
      33674: inst = 32'd203423744;
      33675: inst = 32'd471859200;
      33676: inst = 32'd136314880;
      33677: inst = 32'd268468224;
      33678: inst = 32'd201343534;
      33679: inst = 32'd203423744;
      33680: inst = 32'd471859200;
      33681: inst = 32'd136314880;
      33682: inst = 32'd268468224;
      33683: inst = 32'd201343535;
      33684: inst = 32'd203423744;
      33685: inst = 32'd471859200;
      33686: inst = 32'd136314880;
      33687: inst = 32'd268468224;
      33688: inst = 32'd201343536;
      33689: inst = 32'd203423744;
      33690: inst = 32'd471859200;
      33691: inst = 32'd136314880;
      33692: inst = 32'd268468224;
      33693: inst = 32'd201343537;
      33694: inst = 32'd203423744;
      33695: inst = 32'd471859200;
      33696: inst = 32'd136314880;
      33697: inst = 32'd268468224;
      33698: inst = 32'd201343538;
      33699: inst = 32'd203423744;
      33700: inst = 32'd471859200;
      33701: inst = 32'd136314880;
      33702: inst = 32'd268468224;
      33703: inst = 32'd201343539;
      33704: inst = 32'd203423744;
      33705: inst = 32'd471859200;
      33706: inst = 32'd136314880;
      33707: inst = 32'd268468224;
      33708: inst = 32'd201343540;
      33709: inst = 32'd203423744;
      33710: inst = 32'd471859200;
      33711: inst = 32'd136314880;
      33712: inst = 32'd268468224;
      33713: inst = 32'd201343541;
      33714: inst = 32'd203423744;
      33715: inst = 32'd471859200;
      33716: inst = 32'd136314880;
      33717: inst = 32'd268468224;
      33718: inst = 32'd201343542;
      33719: inst = 32'd203423744;
      33720: inst = 32'd471859200;
      33721: inst = 32'd136314880;
      33722: inst = 32'd268468224;
      33723: inst = 32'd201343543;
      33724: inst = 32'd203423744;
      33725: inst = 32'd471859200;
      33726: inst = 32'd136314880;
      33727: inst = 32'd268468224;
      33728: inst = 32'd201343544;
      33729: inst = 32'd203423744;
      33730: inst = 32'd471859200;
      33731: inst = 32'd136314880;
      33732: inst = 32'd268468224;
      33733: inst = 32'd201343545;
      33734: inst = 32'd203423744;
      33735: inst = 32'd471859200;
      33736: inst = 32'd136314880;
      33737: inst = 32'd268468224;
      33738: inst = 32'd201343546;
      33739: inst = 32'd203423744;
      33740: inst = 32'd471859200;
      33741: inst = 32'd136314880;
      33742: inst = 32'd268468224;
      33743: inst = 32'd201343547;
      33744: inst = 32'd203423744;
      33745: inst = 32'd471859200;
      33746: inst = 32'd136314880;
      33747: inst = 32'd268468224;
      33748: inst = 32'd201343548;
      33749: inst = 32'd203423744;
      33750: inst = 32'd471859200;
      33751: inst = 32'd136314880;
      33752: inst = 32'd268468224;
      33753: inst = 32'd201343549;
      33754: inst = 32'd203423744;
      33755: inst = 32'd471859200;
      33756: inst = 32'd136314880;
      33757: inst = 32'd268468224;
      33758: inst = 32'd201343550;
      33759: inst = 32'd203423744;
      33760: inst = 32'd471859200;
      33761: inst = 32'd136314880;
      33762: inst = 32'd268468224;
      33763: inst = 32'd201343551;
      33764: inst = 32'd203423744;
      33765: inst = 32'd471859200;
      33766: inst = 32'd136314880;
      33767: inst = 32'd268468224;
      33768: inst = 32'd201343552;
      33769: inst = 32'd203423744;
      33770: inst = 32'd471859200;
      33771: inst = 32'd136314880;
      33772: inst = 32'd268468224;
      33773: inst = 32'd201343553;
      33774: inst = 32'd203423744;
      33775: inst = 32'd471859200;
      33776: inst = 32'd136314880;
      33777: inst = 32'd268468224;
      33778: inst = 32'd201343554;
      33779: inst = 32'd203423744;
      33780: inst = 32'd471859200;
      33781: inst = 32'd136314880;
      33782: inst = 32'd268468224;
      33783: inst = 32'd201343555;
      33784: inst = 32'd203423744;
      33785: inst = 32'd471859200;
      33786: inst = 32'd136314880;
      33787: inst = 32'd268468224;
      33788: inst = 32'd201343556;
      33789: inst = 32'd203423744;
      33790: inst = 32'd471859200;
      33791: inst = 32'd136314880;
      33792: inst = 32'd268468224;
      33793: inst = 32'd201343557;
      33794: inst = 32'd203423744;
      33795: inst = 32'd471859200;
      33796: inst = 32'd136314880;
      33797: inst = 32'd268468224;
      33798: inst = 32'd201343558;
      33799: inst = 32'd203423744;
      33800: inst = 32'd471859200;
      33801: inst = 32'd136314880;
      33802: inst = 32'd268468224;
      33803: inst = 32'd201343559;
      33804: inst = 32'd203423744;
      33805: inst = 32'd471859200;
      33806: inst = 32'd136314880;
      33807: inst = 32'd268468224;
      33808: inst = 32'd201343560;
      33809: inst = 32'd203423744;
      33810: inst = 32'd471859200;
      33811: inst = 32'd136314880;
      33812: inst = 32'd268468224;
      33813: inst = 32'd201343561;
      33814: inst = 32'd203423744;
      33815: inst = 32'd471859200;
      33816: inst = 32'd136314880;
      33817: inst = 32'd268468224;
      33818: inst = 32'd201343562;
      33819: inst = 32'd203423744;
      33820: inst = 32'd471859200;
      33821: inst = 32'd136314880;
      33822: inst = 32'd268468224;
      33823: inst = 32'd201343563;
      33824: inst = 32'd203423744;
      33825: inst = 32'd471859200;
      33826: inst = 32'd136314880;
      33827: inst = 32'd268468224;
      33828: inst = 32'd201343564;
      33829: inst = 32'd203423744;
      33830: inst = 32'd471859200;
      33831: inst = 32'd136314880;
      33832: inst = 32'd268468224;
      33833: inst = 32'd201343565;
      33834: inst = 32'd203423744;
      33835: inst = 32'd471859200;
      33836: inst = 32'd136314880;
      33837: inst = 32'd268468224;
      33838: inst = 32'd201343566;
      33839: inst = 32'd203423744;
      33840: inst = 32'd471859200;
      33841: inst = 32'd136314880;
      33842: inst = 32'd268468224;
      33843: inst = 32'd201343567;
      33844: inst = 32'd203423744;
      33845: inst = 32'd471859200;
      33846: inst = 32'd136314880;
      33847: inst = 32'd268468224;
      33848: inst = 32'd201343568;
      33849: inst = 32'd203423744;
      33850: inst = 32'd471859200;
      33851: inst = 32'd136314880;
      33852: inst = 32'd268468224;
      33853: inst = 32'd201343569;
      33854: inst = 32'd203423744;
      33855: inst = 32'd471859200;
      33856: inst = 32'd136314880;
      33857: inst = 32'd268468224;
      33858: inst = 32'd201343570;
      33859: inst = 32'd203423744;
      33860: inst = 32'd471859200;
      33861: inst = 32'd136314880;
      33862: inst = 32'd268468224;
      33863: inst = 32'd201343571;
      33864: inst = 32'd203423744;
      33865: inst = 32'd471859200;
      33866: inst = 32'd136314880;
      33867: inst = 32'd268468224;
      33868: inst = 32'd201343572;
      33869: inst = 32'd203423744;
      33870: inst = 32'd471859200;
      33871: inst = 32'd136314880;
      33872: inst = 32'd268468224;
      33873: inst = 32'd201343573;
      33874: inst = 32'd203423744;
      33875: inst = 32'd471859200;
      33876: inst = 32'd136314880;
      33877: inst = 32'd268468224;
      33878: inst = 32'd201343574;
      33879: inst = 32'd203423744;
      33880: inst = 32'd471859200;
      33881: inst = 32'd136314880;
      33882: inst = 32'd268468224;
      33883: inst = 32'd201343575;
      33884: inst = 32'd203423744;
      33885: inst = 32'd471859200;
      33886: inst = 32'd136314880;
      33887: inst = 32'd268468224;
      33888: inst = 32'd201343576;
      33889: inst = 32'd203423744;
      33890: inst = 32'd471859200;
      33891: inst = 32'd136314880;
      33892: inst = 32'd268468224;
      33893: inst = 32'd201343577;
      33894: inst = 32'd203423744;
      33895: inst = 32'd471859200;
      33896: inst = 32'd136314880;
      33897: inst = 32'd268468224;
      33898: inst = 32'd201343578;
      33899: inst = 32'd203423744;
      33900: inst = 32'd471859200;
      33901: inst = 32'd136314880;
      33902: inst = 32'd268468224;
      33903: inst = 32'd201343579;
      33904: inst = 32'd203423744;
      33905: inst = 32'd471859200;
      33906: inst = 32'd136314880;
      33907: inst = 32'd268468224;
      33908: inst = 32'd201343580;
      33909: inst = 32'd203423744;
      33910: inst = 32'd471859200;
      33911: inst = 32'd136314880;
      33912: inst = 32'd268468224;
      33913: inst = 32'd201343581;
      33914: inst = 32'd203423744;
      33915: inst = 32'd471859200;
      33916: inst = 32'd136314880;
      33917: inst = 32'd268468224;
      33918: inst = 32'd201343582;
      33919: inst = 32'd203423744;
      33920: inst = 32'd471859200;
      33921: inst = 32'd136314880;
      33922: inst = 32'd268468224;
      33923: inst = 32'd201343583;
      33924: inst = 32'd203423744;
      33925: inst = 32'd471859200;
      33926: inst = 32'd136314880;
      33927: inst = 32'd268468224;
      33928: inst = 32'd201343584;
      33929: inst = 32'd203423744;
      33930: inst = 32'd471859200;
      33931: inst = 32'd136314880;
      33932: inst = 32'd268468224;
      33933: inst = 32'd201343585;
      33934: inst = 32'd203423744;
      33935: inst = 32'd471859200;
      33936: inst = 32'd136314880;
      33937: inst = 32'd268468224;
      33938: inst = 32'd201343586;
      33939: inst = 32'd203423744;
      33940: inst = 32'd471859200;
      33941: inst = 32'd136314880;
      33942: inst = 32'd268468224;
      33943: inst = 32'd201343587;
      33944: inst = 32'd203423744;
      33945: inst = 32'd471859200;
      33946: inst = 32'd136314880;
      33947: inst = 32'd268468224;
      33948: inst = 32'd201343588;
      33949: inst = 32'd203423744;
      33950: inst = 32'd471859200;
      33951: inst = 32'd136314880;
      33952: inst = 32'd268468224;
      33953: inst = 32'd201343589;
      33954: inst = 32'd203423744;
      33955: inst = 32'd471859200;
      33956: inst = 32'd136314880;
      33957: inst = 32'd268468224;
      33958: inst = 32'd201343590;
      33959: inst = 32'd203423744;
      33960: inst = 32'd471859200;
      33961: inst = 32'd136314880;
      33962: inst = 32'd268468224;
      33963: inst = 32'd201343591;
      33964: inst = 32'd203423744;
      33965: inst = 32'd471859200;
      33966: inst = 32'd136314880;
      33967: inst = 32'd268468224;
      33968: inst = 32'd201343592;
      33969: inst = 32'd203423744;
      33970: inst = 32'd471859200;
      33971: inst = 32'd136314880;
      33972: inst = 32'd268468224;
      33973: inst = 32'd201343593;
      33974: inst = 32'd203423744;
      33975: inst = 32'd471859200;
      33976: inst = 32'd136314880;
      33977: inst = 32'd268468224;
      33978: inst = 32'd201343594;
      33979: inst = 32'd203423744;
      33980: inst = 32'd471859200;
      33981: inst = 32'd136314880;
      33982: inst = 32'd268468224;
      33983: inst = 32'd201343595;
      33984: inst = 32'd203423744;
      33985: inst = 32'd471859200;
      33986: inst = 32'd136314880;
      33987: inst = 32'd268468224;
      33988: inst = 32'd201343596;
      33989: inst = 32'd203423744;
      33990: inst = 32'd471859200;
      33991: inst = 32'd136314880;
      33992: inst = 32'd268468224;
      33993: inst = 32'd201343597;
      33994: inst = 32'd203423744;
      33995: inst = 32'd471859200;
      33996: inst = 32'd136314880;
      33997: inst = 32'd268468224;
      33998: inst = 32'd201343598;
      33999: inst = 32'd203423744;
      34000: inst = 32'd471859200;
      34001: inst = 32'd136314880;
      34002: inst = 32'd268468224;
      34003: inst = 32'd201343599;
      34004: inst = 32'd203423744;
      34005: inst = 32'd471859200;
      34006: inst = 32'd136314880;
      34007: inst = 32'd268468224;
      34008: inst = 32'd201343600;
      34009: inst = 32'd203423744;
      34010: inst = 32'd471859200;
      34011: inst = 32'd136314880;
      34012: inst = 32'd268468224;
      34013: inst = 32'd201343601;
      34014: inst = 32'd203423744;
      34015: inst = 32'd471859200;
      34016: inst = 32'd136314880;
      34017: inst = 32'd268468224;
      34018: inst = 32'd201343602;
      34019: inst = 32'd203423744;
      34020: inst = 32'd471859200;
      34021: inst = 32'd136314880;
      34022: inst = 32'd268468224;
      34023: inst = 32'd201343603;
      34024: inst = 32'd203423744;
      34025: inst = 32'd471859200;
      34026: inst = 32'd136314880;
      34027: inst = 32'd268468224;
      34028: inst = 32'd201343604;
      34029: inst = 32'd203423744;
      34030: inst = 32'd471859200;
      34031: inst = 32'd136314880;
      34032: inst = 32'd268468224;
      34033: inst = 32'd201343605;
      34034: inst = 32'd203423744;
      34035: inst = 32'd471859200;
      34036: inst = 32'd136314880;
      34037: inst = 32'd268468224;
      34038: inst = 32'd201343606;
      34039: inst = 32'd203423744;
      34040: inst = 32'd471859200;
      34041: inst = 32'd136314880;
      34042: inst = 32'd268468224;
      34043: inst = 32'd201343607;
      34044: inst = 32'd203423744;
      34045: inst = 32'd471859200;
      34046: inst = 32'd136314880;
      34047: inst = 32'd268468224;
      34048: inst = 32'd201343608;
      34049: inst = 32'd203423744;
      34050: inst = 32'd471859200;
      34051: inst = 32'd136314880;
      34052: inst = 32'd268468224;
      34053: inst = 32'd201343609;
      34054: inst = 32'd203423744;
      34055: inst = 32'd471859200;
      34056: inst = 32'd136314880;
      34057: inst = 32'd268468224;
      34058: inst = 32'd201343610;
      34059: inst = 32'd203423744;
      34060: inst = 32'd471859200;
      34061: inst = 32'd136314880;
      34062: inst = 32'd268468224;
      34063: inst = 32'd201343611;
      34064: inst = 32'd203423744;
      34065: inst = 32'd471859200;
      34066: inst = 32'd136314880;
      34067: inst = 32'd268468224;
      34068: inst = 32'd201343612;
      34069: inst = 32'd203423744;
      34070: inst = 32'd471859200;
      34071: inst = 32'd136314880;
      34072: inst = 32'd268468224;
      34073: inst = 32'd201343613;
      34074: inst = 32'd203423744;
      34075: inst = 32'd471859200;
      34076: inst = 32'd136314880;
      34077: inst = 32'd268468224;
      34078: inst = 32'd201343614;
      34079: inst = 32'd203423744;
      34080: inst = 32'd471859200;
      34081: inst = 32'd136314880;
      34082: inst = 32'd268468224;
      34083: inst = 32'd201343615;
      34084: inst = 32'd203423744;
      34085: inst = 32'd471859200;
      34086: inst = 32'd136314880;
      34087: inst = 32'd268468224;
      34088: inst = 32'd201343616;
      34089: inst = 32'd203423744;
      34090: inst = 32'd471859200;
      34091: inst = 32'd136314880;
      34092: inst = 32'd268468224;
      34093: inst = 32'd201343617;
      34094: inst = 32'd203423744;
      34095: inst = 32'd471859200;
      34096: inst = 32'd136314880;
      34097: inst = 32'd268468224;
      34098: inst = 32'd201343618;
      34099: inst = 32'd203423744;
      34100: inst = 32'd471859200;
      34101: inst = 32'd136314880;
      34102: inst = 32'd268468224;
      34103: inst = 32'd201343619;
      34104: inst = 32'd203423744;
      34105: inst = 32'd471859200;
      34106: inst = 32'd136314880;
      34107: inst = 32'd268468224;
      34108: inst = 32'd201343620;
      34109: inst = 32'd203423744;
      34110: inst = 32'd471859200;
      34111: inst = 32'd136314880;
      34112: inst = 32'd268468224;
      34113: inst = 32'd201343621;
      34114: inst = 32'd203423744;
      34115: inst = 32'd471859200;
      34116: inst = 32'd136314880;
      34117: inst = 32'd268468224;
      34118: inst = 32'd201343622;
      34119: inst = 32'd203423744;
      34120: inst = 32'd471859200;
      34121: inst = 32'd136314880;
      34122: inst = 32'd268468224;
      34123: inst = 32'd201343623;
      34124: inst = 32'd203423744;
      34125: inst = 32'd471859200;
      34126: inst = 32'd136314880;
      34127: inst = 32'd268468224;
      34128: inst = 32'd201343624;
      34129: inst = 32'd203423744;
      34130: inst = 32'd471859200;
      34131: inst = 32'd136314880;
      34132: inst = 32'd268468224;
      34133: inst = 32'd201343625;
      34134: inst = 32'd203423744;
      34135: inst = 32'd471859200;
      34136: inst = 32'd136314880;
      34137: inst = 32'd268468224;
      34138: inst = 32'd201343626;
      34139: inst = 32'd203423744;
      34140: inst = 32'd471859200;
      34141: inst = 32'd136314880;
      34142: inst = 32'd268468224;
      34143: inst = 32'd201343627;
      34144: inst = 32'd203423744;
      34145: inst = 32'd471859200;
      34146: inst = 32'd136314880;
      34147: inst = 32'd268468224;
      34148: inst = 32'd201343628;
      34149: inst = 32'd203423744;
      34150: inst = 32'd471859200;
      34151: inst = 32'd136314880;
      34152: inst = 32'd268468224;
      34153: inst = 32'd201343629;
      34154: inst = 32'd203423744;
      34155: inst = 32'd471859200;
      34156: inst = 32'd136314880;
      34157: inst = 32'd268468224;
      34158: inst = 32'd201343630;
      34159: inst = 32'd203423744;
      34160: inst = 32'd471859200;
      34161: inst = 32'd136314880;
      34162: inst = 32'd268468224;
      34163: inst = 32'd201343631;
      34164: inst = 32'd203423744;
      34165: inst = 32'd471859200;
      34166: inst = 32'd136314880;
      34167: inst = 32'd268468224;
      34168: inst = 32'd201343632;
      34169: inst = 32'd203423744;
      34170: inst = 32'd471859200;
      34171: inst = 32'd136314880;
      34172: inst = 32'd268468224;
      34173: inst = 32'd201343633;
      34174: inst = 32'd203423744;
      34175: inst = 32'd471859200;
      34176: inst = 32'd136314880;
      34177: inst = 32'd268468224;
      34178: inst = 32'd201343634;
      34179: inst = 32'd203423744;
      34180: inst = 32'd471859200;
      34181: inst = 32'd136314880;
      34182: inst = 32'd268468224;
      34183: inst = 32'd201343635;
      34184: inst = 32'd203423744;
      34185: inst = 32'd471859200;
      34186: inst = 32'd136314880;
      34187: inst = 32'd268468224;
      34188: inst = 32'd201343636;
      34189: inst = 32'd203423744;
      34190: inst = 32'd471859200;
      34191: inst = 32'd136314880;
      34192: inst = 32'd268468224;
      34193: inst = 32'd201343637;
      34194: inst = 32'd203423744;
      34195: inst = 32'd471859200;
      34196: inst = 32'd136314880;
      34197: inst = 32'd268468224;
      34198: inst = 32'd201343638;
      34199: inst = 32'd203423744;
      34200: inst = 32'd471859200;
      34201: inst = 32'd136314880;
      34202: inst = 32'd268468224;
      34203: inst = 32'd201343639;
      34204: inst = 32'd203423744;
      34205: inst = 32'd471859200;
      34206: inst = 32'd136314880;
      34207: inst = 32'd268468224;
      34208: inst = 32'd201343640;
      34209: inst = 32'd203423744;
      34210: inst = 32'd471859200;
      34211: inst = 32'd136314880;
      34212: inst = 32'd268468224;
      34213: inst = 32'd201343641;
      34214: inst = 32'd203423744;
      34215: inst = 32'd471859200;
      34216: inst = 32'd136314880;
      34217: inst = 32'd268468224;
      34218: inst = 32'd201343642;
      34219: inst = 32'd203423744;
      34220: inst = 32'd471859200;
      34221: inst = 32'd136314880;
      34222: inst = 32'd268468224;
      34223: inst = 32'd201343643;
      34224: inst = 32'd203423744;
      34225: inst = 32'd471859200;
      34226: inst = 32'd136314880;
      34227: inst = 32'd268468224;
      34228: inst = 32'd201343644;
      34229: inst = 32'd203423744;
      34230: inst = 32'd471859200;
      34231: inst = 32'd136314880;
      34232: inst = 32'd268468224;
      34233: inst = 32'd201343645;
      34234: inst = 32'd203423744;
      34235: inst = 32'd471859200;
      34236: inst = 32'd136314880;
      34237: inst = 32'd268468224;
      34238: inst = 32'd201343646;
      34239: inst = 32'd203423744;
      34240: inst = 32'd471859200;
      34241: inst = 32'd136314880;
      34242: inst = 32'd268468224;
      34243: inst = 32'd201343647;
      34244: inst = 32'd203423744;
      34245: inst = 32'd471859200;
      34246: inst = 32'd136314880;
      34247: inst = 32'd268468224;
      34248: inst = 32'd201343648;
      34249: inst = 32'd203423744;
      34250: inst = 32'd471859200;
      34251: inst = 32'd136314880;
      34252: inst = 32'd268468224;
      34253: inst = 32'd201343649;
      34254: inst = 32'd203423744;
      34255: inst = 32'd471859200;
      34256: inst = 32'd136314880;
      34257: inst = 32'd268468224;
      34258: inst = 32'd201343650;
      34259: inst = 32'd203423744;
      34260: inst = 32'd471859200;
      34261: inst = 32'd136314880;
      34262: inst = 32'd268468224;
      34263: inst = 32'd201343651;
      34264: inst = 32'd203423744;
      34265: inst = 32'd471859200;
      34266: inst = 32'd136314880;
      34267: inst = 32'd268468224;
      34268: inst = 32'd201343652;
      34269: inst = 32'd203423744;
      34270: inst = 32'd471859200;
      34271: inst = 32'd136314880;
      34272: inst = 32'd268468224;
      34273: inst = 32'd201343653;
      34274: inst = 32'd203423744;
      34275: inst = 32'd471859200;
      34276: inst = 32'd136314880;
      34277: inst = 32'd268468224;
      34278: inst = 32'd201343654;
      34279: inst = 32'd203423744;
      34280: inst = 32'd471859200;
      34281: inst = 32'd136314880;
      34282: inst = 32'd268468224;
      34283: inst = 32'd201343655;
      34284: inst = 32'd203423744;
      34285: inst = 32'd471859200;
      34286: inst = 32'd136314880;
      34287: inst = 32'd268468224;
      34288: inst = 32'd201343656;
      34289: inst = 32'd203423744;
      34290: inst = 32'd471859200;
      34291: inst = 32'd136314880;
      34292: inst = 32'd268468224;
      34293: inst = 32'd201343657;
      34294: inst = 32'd203423744;
      34295: inst = 32'd471859200;
      34296: inst = 32'd136314880;
      34297: inst = 32'd268468224;
      34298: inst = 32'd201343658;
      34299: inst = 32'd203423744;
      34300: inst = 32'd471859200;
      34301: inst = 32'd136314880;
      34302: inst = 32'd268468224;
      34303: inst = 32'd201343659;
      34304: inst = 32'd203423744;
      34305: inst = 32'd471859200;
      34306: inst = 32'd136314880;
      34307: inst = 32'd268468224;
      34308: inst = 32'd201343660;
      34309: inst = 32'd203423744;
      34310: inst = 32'd471859200;
      34311: inst = 32'd136314880;
      34312: inst = 32'd268468224;
      34313: inst = 32'd201343661;
      34314: inst = 32'd203423744;
      34315: inst = 32'd471859200;
      34316: inst = 32'd136314880;
      34317: inst = 32'd268468224;
      34318: inst = 32'd201343662;
      34319: inst = 32'd203423744;
      34320: inst = 32'd471859200;
      34321: inst = 32'd136314880;
      34322: inst = 32'd268468224;
      34323: inst = 32'd201343663;
      34324: inst = 32'd203423744;
      34325: inst = 32'd471859200;
      34326: inst = 32'd136314880;
      34327: inst = 32'd268468224;
      34328: inst = 32'd201343664;
      34329: inst = 32'd203423744;
      34330: inst = 32'd471859200;
      34331: inst = 32'd136314880;
      34332: inst = 32'd268468224;
      34333: inst = 32'd201343665;
      34334: inst = 32'd203423744;
      34335: inst = 32'd471859200;
      34336: inst = 32'd136314880;
      34337: inst = 32'd268468224;
      34338: inst = 32'd201343666;
      34339: inst = 32'd203423744;
      34340: inst = 32'd471859200;
      34341: inst = 32'd136314880;
      34342: inst = 32'd268468224;
      34343: inst = 32'd201343667;
      34344: inst = 32'd203423744;
      34345: inst = 32'd471859200;
      34346: inst = 32'd136314880;
      34347: inst = 32'd268468224;
      34348: inst = 32'd201343668;
      34349: inst = 32'd203423744;
      34350: inst = 32'd471859200;
      34351: inst = 32'd136314880;
      34352: inst = 32'd268468224;
      34353: inst = 32'd201343669;
      34354: inst = 32'd203423744;
      34355: inst = 32'd471859200;
      34356: inst = 32'd136314880;
      34357: inst = 32'd268468224;
      34358: inst = 32'd201343670;
      34359: inst = 32'd203423744;
      34360: inst = 32'd471859200;
      34361: inst = 32'd136314880;
      34362: inst = 32'd268468224;
      34363: inst = 32'd201343671;
      34364: inst = 32'd203423744;
      34365: inst = 32'd471859200;
      34366: inst = 32'd136314880;
      34367: inst = 32'd268468224;
      34368: inst = 32'd201343672;
      34369: inst = 32'd203423744;
      34370: inst = 32'd471859200;
      34371: inst = 32'd136314880;
      34372: inst = 32'd268468224;
      34373: inst = 32'd201343673;
      34374: inst = 32'd203423744;
      34375: inst = 32'd471859200;
      34376: inst = 32'd136314880;
      34377: inst = 32'd268468224;
      34378: inst = 32'd201343674;
      34379: inst = 32'd203423744;
      34380: inst = 32'd471859200;
      34381: inst = 32'd136314880;
      34382: inst = 32'd268468224;
      34383: inst = 32'd201343675;
      34384: inst = 32'd203423744;
      34385: inst = 32'd471859200;
      34386: inst = 32'd136314880;
      34387: inst = 32'd268468224;
      34388: inst = 32'd201343676;
      34389: inst = 32'd203423744;
      34390: inst = 32'd471859200;
      34391: inst = 32'd136314880;
      34392: inst = 32'd268468224;
      34393: inst = 32'd201343677;
      34394: inst = 32'd203423744;
      34395: inst = 32'd471859200;
      34396: inst = 32'd136314880;
      34397: inst = 32'd268468224;
      34398: inst = 32'd201343678;
      34399: inst = 32'd203423744;
      34400: inst = 32'd471859200;
      34401: inst = 32'd136314880;
      34402: inst = 32'd268468224;
      34403: inst = 32'd201343679;
      34404: inst = 32'd203423744;
      34405: inst = 32'd471859200;
      34406: inst = 32'd136314880;
      34407: inst = 32'd268468224;
      34408: inst = 32'd201343680;
      34409: inst = 32'd203423744;
      34410: inst = 32'd471859200;
      34411: inst = 32'd136314880;
      34412: inst = 32'd268468224;
      34413: inst = 32'd201343681;
      34414: inst = 32'd203423744;
      34415: inst = 32'd471859200;
      34416: inst = 32'd136314880;
      34417: inst = 32'd268468224;
      34418: inst = 32'd201343682;
      34419: inst = 32'd203423744;
      34420: inst = 32'd471859200;
      34421: inst = 32'd136314880;
      34422: inst = 32'd268468224;
      34423: inst = 32'd201343683;
      34424: inst = 32'd203423744;
      34425: inst = 32'd471859200;
      34426: inst = 32'd136314880;
      34427: inst = 32'd268468224;
      34428: inst = 32'd201343684;
      34429: inst = 32'd203423744;
      34430: inst = 32'd471859200;
      34431: inst = 32'd136314880;
      34432: inst = 32'd268468224;
      34433: inst = 32'd201343685;
      34434: inst = 32'd203423744;
      34435: inst = 32'd471859200;
      34436: inst = 32'd136314880;
      34437: inst = 32'd268468224;
      34438: inst = 32'd201343686;
      34439: inst = 32'd203423744;
      34440: inst = 32'd471859200;
      34441: inst = 32'd136314880;
      34442: inst = 32'd268468224;
      34443: inst = 32'd201343687;
      34444: inst = 32'd203423744;
      34445: inst = 32'd471859200;
      34446: inst = 32'd136314880;
      34447: inst = 32'd268468224;
      34448: inst = 32'd201343688;
      34449: inst = 32'd203423744;
      34450: inst = 32'd471859200;
      34451: inst = 32'd136314880;
      34452: inst = 32'd268468224;
      34453: inst = 32'd201343689;
      34454: inst = 32'd203423744;
      34455: inst = 32'd471859200;
      34456: inst = 32'd136314880;
      34457: inst = 32'd268468224;
      34458: inst = 32'd201343690;
      34459: inst = 32'd203423744;
      34460: inst = 32'd471859200;
      34461: inst = 32'd136314880;
      34462: inst = 32'd268468224;
      34463: inst = 32'd201343691;
      34464: inst = 32'd203423744;
      34465: inst = 32'd471859200;
      34466: inst = 32'd136314880;
      34467: inst = 32'd268468224;
      34468: inst = 32'd201343692;
      34469: inst = 32'd203423744;
      34470: inst = 32'd471859200;
      34471: inst = 32'd136314880;
      34472: inst = 32'd268468224;
      34473: inst = 32'd201343693;
      34474: inst = 32'd203423744;
      34475: inst = 32'd471859200;
      34476: inst = 32'd136314880;
      34477: inst = 32'd268468224;
      34478: inst = 32'd201343694;
      34479: inst = 32'd203423744;
      34480: inst = 32'd471859200;
      34481: inst = 32'd136314880;
      34482: inst = 32'd268468224;
      34483: inst = 32'd201343695;
      34484: inst = 32'd203423744;
      34485: inst = 32'd471859200;
      34486: inst = 32'd136314880;
      34487: inst = 32'd268468224;
      34488: inst = 32'd201343696;
      34489: inst = 32'd203423744;
      34490: inst = 32'd471859200;
      34491: inst = 32'd136314880;
      34492: inst = 32'd268468224;
      34493: inst = 32'd201343697;
      34494: inst = 32'd203423744;
      34495: inst = 32'd471859200;
      34496: inst = 32'd136314880;
      34497: inst = 32'd268468224;
      34498: inst = 32'd201343698;
      34499: inst = 32'd203423744;
      34500: inst = 32'd471859200;
      34501: inst = 32'd136314880;
      34502: inst = 32'd268468224;
      34503: inst = 32'd201343699;
      34504: inst = 32'd203423744;
      34505: inst = 32'd471859200;
      34506: inst = 32'd136314880;
      34507: inst = 32'd268468224;
      34508: inst = 32'd201343700;
      34509: inst = 32'd203423744;
      34510: inst = 32'd471859200;
      34511: inst = 32'd136314880;
      34512: inst = 32'd268468224;
      34513: inst = 32'd201343701;
      34514: inst = 32'd203423744;
      34515: inst = 32'd471859200;
      34516: inst = 32'd136314880;
      34517: inst = 32'd268468224;
      34518: inst = 32'd201343702;
      34519: inst = 32'd203423744;
      34520: inst = 32'd471859200;
      34521: inst = 32'd136314880;
      34522: inst = 32'd268468224;
      34523: inst = 32'd201343703;
      34524: inst = 32'd203423744;
      34525: inst = 32'd471859200;
      34526: inst = 32'd136314880;
      34527: inst = 32'd268468224;
      34528: inst = 32'd201343704;
      34529: inst = 32'd203423744;
      34530: inst = 32'd471859200;
      34531: inst = 32'd136314880;
      34532: inst = 32'd268468224;
      34533: inst = 32'd201343705;
      34534: inst = 32'd203423744;
      34535: inst = 32'd471859200;
      34536: inst = 32'd136314880;
      34537: inst = 32'd268468224;
      34538: inst = 32'd201343706;
      34539: inst = 32'd203423744;
      34540: inst = 32'd471859200;
      34541: inst = 32'd136314880;
      34542: inst = 32'd268468224;
      34543: inst = 32'd201343707;
      34544: inst = 32'd203423744;
      34545: inst = 32'd471859200;
      34546: inst = 32'd136314880;
      34547: inst = 32'd268468224;
      34548: inst = 32'd201343708;
      34549: inst = 32'd203423744;
      34550: inst = 32'd471859200;
      34551: inst = 32'd136314880;
      34552: inst = 32'd268468224;
      34553: inst = 32'd201343709;
      34554: inst = 32'd203423744;
      34555: inst = 32'd471859200;
      34556: inst = 32'd136314880;
      34557: inst = 32'd268468224;
      34558: inst = 32'd201343710;
      34559: inst = 32'd203423744;
      34560: inst = 32'd471859200;
      34561: inst = 32'd136314880;
      34562: inst = 32'd268468224;
      34563: inst = 32'd201343711;
      34564: inst = 32'd203423744;
      34565: inst = 32'd471859200;
      34566: inst = 32'd136314880;
      34567: inst = 32'd268468224;
      34568: inst = 32'd201343712;
      34569: inst = 32'd203423744;
      34570: inst = 32'd471859200;
      34571: inst = 32'd136314880;
      34572: inst = 32'd268468224;
      34573: inst = 32'd201343713;
      34574: inst = 32'd203423744;
      34575: inst = 32'd471859200;
      34576: inst = 32'd136314880;
      34577: inst = 32'd268468224;
      34578: inst = 32'd201343714;
      34579: inst = 32'd203423744;
      34580: inst = 32'd471859200;
      34581: inst = 32'd136314880;
      34582: inst = 32'd268468224;
      34583: inst = 32'd201343715;
      34584: inst = 32'd203423744;
      34585: inst = 32'd471859200;
      34586: inst = 32'd136314880;
      34587: inst = 32'd268468224;
      34588: inst = 32'd201343716;
      34589: inst = 32'd203423744;
      34590: inst = 32'd471859200;
      34591: inst = 32'd136314880;
      34592: inst = 32'd268468224;
      34593: inst = 32'd201343717;
      34594: inst = 32'd203423744;
      34595: inst = 32'd471859200;
      34596: inst = 32'd136314880;
      34597: inst = 32'd268468224;
      34598: inst = 32'd201343718;
      34599: inst = 32'd203423744;
      34600: inst = 32'd471859200;
      34601: inst = 32'd136314880;
      34602: inst = 32'd268468224;
      34603: inst = 32'd201343719;
      34604: inst = 32'd203423744;
      34605: inst = 32'd471859200;
      34606: inst = 32'd136314880;
      34607: inst = 32'd268468224;
      34608: inst = 32'd201343720;
      34609: inst = 32'd203423744;
      34610: inst = 32'd471859200;
      34611: inst = 32'd136314880;
      34612: inst = 32'd268468224;
      34613: inst = 32'd201343721;
      34614: inst = 32'd203423744;
      34615: inst = 32'd471859200;
      34616: inst = 32'd136314880;
      34617: inst = 32'd268468224;
      34618: inst = 32'd201343722;
      34619: inst = 32'd203423744;
      34620: inst = 32'd471859200;
      34621: inst = 32'd136314880;
      34622: inst = 32'd268468224;
      34623: inst = 32'd201343723;
      34624: inst = 32'd203423744;
      34625: inst = 32'd471859200;
      34626: inst = 32'd136314880;
      34627: inst = 32'd268468224;
      34628: inst = 32'd201343724;
      34629: inst = 32'd203423744;
      34630: inst = 32'd471859200;
      34631: inst = 32'd136314880;
      34632: inst = 32'd268468224;
      34633: inst = 32'd201343725;
      34634: inst = 32'd203423744;
      34635: inst = 32'd471859200;
      34636: inst = 32'd136314880;
      34637: inst = 32'd268468224;
      34638: inst = 32'd201343726;
      34639: inst = 32'd203423744;
      34640: inst = 32'd471859200;
      34641: inst = 32'd136314880;
      34642: inst = 32'd268468224;
      34643: inst = 32'd201343727;
      34644: inst = 32'd203423744;
      34645: inst = 32'd471859200;
      34646: inst = 32'd136314880;
      34647: inst = 32'd268468224;
      34648: inst = 32'd201343728;
      34649: inst = 32'd203423744;
      34650: inst = 32'd471859200;
      34651: inst = 32'd136314880;
      34652: inst = 32'd268468224;
      34653: inst = 32'd201343729;
      34654: inst = 32'd203423744;
      34655: inst = 32'd471859200;
      34656: inst = 32'd136314880;
      34657: inst = 32'd268468224;
      34658: inst = 32'd201343730;
      34659: inst = 32'd203423744;
      34660: inst = 32'd471859200;
      34661: inst = 32'd136314880;
      34662: inst = 32'd268468224;
      34663: inst = 32'd201343731;
      34664: inst = 32'd203423744;
      34665: inst = 32'd471859200;
      34666: inst = 32'd136314880;
      34667: inst = 32'd268468224;
      34668: inst = 32'd201343732;
      34669: inst = 32'd203423744;
      34670: inst = 32'd471859200;
      34671: inst = 32'd136314880;
      34672: inst = 32'd268468224;
      34673: inst = 32'd201343733;
      34674: inst = 32'd203423744;
      34675: inst = 32'd471859200;
      34676: inst = 32'd136314880;
      34677: inst = 32'd268468224;
      34678: inst = 32'd201343734;
      34679: inst = 32'd203423744;
      34680: inst = 32'd471859200;
      34681: inst = 32'd136314880;
      34682: inst = 32'd268468224;
      34683: inst = 32'd201343735;
      34684: inst = 32'd203423744;
      34685: inst = 32'd471859200;
      34686: inst = 32'd136314880;
      34687: inst = 32'd268468224;
      34688: inst = 32'd201343736;
      34689: inst = 32'd203423744;
      34690: inst = 32'd471859200;
      34691: inst = 32'd136314880;
      34692: inst = 32'd268468224;
      34693: inst = 32'd201343737;
      34694: inst = 32'd203423744;
      34695: inst = 32'd471859200;
      34696: inst = 32'd136314880;
      34697: inst = 32'd268468224;
      34698: inst = 32'd201343738;
      34699: inst = 32'd203423744;
      34700: inst = 32'd471859200;
      34701: inst = 32'd136314880;
      34702: inst = 32'd268468224;
      34703: inst = 32'd201343739;
      34704: inst = 32'd203423744;
      34705: inst = 32'd471859200;
      34706: inst = 32'd136314880;
      34707: inst = 32'd268468224;
      34708: inst = 32'd201343740;
      34709: inst = 32'd203423744;
      34710: inst = 32'd471859200;
      34711: inst = 32'd136314880;
      34712: inst = 32'd268468224;
      34713: inst = 32'd201343741;
      34714: inst = 32'd203423744;
      34715: inst = 32'd471859200;
      34716: inst = 32'd136314880;
      34717: inst = 32'd268468224;
      34718: inst = 32'd201343742;
      34719: inst = 32'd203423744;
      34720: inst = 32'd471859200;
      34721: inst = 32'd136314880;
      34722: inst = 32'd268468224;
      34723: inst = 32'd201343743;
      34724: inst = 32'd203423744;
      34725: inst = 32'd471859200;
      34726: inst = 32'd136314880;
      34727: inst = 32'd268468224;
      34728: inst = 32'd201343744;
      34729: inst = 32'd203423744;
      34730: inst = 32'd471859200;
      34731: inst = 32'd136314880;
      34732: inst = 32'd268468224;
      34733: inst = 32'd201343745;
      34734: inst = 32'd203423744;
      34735: inst = 32'd471859200;
      34736: inst = 32'd136314880;
      34737: inst = 32'd268468224;
      34738: inst = 32'd201343746;
      34739: inst = 32'd203423744;
      34740: inst = 32'd471859200;
      34741: inst = 32'd136314880;
      34742: inst = 32'd268468224;
      34743: inst = 32'd201343747;
      34744: inst = 32'd203423744;
      34745: inst = 32'd471859200;
      34746: inst = 32'd136314880;
      34747: inst = 32'd268468224;
      34748: inst = 32'd201343748;
      34749: inst = 32'd203423744;
      34750: inst = 32'd471859200;
      34751: inst = 32'd136314880;
      34752: inst = 32'd268468224;
      34753: inst = 32'd201343749;
      34754: inst = 32'd203423744;
      34755: inst = 32'd471859200;
      34756: inst = 32'd136314880;
      34757: inst = 32'd268468224;
      34758: inst = 32'd201343750;
      34759: inst = 32'd203423744;
      34760: inst = 32'd471859200;
      34761: inst = 32'd136314880;
      34762: inst = 32'd268468224;
      34763: inst = 32'd201343751;
      34764: inst = 32'd203423744;
      34765: inst = 32'd471859200;
      34766: inst = 32'd136314880;
      34767: inst = 32'd268468224;
      34768: inst = 32'd201343752;
      34769: inst = 32'd203423744;
      34770: inst = 32'd471859200;
      34771: inst = 32'd136314880;
      34772: inst = 32'd268468224;
      34773: inst = 32'd201343753;
      34774: inst = 32'd203423744;
      34775: inst = 32'd471859200;
      34776: inst = 32'd136314880;
      34777: inst = 32'd268468224;
      34778: inst = 32'd201343754;
      34779: inst = 32'd203423744;
      34780: inst = 32'd471859200;
      34781: inst = 32'd136314880;
      34782: inst = 32'd268468224;
      34783: inst = 32'd201343755;
      34784: inst = 32'd203423744;
      34785: inst = 32'd471859200;
      34786: inst = 32'd136314880;
      34787: inst = 32'd268468224;
      34788: inst = 32'd201343756;
      34789: inst = 32'd203423744;
      34790: inst = 32'd471859200;
      34791: inst = 32'd136314880;
      34792: inst = 32'd268468224;
      34793: inst = 32'd201343757;
      34794: inst = 32'd203423744;
      34795: inst = 32'd471859200;
      34796: inst = 32'd136314880;
      34797: inst = 32'd268468224;
      34798: inst = 32'd201343758;
      34799: inst = 32'd203423744;
      34800: inst = 32'd471859200;
      34801: inst = 32'd136314880;
      34802: inst = 32'd268468224;
      34803: inst = 32'd201343759;
      34804: inst = 32'd203423744;
      34805: inst = 32'd471859200;
      34806: inst = 32'd136314880;
      34807: inst = 32'd268468224;
      34808: inst = 32'd201343760;
      34809: inst = 32'd203423744;
      34810: inst = 32'd471859200;
      34811: inst = 32'd136314880;
      34812: inst = 32'd268468224;
      34813: inst = 32'd201343761;
      34814: inst = 32'd203423744;
      34815: inst = 32'd471859200;
      34816: inst = 32'd136314880;
      34817: inst = 32'd268468224;
      34818: inst = 32'd201343762;
      34819: inst = 32'd203423744;
      34820: inst = 32'd471859200;
      34821: inst = 32'd136314880;
      34822: inst = 32'd268468224;
      34823: inst = 32'd201343763;
      34824: inst = 32'd203423744;
      34825: inst = 32'd471859200;
      34826: inst = 32'd136314880;
      34827: inst = 32'd268468224;
      34828: inst = 32'd201343764;
      34829: inst = 32'd203423744;
      34830: inst = 32'd471859200;
      34831: inst = 32'd136314880;
      34832: inst = 32'd268468224;
      34833: inst = 32'd201343765;
      34834: inst = 32'd203423744;
      34835: inst = 32'd471859200;
      34836: inst = 32'd136314880;
      34837: inst = 32'd268468224;
      34838: inst = 32'd201343766;
      34839: inst = 32'd203423744;
      34840: inst = 32'd471859200;
      34841: inst = 32'd136314880;
      34842: inst = 32'd268468224;
      34843: inst = 32'd201343767;
      34844: inst = 32'd203423744;
      34845: inst = 32'd471859200;
      34846: inst = 32'd136314880;
      34847: inst = 32'd268468224;
      34848: inst = 32'd201343768;
      34849: inst = 32'd203423744;
      34850: inst = 32'd471859200;
      34851: inst = 32'd136314880;
      34852: inst = 32'd268468224;
      34853: inst = 32'd201343769;
      34854: inst = 32'd203423744;
      34855: inst = 32'd471859200;
      34856: inst = 32'd136314880;
      34857: inst = 32'd268468224;
      34858: inst = 32'd201343770;
      34859: inst = 32'd203423744;
      34860: inst = 32'd471859200;
      34861: inst = 32'd136314880;
      34862: inst = 32'd268468224;
      34863: inst = 32'd201343771;
      34864: inst = 32'd203423744;
      34865: inst = 32'd471859200;
      34866: inst = 32'd136314880;
      34867: inst = 32'd268468224;
      34868: inst = 32'd201343772;
      34869: inst = 32'd203423744;
      34870: inst = 32'd471859200;
      34871: inst = 32'd136314880;
      34872: inst = 32'd268468224;
      34873: inst = 32'd201343773;
      34874: inst = 32'd203423744;
      34875: inst = 32'd471859200;
      34876: inst = 32'd136314880;
      34877: inst = 32'd268468224;
      34878: inst = 32'd201343774;
      34879: inst = 32'd203423744;
      34880: inst = 32'd471859200;
      34881: inst = 32'd136314880;
      34882: inst = 32'd268468224;
      34883: inst = 32'd201343775;
      34884: inst = 32'd203423744;
      34885: inst = 32'd471859200;
      34886: inst = 32'd136314880;
      34887: inst = 32'd268468224;
      34888: inst = 32'd201343776;
      34889: inst = 32'd203423744;
      34890: inst = 32'd471859200;
      34891: inst = 32'd136314880;
      34892: inst = 32'd268468224;
      34893: inst = 32'd201343777;
      34894: inst = 32'd203423744;
      34895: inst = 32'd471859200;
      34896: inst = 32'd136314880;
      34897: inst = 32'd268468224;
      34898: inst = 32'd201343778;
      34899: inst = 32'd203423744;
      34900: inst = 32'd471859200;
      34901: inst = 32'd136314880;
      34902: inst = 32'd268468224;
      34903: inst = 32'd201343779;
      34904: inst = 32'd203423744;
      34905: inst = 32'd471859200;
      34906: inst = 32'd136314880;
      34907: inst = 32'd268468224;
      34908: inst = 32'd201343780;
      34909: inst = 32'd203423744;
      34910: inst = 32'd471859200;
      34911: inst = 32'd136314880;
      34912: inst = 32'd268468224;
      34913: inst = 32'd201343781;
      34914: inst = 32'd203423744;
      34915: inst = 32'd471859200;
      34916: inst = 32'd136314880;
      34917: inst = 32'd268468224;
      34918: inst = 32'd201343782;
      34919: inst = 32'd203423744;
      34920: inst = 32'd471859200;
      34921: inst = 32'd136314880;
      34922: inst = 32'd268468224;
      34923: inst = 32'd201343783;
      34924: inst = 32'd203423744;
      34925: inst = 32'd471859200;
      34926: inst = 32'd136314880;
      34927: inst = 32'd268468224;
      34928: inst = 32'd201343784;
      34929: inst = 32'd203423744;
      34930: inst = 32'd471859200;
      34931: inst = 32'd136314880;
      34932: inst = 32'd268468224;
      34933: inst = 32'd201343785;
      34934: inst = 32'd203423744;
      34935: inst = 32'd471859200;
      34936: inst = 32'd136314880;
      34937: inst = 32'd268468224;
      34938: inst = 32'd201343786;
      34939: inst = 32'd203423744;
      34940: inst = 32'd471859200;
      34941: inst = 32'd136314880;
      34942: inst = 32'd268468224;
      34943: inst = 32'd201343787;
      34944: inst = 32'd203423744;
      34945: inst = 32'd471859200;
      34946: inst = 32'd136314880;
      34947: inst = 32'd268468224;
      34948: inst = 32'd201343788;
      34949: inst = 32'd203423744;
      34950: inst = 32'd471859200;
      34951: inst = 32'd136314880;
      34952: inst = 32'd268468224;
      34953: inst = 32'd201343789;
      34954: inst = 32'd203423744;
      34955: inst = 32'd471859200;
      34956: inst = 32'd136314880;
      34957: inst = 32'd268468224;
      34958: inst = 32'd201343790;
      34959: inst = 32'd203423744;
      34960: inst = 32'd471859200;
      34961: inst = 32'd136314880;
      34962: inst = 32'd268468224;
      34963: inst = 32'd201343791;
      34964: inst = 32'd203423744;
      34965: inst = 32'd471859200;
      34966: inst = 32'd136314880;
      34967: inst = 32'd268468224;
      34968: inst = 32'd201343792;
      34969: inst = 32'd203423744;
      34970: inst = 32'd471859200;
      34971: inst = 32'd136314880;
      34972: inst = 32'd268468224;
      34973: inst = 32'd201343793;
      34974: inst = 32'd203423744;
      34975: inst = 32'd471859200;
      34976: inst = 32'd136314880;
      34977: inst = 32'd268468224;
      34978: inst = 32'd201343794;
      34979: inst = 32'd203423744;
      34980: inst = 32'd471859200;
      34981: inst = 32'd136314880;
      34982: inst = 32'd268468224;
      34983: inst = 32'd201343795;
      34984: inst = 32'd203423744;
      34985: inst = 32'd471859200;
      34986: inst = 32'd136314880;
      34987: inst = 32'd268468224;
      34988: inst = 32'd201343796;
      34989: inst = 32'd203423744;
      34990: inst = 32'd471859200;
      34991: inst = 32'd136314880;
      34992: inst = 32'd268468224;
      34993: inst = 32'd201343797;
      34994: inst = 32'd203423744;
      34995: inst = 32'd471859200;
      34996: inst = 32'd136314880;
      34997: inst = 32'd268468224;
      34998: inst = 32'd201343798;
      34999: inst = 32'd203423744;
      35000: inst = 32'd471859200;
      35001: inst = 32'd136314880;
      35002: inst = 32'd268468224;
      35003: inst = 32'd201343799;
      35004: inst = 32'd203423744;
      35005: inst = 32'd471859200;
      35006: inst = 32'd136314880;
      35007: inst = 32'd268468224;
      35008: inst = 32'd201343800;
      35009: inst = 32'd203423744;
      35010: inst = 32'd471859200;
      35011: inst = 32'd136314880;
      35012: inst = 32'd268468224;
      35013: inst = 32'd201343801;
      35014: inst = 32'd203423744;
      35015: inst = 32'd471859200;
      35016: inst = 32'd136314880;
      35017: inst = 32'd268468224;
      35018: inst = 32'd201343802;
      35019: inst = 32'd203423744;
      35020: inst = 32'd471859200;
      35021: inst = 32'd136314880;
      35022: inst = 32'd268468224;
      35023: inst = 32'd201343803;
      35024: inst = 32'd203423744;
      35025: inst = 32'd471859200;
      35026: inst = 32'd136314880;
      35027: inst = 32'd268468224;
      35028: inst = 32'd201343804;
      35029: inst = 32'd203423744;
      35030: inst = 32'd471859200;
      35031: inst = 32'd136314880;
      35032: inst = 32'd268468224;
      35033: inst = 32'd201343805;
      35034: inst = 32'd203423744;
      35035: inst = 32'd471859200;
      35036: inst = 32'd136314880;
      35037: inst = 32'd268468224;
      35038: inst = 32'd201343806;
      35039: inst = 32'd203423744;
      35040: inst = 32'd471859200;
      35041: inst = 32'd136314880;
      35042: inst = 32'd268468224;
      35043: inst = 32'd201343807;
      35044: inst = 32'd203423744;
      35045: inst = 32'd471859200;
      35046: inst = 32'd136314880;
      35047: inst = 32'd268468224;
      35048: inst = 32'd201343808;
      35049: inst = 32'd203423744;
      35050: inst = 32'd471859200;
      35051: inst = 32'd136314880;
      35052: inst = 32'd268468224;
      35053: inst = 32'd201343809;
      35054: inst = 32'd203423744;
      35055: inst = 32'd471859200;
      35056: inst = 32'd136314880;
      35057: inst = 32'd268468224;
      35058: inst = 32'd201343810;
      35059: inst = 32'd203423744;
      35060: inst = 32'd471859200;
      35061: inst = 32'd136314880;
      35062: inst = 32'd268468224;
      35063: inst = 32'd201343811;
      35064: inst = 32'd203423744;
      35065: inst = 32'd471859200;
      35066: inst = 32'd136314880;
      35067: inst = 32'd268468224;
      35068: inst = 32'd201343812;
      35069: inst = 32'd203423744;
      35070: inst = 32'd471859200;
      35071: inst = 32'd136314880;
      35072: inst = 32'd268468224;
      35073: inst = 32'd201343813;
      35074: inst = 32'd203423744;
      35075: inst = 32'd471859200;
      35076: inst = 32'd136314880;
      35077: inst = 32'd268468224;
      35078: inst = 32'd201343814;
      35079: inst = 32'd203423744;
      35080: inst = 32'd471859200;
      35081: inst = 32'd136314880;
      35082: inst = 32'd268468224;
      35083: inst = 32'd201343815;
      35084: inst = 32'd203423744;
      35085: inst = 32'd471859200;
      35086: inst = 32'd136314880;
      35087: inst = 32'd268468224;
      35088: inst = 32'd201343816;
      35089: inst = 32'd203423744;
      35090: inst = 32'd471859200;
      35091: inst = 32'd136314880;
      35092: inst = 32'd268468224;
      35093: inst = 32'd201343817;
      35094: inst = 32'd203423744;
      35095: inst = 32'd471859200;
      35096: inst = 32'd136314880;
      35097: inst = 32'd268468224;
      35098: inst = 32'd201343818;
      35099: inst = 32'd203423744;
      35100: inst = 32'd471859200;
      35101: inst = 32'd136314880;
      35102: inst = 32'd268468224;
      35103: inst = 32'd201343819;
      35104: inst = 32'd203423744;
      35105: inst = 32'd471859200;
      35106: inst = 32'd136314880;
      35107: inst = 32'd268468224;
      35108: inst = 32'd201343820;
      35109: inst = 32'd203423744;
      35110: inst = 32'd471859200;
      35111: inst = 32'd136314880;
      35112: inst = 32'd268468224;
      35113: inst = 32'd201343821;
      35114: inst = 32'd203423744;
      35115: inst = 32'd471859200;
      35116: inst = 32'd136314880;
      35117: inst = 32'd268468224;
      35118: inst = 32'd201343822;
      35119: inst = 32'd203423744;
      35120: inst = 32'd471859200;
      35121: inst = 32'd136314880;
      35122: inst = 32'd268468224;
      35123: inst = 32'd201343823;
      35124: inst = 32'd203423744;
      35125: inst = 32'd471859200;
      35126: inst = 32'd136314880;
      35127: inst = 32'd268468224;
      35128: inst = 32'd201343824;
      35129: inst = 32'd203423744;
      35130: inst = 32'd471859200;
      35131: inst = 32'd136314880;
      35132: inst = 32'd268468224;
      35133: inst = 32'd201343825;
      35134: inst = 32'd203423744;
      35135: inst = 32'd471859200;
      35136: inst = 32'd136314880;
      35137: inst = 32'd268468224;
      35138: inst = 32'd201343826;
      35139: inst = 32'd203423744;
      35140: inst = 32'd471859200;
      35141: inst = 32'd136314880;
      35142: inst = 32'd268468224;
      35143: inst = 32'd201343827;
      35144: inst = 32'd203423744;
      35145: inst = 32'd471859200;
      35146: inst = 32'd136314880;
      35147: inst = 32'd268468224;
      35148: inst = 32'd201343828;
      35149: inst = 32'd203423744;
      35150: inst = 32'd471859200;
      35151: inst = 32'd136314880;
      35152: inst = 32'd268468224;
      35153: inst = 32'd201343829;
      35154: inst = 32'd203423744;
      35155: inst = 32'd471859200;
      35156: inst = 32'd136314880;
      35157: inst = 32'd268468224;
      35158: inst = 32'd201343830;
      35159: inst = 32'd203423744;
      35160: inst = 32'd471859200;
      35161: inst = 32'd136314880;
      35162: inst = 32'd268468224;
      35163: inst = 32'd201343831;
      35164: inst = 32'd203423744;
      35165: inst = 32'd471859200;
      35166: inst = 32'd136314880;
      35167: inst = 32'd268468224;
      35168: inst = 32'd201343832;
      35169: inst = 32'd203423744;
      35170: inst = 32'd471859200;
      35171: inst = 32'd136314880;
      35172: inst = 32'd268468224;
      35173: inst = 32'd201343833;
      35174: inst = 32'd203423744;
      35175: inst = 32'd471859200;
      35176: inst = 32'd136314880;
      35177: inst = 32'd268468224;
      35178: inst = 32'd201343834;
      35179: inst = 32'd203423744;
      35180: inst = 32'd471859200;
      35181: inst = 32'd136314880;
      35182: inst = 32'd268468224;
      35183: inst = 32'd201343835;
      35184: inst = 32'd203423744;
      35185: inst = 32'd471859200;
      35186: inst = 32'd136314880;
      35187: inst = 32'd268468224;
      35188: inst = 32'd201343836;
      35189: inst = 32'd203423744;
      35190: inst = 32'd471859200;
      35191: inst = 32'd136314880;
      35192: inst = 32'd268468224;
      35193: inst = 32'd201343837;
      35194: inst = 32'd203423744;
      35195: inst = 32'd471859200;
      35196: inst = 32'd136314880;
      35197: inst = 32'd268468224;
      35198: inst = 32'd201343838;
      35199: inst = 32'd203423744;
      35200: inst = 32'd471859200;
      35201: inst = 32'd136314880;
      35202: inst = 32'd268468224;
      35203: inst = 32'd201343839;
      35204: inst = 32'd203423744;
      35205: inst = 32'd471859200;
      35206: inst = 32'd136314880;
      35207: inst = 32'd268468224;
      35208: inst = 32'd201343840;
      35209: inst = 32'd203423744;
      35210: inst = 32'd471859200;
      35211: inst = 32'd136314880;
      35212: inst = 32'd268468224;
      35213: inst = 32'd201343841;
      35214: inst = 32'd203423744;
      35215: inst = 32'd471859200;
      35216: inst = 32'd136314880;
      35217: inst = 32'd268468224;
      35218: inst = 32'd201343842;
      35219: inst = 32'd203423744;
      35220: inst = 32'd471859200;
      35221: inst = 32'd136314880;
      35222: inst = 32'd268468224;
      35223: inst = 32'd201343843;
      35224: inst = 32'd203423744;
      35225: inst = 32'd471859200;
      35226: inst = 32'd136314880;
      35227: inst = 32'd268468224;
      35228: inst = 32'd201343844;
      35229: inst = 32'd203423744;
      35230: inst = 32'd471859200;
      35231: inst = 32'd136314880;
      35232: inst = 32'd268468224;
      35233: inst = 32'd201343845;
      35234: inst = 32'd203423744;
      35235: inst = 32'd471859200;
      35236: inst = 32'd136314880;
      35237: inst = 32'd268468224;
      35238: inst = 32'd201343846;
      35239: inst = 32'd203423744;
      35240: inst = 32'd471859200;
      35241: inst = 32'd136314880;
      35242: inst = 32'd268468224;
      35243: inst = 32'd201343847;
      35244: inst = 32'd203423744;
      35245: inst = 32'd471859200;
      35246: inst = 32'd136314880;
      35247: inst = 32'd268468224;
      35248: inst = 32'd201343848;
      35249: inst = 32'd203423744;
      35250: inst = 32'd471859200;
      35251: inst = 32'd136314880;
      35252: inst = 32'd268468224;
      35253: inst = 32'd201343849;
      35254: inst = 32'd203423744;
      35255: inst = 32'd471859200;
      35256: inst = 32'd136314880;
      35257: inst = 32'd268468224;
      35258: inst = 32'd201343850;
      35259: inst = 32'd203423744;
      35260: inst = 32'd471859200;
      35261: inst = 32'd136314880;
      35262: inst = 32'd268468224;
      35263: inst = 32'd201343851;
      35264: inst = 32'd203423744;
      35265: inst = 32'd471859200;
      35266: inst = 32'd136314880;
      35267: inst = 32'd268468224;
      35268: inst = 32'd201343852;
      35269: inst = 32'd203423744;
      35270: inst = 32'd471859200;
      35271: inst = 32'd136314880;
      35272: inst = 32'd268468224;
      35273: inst = 32'd201343853;
      35274: inst = 32'd203423744;
      35275: inst = 32'd471859200;
      35276: inst = 32'd136314880;
      35277: inst = 32'd268468224;
      35278: inst = 32'd201343854;
      35279: inst = 32'd203423744;
      35280: inst = 32'd471859200;
      35281: inst = 32'd136314880;
      35282: inst = 32'd268468224;
      35283: inst = 32'd201343855;
      35284: inst = 32'd203423744;
      35285: inst = 32'd471859200;
      35286: inst = 32'd136314880;
      35287: inst = 32'd268468224;
      35288: inst = 32'd201343856;
      35289: inst = 32'd203423744;
      35290: inst = 32'd471859200;
      35291: inst = 32'd136314880;
      35292: inst = 32'd268468224;
      35293: inst = 32'd201343857;
      35294: inst = 32'd203423744;
      35295: inst = 32'd471859200;
      35296: inst = 32'd136314880;
      35297: inst = 32'd268468224;
      35298: inst = 32'd201343858;
      35299: inst = 32'd203423744;
      35300: inst = 32'd471859200;
      35301: inst = 32'd136314880;
      35302: inst = 32'd268468224;
      35303: inst = 32'd201343859;
      35304: inst = 32'd203423744;
      35305: inst = 32'd471859200;
      35306: inst = 32'd136314880;
      35307: inst = 32'd268468224;
      35308: inst = 32'd201343860;
      35309: inst = 32'd203423744;
      35310: inst = 32'd471859200;
      35311: inst = 32'd136314880;
      35312: inst = 32'd268468224;
      35313: inst = 32'd201343861;
      35314: inst = 32'd203423744;
      35315: inst = 32'd471859200;
      35316: inst = 32'd136314880;
      35317: inst = 32'd268468224;
      35318: inst = 32'd201343862;
      35319: inst = 32'd203423744;
      35320: inst = 32'd471859200;
      35321: inst = 32'd136314880;
      35322: inst = 32'd268468224;
      35323: inst = 32'd201343863;
      35324: inst = 32'd203423744;
      35325: inst = 32'd471859200;
      35326: inst = 32'd136314880;
      35327: inst = 32'd268468224;
      35328: inst = 32'd201343864;
      35329: inst = 32'd203423744;
      35330: inst = 32'd471859200;
      35331: inst = 32'd136314880;
      35332: inst = 32'd268468224;
      35333: inst = 32'd201343865;
      35334: inst = 32'd203423744;
      35335: inst = 32'd471859200;
      35336: inst = 32'd136314880;
      35337: inst = 32'd268468224;
      35338: inst = 32'd201343866;
      35339: inst = 32'd203423744;
      35340: inst = 32'd471859200;
      35341: inst = 32'd136314880;
      35342: inst = 32'd268468224;
      35343: inst = 32'd201343867;
      35344: inst = 32'd203423744;
      35345: inst = 32'd471859200;
      35346: inst = 32'd136314880;
      35347: inst = 32'd268468224;
      35348: inst = 32'd201343868;
      35349: inst = 32'd203423744;
      35350: inst = 32'd471859200;
      35351: inst = 32'd136314880;
      35352: inst = 32'd268468224;
      35353: inst = 32'd201343869;
      35354: inst = 32'd203423744;
      35355: inst = 32'd471859200;
      35356: inst = 32'd136314880;
      35357: inst = 32'd268468224;
      35358: inst = 32'd201343870;
      35359: inst = 32'd203423744;
      35360: inst = 32'd471859200;
      35361: inst = 32'd136314880;
      35362: inst = 32'd268468224;
      35363: inst = 32'd201343871;
      35364: inst = 32'd203423744;
      35365: inst = 32'd471859200;
      35366: inst = 32'd136314880;
      35367: inst = 32'd268468224;
      35368: inst = 32'd201343872;
      35369: inst = 32'd203423744;
      35370: inst = 32'd471859200;
      35371: inst = 32'd136314880;
      35372: inst = 32'd268468224;
      35373: inst = 32'd201343873;
      35374: inst = 32'd203423744;
      35375: inst = 32'd471859200;
      35376: inst = 32'd136314880;
      35377: inst = 32'd268468224;
      35378: inst = 32'd201343874;
      35379: inst = 32'd203423744;
      35380: inst = 32'd471859200;
      35381: inst = 32'd136314880;
      35382: inst = 32'd268468224;
      35383: inst = 32'd201343875;
      35384: inst = 32'd203423744;
      35385: inst = 32'd471859200;
      35386: inst = 32'd136314880;
      35387: inst = 32'd268468224;
      35388: inst = 32'd201343876;
      35389: inst = 32'd203423744;
      35390: inst = 32'd471859200;
      35391: inst = 32'd136314880;
      35392: inst = 32'd268468224;
      35393: inst = 32'd201343877;
      35394: inst = 32'd203423744;
      35395: inst = 32'd471859200;
      35396: inst = 32'd136314880;
      35397: inst = 32'd268468224;
      35398: inst = 32'd201343878;
      35399: inst = 32'd203423744;
      35400: inst = 32'd471859200;
      35401: inst = 32'd136314880;
      35402: inst = 32'd268468224;
      35403: inst = 32'd201343879;
      35404: inst = 32'd203423744;
      35405: inst = 32'd471859200;
      35406: inst = 32'd136314880;
      35407: inst = 32'd268468224;
      35408: inst = 32'd201343880;
      35409: inst = 32'd203423744;
      35410: inst = 32'd471859200;
      35411: inst = 32'd136314880;
      35412: inst = 32'd268468224;
      35413: inst = 32'd201343881;
      35414: inst = 32'd203423744;
      35415: inst = 32'd471859200;
      35416: inst = 32'd136314880;
      35417: inst = 32'd268468224;
      35418: inst = 32'd201343882;
      35419: inst = 32'd203423744;
      35420: inst = 32'd471859200;
      35421: inst = 32'd136314880;
      35422: inst = 32'd268468224;
      35423: inst = 32'd201343883;
      35424: inst = 32'd203423744;
      35425: inst = 32'd471859200;
      35426: inst = 32'd136314880;
      35427: inst = 32'd268468224;
      35428: inst = 32'd201343884;
      35429: inst = 32'd203423744;
      35430: inst = 32'd471859200;
      35431: inst = 32'd136314880;
      35432: inst = 32'd268468224;
      35433: inst = 32'd201343885;
      35434: inst = 32'd203423744;
      35435: inst = 32'd471859200;
      35436: inst = 32'd136314880;
      35437: inst = 32'd268468224;
      35438: inst = 32'd201343886;
      35439: inst = 32'd203423744;
      35440: inst = 32'd471859200;
      35441: inst = 32'd136314880;
      35442: inst = 32'd268468224;
      35443: inst = 32'd201343887;
      35444: inst = 32'd203423744;
      35445: inst = 32'd471859200;
      35446: inst = 32'd136314880;
      35447: inst = 32'd268468224;
      35448: inst = 32'd201343888;
      35449: inst = 32'd203423744;
      35450: inst = 32'd471859200;
      35451: inst = 32'd136314880;
      35452: inst = 32'd268468224;
      35453: inst = 32'd201343889;
      35454: inst = 32'd203423744;
      35455: inst = 32'd471859200;
      35456: inst = 32'd136314880;
      35457: inst = 32'd268468224;
      35458: inst = 32'd201343890;
      35459: inst = 32'd203423744;
      35460: inst = 32'd471859200;
      35461: inst = 32'd136314880;
      35462: inst = 32'd268468224;
      35463: inst = 32'd201343891;
      35464: inst = 32'd203423744;
      35465: inst = 32'd471859200;
      35466: inst = 32'd136314880;
      35467: inst = 32'd268468224;
      35468: inst = 32'd201343892;
      35469: inst = 32'd203423744;
      35470: inst = 32'd471859200;
      35471: inst = 32'd136314880;
      35472: inst = 32'd268468224;
      35473: inst = 32'd201343893;
      35474: inst = 32'd203423744;
      35475: inst = 32'd471859200;
      35476: inst = 32'd136314880;
      35477: inst = 32'd268468224;
      35478: inst = 32'd201343894;
      35479: inst = 32'd203423744;
      35480: inst = 32'd471859200;
      35481: inst = 32'd136314880;
      35482: inst = 32'd268468224;
      35483: inst = 32'd201343895;
      35484: inst = 32'd203423744;
      35485: inst = 32'd471859200;
      35486: inst = 32'd136314880;
      35487: inst = 32'd268468224;
      35488: inst = 32'd201343896;
      35489: inst = 32'd203423744;
      35490: inst = 32'd471859200;
      35491: inst = 32'd136314880;
      35492: inst = 32'd268468224;
      35493: inst = 32'd201343897;
      35494: inst = 32'd203423744;
      35495: inst = 32'd471859200;
      35496: inst = 32'd136314880;
      35497: inst = 32'd268468224;
      35498: inst = 32'd201343898;
      35499: inst = 32'd203423744;
      35500: inst = 32'd471859200;
      35501: inst = 32'd136314880;
      35502: inst = 32'd268468224;
      35503: inst = 32'd201343899;
      35504: inst = 32'd203423744;
      35505: inst = 32'd471859200;
      35506: inst = 32'd136314880;
      35507: inst = 32'd268468224;
      35508: inst = 32'd201343900;
      35509: inst = 32'd203423744;
      35510: inst = 32'd471859200;
      35511: inst = 32'd136314880;
      35512: inst = 32'd268468224;
      35513: inst = 32'd201343901;
      35514: inst = 32'd203423744;
      35515: inst = 32'd471859200;
      35516: inst = 32'd136314880;
      35517: inst = 32'd268468224;
      35518: inst = 32'd201343902;
      35519: inst = 32'd203423744;
      35520: inst = 32'd471859200;
      35521: inst = 32'd136314880;
      35522: inst = 32'd268468224;
      35523: inst = 32'd201343903;
      35524: inst = 32'd203423744;
      35525: inst = 32'd471859200;
      35526: inst = 32'd136314880;
      35527: inst = 32'd268468224;
      35528: inst = 32'd201343904;
      35529: inst = 32'd203423744;
      35530: inst = 32'd471859200;
      35531: inst = 32'd136314880;
      35532: inst = 32'd268468224;
      35533: inst = 32'd201343905;
      35534: inst = 32'd203423744;
      35535: inst = 32'd471859200;
      35536: inst = 32'd136314880;
      35537: inst = 32'd268468224;
      35538: inst = 32'd201343906;
      35539: inst = 32'd203423744;
      35540: inst = 32'd471859200;
      35541: inst = 32'd136314880;
      35542: inst = 32'd268468224;
      35543: inst = 32'd201343907;
      35544: inst = 32'd203423744;
      35545: inst = 32'd471859200;
      35546: inst = 32'd136314880;
      35547: inst = 32'd268468224;
      35548: inst = 32'd201343908;
      35549: inst = 32'd203423744;
      35550: inst = 32'd471859200;
      35551: inst = 32'd136314880;
      35552: inst = 32'd268468224;
      35553: inst = 32'd201343909;
      35554: inst = 32'd203423744;
      35555: inst = 32'd471859200;
      35556: inst = 32'd136314880;
      35557: inst = 32'd268468224;
      35558: inst = 32'd201343910;
      35559: inst = 32'd203423744;
      35560: inst = 32'd471859200;
      35561: inst = 32'd136314880;
      35562: inst = 32'd268468224;
      35563: inst = 32'd201343911;
      35564: inst = 32'd203423744;
      35565: inst = 32'd471859200;
      35566: inst = 32'd136314880;
      35567: inst = 32'd268468224;
      35568: inst = 32'd201343912;
      35569: inst = 32'd203423744;
      35570: inst = 32'd471859200;
      35571: inst = 32'd136314880;
      35572: inst = 32'd268468224;
      35573: inst = 32'd201343913;
      35574: inst = 32'd203423744;
      35575: inst = 32'd471859200;
      35576: inst = 32'd136314880;
      35577: inst = 32'd268468224;
      35578: inst = 32'd201343914;
      35579: inst = 32'd203423744;
      35580: inst = 32'd471859200;
      35581: inst = 32'd136314880;
      35582: inst = 32'd268468224;
      35583: inst = 32'd201343915;
      35584: inst = 32'd203423744;
      35585: inst = 32'd471859200;
      35586: inst = 32'd136314880;
      35587: inst = 32'd268468224;
      35588: inst = 32'd201343916;
      35589: inst = 32'd203423744;
      35590: inst = 32'd471859200;
      35591: inst = 32'd136314880;
      35592: inst = 32'd268468224;
      35593: inst = 32'd201343917;
      35594: inst = 32'd203423744;
      35595: inst = 32'd471859200;
      35596: inst = 32'd136314880;
      35597: inst = 32'd268468224;
      35598: inst = 32'd201343918;
      35599: inst = 32'd203423744;
      35600: inst = 32'd471859200;
      35601: inst = 32'd136314880;
      35602: inst = 32'd268468224;
      35603: inst = 32'd201343919;
      35604: inst = 32'd203423744;
      35605: inst = 32'd471859200;
      35606: inst = 32'd136314880;
      35607: inst = 32'd268468224;
      35608: inst = 32'd201343920;
      35609: inst = 32'd203423744;
      35610: inst = 32'd471859200;
      35611: inst = 32'd136314880;
      35612: inst = 32'd268468224;
      35613: inst = 32'd201343921;
      35614: inst = 32'd203423744;
      35615: inst = 32'd471859200;
      35616: inst = 32'd136314880;
      35617: inst = 32'd268468224;
      35618: inst = 32'd201343922;
      35619: inst = 32'd203423744;
      35620: inst = 32'd471859200;
      35621: inst = 32'd136314880;
      35622: inst = 32'd268468224;
      35623: inst = 32'd201343923;
      35624: inst = 32'd203423744;
      35625: inst = 32'd471859200;
      35626: inst = 32'd136314880;
      35627: inst = 32'd268468224;
      35628: inst = 32'd201343924;
      35629: inst = 32'd203423744;
      35630: inst = 32'd471859200;
      35631: inst = 32'd136314880;
      35632: inst = 32'd268468224;
      35633: inst = 32'd201343925;
      35634: inst = 32'd203423744;
      35635: inst = 32'd471859200;
      35636: inst = 32'd136314880;
      35637: inst = 32'd268468224;
      35638: inst = 32'd201343926;
      35639: inst = 32'd203423744;
      35640: inst = 32'd471859200;
      35641: inst = 32'd136314880;
      35642: inst = 32'd268468224;
      35643: inst = 32'd201343927;
      35644: inst = 32'd203423744;
      35645: inst = 32'd471859200;
      35646: inst = 32'd136314880;
      35647: inst = 32'd268468224;
      35648: inst = 32'd201343928;
      35649: inst = 32'd203423744;
      35650: inst = 32'd471859200;
      35651: inst = 32'd136314880;
      35652: inst = 32'd268468224;
      35653: inst = 32'd201343929;
      35654: inst = 32'd203423744;
      35655: inst = 32'd471859200;
      35656: inst = 32'd136314880;
      35657: inst = 32'd268468224;
      35658: inst = 32'd201343930;
      35659: inst = 32'd203423744;
      35660: inst = 32'd471859200;
      35661: inst = 32'd136314880;
      35662: inst = 32'd268468224;
      35663: inst = 32'd201343931;
      35664: inst = 32'd203423744;
      35665: inst = 32'd471859200;
      35666: inst = 32'd136314880;
      35667: inst = 32'd268468224;
      35668: inst = 32'd201343932;
      35669: inst = 32'd203423744;
      35670: inst = 32'd471859200;
      35671: inst = 32'd136314880;
      35672: inst = 32'd268468224;
      35673: inst = 32'd201343933;
      35674: inst = 32'd203423744;
      35675: inst = 32'd471859200;
      35676: inst = 32'd136314880;
      35677: inst = 32'd268468224;
      35678: inst = 32'd201343934;
      35679: inst = 32'd203423744;
      35680: inst = 32'd471859200;
      35681: inst = 32'd136314880;
      35682: inst = 32'd268468224;
      35683: inst = 32'd201343935;
      35684: inst = 32'd203423744;
      35685: inst = 32'd471859200;
      35686: inst = 32'd136314880;
      35687: inst = 32'd268468224;
      35688: inst = 32'd201343936;
      35689: inst = 32'd203423744;
      35690: inst = 32'd471859200;
      35691: inst = 32'd136314880;
      35692: inst = 32'd268468224;
      35693: inst = 32'd201343937;
      35694: inst = 32'd203423744;
      35695: inst = 32'd471859200;
      35696: inst = 32'd136314880;
      35697: inst = 32'd268468224;
      35698: inst = 32'd201343938;
      35699: inst = 32'd203423744;
      35700: inst = 32'd471859200;
      35701: inst = 32'd136314880;
      35702: inst = 32'd268468224;
      35703: inst = 32'd201343939;
      35704: inst = 32'd203423744;
      35705: inst = 32'd471859200;
      35706: inst = 32'd136314880;
      35707: inst = 32'd268468224;
      35708: inst = 32'd201343940;
      35709: inst = 32'd203423744;
      35710: inst = 32'd471859200;
      35711: inst = 32'd136314880;
      35712: inst = 32'd268468224;
      35713: inst = 32'd201343941;
      35714: inst = 32'd203423744;
      35715: inst = 32'd471859200;
      35716: inst = 32'd136314880;
      35717: inst = 32'd268468224;
      35718: inst = 32'd201343942;
      35719: inst = 32'd203423744;
      35720: inst = 32'd471859200;
      35721: inst = 32'd136314880;
      35722: inst = 32'd268468224;
      35723: inst = 32'd201343943;
      35724: inst = 32'd203423744;
      35725: inst = 32'd471859200;
      35726: inst = 32'd136314880;
      35727: inst = 32'd268468224;
      35728: inst = 32'd201343944;
      35729: inst = 32'd203423744;
      35730: inst = 32'd471859200;
      35731: inst = 32'd136314880;
      35732: inst = 32'd268468224;
      35733: inst = 32'd201343945;
      35734: inst = 32'd203423744;
      35735: inst = 32'd471859200;
      35736: inst = 32'd136314880;
      35737: inst = 32'd268468224;
      35738: inst = 32'd201343946;
      35739: inst = 32'd203423744;
      35740: inst = 32'd471859200;
      35741: inst = 32'd136314880;
      35742: inst = 32'd268468224;
      35743: inst = 32'd201343947;
      35744: inst = 32'd203423744;
      35745: inst = 32'd471859200;
      35746: inst = 32'd136314880;
      35747: inst = 32'd268468224;
      35748: inst = 32'd201343948;
      35749: inst = 32'd203423744;
      35750: inst = 32'd471859200;
      35751: inst = 32'd136314880;
      35752: inst = 32'd268468224;
      35753: inst = 32'd201343949;
      35754: inst = 32'd203423744;
      35755: inst = 32'd471859200;
      35756: inst = 32'd136314880;
      35757: inst = 32'd268468224;
      35758: inst = 32'd201343950;
      35759: inst = 32'd203423744;
      35760: inst = 32'd471859200;
      35761: inst = 32'd136314880;
      35762: inst = 32'd268468224;
      35763: inst = 32'd201343951;
      35764: inst = 32'd203423744;
      35765: inst = 32'd471859200;
      35766: inst = 32'd136314880;
      35767: inst = 32'd268468224;
      35768: inst = 32'd201343952;
      35769: inst = 32'd203423744;
      35770: inst = 32'd471859200;
      35771: inst = 32'd136314880;
      35772: inst = 32'd268468224;
      35773: inst = 32'd201343953;
      35774: inst = 32'd203423744;
      35775: inst = 32'd471859200;
      35776: inst = 32'd136314880;
      35777: inst = 32'd268468224;
      35778: inst = 32'd201343954;
      35779: inst = 32'd203423744;
      35780: inst = 32'd471859200;
      35781: inst = 32'd136314880;
      35782: inst = 32'd268468224;
      35783: inst = 32'd201343955;
      35784: inst = 32'd203423744;
      35785: inst = 32'd471859200;
      35786: inst = 32'd136314880;
      35787: inst = 32'd268468224;
      35788: inst = 32'd201343956;
      35789: inst = 32'd203423744;
      35790: inst = 32'd471859200;
      35791: inst = 32'd136314880;
      35792: inst = 32'd268468224;
      35793: inst = 32'd201343957;
      35794: inst = 32'd203423744;
      35795: inst = 32'd471859200;
      35796: inst = 32'd136314880;
      35797: inst = 32'd268468224;
      35798: inst = 32'd201343958;
      35799: inst = 32'd203423744;
      35800: inst = 32'd471859200;
      35801: inst = 32'd136314880;
      35802: inst = 32'd268468224;
      35803: inst = 32'd201343959;
      35804: inst = 32'd203423744;
      35805: inst = 32'd471859200;
      35806: inst = 32'd136314880;
      35807: inst = 32'd268468224;
      35808: inst = 32'd201343960;
      35809: inst = 32'd203423744;
      35810: inst = 32'd471859200;
      35811: inst = 32'd136314880;
      35812: inst = 32'd268468224;
      35813: inst = 32'd201343961;
      35814: inst = 32'd203423744;
      35815: inst = 32'd471859200;
      35816: inst = 32'd136314880;
      35817: inst = 32'd268468224;
      35818: inst = 32'd201343962;
      35819: inst = 32'd203423744;
      35820: inst = 32'd471859200;
      35821: inst = 32'd136314880;
      35822: inst = 32'd268468224;
      35823: inst = 32'd201343963;
      35824: inst = 32'd203423744;
      35825: inst = 32'd471859200;
      35826: inst = 32'd136314880;
      35827: inst = 32'd268468224;
      35828: inst = 32'd201343964;
      35829: inst = 32'd203423744;
      35830: inst = 32'd471859200;
      35831: inst = 32'd136314880;
      35832: inst = 32'd268468224;
      35833: inst = 32'd201343965;
      35834: inst = 32'd203423744;
      35835: inst = 32'd471859200;
      35836: inst = 32'd136314880;
      35837: inst = 32'd268468224;
      35838: inst = 32'd201343966;
      35839: inst = 32'd203423744;
      35840: inst = 32'd471859200;
      35841: inst = 32'd136314880;
      35842: inst = 32'd268468224;
      35843: inst = 32'd201343967;
      35844: inst = 32'd203423744;
      35845: inst = 32'd471859200;
      35846: inst = 32'd136314880;
      35847: inst = 32'd268468224;
      35848: inst = 32'd201343968;
      35849: inst = 32'd203423744;
      35850: inst = 32'd471859200;
      35851: inst = 32'd136314880;
      35852: inst = 32'd268468224;
      35853: inst = 32'd201343969;
      35854: inst = 32'd203423744;
      35855: inst = 32'd471859200;
      35856: inst = 32'd136314880;
      35857: inst = 32'd268468224;
      35858: inst = 32'd201343970;
      35859: inst = 32'd203423744;
      35860: inst = 32'd471859200;
      35861: inst = 32'd136314880;
      35862: inst = 32'd268468224;
      35863: inst = 32'd201343971;
      35864: inst = 32'd203423744;
      35865: inst = 32'd471859200;
      35866: inst = 32'd136314880;
      35867: inst = 32'd268468224;
      35868: inst = 32'd201343972;
      35869: inst = 32'd203423744;
      35870: inst = 32'd471859200;
      35871: inst = 32'd136314880;
      35872: inst = 32'd268468224;
      35873: inst = 32'd201343973;
      35874: inst = 32'd203423744;
      35875: inst = 32'd471859200;
      35876: inst = 32'd136314880;
      35877: inst = 32'd268468224;
      35878: inst = 32'd201343974;
      35879: inst = 32'd203423744;
      35880: inst = 32'd471859200;
      35881: inst = 32'd136314880;
      35882: inst = 32'd268468224;
      35883: inst = 32'd201343975;
      35884: inst = 32'd203423744;
      35885: inst = 32'd471859200;
      35886: inst = 32'd136314880;
      35887: inst = 32'd268468224;
      35888: inst = 32'd201343976;
      35889: inst = 32'd203423744;
      35890: inst = 32'd471859200;
      35891: inst = 32'd136314880;
      35892: inst = 32'd268468224;
      35893: inst = 32'd201343977;
      35894: inst = 32'd203423744;
      35895: inst = 32'd471859200;
      35896: inst = 32'd136314880;
      35897: inst = 32'd268468224;
      35898: inst = 32'd201343978;
      35899: inst = 32'd203423744;
      35900: inst = 32'd471859200;
      35901: inst = 32'd136314880;
      35902: inst = 32'd268468224;
      35903: inst = 32'd201343979;
      35904: inst = 32'd203423744;
      35905: inst = 32'd471859200;
      35906: inst = 32'd136314880;
      35907: inst = 32'd268468224;
      35908: inst = 32'd201343980;
      35909: inst = 32'd203423744;
      35910: inst = 32'd471859200;
      35911: inst = 32'd136314880;
      35912: inst = 32'd268468224;
      35913: inst = 32'd201343981;
      35914: inst = 32'd203423744;
      35915: inst = 32'd471859200;
      35916: inst = 32'd136314880;
      35917: inst = 32'd268468224;
      35918: inst = 32'd201343982;
      35919: inst = 32'd203423744;
      35920: inst = 32'd471859200;
      35921: inst = 32'd136314880;
      35922: inst = 32'd268468224;
      35923: inst = 32'd201343983;
      35924: inst = 32'd203423744;
      35925: inst = 32'd471859200;
      35926: inst = 32'd136314880;
      35927: inst = 32'd268468224;
      35928: inst = 32'd201343984;
      35929: inst = 32'd203423744;
      35930: inst = 32'd471859200;
      35931: inst = 32'd136314880;
      35932: inst = 32'd268468224;
      35933: inst = 32'd201343985;
      35934: inst = 32'd203423744;
      35935: inst = 32'd471859200;
      35936: inst = 32'd136314880;
      35937: inst = 32'd268468224;
      35938: inst = 32'd201343986;
      35939: inst = 32'd203423744;
      35940: inst = 32'd471859200;
      35941: inst = 32'd136314880;
      35942: inst = 32'd268468224;
      35943: inst = 32'd201343987;
      35944: inst = 32'd203423744;
      35945: inst = 32'd471859200;
      35946: inst = 32'd136314880;
      35947: inst = 32'd268468224;
      35948: inst = 32'd201343988;
      35949: inst = 32'd203423744;
      35950: inst = 32'd471859200;
      35951: inst = 32'd136314880;
      35952: inst = 32'd268468224;
      35953: inst = 32'd201343989;
      35954: inst = 32'd203423744;
      35955: inst = 32'd471859200;
      35956: inst = 32'd136314880;
      35957: inst = 32'd268468224;
      35958: inst = 32'd201343990;
      35959: inst = 32'd203423744;
      35960: inst = 32'd471859200;
      35961: inst = 32'd136314880;
      35962: inst = 32'd268468224;
      35963: inst = 32'd201343991;
      35964: inst = 32'd203423744;
      35965: inst = 32'd471859200;
      35966: inst = 32'd136314880;
      35967: inst = 32'd268468224;
      35968: inst = 32'd201343992;
      35969: inst = 32'd203423744;
      35970: inst = 32'd471859200;
      35971: inst = 32'd136314880;
      35972: inst = 32'd268468224;
      35973: inst = 32'd201343993;
      35974: inst = 32'd203423744;
      35975: inst = 32'd471859200;
      35976: inst = 32'd136314880;
      35977: inst = 32'd268468224;
      35978: inst = 32'd201343994;
      35979: inst = 32'd203423744;
      35980: inst = 32'd471859200;
      35981: inst = 32'd136314880;
      35982: inst = 32'd268468224;
      35983: inst = 32'd201343995;
      35984: inst = 32'd203423744;
      35985: inst = 32'd471859200;
      35986: inst = 32'd136314880;
      35987: inst = 32'd268468224;
      35988: inst = 32'd201343996;
      35989: inst = 32'd203423744;
      35990: inst = 32'd471859200;
      35991: inst = 32'd136314880;
      35992: inst = 32'd268468224;
      35993: inst = 32'd201343997;
      35994: inst = 32'd203423744;
      35995: inst = 32'd471859200;
      35996: inst = 32'd136314880;
      35997: inst = 32'd268468224;
      35998: inst = 32'd201343998;
      35999: inst = 32'd203423744;
      36000: inst = 32'd471859200;
      36001: inst = 32'd136314880;
      36002: inst = 32'd268468224;
      36003: inst = 32'd201343999;
      36004: inst = 32'd203423744;
      36005: inst = 32'd471859200;
      36006: inst = 32'd136314880;
      36007: inst = 32'd268468224;
      36008: inst = 32'd201344000;
      36009: inst = 32'd203423744;
      36010: inst = 32'd471859200;
      36011: inst = 32'd136314880;
      36012: inst = 32'd268468224;
      36013: inst = 32'd201344001;
      36014: inst = 32'd203423744;
      36015: inst = 32'd471859200;
      36016: inst = 32'd136314880;
      36017: inst = 32'd268468224;
      36018: inst = 32'd201344002;
      36019: inst = 32'd203423744;
      36020: inst = 32'd471859200;
      36021: inst = 32'd136314880;
      36022: inst = 32'd268468224;
      36023: inst = 32'd201344003;
      36024: inst = 32'd203423744;
      36025: inst = 32'd471859200;
      36026: inst = 32'd136314880;
      36027: inst = 32'd268468224;
      36028: inst = 32'd201344004;
      36029: inst = 32'd203423744;
      36030: inst = 32'd471859200;
      36031: inst = 32'd136314880;
      36032: inst = 32'd268468224;
      36033: inst = 32'd201344005;
      36034: inst = 32'd203423744;
      36035: inst = 32'd471859200;
      36036: inst = 32'd136314880;
      36037: inst = 32'd268468224;
      36038: inst = 32'd201344006;
      36039: inst = 32'd203423744;
      36040: inst = 32'd471859200;
      36041: inst = 32'd136314880;
      36042: inst = 32'd268468224;
      36043: inst = 32'd201344007;
      36044: inst = 32'd203423744;
      36045: inst = 32'd471859200;
      36046: inst = 32'd136314880;
      36047: inst = 32'd268468224;
      36048: inst = 32'd201344008;
      36049: inst = 32'd203423744;
      36050: inst = 32'd471859200;
      36051: inst = 32'd136314880;
      36052: inst = 32'd268468224;
      36053: inst = 32'd201344009;
      36054: inst = 32'd203423744;
      36055: inst = 32'd471859200;
      36056: inst = 32'd136314880;
      36057: inst = 32'd268468224;
      36058: inst = 32'd201344010;
      36059: inst = 32'd203423744;
      36060: inst = 32'd471859200;
      36061: inst = 32'd136314880;
      36062: inst = 32'd268468224;
      36063: inst = 32'd201344011;
      36064: inst = 32'd203423744;
      36065: inst = 32'd471859200;
      36066: inst = 32'd136314880;
      36067: inst = 32'd268468224;
      36068: inst = 32'd201344012;
      36069: inst = 32'd203423744;
      36070: inst = 32'd471859200;
      36071: inst = 32'd136314880;
      36072: inst = 32'd268468224;
      36073: inst = 32'd201344013;
      36074: inst = 32'd203423744;
      36075: inst = 32'd471859200;
      36076: inst = 32'd136314880;
      36077: inst = 32'd268468224;
      36078: inst = 32'd201344014;
      36079: inst = 32'd203423744;
      36080: inst = 32'd471859200;
      36081: inst = 32'd136314880;
      36082: inst = 32'd268468224;
      36083: inst = 32'd201344015;
      36084: inst = 32'd203423744;
      36085: inst = 32'd471859200;
      36086: inst = 32'd136314880;
      36087: inst = 32'd268468224;
      36088: inst = 32'd201344016;
      36089: inst = 32'd203423744;
      36090: inst = 32'd471859200;
      36091: inst = 32'd136314880;
      36092: inst = 32'd268468224;
      36093: inst = 32'd201344017;
      36094: inst = 32'd203423744;
      36095: inst = 32'd471859200;
      36096: inst = 32'd136314880;
      36097: inst = 32'd268468224;
      36098: inst = 32'd201344018;
      36099: inst = 32'd203423744;
      36100: inst = 32'd471859200;
      36101: inst = 32'd136314880;
      36102: inst = 32'd268468224;
      36103: inst = 32'd201344019;
      36104: inst = 32'd203423744;
      36105: inst = 32'd471859200;
      36106: inst = 32'd136314880;
      36107: inst = 32'd268468224;
      36108: inst = 32'd201344020;
      36109: inst = 32'd203423744;
      36110: inst = 32'd471859200;
      36111: inst = 32'd136314880;
      36112: inst = 32'd268468224;
      36113: inst = 32'd201344021;
      36114: inst = 32'd203423744;
      36115: inst = 32'd471859200;
      36116: inst = 32'd136314880;
      36117: inst = 32'd268468224;
      36118: inst = 32'd201344022;
      36119: inst = 32'd203423744;
      36120: inst = 32'd471859200;
      36121: inst = 32'd136314880;
      36122: inst = 32'd268468224;
      36123: inst = 32'd201344023;
      36124: inst = 32'd203423744;
      36125: inst = 32'd471859200;
      36126: inst = 32'd136314880;
      36127: inst = 32'd268468224;
      36128: inst = 32'd201344024;
      36129: inst = 32'd203423744;
      36130: inst = 32'd471859200;
      36131: inst = 32'd136314880;
      36132: inst = 32'd268468224;
      36133: inst = 32'd201344025;
      36134: inst = 32'd203423744;
      36135: inst = 32'd471859200;
      36136: inst = 32'd136314880;
      36137: inst = 32'd268468224;
      36138: inst = 32'd201344026;
      36139: inst = 32'd203423744;
      36140: inst = 32'd471859200;
      36141: inst = 32'd136314880;
      36142: inst = 32'd268468224;
      36143: inst = 32'd201344027;
      36144: inst = 32'd203423744;
      36145: inst = 32'd471859200;
      36146: inst = 32'd136314880;
      36147: inst = 32'd268468224;
      36148: inst = 32'd201344028;
      36149: inst = 32'd203423744;
      36150: inst = 32'd471859200;
      36151: inst = 32'd136314880;
      36152: inst = 32'd268468224;
      36153: inst = 32'd201344029;
      36154: inst = 32'd203423744;
      36155: inst = 32'd471859200;
      36156: inst = 32'd136314880;
      36157: inst = 32'd268468224;
      36158: inst = 32'd201344030;
      36159: inst = 32'd203423744;
      36160: inst = 32'd471859200;
      36161: inst = 32'd136314880;
      36162: inst = 32'd268468224;
      36163: inst = 32'd201344031;
      36164: inst = 32'd203423744;
      36165: inst = 32'd471859200;
      36166: inst = 32'd136314880;
      36167: inst = 32'd268468224;
      36168: inst = 32'd201344032;
      36169: inst = 32'd203423744;
      36170: inst = 32'd471859200;
      36171: inst = 32'd136314880;
      36172: inst = 32'd268468224;
      36173: inst = 32'd201344033;
      36174: inst = 32'd203423744;
      36175: inst = 32'd471859200;
      36176: inst = 32'd136314880;
      36177: inst = 32'd268468224;
      36178: inst = 32'd201344034;
      36179: inst = 32'd203423744;
      36180: inst = 32'd471859200;
      36181: inst = 32'd136314880;
      36182: inst = 32'd268468224;
      36183: inst = 32'd201344035;
      36184: inst = 32'd203423744;
      36185: inst = 32'd471859200;
      36186: inst = 32'd136314880;
      36187: inst = 32'd268468224;
      36188: inst = 32'd201344036;
      36189: inst = 32'd203423744;
      36190: inst = 32'd471859200;
      36191: inst = 32'd136314880;
      36192: inst = 32'd268468224;
      36193: inst = 32'd201344037;
      36194: inst = 32'd203423744;
      36195: inst = 32'd471859200;
      36196: inst = 32'd136314880;
      36197: inst = 32'd268468224;
      36198: inst = 32'd201344038;
      36199: inst = 32'd203423744;
      36200: inst = 32'd471859200;
      36201: inst = 32'd136314880;
      36202: inst = 32'd268468224;
      36203: inst = 32'd201344039;
      36204: inst = 32'd203423744;
      36205: inst = 32'd471859200;
      36206: inst = 32'd136314880;
      36207: inst = 32'd268468224;
      36208: inst = 32'd201344040;
      36209: inst = 32'd203423744;
      36210: inst = 32'd471859200;
      36211: inst = 32'd136314880;
      36212: inst = 32'd268468224;
      36213: inst = 32'd201344041;
      36214: inst = 32'd203423744;
      36215: inst = 32'd471859200;
      36216: inst = 32'd136314880;
      36217: inst = 32'd268468224;
      36218: inst = 32'd201344042;
      36219: inst = 32'd203423744;
      36220: inst = 32'd471859200;
      36221: inst = 32'd136314880;
      36222: inst = 32'd268468224;
      36223: inst = 32'd201344043;
      36224: inst = 32'd203423744;
      36225: inst = 32'd471859200;
      36226: inst = 32'd136314880;
      36227: inst = 32'd268468224;
      36228: inst = 32'd201344044;
      36229: inst = 32'd203423744;
      36230: inst = 32'd471859200;
      36231: inst = 32'd136314880;
      36232: inst = 32'd268468224;
      36233: inst = 32'd201344045;
      36234: inst = 32'd203423744;
      36235: inst = 32'd471859200;
      36236: inst = 32'd136314880;
      36237: inst = 32'd268468224;
      36238: inst = 32'd201344046;
      36239: inst = 32'd203423744;
      36240: inst = 32'd471859200;
      36241: inst = 32'd136314880;
      36242: inst = 32'd268468224;
      36243: inst = 32'd201344047;
      36244: inst = 32'd203423744;
      36245: inst = 32'd471859200;
      36246: inst = 32'd136314880;
      36247: inst = 32'd268468224;
      36248: inst = 32'd201344048;
      36249: inst = 32'd203423744;
      36250: inst = 32'd471859200;
      36251: inst = 32'd136314880;
      36252: inst = 32'd268468224;
      36253: inst = 32'd201344049;
      36254: inst = 32'd203423744;
      36255: inst = 32'd471859200;
      36256: inst = 32'd136314880;
      36257: inst = 32'd268468224;
      36258: inst = 32'd201344050;
      36259: inst = 32'd203423744;
      36260: inst = 32'd471859200;
      36261: inst = 32'd136314880;
      36262: inst = 32'd268468224;
      36263: inst = 32'd201344051;
      36264: inst = 32'd203423744;
      36265: inst = 32'd471859200;
      36266: inst = 32'd136314880;
      36267: inst = 32'd268468224;
      36268: inst = 32'd201344052;
      36269: inst = 32'd203423744;
      36270: inst = 32'd471859200;
      36271: inst = 32'd136314880;
      36272: inst = 32'd268468224;
      36273: inst = 32'd201344053;
      36274: inst = 32'd203423744;
      36275: inst = 32'd471859200;
      36276: inst = 32'd136314880;
      36277: inst = 32'd268468224;
      36278: inst = 32'd201344054;
      36279: inst = 32'd203423744;
      36280: inst = 32'd471859200;
      36281: inst = 32'd136314880;
      36282: inst = 32'd268468224;
      36283: inst = 32'd201344055;
      36284: inst = 32'd203423744;
      36285: inst = 32'd471859200;
      36286: inst = 32'd136314880;
      36287: inst = 32'd268468224;
      36288: inst = 32'd201344056;
      36289: inst = 32'd203423744;
      36290: inst = 32'd471859200;
      36291: inst = 32'd136314880;
      36292: inst = 32'd268468224;
      36293: inst = 32'd201344057;
      36294: inst = 32'd203423744;
      36295: inst = 32'd471859200;
      36296: inst = 32'd136314880;
      36297: inst = 32'd268468224;
      36298: inst = 32'd201344058;
      36299: inst = 32'd203423744;
      36300: inst = 32'd471859200;
      36301: inst = 32'd136314880;
      36302: inst = 32'd268468224;
      36303: inst = 32'd201344059;
      36304: inst = 32'd203423744;
      36305: inst = 32'd471859200;
      36306: inst = 32'd136314880;
      36307: inst = 32'd268468224;
      36308: inst = 32'd201344060;
      36309: inst = 32'd203423744;
      36310: inst = 32'd471859200;
      36311: inst = 32'd136314880;
      36312: inst = 32'd268468224;
      36313: inst = 32'd201344061;
      36314: inst = 32'd203423744;
      36315: inst = 32'd471859200;
      36316: inst = 32'd136314880;
      36317: inst = 32'd268468224;
      36318: inst = 32'd201344062;
      36319: inst = 32'd203423744;
      36320: inst = 32'd471859200;
      36321: inst = 32'd136314880;
      36322: inst = 32'd268468224;
      36323: inst = 32'd201344063;
      36324: inst = 32'd203423744;
      36325: inst = 32'd471859200;
      36326: inst = 32'd136314880;
      36327: inst = 32'd268468224;
      36328: inst = 32'd201344064;
      36329: inst = 32'd203423744;
      36330: inst = 32'd471859200;
      36331: inst = 32'd136314880;
      36332: inst = 32'd268468224;
      36333: inst = 32'd201344065;
      36334: inst = 32'd203423744;
      36335: inst = 32'd471859200;
      36336: inst = 32'd136314880;
      36337: inst = 32'd268468224;
      36338: inst = 32'd201344066;
      36339: inst = 32'd203423744;
      36340: inst = 32'd471859200;
      36341: inst = 32'd136314880;
      36342: inst = 32'd268468224;
      36343: inst = 32'd201344067;
      36344: inst = 32'd203423744;
      36345: inst = 32'd471859200;
      36346: inst = 32'd136314880;
      36347: inst = 32'd268468224;
      36348: inst = 32'd201344068;
      36349: inst = 32'd203423744;
      36350: inst = 32'd471859200;
      36351: inst = 32'd136314880;
      36352: inst = 32'd268468224;
      36353: inst = 32'd201344069;
      36354: inst = 32'd203423744;
      36355: inst = 32'd471859200;
      36356: inst = 32'd136314880;
      36357: inst = 32'd268468224;
      36358: inst = 32'd201344070;
      36359: inst = 32'd203423744;
      36360: inst = 32'd471859200;
      36361: inst = 32'd136314880;
      36362: inst = 32'd268468224;
      36363: inst = 32'd201344071;
      36364: inst = 32'd203423744;
      36365: inst = 32'd471859200;
      36366: inst = 32'd136314880;
      36367: inst = 32'd268468224;
      36368: inst = 32'd201344072;
      36369: inst = 32'd203423744;
      36370: inst = 32'd471859200;
      36371: inst = 32'd136314880;
      36372: inst = 32'd268468224;
      36373: inst = 32'd201344073;
      36374: inst = 32'd203423744;
      36375: inst = 32'd471859200;
      36376: inst = 32'd136314880;
      36377: inst = 32'd268468224;
      36378: inst = 32'd201344074;
      36379: inst = 32'd203423744;
      36380: inst = 32'd471859200;
      36381: inst = 32'd136314880;
      36382: inst = 32'd268468224;
      36383: inst = 32'd201344075;
      36384: inst = 32'd203423744;
      36385: inst = 32'd471859200;
      36386: inst = 32'd136314880;
      36387: inst = 32'd268468224;
      36388: inst = 32'd201344076;
      36389: inst = 32'd203423744;
      36390: inst = 32'd471859200;
      36391: inst = 32'd136314880;
      36392: inst = 32'd268468224;
      36393: inst = 32'd201344077;
      36394: inst = 32'd203423744;
      36395: inst = 32'd471859200;
      36396: inst = 32'd136314880;
      36397: inst = 32'd268468224;
      36398: inst = 32'd201344078;
      36399: inst = 32'd203423744;
      36400: inst = 32'd471859200;
      36401: inst = 32'd136314880;
      36402: inst = 32'd268468224;
      36403: inst = 32'd201344079;
      36404: inst = 32'd203423744;
      36405: inst = 32'd471859200;
      36406: inst = 32'd136314880;
      36407: inst = 32'd268468224;
      36408: inst = 32'd201344080;
      36409: inst = 32'd203423744;
      36410: inst = 32'd471859200;
      36411: inst = 32'd136314880;
      36412: inst = 32'd268468224;
      36413: inst = 32'd201344081;
      36414: inst = 32'd203423744;
      36415: inst = 32'd471859200;
      36416: inst = 32'd136314880;
      36417: inst = 32'd268468224;
      36418: inst = 32'd201344082;
      36419: inst = 32'd203423744;
      36420: inst = 32'd471859200;
      36421: inst = 32'd136314880;
      36422: inst = 32'd268468224;
      36423: inst = 32'd201344083;
      36424: inst = 32'd203423744;
      36425: inst = 32'd471859200;
      36426: inst = 32'd136314880;
      36427: inst = 32'd268468224;
      36428: inst = 32'd201344084;
      36429: inst = 32'd203423744;
      36430: inst = 32'd471859200;
      36431: inst = 32'd136314880;
      36432: inst = 32'd268468224;
      36433: inst = 32'd201344085;
      36434: inst = 32'd203423744;
      36435: inst = 32'd471859200;
      36436: inst = 32'd136314880;
      36437: inst = 32'd268468224;
      36438: inst = 32'd201344086;
      36439: inst = 32'd203423744;
      36440: inst = 32'd471859200;
      36441: inst = 32'd136314880;
      36442: inst = 32'd268468224;
      36443: inst = 32'd201344087;
      36444: inst = 32'd203423744;
      36445: inst = 32'd471859200;
      36446: inst = 32'd136314880;
      36447: inst = 32'd268468224;
      36448: inst = 32'd201344088;
      36449: inst = 32'd203423744;
      36450: inst = 32'd471859200;
      36451: inst = 32'd136314880;
      36452: inst = 32'd268468224;
      36453: inst = 32'd201344089;
      36454: inst = 32'd203423744;
      36455: inst = 32'd471859200;
      36456: inst = 32'd136314880;
      36457: inst = 32'd268468224;
      36458: inst = 32'd201344090;
      36459: inst = 32'd203423744;
      36460: inst = 32'd471859200;
      36461: inst = 32'd136314880;
      36462: inst = 32'd268468224;
      36463: inst = 32'd201344091;
      36464: inst = 32'd203423744;
      36465: inst = 32'd471859200;
      36466: inst = 32'd136314880;
      36467: inst = 32'd268468224;
      36468: inst = 32'd201344092;
      36469: inst = 32'd203423744;
      36470: inst = 32'd471859200;
      36471: inst = 32'd136314880;
      36472: inst = 32'd268468224;
      36473: inst = 32'd201344093;
      36474: inst = 32'd203423744;
      36475: inst = 32'd471859200;
      36476: inst = 32'd136314880;
      36477: inst = 32'd268468224;
      36478: inst = 32'd201344094;
      36479: inst = 32'd203423744;
      36480: inst = 32'd471859200;
      36481: inst = 32'd136314880;
      36482: inst = 32'd268468224;
      36483: inst = 32'd201344095;
      36484: inst = 32'd203423744;
      36485: inst = 32'd471859200;
      36486: inst = 32'd136314880;
      36487: inst = 32'd268468224;
      36488: inst = 32'd201344096;
      36489: inst = 32'd203423744;
      36490: inst = 32'd471859200;
      36491: inst = 32'd136314880;
      36492: inst = 32'd268468224;
      36493: inst = 32'd201344097;
      36494: inst = 32'd203423744;
      36495: inst = 32'd471859200;
      36496: inst = 32'd136314880;
      36497: inst = 32'd268468224;
      36498: inst = 32'd201344098;
      36499: inst = 32'd203423744;
      36500: inst = 32'd471859200;
      36501: inst = 32'd136314880;
      36502: inst = 32'd268468224;
      36503: inst = 32'd201344099;
      36504: inst = 32'd203423744;
      36505: inst = 32'd471859200;
      36506: inst = 32'd136314880;
      36507: inst = 32'd268468224;
      36508: inst = 32'd201344100;
      36509: inst = 32'd203423744;
      36510: inst = 32'd471859200;
      36511: inst = 32'd136314880;
      36512: inst = 32'd268468224;
      36513: inst = 32'd201344101;
      36514: inst = 32'd203423744;
      36515: inst = 32'd471859200;
      36516: inst = 32'd136314880;
      36517: inst = 32'd268468224;
      36518: inst = 32'd201344102;
      36519: inst = 32'd203423744;
      36520: inst = 32'd471859200;
      36521: inst = 32'd136314880;
      36522: inst = 32'd268468224;
      36523: inst = 32'd201344103;
      36524: inst = 32'd203423744;
      36525: inst = 32'd471859200;
      36526: inst = 32'd136314880;
      36527: inst = 32'd268468224;
      36528: inst = 32'd201344104;
      36529: inst = 32'd203423744;
      36530: inst = 32'd471859200;
      36531: inst = 32'd136314880;
      36532: inst = 32'd268468224;
      36533: inst = 32'd201344105;
      36534: inst = 32'd203423744;
      36535: inst = 32'd471859200;
      36536: inst = 32'd136314880;
      36537: inst = 32'd268468224;
      36538: inst = 32'd201344106;
      36539: inst = 32'd203423744;
      36540: inst = 32'd471859200;
      36541: inst = 32'd136314880;
      36542: inst = 32'd268468224;
      36543: inst = 32'd201344107;
      36544: inst = 32'd203423744;
      36545: inst = 32'd471859200;
      36546: inst = 32'd136314880;
      36547: inst = 32'd268468224;
      36548: inst = 32'd201344108;
      36549: inst = 32'd203423744;
      36550: inst = 32'd471859200;
      36551: inst = 32'd136314880;
      36552: inst = 32'd268468224;
      36553: inst = 32'd201344109;
      36554: inst = 32'd203423744;
      36555: inst = 32'd471859200;
      36556: inst = 32'd136314880;
      36557: inst = 32'd268468224;
      36558: inst = 32'd201344110;
      36559: inst = 32'd203483685;
      36560: inst = 32'd471859200;
      36561: inst = 32'd136314880;
      36562: inst = 32'd268468224;
      36563: inst = 32'd201344111;
      36564: inst = 32'd203483685;
      36565: inst = 32'd471859200;
      36566: inst = 32'd136314880;
      36567: inst = 32'd268468224;
      36568: inst = 32'd201344112;
      36569: inst = 32'd203483685;
      36570: inst = 32'd471859200;
      36571: inst = 32'd136314880;
      36572: inst = 32'd268468224;
      36573: inst = 32'd201344113;
      36574: inst = 32'd203483685;
      36575: inst = 32'd471859200;
      36576: inst = 32'd136314880;
      36577: inst = 32'd268468224;
      36578: inst = 32'd201344114;
      36579: inst = 32'd203483685;
      36580: inst = 32'd471859200;
      36581: inst = 32'd136314880;
      36582: inst = 32'd268468224;
      36583: inst = 32'd201344115;
      36584: inst = 32'd203483685;
      36585: inst = 32'd471859200;
      36586: inst = 32'd136314880;
      36587: inst = 32'd268468224;
      36588: inst = 32'd201344116;
      36589: inst = 32'd203483685;
      36590: inst = 32'd471859200;
      36591: inst = 32'd136314880;
      36592: inst = 32'd268468224;
      36593: inst = 32'd201344117;
      36594: inst = 32'd203483685;
      36595: inst = 32'd471859200;
      36596: inst = 32'd136314880;
      36597: inst = 32'd268468224;
      36598: inst = 32'd201344118;
      36599: inst = 32'd203483685;
      36600: inst = 32'd471859200;
      36601: inst = 32'd136314880;
      36602: inst = 32'd268468224;
      36603: inst = 32'd201344119;
      36604: inst = 32'd203483685;
      36605: inst = 32'd471859200;
      36606: inst = 32'd136314880;
      36607: inst = 32'd268468224;
      36608: inst = 32'd201344120;
      36609: inst = 32'd203483685;
      36610: inst = 32'd471859200;
      36611: inst = 32'd136314880;
      36612: inst = 32'd268468224;
      36613: inst = 32'd201344121;
      36614: inst = 32'd203423744;
      36615: inst = 32'd471859200;
      36616: inst = 32'd136314880;
      36617: inst = 32'd268468224;
      36618: inst = 32'd201344122;
      36619: inst = 32'd203483685;
      36620: inst = 32'd471859200;
      36621: inst = 32'd136314880;
      36622: inst = 32'd268468224;
      36623: inst = 32'd201344123;
      36624: inst = 32'd203483685;
      36625: inst = 32'd471859200;
      36626: inst = 32'd136314880;
      36627: inst = 32'd268468224;
      36628: inst = 32'd201344124;
      36629: inst = 32'd203483685;
      36630: inst = 32'd471859200;
      36631: inst = 32'd136314880;
      36632: inst = 32'd268468224;
      36633: inst = 32'd201344125;
      36634: inst = 32'd203483685;
      36635: inst = 32'd471859200;
      36636: inst = 32'd136314880;
      36637: inst = 32'd268468224;
      36638: inst = 32'd201344126;
      36639: inst = 32'd203483685;
      36640: inst = 32'd471859200;
      36641: inst = 32'd136314880;
      36642: inst = 32'd268468224;
      36643: inst = 32'd201344127;
      36644: inst = 32'd203483685;
      36645: inst = 32'd471859200;
      36646: inst = 32'd136314880;
      36647: inst = 32'd268468224;
      36648: inst = 32'd201344128;
      36649: inst = 32'd203483685;
      36650: inst = 32'd471859200;
      36651: inst = 32'd136314880;
      36652: inst = 32'd268468224;
      36653: inst = 32'd201344129;
      36654: inst = 32'd203483685;
      36655: inst = 32'd471859200;
      36656: inst = 32'd136314880;
      36657: inst = 32'd268468224;
      36658: inst = 32'd201344130;
      36659: inst = 32'd203483685;
      36660: inst = 32'd471859200;
      36661: inst = 32'd136314880;
      36662: inst = 32'd268468224;
      36663: inst = 32'd201344131;
      36664: inst = 32'd203483685;
      36665: inst = 32'd471859200;
      36666: inst = 32'd136314880;
      36667: inst = 32'd268468224;
      36668: inst = 32'd201344132;
      36669: inst = 32'd203483685;
      36670: inst = 32'd471859200;
      36671: inst = 32'd136314880;
      36672: inst = 32'd268468224;
      36673: inst = 32'd201344133;
      36674: inst = 32'd203483685;
      36675: inst = 32'd471859200;
      36676: inst = 32'd136314880;
      36677: inst = 32'd268468224;
      36678: inst = 32'd201344134;
      36679: inst = 32'd203483685;
      36680: inst = 32'd471859200;
      36681: inst = 32'd136314880;
      36682: inst = 32'd268468224;
      36683: inst = 32'd201344135;
      36684: inst = 32'd203483685;
      36685: inst = 32'd471859200;
      36686: inst = 32'd136314880;
      36687: inst = 32'd268468224;
      36688: inst = 32'd201344136;
      36689: inst = 32'd203483685;
      36690: inst = 32'd471859200;
      36691: inst = 32'd136314880;
      36692: inst = 32'd268468224;
      36693: inst = 32'd201344137;
      36694: inst = 32'd203483685;
      36695: inst = 32'd471859200;
      36696: inst = 32'd136314880;
      36697: inst = 32'd268468224;
      36698: inst = 32'd201344138;
      36699: inst = 32'd203483685;
      36700: inst = 32'd471859200;
      36701: inst = 32'd136314880;
      36702: inst = 32'd268468224;
      36703: inst = 32'd201344139;
      36704: inst = 32'd203483685;
      36705: inst = 32'd471859200;
      36706: inst = 32'd136314880;
      36707: inst = 32'd268468224;
      36708: inst = 32'd201344140;
      36709: inst = 32'd203483685;
      36710: inst = 32'd471859200;
      36711: inst = 32'd136314880;
      36712: inst = 32'd268468224;
      36713: inst = 32'd201344141;
      36714: inst = 32'd203483685;
      36715: inst = 32'd471859200;
      36716: inst = 32'd136314880;
      36717: inst = 32'd268468224;
      36718: inst = 32'd201344142;
      36719: inst = 32'd203483685;
      36720: inst = 32'd471859200;
      36721: inst = 32'd136314880;
      36722: inst = 32'd268468224;
      36723: inst = 32'd201344143;
      36724: inst = 32'd203423744;
      36725: inst = 32'd471859200;
      36726: inst = 32'd136314880;
      36727: inst = 32'd268468224;
      36728: inst = 32'd201344144;
      36729: inst = 32'd203423744;
      36730: inst = 32'd471859200;
      36731: inst = 32'd136314880;
      36732: inst = 32'd268468224;
      36733: inst = 32'd201344145;
      36734: inst = 32'd203423744;
      36735: inst = 32'd471859200;
      36736: inst = 32'd136314880;
      36737: inst = 32'd268468224;
      36738: inst = 32'd201344146;
      36739: inst = 32'd203483685;
      36740: inst = 32'd471859200;
      36741: inst = 32'd136314880;
      36742: inst = 32'd268468224;
      36743: inst = 32'd201344147;
      36744: inst = 32'd203483685;
      36745: inst = 32'd471859200;
      36746: inst = 32'd136314880;
      36747: inst = 32'd268468224;
      36748: inst = 32'd201344148;
      36749: inst = 32'd203483685;
      36750: inst = 32'd471859200;
      36751: inst = 32'd136314880;
      36752: inst = 32'd268468224;
      36753: inst = 32'd201344149;
      36754: inst = 32'd203483685;
      36755: inst = 32'd471859200;
      36756: inst = 32'd136314880;
      36757: inst = 32'd268468224;
      36758: inst = 32'd201344150;
      36759: inst = 32'd203483685;
      36760: inst = 32'd471859200;
      36761: inst = 32'd136314880;
      36762: inst = 32'd268468224;
      36763: inst = 32'd201344151;
      36764: inst = 32'd203483685;
      36765: inst = 32'd471859200;
      36766: inst = 32'd136314880;
      36767: inst = 32'd268468224;
      36768: inst = 32'd201344152;
      36769: inst = 32'd203483685;
      36770: inst = 32'd471859200;
      36771: inst = 32'd136314880;
      36772: inst = 32'd268468224;
      36773: inst = 32'd201344153;
      36774: inst = 32'd203483685;
      36775: inst = 32'd471859200;
      36776: inst = 32'd136314880;
      36777: inst = 32'd268468224;
      36778: inst = 32'd201344154;
      36779: inst = 32'd203483685;
      36780: inst = 32'd471859200;
      36781: inst = 32'd136314880;
      36782: inst = 32'd268468224;
      36783: inst = 32'd201344155;
      36784: inst = 32'd203483685;
      36785: inst = 32'd471859200;
      36786: inst = 32'd136314880;
      36787: inst = 32'd268468224;
      36788: inst = 32'd201344156;
      36789: inst = 32'd203483685;
      36790: inst = 32'd471859200;
      36791: inst = 32'd136314880;
      36792: inst = 32'd268468224;
      36793: inst = 32'd201344157;
      36794: inst = 32'd203483685;
      36795: inst = 32'd471859200;
      36796: inst = 32'd136314880;
      36797: inst = 32'd268468224;
      36798: inst = 32'd201344158;
      36799: inst = 32'd203483685;
      36800: inst = 32'd471859200;
      36801: inst = 32'd136314880;
      36802: inst = 32'd268468224;
      36803: inst = 32'd201344159;
      36804: inst = 32'd203483685;
      36805: inst = 32'd471859200;
      36806: inst = 32'd136314880;
      36807: inst = 32'd268468224;
      36808: inst = 32'd201344160;
      36809: inst = 32'd203483685;
      36810: inst = 32'd471859200;
      36811: inst = 32'd136314880;
      36812: inst = 32'd268468224;
      36813: inst = 32'd201344161;
      36814: inst = 32'd203483685;
      36815: inst = 32'd471859200;
      36816: inst = 32'd136314880;
      36817: inst = 32'd268468224;
      36818: inst = 32'd201344162;
      36819: inst = 32'd203483685;
      36820: inst = 32'd471859200;
      36821: inst = 32'd136314880;
      36822: inst = 32'd268468224;
      36823: inst = 32'd201344163;
      36824: inst = 32'd203483685;
      36825: inst = 32'd471859200;
      36826: inst = 32'd136314880;
      36827: inst = 32'd268468224;
      36828: inst = 32'd201344164;
      36829: inst = 32'd203483685;
      36830: inst = 32'd471859200;
      36831: inst = 32'd136314880;
      36832: inst = 32'd268468224;
      36833: inst = 32'd201344165;
      36834: inst = 32'd203483685;
      36835: inst = 32'd471859200;
      36836: inst = 32'd136314880;
      36837: inst = 32'd268468224;
      36838: inst = 32'd201344166;
      36839: inst = 32'd203483685;
      36840: inst = 32'd471859200;
      36841: inst = 32'd136314880;
      36842: inst = 32'd268468224;
      36843: inst = 32'd201344167;
      36844: inst = 32'd203483685;
      36845: inst = 32'd471859200;
      36846: inst = 32'd136314880;
      36847: inst = 32'd268468224;
      36848: inst = 32'd201344168;
      36849: inst = 32'd203483685;
      36850: inst = 32'd471859200;
      36851: inst = 32'd136314880;
      36852: inst = 32'd268468224;
      36853: inst = 32'd201344169;
      36854: inst = 32'd203423744;
      36855: inst = 32'd471859200;
      36856: inst = 32'd136314880;
      36857: inst = 32'd268468224;
      36858: inst = 32'd201344170;
      36859: inst = 32'd203423744;
      36860: inst = 32'd471859200;
      36861: inst = 32'd136314880;
      36862: inst = 32'd268468224;
      36863: inst = 32'd201344171;
      36864: inst = 32'd203423744;
      36865: inst = 32'd471859200;
      36866: inst = 32'd136314880;
      36867: inst = 32'd268468224;
      36868: inst = 32'd201344172;
      36869: inst = 32'd203483685;
      36870: inst = 32'd471859200;
      36871: inst = 32'd136314880;
      36872: inst = 32'd268468224;
      36873: inst = 32'd201344173;
      36874: inst = 32'd203483685;
      36875: inst = 32'd471859200;
      36876: inst = 32'd136314880;
      36877: inst = 32'd268468224;
      36878: inst = 32'd201344174;
      36879: inst = 32'd203483685;
      36880: inst = 32'd471859200;
      36881: inst = 32'd136314880;
      36882: inst = 32'd268468224;
      36883: inst = 32'd201344175;
      36884: inst = 32'd203483685;
      36885: inst = 32'd471859200;
      36886: inst = 32'd136314880;
      36887: inst = 32'd268468224;
      36888: inst = 32'd201344176;
      36889: inst = 32'd203483685;
      36890: inst = 32'd471859200;
      36891: inst = 32'd136314880;
      36892: inst = 32'd268468224;
      36893: inst = 32'd201344177;
      36894: inst = 32'd203483685;
      36895: inst = 32'd471859200;
      36896: inst = 32'd136314880;
      36897: inst = 32'd268468224;
      36898: inst = 32'd201344178;
      36899: inst = 32'd203483685;
      36900: inst = 32'd471859200;
      36901: inst = 32'd136314880;
      36902: inst = 32'd268468224;
      36903: inst = 32'd201344179;
      36904: inst = 32'd203483685;
      36905: inst = 32'd471859200;
      36906: inst = 32'd136314880;
      36907: inst = 32'd268468224;
      36908: inst = 32'd201344180;
      36909: inst = 32'd203483685;
      36910: inst = 32'd471859200;
      36911: inst = 32'd136314880;
      36912: inst = 32'd268468224;
      36913: inst = 32'd201344181;
      36914: inst = 32'd203483685;
      36915: inst = 32'd471859200;
      36916: inst = 32'd136314880;
      36917: inst = 32'd268468224;
      36918: inst = 32'd201344182;
      36919: inst = 32'd203423744;
      36920: inst = 32'd471859200;
      36921: inst = 32'd136314880;
      36922: inst = 32'd268468224;
      36923: inst = 32'd201344183;
      36924: inst = 32'd203423744;
      36925: inst = 32'd471859200;
      36926: inst = 32'd136314880;
      36927: inst = 32'd268468224;
      36928: inst = 32'd201344184;
      36929: inst = 32'd203423744;
      36930: inst = 32'd471859200;
      36931: inst = 32'd136314880;
      36932: inst = 32'd268468224;
      36933: inst = 32'd201344185;
      36934: inst = 32'd203423744;
      36935: inst = 32'd471859200;
      36936: inst = 32'd136314880;
      36937: inst = 32'd268468224;
      36938: inst = 32'd201344186;
      36939: inst = 32'd203423744;
      36940: inst = 32'd471859200;
      36941: inst = 32'd136314880;
      36942: inst = 32'd268468224;
      36943: inst = 32'd201344187;
      36944: inst = 32'd203423744;
      36945: inst = 32'd471859200;
      36946: inst = 32'd136314880;
      36947: inst = 32'd268468224;
      36948: inst = 32'd201344188;
      36949: inst = 32'd203423744;
      36950: inst = 32'd471859200;
      36951: inst = 32'd136314880;
      36952: inst = 32'd268468224;
      36953: inst = 32'd201344189;
      36954: inst = 32'd203423744;
      36955: inst = 32'd471859200;
      36956: inst = 32'd136314880;
      36957: inst = 32'd268468224;
      36958: inst = 32'd201344190;
      36959: inst = 32'd203423744;
      36960: inst = 32'd471859200;
      36961: inst = 32'd136314880;
      36962: inst = 32'd268468224;
      36963: inst = 32'd201344191;
      36964: inst = 32'd203423744;
      36965: inst = 32'd471859200;
      36966: inst = 32'd136314880;
      36967: inst = 32'd268468224;
      36968: inst = 32'd201344192;
      36969: inst = 32'd203423744;
      36970: inst = 32'd471859200;
      36971: inst = 32'd136314880;
      36972: inst = 32'd268468224;
      36973: inst = 32'd201344193;
      36974: inst = 32'd203423744;
      36975: inst = 32'd471859200;
      36976: inst = 32'd136314880;
      36977: inst = 32'd268468224;
      36978: inst = 32'd201344194;
      36979: inst = 32'd203423744;
      36980: inst = 32'd471859200;
      36981: inst = 32'd136314880;
      36982: inst = 32'd268468224;
      36983: inst = 32'd201344195;
      36984: inst = 32'd203423744;
      36985: inst = 32'd471859200;
      36986: inst = 32'd136314880;
      36987: inst = 32'd268468224;
      36988: inst = 32'd201344196;
      36989: inst = 32'd203423744;
      36990: inst = 32'd471859200;
      36991: inst = 32'd136314880;
      36992: inst = 32'd268468224;
      36993: inst = 32'd201344197;
      36994: inst = 32'd203423744;
      36995: inst = 32'd471859200;
      36996: inst = 32'd136314880;
      36997: inst = 32'd268468224;
      36998: inst = 32'd201344198;
      36999: inst = 32'd203423744;
      37000: inst = 32'd471859200;
      37001: inst = 32'd136314880;
      37002: inst = 32'd268468224;
      37003: inst = 32'd201344199;
      37004: inst = 32'd203423744;
      37005: inst = 32'd471859200;
      37006: inst = 32'd136314880;
      37007: inst = 32'd268468224;
      37008: inst = 32'd201344200;
      37009: inst = 32'd203423744;
      37010: inst = 32'd471859200;
      37011: inst = 32'd136314880;
      37012: inst = 32'd268468224;
      37013: inst = 32'd201344201;
      37014: inst = 32'd203423744;
      37015: inst = 32'd471859200;
      37016: inst = 32'd136314880;
      37017: inst = 32'd268468224;
      37018: inst = 32'd201344202;
      37019: inst = 32'd203423744;
      37020: inst = 32'd471859200;
      37021: inst = 32'd136314880;
      37022: inst = 32'd268468224;
      37023: inst = 32'd201344203;
      37024: inst = 32'd203423744;
      37025: inst = 32'd471859200;
      37026: inst = 32'd136314880;
      37027: inst = 32'd268468224;
      37028: inst = 32'd201344204;
      37029: inst = 32'd203423744;
      37030: inst = 32'd471859200;
      37031: inst = 32'd136314880;
      37032: inst = 32'd268468224;
      37033: inst = 32'd201344205;
      37034: inst = 32'd203483685;
      37035: inst = 32'd471859200;
      37036: inst = 32'd136314880;
      37037: inst = 32'd268468224;
      37038: inst = 32'd201344206;
      37039: inst = 32'd203483685;
      37040: inst = 32'd471859200;
      37041: inst = 32'd136314880;
      37042: inst = 32'd268468224;
      37043: inst = 32'd201344207;
      37044: inst = 32'd203483685;
      37045: inst = 32'd471859200;
      37046: inst = 32'd136314880;
      37047: inst = 32'd268468224;
      37048: inst = 32'd201344208;
      37049: inst = 32'd203483685;
      37050: inst = 32'd471859200;
      37051: inst = 32'd136314880;
      37052: inst = 32'd268468224;
      37053: inst = 32'd201344209;
      37054: inst = 32'd203483685;
      37055: inst = 32'd471859200;
      37056: inst = 32'd136314880;
      37057: inst = 32'd268468224;
      37058: inst = 32'd201344210;
      37059: inst = 32'd203483685;
      37060: inst = 32'd471859200;
      37061: inst = 32'd136314880;
      37062: inst = 32'd268468224;
      37063: inst = 32'd201344211;
      37064: inst = 32'd203483685;
      37065: inst = 32'd471859200;
      37066: inst = 32'd136314880;
      37067: inst = 32'd268468224;
      37068: inst = 32'd201344212;
      37069: inst = 32'd203483685;
      37070: inst = 32'd471859200;
      37071: inst = 32'd136314880;
      37072: inst = 32'd268468224;
      37073: inst = 32'd201344213;
      37074: inst = 32'd203483685;
      37075: inst = 32'd471859200;
      37076: inst = 32'd136314880;
      37077: inst = 32'd268468224;
      37078: inst = 32'd201344214;
      37079: inst = 32'd203483685;
      37080: inst = 32'd471859200;
      37081: inst = 32'd136314880;
      37082: inst = 32'd268468224;
      37083: inst = 32'd201344215;
      37084: inst = 32'd203483685;
      37085: inst = 32'd471859200;
      37086: inst = 32'd136314880;
      37087: inst = 32'd268468224;
      37088: inst = 32'd201344216;
      37089: inst = 32'd203483685;
      37090: inst = 32'd471859200;
      37091: inst = 32'd136314880;
      37092: inst = 32'd268468224;
      37093: inst = 32'd201344217;
      37094: inst = 32'd203483685;
      37095: inst = 32'd471859200;
      37096: inst = 32'd136314880;
      37097: inst = 32'd268468224;
      37098: inst = 32'd201344218;
      37099: inst = 32'd203483685;
      37100: inst = 32'd471859200;
      37101: inst = 32'd136314880;
      37102: inst = 32'd268468224;
      37103: inst = 32'd201344219;
      37104: inst = 32'd203483685;
      37105: inst = 32'd471859200;
      37106: inst = 32'd136314880;
      37107: inst = 32'd268468224;
      37108: inst = 32'd201344220;
      37109: inst = 32'd203483685;
      37110: inst = 32'd471859200;
      37111: inst = 32'd136314880;
      37112: inst = 32'd268468224;
      37113: inst = 32'd201344221;
      37114: inst = 32'd203483685;
      37115: inst = 32'd471859200;
      37116: inst = 32'd136314880;
      37117: inst = 32'd268468224;
      37118: inst = 32'd201344222;
      37119: inst = 32'd203483685;
      37120: inst = 32'd471859200;
      37121: inst = 32'd136314880;
      37122: inst = 32'd268468224;
      37123: inst = 32'd201344223;
      37124: inst = 32'd203483685;
      37125: inst = 32'd471859200;
      37126: inst = 32'd136314880;
      37127: inst = 32'd268468224;
      37128: inst = 32'd201344224;
      37129: inst = 32'd203483685;
      37130: inst = 32'd471859200;
      37131: inst = 32'd136314880;
      37132: inst = 32'd268468224;
      37133: inst = 32'd201344225;
      37134: inst = 32'd203483685;
      37135: inst = 32'd471859200;
      37136: inst = 32'd136314880;
      37137: inst = 32'd268468224;
      37138: inst = 32'd201344226;
      37139: inst = 32'd203483685;
      37140: inst = 32'd471859200;
      37141: inst = 32'd136314880;
      37142: inst = 32'd268468224;
      37143: inst = 32'd201344227;
      37144: inst = 32'd203483685;
      37145: inst = 32'd471859200;
      37146: inst = 32'd136314880;
      37147: inst = 32'd268468224;
      37148: inst = 32'd201344228;
      37149: inst = 32'd203483685;
      37150: inst = 32'd471859200;
      37151: inst = 32'd136314880;
      37152: inst = 32'd268468224;
      37153: inst = 32'd201344229;
      37154: inst = 32'd203483685;
      37155: inst = 32'd471859200;
      37156: inst = 32'd136314880;
      37157: inst = 32'd268468224;
      37158: inst = 32'd201344230;
      37159: inst = 32'd203483685;
      37160: inst = 32'd471859200;
      37161: inst = 32'd136314880;
      37162: inst = 32'd268468224;
      37163: inst = 32'd201344231;
      37164: inst = 32'd203483685;
      37165: inst = 32'd471859200;
      37166: inst = 32'd136314880;
      37167: inst = 32'd268468224;
      37168: inst = 32'd201344232;
      37169: inst = 32'd203483685;
      37170: inst = 32'd471859200;
      37171: inst = 32'd136314880;
      37172: inst = 32'd268468224;
      37173: inst = 32'd201344233;
      37174: inst = 32'd203483685;
      37175: inst = 32'd471859200;
      37176: inst = 32'd136314880;
      37177: inst = 32'd268468224;
      37178: inst = 32'd201344234;
      37179: inst = 32'd203483685;
      37180: inst = 32'd471859200;
      37181: inst = 32'd136314880;
      37182: inst = 32'd268468224;
      37183: inst = 32'd201344235;
      37184: inst = 32'd203483685;
      37185: inst = 32'd471859200;
      37186: inst = 32'd136314880;
      37187: inst = 32'd268468224;
      37188: inst = 32'd201344236;
      37189: inst = 32'd203483685;
      37190: inst = 32'd471859200;
      37191: inst = 32'd136314880;
      37192: inst = 32'd268468224;
      37193: inst = 32'd201344237;
      37194: inst = 32'd203483685;
      37195: inst = 32'd471859200;
      37196: inst = 32'd136314880;
      37197: inst = 32'd268468224;
      37198: inst = 32'd201344238;
      37199: inst = 32'd203483685;
      37200: inst = 32'd471859200;
      37201: inst = 32'd136314880;
      37202: inst = 32'd268468224;
      37203: inst = 32'd201344239;
      37204: inst = 32'd203423744;
      37205: inst = 32'd471859200;
      37206: inst = 32'd136314880;
      37207: inst = 32'd268468224;
      37208: inst = 32'd201344240;
      37209: inst = 32'd203423744;
      37210: inst = 32'd471859200;
      37211: inst = 32'd136314880;
      37212: inst = 32'd268468224;
      37213: inst = 32'd201344241;
      37214: inst = 32'd203483685;
      37215: inst = 32'd471859200;
      37216: inst = 32'd136314880;
      37217: inst = 32'd268468224;
      37218: inst = 32'd201344242;
      37219: inst = 32'd203483685;
      37220: inst = 32'd471859200;
      37221: inst = 32'd136314880;
      37222: inst = 32'd268468224;
      37223: inst = 32'd201344243;
      37224: inst = 32'd203483685;
      37225: inst = 32'd471859200;
      37226: inst = 32'd136314880;
      37227: inst = 32'd268468224;
      37228: inst = 32'd201344244;
      37229: inst = 32'd203483685;
      37230: inst = 32'd471859200;
      37231: inst = 32'd136314880;
      37232: inst = 32'd268468224;
      37233: inst = 32'd201344245;
      37234: inst = 32'd203483685;
      37235: inst = 32'd471859200;
      37236: inst = 32'd136314880;
      37237: inst = 32'd268468224;
      37238: inst = 32'd201344246;
      37239: inst = 32'd203483685;
      37240: inst = 32'd471859200;
      37241: inst = 32'd136314880;
      37242: inst = 32'd268468224;
      37243: inst = 32'd201344247;
      37244: inst = 32'd203483685;
      37245: inst = 32'd471859200;
      37246: inst = 32'd136314880;
      37247: inst = 32'd268468224;
      37248: inst = 32'd201344248;
      37249: inst = 32'd203483685;
      37250: inst = 32'd471859200;
      37251: inst = 32'd136314880;
      37252: inst = 32'd268468224;
      37253: inst = 32'd201344249;
      37254: inst = 32'd203483685;
      37255: inst = 32'd471859200;
      37256: inst = 32'd136314880;
      37257: inst = 32'd268468224;
      37258: inst = 32'd201344250;
      37259: inst = 32'd203483685;
      37260: inst = 32'd471859200;
      37261: inst = 32'd136314880;
      37262: inst = 32'd268468224;
      37263: inst = 32'd201344251;
      37264: inst = 32'd203483685;
      37265: inst = 32'd471859200;
      37266: inst = 32'd136314880;
      37267: inst = 32'd268468224;
      37268: inst = 32'd201344252;
      37269: inst = 32'd203483685;
      37270: inst = 32'd471859200;
      37271: inst = 32'd136314880;
      37272: inst = 32'd268468224;
      37273: inst = 32'd201344253;
      37274: inst = 32'd203483685;
      37275: inst = 32'd471859200;
      37276: inst = 32'd136314880;
      37277: inst = 32'd268468224;
      37278: inst = 32'd201344254;
      37279: inst = 32'd203483685;
      37280: inst = 32'd471859200;
      37281: inst = 32'd136314880;
      37282: inst = 32'd268468224;
      37283: inst = 32'd201344255;
      37284: inst = 32'd203483685;
      37285: inst = 32'd471859200;
      37286: inst = 32'd136314880;
      37287: inst = 32'd268468224;
      37288: inst = 32'd201344256;
      37289: inst = 32'd203483685;
      37290: inst = 32'd471859200;
      37291: inst = 32'd136314880;
      37292: inst = 32'd268468224;
      37293: inst = 32'd201344257;
      37294: inst = 32'd203483685;
      37295: inst = 32'd471859200;
      37296: inst = 32'd136314880;
      37297: inst = 32'd268468224;
      37298: inst = 32'd201344258;
      37299: inst = 32'd203483685;
      37300: inst = 32'd471859200;
      37301: inst = 32'd136314880;
      37302: inst = 32'd268468224;
      37303: inst = 32'd201344259;
      37304: inst = 32'd203483685;
      37305: inst = 32'd471859200;
      37306: inst = 32'd136314880;
      37307: inst = 32'd268468224;
      37308: inst = 32'd201344260;
      37309: inst = 32'd203483685;
      37310: inst = 32'd471859200;
      37311: inst = 32'd136314880;
      37312: inst = 32'd268468224;
      37313: inst = 32'd201344261;
      37314: inst = 32'd203483685;
      37315: inst = 32'd471859200;
      37316: inst = 32'd136314880;
      37317: inst = 32'd268468224;
      37318: inst = 32'd201344262;
      37319: inst = 32'd203483685;
      37320: inst = 32'd471859200;
      37321: inst = 32'd136314880;
      37322: inst = 32'd268468224;
      37323: inst = 32'd201344263;
      37324: inst = 32'd203483685;
      37325: inst = 32'd471859200;
      37326: inst = 32'd136314880;
      37327: inst = 32'd268468224;
      37328: inst = 32'd201344264;
      37329: inst = 32'd203483685;
      37330: inst = 32'd471859200;
      37331: inst = 32'd136314880;
      37332: inst = 32'd268468224;
      37333: inst = 32'd201344265;
      37334: inst = 32'd203423744;
      37335: inst = 32'd471859200;
      37336: inst = 32'd136314880;
      37337: inst = 32'd268468224;
      37338: inst = 32'd201344266;
      37339: inst = 32'd203423744;
      37340: inst = 32'd471859200;
      37341: inst = 32'd136314880;
      37342: inst = 32'd268468224;
      37343: inst = 32'd201344267;
      37344: inst = 32'd203483685;
      37345: inst = 32'd471859200;
      37346: inst = 32'd136314880;
      37347: inst = 32'd268468224;
      37348: inst = 32'd201344268;
      37349: inst = 32'd203483685;
      37350: inst = 32'd471859200;
      37351: inst = 32'd136314880;
      37352: inst = 32'd268468224;
      37353: inst = 32'd201344269;
      37354: inst = 32'd203483685;
      37355: inst = 32'd471859200;
      37356: inst = 32'd136314880;
      37357: inst = 32'd268468224;
      37358: inst = 32'd201344270;
      37359: inst = 32'd203483685;
      37360: inst = 32'd471859200;
      37361: inst = 32'd136314880;
      37362: inst = 32'd268468224;
      37363: inst = 32'd201344271;
      37364: inst = 32'd203483685;
      37365: inst = 32'd471859200;
      37366: inst = 32'd136314880;
      37367: inst = 32'd268468224;
      37368: inst = 32'd201344272;
      37369: inst = 32'd203483685;
      37370: inst = 32'd471859200;
      37371: inst = 32'd136314880;
      37372: inst = 32'd268468224;
      37373: inst = 32'd201344273;
      37374: inst = 32'd203483685;
      37375: inst = 32'd471859200;
      37376: inst = 32'd136314880;
      37377: inst = 32'd268468224;
      37378: inst = 32'd201344274;
      37379: inst = 32'd203483685;
      37380: inst = 32'd471859200;
      37381: inst = 32'd136314880;
      37382: inst = 32'd268468224;
      37383: inst = 32'd201344275;
      37384: inst = 32'd203483685;
      37385: inst = 32'd471859200;
      37386: inst = 32'd136314880;
      37387: inst = 32'd268468224;
      37388: inst = 32'd201344276;
      37389: inst = 32'd203483685;
      37390: inst = 32'd471859200;
      37391: inst = 32'd136314880;
      37392: inst = 32'd268468224;
      37393: inst = 32'd201344277;
      37394: inst = 32'd203483685;
      37395: inst = 32'd471859200;
      37396: inst = 32'd136314880;
      37397: inst = 32'd268468224;
      37398: inst = 32'd201344278;
      37399: inst = 32'd203423744;
      37400: inst = 32'd471859200;
      37401: inst = 32'd136314880;
      37402: inst = 32'd268468224;
      37403: inst = 32'd201344279;
      37404: inst = 32'd203423744;
      37405: inst = 32'd471859200;
      37406: inst = 32'd136314880;
      37407: inst = 32'd268468224;
      37408: inst = 32'd201344280;
      37409: inst = 32'd203423744;
      37410: inst = 32'd471859200;
      37411: inst = 32'd136314880;
      37412: inst = 32'd268468224;
      37413: inst = 32'd201344281;
      37414: inst = 32'd203423744;
      37415: inst = 32'd471859200;
      37416: inst = 32'd136314880;
      37417: inst = 32'd268468224;
      37418: inst = 32'd201344282;
      37419: inst = 32'd203423744;
      37420: inst = 32'd471859200;
      37421: inst = 32'd136314880;
      37422: inst = 32'd268468224;
      37423: inst = 32'd201344283;
      37424: inst = 32'd203423744;
      37425: inst = 32'd471859200;
      37426: inst = 32'd136314880;
      37427: inst = 32'd268468224;
      37428: inst = 32'd201344284;
      37429: inst = 32'd203423744;
      37430: inst = 32'd471859200;
      37431: inst = 32'd136314880;
      37432: inst = 32'd268468224;
      37433: inst = 32'd201344285;
      37434: inst = 32'd203423744;
      37435: inst = 32'd471859200;
      37436: inst = 32'd136314880;
      37437: inst = 32'd268468224;
      37438: inst = 32'd201344286;
      37439: inst = 32'd203423744;
      37440: inst = 32'd471859200;
      37441: inst = 32'd136314880;
      37442: inst = 32'd268468224;
      37443: inst = 32'd201344287;
      37444: inst = 32'd203423744;
      37445: inst = 32'd471859200;
      37446: inst = 32'd136314880;
      37447: inst = 32'd268468224;
      37448: inst = 32'd201344288;
      37449: inst = 32'd203423744;
      37450: inst = 32'd471859200;
      37451: inst = 32'd136314880;
      37452: inst = 32'd268468224;
      37453: inst = 32'd201344289;
      37454: inst = 32'd203423744;
      37455: inst = 32'd471859200;
      37456: inst = 32'd136314880;
      37457: inst = 32'd268468224;
      37458: inst = 32'd201344290;
      37459: inst = 32'd203423744;
      37460: inst = 32'd471859200;
      37461: inst = 32'd136314880;
      37462: inst = 32'd268468224;
      37463: inst = 32'd201344291;
      37464: inst = 32'd203423744;
      37465: inst = 32'd471859200;
      37466: inst = 32'd136314880;
      37467: inst = 32'd268468224;
      37468: inst = 32'd201344292;
      37469: inst = 32'd203423744;
      37470: inst = 32'd471859200;
      37471: inst = 32'd136314880;
      37472: inst = 32'd268468224;
      37473: inst = 32'd201344293;
      37474: inst = 32'd203423744;
      37475: inst = 32'd471859200;
      37476: inst = 32'd136314880;
      37477: inst = 32'd268468224;
      37478: inst = 32'd201344294;
      37479: inst = 32'd203423744;
      37480: inst = 32'd471859200;
      37481: inst = 32'd136314880;
      37482: inst = 32'd268468224;
      37483: inst = 32'd201344295;
      37484: inst = 32'd203423744;
      37485: inst = 32'd471859200;
      37486: inst = 32'd136314880;
      37487: inst = 32'd268468224;
      37488: inst = 32'd201344296;
      37489: inst = 32'd203423744;
      37490: inst = 32'd471859200;
      37491: inst = 32'd136314880;
      37492: inst = 32'd268468224;
      37493: inst = 32'd201344297;
      37494: inst = 32'd203423744;
      37495: inst = 32'd471859200;
      37496: inst = 32'd136314880;
      37497: inst = 32'd268468224;
      37498: inst = 32'd201344298;
      37499: inst = 32'd203423744;
      37500: inst = 32'd471859200;
      37501: inst = 32'd136314880;
      37502: inst = 32'd268468224;
      37503: inst = 32'd201344299;
      37504: inst = 32'd203423744;
      37505: inst = 32'd471859200;
      37506: inst = 32'd136314880;
      37507: inst = 32'd268468224;
      37508: inst = 32'd201344300;
      37509: inst = 32'd203423744;
      37510: inst = 32'd471859200;
      37511: inst = 32'd136314880;
      37512: inst = 32'd268468224;
      37513: inst = 32'd201344301;
      37514: inst = 32'd203483685;
      37515: inst = 32'd471859200;
      37516: inst = 32'd136314880;
      37517: inst = 32'd268468224;
      37518: inst = 32'd201344302;
      37519: inst = 32'd203483685;
      37520: inst = 32'd471859200;
      37521: inst = 32'd136314880;
      37522: inst = 32'd268468224;
      37523: inst = 32'd201344303;
      37524: inst = 32'd203483685;
      37525: inst = 32'd471859200;
      37526: inst = 32'd136314880;
      37527: inst = 32'd268468224;
      37528: inst = 32'd201344304;
      37529: inst = 32'd203483685;
      37530: inst = 32'd471859200;
      37531: inst = 32'd136314880;
      37532: inst = 32'd268468224;
      37533: inst = 32'd201344305;
      37534: inst = 32'd203483685;
      37535: inst = 32'd471859200;
      37536: inst = 32'd136314880;
      37537: inst = 32'd268468224;
      37538: inst = 32'd201344306;
      37539: inst = 32'd203483685;
      37540: inst = 32'd471859200;
      37541: inst = 32'd136314880;
      37542: inst = 32'd268468224;
      37543: inst = 32'd201344307;
      37544: inst = 32'd203483685;
      37545: inst = 32'd471859200;
      37546: inst = 32'd136314880;
      37547: inst = 32'd268468224;
      37548: inst = 32'd201344308;
      37549: inst = 32'd203483685;
      37550: inst = 32'd471859200;
      37551: inst = 32'd136314880;
      37552: inst = 32'd268468224;
      37553: inst = 32'd201344309;
      37554: inst = 32'd203483685;
      37555: inst = 32'd471859200;
      37556: inst = 32'd136314880;
      37557: inst = 32'd268468224;
      37558: inst = 32'd201344310;
      37559: inst = 32'd203483685;
      37560: inst = 32'd471859200;
      37561: inst = 32'd136314880;
      37562: inst = 32'd268468224;
      37563: inst = 32'd201344311;
      37564: inst = 32'd203483685;
      37565: inst = 32'd471859200;
      37566: inst = 32'd136314880;
      37567: inst = 32'd268468224;
      37568: inst = 32'd201344312;
      37569: inst = 32'd203483685;
      37570: inst = 32'd471859200;
      37571: inst = 32'd136314880;
      37572: inst = 32'd268468224;
      37573: inst = 32'd201344313;
      37574: inst = 32'd203483685;
      37575: inst = 32'd471859200;
      37576: inst = 32'd136314880;
      37577: inst = 32'd268468224;
      37578: inst = 32'd201344314;
      37579: inst = 32'd203483685;
      37580: inst = 32'd471859200;
      37581: inst = 32'd136314880;
      37582: inst = 32'd268468224;
      37583: inst = 32'd201344315;
      37584: inst = 32'd203483685;
      37585: inst = 32'd471859200;
      37586: inst = 32'd136314880;
      37587: inst = 32'd268468224;
      37588: inst = 32'd201344316;
      37589: inst = 32'd203483685;
      37590: inst = 32'd471859200;
      37591: inst = 32'd136314880;
      37592: inst = 32'd268468224;
      37593: inst = 32'd201344317;
      37594: inst = 32'd203483685;
      37595: inst = 32'd471859200;
      37596: inst = 32'd136314880;
      37597: inst = 32'd268468224;
      37598: inst = 32'd201344318;
      37599: inst = 32'd203483685;
      37600: inst = 32'd471859200;
      37601: inst = 32'd136314880;
      37602: inst = 32'd268468224;
      37603: inst = 32'd201344319;
      37604: inst = 32'd203483685;
      37605: inst = 32'd471859200;
      37606: inst = 32'd136314880;
      37607: inst = 32'd268468224;
      37608: inst = 32'd201344320;
      37609: inst = 32'd203483685;
      37610: inst = 32'd471859200;
      37611: inst = 32'd136314880;
      37612: inst = 32'd268468224;
      37613: inst = 32'd201344321;
      37614: inst = 32'd203483685;
      37615: inst = 32'd471859200;
      37616: inst = 32'd136314880;
      37617: inst = 32'd268468224;
      37618: inst = 32'd201344322;
      37619: inst = 32'd203483685;
      37620: inst = 32'd471859200;
      37621: inst = 32'd136314880;
      37622: inst = 32'd268468224;
      37623: inst = 32'd201344323;
      37624: inst = 32'd203483685;
      37625: inst = 32'd471859200;
      37626: inst = 32'd136314880;
      37627: inst = 32'd268468224;
      37628: inst = 32'd201344324;
      37629: inst = 32'd203483685;
      37630: inst = 32'd471859200;
      37631: inst = 32'd136314880;
      37632: inst = 32'd268468224;
      37633: inst = 32'd201344325;
      37634: inst = 32'd203483685;
      37635: inst = 32'd471859200;
      37636: inst = 32'd136314880;
      37637: inst = 32'd268468224;
      37638: inst = 32'd201344326;
      37639: inst = 32'd203483685;
      37640: inst = 32'd471859200;
      37641: inst = 32'd136314880;
      37642: inst = 32'd268468224;
      37643: inst = 32'd201344327;
      37644: inst = 32'd203483685;
      37645: inst = 32'd471859200;
      37646: inst = 32'd136314880;
      37647: inst = 32'd268468224;
      37648: inst = 32'd201344328;
      37649: inst = 32'd203483685;
      37650: inst = 32'd471859200;
      37651: inst = 32'd136314880;
      37652: inst = 32'd268468224;
      37653: inst = 32'd201344329;
      37654: inst = 32'd203483685;
      37655: inst = 32'd471859200;
      37656: inst = 32'd136314880;
      37657: inst = 32'd268468224;
      37658: inst = 32'd201344330;
      37659: inst = 32'd203483685;
      37660: inst = 32'd471859200;
      37661: inst = 32'd136314880;
      37662: inst = 32'd268468224;
      37663: inst = 32'd201344331;
      37664: inst = 32'd203483685;
      37665: inst = 32'd471859200;
      37666: inst = 32'd136314880;
      37667: inst = 32'd268468224;
      37668: inst = 32'd201344332;
      37669: inst = 32'd203483685;
      37670: inst = 32'd471859200;
      37671: inst = 32'd136314880;
      37672: inst = 32'd268468224;
      37673: inst = 32'd201344333;
      37674: inst = 32'd203483685;
      37675: inst = 32'd471859200;
      37676: inst = 32'd136314880;
      37677: inst = 32'd268468224;
      37678: inst = 32'd201344334;
      37679: inst = 32'd203483685;
      37680: inst = 32'd471859200;
      37681: inst = 32'd136314880;
      37682: inst = 32'd268468224;
      37683: inst = 32'd201344335;
      37684: inst = 32'd203423744;
      37685: inst = 32'd471859200;
      37686: inst = 32'd136314880;
      37687: inst = 32'd268468224;
      37688: inst = 32'd201344336;
      37689: inst = 32'd203423744;
      37690: inst = 32'd471859200;
      37691: inst = 32'd136314880;
      37692: inst = 32'd268468224;
      37693: inst = 32'd201344337;
      37694: inst = 32'd203483685;
      37695: inst = 32'd471859200;
      37696: inst = 32'd136314880;
      37697: inst = 32'd268468224;
      37698: inst = 32'd201344338;
      37699: inst = 32'd203483685;
      37700: inst = 32'd471859200;
      37701: inst = 32'd136314880;
      37702: inst = 32'd268468224;
      37703: inst = 32'd201344339;
      37704: inst = 32'd203483685;
      37705: inst = 32'd471859200;
      37706: inst = 32'd136314880;
      37707: inst = 32'd268468224;
      37708: inst = 32'd201344340;
      37709: inst = 32'd203483685;
      37710: inst = 32'd471859200;
      37711: inst = 32'd136314880;
      37712: inst = 32'd268468224;
      37713: inst = 32'd201344341;
      37714: inst = 32'd203483685;
      37715: inst = 32'd471859200;
      37716: inst = 32'd136314880;
      37717: inst = 32'd268468224;
      37718: inst = 32'd201344342;
      37719: inst = 32'd203483685;
      37720: inst = 32'd471859200;
      37721: inst = 32'd136314880;
      37722: inst = 32'd268468224;
      37723: inst = 32'd201344343;
      37724: inst = 32'd203483685;
      37725: inst = 32'd471859200;
      37726: inst = 32'd136314880;
      37727: inst = 32'd268468224;
      37728: inst = 32'd201344344;
      37729: inst = 32'd203483685;
      37730: inst = 32'd471859200;
      37731: inst = 32'd136314880;
      37732: inst = 32'd268468224;
      37733: inst = 32'd201344345;
      37734: inst = 32'd203483685;
      37735: inst = 32'd471859200;
      37736: inst = 32'd136314880;
      37737: inst = 32'd268468224;
      37738: inst = 32'd201344346;
      37739: inst = 32'd203483685;
      37740: inst = 32'd471859200;
      37741: inst = 32'd136314880;
      37742: inst = 32'd268468224;
      37743: inst = 32'd201344347;
      37744: inst = 32'd203483685;
      37745: inst = 32'd471859200;
      37746: inst = 32'd136314880;
      37747: inst = 32'd268468224;
      37748: inst = 32'd201344348;
      37749: inst = 32'd203483685;
      37750: inst = 32'd471859200;
      37751: inst = 32'd136314880;
      37752: inst = 32'd268468224;
      37753: inst = 32'd201344349;
      37754: inst = 32'd203483685;
      37755: inst = 32'd471859200;
      37756: inst = 32'd136314880;
      37757: inst = 32'd268468224;
      37758: inst = 32'd201344350;
      37759: inst = 32'd203483685;
      37760: inst = 32'd471859200;
      37761: inst = 32'd136314880;
      37762: inst = 32'd268468224;
      37763: inst = 32'd201344351;
      37764: inst = 32'd203483685;
      37765: inst = 32'd471859200;
      37766: inst = 32'd136314880;
      37767: inst = 32'd268468224;
      37768: inst = 32'd201344352;
      37769: inst = 32'd203483685;
      37770: inst = 32'd471859200;
      37771: inst = 32'd136314880;
      37772: inst = 32'd268468224;
      37773: inst = 32'd201344353;
      37774: inst = 32'd203483685;
      37775: inst = 32'd471859200;
      37776: inst = 32'd136314880;
      37777: inst = 32'd268468224;
      37778: inst = 32'd201344354;
      37779: inst = 32'd203483685;
      37780: inst = 32'd471859200;
      37781: inst = 32'd136314880;
      37782: inst = 32'd268468224;
      37783: inst = 32'd201344355;
      37784: inst = 32'd203483685;
      37785: inst = 32'd471859200;
      37786: inst = 32'd136314880;
      37787: inst = 32'd268468224;
      37788: inst = 32'd201344356;
      37789: inst = 32'd203483685;
      37790: inst = 32'd471859200;
      37791: inst = 32'd136314880;
      37792: inst = 32'd268468224;
      37793: inst = 32'd201344357;
      37794: inst = 32'd203483685;
      37795: inst = 32'd471859200;
      37796: inst = 32'd136314880;
      37797: inst = 32'd268468224;
      37798: inst = 32'd201344358;
      37799: inst = 32'd203483685;
      37800: inst = 32'd471859200;
      37801: inst = 32'd136314880;
      37802: inst = 32'd268468224;
      37803: inst = 32'd201344359;
      37804: inst = 32'd203483685;
      37805: inst = 32'd471859200;
      37806: inst = 32'd136314880;
      37807: inst = 32'd268468224;
      37808: inst = 32'd201344360;
      37809: inst = 32'd203483685;
      37810: inst = 32'd471859200;
      37811: inst = 32'd136314880;
      37812: inst = 32'd268468224;
      37813: inst = 32'd201344361;
      37814: inst = 32'd203423744;
      37815: inst = 32'd471859200;
      37816: inst = 32'd136314880;
      37817: inst = 32'd268468224;
      37818: inst = 32'd201344362;
      37819: inst = 32'd203483685;
      37820: inst = 32'd471859200;
      37821: inst = 32'd136314880;
      37822: inst = 32'd268468224;
      37823: inst = 32'd201344363;
      37824: inst = 32'd203483685;
      37825: inst = 32'd471859200;
      37826: inst = 32'd136314880;
      37827: inst = 32'd268468224;
      37828: inst = 32'd201344364;
      37829: inst = 32'd203483685;
      37830: inst = 32'd471859200;
      37831: inst = 32'd136314880;
      37832: inst = 32'd268468224;
      37833: inst = 32'd201344365;
      37834: inst = 32'd203483685;
      37835: inst = 32'd471859200;
      37836: inst = 32'd136314880;
      37837: inst = 32'd268468224;
      37838: inst = 32'd201344366;
      37839: inst = 32'd203483685;
      37840: inst = 32'd471859200;
      37841: inst = 32'd136314880;
      37842: inst = 32'd268468224;
      37843: inst = 32'd201344367;
      37844: inst = 32'd203483685;
      37845: inst = 32'd471859200;
      37846: inst = 32'd136314880;
      37847: inst = 32'd268468224;
      37848: inst = 32'd201344368;
      37849: inst = 32'd203483685;
      37850: inst = 32'd471859200;
      37851: inst = 32'd136314880;
      37852: inst = 32'd268468224;
      37853: inst = 32'd201344369;
      37854: inst = 32'd203483685;
      37855: inst = 32'd471859200;
      37856: inst = 32'd136314880;
      37857: inst = 32'd268468224;
      37858: inst = 32'd201344370;
      37859: inst = 32'd203483685;
      37860: inst = 32'd471859200;
      37861: inst = 32'd136314880;
      37862: inst = 32'd268468224;
      37863: inst = 32'd201344371;
      37864: inst = 32'd203483685;
      37865: inst = 32'd471859200;
      37866: inst = 32'd136314880;
      37867: inst = 32'd268468224;
      37868: inst = 32'd201344372;
      37869: inst = 32'd203483685;
      37870: inst = 32'd471859200;
      37871: inst = 32'd136314880;
      37872: inst = 32'd268468224;
      37873: inst = 32'd201344373;
      37874: inst = 32'd203483685;
      37875: inst = 32'd471859200;
      37876: inst = 32'd136314880;
      37877: inst = 32'd268468224;
      37878: inst = 32'd201344374;
      37879: inst = 32'd203423744;
      37880: inst = 32'd471859200;
      37881: inst = 32'd136314880;
      37882: inst = 32'd268468224;
      37883: inst = 32'd201344375;
      37884: inst = 32'd203423744;
      37885: inst = 32'd471859200;
      37886: inst = 32'd136314880;
      37887: inst = 32'd268468224;
      37888: inst = 32'd201344376;
      37889: inst = 32'd203423744;
      37890: inst = 32'd471859200;
      37891: inst = 32'd136314880;
      37892: inst = 32'd268468224;
      37893: inst = 32'd201344377;
      37894: inst = 32'd203423744;
      37895: inst = 32'd471859200;
      37896: inst = 32'd136314880;
      37897: inst = 32'd268468224;
      37898: inst = 32'd201344378;
      37899: inst = 32'd203423744;
      37900: inst = 32'd471859200;
      37901: inst = 32'd136314880;
      37902: inst = 32'd268468224;
      37903: inst = 32'd201344379;
      37904: inst = 32'd203423744;
      37905: inst = 32'd471859200;
      37906: inst = 32'd136314880;
      37907: inst = 32'd268468224;
      37908: inst = 32'd201344380;
      37909: inst = 32'd203423744;
      37910: inst = 32'd471859200;
      37911: inst = 32'd136314880;
      37912: inst = 32'd268468224;
      37913: inst = 32'd201344381;
      37914: inst = 32'd203423744;
      37915: inst = 32'd471859200;
      37916: inst = 32'd136314880;
      37917: inst = 32'd268468224;
      37918: inst = 32'd201344382;
      37919: inst = 32'd203423744;
      37920: inst = 32'd471859200;
      37921: inst = 32'd136314880;
      37922: inst = 32'd268468224;
      37923: inst = 32'd201344383;
      37924: inst = 32'd203423744;
      37925: inst = 32'd471859200;
      37926: inst = 32'd136314880;
      37927: inst = 32'd268468224;
      37928: inst = 32'd201344384;
      37929: inst = 32'd203423744;
      37930: inst = 32'd471859200;
      37931: inst = 32'd136314880;
      37932: inst = 32'd268468224;
      37933: inst = 32'd201344385;
      37934: inst = 32'd203423744;
      37935: inst = 32'd471859200;
      37936: inst = 32'd136314880;
      37937: inst = 32'd268468224;
      37938: inst = 32'd201344386;
      37939: inst = 32'd203423744;
      37940: inst = 32'd471859200;
      37941: inst = 32'd136314880;
      37942: inst = 32'd268468224;
      37943: inst = 32'd201344387;
      37944: inst = 32'd203423744;
      37945: inst = 32'd471859200;
      37946: inst = 32'd136314880;
      37947: inst = 32'd268468224;
      37948: inst = 32'd201344388;
      37949: inst = 32'd203423744;
      37950: inst = 32'd471859200;
      37951: inst = 32'd136314880;
      37952: inst = 32'd268468224;
      37953: inst = 32'd201344389;
      37954: inst = 32'd203423744;
      37955: inst = 32'd471859200;
      37956: inst = 32'd136314880;
      37957: inst = 32'd268468224;
      37958: inst = 32'd201344390;
      37959: inst = 32'd203423744;
      37960: inst = 32'd471859200;
      37961: inst = 32'd136314880;
      37962: inst = 32'd268468224;
      37963: inst = 32'd201344391;
      37964: inst = 32'd203423744;
      37965: inst = 32'd471859200;
      37966: inst = 32'd136314880;
      37967: inst = 32'd268468224;
      37968: inst = 32'd201344392;
      37969: inst = 32'd203423744;
      37970: inst = 32'd471859200;
      37971: inst = 32'd136314880;
      37972: inst = 32'd268468224;
      37973: inst = 32'd201344393;
      37974: inst = 32'd203423744;
      37975: inst = 32'd471859200;
      37976: inst = 32'd136314880;
      37977: inst = 32'd268468224;
      37978: inst = 32'd201344394;
      37979: inst = 32'd203423744;
      37980: inst = 32'd471859200;
      37981: inst = 32'd136314880;
      37982: inst = 32'd268468224;
      37983: inst = 32'd201344395;
      37984: inst = 32'd203423744;
      37985: inst = 32'd471859200;
      37986: inst = 32'd136314880;
      37987: inst = 32'd268468224;
      37988: inst = 32'd201344396;
      37989: inst = 32'd203423744;
      37990: inst = 32'd471859200;
      37991: inst = 32'd136314880;
      37992: inst = 32'd268468224;
      37993: inst = 32'd201344397;
      37994: inst = 32'd203483685;
      37995: inst = 32'd471859200;
      37996: inst = 32'd136314880;
      37997: inst = 32'd268468224;
      37998: inst = 32'd201344398;
      37999: inst = 32'd203483685;
      38000: inst = 32'd471859200;
      38001: inst = 32'd136314880;
      38002: inst = 32'd268468224;
      38003: inst = 32'd201344399;
      38004: inst = 32'd203483685;
      38005: inst = 32'd471859200;
      38006: inst = 32'd136314880;
      38007: inst = 32'd268468224;
      38008: inst = 32'd201344400;
      38009: inst = 32'd203423744;
      38010: inst = 32'd471859200;
      38011: inst = 32'd136314880;
      38012: inst = 32'd268468224;
      38013: inst = 32'd201344401;
      38014: inst = 32'd203423744;
      38015: inst = 32'd471859200;
      38016: inst = 32'd136314880;
      38017: inst = 32'd268468224;
      38018: inst = 32'd201344402;
      38019: inst = 32'd203423744;
      38020: inst = 32'd471859200;
      38021: inst = 32'd136314880;
      38022: inst = 32'd268468224;
      38023: inst = 32'd201344403;
      38024: inst = 32'd203423744;
      38025: inst = 32'd471859200;
      38026: inst = 32'd136314880;
      38027: inst = 32'd268468224;
      38028: inst = 32'd201344404;
      38029: inst = 32'd203423744;
      38030: inst = 32'd471859200;
      38031: inst = 32'd136314880;
      38032: inst = 32'd268468224;
      38033: inst = 32'd201344405;
      38034: inst = 32'd203423744;
      38035: inst = 32'd471859200;
      38036: inst = 32'd136314880;
      38037: inst = 32'd268468224;
      38038: inst = 32'd201344406;
      38039: inst = 32'd203423744;
      38040: inst = 32'd471859200;
      38041: inst = 32'd136314880;
      38042: inst = 32'd268468224;
      38043: inst = 32'd201344407;
      38044: inst = 32'd203423744;
      38045: inst = 32'd471859200;
      38046: inst = 32'd136314880;
      38047: inst = 32'd268468224;
      38048: inst = 32'd201344408;
      38049: inst = 32'd203483685;
      38050: inst = 32'd471859200;
      38051: inst = 32'd136314880;
      38052: inst = 32'd268468224;
      38053: inst = 32'd201344409;
      38054: inst = 32'd203483685;
      38055: inst = 32'd471859200;
      38056: inst = 32'd136314880;
      38057: inst = 32'd268468224;
      38058: inst = 32'd201344410;
      38059: inst = 32'd203483685;
      38060: inst = 32'd471859200;
      38061: inst = 32'd136314880;
      38062: inst = 32'd268468224;
      38063: inst = 32'd201344411;
      38064: inst = 32'd203483685;
      38065: inst = 32'd471859200;
      38066: inst = 32'd136314880;
      38067: inst = 32'd268468224;
      38068: inst = 32'd201344412;
      38069: inst = 32'd203423744;
      38070: inst = 32'd471859200;
      38071: inst = 32'd136314880;
      38072: inst = 32'd268468224;
      38073: inst = 32'd201344413;
      38074: inst = 32'd203423744;
      38075: inst = 32'd471859200;
      38076: inst = 32'd136314880;
      38077: inst = 32'd268468224;
      38078: inst = 32'd201344414;
      38079: inst = 32'd203423744;
      38080: inst = 32'd471859200;
      38081: inst = 32'd136314880;
      38082: inst = 32'd268468224;
      38083: inst = 32'd201344415;
      38084: inst = 32'd203423744;
      38085: inst = 32'd471859200;
      38086: inst = 32'd136314880;
      38087: inst = 32'd268468224;
      38088: inst = 32'd201344416;
      38089: inst = 32'd203423744;
      38090: inst = 32'd471859200;
      38091: inst = 32'd136314880;
      38092: inst = 32'd268468224;
      38093: inst = 32'd201344417;
      38094: inst = 32'd203423744;
      38095: inst = 32'd471859200;
      38096: inst = 32'd136314880;
      38097: inst = 32'd268468224;
      38098: inst = 32'd201344418;
      38099: inst = 32'd203423744;
      38100: inst = 32'd471859200;
      38101: inst = 32'd136314880;
      38102: inst = 32'd268468224;
      38103: inst = 32'd201344419;
      38104: inst = 32'd203423744;
      38105: inst = 32'd471859200;
      38106: inst = 32'd136314880;
      38107: inst = 32'd268468224;
      38108: inst = 32'd201344420;
      38109: inst = 32'd203423744;
      38110: inst = 32'd471859200;
      38111: inst = 32'd136314880;
      38112: inst = 32'd268468224;
      38113: inst = 32'd201344421;
      38114: inst = 32'd203423744;
      38115: inst = 32'd471859200;
      38116: inst = 32'd136314880;
      38117: inst = 32'd268468224;
      38118: inst = 32'd201344422;
      38119: inst = 32'd203423744;
      38120: inst = 32'd471859200;
      38121: inst = 32'd136314880;
      38122: inst = 32'd268468224;
      38123: inst = 32'd201344423;
      38124: inst = 32'd203423744;
      38125: inst = 32'd471859200;
      38126: inst = 32'd136314880;
      38127: inst = 32'd268468224;
      38128: inst = 32'd201344424;
      38129: inst = 32'd203423744;
      38130: inst = 32'd471859200;
      38131: inst = 32'd136314880;
      38132: inst = 32'd268468224;
      38133: inst = 32'd201344425;
      38134: inst = 32'd203483685;
      38135: inst = 32'd471859200;
      38136: inst = 32'd136314880;
      38137: inst = 32'd268468224;
      38138: inst = 32'd201344426;
      38139: inst = 32'd203483685;
      38140: inst = 32'd471859200;
      38141: inst = 32'd136314880;
      38142: inst = 32'd268468224;
      38143: inst = 32'd201344427;
      38144: inst = 32'd203483685;
      38145: inst = 32'd471859200;
      38146: inst = 32'd136314880;
      38147: inst = 32'd268468224;
      38148: inst = 32'd201344428;
      38149: inst = 32'd203483685;
      38150: inst = 32'd471859200;
      38151: inst = 32'd136314880;
      38152: inst = 32'd268468224;
      38153: inst = 32'd201344429;
      38154: inst = 32'd203483685;
      38155: inst = 32'd471859200;
      38156: inst = 32'd136314880;
      38157: inst = 32'd268468224;
      38158: inst = 32'd201344430;
      38159: inst = 32'd203423744;
      38160: inst = 32'd471859200;
      38161: inst = 32'd136314880;
      38162: inst = 32'd268468224;
      38163: inst = 32'd201344431;
      38164: inst = 32'd203423744;
      38165: inst = 32'd471859200;
      38166: inst = 32'd136314880;
      38167: inst = 32'd268468224;
      38168: inst = 32'd201344432;
      38169: inst = 32'd203423744;
      38170: inst = 32'd471859200;
      38171: inst = 32'd136314880;
      38172: inst = 32'd268468224;
      38173: inst = 32'd201344433;
      38174: inst = 32'd203483685;
      38175: inst = 32'd471859200;
      38176: inst = 32'd136314880;
      38177: inst = 32'd268468224;
      38178: inst = 32'd201344434;
      38179: inst = 32'd203483685;
      38180: inst = 32'd471859200;
      38181: inst = 32'd136314880;
      38182: inst = 32'd268468224;
      38183: inst = 32'd201344435;
      38184: inst = 32'd203483685;
      38185: inst = 32'd471859200;
      38186: inst = 32'd136314880;
      38187: inst = 32'd268468224;
      38188: inst = 32'd201344436;
      38189: inst = 32'd203423744;
      38190: inst = 32'd471859200;
      38191: inst = 32'd136314880;
      38192: inst = 32'd268468224;
      38193: inst = 32'd201344437;
      38194: inst = 32'd203423744;
      38195: inst = 32'd471859200;
      38196: inst = 32'd136314880;
      38197: inst = 32'd268468224;
      38198: inst = 32'd201344438;
      38199: inst = 32'd203483685;
      38200: inst = 32'd471859200;
      38201: inst = 32'd136314880;
      38202: inst = 32'd268468224;
      38203: inst = 32'd201344439;
      38204: inst = 32'd203483685;
      38205: inst = 32'd471859200;
      38206: inst = 32'd136314880;
      38207: inst = 32'd268468224;
      38208: inst = 32'd201344440;
      38209: inst = 32'd203483685;
      38210: inst = 32'd471859200;
      38211: inst = 32'd136314880;
      38212: inst = 32'd268468224;
      38213: inst = 32'd201344441;
      38214: inst = 32'd203483685;
      38215: inst = 32'd471859200;
      38216: inst = 32'd136314880;
      38217: inst = 32'd268468224;
      38218: inst = 32'd201344442;
      38219: inst = 32'd203483685;
      38220: inst = 32'd471859200;
      38221: inst = 32'd136314880;
      38222: inst = 32'd268468224;
      38223: inst = 32'd201344443;
      38224: inst = 32'd203483685;
      38225: inst = 32'd471859200;
      38226: inst = 32'd136314880;
      38227: inst = 32'd268468224;
      38228: inst = 32'd201344444;
      38229: inst = 32'd203483685;
      38230: inst = 32'd471859200;
      38231: inst = 32'd136314880;
      38232: inst = 32'd268468224;
      38233: inst = 32'd201344445;
      38234: inst = 32'd203483685;
      38235: inst = 32'd471859200;
      38236: inst = 32'd136314880;
      38237: inst = 32'd268468224;
      38238: inst = 32'd201344446;
      38239: inst = 32'd203423744;
      38240: inst = 32'd471859200;
      38241: inst = 32'd136314880;
      38242: inst = 32'd268468224;
      38243: inst = 32'd201344447;
      38244: inst = 32'd203423744;
      38245: inst = 32'd471859200;
      38246: inst = 32'd136314880;
      38247: inst = 32'd268468224;
      38248: inst = 32'd201344448;
      38249: inst = 32'd203423744;
      38250: inst = 32'd471859200;
      38251: inst = 32'd136314880;
      38252: inst = 32'd268468224;
      38253: inst = 32'd201344449;
      38254: inst = 32'd203423744;
      38255: inst = 32'd471859200;
      38256: inst = 32'd136314880;
      38257: inst = 32'd268468224;
      38258: inst = 32'd201344450;
      38259: inst = 32'd203483685;
      38260: inst = 32'd471859200;
      38261: inst = 32'd136314880;
      38262: inst = 32'd268468224;
      38263: inst = 32'd201344451;
      38264: inst = 32'd203483685;
      38265: inst = 32'd471859200;
      38266: inst = 32'd136314880;
      38267: inst = 32'd268468224;
      38268: inst = 32'd201344452;
      38269: inst = 32'd203483685;
      38270: inst = 32'd471859200;
      38271: inst = 32'd136314880;
      38272: inst = 32'd268468224;
      38273: inst = 32'd201344453;
      38274: inst = 32'd203483685;
      38275: inst = 32'd471859200;
      38276: inst = 32'd136314880;
      38277: inst = 32'd268468224;
      38278: inst = 32'd201344454;
      38279: inst = 32'd203483685;
      38280: inst = 32'd471859200;
      38281: inst = 32'd136314880;
      38282: inst = 32'd268468224;
      38283: inst = 32'd201344455;
      38284: inst = 32'd203483685;
      38285: inst = 32'd471859200;
      38286: inst = 32'd136314880;
      38287: inst = 32'd268468224;
      38288: inst = 32'd201344456;
      38289: inst = 32'd203423744;
      38290: inst = 32'd471859200;
      38291: inst = 32'd136314880;
      38292: inst = 32'd268468224;
      38293: inst = 32'd201344457;
      38294: inst = 32'd203423744;
      38295: inst = 32'd471859200;
      38296: inst = 32'd136314880;
      38297: inst = 32'd268468224;
      38298: inst = 32'd201344458;
      38299: inst = 32'd203483685;
      38300: inst = 32'd471859200;
      38301: inst = 32'd136314880;
      38302: inst = 32'd268468224;
      38303: inst = 32'd201344459;
      38304: inst = 32'd203483685;
      38305: inst = 32'd471859200;
      38306: inst = 32'd136314880;
      38307: inst = 32'd268468224;
      38308: inst = 32'd201344460;
      38309: inst = 32'd203483685;
      38310: inst = 32'd471859200;
      38311: inst = 32'd136314880;
      38312: inst = 32'd268468224;
      38313: inst = 32'd201344461;
      38314: inst = 32'd203483685;
      38315: inst = 32'd471859200;
      38316: inst = 32'd136314880;
      38317: inst = 32'd268468224;
      38318: inst = 32'd201344462;
      38319: inst = 32'd203423744;
      38320: inst = 32'd471859200;
      38321: inst = 32'd136314880;
      38322: inst = 32'd268468224;
      38323: inst = 32'd201344463;
      38324: inst = 32'd203423744;
      38325: inst = 32'd471859200;
      38326: inst = 32'd136314880;
      38327: inst = 32'd268468224;
      38328: inst = 32'd201344464;
      38329: inst = 32'd203423744;
      38330: inst = 32'd471859200;
      38331: inst = 32'd136314880;
      38332: inst = 32'd268468224;
      38333: inst = 32'd201344465;
      38334: inst = 32'd203423744;
      38335: inst = 32'd471859200;
      38336: inst = 32'd136314880;
      38337: inst = 32'd268468224;
      38338: inst = 32'd201344466;
      38339: inst = 32'd203423744;
      38340: inst = 32'd471859200;
      38341: inst = 32'd136314880;
      38342: inst = 32'd268468224;
      38343: inst = 32'd201344467;
      38344: inst = 32'd203423744;
      38345: inst = 32'd471859200;
      38346: inst = 32'd136314880;
      38347: inst = 32'd268468224;
      38348: inst = 32'd201344468;
      38349: inst = 32'd203423744;
      38350: inst = 32'd471859200;
      38351: inst = 32'd136314880;
      38352: inst = 32'd268468224;
      38353: inst = 32'd201344469;
      38354: inst = 32'd203423744;
      38355: inst = 32'd471859200;
      38356: inst = 32'd136314880;
      38357: inst = 32'd268468224;
      38358: inst = 32'd201344470;
      38359: inst = 32'd203423744;
      38360: inst = 32'd471859200;
      38361: inst = 32'd136314880;
      38362: inst = 32'd268468224;
      38363: inst = 32'd201344471;
      38364: inst = 32'd203423744;
      38365: inst = 32'd471859200;
      38366: inst = 32'd136314880;
      38367: inst = 32'd268468224;
      38368: inst = 32'd201344472;
      38369: inst = 32'd203423744;
      38370: inst = 32'd471859200;
      38371: inst = 32'd136314880;
      38372: inst = 32'd268468224;
      38373: inst = 32'd201344473;
      38374: inst = 32'd203423744;
      38375: inst = 32'd471859200;
      38376: inst = 32'd136314880;
      38377: inst = 32'd268468224;
      38378: inst = 32'd201344474;
      38379: inst = 32'd203423744;
      38380: inst = 32'd471859200;
      38381: inst = 32'd136314880;
      38382: inst = 32'd268468224;
      38383: inst = 32'd201344475;
      38384: inst = 32'd203423744;
      38385: inst = 32'd471859200;
      38386: inst = 32'd136314880;
      38387: inst = 32'd268468224;
      38388: inst = 32'd201344476;
      38389: inst = 32'd203423744;
      38390: inst = 32'd471859200;
      38391: inst = 32'd136314880;
      38392: inst = 32'd268468224;
      38393: inst = 32'd201344477;
      38394: inst = 32'd203423744;
      38395: inst = 32'd471859200;
      38396: inst = 32'd136314880;
      38397: inst = 32'd268468224;
      38398: inst = 32'd201344478;
      38399: inst = 32'd203423744;
      38400: inst = 32'd471859200;
      38401: inst = 32'd136314880;
      38402: inst = 32'd268468224;
      38403: inst = 32'd201344479;
      38404: inst = 32'd203423744;
      38405: inst = 32'd471859200;
      38406: inst = 32'd136314880;
      38407: inst = 32'd268468224;
      38408: inst = 32'd201344480;
      38409: inst = 32'd203423744;
      38410: inst = 32'd471859200;
      38411: inst = 32'd136314880;
      38412: inst = 32'd268468224;
      38413: inst = 32'd201344481;
      38414: inst = 32'd203423744;
      38415: inst = 32'd471859200;
      38416: inst = 32'd136314880;
      38417: inst = 32'd268468224;
      38418: inst = 32'd201344482;
      38419: inst = 32'd203423744;
      38420: inst = 32'd471859200;
      38421: inst = 32'd136314880;
      38422: inst = 32'd268468224;
      38423: inst = 32'd201344483;
      38424: inst = 32'd203423744;
      38425: inst = 32'd471859200;
      38426: inst = 32'd136314880;
      38427: inst = 32'd268468224;
      38428: inst = 32'd201344484;
      38429: inst = 32'd203423744;
      38430: inst = 32'd471859200;
      38431: inst = 32'd136314880;
      38432: inst = 32'd268468224;
      38433: inst = 32'd201344485;
      38434: inst = 32'd203423744;
      38435: inst = 32'd471859200;
      38436: inst = 32'd136314880;
      38437: inst = 32'd268468224;
      38438: inst = 32'd201344486;
      38439: inst = 32'd203423744;
      38440: inst = 32'd471859200;
      38441: inst = 32'd136314880;
      38442: inst = 32'd268468224;
      38443: inst = 32'd201344487;
      38444: inst = 32'd203423744;
      38445: inst = 32'd471859200;
      38446: inst = 32'd136314880;
      38447: inst = 32'd268468224;
      38448: inst = 32'd201344488;
      38449: inst = 32'd203423744;
      38450: inst = 32'd471859200;
      38451: inst = 32'd136314880;
      38452: inst = 32'd268468224;
      38453: inst = 32'd201344489;
      38454: inst = 32'd203423744;
      38455: inst = 32'd471859200;
      38456: inst = 32'd136314880;
      38457: inst = 32'd268468224;
      38458: inst = 32'd201344490;
      38459: inst = 32'd203423744;
      38460: inst = 32'd471859200;
      38461: inst = 32'd136314880;
      38462: inst = 32'd268468224;
      38463: inst = 32'd201344491;
      38464: inst = 32'd203423744;
      38465: inst = 32'd471859200;
      38466: inst = 32'd136314880;
      38467: inst = 32'd268468224;
      38468: inst = 32'd201344492;
      38469: inst = 32'd203423744;
      38470: inst = 32'd471859200;
      38471: inst = 32'd136314880;
      38472: inst = 32'd268468224;
      38473: inst = 32'd201344493;
      38474: inst = 32'd203483685;
      38475: inst = 32'd471859200;
      38476: inst = 32'd136314880;
      38477: inst = 32'd268468224;
      38478: inst = 32'd201344494;
      38479: inst = 32'd203483685;
      38480: inst = 32'd471859200;
      38481: inst = 32'd136314880;
      38482: inst = 32'd268468224;
      38483: inst = 32'd201344495;
      38484: inst = 32'd203483685;
      38485: inst = 32'd471859200;
      38486: inst = 32'd136314880;
      38487: inst = 32'd268468224;
      38488: inst = 32'd201344496;
      38489: inst = 32'd203483685;
      38490: inst = 32'd471859200;
      38491: inst = 32'd136314880;
      38492: inst = 32'd268468224;
      38493: inst = 32'd201344497;
      38494: inst = 32'd203483685;
      38495: inst = 32'd471859200;
      38496: inst = 32'd136314880;
      38497: inst = 32'd268468224;
      38498: inst = 32'd201344498;
      38499: inst = 32'd203483685;
      38500: inst = 32'd471859200;
      38501: inst = 32'd136314880;
      38502: inst = 32'd268468224;
      38503: inst = 32'd201344499;
      38504: inst = 32'd203483685;
      38505: inst = 32'd471859200;
      38506: inst = 32'd136314880;
      38507: inst = 32'd268468224;
      38508: inst = 32'd201344500;
      38509: inst = 32'd203483685;
      38510: inst = 32'd471859200;
      38511: inst = 32'd136314880;
      38512: inst = 32'd268468224;
      38513: inst = 32'd201344501;
      38514: inst = 32'd203423744;
      38515: inst = 32'd471859200;
      38516: inst = 32'd136314880;
      38517: inst = 32'd268468224;
      38518: inst = 32'd201344502;
      38519: inst = 32'd203423744;
      38520: inst = 32'd471859200;
      38521: inst = 32'd136314880;
      38522: inst = 32'd268468224;
      38523: inst = 32'd201344503;
      38524: inst = 32'd203423744;
      38525: inst = 32'd471859200;
      38526: inst = 32'd136314880;
      38527: inst = 32'd268468224;
      38528: inst = 32'd201344504;
      38529: inst = 32'd203483685;
      38530: inst = 32'd471859200;
      38531: inst = 32'd136314880;
      38532: inst = 32'd268468224;
      38533: inst = 32'd201344505;
      38534: inst = 32'd203483685;
      38535: inst = 32'd471859200;
      38536: inst = 32'd136314880;
      38537: inst = 32'd268468224;
      38538: inst = 32'd201344506;
      38539: inst = 32'd203483685;
      38540: inst = 32'd471859200;
      38541: inst = 32'd136314880;
      38542: inst = 32'd268468224;
      38543: inst = 32'd201344507;
      38544: inst = 32'd203483685;
      38545: inst = 32'd471859200;
      38546: inst = 32'd136314880;
      38547: inst = 32'd268468224;
      38548: inst = 32'd201344508;
      38549: inst = 32'd203483685;
      38550: inst = 32'd471859200;
      38551: inst = 32'd136314880;
      38552: inst = 32'd268468224;
      38553: inst = 32'd201344509;
      38554: inst = 32'd203483685;
      38555: inst = 32'd471859200;
      38556: inst = 32'd136314880;
      38557: inst = 32'd268468224;
      38558: inst = 32'd201344510;
      38559: inst = 32'd203483685;
      38560: inst = 32'd471859200;
      38561: inst = 32'd136314880;
      38562: inst = 32'd268468224;
      38563: inst = 32'd201344511;
      38564: inst = 32'd203483685;
      38565: inst = 32'd471859200;
      38566: inst = 32'd136314880;
      38567: inst = 32'd268468224;
      38568: inst = 32'd201344512;
      38569: inst = 32'd203483685;
      38570: inst = 32'd471859200;
      38571: inst = 32'd136314880;
      38572: inst = 32'd268468224;
      38573: inst = 32'd201344513;
      38574: inst = 32'd203423744;
      38575: inst = 32'd471859200;
      38576: inst = 32'd136314880;
      38577: inst = 32'd268468224;
      38578: inst = 32'd201344514;
      38579: inst = 32'd203423744;
      38580: inst = 32'd471859200;
      38581: inst = 32'd136314880;
      38582: inst = 32'd268468224;
      38583: inst = 32'd201344515;
      38584: inst = 32'd203423744;
      38585: inst = 32'd471859200;
      38586: inst = 32'd136314880;
      38587: inst = 32'd268468224;
      38588: inst = 32'd201344516;
      38589: inst = 32'd203423744;
      38590: inst = 32'd471859200;
      38591: inst = 32'd136314880;
      38592: inst = 32'd268468224;
      38593: inst = 32'd201344517;
      38594: inst = 32'd203423744;
      38595: inst = 32'd471859200;
      38596: inst = 32'd136314880;
      38597: inst = 32'd268468224;
      38598: inst = 32'd201344518;
      38599: inst = 32'd203423744;
      38600: inst = 32'd471859200;
      38601: inst = 32'd136314880;
      38602: inst = 32'd268468224;
      38603: inst = 32'd201344519;
      38604: inst = 32'd203423744;
      38605: inst = 32'd471859200;
      38606: inst = 32'd136314880;
      38607: inst = 32'd268468224;
      38608: inst = 32'd201344520;
      38609: inst = 32'd203483685;
      38610: inst = 32'd471859200;
      38611: inst = 32'd136314880;
      38612: inst = 32'd268468224;
      38613: inst = 32'd201344521;
      38614: inst = 32'd203483685;
      38615: inst = 32'd471859200;
      38616: inst = 32'd136314880;
      38617: inst = 32'd268468224;
      38618: inst = 32'd201344522;
      38619: inst = 32'd203483685;
      38620: inst = 32'd471859200;
      38621: inst = 32'd136314880;
      38622: inst = 32'd268468224;
      38623: inst = 32'd201344523;
      38624: inst = 32'd203483685;
      38625: inst = 32'd471859200;
      38626: inst = 32'd136314880;
      38627: inst = 32'd268468224;
      38628: inst = 32'd201344524;
      38629: inst = 32'd203483685;
      38630: inst = 32'd471859200;
      38631: inst = 32'd136314880;
      38632: inst = 32'd268468224;
      38633: inst = 32'd201344525;
      38634: inst = 32'd203423744;
      38635: inst = 32'd471859200;
      38636: inst = 32'd136314880;
      38637: inst = 32'd268468224;
      38638: inst = 32'd201344526;
      38639: inst = 32'd203423744;
      38640: inst = 32'd471859200;
      38641: inst = 32'd136314880;
      38642: inst = 32'd268468224;
      38643: inst = 32'd201344527;
      38644: inst = 32'd203423744;
      38645: inst = 32'd471859200;
      38646: inst = 32'd136314880;
      38647: inst = 32'd268468224;
      38648: inst = 32'd201344528;
      38649: inst = 32'd203423744;
      38650: inst = 32'd471859200;
      38651: inst = 32'd136314880;
      38652: inst = 32'd268468224;
      38653: inst = 32'd201344529;
      38654: inst = 32'd203483685;
      38655: inst = 32'd471859200;
      38656: inst = 32'd136314880;
      38657: inst = 32'd268468224;
      38658: inst = 32'd201344530;
      38659: inst = 32'd203483685;
      38660: inst = 32'd471859200;
      38661: inst = 32'd136314880;
      38662: inst = 32'd268468224;
      38663: inst = 32'd201344531;
      38664: inst = 32'd203483685;
      38665: inst = 32'd471859200;
      38666: inst = 32'd136314880;
      38667: inst = 32'd268468224;
      38668: inst = 32'd201344532;
      38669: inst = 32'd203423744;
      38670: inst = 32'd471859200;
      38671: inst = 32'd136314880;
      38672: inst = 32'd268468224;
      38673: inst = 32'd201344533;
      38674: inst = 32'd203423744;
      38675: inst = 32'd471859200;
      38676: inst = 32'd136314880;
      38677: inst = 32'd268468224;
      38678: inst = 32'd201344534;
      38679: inst = 32'd203423744;
      38680: inst = 32'd471859200;
      38681: inst = 32'd136314880;
      38682: inst = 32'd268468224;
      38683: inst = 32'd201344535;
      38684: inst = 32'd203423744;
      38685: inst = 32'd471859200;
      38686: inst = 32'd136314880;
      38687: inst = 32'd268468224;
      38688: inst = 32'd201344536;
      38689: inst = 32'd203423744;
      38690: inst = 32'd471859200;
      38691: inst = 32'd136314880;
      38692: inst = 32'd268468224;
      38693: inst = 32'd201344537;
      38694: inst = 32'd203423744;
      38695: inst = 32'd471859200;
      38696: inst = 32'd136314880;
      38697: inst = 32'd268468224;
      38698: inst = 32'd201344538;
      38699: inst = 32'd203483685;
      38700: inst = 32'd471859200;
      38701: inst = 32'd136314880;
      38702: inst = 32'd268468224;
      38703: inst = 32'd201344539;
      38704: inst = 32'd203483685;
      38705: inst = 32'd471859200;
      38706: inst = 32'd136314880;
      38707: inst = 32'd268468224;
      38708: inst = 32'd201344540;
      38709: inst = 32'd203483685;
      38710: inst = 32'd471859200;
      38711: inst = 32'd136314880;
      38712: inst = 32'd268468224;
      38713: inst = 32'd201344541;
      38714: inst = 32'd203483685;
      38715: inst = 32'd471859200;
      38716: inst = 32'd136314880;
      38717: inst = 32'd268468224;
      38718: inst = 32'd201344542;
      38719: inst = 32'd203423744;
      38720: inst = 32'd471859200;
      38721: inst = 32'd136314880;
      38722: inst = 32'd268468224;
      38723: inst = 32'd201344543;
      38724: inst = 32'd203423744;
      38725: inst = 32'd471859200;
      38726: inst = 32'd136314880;
      38727: inst = 32'd268468224;
      38728: inst = 32'd201344544;
      38729: inst = 32'd203423744;
      38730: inst = 32'd471859200;
      38731: inst = 32'd136314880;
      38732: inst = 32'd268468224;
      38733: inst = 32'd201344545;
      38734: inst = 32'd203483685;
      38735: inst = 32'd471859200;
      38736: inst = 32'd136314880;
      38737: inst = 32'd268468224;
      38738: inst = 32'd201344546;
      38739: inst = 32'd203483685;
      38740: inst = 32'd471859200;
      38741: inst = 32'd136314880;
      38742: inst = 32'd268468224;
      38743: inst = 32'd201344547;
      38744: inst = 32'd203483685;
      38745: inst = 32'd471859200;
      38746: inst = 32'd136314880;
      38747: inst = 32'd268468224;
      38748: inst = 32'd201344548;
      38749: inst = 32'd203483685;
      38750: inst = 32'd471859200;
      38751: inst = 32'd136314880;
      38752: inst = 32'd268468224;
      38753: inst = 32'd201344549;
      38754: inst = 32'd203483685;
      38755: inst = 32'd471859200;
      38756: inst = 32'd136314880;
      38757: inst = 32'd268468224;
      38758: inst = 32'd201344550;
      38759: inst = 32'd203483685;
      38760: inst = 32'd471859200;
      38761: inst = 32'd136314880;
      38762: inst = 32'd268468224;
      38763: inst = 32'd201344551;
      38764: inst = 32'd203423744;
      38765: inst = 32'd471859200;
      38766: inst = 32'd136314880;
      38767: inst = 32'd268468224;
      38768: inst = 32'd201344552;
      38769: inst = 32'd203423744;
      38770: inst = 32'd471859200;
      38771: inst = 32'd136314880;
      38772: inst = 32'd268468224;
      38773: inst = 32'd201344553;
      38774: inst = 32'd203423744;
      38775: inst = 32'd471859200;
      38776: inst = 32'd136314880;
      38777: inst = 32'd268468224;
      38778: inst = 32'd201344554;
      38779: inst = 32'd203483685;
      38780: inst = 32'd471859200;
      38781: inst = 32'd136314880;
      38782: inst = 32'd268468224;
      38783: inst = 32'd201344555;
      38784: inst = 32'd203483685;
      38785: inst = 32'd471859200;
      38786: inst = 32'd136314880;
      38787: inst = 32'd268468224;
      38788: inst = 32'd201344556;
      38789: inst = 32'd203483685;
      38790: inst = 32'd471859200;
      38791: inst = 32'd136314880;
      38792: inst = 32'd268468224;
      38793: inst = 32'd201344557;
      38794: inst = 32'd203483685;
      38795: inst = 32'd471859200;
      38796: inst = 32'd136314880;
      38797: inst = 32'd268468224;
      38798: inst = 32'd201344558;
      38799: inst = 32'd203483685;
      38800: inst = 32'd471859200;
      38801: inst = 32'd136314880;
      38802: inst = 32'd268468224;
      38803: inst = 32'd201344559;
      38804: inst = 32'd203483685;
      38805: inst = 32'd471859200;
      38806: inst = 32'd136314880;
      38807: inst = 32'd268468224;
      38808: inst = 32'd201344560;
      38809: inst = 32'd203483685;
      38810: inst = 32'd471859200;
      38811: inst = 32'd136314880;
      38812: inst = 32'd268468224;
      38813: inst = 32'd201344561;
      38814: inst = 32'd203483685;
      38815: inst = 32'd471859200;
      38816: inst = 32'd136314880;
      38817: inst = 32'd268468224;
      38818: inst = 32'd201344562;
      38819: inst = 32'd203483685;
      38820: inst = 32'd471859200;
      38821: inst = 32'd136314880;
      38822: inst = 32'd268468224;
      38823: inst = 32'd201344563;
      38824: inst = 32'd203483685;
      38825: inst = 32'd471859200;
      38826: inst = 32'd136314880;
      38827: inst = 32'd268468224;
      38828: inst = 32'd201344564;
      38829: inst = 32'd203483685;
      38830: inst = 32'd471859200;
      38831: inst = 32'd136314880;
      38832: inst = 32'd268468224;
      38833: inst = 32'd201344565;
      38834: inst = 32'd203423744;
      38835: inst = 32'd471859200;
      38836: inst = 32'd136314880;
      38837: inst = 32'd268468224;
      38838: inst = 32'd201344566;
      38839: inst = 32'd203423744;
      38840: inst = 32'd471859200;
      38841: inst = 32'd136314880;
      38842: inst = 32'd268468224;
      38843: inst = 32'd201344567;
      38844: inst = 32'd203423744;
      38845: inst = 32'd471859200;
      38846: inst = 32'd136314880;
      38847: inst = 32'd268468224;
      38848: inst = 32'd201344568;
      38849: inst = 32'd203423744;
      38850: inst = 32'd471859200;
      38851: inst = 32'd136314880;
      38852: inst = 32'd268468224;
      38853: inst = 32'd201344569;
      38854: inst = 32'd203423744;
      38855: inst = 32'd471859200;
      38856: inst = 32'd136314880;
      38857: inst = 32'd268468224;
      38858: inst = 32'd201344570;
      38859: inst = 32'd203423744;
      38860: inst = 32'd471859200;
      38861: inst = 32'd136314880;
      38862: inst = 32'd268468224;
      38863: inst = 32'd201344571;
      38864: inst = 32'd203423744;
      38865: inst = 32'd471859200;
      38866: inst = 32'd136314880;
      38867: inst = 32'd268468224;
      38868: inst = 32'd201344572;
      38869: inst = 32'd203423744;
      38870: inst = 32'd471859200;
      38871: inst = 32'd136314880;
      38872: inst = 32'd268468224;
      38873: inst = 32'd201344573;
      38874: inst = 32'd203423744;
      38875: inst = 32'd471859200;
      38876: inst = 32'd136314880;
      38877: inst = 32'd268468224;
      38878: inst = 32'd201344574;
      38879: inst = 32'd203423744;
      38880: inst = 32'd471859200;
      38881: inst = 32'd136314880;
      38882: inst = 32'd268468224;
      38883: inst = 32'd201344575;
      38884: inst = 32'd203423744;
      38885: inst = 32'd471859200;
      38886: inst = 32'd136314880;
      38887: inst = 32'd268468224;
      38888: inst = 32'd201344576;
      38889: inst = 32'd203423744;
      38890: inst = 32'd471859200;
      38891: inst = 32'd136314880;
      38892: inst = 32'd268468224;
      38893: inst = 32'd201344577;
      38894: inst = 32'd203423744;
      38895: inst = 32'd471859200;
      38896: inst = 32'd136314880;
      38897: inst = 32'd268468224;
      38898: inst = 32'd201344578;
      38899: inst = 32'd203423744;
      38900: inst = 32'd471859200;
      38901: inst = 32'd136314880;
      38902: inst = 32'd268468224;
      38903: inst = 32'd201344579;
      38904: inst = 32'd203423744;
      38905: inst = 32'd471859200;
      38906: inst = 32'd136314880;
      38907: inst = 32'd268468224;
      38908: inst = 32'd201344580;
      38909: inst = 32'd203423744;
      38910: inst = 32'd471859200;
      38911: inst = 32'd136314880;
      38912: inst = 32'd268468224;
      38913: inst = 32'd201344581;
      38914: inst = 32'd203423744;
      38915: inst = 32'd471859200;
      38916: inst = 32'd136314880;
      38917: inst = 32'd268468224;
      38918: inst = 32'd201344582;
      38919: inst = 32'd203423744;
      38920: inst = 32'd471859200;
      38921: inst = 32'd136314880;
      38922: inst = 32'd268468224;
      38923: inst = 32'd201344583;
      38924: inst = 32'd203423744;
      38925: inst = 32'd471859200;
      38926: inst = 32'd136314880;
      38927: inst = 32'd268468224;
      38928: inst = 32'd201344584;
      38929: inst = 32'd203423744;
      38930: inst = 32'd471859200;
      38931: inst = 32'd136314880;
      38932: inst = 32'd268468224;
      38933: inst = 32'd201344585;
      38934: inst = 32'd203423744;
      38935: inst = 32'd471859200;
      38936: inst = 32'd136314880;
      38937: inst = 32'd268468224;
      38938: inst = 32'd201344586;
      38939: inst = 32'd203423744;
      38940: inst = 32'd471859200;
      38941: inst = 32'd136314880;
      38942: inst = 32'd268468224;
      38943: inst = 32'd201344587;
      38944: inst = 32'd203423744;
      38945: inst = 32'd471859200;
      38946: inst = 32'd136314880;
      38947: inst = 32'd268468224;
      38948: inst = 32'd201344588;
      38949: inst = 32'd203423744;
      38950: inst = 32'd471859200;
      38951: inst = 32'd136314880;
      38952: inst = 32'd268468224;
      38953: inst = 32'd201344589;
      38954: inst = 32'd203483685;
      38955: inst = 32'd471859200;
      38956: inst = 32'd136314880;
      38957: inst = 32'd268468224;
      38958: inst = 32'd201344590;
      38959: inst = 32'd203483685;
      38960: inst = 32'd471859200;
      38961: inst = 32'd136314880;
      38962: inst = 32'd268468224;
      38963: inst = 32'd201344591;
      38964: inst = 32'd203483685;
      38965: inst = 32'd471859200;
      38966: inst = 32'd136314880;
      38967: inst = 32'd268468224;
      38968: inst = 32'd201344592;
      38969: inst = 32'd203483685;
      38970: inst = 32'd471859200;
      38971: inst = 32'd136314880;
      38972: inst = 32'd268468224;
      38973: inst = 32'd201344593;
      38974: inst = 32'd203483685;
      38975: inst = 32'd471859200;
      38976: inst = 32'd136314880;
      38977: inst = 32'd268468224;
      38978: inst = 32'd201344594;
      38979: inst = 32'd203483685;
      38980: inst = 32'd471859200;
      38981: inst = 32'd136314880;
      38982: inst = 32'd268468224;
      38983: inst = 32'd201344595;
      38984: inst = 32'd203483685;
      38985: inst = 32'd471859200;
      38986: inst = 32'd136314880;
      38987: inst = 32'd268468224;
      38988: inst = 32'd201344596;
      38989: inst = 32'd203483685;
      38990: inst = 32'd471859200;
      38991: inst = 32'd136314880;
      38992: inst = 32'd268468224;
      38993: inst = 32'd201344597;
      38994: inst = 32'd203423744;
      38995: inst = 32'd471859200;
      38996: inst = 32'd136314880;
      38997: inst = 32'd268468224;
      38998: inst = 32'd201344598;
      38999: inst = 32'd203423744;
      39000: inst = 32'd471859200;
      39001: inst = 32'd136314880;
      39002: inst = 32'd268468224;
      39003: inst = 32'd201344599;
      39004: inst = 32'd203423744;
      39005: inst = 32'd471859200;
      39006: inst = 32'd136314880;
      39007: inst = 32'd268468224;
      39008: inst = 32'd201344600;
      39009: inst = 32'd203483685;
      39010: inst = 32'd471859200;
      39011: inst = 32'd136314880;
      39012: inst = 32'd268468224;
      39013: inst = 32'd201344601;
      39014: inst = 32'd203483685;
      39015: inst = 32'd471859200;
      39016: inst = 32'd136314880;
      39017: inst = 32'd268468224;
      39018: inst = 32'd201344602;
      39019: inst = 32'd203483685;
      39020: inst = 32'd471859200;
      39021: inst = 32'd136314880;
      39022: inst = 32'd268468224;
      39023: inst = 32'd201344603;
      39024: inst = 32'd203483685;
      39025: inst = 32'd471859200;
      39026: inst = 32'd136314880;
      39027: inst = 32'd268468224;
      39028: inst = 32'd201344604;
      39029: inst = 32'd203483685;
      39030: inst = 32'd471859200;
      39031: inst = 32'd136314880;
      39032: inst = 32'd268468224;
      39033: inst = 32'd201344605;
      39034: inst = 32'd203483685;
      39035: inst = 32'd471859200;
      39036: inst = 32'd136314880;
      39037: inst = 32'd268468224;
      39038: inst = 32'd201344606;
      39039: inst = 32'd203483685;
      39040: inst = 32'd471859200;
      39041: inst = 32'd136314880;
      39042: inst = 32'd268468224;
      39043: inst = 32'd201344607;
      39044: inst = 32'd203483685;
      39045: inst = 32'd471859200;
      39046: inst = 32'd136314880;
      39047: inst = 32'd268468224;
      39048: inst = 32'd201344608;
      39049: inst = 32'd203483685;
      39050: inst = 32'd471859200;
      39051: inst = 32'd136314880;
      39052: inst = 32'd268468224;
      39053: inst = 32'd201344609;
      39054: inst = 32'd203423744;
      39055: inst = 32'd471859200;
      39056: inst = 32'd136314880;
      39057: inst = 32'd268468224;
      39058: inst = 32'd201344610;
      39059: inst = 32'd203423744;
      39060: inst = 32'd471859200;
      39061: inst = 32'd136314880;
      39062: inst = 32'd268468224;
      39063: inst = 32'd201344611;
      39064: inst = 32'd203423744;
      39065: inst = 32'd471859200;
      39066: inst = 32'd136314880;
      39067: inst = 32'd268468224;
      39068: inst = 32'd201344612;
      39069: inst = 32'd203423744;
      39070: inst = 32'd471859200;
      39071: inst = 32'd136314880;
      39072: inst = 32'd268468224;
      39073: inst = 32'd201344613;
      39074: inst = 32'd203423744;
      39075: inst = 32'd471859200;
      39076: inst = 32'd136314880;
      39077: inst = 32'd268468224;
      39078: inst = 32'd201344614;
      39079: inst = 32'd203423744;
      39080: inst = 32'd471859200;
      39081: inst = 32'd136314880;
      39082: inst = 32'd268468224;
      39083: inst = 32'd201344615;
      39084: inst = 32'd203483685;
      39085: inst = 32'd471859200;
      39086: inst = 32'd136314880;
      39087: inst = 32'd268468224;
      39088: inst = 32'd201344616;
      39089: inst = 32'd203483685;
      39090: inst = 32'd471859200;
      39091: inst = 32'd136314880;
      39092: inst = 32'd268468224;
      39093: inst = 32'd201344617;
      39094: inst = 32'd203483685;
      39095: inst = 32'd471859200;
      39096: inst = 32'd136314880;
      39097: inst = 32'd268468224;
      39098: inst = 32'd201344618;
      39099: inst = 32'd203483685;
      39100: inst = 32'd471859200;
      39101: inst = 32'd136314880;
      39102: inst = 32'd268468224;
      39103: inst = 32'd201344619;
      39104: inst = 32'd203483685;
      39105: inst = 32'd471859200;
      39106: inst = 32'd136314880;
      39107: inst = 32'd268468224;
      39108: inst = 32'd201344620;
      39109: inst = 32'd203423744;
      39110: inst = 32'd471859200;
      39111: inst = 32'd136314880;
      39112: inst = 32'd268468224;
      39113: inst = 32'd201344621;
      39114: inst = 32'd203423744;
      39115: inst = 32'd471859200;
      39116: inst = 32'd136314880;
      39117: inst = 32'd268468224;
      39118: inst = 32'd201344622;
      39119: inst = 32'd203423744;
      39120: inst = 32'd471859200;
      39121: inst = 32'd136314880;
      39122: inst = 32'd268468224;
      39123: inst = 32'd201344623;
      39124: inst = 32'd203423744;
      39125: inst = 32'd471859200;
      39126: inst = 32'd136314880;
      39127: inst = 32'd268468224;
      39128: inst = 32'd201344624;
      39129: inst = 32'd203423744;
      39130: inst = 32'd471859200;
      39131: inst = 32'd136314880;
      39132: inst = 32'd268468224;
      39133: inst = 32'd201344625;
      39134: inst = 32'd203483685;
      39135: inst = 32'd471859200;
      39136: inst = 32'd136314880;
      39137: inst = 32'd268468224;
      39138: inst = 32'd201344626;
      39139: inst = 32'd203483685;
      39140: inst = 32'd471859200;
      39141: inst = 32'd136314880;
      39142: inst = 32'd268468224;
      39143: inst = 32'd201344627;
      39144: inst = 32'd203483685;
      39145: inst = 32'd471859200;
      39146: inst = 32'd136314880;
      39147: inst = 32'd268468224;
      39148: inst = 32'd201344628;
      39149: inst = 32'd203423744;
      39150: inst = 32'd471859200;
      39151: inst = 32'd136314880;
      39152: inst = 32'd268468224;
      39153: inst = 32'd201344629;
      39154: inst = 32'd203423744;
      39155: inst = 32'd471859200;
      39156: inst = 32'd136314880;
      39157: inst = 32'd268468224;
      39158: inst = 32'd201344630;
      39159: inst = 32'd203423744;
      39160: inst = 32'd471859200;
      39161: inst = 32'd136314880;
      39162: inst = 32'd268468224;
      39163: inst = 32'd201344631;
      39164: inst = 32'd203423744;
      39165: inst = 32'd471859200;
      39166: inst = 32'd136314880;
      39167: inst = 32'd268468224;
      39168: inst = 32'd201344632;
      39169: inst = 32'd203423744;
      39170: inst = 32'd471859200;
      39171: inst = 32'd136314880;
      39172: inst = 32'd268468224;
      39173: inst = 32'd201344633;
      39174: inst = 32'd203423744;
      39175: inst = 32'd471859200;
      39176: inst = 32'd136314880;
      39177: inst = 32'd268468224;
      39178: inst = 32'd201344634;
      39179: inst = 32'd203483685;
      39180: inst = 32'd471859200;
      39181: inst = 32'd136314880;
      39182: inst = 32'd268468224;
      39183: inst = 32'd201344635;
      39184: inst = 32'd203483685;
      39185: inst = 32'd471859200;
      39186: inst = 32'd136314880;
      39187: inst = 32'd268468224;
      39188: inst = 32'd201344636;
      39189: inst = 32'd203483685;
      39190: inst = 32'd471859200;
      39191: inst = 32'd136314880;
      39192: inst = 32'd268468224;
      39193: inst = 32'd201344637;
      39194: inst = 32'd203483685;
      39195: inst = 32'd471859200;
      39196: inst = 32'd136314880;
      39197: inst = 32'd268468224;
      39198: inst = 32'd201344638;
      39199: inst = 32'd203423744;
      39200: inst = 32'd471859200;
      39201: inst = 32'd136314880;
      39202: inst = 32'd268468224;
      39203: inst = 32'd201344639;
      39204: inst = 32'd203423744;
      39205: inst = 32'd471859200;
      39206: inst = 32'd136314880;
      39207: inst = 32'd268468224;
      39208: inst = 32'd201344640;
      39209: inst = 32'd203423744;
      39210: inst = 32'd471859200;
      39211: inst = 32'd136314880;
      39212: inst = 32'd268468224;
      39213: inst = 32'd201344641;
      39214: inst = 32'd203483685;
      39215: inst = 32'd471859200;
      39216: inst = 32'd136314880;
      39217: inst = 32'd268468224;
      39218: inst = 32'd201344642;
      39219: inst = 32'd203483685;
      39220: inst = 32'd471859200;
      39221: inst = 32'd136314880;
      39222: inst = 32'd268468224;
      39223: inst = 32'd201344643;
      39224: inst = 32'd203483685;
      39225: inst = 32'd471859200;
      39226: inst = 32'd136314880;
      39227: inst = 32'd268468224;
      39228: inst = 32'd201344644;
      39229: inst = 32'd203483685;
      39230: inst = 32'd471859200;
      39231: inst = 32'd136314880;
      39232: inst = 32'd268468224;
      39233: inst = 32'd201344645;
      39234: inst = 32'd203483685;
      39235: inst = 32'd471859200;
      39236: inst = 32'd136314880;
      39237: inst = 32'd268468224;
      39238: inst = 32'd201344646;
      39239: inst = 32'd203423744;
      39240: inst = 32'd471859200;
      39241: inst = 32'd136314880;
      39242: inst = 32'd268468224;
      39243: inst = 32'd201344647;
      39244: inst = 32'd203423744;
      39245: inst = 32'd471859200;
      39246: inst = 32'd136314880;
      39247: inst = 32'd268468224;
      39248: inst = 32'd201344648;
      39249: inst = 32'd203423744;
      39250: inst = 32'd471859200;
      39251: inst = 32'd136314880;
      39252: inst = 32'd268468224;
      39253: inst = 32'd201344649;
      39254: inst = 32'd203423744;
      39255: inst = 32'd471859200;
      39256: inst = 32'd136314880;
      39257: inst = 32'd268468224;
      39258: inst = 32'd201344650;
      39259: inst = 32'd203483685;
      39260: inst = 32'd471859200;
      39261: inst = 32'd136314880;
      39262: inst = 32'd268468224;
      39263: inst = 32'd201344651;
      39264: inst = 32'd203483685;
      39265: inst = 32'd471859200;
      39266: inst = 32'd136314880;
      39267: inst = 32'd268468224;
      39268: inst = 32'd201344652;
      39269: inst = 32'd203483685;
      39270: inst = 32'd471859200;
      39271: inst = 32'd136314880;
      39272: inst = 32'd268468224;
      39273: inst = 32'd201344653;
      39274: inst = 32'd203483685;
      39275: inst = 32'd471859200;
      39276: inst = 32'd136314880;
      39277: inst = 32'd268468224;
      39278: inst = 32'd201344654;
      39279: inst = 32'd203483685;
      39280: inst = 32'd471859200;
      39281: inst = 32'd136314880;
      39282: inst = 32'd268468224;
      39283: inst = 32'd201344655;
      39284: inst = 32'd203483685;
      39285: inst = 32'd471859200;
      39286: inst = 32'd136314880;
      39287: inst = 32'd268468224;
      39288: inst = 32'd201344656;
      39289: inst = 32'd203483685;
      39290: inst = 32'd471859200;
      39291: inst = 32'd136314880;
      39292: inst = 32'd268468224;
      39293: inst = 32'd201344657;
      39294: inst = 32'd203483685;
      39295: inst = 32'd471859200;
      39296: inst = 32'd136314880;
      39297: inst = 32'd268468224;
      39298: inst = 32'd201344658;
      39299: inst = 32'd203483685;
      39300: inst = 32'd471859200;
      39301: inst = 32'd136314880;
      39302: inst = 32'd268468224;
      39303: inst = 32'd201344659;
      39304: inst = 32'd203483685;
      39305: inst = 32'd471859200;
      39306: inst = 32'd136314880;
      39307: inst = 32'd268468224;
      39308: inst = 32'd201344660;
      39309: inst = 32'd203483685;
      39310: inst = 32'd471859200;
      39311: inst = 32'd136314880;
      39312: inst = 32'd268468224;
      39313: inst = 32'd201344661;
      39314: inst = 32'd203483685;
      39315: inst = 32'd471859200;
      39316: inst = 32'd136314880;
      39317: inst = 32'd268468224;
      39318: inst = 32'd201344662;
      39319: inst = 32'd203423744;
      39320: inst = 32'd471859200;
      39321: inst = 32'd136314880;
      39322: inst = 32'd268468224;
      39323: inst = 32'd201344663;
      39324: inst = 32'd203423744;
      39325: inst = 32'd471859200;
      39326: inst = 32'd136314880;
      39327: inst = 32'd268468224;
      39328: inst = 32'd201344664;
      39329: inst = 32'd203423744;
      39330: inst = 32'd471859200;
      39331: inst = 32'd136314880;
      39332: inst = 32'd268468224;
      39333: inst = 32'd201344665;
      39334: inst = 32'd203423744;
      39335: inst = 32'd471859200;
      39336: inst = 32'd136314880;
      39337: inst = 32'd268468224;
      39338: inst = 32'd201344666;
      39339: inst = 32'd203423744;
      39340: inst = 32'd471859200;
      39341: inst = 32'd136314880;
      39342: inst = 32'd268468224;
      39343: inst = 32'd201344667;
      39344: inst = 32'd203423744;
      39345: inst = 32'd471859200;
      39346: inst = 32'd136314880;
      39347: inst = 32'd268468224;
      39348: inst = 32'd201344668;
      39349: inst = 32'd203423744;
      39350: inst = 32'd471859200;
      39351: inst = 32'd136314880;
      39352: inst = 32'd268468224;
      39353: inst = 32'd201344669;
      39354: inst = 32'd203423744;
      39355: inst = 32'd471859200;
      39356: inst = 32'd136314880;
      39357: inst = 32'd268468224;
      39358: inst = 32'd201344670;
      39359: inst = 32'd203423744;
      39360: inst = 32'd471859200;
      39361: inst = 32'd136314880;
      39362: inst = 32'd268468224;
      39363: inst = 32'd201344671;
      39364: inst = 32'd203423744;
      39365: inst = 32'd471859200;
      39366: inst = 32'd136314880;
      39367: inst = 32'd268468224;
      39368: inst = 32'd201344672;
      39369: inst = 32'd203423744;
      39370: inst = 32'd471859200;
      39371: inst = 32'd136314880;
      39372: inst = 32'd268468224;
      39373: inst = 32'd201344673;
      39374: inst = 32'd203423744;
      39375: inst = 32'd471859200;
      39376: inst = 32'd136314880;
      39377: inst = 32'd268468224;
      39378: inst = 32'd201344674;
      39379: inst = 32'd203423744;
      39380: inst = 32'd471859200;
      39381: inst = 32'd136314880;
      39382: inst = 32'd268468224;
      39383: inst = 32'd201344675;
      39384: inst = 32'd203423744;
      39385: inst = 32'd471859200;
      39386: inst = 32'd136314880;
      39387: inst = 32'd268468224;
      39388: inst = 32'd201344676;
      39389: inst = 32'd203423744;
      39390: inst = 32'd471859200;
      39391: inst = 32'd136314880;
      39392: inst = 32'd268468224;
      39393: inst = 32'd201344677;
      39394: inst = 32'd203423744;
      39395: inst = 32'd471859200;
      39396: inst = 32'd136314880;
      39397: inst = 32'd268468224;
      39398: inst = 32'd201344678;
      39399: inst = 32'd203423744;
      39400: inst = 32'd471859200;
      39401: inst = 32'd136314880;
      39402: inst = 32'd268468224;
      39403: inst = 32'd201344679;
      39404: inst = 32'd203423744;
      39405: inst = 32'd471859200;
      39406: inst = 32'd136314880;
      39407: inst = 32'd268468224;
      39408: inst = 32'd201344680;
      39409: inst = 32'd203423744;
      39410: inst = 32'd471859200;
      39411: inst = 32'd136314880;
      39412: inst = 32'd268468224;
      39413: inst = 32'd201344681;
      39414: inst = 32'd203423744;
      39415: inst = 32'd471859200;
      39416: inst = 32'd136314880;
      39417: inst = 32'd268468224;
      39418: inst = 32'd201344682;
      39419: inst = 32'd203423744;
      39420: inst = 32'd471859200;
      39421: inst = 32'd136314880;
      39422: inst = 32'd268468224;
      39423: inst = 32'd201344683;
      39424: inst = 32'd203423744;
      39425: inst = 32'd471859200;
      39426: inst = 32'd136314880;
      39427: inst = 32'd268468224;
      39428: inst = 32'd201344684;
      39429: inst = 32'd203423744;
      39430: inst = 32'd471859200;
      39431: inst = 32'd136314880;
      39432: inst = 32'd268468224;
      39433: inst = 32'd201344685;
      39434: inst = 32'd203483685;
      39435: inst = 32'd471859200;
      39436: inst = 32'd136314880;
      39437: inst = 32'd268468224;
      39438: inst = 32'd201344686;
      39439: inst = 32'd203483685;
      39440: inst = 32'd471859200;
      39441: inst = 32'd136314880;
      39442: inst = 32'd268468224;
      39443: inst = 32'd201344687;
      39444: inst = 32'd203483685;
      39445: inst = 32'd471859200;
      39446: inst = 32'd136314880;
      39447: inst = 32'd268468224;
      39448: inst = 32'd201344688;
      39449: inst = 32'd203483685;
      39450: inst = 32'd471859200;
      39451: inst = 32'd136314880;
      39452: inst = 32'd268468224;
      39453: inst = 32'd201344689;
      39454: inst = 32'd203483685;
      39455: inst = 32'd471859200;
      39456: inst = 32'd136314880;
      39457: inst = 32'd268468224;
      39458: inst = 32'd201344690;
      39459: inst = 32'd203483685;
      39460: inst = 32'd471859200;
      39461: inst = 32'd136314880;
      39462: inst = 32'd268468224;
      39463: inst = 32'd201344691;
      39464: inst = 32'd203483685;
      39465: inst = 32'd471859200;
      39466: inst = 32'd136314880;
      39467: inst = 32'd268468224;
      39468: inst = 32'd201344692;
      39469: inst = 32'd203483685;
      39470: inst = 32'd471859200;
      39471: inst = 32'd136314880;
      39472: inst = 32'd268468224;
      39473: inst = 32'd201344693;
      39474: inst = 32'd203423744;
      39475: inst = 32'd471859200;
      39476: inst = 32'd136314880;
      39477: inst = 32'd268468224;
      39478: inst = 32'd201344694;
      39479: inst = 32'd203423744;
      39480: inst = 32'd471859200;
      39481: inst = 32'd136314880;
      39482: inst = 32'd268468224;
      39483: inst = 32'd201344695;
      39484: inst = 32'd203423744;
      39485: inst = 32'd471859200;
      39486: inst = 32'd136314880;
      39487: inst = 32'd268468224;
      39488: inst = 32'd201344696;
      39489: inst = 32'd203483685;
      39490: inst = 32'd471859200;
      39491: inst = 32'd136314880;
      39492: inst = 32'd268468224;
      39493: inst = 32'd201344697;
      39494: inst = 32'd203483685;
      39495: inst = 32'd471859200;
      39496: inst = 32'd136314880;
      39497: inst = 32'd268468224;
      39498: inst = 32'd201344698;
      39499: inst = 32'd203483685;
      39500: inst = 32'd471859200;
      39501: inst = 32'd136314880;
      39502: inst = 32'd268468224;
      39503: inst = 32'd201344699;
      39504: inst = 32'd203483685;
      39505: inst = 32'd471859200;
      39506: inst = 32'd136314880;
      39507: inst = 32'd268468224;
      39508: inst = 32'd201344700;
      39509: inst = 32'd203483685;
      39510: inst = 32'd471859200;
      39511: inst = 32'd136314880;
      39512: inst = 32'd268468224;
      39513: inst = 32'd201344701;
      39514: inst = 32'd203483685;
      39515: inst = 32'd471859200;
      39516: inst = 32'd136314880;
      39517: inst = 32'd268468224;
      39518: inst = 32'd201344702;
      39519: inst = 32'd203483685;
      39520: inst = 32'd471859200;
      39521: inst = 32'd136314880;
      39522: inst = 32'd268468224;
      39523: inst = 32'd201344703;
      39524: inst = 32'd203483685;
      39525: inst = 32'd471859200;
      39526: inst = 32'd136314880;
      39527: inst = 32'd268468224;
      39528: inst = 32'd201344704;
      39529: inst = 32'd203483685;
      39530: inst = 32'd471859200;
      39531: inst = 32'd136314880;
      39532: inst = 32'd268468224;
      39533: inst = 32'd201344705;
      39534: inst = 32'd203423744;
      39535: inst = 32'd471859200;
      39536: inst = 32'd136314880;
      39537: inst = 32'd268468224;
      39538: inst = 32'd201344706;
      39539: inst = 32'd203423744;
      39540: inst = 32'd471859200;
      39541: inst = 32'd136314880;
      39542: inst = 32'd268468224;
      39543: inst = 32'd201344707;
      39544: inst = 32'd203423744;
      39545: inst = 32'd471859200;
      39546: inst = 32'd136314880;
      39547: inst = 32'd268468224;
      39548: inst = 32'd201344708;
      39549: inst = 32'd203423744;
      39550: inst = 32'd471859200;
      39551: inst = 32'd136314880;
      39552: inst = 32'd268468224;
      39553: inst = 32'd201344709;
      39554: inst = 32'd203423744;
      39555: inst = 32'd471859200;
      39556: inst = 32'd136314880;
      39557: inst = 32'd268468224;
      39558: inst = 32'd201344710;
      39559: inst = 32'd203423744;
      39560: inst = 32'd471859200;
      39561: inst = 32'd136314880;
      39562: inst = 32'd268468224;
      39563: inst = 32'd201344711;
      39564: inst = 32'd203483685;
      39565: inst = 32'd471859200;
      39566: inst = 32'd136314880;
      39567: inst = 32'd268468224;
      39568: inst = 32'd201344712;
      39569: inst = 32'd203483685;
      39570: inst = 32'd471859200;
      39571: inst = 32'd136314880;
      39572: inst = 32'd268468224;
      39573: inst = 32'd201344713;
      39574: inst = 32'd203423744;
      39575: inst = 32'd471859200;
      39576: inst = 32'd136314880;
      39577: inst = 32'd268468224;
      39578: inst = 32'd201344714;
      39579: inst = 32'd203423744;
      39580: inst = 32'd471859200;
      39581: inst = 32'd136314880;
      39582: inst = 32'd268468224;
      39583: inst = 32'd201344715;
      39584: inst = 32'd203423744;
      39585: inst = 32'd471859200;
      39586: inst = 32'd136314880;
      39587: inst = 32'd268468224;
      39588: inst = 32'd201344716;
      39589: inst = 32'd203423744;
      39590: inst = 32'd471859200;
      39591: inst = 32'd136314880;
      39592: inst = 32'd268468224;
      39593: inst = 32'd201344717;
      39594: inst = 32'd203423744;
      39595: inst = 32'd471859200;
      39596: inst = 32'd136314880;
      39597: inst = 32'd268468224;
      39598: inst = 32'd201344718;
      39599: inst = 32'd203423744;
      39600: inst = 32'd471859200;
      39601: inst = 32'd136314880;
      39602: inst = 32'd268468224;
      39603: inst = 32'd201344719;
      39604: inst = 32'd203423744;
      39605: inst = 32'd471859200;
      39606: inst = 32'd136314880;
      39607: inst = 32'd268468224;
      39608: inst = 32'd201344720;
      39609: inst = 32'd203423744;
      39610: inst = 32'd471859200;
      39611: inst = 32'd136314880;
      39612: inst = 32'd268468224;
      39613: inst = 32'd201344721;
      39614: inst = 32'd203483685;
      39615: inst = 32'd471859200;
      39616: inst = 32'd136314880;
      39617: inst = 32'd268468224;
      39618: inst = 32'd201344722;
      39619: inst = 32'd203483685;
      39620: inst = 32'd471859200;
      39621: inst = 32'd136314880;
      39622: inst = 32'd268468224;
      39623: inst = 32'd201344723;
      39624: inst = 32'd203483685;
      39625: inst = 32'd471859200;
      39626: inst = 32'd136314880;
      39627: inst = 32'd268468224;
      39628: inst = 32'd201344724;
      39629: inst = 32'd203483685;
      39630: inst = 32'd471859200;
      39631: inst = 32'd136314880;
      39632: inst = 32'd268468224;
      39633: inst = 32'd201344725;
      39634: inst = 32'd203483685;
      39635: inst = 32'd471859200;
      39636: inst = 32'd136314880;
      39637: inst = 32'd268468224;
      39638: inst = 32'd201344726;
      39639: inst = 32'd203483685;
      39640: inst = 32'd471859200;
      39641: inst = 32'd136314880;
      39642: inst = 32'd268468224;
      39643: inst = 32'd201344727;
      39644: inst = 32'd203483685;
      39645: inst = 32'd471859200;
      39646: inst = 32'd136314880;
      39647: inst = 32'd268468224;
      39648: inst = 32'd201344728;
      39649: inst = 32'd203483685;
      39650: inst = 32'd471859200;
      39651: inst = 32'd136314880;
      39652: inst = 32'd268468224;
      39653: inst = 32'd201344729;
      39654: inst = 32'd203423744;
      39655: inst = 32'd471859200;
      39656: inst = 32'd136314880;
      39657: inst = 32'd268468224;
      39658: inst = 32'd201344730;
      39659: inst = 32'd203483685;
      39660: inst = 32'd471859200;
      39661: inst = 32'd136314880;
      39662: inst = 32'd268468224;
      39663: inst = 32'd201344731;
      39664: inst = 32'd203483685;
      39665: inst = 32'd471859200;
      39666: inst = 32'd136314880;
      39667: inst = 32'd268468224;
      39668: inst = 32'd201344732;
      39669: inst = 32'd203483685;
      39670: inst = 32'd471859200;
      39671: inst = 32'd136314880;
      39672: inst = 32'd268468224;
      39673: inst = 32'd201344733;
      39674: inst = 32'd203483685;
      39675: inst = 32'd471859200;
      39676: inst = 32'd136314880;
      39677: inst = 32'd268468224;
      39678: inst = 32'd201344734;
      39679: inst = 32'd203423744;
      39680: inst = 32'd471859200;
      39681: inst = 32'd136314880;
      39682: inst = 32'd268468224;
      39683: inst = 32'd201344735;
      39684: inst = 32'd203423744;
      39685: inst = 32'd471859200;
      39686: inst = 32'd136314880;
      39687: inst = 32'd268468224;
      39688: inst = 32'd201344736;
      39689: inst = 32'd203423744;
      39690: inst = 32'd471859200;
      39691: inst = 32'd136314880;
      39692: inst = 32'd268468224;
      39693: inst = 32'd201344737;
      39694: inst = 32'd203483685;
      39695: inst = 32'd471859200;
      39696: inst = 32'd136314880;
      39697: inst = 32'd268468224;
      39698: inst = 32'd201344738;
      39699: inst = 32'd203423744;
      39700: inst = 32'd471859200;
      39701: inst = 32'd136314880;
      39702: inst = 32'd268468224;
      39703: inst = 32'd201344739;
      39704: inst = 32'd203423744;
      39705: inst = 32'd471859200;
      39706: inst = 32'd136314880;
      39707: inst = 32'd268468224;
      39708: inst = 32'd201344740;
      39709: inst = 32'd203423744;
      39710: inst = 32'd471859200;
      39711: inst = 32'd136314880;
      39712: inst = 32'd268468224;
      39713: inst = 32'd201344741;
      39714: inst = 32'd203423744;
      39715: inst = 32'd471859200;
      39716: inst = 32'd136314880;
      39717: inst = 32'd268468224;
      39718: inst = 32'd201344742;
      39719: inst = 32'd203423744;
      39720: inst = 32'd471859200;
      39721: inst = 32'd136314880;
      39722: inst = 32'd268468224;
      39723: inst = 32'd201344743;
      39724: inst = 32'd203423744;
      39725: inst = 32'd471859200;
      39726: inst = 32'd136314880;
      39727: inst = 32'd268468224;
      39728: inst = 32'd201344744;
      39729: inst = 32'd203423744;
      39730: inst = 32'd471859200;
      39731: inst = 32'd136314880;
      39732: inst = 32'd268468224;
      39733: inst = 32'd201344745;
      39734: inst = 32'd203423744;
      39735: inst = 32'd471859200;
      39736: inst = 32'd136314880;
      39737: inst = 32'd268468224;
      39738: inst = 32'd201344746;
      39739: inst = 32'd203483685;
      39740: inst = 32'd471859200;
      39741: inst = 32'd136314880;
      39742: inst = 32'd268468224;
      39743: inst = 32'd201344747;
      39744: inst = 32'd203483685;
      39745: inst = 32'd471859200;
      39746: inst = 32'd136314880;
      39747: inst = 32'd268468224;
      39748: inst = 32'd201344748;
      39749: inst = 32'd203483685;
      39750: inst = 32'd471859200;
      39751: inst = 32'd136314880;
      39752: inst = 32'd268468224;
      39753: inst = 32'd201344749;
      39754: inst = 32'd203483685;
      39755: inst = 32'd471859200;
      39756: inst = 32'd136314880;
      39757: inst = 32'd268468224;
      39758: inst = 32'd201344750;
      39759: inst = 32'd203483685;
      39760: inst = 32'd471859200;
      39761: inst = 32'd136314880;
      39762: inst = 32'd268468224;
      39763: inst = 32'd201344751;
      39764: inst = 32'd203483685;
      39765: inst = 32'd471859200;
      39766: inst = 32'd136314880;
      39767: inst = 32'd268468224;
      39768: inst = 32'd201344752;
      39769: inst = 32'd203483685;
      39770: inst = 32'd471859200;
      39771: inst = 32'd136314880;
      39772: inst = 32'd268468224;
      39773: inst = 32'd201344753;
      39774: inst = 32'd203483685;
      39775: inst = 32'd471859200;
      39776: inst = 32'd136314880;
      39777: inst = 32'd268468224;
      39778: inst = 32'd201344754;
      39779: inst = 32'd203483685;
      39780: inst = 32'd471859200;
      39781: inst = 32'd136314880;
      39782: inst = 32'd268468224;
      39783: inst = 32'd201344755;
      39784: inst = 32'd203483685;
      39785: inst = 32'd471859200;
      39786: inst = 32'd136314880;
      39787: inst = 32'd268468224;
      39788: inst = 32'd201344756;
      39789: inst = 32'd203483685;
      39790: inst = 32'd471859200;
      39791: inst = 32'd136314880;
      39792: inst = 32'd268468224;
      39793: inst = 32'd201344757;
      39794: inst = 32'd203483685;
      39795: inst = 32'd471859200;
      39796: inst = 32'd136314880;
      39797: inst = 32'd268468224;
      39798: inst = 32'd201344758;
      39799: inst = 32'd203423744;
      39800: inst = 32'd471859200;
      39801: inst = 32'd136314880;
      39802: inst = 32'd268468224;
      39803: inst = 32'd201344759;
      39804: inst = 32'd203423744;
      39805: inst = 32'd471859200;
      39806: inst = 32'd136314880;
      39807: inst = 32'd268468224;
      39808: inst = 32'd201344760;
      39809: inst = 32'd203423744;
      39810: inst = 32'd471859200;
      39811: inst = 32'd136314880;
      39812: inst = 32'd268468224;
      39813: inst = 32'd201344761;
      39814: inst = 32'd203423744;
      39815: inst = 32'd471859200;
      39816: inst = 32'd136314880;
      39817: inst = 32'd268468224;
      39818: inst = 32'd201344762;
      39819: inst = 32'd203423744;
      39820: inst = 32'd471859200;
      39821: inst = 32'd136314880;
      39822: inst = 32'd268468224;
      39823: inst = 32'd201344763;
      39824: inst = 32'd203423744;
      39825: inst = 32'd471859200;
      39826: inst = 32'd136314880;
      39827: inst = 32'd268468224;
      39828: inst = 32'd201344764;
      39829: inst = 32'd203423744;
      39830: inst = 32'd471859200;
      39831: inst = 32'd136314880;
      39832: inst = 32'd268468224;
      39833: inst = 32'd201344765;
      39834: inst = 32'd203423744;
      39835: inst = 32'd471859200;
      39836: inst = 32'd136314880;
      39837: inst = 32'd268468224;
      39838: inst = 32'd201344766;
      39839: inst = 32'd203423744;
      39840: inst = 32'd471859200;
      39841: inst = 32'd136314880;
      39842: inst = 32'd268468224;
      39843: inst = 32'd201344767;
      39844: inst = 32'd203423744;
      39845: inst = 32'd471859200;
      39846: inst = 32'd136314880;
      39847: inst = 32'd268468224;
      39848: inst = 32'd201344768;
      39849: inst = 32'd203423744;
      39850: inst = 32'd471859200;
      39851: inst = 32'd136314880;
      39852: inst = 32'd268468224;
      39853: inst = 32'd201344769;
      39854: inst = 32'd203423744;
      39855: inst = 32'd471859200;
      39856: inst = 32'd136314880;
      39857: inst = 32'd268468224;
      39858: inst = 32'd201344770;
      39859: inst = 32'd203423744;
      39860: inst = 32'd471859200;
      39861: inst = 32'd136314880;
      39862: inst = 32'd268468224;
      39863: inst = 32'd201344771;
      39864: inst = 32'd203423744;
      39865: inst = 32'd471859200;
      39866: inst = 32'd136314880;
      39867: inst = 32'd268468224;
      39868: inst = 32'd201344772;
      39869: inst = 32'd203423744;
      39870: inst = 32'd471859200;
      39871: inst = 32'd136314880;
      39872: inst = 32'd268468224;
      39873: inst = 32'd201344773;
      39874: inst = 32'd203423744;
      39875: inst = 32'd471859200;
      39876: inst = 32'd136314880;
      39877: inst = 32'd268468224;
      39878: inst = 32'd201344774;
      39879: inst = 32'd203423744;
      39880: inst = 32'd471859200;
      39881: inst = 32'd136314880;
      39882: inst = 32'd268468224;
      39883: inst = 32'd201344775;
      39884: inst = 32'd203423744;
      39885: inst = 32'd471859200;
      39886: inst = 32'd136314880;
      39887: inst = 32'd268468224;
      39888: inst = 32'd201344776;
      39889: inst = 32'd203423744;
      39890: inst = 32'd471859200;
      39891: inst = 32'd136314880;
      39892: inst = 32'd268468224;
      39893: inst = 32'd201344777;
      39894: inst = 32'd203423744;
      39895: inst = 32'd471859200;
      39896: inst = 32'd136314880;
      39897: inst = 32'd268468224;
      39898: inst = 32'd201344778;
      39899: inst = 32'd203423744;
      39900: inst = 32'd471859200;
      39901: inst = 32'd136314880;
      39902: inst = 32'd268468224;
      39903: inst = 32'd201344779;
      39904: inst = 32'd203423744;
      39905: inst = 32'd471859200;
      39906: inst = 32'd136314880;
      39907: inst = 32'd268468224;
      39908: inst = 32'd201344780;
      39909: inst = 32'd203423744;
      39910: inst = 32'd471859200;
      39911: inst = 32'd136314880;
      39912: inst = 32'd268468224;
      39913: inst = 32'd201344781;
      39914: inst = 32'd203483685;
      39915: inst = 32'd471859200;
      39916: inst = 32'd136314880;
      39917: inst = 32'd268468224;
      39918: inst = 32'd201344782;
      39919: inst = 32'd203483685;
      39920: inst = 32'd471859200;
      39921: inst = 32'd136314880;
      39922: inst = 32'd268468224;
      39923: inst = 32'd201344783;
      39924: inst = 32'd203483685;
      39925: inst = 32'd471859200;
      39926: inst = 32'd136314880;
      39927: inst = 32'd268468224;
      39928: inst = 32'd201344784;
      39929: inst = 32'd203483685;
      39930: inst = 32'd471859200;
      39931: inst = 32'd136314880;
      39932: inst = 32'd268468224;
      39933: inst = 32'd201344785;
      39934: inst = 32'd203483685;
      39935: inst = 32'd471859200;
      39936: inst = 32'd136314880;
      39937: inst = 32'd268468224;
      39938: inst = 32'd201344786;
      39939: inst = 32'd203483685;
      39940: inst = 32'd471859200;
      39941: inst = 32'd136314880;
      39942: inst = 32'd268468224;
      39943: inst = 32'd201344787;
      39944: inst = 32'd203483685;
      39945: inst = 32'd471859200;
      39946: inst = 32'd136314880;
      39947: inst = 32'd268468224;
      39948: inst = 32'd201344788;
      39949: inst = 32'd203483685;
      39950: inst = 32'd471859200;
      39951: inst = 32'd136314880;
      39952: inst = 32'd268468224;
      39953: inst = 32'd201344789;
      39954: inst = 32'd203483685;
      39955: inst = 32'd471859200;
      39956: inst = 32'd136314880;
      39957: inst = 32'd268468224;
      39958: inst = 32'd201344790;
      39959: inst = 32'd203483685;
      39960: inst = 32'd471859200;
      39961: inst = 32'd136314880;
      39962: inst = 32'd268468224;
      39963: inst = 32'd201344791;
      39964: inst = 32'd203483685;
      39965: inst = 32'd471859200;
      39966: inst = 32'd136314880;
      39967: inst = 32'd268468224;
      39968: inst = 32'd201344792;
      39969: inst = 32'd203483685;
      39970: inst = 32'd471859200;
      39971: inst = 32'd136314880;
      39972: inst = 32'd268468224;
      39973: inst = 32'd201344793;
      39974: inst = 32'd203483685;
      39975: inst = 32'd471859200;
      39976: inst = 32'd136314880;
      39977: inst = 32'd268468224;
      39978: inst = 32'd201344794;
      39979: inst = 32'd203483685;
      39980: inst = 32'd471859200;
      39981: inst = 32'd136314880;
      39982: inst = 32'd268468224;
      39983: inst = 32'd201344795;
      39984: inst = 32'd203483685;
      39985: inst = 32'd471859200;
      39986: inst = 32'd136314880;
      39987: inst = 32'd268468224;
      39988: inst = 32'd201344796;
      39989: inst = 32'd203483685;
      39990: inst = 32'd471859200;
      39991: inst = 32'd136314880;
      39992: inst = 32'd268468224;
      39993: inst = 32'd201344797;
      39994: inst = 32'd203483685;
      39995: inst = 32'd471859200;
      39996: inst = 32'd136314880;
      39997: inst = 32'd268468224;
      39998: inst = 32'd201344798;
      39999: inst = 32'd203483685;
      40000: inst = 32'd471859200;
      40001: inst = 32'd136314880;
      40002: inst = 32'd268468224;
      40003: inst = 32'd201344799;
      40004: inst = 32'd203483685;
      40005: inst = 32'd471859200;
      40006: inst = 32'd136314880;
      40007: inst = 32'd268468224;
      40008: inst = 32'd201344800;
      40009: inst = 32'd203483685;
      40010: inst = 32'd471859200;
      40011: inst = 32'd136314880;
      40012: inst = 32'd268468224;
      40013: inst = 32'd201344801;
      40014: inst = 32'd203483685;
      40015: inst = 32'd471859200;
      40016: inst = 32'd136314880;
      40017: inst = 32'd268468224;
      40018: inst = 32'd201344802;
      40019: inst = 32'd203483685;
      40020: inst = 32'd471859200;
      40021: inst = 32'd136314880;
      40022: inst = 32'd268468224;
      40023: inst = 32'd201344803;
      40024: inst = 32'd203483685;
      40025: inst = 32'd471859200;
      40026: inst = 32'd136314880;
      40027: inst = 32'd268468224;
      40028: inst = 32'd201344804;
      40029: inst = 32'd203423744;
      40030: inst = 32'd471859200;
      40031: inst = 32'd136314880;
      40032: inst = 32'd268468224;
      40033: inst = 32'd201344805;
      40034: inst = 32'd203483685;
      40035: inst = 32'd471859200;
      40036: inst = 32'd136314880;
      40037: inst = 32'd268468224;
      40038: inst = 32'd201344806;
      40039: inst = 32'd203483685;
      40040: inst = 32'd471859200;
      40041: inst = 32'd136314880;
      40042: inst = 32'd268468224;
      40043: inst = 32'd201344807;
      40044: inst = 32'd203483685;
      40045: inst = 32'd471859200;
      40046: inst = 32'd136314880;
      40047: inst = 32'd268468224;
      40048: inst = 32'd201344808;
      40049: inst = 32'd203483685;
      40050: inst = 32'd471859200;
      40051: inst = 32'd136314880;
      40052: inst = 32'd268468224;
      40053: inst = 32'd201344809;
      40054: inst = 32'd203483685;
      40055: inst = 32'd471859200;
      40056: inst = 32'd136314880;
      40057: inst = 32'd268468224;
      40058: inst = 32'd201344810;
      40059: inst = 32'd203483685;
      40060: inst = 32'd471859200;
      40061: inst = 32'd136314880;
      40062: inst = 32'd268468224;
      40063: inst = 32'd201344811;
      40064: inst = 32'd203483685;
      40065: inst = 32'd471859200;
      40066: inst = 32'd136314880;
      40067: inst = 32'd268468224;
      40068: inst = 32'd201344812;
      40069: inst = 32'd203483685;
      40070: inst = 32'd471859200;
      40071: inst = 32'd136314880;
      40072: inst = 32'd268468224;
      40073: inst = 32'd201344813;
      40074: inst = 32'd203483685;
      40075: inst = 32'd471859200;
      40076: inst = 32'd136314880;
      40077: inst = 32'd268468224;
      40078: inst = 32'd201344814;
      40079: inst = 32'd203483685;
      40080: inst = 32'd471859200;
      40081: inst = 32'd136314880;
      40082: inst = 32'd268468224;
      40083: inst = 32'd201344815;
      40084: inst = 32'd203483685;
      40085: inst = 32'd471859200;
      40086: inst = 32'd136314880;
      40087: inst = 32'd268468224;
      40088: inst = 32'd201344816;
      40089: inst = 32'd203483685;
      40090: inst = 32'd471859200;
      40091: inst = 32'd136314880;
      40092: inst = 32'd268468224;
      40093: inst = 32'd201344817;
      40094: inst = 32'd203483685;
      40095: inst = 32'd471859200;
      40096: inst = 32'd136314880;
      40097: inst = 32'd268468224;
      40098: inst = 32'd201344818;
      40099: inst = 32'd203483685;
      40100: inst = 32'd471859200;
      40101: inst = 32'd136314880;
      40102: inst = 32'd268468224;
      40103: inst = 32'd201344819;
      40104: inst = 32'd203483685;
      40105: inst = 32'd471859200;
      40106: inst = 32'd136314880;
      40107: inst = 32'd268468224;
      40108: inst = 32'd201344820;
      40109: inst = 32'd203483685;
      40110: inst = 32'd471859200;
      40111: inst = 32'd136314880;
      40112: inst = 32'd268468224;
      40113: inst = 32'd201344821;
      40114: inst = 32'd203483685;
      40115: inst = 32'd471859200;
      40116: inst = 32'd136314880;
      40117: inst = 32'd268468224;
      40118: inst = 32'd201344822;
      40119: inst = 32'd203483685;
      40120: inst = 32'd471859200;
      40121: inst = 32'd136314880;
      40122: inst = 32'd268468224;
      40123: inst = 32'd201344823;
      40124: inst = 32'd203483685;
      40125: inst = 32'd471859200;
      40126: inst = 32'd136314880;
      40127: inst = 32'd268468224;
      40128: inst = 32'd201344824;
      40129: inst = 32'd203483685;
      40130: inst = 32'd471859200;
      40131: inst = 32'd136314880;
      40132: inst = 32'd268468224;
      40133: inst = 32'd201344825;
      40134: inst = 32'd203483685;
      40135: inst = 32'd471859200;
      40136: inst = 32'd136314880;
      40137: inst = 32'd268468224;
      40138: inst = 32'd201344826;
      40139: inst = 32'd203483685;
      40140: inst = 32'd471859200;
      40141: inst = 32'd136314880;
      40142: inst = 32'd268468224;
      40143: inst = 32'd201344827;
      40144: inst = 32'd203483685;
      40145: inst = 32'd471859200;
      40146: inst = 32'd136314880;
      40147: inst = 32'd268468224;
      40148: inst = 32'd201344828;
      40149: inst = 32'd203483685;
      40150: inst = 32'd471859200;
      40151: inst = 32'd136314880;
      40152: inst = 32'd268468224;
      40153: inst = 32'd201344829;
      40154: inst = 32'd203483685;
      40155: inst = 32'd471859200;
      40156: inst = 32'd136314880;
      40157: inst = 32'd268468224;
      40158: inst = 32'd201344830;
      40159: inst = 32'd203423744;
      40160: inst = 32'd471859200;
      40161: inst = 32'd136314880;
      40162: inst = 32'd268468224;
      40163: inst = 32'd201344831;
      40164: inst = 32'd203483685;
      40165: inst = 32'd471859200;
      40166: inst = 32'd136314880;
      40167: inst = 32'd268468224;
      40168: inst = 32'd201344832;
      40169: inst = 32'd203483685;
      40170: inst = 32'd471859200;
      40171: inst = 32'd136314880;
      40172: inst = 32'd268468224;
      40173: inst = 32'd201344833;
      40174: inst = 32'd203483685;
      40175: inst = 32'd471859200;
      40176: inst = 32'd136314880;
      40177: inst = 32'd268468224;
      40178: inst = 32'd201344834;
      40179: inst = 32'd203483685;
      40180: inst = 32'd471859200;
      40181: inst = 32'd136314880;
      40182: inst = 32'd268468224;
      40183: inst = 32'd201344835;
      40184: inst = 32'd203483685;
      40185: inst = 32'd471859200;
      40186: inst = 32'd136314880;
      40187: inst = 32'd268468224;
      40188: inst = 32'd201344836;
      40189: inst = 32'd203483685;
      40190: inst = 32'd471859200;
      40191: inst = 32'd136314880;
      40192: inst = 32'd268468224;
      40193: inst = 32'd201344837;
      40194: inst = 32'd203483685;
      40195: inst = 32'd471859200;
      40196: inst = 32'd136314880;
      40197: inst = 32'd268468224;
      40198: inst = 32'd201344838;
      40199: inst = 32'd203483685;
      40200: inst = 32'd471859200;
      40201: inst = 32'd136314880;
      40202: inst = 32'd268468224;
      40203: inst = 32'd201344839;
      40204: inst = 32'd203483685;
      40205: inst = 32'd471859200;
      40206: inst = 32'd136314880;
      40207: inst = 32'd268468224;
      40208: inst = 32'd201344840;
      40209: inst = 32'd203483685;
      40210: inst = 32'd471859200;
      40211: inst = 32'd136314880;
      40212: inst = 32'd268468224;
      40213: inst = 32'd201344841;
      40214: inst = 32'd203483685;
      40215: inst = 32'd471859200;
      40216: inst = 32'd136314880;
      40217: inst = 32'd268468224;
      40218: inst = 32'd201344842;
      40219: inst = 32'd203483685;
      40220: inst = 32'd471859200;
      40221: inst = 32'd136314880;
      40222: inst = 32'd268468224;
      40223: inst = 32'd201344843;
      40224: inst = 32'd203483685;
      40225: inst = 32'd471859200;
      40226: inst = 32'd136314880;
      40227: inst = 32'd268468224;
      40228: inst = 32'd201344844;
      40229: inst = 32'd203483685;
      40230: inst = 32'd471859200;
      40231: inst = 32'd136314880;
      40232: inst = 32'd268468224;
      40233: inst = 32'd201344845;
      40234: inst = 32'd203483685;
      40235: inst = 32'd471859200;
      40236: inst = 32'd136314880;
      40237: inst = 32'd268468224;
      40238: inst = 32'd201344846;
      40239: inst = 32'd203483685;
      40240: inst = 32'd471859200;
      40241: inst = 32'd136314880;
      40242: inst = 32'd268468224;
      40243: inst = 32'd201344847;
      40244: inst = 32'd203483685;
      40245: inst = 32'd471859200;
      40246: inst = 32'd136314880;
      40247: inst = 32'd268468224;
      40248: inst = 32'd201344848;
      40249: inst = 32'd203483685;
      40250: inst = 32'd471859200;
      40251: inst = 32'd136314880;
      40252: inst = 32'd268468224;
      40253: inst = 32'd201344849;
      40254: inst = 32'd203483685;
      40255: inst = 32'd471859200;
      40256: inst = 32'd136314880;
      40257: inst = 32'd268468224;
      40258: inst = 32'd201344850;
      40259: inst = 32'd203483685;
      40260: inst = 32'd471859200;
      40261: inst = 32'd136314880;
      40262: inst = 32'd268468224;
      40263: inst = 32'd201344851;
      40264: inst = 32'd203483685;
      40265: inst = 32'd471859200;
      40266: inst = 32'd136314880;
      40267: inst = 32'd268468224;
      40268: inst = 32'd201344852;
      40269: inst = 32'd203483685;
      40270: inst = 32'd471859200;
      40271: inst = 32'd136314880;
      40272: inst = 32'd268468224;
      40273: inst = 32'd201344853;
      40274: inst = 32'd203483685;
      40275: inst = 32'd471859200;
      40276: inst = 32'd136314880;
      40277: inst = 32'd268468224;
      40278: inst = 32'd201344854;
      40279: inst = 32'd203423744;
      40280: inst = 32'd471859200;
      40281: inst = 32'd136314880;
      40282: inst = 32'd268468224;
      40283: inst = 32'd201344855;
      40284: inst = 32'd203423744;
      40285: inst = 32'd471859200;
      40286: inst = 32'd136314880;
      40287: inst = 32'd268468224;
      40288: inst = 32'd201344856;
      40289: inst = 32'd203423744;
      40290: inst = 32'd471859200;
      40291: inst = 32'd136314880;
      40292: inst = 32'd268468224;
      40293: inst = 32'd201344857;
      40294: inst = 32'd203423744;
      40295: inst = 32'd471859200;
      40296: inst = 32'd136314880;
      40297: inst = 32'd268468224;
      40298: inst = 32'd201344858;
      40299: inst = 32'd203423744;
      40300: inst = 32'd471859200;
      40301: inst = 32'd136314880;
      40302: inst = 32'd268468224;
      40303: inst = 32'd201344859;
      40304: inst = 32'd203423744;
      40305: inst = 32'd471859200;
      40306: inst = 32'd136314880;
      40307: inst = 32'd268468224;
      40308: inst = 32'd201344860;
      40309: inst = 32'd203423744;
      40310: inst = 32'd471859200;
      40311: inst = 32'd136314880;
      40312: inst = 32'd268468224;
      40313: inst = 32'd201344861;
      40314: inst = 32'd203423744;
      40315: inst = 32'd471859200;
      40316: inst = 32'd136314880;
      40317: inst = 32'd268468224;
      40318: inst = 32'd201344862;
      40319: inst = 32'd203423744;
      40320: inst = 32'd471859200;
      40321: inst = 32'd136314880;
      40322: inst = 32'd268468224;
      40323: inst = 32'd201344863;
      40324: inst = 32'd203423744;
      40325: inst = 32'd471859200;
      40326: inst = 32'd136314880;
      40327: inst = 32'd268468224;
      40328: inst = 32'd201344864;
      40329: inst = 32'd203423744;
      40330: inst = 32'd471859200;
      40331: inst = 32'd136314880;
      40332: inst = 32'd268468224;
      40333: inst = 32'd201344865;
      40334: inst = 32'd203423744;
      40335: inst = 32'd471859200;
      40336: inst = 32'd136314880;
      40337: inst = 32'd268468224;
      40338: inst = 32'd201344866;
      40339: inst = 32'd203423744;
      40340: inst = 32'd471859200;
      40341: inst = 32'd136314880;
      40342: inst = 32'd268468224;
      40343: inst = 32'd201344867;
      40344: inst = 32'd203423744;
      40345: inst = 32'd471859200;
      40346: inst = 32'd136314880;
      40347: inst = 32'd268468224;
      40348: inst = 32'd201344868;
      40349: inst = 32'd203423744;
      40350: inst = 32'd471859200;
      40351: inst = 32'd136314880;
      40352: inst = 32'd268468224;
      40353: inst = 32'd201344869;
      40354: inst = 32'd203423744;
      40355: inst = 32'd471859200;
      40356: inst = 32'd136314880;
      40357: inst = 32'd268468224;
      40358: inst = 32'd201344870;
      40359: inst = 32'd203423744;
      40360: inst = 32'd471859200;
      40361: inst = 32'd136314880;
      40362: inst = 32'd268468224;
      40363: inst = 32'd201344871;
      40364: inst = 32'd203423744;
      40365: inst = 32'd471859200;
      40366: inst = 32'd136314880;
      40367: inst = 32'd268468224;
      40368: inst = 32'd201344872;
      40369: inst = 32'd203423744;
      40370: inst = 32'd471859200;
      40371: inst = 32'd136314880;
      40372: inst = 32'd268468224;
      40373: inst = 32'd201344873;
      40374: inst = 32'd203423744;
      40375: inst = 32'd471859200;
      40376: inst = 32'd136314880;
      40377: inst = 32'd268468224;
      40378: inst = 32'd201344874;
      40379: inst = 32'd203423744;
      40380: inst = 32'd471859200;
      40381: inst = 32'd136314880;
      40382: inst = 32'd268468224;
      40383: inst = 32'd201344875;
      40384: inst = 32'd203423744;
      40385: inst = 32'd471859200;
      40386: inst = 32'd136314880;
      40387: inst = 32'd268468224;
      40388: inst = 32'd201344876;
      40389: inst = 32'd203423744;
      40390: inst = 32'd471859200;
      40391: inst = 32'd136314880;
      40392: inst = 32'd268468224;
      40393: inst = 32'd201344877;
      40394: inst = 32'd203483685;
      40395: inst = 32'd471859200;
      40396: inst = 32'd136314880;
      40397: inst = 32'd268468224;
      40398: inst = 32'd201344878;
      40399: inst = 32'd203483685;
      40400: inst = 32'd471859200;
      40401: inst = 32'd136314880;
      40402: inst = 32'd268468224;
      40403: inst = 32'd201344879;
      40404: inst = 32'd203483685;
      40405: inst = 32'd471859200;
      40406: inst = 32'd136314880;
      40407: inst = 32'd268468224;
      40408: inst = 32'd201344880;
      40409: inst = 32'd203483685;
      40410: inst = 32'd471859200;
      40411: inst = 32'd136314880;
      40412: inst = 32'd268468224;
      40413: inst = 32'd201344881;
      40414: inst = 32'd203483685;
      40415: inst = 32'd471859200;
      40416: inst = 32'd136314880;
      40417: inst = 32'd268468224;
      40418: inst = 32'd201344882;
      40419: inst = 32'd203483685;
      40420: inst = 32'd471859200;
      40421: inst = 32'd136314880;
      40422: inst = 32'd268468224;
      40423: inst = 32'd201344883;
      40424: inst = 32'd203483685;
      40425: inst = 32'd471859200;
      40426: inst = 32'd136314880;
      40427: inst = 32'd268468224;
      40428: inst = 32'd201344884;
      40429: inst = 32'd203483685;
      40430: inst = 32'd471859200;
      40431: inst = 32'd136314880;
      40432: inst = 32'd268468224;
      40433: inst = 32'd201344885;
      40434: inst = 32'd203483685;
      40435: inst = 32'd471859200;
      40436: inst = 32'd136314880;
      40437: inst = 32'd268468224;
      40438: inst = 32'd201344886;
      40439: inst = 32'd203483685;
      40440: inst = 32'd471859200;
      40441: inst = 32'd136314880;
      40442: inst = 32'd268468224;
      40443: inst = 32'd201344887;
      40444: inst = 32'd203483685;
      40445: inst = 32'd471859200;
      40446: inst = 32'd136314880;
      40447: inst = 32'd268468224;
      40448: inst = 32'd201344888;
      40449: inst = 32'd203483685;
      40450: inst = 32'd471859200;
      40451: inst = 32'd136314880;
      40452: inst = 32'd268468224;
      40453: inst = 32'd201344889;
      40454: inst = 32'd203483685;
      40455: inst = 32'd471859200;
      40456: inst = 32'd136314880;
      40457: inst = 32'd268468224;
      40458: inst = 32'd201344890;
      40459: inst = 32'd203483685;
      40460: inst = 32'd471859200;
      40461: inst = 32'd136314880;
      40462: inst = 32'd268468224;
      40463: inst = 32'd201344891;
      40464: inst = 32'd203483685;
      40465: inst = 32'd471859200;
      40466: inst = 32'd136314880;
      40467: inst = 32'd268468224;
      40468: inst = 32'd201344892;
      40469: inst = 32'd203483685;
      40470: inst = 32'd471859200;
      40471: inst = 32'd136314880;
      40472: inst = 32'd268468224;
      40473: inst = 32'd201344893;
      40474: inst = 32'd203483685;
      40475: inst = 32'd471859200;
      40476: inst = 32'd136314880;
      40477: inst = 32'd268468224;
      40478: inst = 32'd201344894;
      40479: inst = 32'd203483685;
      40480: inst = 32'd471859200;
      40481: inst = 32'd136314880;
      40482: inst = 32'd268468224;
      40483: inst = 32'd201344895;
      40484: inst = 32'd203483685;
      40485: inst = 32'd471859200;
      40486: inst = 32'd136314880;
      40487: inst = 32'd268468224;
      40488: inst = 32'd201344896;
      40489: inst = 32'd203483685;
      40490: inst = 32'd471859200;
      40491: inst = 32'd136314880;
      40492: inst = 32'd268468224;
      40493: inst = 32'd201344897;
      40494: inst = 32'd203483685;
      40495: inst = 32'd471859200;
      40496: inst = 32'd136314880;
      40497: inst = 32'd268468224;
      40498: inst = 32'd201344898;
      40499: inst = 32'd203483685;
      40500: inst = 32'd471859200;
      40501: inst = 32'd136314880;
      40502: inst = 32'd268468224;
      40503: inst = 32'd201344899;
      40504: inst = 32'd203483685;
      40505: inst = 32'd471859200;
      40506: inst = 32'd136314880;
      40507: inst = 32'd268468224;
      40508: inst = 32'd201344900;
      40509: inst = 32'd203483685;
      40510: inst = 32'd471859200;
      40511: inst = 32'd136314880;
      40512: inst = 32'd268468224;
      40513: inst = 32'd201344901;
      40514: inst = 32'd203483685;
      40515: inst = 32'd471859200;
      40516: inst = 32'd136314880;
      40517: inst = 32'd268468224;
      40518: inst = 32'd201344902;
      40519: inst = 32'd203483685;
      40520: inst = 32'd471859200;
      40521: inst = 32'd136314880;
      40522: inst = 32'd268468224;
      40523: inst = 32'd201344903;
      40524: inst = 32'd203483685;
      40525: inst = 32'd471859200;
      40526: inst = 32'd136314880;
      40527: inst = 32'd268468224;
      40528: inst = 32'd201344904;
      40529: inst = 32'd203483685;
      40530: inst = 32'd471859200;
      40531: inst = 32'd136314880;
      40532: inst = 32'd268468224;
      40533: inst = 32'd201344905;
      40534: inst = 32'd203483685;
      40535: inst = 32'd471859200;
      40536: inst = 32'd136314880;
      40537: inst = 32'd268468224;
      40538: inst = 32'd201344906;
      40539: inst = 32'd203483685;
      40540: inst = 32'd471859200;
      40541: inst = 32'd136314880;
      40542: inst = 32'd268468224;
      40543: inst = 32'd201344907;
      40544: inst = 32'd203483685;
      40545: inst = 32'd471859200;
      40546: inst = 32'd136314880;
      40547: inst = 32'd268468224;
      40548: inst = 32'd201344908;
      40549: inst = 32'd203483685;
      40550: inst = 32'd471859200;
      40551: inst = 32'd136314880;
      40552: inst = 32'd268468224;
      40553: inst = 32'd201344909;
      40554: inst = 32'd203483685;
      40555: inst = 32'd471859200;
      40556: inst = 32'd136314880;
      40557: inst = 32'd268468224;
      40558: inst = 32'd201344910;
      40559: inst = 32'd203483685;
      40560: inst = 32'd471859200;
      40561: inst = 32'd136314880;
      40562: inst = 32'd268468224;
      40563: inst = 32'd201344911;
      40564: inst = 32'd203483685;
      40565: inst = 32'd471859200;
      40566: inst = 32'd136314880;
      40567: inst = 32'd268468224;
      40568: inst = 32'd201344912;
      40569: inst = 32'd203483685;
      40570: inst = 32'd471859200;
      40571: inst = 32'd136314880;
      40572: inst = 32'd268468224;
      40573: inst = 32'd201344913;
      40574: inst = 32'd203483685;
      40575: inst = 32'd471859200;
      40576: inst = 32'd136314880;
      40577: inst = 32'd268468224;
      40578: inst = 32'd201344914;
      40579: inst = 32'd203483685;
      40580: inst = 32'd471859200;
      40581: inst = 32'd136314880;
      40582: inst = 32'd268468224;
      40583: inst = 32'd201344915;
      40584: inst = 32'd203483685;
      40585: inst = 32'd471859200;
      40586: inst = 32'd136314880;
      40587: inst = 32'd268468224;
      40588: inst = 32'd201344916;
      40589: inst = 32'd203483685;
      40590: inst = 32'd471859200;
      40591: inst = 32'd136314880;
      40592: inst = 32'd268468224;
      40593: inst = 32'd201344917;
      40594: inst = 32'd203483685;
      40595: inst = 32'd471859200;
      40596: inst = 32'd136314880;
      40597: inst = 32'd268468224;
      40598: inst = 32'd201344918;
      40599: inst = 32'd203483685;
      40600: inst = 32'd471859200;
      40601: inst = 32'd136314880;
      40602: inst = 32'd268468224;
      40603: inst = 32'd201344919;
      40604: inst = 32'd203483685;
      40605: inst = 32'd471859200;
      40606: inst = 32'd136314880;
      40607: inst = 32'd268468224;
      40608: inst = 32'd201344920;
      40609: inst = 32'd203483685;
      40610: inst = 32'd471859200;
      40611: inst = 32'd136314880;
      40612: inst = 32'd268468224;
      40613: inst = 32'd201344921;
      40614: inst = 32'd203483685;
      40615: inst = 32'd471859200;
      40616: inst = 32'd136314880;
      40617: inst = 32'd268468224;
      40618: inst = 32'd201344922;
      40619: inst = 32'd203483685;
      40620: inst = 32'd471859200;
      40621: inst = 32'd136314880;
      40622: inst = 32'd268468224;
      40623: inst = 32'd201344923;
      40624: inst = 32'd203483685;
      40625: inst = 32'd471859200;
      40626: inst = 32'd136314880;
      40627: inst = 32'd268468224;
      40628: inst = 32'd201344924;
      40629: inst = 32'd203483685;
      40630: inst = 32'd471859200;
      40631: inst = 32'd136314880;
      40632: inst = 32'd268468224;
      40633: inst = 32'd201344925;
      40634: inst = 32'd203423744;
      40635: inst = 32'd471859200;
      40636: inst = 32'd136314880;
      40637: inst = 32'd268468224;
      40638: inst = 32'd201344926;
      40639: inst = 32'd203483685;
      40640: inst = 32'd471859200;
      40641: inst = 32'd136314880;
      40642: inst = 32'd268468224;
      40643: inst = 32'd201344927;
      40644: inst = 32'd203483685;
      40645: inst = 32'd471859200;
      40646: inst = 32'd136314880;
      40647: inst = 32'd268468224;
      40648: inst = 32'd201344928;
      40649: inst = 32'd203483685;
      40650: inst = 32'd471859200;
      40651: inst = 32'd136314880;
      40652: inst = 32'd268468224;
      40653: inst = 32'd201344929;
      40654: inst = 32'd203483685;
      40655: inst = 32'd471859200;
      40656: inst = 32'd136314880;
      40657: inst = 32'd268468224;
      40658: inst = 32'd201344930;
      40659: inst = 32'd203483685;
      40660: inst = 32'd471859200;
      40661: inst = 32'd136314880;
      40662: inst = 32'd268468224;
      40663: inst = 32'd201344931;
      40664: inst = 32'd203483685;
      40665: inst = 32'd471859200;
      40666: inst = 32'd136314880;
      40667: inst = 32'd268468224;
      40668: inst = 32'd201344932;
      40669: inst = 32'd203483685;
      40670: inst = 32'd471859200;
      40671: inst = 32'd136314880;
      40672: inst = 32'd268468224;
      40673: inst = 32'd201344933;
      40674: inst = 32'd203483685;
      40675: inst = 32'd471859200;
      40676: inst = 32'd136314880;
      40677: inst = 32'd268468224;
      40678: inst = 32'd201344934;
      40679: inst = 32'd203483685;
      40680: inst = 32'd471859200;
      40681: inst = 32'd136314880;
      40682: inst = 32'd268468224;
      40683: inst = 32'd201344935;
      40684: inst = 32'd203483685;
      40685: inst = 32'd471859200;
      40686: inst = 32'd136314880;
      40687: inst = 32'd268468224;
      40688: inst = 32'd201344936;
      40689: inst = 32'd203483685;
      40690: inst = 32'd471859200;
      40691: inst = 32'd136314880;
      40692: inst = 32'd268468224;
      40693: inst = 32'd201344937;
      40694: inst = 32'd203483685;
      40695: inst = 32'd471859200;
      40696: inst = 32'd136314880;
      40697: inst = 32'd268468224;
      40698: inst = 32'd201344938;
      40699: inst = 32'd203483685;
      40700: inst = 32'd471859200;
      40701: inst = 32'd136314880;
      40702: inst = 32'd268468224;
      40703: inst = 32'd201344939;
      40704: inst = 32'd203483685;
      40705: inst = 32'd471859200;
      40706: inst = 32'd136314880;
      40707: inst = 32'd268468224;
      40708: inst = 32'd201344940;
      40709: inst = 32'd203483685;
      40710: inst = 32'd471859200;
      40711: inst = 32'd136314880;
      40712: inst = 32'd268468224;
      40713: inst = 32'd201344941;
      40714: inst = 32'd203483685;
      40715: inst = 32'd471859200;
      40716: inst = 32'd136314880;
      40717: inst = 32'd268468224;
      40718: inst = 32'd201344942;
      40719: inst = 32'd203483685;
      40720: inst = 32'd471859200;
      40721: inst = 32'd136314880;
      40722: inst = 32'd268468224;
      40723: inst = 32'd201344943;
      40724: inst = 32'd203483685;
      40725: inst = 32'd471859200;
      40726: inst = 32'd136314880;
      40727: inst = 32'd268468224;
      40728: inst = 32'd201344944;
      40729: inst = 32'd203483685;
      40730: inst = 32'd471859200;
      40731: inst = 32'd136314880;
      40732: inst = 32'd268468224;
      40733: inst = 32'd201344945;
      40734: inst = 32'd203483685;
      40735: inst = 32'd471859200;
      40736: inst = 32'd136314880;
      40737: inst = 32'd268468224;
      40738: inst = 32'd201344946;
      40739: inst = 32'd203483685;
      40740: inst = 32'd471859200;
      40741: inst = 32'd136314880;
      40742: inst = 32'd268468224;
      40743: inst = 32'd201344947;
      40744: inst = 32'd203483685;
      40745: inst = 32'd471859200;
      40746: inst = 32'd136314880;
      40747: inst = 32'd268468224;
      40748: inst = 32'd201344948;
      40749: inst = 32'd203483685;
      40750: inst = 32'd471859200;
      40751: inst = 32'd136314880;
      40752: inst = 32'd268468224;
      40753: inst = 32'd201344949;
      40754: inst = 32'd203483685;
      40755: inst = 32'd471859200;
      40756: inst = 32'd136314880;
      40757: inst = 32'd268468224;
      40758: inst = 32'd201344950;
      40759: inst = 32'd203423744;
      40760: inst = 32'd471859200;
      40761: inst = 32'd136314880;
      40762: inst = 32'd268468224;
      40763: inst = 32'd201344951;
      40764: inst = 32'd203423744;
      40765: inst = 32'd471859200;
      40766: inst = 32'd136314880;
      40767: inst = 32'd268468224;
      40768: inst = 32'd201344952;
      40769: inst = 32'd203423744;
      40770: inst = 32'd471859200;
      40771: inst = 32'd136314880;
      40772: inst = 32'd268468224;
      40773: inst = 32'd201344953;
      40774: inst = 32'd203423744;
      40775: inst = 32'd471859200;
      40776: inst = 32'd136314880;
      40777: inst = 32'd268468224;
      40778: inst = 32'd201344954;
      40779: inst = 32'd203423744;
      40780: inst = 32'd471859200;
      40781: inst = 32'd136314880;
      40782: inst = 32'd268468224;
      40783: inst = 32'd201344955;
      40784: inst = 32'd203423744;
      40785: inst = 32'd471859200;
      40786: inst = 32'd136314880;
      40787: inst = 32'd268468224;
      40788: inst = 32'd201344956;
      40789: inst = 32'd203423744;
      40790: inst = 32'd471859200;
      40791: inst = 32'd136314880;
      40792: inst = 32'd268468224;
      40793: inst = 32'd201344957;
      40794: inst = 32'd203423744;
      40795: inst = 32'd471859200;
      40796: inst = 32'd136314880;
      40797: inst = 32'd268468224;
      40798: inst = 32'd201344958;
      40799: inst = 32'd203423744;
      40800: inst = 32'd471859200;
      40801: inst = 32'd136314880;
      40802: inst = 32'd268468224;
      40803: inst = 32'd201344959;
      40804: inst = 32'd203423744;
      40805: inst = 32'd471859200;
      40806: inst = 32'd136314880;
      40807: inst = 32'd268468224;
      40808: inst = 32'd201344960;
      40809: inst = 32'd203423744;
      40810: inst = 32'd471859200;
      40811: inst = 32'd136314880;
      40812: inst = 32'd268468224;
      40813: inst = 32'd201344961;
      40814: inst = 32'd203423744;
      40815: inst = 32'd471859200;
      40816: inst = 32'd136314880;
      40817: inst = 32'd268468224;
      40818: inst = 32'd201344962;
      40819: inst = 32'd203423744;
      40820: inst = 32'd471859200;
      40821: inst = 32'd136314880;
      40822: inst = 32'd268468224;
      40823: inst = 32'd201344963;
      40824: inst = 32'd203423744;
      40825: inst = 32'd471859200;
      40826: inst = 32'd136314880;
      40827: inst = 32'd268468224;
      40828: inst = 32'd201344964;
      40829: inst = 32'd203423744;
      40830: inst = 32'd471859200;
      40831: inst = 32'd136314880;
      40832: inst = 32'd268468224;
      40833: inst = 32'd201344965;
      40834: inst = 32'd203423744;
      40835: inst = 32'd471859200;
      40836: inst = 32'd136314880;
      40837: inst = 32'd268468224;
      40838: inst = 32'd201344966;
      40839: inst = 32'd203423744;
      40840: inst = 32'd471859200;
      40841: inst = 32'd136314880;
      40842: inst = 32'd268468224;
      40843: inst = 32'd201344967;
      40844: inst = 32'd203423744;
      40845: inst = 32'd471859200;
      40846: inst = 32'd136314880;
      40847: inst = 32'd268468224;
      40848: inst = 32'd201344968;
      40849: inst = 32'd203423744;
      40850: inst = 32'd471859200;
      40851: inst = 32'd136314880;
      40852: inst = 32'd268468224;
      40853: inst = 32'd201344969;
      40854: inst = 32'd203423744;
      40855: inst = 32'd471859200;
      40856: inst = 32'd136314880;
      40857: inst = 32'd268468224;
      40858: inst = 32'd201344970;
      40859: inst = 32'd203423744;
      40860: inst = 32'd471859200;
      40861: inst = 32'd136314880;
      40862: inst = 32'd268468224;
      40863: inst = 32'd201344971;
      40864: inst = 32'd203423744;
      40865: inst = 32'd471859200;
      40866: inst = 32'd136314880;
      40867: inst = 32'd268468224;
      40868: inst = 32'd201344972;
      40869: inst = 32'd203423744;
      40870: inst = 32'd471859200;
      40871: inst = 32'd136314880;
      40872: inst = 32'd268468224;
      40873: inst = 32'd201344973;
      40874: inst = 32'd203483685;
      40875: inst = 32'd471859200;
      40876: inst = 32'd136314880;
      40877: inst = 32'd268468224;
      40878: inst = 32'd201344974;
      40879: inst = 32'd203483685;
      40880: inst = 32'd471859200;
      40881: inst = 32'd136314880;
      40882: inst = 32'd268468224;
      40883: inst = 32'd201344975;
      40884: inst = 32'd203483685;
      40885: inst = 32'd471859200;
      40886: inst = 32'd136314880;
      40887: inst = 32'd268468224;
      40888: inst = 32'd201344976;
      40889: inst = 32'd203483685;
      40890: inst = 32'd471859200;
      40891: inst = 32'd136314880;
      40892: inst = 32'd268468224;
      40893: inst = 32'd201344977;
      40894: inst = 32'd203483685;
      40895: inst = 32'd471859200;
      40896: inst = 32'd136314880;
      40897: inst = 32'd268468224;
      40898: inst = 32'd201344978;
      40899: inst = 32'd203483685;
      40900: inst = 32'd471859200;
      40901: inst = 32'd136314880;
      40902: inst = 32'd268468224;
      40903: inst = 32'd201344979;
      40904: inst = 32'd203483685;
      40905: inst = 32'd471859200;
      40906: inst = 32'd136314880;
      40907: inst = 32'd268468224;
      40908: inst = 32'd201344980;
      40909: inst = 32'd203483685;
      40910: inst = 32'd471859200;
      40911: inst = 32'd136314880;
      40912: inst = 32'd268468224;
      40913: inst = 32'd201344981;
      40914: inst = 32'd203483685;
      40915: inst = 32'd471859200;
      40916: inst = 32'd136314880;
      40917: inst = 32'd268468224;
      40918: inst = 32'd201344982;
      40919: inst = 32'd203483685;
      40920: inst = 32'd471859200;
      40921: inst = 32'd136314880;
      40922: inst = 32'd268468224;
      40923: inst = 32'd201344983;
      40924: inst = 32'd203423744;
      40925: inst = 32'd471859200;
      40926: inst = 32'd136314880;
      40927: inst = 32'd268468224;
      40928: inst = 32'd201344984;
      40929: inst = 32'd203483685;
      40930: inst = 32'd471859200;
      40931: inst = 32'd136314880;
      40932: inst = 32'd268468224;
      40933: inst = 32'd201344985;
      40934: inst = 32'd203483685;
      40935: inst = 32'd471859200;
      40936: inst = 32'd136314880;
      40937: inst = 32'd268468224;
      40938: inst = 32'd201344986;
      40939: inst = 32'd203483685;
      40940: inst = 32'd471859200;
      40941: inst = 32'd136314880;
      40942: inst = 32'd268468224;
      40943: inst = 32'd201344987;
      40944: inst = 32'd203483685;
      40945: inst = 32'd471859200;
      40946: inst = 32'd136314880;
      40947: inst = 32'd268468224;
      40948: inst = 32'd201344988;
      40949: inst = 32'd203483685;
      40950: inst = 32'd471859200;
      40951: inst = 32'd136314880;
      40952: inst = 32'd268468224;
      40953: inst = 32'd201344989;
      40954: inst = 32'd203483685;
      40955: inst = 32'd471859200;
      40956: inst = 32'd136314880;
      40957: inst = 32'd268468224;
      40958: inst = 32'd201344990;
      40959: inst = 32'd203483685;
      40960: inst = 32'd471859200;
      40961: inst = 32'd136314880;
      40962: inst = 32'd268468224;
      40963: inst = 32'd201344991;
      40964: inst = 32'd203483685;
      40965: inst = 32'd471859200;
      40966: inst = 32'd136314880;
      40967: inst = 32'd268468224;
      40968: inst = 32'd201344992;
      40969: inst = 32'd203483685;
      40970: inst = 32'd471859200;
      40971: inst = 32'd136314880;
      40972: inst = 32'd268468224;
      40973: inst = 32'd201344993;
      40974: inst = 32'd203483685;
      40975: inst = 32'd471859200;
      40976: inst = 32'd136314880;
      40977: inst = 32'd268468224;
      40978: inst = 32'd201344994;
      40979: inst = 32'd203423744;
      40980: inst = 32'd471859200;
      40981: inst = 32'd136314880;
      40982: inst = 32'd268468224;
      40983: inst = 32'd201344995;
      40984: inst = 32'd203423744;
      40985: inst = 32'd471859200;
      40986: inst = 32'd136314880;
      40987: inst = 32'd268468224;
      40988: inst = 32'd201344996;
      40989: inst = 32'd203483685;
      40990: inst = 32'd471859200;
      40991: inst = 32'd136314880;
      40992: inst = 32'd268468224;
      40993: inst = 32'd201344997;
      40994: inst = 32'd203483685;
      40995: inst = 32'd471859200;
      40996: inst = 32'd136314880;
      40997: inst = 32'd268468224;
      40998: inst = 32'd201344998;
      40999: inst = 32'd203483685;
      41000: inst = 32'd471859200;
      41001: inst = 32'd136314880;
      41002: inst = 32'd268468224;
      41003: inst = 32'd201344999;
      41004: inst = 32'd203483685;
      41005: inst = 32'd471859200;
      41006: inst = 32'd136314880;
      41007: inst = 32'd268468224;
      41008: inst = 32'd201345000;
      41009: inst = 32'd203483685;
      41010: inst = 32'd471859200;
      41011: inst = 32'd136314880;
      41012: inst = 32'd268468224;
      41013: inst = 32'd201345001;
      41014: inst = 32'd203483685;
      41015: inst = 32'd471859200;
      41016: inst = 32'd136314880;
      41017: inst = 32'd268468224;
      41018: inst = 32'd201345002;
      41019: inst = 32'd203483685;
      41020: inst = 32'd471859200;
      41021: inst = 32'd136314880;
      41022: inst = 32'd268468224;
      41023: inst = 32'd201345003;
      41024: inst = 32'd203483685;
      41025: inst = 32'd471859200;
      41026: inst = 32'd136314880;
      41027: inst = 32'd268468224;
      41028: inst = 32'd201345004;
      41029: inst = 32'd203483685;
      41030: inst = 32'd471859200;
      41031: inst = 32'd136314880;
      41032: inst = 32'd268468224;
      41033: inst = 32'd201345005;
      41034: inst = 32'd203483685;
      41035: inst = 32'd471859200;
      41036: inst = 32'd136314880;
      41037: inst = 32'd268468224;
      41038: inst = 32'd201345006;
      41039: inst = 32'd203483685;
      41040: inst = 32'd471859200;
      41041: inst = 32'd136314880;
      41042: inst = 32'd268468224;
      41043: inst = 32'd201345007;
      41044: inst = 32'd203483685;
      41045: inst = 32'd471859200;
      41046: inst = 32'd136314880;
      41047: inst = 32'd268468224;
      41048: inst = 32'd201345008;
      41049: inst = 32'd203483685;
      41050: inst = 32'd471859200;
      41051: inst = 32'd136314880;
      41052: inst = 32'd268468224;
      41053: inst = 32'd201345009;
      41054: inst = 32'd203483685;
      41055: inst = 32'd471859200;
      41056: inst = 32'd136314880;
      41057: inst = 32'd268468224;
      41058: inst = 32'd201345010;
      41059: inst = 32'd203483685;
      41060: inst = 32'd471859200;
      41061: inst = 32'd136314880;
      41062: inst = 32'd268468224;
      41063: inst = 32'd201345011;
      41064: inst = 32'd203483685;
      41065: inst = 32'd471859200;
      41066: inst = 32'd136314880;
      41067: inst = 32'd268468224;
      41068: inst = 32'd201345012;
      41069: inst = 32'd203483685;
      41070: inst = 32'd471859200;
      41071: inst = 32'd136314880;
      41072: inst = 32'd268468224;
      41073: inst = 32'd201345013;
      41074: inst = 32'd203483685;
      41075: inst = 32'd471859200;
      41076: inst = 32'd136314880;
      41077: inst = 32'd268468224;
      41078: inst = 32'd201345014;
      41079: inst = 32'd203483685;
      41080: inst = 32'd471859200;
      41081: inst = 32'd136314880;
      41082: inst = 32'd268468224;
      41083: inst = 32'd201345015;
      41084: inst = 32'd203483685;
      41085: inst = 32'd471859200;
      41086: inst = 32'd136314880;
      41087: inst = 32'd268468224;
      41088: inst = 32'd201345016;
      41089: inst = 32'd203483685;
      41090: inst = 32'd471859200;
      41091: inst = 32'd136314880;
      41092: inst = 32'd268468224;
      41093: inst = 32'd201345017;
      41094: inst = 32'd203483685;
      41095: inst = 32'd471859200;
      41096: inst = 32'd136314880;
      41097: inst = 32'd268468224;
      41098: inst = 32'd201345018;
      41099: inst = 32'd203483685;
      41100: inst = 32'd471859200;
      41101: inst = 32'd136314880;
      41102: inst = 32'd268468224;
      41103: inst = 32'd201345019;
      41104: inst = 32'd203483685;
      41105: inst = 32'd471859200;
      41106: inst = 32'd136314880;
      41107: inst = 32'd268468224;
      41108: inst = 32'd201345020;
      41109: inst = 32'd203423744;
      41110: inst = 32'd471859200;
      41111: inst = 32'd136314880;
      41112: inst = 32'd268468224;
      41113: inst = 32'd201345021;
      41114: inst = 32'd203423744;
      41115: inst = 32'd471859200;
      41116: inst = 32'd136314880;
      41117: inst = 32'd268468224;
      41118: inst = 32'd201345022;
      41119: inst = 32'd203483685;
      41120: inst = 32'd471859200;
      41121: inst = 32'd136314880;
      41122: inst = 32'd268468224;
      41123: inst = 32'd201345023;
      41124: inst = 32'd203483685;
      41125: inst = 32'd471859200;
      41126: inst = 32'd136314880;
      41127: inst = 32'd268468224;
      41128: inst = 32'd201345024;
      41129: inst = 32'd203483685;
      41130: inst = 32'd471859200;
      41131: inst = 32'd136314880;
      41132: inst = 32'd268468224;
      41133: inst = 32'd201345025;
      41134: inst = 32'd203483685;
      41135: inst = 32'd471859200;
      41136: inst = 32'd136314880;
      41137: inst = 32'd268468224;
      41138: inst = 32'd201345026;
      41139: inst = 32'd203483685;
      41140: inst = 32'd471859200;
      41141: inst = 32'd136314880;
      41142: inst = 32'd268468224;
      41143: inst = 32'd201345027;
      41144: inst = 32'd203483685;
      41145: inst = 32'd471859200;
      41146: inst = 32'd136314880;
      41147: inst = 32'd268468224;
      41148: inst = 32'd201345028;
      41149: inst = 32'd203483685;
      41150: inst = 32'd471859200;
      41151: inst = 32'd136314880;
      41152: inst = 32'd268468224;
      41153: inst = 32'd201345029;
      41154: inst = 32'd203483685;
      41155: inst = 32'd471859200;
      41156: inst = 32'd136314880;
      41157: inst = 32'd268468224;
      41158: inst = 32'd201345030;
      41159: inst = 32'd203483685;
      41160: inst = 32'd471859200;
      41161: inst = 32'd136314880;
      41162: inst = 32'd268468224;
      41163: inst = 32'd201345031;
      41164: inst = 32'd203483685;
      41165: inst = 32'd471859200;
      41166: inst = 32'd136314880;
      41167: inst = 32'd268468224;
      41168: inst = 32'd201345032;
      41169: inst = 32'd203483685;
      41170: inst = 32'd471859200;
      41171: inst = 32'd136314880;
      41172: inst = 32'd268468224;
      41173: inst = 32'd201345033;
      41174: inst = 32'd203483685;
      41175: inst = 32'd471859200;
      41176: inst = 32'd136314880;
      41177: inst = 32'd268468224;
      41178: inst = 32'd201345034;
      41179: inst = 32'd203483685;
      41180: inst = 32'd471859200;
      41181: inst = 32'd136314880;
      41182: inst = 32'd268468224;
      41183: inst = 32'd201345035;
      41184: inst = 32'd203483685;
      41185: inst = 32'd471859200;
      41186: inst = 32'd136314880;
      41187: inst = 32'd268468224;
      41188: inst = 32'd201345036;
      41189: inst = 32'd203483685;
      41190: inst = 32'd471859200;
      41191: inst = 32'd136314880;
      41192: inst = 32'd268468224;
      41193: inst = 32'd201345037;
      41194: inst = 32'd203483685;
      41195: inst = 32'd471859200;
      41196: inst = 32'd136314880;
      41197: inst = 32'd268468224;
      41198: inst = 32'd201345038;
      41199: inst = 32'd203483685;
      41200: inst = 32'd471859200;
      41201: inst = 32'd136314880;
      41202: inst = 32'd268468224;
      41203: inst = 32'd201345039;
      41204: inst = 32'd203483685;
      41205: inst = 32'd471859200;
      41206: inst = 32'd136314880;
      41207: inst = 32'd268468224;
      41208: inst = 32'd201345040;
      41209: inst = 32'd203483685;
      41210: inst = 32'd471859200;
      41211: inst = 32'd136314880;
      41212: inst = 32'd268468224;
      41213: inst = 32'd201345041;
      41214: inst = 32'd203483685;
      41215: inst = 32'd471859200;
      41216: inst = 32'd136314880;
      41217: inst = 32'd268468224;
      41218: inst = 32'd201345042;
      41219: inst = 32'd203483685;
      41220: inst = 32'd471859200;
      41221: inst = 32'd136314880;
      41222: inst = 32'd268468224;
      41223: inst = 32'd201345043;
      41224: inst = 32'd203483685;
      41225: inst = 32'd471859200;
      41226: inst = 32'd136314880;
      41227: inst = 32'd268468224;
      41228: inst = 32'd201345044;
      41229: inst = 32'd203483685;
      41230: inst = 32'd471859200;
      41231: inst = 32'd136314880;
      41232: inst = 32'd268468224;
      41233: inst = 32'd201345045;
      41234: inst = 32'd203483685;
      41235: inst = 32'd471859200;
      41236: inst = 32'd136314880;
      41237: inst = 32'd268468224;
      41238: inst = 32'd201345046;
      41239: inst = 32'd203423744;
      41240: inst = 32'd471859200;
      41241: inst = 32'd136314880;
      41242: inst = 32'd268468224;
      41243: inst = 32'd201345047;
      41244: inst = 32'd203423744;
      41245: inst = 32'd471859200;
      41246: inst = 32'd136314880;
      41247: inst = 32'd268468224;
      41248: inst = 32'd201345048;
      41249: inst = 32'd203423744;
      41250: inst = 32'd471859200;
      41251: inst = 32'd136314880;
      41252: inst = 32'd268468224;
      41253: inst = 32'd201345049;
      41254: inst = 32'd203423744;
      41255: inst = 32'd471859200;
      41256: inst = 32'd136314880;
      41257: inst = 32'd268468224;
      41258: inst = 32'd201345050;
      41259: inst = 32'd203423744;
      41260: inst = 32'd471859200;
      41261: inst = 32'd136314880;
      41262: inst = 32'd268468224;
      41263: inst = 32'd201345051;
      41264: inst = 32'd203423744;
      41265: inst = 32'd471859200;
      41266: inst = 32'd136314880;
      41267: inst = 32'd268468224;
      41268: inst = 32'd201345052;
      41269: inst = 32'd203423744;
      41270: inst = 32'd471859200;
      41271: inst = 32'd136314880;
      41272: inst = 32'd268468224;
      41273: inst = 32'd201345053;
      41274: inst = 32'd203423744;
      41275: inst = 32'd471859200;
      41276: inst = 32'd136314880;
      41277: inst = 32'd268468224;
      41278: inst = 32'd201345054;
      41279: inst = 32'd203423744;
      41280: inst = 32'd471859200;
      41281: inst = 32'd136314880;
      41282: inst = 32'd268468224;
      41283: inst = 32'd201345055;
      41284: inst = 32'd203423744;
      41285: inst = 32'd471859200;
      41286: inst = 32'd136314880;
      41287: inst = 32'd268468224;
      41288: inst = 32'd201345056;
      41289: inst = 32'd203423744;
      41290: inst = 32'd471859200;
      41291: inst = 32'd136314880;
      41292: inst = 32'd268468224;
      41293: inst = 32'd201345057;
      41294: inst = 32'd203423744;
      41295: inst = 32'd471859200;
      41296: inst = 32'd136314880;
      41297: inst = 32'd268468224;
      41298: inst = 32'd201345058;
      41299: inst = 32'd203423744;
      41300: inst = 32'd471859200;
      41301: inst = 32'd136314880;
      41302: inst = 32'd268468224;
      41303: inst = 32'd201345059;
      41304: inst = 32'd203423744;
      41305: inst = 32'd471859200;
      41306: inst = 32'd136314880;
      41307: inst = 32'd268468224;
      41308: inst = 32'd201345060;
      41309: inst = 32'd203423744;
      41310: inst = 32'd471859200;
      41311: inst = 32'd136314880;
      41312: inst = 32'd268468224;
      41313: inst = 32'd201345061;
      41314: inst = 32'd203423744;
      41315: inst = 32'd471859200;
      41316: inst = 32'd136314880;
      41317: inst = 32'd268468224;
      41318: inst = 32'd201345062;
      41319: inst = 32'd203423744;
      41320: inst = 32'd471859200;
      41321: inst = 32'd136314880;
      41322: inst = 32'd268468224;
      41323: inst = 32'd201345063;
      41324: inst = 32'd203423744;
      41325: inst = 32'd471859200;
      41326: inst = 32'd136314880;
      41327: inst = 32'd268468224;
      41328: inst = 32'd201345064;
      41329: inst = 32'd203423744;
      41330: inst = 32'd471859200;
      41331: inst = 32'd136314880;
      41332: inst = 32'd268468224;
      41333: inst = 32'd201345065;
      41334: inst = 32'd203423744;
      41335: inst = 32'd471859200;
      41336: inst = 32'd136314880;
      41337: inst = 32'd268468224;
      41338: inst = 32'd201345066;
      41339: inst = 32'd203423744;
      41340: inst = 32'd471859200;
      41341: inst = 32'd136314880;
      41342: inst = 32'd268468224;
      41343: inst = 32'd201345067;
      41344: inst = 32'd203423744;
      41345: inst = 32'd471859200;
      41346: inst = 32'd136314880;
      41347: inst = 32'd268468224;
      41348: inst = 32'd201345068;
      41349: inst = 32'd203423744;
      41350: inst = 32'd471859200;
      41351: inst = 32'd136314880;
      41352: inst = 32'd268468224;
      41353: inst = 32'd201345069;
      41354: inst = 32'd203423744;
      41355: inst = 32'd471859200;
      41356: inst = 32'd136314880;
      41357: inst = 32'd268468224;
      41358: inst = 32'd201345070;
      41359: inst = 32'd203423744;
      41360: inst = 32'd471859200;
      41361: inst = 32'd136314880;
      41362: inst = 32'd268468224;
      41363: inst = 32'd201345071;
      41364: inst = 32'd203423744;
      41365: inst = 32'd471859200;
      41366: inst = 32'd136314880;
      41367: inst = 32'd268468224;
      41368: inst = 32'd201345072;
      41369: inst = 32'd203423744;
      41370: inst = 32'd471859200;
      41371: inst = 32'd136314880;
      41372: inst = 32'd268468224;
      41373: inst = 32'd201345073;
      41374: inst = 32'd203423744;
      41375: inst = 32'd471859200;
      41376: inst = 32'd136314880;
      41377: inst = 32'd268468224;
      41378: inst = 32'd201345074;
      41379: inst = 32'd203423744;
      41380: inst = 32'd471859200;
      41381: inst = 32'd136314880;
      41382: inst = 32'd268468224;
      41383: inst = 32'd201345075;
      41384: inst = 32'd203423744;
      41385: inst = 32'd471859200;
      41386: inst = 32'd136314880;
      41387: inst = 32'd268468224;
      41388: inst = 32'd201345076;
      41389: inst = 32'd203423744;
      41390: inst = 32'd471859200;
      41391: inst = 32'd136314880;
      41392: inst = 32'd268468224;
      41393: inst = 32'd201345077;
      41394: inst = 32'd203423744;
      41395: inst = 32'd471859200;
      41396: inst = 32'd136314880;
      41397: inst = 32'd268468224;
      41398: inst = 32'd201345078;
      41399: inst = 32'd203423744;
      41400: inst = 32'd471859200;
      41401: inst = 32'd136314880;
      41402: inst = 32'd268468224;
      41403: inst = 32'd201345079;
      41404: inst = 32'd203423744;
      41405: inst = 32'd471859200;
      41406: inst = 32'd136314880;
      41407: inst = 32'd268468224;
      41408: inst = 32'd201345080;
      41409: inst = 32'd203423744;
      41410: inst = 32'd471859200;
      41411: inst = 32'd136314880;
      41412: inst = 32'd268468224;
      41413: inst = 32'd201345081;
      41414: inst = 32'd203423744;
      41415: inst = 32'd471859200;
      41416: inst = 32'd136314880;
      41417: inst = 32'd268468224;
      41418: inst = 32'd201345082;
      41419: inst = 32'd203423744;
      41420: inst = 32'd471859200;
      41421: inst = 32'd136314880;
      41422: inst = 32'd268468224;
      41423: inst = 32'd201345083;
      41424: inst = 32'd203423744;
      41425: inst = 32'd471859200;
      41426: inst = 32'd136314880;
      41427: inst = 32'd268468224;
      41428: inst = 32'd201345084;
      41429: inst = 32'd203423744;
      41430: inst = 32'd471859200;
      41431: inst = 32'd136314880;
      41432: inst = 32'd268468224;
      41433: inst = 32'd201345085;
      41434: inst = 32'd203423744;
      41435: inst = 32'd471859200;
      41436: inst = 32'd136314880;
      41437: inst = 32'd268468224;
      41438: inst = 32'd201345086;
      41439: inst = 32'd203423744;
      41440: inst = 32'd471859200;
      41441: inst = 32'd136314880;
      41442: inst = 32'd268468224;
      41443: inst = 32'd201345087;
      41444: inst = 32'd203423744;
      41445: inst = 32'd471859200;
      41446: inst = 32'd136314880;
      41447: inst = 32'd268468224;
      41448: inst = 32'd201345088;
      41449: inst = 32'd203423744;
      41450: inst = 32'd471859200;
      41451: inst = 32'd136314880;
      41452: inst = 32'd268468224;
      41453: inst = 32'd201345089;
      41454: inst = 32'd203423744;
      41455: inst = 32'd471859200;
      41456: inst = 32'd136314880;
      41457: inst = 32'd268468224;
      41458: inst = 32'd201345090;
      41459: inst = 32'd203423744;
      41460: inst = 32'd471859200;
      41461: inst = 32'd136314880;
      41462: inst = 32'd268468224;
      41463: inst = 32'd201345091;
      41464: inst = 32'd203423744;
      41465: inst = 32'd471859200;
      41466: inst = 32'd136314880;
      41467: inst = 32'd268468224;
      41468: inst = 32'd201345092;
      41469: inst = 32'd203423744;
      41470: inst = 32'd471859200;
      41471: inst = 32'd136314880;
      41472: inst = 32'd268468224;
      41473: inst = 32'd201345093;
      41474: inst = 32'd203423744;
      41475: inst = 32'd471859200;
      41476: inst = 32'd136314880;
      41477: inst = 32'd268468224;
      41478: inst = 32'd201345094;
      41479: inst = 32'd203423744;
      41480: inst = 32'd471859200;
      41481: inst = 32'd136314880;
      41482: inst = 32'd268468224;
      41483: inst = 32'd201345095;
      41484: inst = 32'd203423744;
      41485: inst = 32'd471859200;
      41486: inst = 32'd136314880;
      41487: inst = 32'd268468224;
      41488: inst = 32'd201345096;
      41489: inst = 32'd203423744;
      41490: inst = 32'd471859200;
      41491: inst = 32'd136314880;
      41492: inst = 32'd268468224;
      41493: inst = 32'd201345097;
      41494: inst = 32'd203423744;
      41495: inst = 32'd471859200;
      41496: inst = 32'd136314880;
      41497: inst = 32'd268468224;
      41498: inst = 32'd201345098;
      41499: inst = 32'd203423744;
      41500: inst = 32'd471859200;
      41501: inst = 32'd136314880;
      41502: inst = 32'd268468224;
      41503: inst = 32'd201345099;
      41504: inst = 32'd203423744;
      41505: inst = 32'd471859200;
      41506: inst = 32'd136314880;
      41507: inst = 32'd268468224;
      41508: inst = 32'd201345100;
      41509: inst = 32'd203423744;
      41510: inst = 32'd471859200;
      41511: inst = 32'd136314880;
      41512: inst = 32'd268468224;
      41513: inst = 32'd201345101;
      41514: inst = 32'd203423744;
      41515: inst = 32'd471859200;
      41516: inst = 32'd136314880;
      41517: inst = 32'd268468224;
      41518: inst = 32'd201345102;
      41519: inst = 32'd203423744;
      41520: inst = 32'd471859200;
      41521: inst = 32'd136314880;
      41522: inst = 32'd268468224;
      41523: inst = 32'd201345103;
      41524: inst = 32'd203423744;
      41525: inst = 32'd471859200;
      41526: inst = 32'd136314880;
      41527: inst = 32'd268468224;
      41528: inst = 32'd201345104;
      41529: inst = 32'd203423744;
      41530: inst = 32'd471859200;
      41531: inst = 32'd136314880;
      41532: inst = 32'd268468224;
      41533: inst = 32'd201345105;
      41534: inst = 32'd203423744;
      41535: inst = 32'd471859200;
      41536: inst = 32'd136314880;
      41537: inst = 32'd268468224;
      41538: inst = 32'd201345106;
      41539: inst = 32'd203423744;
      41540: inst = 32'd471859200;
      41541: inst = 32'd136314880;
      41542: inst = 32'd268468224;
      41543: inst = 32'd201345107;
      41544: inst = 32'd203423744;
      41545: inst = 32'd471859200;
      41546: inst = 32'd136314880;
      41547: inst = 32'd268468224;
      41548: inst = 32'd201345108;
      41549: inst = 32'd203423744;
      41550: inst = 32'd471859200;
      41551: inst = 32'd136314880;
      41552: inst = 32'd268468224;
      41553: inst = 32'd201345109;
      41554: inst = 32'd203423744;
      41555: inst = 32'd471859200;
      41556: inst = 32'd136314880;
      41557: inst = 32'd268468224;
      41558: inst = 32'd201345110;
      41559: inst = 32'd203423744;
      41560: inst = 32'd471859200;
      41561: inst = 32'd136314880;
      41562: inst = 32'd268468224;
      41563: inst = 32'd201345111;
      41564: inst = 32'd203423744;
      41565: inst = 32'd471859200;
      41566: inst = 32'd136314880;
      41567: inst = 32'd268468224;
      41568: inst = 32'd201345112;
      41569: inst = 32'd203423744;
      41570: inst = 32'd471859200;
      41571: inst = 32'd136314880;
      41572: inst = 32'd268468224;
      41573: inst = 32'd201345113;
      41574: inst = 32'd203423744;
      41575: inst = 32'd471859200;
      41576: inst = 32'd136314880;
      41577: inst = 32'd268468224;
      41578: inst = 32'd201345114;
      41579: inst = 32'd203423744;
      41580: inst = 32'd471859200;
      41581: inst = 32'd136314880;
      41582: inst = 32'd268468224;
      41583: inst = 32'd201345115;
      41584: inst = 32'd203423744;
      41585: inst = 32'd471859200;
      41586: inst = 32'd136314880;
      41587: inst = 32'd268468224;
      41588: inst = 32'd201345116;
      41589: inst = 32'd203423744;
      41590: inst = 32'd471859200;
      41591: inst = 32'd136314880;
      41592: inst = 32'd268468224;
      41593: inst = 32'd201345117;
      41594: inst = 32'd203423744;
      41595: inst = 32'd471859200;
      41596: inst = 32'd136314880;
      41597: inst = 32'd268468224;
      41598: inst = 32'd201345118;
      41599: inst = 32'd203423744;
      41600: inst = 32'd471859200;
      41601: inst = 32'd136314880;
      41602: inst = 32'd268468224;
      41603: inst = 32'd201345119;
      41604: inst = 32'd203423744;
      41605: inst = 32'd471859200;
      41606: inst = 32'd136314880;
      41607: inst = 32'd268468224;
      41608: inst = 32'd201345120;
      41609: inst = 32'd203423744;
      41610: inst = 32'd471859200;
      41611: inst = 32'd136314880;
      41612: inst = 32'd268468224;
      41613: inst = 32'd201345121;
      41614: inst = 32'd203423744;
      41615: inst = 32'd471859200;
      41616: inst = 32'd136314880;
      41617: inst = 32'd268468224;
      41618: inst = 32'd201345122;
      41619: inst = 32'd203423744;
      41620: inst = 32'd471859200;
      41621: inst = 32'd136314880;
      41622: inst = 32'd268468224;
      41623: inst = 32'd201345123;
      41624: inst = 32'd203423744;
      41625: inst = 32'd471859200;
      41626: inst = 32'd136314880;
      41627: inst = 32'd268468224;
      41628: inst = 32'd201345124;
      41629: inst = 32'd203423744;
      41630: inst = 32'd471859200;
      41631: inst = 32'd136314880;
      41632: inst = 32'd268468224;
      41633: inst = 32'd201345125;
      41634: inst = 32'd203423744;
      41635: inst = 32'd471859200;
      41636: inst = 32'd136314880;
      41637: inst = 32'd268468224;
      41638: inst = 32'd201345126;
      41639: inst = 32'd203423744;
      41640: inst = 32'd471859200;
      41641: inst = 32'd136314880;
      41642: inst = 32'd268468224;
      41643: inst = 32'd201345127;
      41644: inst = 32'd203423744;
      41645: inst = 32'd471859200;
      41646: inst = 32'd136314880;
      41647: inst = 32'd268468224;
      41648: inst = 32'd201345128;
      41649: inst = 32'd203423744;
      41650: inst = 32'd471859200;
      41651: inst = 32'd136314880;
      41652: inst = 32'd268468224;
      41653: inst = 32'd201345129;
      41654: inst = 32'd203423744;
      41655: inst = 32'd471859200;
      41656: inst = 32'd136314880;
      41657: inst = 32'd268468224;
      41658: inst = 32'd201345130;
      41659: inst = 32'd203423744;
      41660: inst = 32'd471859200;
      41661: inst = 32'd136314880;
      41662: inst = 32'd268468224;
      41663: inst = 32'd201345131;
      41664: inst = 32'd203423744;
      41665: inst = 32'd471859200;
      41666: inst = 32'd136314880;
      41667: inst = 32'd268468224;
      41668: inst = 32'd201345132;
      41669: inst = 32'd203423744;
      41670: inst = 32'd471859200;
      41671: inst = 32'd136314880;
      41672: inst = 32'd268468224;
      41673: inst = 32'd201345133;
      41674: inst = 32'd203423744;
      41675: inst = 32'd471859200;
      41676: inst = 32'd136314880;
      41677: inst = 32'd268468224;
      41678: inst = 32'd201345134;
      41679: inst = 32'd203423744;
      41680: inst = 32'd471859200;
      41681: inst = 32'd136314880;
      41682: inst = 32'd268468224;
      41683: inst = 32'd201345135;
      41684: inst = 32'd203423744;
      41685: inst = 32'd471859200;
      41686: inst = 32'd136314880;
      41687: inst = 32'd268468224;
      41688: inst = 32'd201345136;
      41689: inst = 32'd203423744;
      41690: inst = 32'd471859200;
      41691: inst = 32'd136314880;
      41692: inst = 32'd268468224;
      41693: inst = 32'd201345137;
      41694: inst = 32'd203423744;
      41695: inst = 32'd471859200;
      41696: inst = 32'd136314880;
      41697: inst = 32'd268468224;
      41698: inst = 32'd201345138;
      41699: inst = 32'd203423744;
      41700: inst = 32'd471859200;
      41701: inst = 32'd136314880;
      41702: inst = 32'd268468224;
      41703: inst = 32'd201345139;
      41704: inst = 32'd203423744;
      41705: inst = 32'd471859200;
      41706: inst = 32'd136314880;
      41707: inst = 32'd268468224;
      41708: inst = 32'd201345140;
      41709: inst = 32'd203423744;
      41710: inst = 32'd471859200;
      41711: inst = 32'd136314880;
      41712: inst = 32'd268468224;
      41713: inst = 32'd201345141;
      41714: inst = 32'd203423744;
      41715: inst = 32'd471859200;
      41716: inst = 32'd136314880;
      41717: inst = 32'd268468224;
      41718: inst = 32'd201345142;
      41719: inst = 32'd203423744;
      41720: inst = 32'd471859200;
      41721: inst = 32'd136314880;
      41722: inst = 32'd268468224;
      41723: inst = 32'd201345143;
      41724: inst = 32'd203423744;
      41725: inst = 32'd471859200;
      41726: inst = 32'd136314880;
      41727: inst = 32'd268468224;
      41728: inst = 32'd201345144;
      41729: inst = 32'd203423744;
      41730: inst = 32'd471859200;
      41731: inst = 32'd136314880;
      41732: inst = 32'd268468224;
      41733: inst = 32'd201345145;
      41734: inst = 32'd203423744;
      41735: inst = 32'd471859200;
      41736: inst = 32'd136314880;
      41737: inst = 32'd268468224;
      41738: inst = 32'd201345146;
      41739: inst = 32'd203423744;
      41740: inst = 32'd471859200;
      41741: inst = 32'd136314880;
      41742: inst = 32'd268468224;
      41743: inst = 32'd201345147;
      41744: inst = 32'd203423744;
      41745: inst = 32'd471859200;
      41746: inst = 32'd136314880;
      41747: inst = 32'd268468224;
      41748: inst = 32'd201345148;
      41749: inst = 32'd203423744;
      41750: inst = 32'd471859200;
      41751: inst = 32'd136314880;
      41752: inst = 32'd268468224;
      41753: inst = 32'd201345149;
      41754: inst = 32'd203423744;
      41755: inst = 32'd471859200;
      41756: inst = 32'd136314880;
      41757: inst = 32'd268468224;
      41758: inst = 32'd201345150;
      41759: inst = 32'd203423744;
      41760: inst = 32'd471859200;
      41761: inst = 32'd136314880;
      41762: inst = 32'd268468224;
      41763: inst = 32'd201345151;
      41764: inst = 32'd203423744;
      41765: inst = 32'd471859200;
      41766: inst = 32'd136314880;
      41767: inst = 32'd268468224;
      41768: inst = 32'd201345152;
      41769: inst = 32'd203423744;
      41770: inst = 32'd471859200;
      41771: inst = 32'd136314880;
      41772: inst = 32'd268468224;
      41773: inst = 32'd201345153;
      41774: inst = 32'd203423744;
      41775: inst = 32'd471859200;
      41776: inst = 32'd136314880;
      41777: inst = 32'd268468224;
      41778: inst = 32'd201345154;
      41779: inst = 32'd203423744;
      41780: inst = 32'd471859200;
      41781: inst = 32'd136314880;
      41782: inst = 32'd268468224;
      41783: inst = 32'd201345155;
      41784: inst = 32'd203423744;
      41785: inst = 32'd471859200;
      41786: inst = 32'd136314880;
      41787: inst = 32'd268468224;
      41788: inst = 32'd201345156;
      41789: inst = 32'd203423744;
      41790: inst = 32'd471859200;
      41791: inst = 32'd136314880;
      41792: inst = 32'd268468224;
      41793: inst = 32'd201345157;
      41794: inst = 32'd203423744;
      41795: inst = 32'd471859200;
      41796: inst = 32'd136314880;
      41797: inst = 32'd268468224;
      41798: inst = 32'd201345158;
      41799: inst = 32'd203423744;
      41800: inst = 32'd471859200;
      41801: inst = 32'd136314880;
      41802: inst = 32'd268468224;
      41803: inst = 32'd201345159;
      41804: inst = 32'd203423744;
      41805: inst = 32'd471859200;
      41806: inst = 32'd136314880;
      41807: inst = 32'd268468224;
      41808: inst = 32'd201345160;
      41809: inst = 32'd203423744;
      41810: inst = 32'd471859200;
      41811: inst = 32'd136314880;
      41812: inst = 32'd268468224;
      41813: inst = 32'd201345161;
      41814: inst = 32'd203423744;
      41815: inst = 32'd471859200;
      41816: inst = 32'd136314880;
      41817: inst = 32'd268468224;
      41818: inst = 32'd201345162;
      41819: inst = 32'd203423744;
      41820: inst = 32'd471859200;
      41821: inst = 32'd136314880;
      41822: inst = 32'd268468224;
      41823: inst = 32'd201345163;
      41824: inst = 32'd203423744;
      41825: inst = 32'd471859200;
      41826: inst = 32'd136314880;
      41827: inst = 32'd268468224;
      41828: inst = 32'd201345164;
      41829: inst = 32'd203423744;
      41830: inst = 32'd471859200;
      41831: inst = 32'd136314880;
      41832: inst = 32'd268468224;
      41833: inst = 32'd201345165;
      41834: inst = 32'd203423744;
      41835: inst = 32'd471859200;
      41836: inst = 32'd136314880;
      41837: inst = 32'd268468224;
      41838: inst = 32'd201345166;
      41839: inst = 32'd203423744;
      41840: inst = 32'd471859200;
      41841: inst = 32'd136314880;
      41842: inst = 32'd268468224;
      41843: inst = 32'd201345167;
      41844: inst = 32'd203423744;
      41845: inst = 32'd471859200;
      41846: inst = 32'd136314880;
      41847: inst = 32'd268468224;
      41848: inst = 32'd201345168;
      41849: inst = 32'd203423744;
      41850: inst = 32'd471859200;
      41851: inst = 32'd136314880;
      41852: inst = 32'd268468224;
      41853: inst = 32'd201345169;
      41854: inst = 32'd203423744;
      41855: inst = 32'd471859200;
      41856: inst = 32'd136314880;
      41857: inst = 32'd268468224;
      41858: inst = 32'd201345170;
      41859: inst = 32'd203423744;
      41860: inst = 32'd471859200;
      41861: inst = 32'd136314880;
      41862: inst = 32'd268468224;
      41863: inst = 32'd201345171;
      41864: inst = 32'd203423744;
      41865: inst = 32'd471859200;
      41866: inst = 32'd136314880;
      41867: inst = 32'd268468224;
      41868: inst = 32'd201345172;
      41869: inst = 32'd203423744;
      41870: inst = 32'd471859200;
      41871: inst = 32'd136314880;
      41872: inst = 32'd268468224;
      41873: inst = 32'd201345173;
      41874: inst = 32'd203423744;
      41875: inst = 32'd471859200;
      41876: inst = 32'd136314880;
      41877: inst = 32'd268468224;
      41878: inst = 32'd201345174;
      41879: inst = 32'd203423744;
      41880: inst = 32'd471859200;
      41881: inst = 32'd136314880;
      41882: inst = 32'd268468224;
      41883: inst = 32'd201345175;
      41884: inst = 32'd203423744;
      41885: inst = 32'd471859200;
      41886: inst = 32'd136314880;
      41887: inst = 32'd268468224;
      41888: inst = 32'd201345176;
      41889: inst = 32'd203423744;
      41890: inst = 32'd471859200;
      41891: inst = 32'd136314880;
      41892: inst = 32'd268468224;
      41893: inst = 32'd201345177;
      41894: inst = 32'd203423744;
      41895: inst = 32'd471859200;
      41896: inst = 32'd136314880;
      41897: inst = 32'd268468224;
      41898: inst = 32'd201345178;
      41899: inst = 32'd203423744;
      41900: inst = 32'd471859200;
      41901: inst = 32'd136314880;
      41902: inst = 32'd268468224;
      41903: inst = 32'd201345179;
      41904: inst = 32'd203423744;
      41905: inst = 32'd471859200;
      41906: inst = 32'd136314880;
      41907: inst = 32'd268468224;
      41908: inst = 32'd201345180;
      41909: inst = 32'd203423744;
      41910: inst = 32'd471859200;
      41911: inst = 32'd136314880;
      41912: inst = 32'd268468224;
      41913: inst = 32'd201345181;
      41914: inst = 32'd203423744;
      41915: inst = 32'd471859200;
      41916: inst = 32'd136314880;
      41917: inst = 32'd268468224;
      41918: inst = 32'd201345182;
      41919: inst = 32'd203423744;
      41920: inst = 32'd471859200;
      41921: inst = 32'd136314880;
      41922: inst = 32'd268468224;
      41923: inst = 32'd201345183;
      41924: inst = 32'd203423744;
      41925: inst = 32'd471859200;
      41926: inst = 32'd136314880;
      41927: inst = 32'd268468224;
      41928: inst = 32'd201345184;
      41929: inst = 32'd203423744;
      41930: inst = 32'd471859200;
      41931: inst = 32'd136314880;
      41932: inst = 32'd268468224;
      41933: inst = 32'd201345185;
      41934: inst = 32'd203423744;
      41935: inst = 32'd471859200;
      41936: inst = 32'd136314880;
      41937: inst = 32'd268468224;
      41938: inst = 32'd201345186;
      41939: inst = 32'd203423744;
      41940: inst = 32'd471859200;
      41941: inst = 32'd136314880;
      41942: inst = 32'd268468224;
      41943: inst = 32'd201345187;
      41944: inst = 32'd203423744;
      41945: inst = 32'd471859200;
      41946: inst = 32'd136314880;
      41947: inst = 32'd268468224;
      41948: inst = 32'd201345188;
      41949: inst = 32'd203423744;
      41950: inst = 32'd471859200;
      41951: inst = 32'd136314880;
      41952: inst = 32'd268468224;
      41953: inst = 32'd201345189;
      41954: inst = 32'd203423744;
      41955: inst = 32'd471859200;
      41956: inst = 32'd136314880;
      41957: inst = 32'd268468224;
      41958: inst = 32'd201345190;
      41959: inst = 32'd203423744;
      41960: inst = 32'd471859200;
      41961: inst = 32'd136314880;
      41962: inst = 32'd268468224;
      41963: inst = 32'd201345191;
      41964: inst = 32'd203423744;
      41965: inst = 32'd471859200;
      41966: inst = 32'd136314880;
      41967: inst = 32'd268468224;
      41968: inst = 32'd201345192;
      41969: inst = 32'd203423744;
      41970: inst = 32'd471859200;
      41971: inst = 32'd136314880;
      41972: inst = 32'd268468224;
      41973: inst = 32'd201345193;
      41974: inst = 32'd203423744;
      41975: inst = 32'd471859200;
      41976: inst = 32'd136314880;
      41977: inst = 32'd268468224;
      41978: inst = 32'd201345194;
      41979: inst = 32'd203423744;
      41980: inst = 32'd471859200;
      41981: inst = 32'd136314880;
      41982: inst = 32'd268468224;
      41983: inst = 32'd201345195;
      41984: inst = 32'd203423744;
      41985: inst = 32'd471859200;
      41986: inst = 32'd136314880;
      41987: inst = 32'd268468224;
      41988: inst = 32'd201345196;
      41989: inst = 32'd203423744;
      41990: inst = 32'd471859200;
      41991: inst = 32'd136314880;
      41992: inst = 32'd268468224;
      41993: inst = 32'd201345197;
      41994: inst = 32'd203423744;
      41995: inst = 32'd471859200;
      41996: inst = 32'd136314880;
      41997: inst = 32'd268468224;
      41998: inst = 32'd201345198;
      41999: inst = 32'd203423744;
      42000: inst = 32'd471859200;
      42001: inst = 32'd136314880;
      42002: inst = 32'd268468224;
      42003: inst = 32'd201345199;
      42004: inst = 32'd203423744;
      42005: inst = 32'd471859200;
      42006: inst = 32'd136314880;
      42007: inst = 32'd268468224;
      42008: inst = 32'd201345200;
      42009: inst = 32'd203423744;
      42010: inst = 32'd471859200;
      42011: inst = 32'd136314880;
      42012: inst = 32'd268468224;
      42013: inst = 32'd201345201;
      42014: inst = 32'd203423744;
      42015: inst = 32'd471859200;
      42016: inst = 32'd136314880;
      42017: inst = 32'd268468224;
      42018: inst = 32'd201345202;
      42019: inst = 32'd203423744;
      42020: inst = 32'd471859200;
      42021: inst = 32'd136314880;
      42022: inst = 32'd268468224;
      42023: inst = 32'd201345203;
      42024: inst = 32'd203423744;
      42025: inst = 32'd471859200;
      42026: inst = 32'd136314880;
      42027: inst = 32'd268468224;
      42028: inst = 32'd201345204;
      42029: inst = 32'd203423744;
      42030: inst = 32'd471859200;
      42031: inst = 32'd136314880;
      42032: inst = 32'd268468224;
      42033: inst = 32'd201345205;
      42034: inst = 32'd203423744;
      42035: inst = 32'd471859200;
      42036: inst = 32'd136314880;
      42037: inst = 32'd268468224;
      42038: inst = 32'd201345206;
      42039: inst = 32'd203423744;
      42040: inst = 32'd471859200;
      42041: inst = 32'd136314880;
      42042: inst = 32'd268468224;
      42043: inst = 32'd201345207;
      42044: inst = 32'd203423744;
      42045: inst = 32'd471859200;
      42046: inst = 32'd136314880;
      42047: inst = 32'd268468224;
      42048: inst = 32'd201345208;
      42049: inst = 32'd203423744;
      42050: inst = 32'd471859200;
      42051: inst = 32'd136314880;
      42052: inst = 32'd268468224;
      42053: inst = 32'd201345209;
      42054: inst = 32'd203423744;
      42055: inst = 32'd471859200;
      42056: inst = 32'd136314880;
      42057: inst = 32'd268468224;
      42058: inst = 32'd201345210;
      42059: inst = 32'd203423744;
      42060: inst = 32'd471859200;
      42061: inst = 32'd136314880;
      42062: inst = 32'd268468224;
      42063: inst = 32'd201345211;
      42064: inst = 32'd203423744;
      42065: inst = 32'd471859200;
      42066: inst = 32'd136314880;
      42067: inst = 32'd268468224;
      42068: inst = 32'd201345212;
      42069: inst = 32'd203423744;
      42070: inst = 32'd471859200;
      42071: inst = 32'd136314880;
      42072: inst = 32'd268468224;
      42073: inst = 32'd201345213;
      42074: inst = 32'd203423744;
      42075: inst = 32'd471859200;
      42076: inst = 32'd136314880;
      42077: inst = 32'd268468224;
      42078: inst = 32'd201345214;
      42079: inst = 32'd203423744;
      42080: inst = 32'd471859200;
      42081: inst = 32'd136314880;
      42082: inst = 32'd268468224;
      42083: inst = 32'd201345215;
      42084: inst = 32'd203423744;
      42085: inst = 32'd471859200;
      42086: inst = 32'd136314880;
      42087: inst = 32'd268468224;
      42088: inst = 32'd201345216;
      42089: inst = 32'd203423744;
      42090: inst = 32'd471859200;
      42091: inst = 32'd136314880;
      42092: inst = 32'd268468224;
      42093: inst = 32'd201345217;
      42094: inst = 32'd203423744;
      42095: inst = 32'd471859200;
      42096: inst = 32'd136314880;
      42097: inst = 32'd268468224;
      42098: inst = 32'd201345218;
      42099: inst = 32'd203423744;
      42100: inst = 32'd471859200;
      42101: inst = 32'd136314880;
      42102: inst = 32'd268468224;
      42103: inst = 32'd201345219;
      42104: inst = 32'd203423744;
      42105: inst = 32'd471859200;
      42106: inst = 32'd136314880;
      42107: inst = 32'd268468224;
      42108: inst = 32'd201345220;
      42109: inst = 32'd203423744;
      42110: inst = 32'd471859200;
      42111: inst = 32'd136314880;
      42112: inst = 32'd268468224;
      42113: inst = 32'd201345221;
      42114: inst = 32'd203423744;
      42115: inst = 32'd471859200;
      42116: inst = 32'd136314880;
      42117: inst = 32'd268468224;
      42118: inst = 32'd201345222;
      42119: inst = 32'd203423744;
      42120: inst = 32'd471859200;
      42121: inst = 32'd136314880;
      42122: inst = 32'd268468224;
      42123: inst = 32'd201345223;
      42124: inst = 32'd203423744;
      42125: inst = 32'd471859200;
      42126: inst = 32'd136314880;
      42127: inst = 32'd268468224;
      42128: inst = 32'd201345224;
      42129: inst = 32'd203423744;
      42130: inst = 32'd471859200;
      42131: inst = 32'd136314880;
      42132: inst = 32'd268468224;
      42133: inst = 32'd201345225;
      42134: inst = 32'd203423744;
      42135: inst = 32'd471859200;
      42136: inst = 32'd136314880;
      42137: inst = 32'd268468224;
      42138: inst = 32'd201345226;
      42139: inst = 32'd203423744;
      42140: inst = 32'd471859200;
      42141: inst = 32'd136314880;
      42142: inst = 32'd268468224;
      42143: inst = 32'd201345227;
      42144: inst = 32'd203423744;
      42145: inst = 32'd471859200;
      42146: inst = 32'd136314880;
      42147: inst = 32'd268468224;
      42148: inst = 32'd201345228;
      42149: inst = 32'd203423744;
      42150: inst = 32'd471859200;
      42151: inst = 32'd136314880;
      42152: inst = 32'd268468224;
      42153: inst = 32'd201345229;
      42154: inst = 32'd203423744;
      42155: inst = 32'd471859200;
      42156: inst = 32'd136314880;
      42157: inst = 32'd268468224;
      42158: inst = 32'd201345230;
      42159: inst = 32'd203423744;
      42160: inst = 32'd471859200;
      42161: inst = 32'd136314880;
      42162: inst = 32'd268468224;
      42163: inst = 32'd201345231;
      42164: inst = 32'd203423744;
      42165: inst = 32'd471859200;
      42166: inst = 32'd136314880;
      42167: inst = 32'd268468224;
      42168: inst = 32'd201345232;
      42169: inst = 32'd203423744;
      42170: inst = 32'd471859200;
      42171: inst = 32'd136314880;
      42172: inst = 32'd268468224;
      42173: inst = 32'd201345233;
      42174: inst = 32'd203423744;
      42175: inst = 32'd471859200;
      42176: inst = 32'd136314880;
      42177: inst = 32'd268468224;
      42178: inst = 32'd201345234;
      42179: inst = 32'd203423744;
      42180: inst = 32'd471859200;
      42181: inst = 32'd136314880;
      42182: inst = 32'd268468224;
      42183: inst = 32'd201345235;
      42184: inst = 32'd203423744;
      42185: inst = 32'd471859200;
      42186: inst = 32'd136314880;
      42187: inst = 32'd268468224;
      42188: inst = 32'd201345236;
      42189: inst = 32'd203423744;
      42190: inst = 32'd471859200;
      42191: inst = 32'd136314880;
      42192: inst = 32'd268468224;
      42193: inst = 32'd201345237;
      42194: inst = 32'd203423744;
      42195: inst = 32'd471859200;
      42196: inst = 32'd136314880;
      42197: inst = 32'd268468224;
      42198: inst = 32'd201345238;
      42199: inst = 32'd203423744;
      42200: inst = 32'd471859200;
      42201: inst = 32'd136314880;
      42202: inst = 32'd268468224;
      42203: inst = 32'd201345239;
      42204: inst = 32'd203423744;
      42205: inst = 32'd471859200;
      42206: inst = 32'd136314880;
      42207: inst = 32'd268468224;
      42208: inst = 32'd201345240;
      42209: inst = 32'd203423744;
      42210: inst = 32'd471859200;
      42211: inst = 32'd136314880;
      42212: inst = 32'd268468224;
      42213: inst = 32'd201345241;
      42214: inst = 32'd203423744;
      42215: inst = 32'd471859200;
      42216: inst = 32'd136314880;
      42217: inst = 32'd268468224;
      42218: inst = 32'd201345242;
      42219: inst = 32'd203423744;
      42220: inst = 32'd471859200;
      42221: inst = 32'd136314880;
      42222: inst = 32'd268468224;
      42223: inst = 32'd201345243;
      42224: inst = 32'd203423744;
      42225: inst = 32'd471859200;
      42226: inst = 32'd136314880;
      42227: inst = 32'd268468224;
      42228: inst = 32'd201345244;
      42229: inst = 32'd203423744;
      42230: inst = 32'd471859200;
      42231: inst = 32'd136314880;
      42232: inst = 32'd268468224;
      42233: inst = 32'd201345245;
      42234: inst = 32'd203423744;
      42235: inst = 32'd471859200;
      42236: inst = 32'd136314880;
      42237: inst = 32'd268468224;
      42238: inst = 32'd201345246;
      42239: inst = 32'd203423744;
      42240: inst = 32'd471859200;
      42241: inst = 32'd136314880;
      42242: inst = 32'd268468224;
      42243: inst = 32'd201345247;
      42244: inst = 32'd203423744;
      42245: inst = 32'd471859200;
      42246: inst = 32'd136314880;
      42247: inst = 32'd268468224;
      42248: inst = 32'd201345248;
      42249: inst = 32'd203423744;
      42250: inst = 32'd471859200;
      42251: inst = 32'd136314880;
      42252: inst = 32'd268468224;
      42253: inst = 32'd201345249;
      42254: inst = 32'd203423744;
      42255: inst = 32'd471859200;
      42256: inst = 32'd136314880;
      42257: inst = 32'd268468224;
      42258: inst = 32'd201345250;
      42259: inst = 32'd203423744;
      42260: inst = 32'd471859200;
      42261: inst = 32'd136314880;
      42262: inst = 32'd268468224;
      42263: inst = 32'd201345251;
      42264: inst = 32'd203423744;
      42265: inst = 32'd471859200;
      42266: inst = 32'd136314880;
      42267: inst = 32'd268468224;
      42268: inst = 32'd201345252;
      42269: inst = 32'd203423744;
      42270: inst = 32'd471859200;
      42271: inst = 32'd136314880;
      42272: inst = 32'd268468224;
      42273: inst = 32'd201345253;
      42274: inst = 32'd203423744;
      42275: inst = 32'd471859200;
      42276: inst = 32'd136314880;
      42277: inst = 32'd268468224;
      42278: inst = 32'd201345254;
      42279: inst = 32'd203423744;
      42280: inst = 32'd471859200;
      42281: inst = 32'd136314880;
      42282: inst = 32'd268468224;
      42283: inst = 32'd201345255;
      42284: inst = 32'd203423744;
      42285: inst = 32'd471859200;
      42286: inst = 32'd136314880;
      42287: inst = 32'd268468224;
      42288: inst = 32'd201345256;
      42289: inst = 32'd203423744;
      42290: inst = 32'd471859200;
      42291: inst = 32'd136314880;
      42292: inst = 32'd268468224;
      42293: inst = 32'd201345257;
      42294: inst = 32'd203423744;
      42295: inst = 32'd471859200;
      42296: inst = 32'd136314880;
      42297: inst = 32'd268468224;
      42298: inst = 32'd201345258;
      42299: inst = 32'd203423744;
      42300: inst = 32'd471859200;
      42301: inst = 32'd136314880;
      42302: inst = 32'd268468224;
      42303: inst = 32'd201345259;
      42304: inst = 32'd203423744;
      42305: inst = 32'd471859200;
      42306: inst = 32'd136314880;
      42307: inst = 32'd268468224;
      42308: inst = 32'd201345260;
      42309: inst = 32'd203423744;
      42310: inst = 32'd471859200;
      42311: inst = 32'd136314880;
      42312: inst = 32'd268468224;
      42313: inst = 32'd201345261;
      42314: inst = 32'd203423744;
      42315: inst = 32'd471859200;
      42316: inst = 32'd136314880;
      42317: inst = 32'd268468224;
      42318: inst = 32'd201345262;
      42319: inst = 32'd203423744;
      42320: inst = 32'd471859200;
      42321: inst = 32'd136314880;
      42322: inst = 32'd268468224;
      42323: inst = 32'd201345263;
      42324: inst = 32'd203423744;
      42325: inst = 32'd471859200;
      42326: inst = 32'd136314880;
      42327: inst = 32'd268468224;
      42328: inst = 32'd201345264;
      42329: inst = 32'd203423744;
      42330: inst = 32'd471859200;
      42331: inst = 32'd136314880;
      42332: inst = 32'd268468224;
      42333: inst = 32'd201345265;
      42334: inst = 32'd203423744;
      42335: inst = 32'd471859200;
      42336: inst = 32'd136314880;
      42337: inst = 32'd268468224;
      42338: inst = 32'd201345266;
      42339: inst = 32'd203423744;
      42340: inst = 32'd471859200;
      42341: inst = 32'd136314880;
      42342: inst = 32'd268468224;
      42343: inst = 32'd201345267;
      42344: inst = 32'd203423744;
      42345: inst = 32'd471859200;
      42346: inst = 32'd136314880;
      42347: inst = 32'd268468224;
      42348: inst = 32'd201345268;
      42349: inst = 32'd203423744;
      42350: inst = 32'd471859200;
      42351: inst = 32'd136314880;
      42352: inst = 32'd268468224;
      42353: inst = 32'd201345269;
      42354: inst = 32'd203423744;
      42355: inst = 32'd471859200;
      42356: inst = 32'd136314880;
      42357: inst = 32'd268468224;
      42358: inst = 32'd201345270;
      42359: inst = 32'd203423744;
      42360: inst = 32'd471859200;
      42361: inst = 32'd136314880;
      42362: inst = 32'd268468224;
      42363: inst = 32'd201345271;
      42364: inst = 32'd203423744;
      42365: inst = 32'd471859200;
      42366: inst = 32'd136314880;
      42367: inst = 32'd268468224;
      42368: inst = 32'd201345272;
      42369: inst = 32'd203423744;
      42370: inst = 32'd471859200;
      42371: inst = 32'd136314880;
      42372: inst = 32'd268468224;
      42373: inst = 32'd201345273;
      42374: inst = 32'd203423744;
      42375: inst = 32'd471859200;
      42376: inst = 32'd136314880;
      42377: inst = 32'd268468224;
      42378: inst = 32'd201345274;
      42379: inst = 32'd203423744;
      42380: inst = 32'd471859200;
      42381: inst = 32'd136314880;
      42382: inst = 32'd268468224;
      42383: inst = 32'd201345275;
      42384: inst = 32'd203423744;
      42385: inst = 32'd471859200;
      42386: inst = 32'd136314880;
      42387: inst = 32'd268468224;
      42388: inst = 32'd201345276;
      42389: inst = 32'd203423744;
      42390: inst = 32'd471859200;
      42391: inst = 32'd136314880;
      42392: inst = 32'd268468224;
      42393: inst = 32'd201345277;
      42394: inst = 32'd203423744;
      42395: inst = 32'd471859200;
      42396: inst = 32'd136314880;
      42397: inst = 32'd268468224;
      42398: inst = 32'd201345278;
      42399: inst = 32'd203423744;
      42400: inst = 32'd471859200;
      42401: inst = 32'd136314880;
      42402: inst = 32'd268468224;
      42403: inst = 32'd201345279;
      42404: inst = 32'd203423744;
      42405: inst = 32'd471859200;
      42406: inst = 32'd136314880;
      42407: inst = 32'd268468224;
      42408: inst = 32'd201345280;
      42409: inst = 32'd203423744;
      42410: inst = 32'd471859200;
      42411: inst = 32'd136314880;
      42412: inst = 32'd268468224;
      42413: inst = 32'd201345281;
      42414: inst = 32'd203423744;
      42415: inst = 32'd471859200;
      42416: inst = 32'd136314880;
      42417: inst = 32'd268468224;
      42418: inst = 32'd201345282;
      42419: inst = 32'd203423744;
      42420: inst = 32'd471859200;
      42421: inst = 32'd136314880;
      42422: inst = 32'd268468224;
      42423: inst = 32'd201345283;
      42424: inst = 32'd203423744;
      42425: inst = 32'd471859200;
      42426: inst = 32'd136314880;
      42427: inst = 32'd268468224;
      42428: inst = 32'd201345284;
      42429: inst = 32'd203423744;
      42430: inst = 32'd471859200;
      42431: inst = 32'd136314880;
      42432: inst = 32'd268468224;
      42433: inst = 32'd201345285;
      42434: inst = 32'd203423744;
      42435: inst = 32'd471859200;
      42436: inst = 32'd136314880;
      42437: inst = 32'd268468224;
      42438: inst = 32'd201345286;
      42439: inst = 32'd203423744;
      42440: inst = 32'd471859200;
      42441: inst = 32'd136314880;
      42442: inst = 32'd268468224;
      42443: inst = 32'd201345287;
      42444: inst = 32'd203423744;
      42445: inst = 32'd471859200;
      42446: inst = 32'd136314880;
      42447: inst = 32'd268468224;
      42448: inst = 32'd201345288;
      42449: inst = 32'd203423744;
      42450: inst = 32'd471859200;
      42451: inst = 32'd136314880;
      42452: inst = 32'd268468224;
      42453: inst = 32'd201345289;
      42454: inst = 32'd203423744;
      42455: inst = 32'd471859200;
      42456: inst = 32'd136314880;
      42457: inst = 32'd268468224;
      42458: inst = 32'd201345290;
      42459: inst = 32'd203423744;
      42460: inst = 32'd471859200;
      42461: inst = 32'd136314880;
      42462: inst = 32'd268468224;
      42463: inst = 32'd201345291;
      42464: inst = 32'd203423744;
      42465: inst = 32'd471859200;
      42466: inst = 32'd136314880;
      42467: inst = 32'd268468224;
      42468: inst = 32'd201345292;
      42469: inst = 32'd203423744;
      42470: inst = 32'd471859200;
      42471: inst = 32'd136314880;
      42472: inst = 32'd268468224;
      42473: inst = 32'd201345293;
      42474: inst = 32'd203423744;
      42475: inst = 32'd471859200;
      42476: inst = 32'd136314880;
      42477: inst = 32'd268468224;
      42478: inst = 32'd201345294;
      42479: inst = 32'd203423744;
      42480: inst = 32'd471859200;
      42481: inst = 32'd136314880;
      42482: inst = 32'd268468224;
      42483: inst = 32'd201345295;
      42484: inst = 32'd203423744;
      42485: inst = 32'd471859200;
      42486: inst = 32'd136314880;
      42487: inst = 32'd268468224;
      42488: inst = 32'd201345296;
      42489: inst = 32'd203423744;
      42490: inst = 32'd471859200;
      42491: inst = 32'd136314880;
      42492: inst = 32'd268468224;
      42493: inst = 32'd201345297;
      42494: inst = 32'd203423744;
      42495: inst = 32'd471859200;
      42496: inst = 32'd136314880;
      42497: inst = 32'd268468224;
      42498: inst = 32'd201345298;
      42499: inst = 32'd203423744;
      42500: inst = 32'd471859200;
      42501: inst = 32'd136314880;
      42502: inst = 32'd268468224;
      42503: inst = 32'd201345299;
      42504: inst = 32'd203423744;
      42505: inst = 32'd471859200;
      42506: inst = 32'd136314880;
      42507: inst = 32'd268468224;
      42508: inst = 32'd201345300;
      42509: inst = 32'd203423744;
      42510: inst = 32'd471859200;
      42511: inst = 32'd136314880;
      42512: inst = 32'd268468224;
      42513: inst = 32'd201345301;
      42514: inst = 32'd203423744;
      42515: inst = 32'd471859200;
      42516: inst = 32'd136314880;
      42517: inst = 32'd268468224;
      42518: inst = 32'd201345302;
      42519: inst = 32'd203423744;
      42520: inst = 32'd471859200;
      42521: inst = 32'd136314880;
      42522: inst = 32'd268468224;
      42523: inst = 32'd201345303;
      42524: inst = 32'd203423744;
      42525: inst = 32'd471859200;
      42526: inst = 32'd136314880;
      42527: inst = 32'd268468224;
      42528: inst = 32'd201345304;
      42529: inst = 32'd203423744;
      42530: inst = 32'd471859200;
      42531: inst = 32'd136314880;
      42532: inst = 32'd268468224;
      42533: inst = 32'd201345305;
      42534: inst = 32'd203423744;
      42535: inst = 32'd471859200;
      42536: inst = 32'd136314880;
      42537: inst = 32'd268468224;
      42538: inst = 32'd201345306;
      42539: inst = 32'd203423744;
      42540: inst = 32'd471859200;
      42541: inst = 32'd136314880;
      42542: inst = 32'd268468224;
      42543: inst = 32'd201345307;
      42544: inst = 32'd203423744;
      42545: inst = 32'd471859200;
      42546: inst = 32'd136314880;
      42547: inst = 32'd268468224;
      42548: inst = 32'd201345308;
      42549: inst = 32'd203423744;
      42550: inst = 32'd471859200;
      42551: inst = 32'd136314880;
      42552: inst = 32'd268468224;
      42553: inst = 32'd201345309;
      42554: inst = 32'd203423744;
      42555: inst = 32'd471859200;
      42556: inst = 32'd136314880;
      42557: inst = 32'd268468224;
      42558: inst = 32'd201345310;
      42559: inst = 32'd203423744;
      42560: inst = 32'd471859200;
      42561: inst = 32'd136314880;
      42562: inst = 32'd268468224;
      42563: inst = 32'd201345311;
      42564: inst = 32'd203423744;
      42565: inst = 32'd471859200;
      42566: inst = 32'd136314880;
      42567: inst = 32'd268468224;
      42568: inst = 32'd201345312;
      42569: inst = 32'd203423744;
      42570: inst = 32'd471859200;
      42571: inst = 32'd136314880;
      42572: inst = 32'd268468224;
      42573: inst = 32'd201345313;
      42574: inst = 32'd203423744;
      42575: inst = 32'd471859200;
      42576: inst = 32'd136314880;
      42577: inst = 32'd268468224;
      42578: inst = 32'd201345314;
      42579: inst = 32'd203423744;
      42580: inst = 32'd471859200;
      42581: inst = 32'd136314880;
      42582: inst = 32'd268468224;
      42583: inst = 32'd201345315;
      42584: inst = 32'd203423744;
      42585: inst = 32'd471859200;
      42586: inst = 32'd136314880;
      42587: inst = 32'd268468224;
      42588: inst = 32'd201345316;
      42589: inst = 32'd203423744;
      42590: inst = 32'd471859200;
      42591: inst = 32'd136314880;
      42592: inst = 32'd268468224;
      42593: inst = 32'd201345317;
      42594: inst = 32'd203423744;
      42595: inst = 32'd471859200;
      42596: inst = 32'd136314880;
      42597: inst = 32'd268468224;
      42598: inst = 32'd201345318;
      42599: inst = 32'd203423744;
      42600: inst = 32'd471859200;
      42601: inst = 32'd136314880;
      42602: inst = 32'd268468224;
      42603: inst = 32'd201345319;
      42604: inst = 32'd203423744;
      42605: inst = 32'd471859200;
      42606: inst = 32'd136314880;
      42607: inst = 32'd268468224;
      42608: inst = 32'd201345320;
      42609: inst = 32'd203423744;
      42610: inst = 32'd471859200;
      42611: inst = 32'd136314880;
      42612: inst = 32'd268468224;
      42613: inst = 32'd201345321;
      42614: inst = 32'd203423744;
      42615: inst = 32'd471859200;
      42616: inst = 32'd136314880;
      42617: inst = 32'd268468224;
      42618: inst = 32'd201345322;
      42619: inst = 32'd203423744;
      42620: inst = 32'd471859200;
      42621: inst = 32'd136314880;
      42622: inst = 32'd268468224;
      42623: inst = 32'd201345323;
      42624: inst = 32'd203423744;
      42625: inst = 32'd471859200;
      42626: inst = 32'd136314880;
      42627: inst = 32'd268468224;
      42628: inst = 32'd201345324;
      42629: inst = 32'd203423744;
      42630: inst = 32'd471859200;
      42631: inst = 32'd136314880;
      42632: inst = 32'd268468224;
      42633: inst = 32'd201345325;
      42634: inst = 32'd203423744;
      42635: inst = 32'd471859200;
      42636: inst = 32'd136314880;
      42637: inst = 32'd268468224;
      42638: inst = 32'd201345326;
      42639: inst = 32'd203423744;
      42640: inst = 32'd471859200;
      42641: inst = 32'd136314880;
      42642: inst = 32'd268468224;
      42643: inst = 32'd201345327;
      42644: inst = 32'd203423744;
      42645: inst = 32'd471859200;
      42646: inst = 32'd136314880;
      42647: inst = 32'd268468224;
      42648: inst = 32'd201345328;
      42649: inst = 32'd203423744;
      42650: inst = 32'd471859200;
      42651: inst = 32'd136314880;
      42652: inst = 32'd268468224;
      42653: inst = 32'd201345329;
      42654: inst = 32'd203423744;
      42655: inst = 32'd471859200;
      42656: inst = 32'd136314880;
      42657: inst = 32'd268468224;
      42658: inst = 32'd201345330;
      42659: inst = 32'd203423744;
      42660: inst = 32'd471859200;
      42661: inst = 32'd136314880;
      42662: inst = 32'd268468224;
      42663: inst = 32'd201345331;
      42664: inst = 32'd203423744;
      42665: inst = 32'd471859200;
      42666: inst = 32'd136314880;
      42667: inst = 32'd268468224;
      42668: inst = 32'd201345332;
      42669: inst = 32'd203423744;
      42670: inst = 32'd471859200;
      42671: inst = 32'd136314880;
      42672: inst = 32'd268468224;
      42673: inst = 32'd201345333;
      42674: inst = 32'd203423744;
      42675: inst = 32'd471859200;
      42676: inst = 32'd136314880;
      42677: inst = 32'd268468224;
      42678: inst = 32'd201345334;
      42679: inst = 32'd203423744;
      42680: inst = 32'd471859200;
      42681: inst = 32'd136314880;
      42682: inst = 32'd268468224;
      42683: inst = 32'd201345335;
      42684: inst = 32'd203423744;
      42685: inst = 32'd471859200;
      42686: inst = 32'd136314880;
      42687: inst = 32'd268468224;
      42688: inst = 32'd201345336;
      42689: inst = 32'd203423744;
      42690: inst = 32'd471859200;
      42691: inst = 32'd136314880;
      42692: inst = 32'd268468224;
      42693: inst = 32'd201345337;
      42694: inst = 32'd203423744;
      42695: inst = 32'd471859200;
      42696: inst = 32'd136314880;
      42697: inst = 32'd268468224;
      42698: inst = 32'd201345338;
      42699: inst = 32'd203423744;
      42700: inst = 32'd471859200;
      42701: inst = 32'd136314880;
      42702: inst = 32'd268468224;
      42703: inst = 32'd201345339;
      42704: inst = 32'd203423744;
      42705: inst = 32'd471859200;
      42706: inst = 32'd136314880;
      42707: inst = 32'd268468224;
      42708: inst = 32'd201345340;
      42709: inst = 32'd203423744;
      42710: inst = 32'd471859200;
      42711: inst = 32'd136314880;
      42712: inst = 32'd268468224;
      42713: inst = 32'd201345341;
      42714: inst = 32'd203423744;
      42715: inst = 32'd471859200;
      42716: inst = 32'd136314880;
      42717: inst = 32'd268468224;
      42718: inst = 32'd201345342;
      42719: inst = 32'd203423744;
      42720: inst = 32'd471859200;
      42721: inst = 32'd136314880;
      42722: inst = 32'd268468224;
      42723: inst = 32'd201345343;
      42724: inst = 32'd203423744;
      42725: inst = 32'd471859200;
      42726: inst = 32'd136314880;
      42727: inst = 32'd268468224;
      42728: inst = 32'd201345344;
      42729: inst = 32'd203423744;
      42730: inst = 32'd471859200;
      42731: inst = 32'd136314880;
      42732: inst = 32'd268468224;
      42733: inst = 32'd201345345;
      42734: inst = 32'd203423744;
      42735: inst = 32'd471859200;
      42736: inst = 32'd136314880;
      42737: inst = 32'd268468224;
      42738: inst = 32'd201345346;
      42739: inst = 32'd203423744;
      42740: inst = 32'd471859200;
      42741: inst = 32'd136314880;
      42742: inst = 32'd268468224;
      42743: inst = 32'd201345347;
      42744: inst = 32'd203423744;
      42745: inst = 32'd471859200;
      42746: inst = 32'd136314880;
      42747: inst = 32'd268468224;
      42748: inst = 32'd201345348;
      42749: inst = 32'd203423744;
      42750: inst = 32'd471859200;
      42751: inst = 32'd136314880;
      42752: inst = 32'd268468224;
      42753: inst = 32'd201345349;
      42754: inst = 32'd203423744;
      42755: inst = 32'd471859200;
      42756: inst = 32'd136314880;
      42757: inst = 32'd268468224;
      42758: inst = 32'd201345350;
      42759: inst = 32'd203423744;
      42760: inst = 32'd471859200;
      42761: inst = 32'd136314880;
      42762: inst = 32'd268468224;
      42763: inst = 32'd201345351;
      42764: inst = 32'd203423744;
      42765: inst = 32'd471859200;
      42766: inst = 32'd136314880;
      42767: inst = 32'd268468224;
      42768: inst = 32'd201345352;
      42769: inst = 32'd203423744;
      42770: inst = 32'd471859200;
      42771: inst = 32'd136314880;
      42772: inst = 32'd268468224;
      42773: inst = 32'd201345353;
      42774: inst = 32'd203423744;
      42775: inst = 32'd471859200;
      42776: inst = 32'd136314880;
      42777: inst = 32'd268468224;
      42778: inst = 32'd201345354;
      42779: inst = 32'd203423744;
      42780: inst = 32'd471859200;
      42781: inst = 32'd136314880;
      42782: inst = 32'd268468224;
      42783: inst = 32'd201345355;
      42784: inst = 32'd203423744;
      42785: inst = 32'd471859200;
      42786: inst = 32'd136314880;
      42787: inst = 32'd268468224;
      42788: inst = 32'd201345356;
      42789: inst = 32'd203423744;
      42790: inst = 32'd471859200;
      42791: inst = 32'd136314880;
      42792: inst = 32'd268468224;
      42793: inst = 32'd201345357;
      42794: inst = 32'd203423744;
      42795: inst = 32'd471859200;
      42796: inst = 32'd136314880;
      42797: inst = 32'd268468224;
      42798: inst = 32'd201345358;
      42799: inst = 32'd203423744;
      42800: inst = 32'd471859200;
      42801: inst = 32'd136314880;
      42802: inst = 32'd268468224;
      42803: inst = 32'd201345359;
      42804: inst = 32'd203423744;
      42805: inst = 32'd471859200;
      42806: inst = 32'd136314880;
      42807: inst = 32'd268468224;
      42808: inst = 32'd201345360;
      42809: inst = 32'd203423744;
      42810: inst = 32'd471859200;
      42811: inst = 32'd136314880;
      42812: inst = 32'd268468224;
      42813: inst = 32'd201345361;
      42814: inst = 32'd203423744;
      42815: inst = 32'd471859200;
      42816: inst = 32'd136314880;
      42817: inst = 32'd268468224;
      42818: inst = 32'd201345362;
      42819: inst = 32'd203423744;
      42820: inst = 32'd471859200;
      42821: inst = 32'd136314880;
      42822: inst = 32'd268468224;
      42823: inst = 32'd201345363;
      42824: inst = 32'd203423744;
      42825: inst = 32'd471859200;
      42826: inst = 32'd136314880;
      42827: inst = 32'd268468224;
      42828: inst = 32'd201345364;
      42829: inst = 32'd203423744;
      42830: inst = 32'd471859200;
      42831: inst = 32'd136314880;
      42832: inst = 32'd268468224;
      42833: inst = 32'd201345365;
      42834: inst = 32'd203423744;
      42835: inst = 32'd471859200;
      42836: inst = 32'd136314880;
      42837: inst = 32'd268468224;
      42838: inst = 32'd201345366;
      42839: inst = 32'd203423744;
      42840: inst = 32'd471859200;
      42841: inst = 32'd136314880;
      42842: inst = 32'd268468224;
      42843: inst = 32'd201345367;
      42844: inst = 32'd203423744;
      42845: inst = 32'd471859200;
      42846: inst = 32'd136314880;
      42847: inst = 32'd268468224;
      42848: inst = 32'd201345368;
      42849: inst = 32'd203423744;
      42850: inst = 32'd471859200;
      42851: inst = 32'd136314880;
      42852: inst = 32'd268468224;
      42853: inst = 32'd201345369;
      42854: inst = 32'd203423744;
      42855: inst = 32'd471859200;
      42856: inst = 32'd136314880;
      42857: inst = 32'd268468224;
      42858: inst = 32'd201345370;
      42859: inst = 32'd203423744;
      42860: inst = 32'd471859200;
      42861: inst = 32'd136314880;
      42862: inst = 32'd268468224;
      42863: inst = 32'd201345371;
      42864: inst = 32'd203423744;
      42865: inst = 32'd471859200;
      42866: inst = 32'd136314880;
      42867: inst = 32'd268468224;
      42868: inst = 32'd201345372;
      42869: inst = 32'd203423744;
      42870: inst = 32'd471859200;
      42871: inst = 32'd136314880;
      42872: inst = 32'd268468224;
      42873: inst = 32'd201345373;
      42874: inst = 32'd203423744;
      42875: inst = 32'd471859200;
      42876: inst = 32'd136314880;
      42877: inst = 32'd268468224;
      42878: inst = 32'd201345374;
      42879: inst = 32'd203423744;
      42880: inst = 32'd471859200;
      42881: inst = 32'd136314880;
      42882: inst = 32'd268468224;
      42883: inst = 32'd201345375;
      42884: inst = 32'd203423744;
      42885: inst = 32'd471859200;
      42886: inst = 32'd136314880;
      42887: inst = 32'd268468224;
      42888: inst = 32'd201345376;
      42889: inst = 32'd203423744;
      42890: inst = 32'd471859200;
      42891: inst = 32'd136314880;
      42892: inst = 32'd268468224;
      42893: inst = 32'd201345377;
      42894: inst = 32'd203423744;
      42895: inst = 32'd471859200;
      42896: inst = 32'd136314880;
      42897: inst = 32'd268468224;
      42898: inst = 32'd201345378;
      42899: inst = 32'd203423744;
      42900: inst = 32'd471859200;
      42901: inst = 32'd136314880;
      42902: inst = 32'd268468224;
      42903: inst = 32'd201345379;
      42904: inst = 32'd203423744;
      42905: inst = 32'd471859200;
      42906: inst = 32'd136314880;
      42907: inst = 32'd268468224;
      42908: inst = 32'd201345380;
      42909: inst = 32'd203423744;
      42910: inst = 32'd471859200;
      42911: inst = 32'd136314880;
      42912: inst = 32'd268468224;
      42913: inst = 32'd201345381;
      42914: inst = 32'd203423744;
      42915: inst = 32'd471859200;
      42916: inst = 32'd136314880;
      42917: inst = 32'd268468224;
      42918: inst = 32'd201345382;
      42919: inst = 32'd203423744;
      42920: inst = 32'd471859200;
      42921: inst = 32'd136314880;
      42922: inst = 32'd268468224;
      42923: inst = 32'd201345383;
      42924: inst = 32'd203423744;
      42925: inst = 32'd471859200;
      42926: inst = 32'd136314880;
      42927: inst = 32'd268468224;
      42928: inst = 32'd201345384;
      42929: inst = 32'd203423744;
      42930: inst = 32'd471859200;
      42931: inst = 32'd136314880;
      42932: inst = 32'd268468224;
      42933: inst = 32'd201345385;
      42934: inst = 32'd203423744;
      42935: inst = 32'd471859200;
      42936: inst = 32'd136314880;
      42937: inst = 32'd268468224;
      42938: inst = 32'd201345386;
      42939: inst = 32'd203423744;
      42940: inst = 32'd471859200;
      42941: inst = 32'd136314880;
      42942: inst = 32'd268468224;
      42943: inst = 32'd201345387;
      42944: inst = 32'd203423744;
      42945: inst = 32'd471859200;
      42946: inst = 32'd136314880;
      42947: inst = 32'd268468224;
      42948: inst = 32'd201345388;
      42949: inst = 32'd203423744;
      42950: inst = 32'd471859200;
      42951: inst = 32'd136314880;
      42952: inst = 32'd268468224;
      42953: inst = 32'd201345389;
      42954: inst = 32'd203423744;
      42955: inst = 32'd471859200;
      42956: inst = 32'd136314880;
      42957: inst = 32'd268468224;
      42958: inst = 32'd201345390;
      42959: inst = 32'd203423744;
      42960: inst = 32'd471859200;
      42961: inst = 32'd136314880;
      42962: inst = 32'd268468224;
      42963: inst = 32'd201345391;
      42964: inst = 32'd203423744;
      42965: inst = 32'd471859200;
      42966: inst = 32'd136314880;
      42967: inst = 32'd268468224;
      42968: inst = 32'd201345392;
      42969: inst = 32'd203423744;
      42970: inst = 32'd471859200;
      42971: inst = 32'd136314880;
      42972: inst = 32'd268468224;
      42973: inst = 32'd201345393;
      42974: inst = 32'd203423744;
      42975: inst = 32'd471859200;
      42976: inst = 32'd136314880;
      42977: inst = 32'd268468224;
      42978: inst = 32'd201345394;
      42979: inst = 32'd203423744;
      42980: inst = 32'd471859200;
      42981: inst = 32'd136314880;
      42982: inst = 32'd268468224;
      42983: inst = 32'd201345395;
      42984: inst = 32'd203423744;
      42985: inst = 32'd471859200;
      42986: inst = 32'd136314880;
      42987: inst = 32'd268468224;
      42988: inst = 32'd201345396;
      42989: inst = 32'd203423744;
      42990: inst = 32'd471859200;
      42991: inst = 32'd136314880;
      42992: inst = 32'd268468224;
      42993: inst = 32'd201345397;
      42994: inst = 32'd203423744;
      42995: inst = 32'd471859200;
      42996: inst = 32'd136314880;
      42997: inst = 32'd268468224;
      42998: inst = 32'd201345398;
      42999: inst = 32'd203423744;
      43000: inst = 32'd471859200;
      43001: inst = 32'd136314880;
      43002: inst = 32'd268468224;
      43003: inst = 32'd201345399;
      43004: inst = 32'd203423744;
      43005: inst = 32'd471859200;
      43006: inst = 32'd136314880;
      43007: inst = 32'd268468224;
      43008: inst = 32'd201345400;
      43009: inst = 32'd203423744;
      43010: inst = 32'd471859200;
      43011: inst = 32'd136314880;
      43012: inst = 32'd268468224;
      43013: inst = 32'd201345401;
      43014: inst = 32'd203423744;
      43015: inst = 32'd471859200;
      43016: inst = 32'd136314880;
      43017: inst = 32'd268468224;
      43018: inst = 32'd201345402;
      43019: inst = 32'd203423744;
      43020: inst = 32'd471859200;
      43021: inst = 32'd136314880;
      43022: inst = 32'd268468224;
      43023: inst = 32'd201345403;
      43024: inst = 32'd203423744;
      43025: inst = 32'd471859200;
      43026: inst = 32'd136314880;
      43027: inst = 32'd268468224;
      43028: inst = 32'd201345404;
      43029: inst = 32'd203423744;
      43030: inst = 32'd471859200;
      43031: inst = 32'd136314880;
      43032: inst = 32'd268468224;
      43033: inst = 32'd201345405;
      43034: inst = 32'd203423744;
      43035: inst = 32'd471859200;
      43036: inst = 32'd136314880;
      43037: inst = 32'd268468224;
      43038: inst = 32'd201345406;
      43039: inst = 32'd203423744;
      43040: inst = 32'd471859200;
      43041: inst = 32'd136314880;
      43042: inst = 32'd268468224;
      43043: inst = 32'd201345407;
      43044: inst = 32'd203423744;
      43045: inst = 32'd471859200;
      43046: inst = 32'd136314880;
      43047: inst = 32'd268468224;
      43048: inst = 32'd201345408;
      43049: inst = 32'd203423744;
      43050: inst = 32'd471859200;
      43051: inst = 32'd136314880;
      43052: inst = 32'd268468224;
      43053: inst = 32'd201345409;
      43054: inst = 32'd203423744;
      43055: inst = 32'd471859200;
      43056: inst = 32'd136314880;
      43057: inst = 32'd268468224;
      43058: inst = 32'd201345410;
      43059: inst = 32'd203423744;
      43060: inst = 32'd471859200;
      43061: inst = 32'd136314880;
      43062: inst = 32'd268468224;
      43063: inst = 32'd201345411;
      43064: inst = 32'd203423744;
      43065: inst = 32'd471859200;
      43066: inst = 32'd136314880;
      43067: inst = 32'd268468224;
      43068: inst = 32'd201345412;
      43069: inst = 32'd203423744;
      43070: inst = 32'd471859200;
      43071: inst = 32'd136314880;
      43072: inst = 32'd268468224;
      43073: inst = 32'd201345413;
      43074: inst = 32'd203423744;
      43075: inst = 32'd471859200;
      43076: inst = 32'd136314880;
      43077: inst = 32'd268468224;
      43078: inst = 32'd201345414;
      43079: inst = 32'd203423744;
      43080: inst = 32'd471859200;
      43081: inst = 32'd136314880;
      43082: inst = 32'd268468224;
      43083: inst = 32'd201345415;
      43084: inst = 32'd203423744;
      43085: inst = 32'd471859200;
      43086: inst = 32'd136314880;
      43087: inst = 32'd268468224;
      43088: inst = 32'd201345416;
      43089: inst = 32'd203423744;
      43090: inst = 32'd471859200;
      43091: inst = 32'd136314880;
      43092: inst = 32'd268468224;
      43093: inst = 32'd201345417;
      43094: inst = 32'd203423744;
      43095: inst = 32'd471859200;
      43096: inst = 32'd136314880;
      43097: inst = 32'd268468224;
      43098: inst = 32'd201345418;
      43099: inst = 32'd203423744;
      43100: inst = 32'd471859200;
      43101: inst = 32'd136314880;
      43102: inst = 32'd268468224;
      43103: inst = 32'd201345419;
      43104: inst = 32'd203423744;
      43105: inst = 32'd471859200;
      43106: inst = 32'd136314880;
      43107: inst = 32'd268468224;
      43108: inst = 32'd201345420;
      43109: inst = 32'd203423744;
      43110: inst = 32'd471859200;
      43111: inst = 32'd136314880;
      43112: inst = 32'd268468224;
      43113: inst = 32'd201345421;
      43114: inst = 32'd203423744;
      43115: inst = 32'd471859200;
      43116: inst = 32'd136314880;
      43117: inst = 32'd268468224;
      43118: inst = 32'd201345422;
      43119: inst = 32'd203423744;
      43120: inst = 32'd471859200;
      43121: inst = 32'd136314880;
      43122: inst = 32'd268468224;
      43123: inst = 32'd201345423;
      43124: inst = 32'd203423744;
      43125: inst = 32'd471859200;
      43126: inst = 32'd136314880;
      43127: inst = 32'd268468224;
      43128: inst = 32'd201345424;
      43129: inst = 32'd203423744;
      43130: inst = 32'd471859200;
      43131: inst = 32'd136314880;
      43132: inst = 32'd268468224;
      43133: inst = 32'd201345425;
      43134: inst = 32'd203423744;
      43135: inst = 32'd471859200;
      43136: inst = 32'd136314880;
      43137: inst = 32'd268468224;
      43138: inst = 32'd201345426;
      43139: inst = 32'd203423744;
      43140: inst = 32'd471859200;
      43141: inst = 32'd136314880;
      43142: inst = 32'd268468224;
      43143: inst = 32'd201345427;
      43144: inst = 32'd203423744;
      43145: inst = 32'd471859200;
      43146: inst = 32'd136314880;
      43147: inst = 32'd268468224;
      43148: inst = 32'd201345428;
      43149: inst = 32'd203423744;
      43150: inst = 32'd471859200;
      43151: inst = 32'd136314880;
      43152: inst = 32'd268468224;
      43153: inst = 32'd201345429;
      43154: inst = 32'd203423744;
      43155: inst = 32'd471859200;
      43156: inst = 32'd136314880;
      43157: inst = 32'd268468224;
      43158: inst = 32'd201345430;
      43159: inst = 32'd203423744;
      43160: inst = 32'd471859200;
      43161: inst = 32'd136314880;
      43162: inst = 32'd268468224;
      43163: inst = 32'd201345431;
      43164: inst = 32'd203423744;
      43165: inst = 32'd471859200;
      43166: inst = 32'd136314880;
      43167: inst = 32'd268468224;
      43168: inst = 32'd201345432;
      43169: inst = 32'd203423744;
      43170: inst = 32'd471859200;
      43171: inst = 32'd136314880;
      43172: inst = 32'd268468224;
      43173: inst = 32'd201345433;
      43174: inst = 32'd203423744;
      43175: inst = 32'd471859200;
      43176: inst = 32'd136314880;
      43177: inst = 32'd268468224;
      43178: inst = 32'd201345434;
      43179: inst = 32'd203423744;
      43180: inst = 32'd471859200;
      43181: inst = 32'd136314880;
      43182: inst = 32'd268468224;
      43183: inst = 32'd201345435;
      43184: inst = 32'd203423744;
      43185: inst = 32'd471859200;
      43186: inst = 32'd136314880;
      43187: inst = 32'd268468224;
      43188: inst = 32'd201345436;
      43189: inst = 32'd203423744;
      43190: inst = 32'd471859200;
      43191: inst = 32'd136314880;
      43192: inst = 32'd268468224;
      43193: inst = 32'd201345437;
      43194: inst = 32'd203423744;
      43195: inst = 32'd471859200;
      43196: inst = 32'd136314880;
      43197: inst = 32'd268468224;
      43198: inst = 32'd201345438;
      43199: inst = 32'd203423744;
      43200: inst = 32'd471859200;
      43201: inst = 32'd136314880;
      43202: inst = 32'd268468224;
      43203: inst = 32'd201345439;
      43204: inst = 32'd203423744;
      43205: inst = 32'd471859200;
      43206: inst = 32'd136314880;
      43207: inst = 32'd268468224;
      43208: inst = 32'd201345440;
      43209: inst = 32'd203423744;
      43210: inst = 32'd471859200;
      43211: inst = 32'd136314880;
      43212: inst = 32'd268468224;
      43213: inst = 32'd201345441;
      43214: inst = 32'd203423744;
      43215: inst = 32'd471859200;
      43216: inst = 32'd136314880;
      43217: inst = 32'd268468224;
      43218: inst = 32'd201345442;
      43219: inst = 32'd203423744;
      43220: inst = 32'd471859200;
      43221: inst = 32'd136314880;
      43222: inst = 32'd268468224;
      43223: inst = 32'd201345443;
      43224: inst = 32'd203423744;
      43225: inst = 32'd471859200;
      43226: inst = 32'd136314880;
      43227: inst = 32'd268468224;
      43228: inst = 32'd201345444;
      43229: inst = 32'd203423744;
      43230: inst = 32'd471859200;
      43231: inst = 32'd136314880;
      43232: inst = 32'd268468224;
      43233: inst = 32'd201345445;
      43234: inst = 32'd203423744;
      43235: inst = 32'd471859200;
      43236: inst = 32'd136314880;
      43237: inst = 32'd268468224;
      43238: inst = 32'd201345446;
      43239: inst = 32'd203423744;
      43240: inst = 32'd471859200;
      43241: inst = 32'd136314880;
      43242: inst = 32'd268468224;
      43243: inst = 32'd201345447;
      43244: inst = 32'd203423744;
      43245: inst = 32'd471859200;
      43246: inst = 32'd136314880;
      43247: inst = 32'd268468224;
      43248: inst = 32'd201345448;
      43249: inst = 32'd203423744;
      43250: inst = 32'd471859200;
      43251: inst = 32'd136314880;
      43252: inst = 32'd268468224;
      43253: inst = 32'd201345449;
      43254: inst = 32'd203423744;
      43255: inst = 32'd471859200;
      43256: inst = 32'd136314880;
      43257: inst = 32'd268468224;
      43258: inst = 32'd201345450;
      43259: inst = 32'd203423744;
      43260: inst = 32'd471859200;
      43261: inst = 32'd136314880;
      43262: inst = 32'd268468224;
      43263: inst = 32'd201345451;
      43264: inst = 32'd203423744;
      43265: inst = 32'd471859200;
      43266: inst = 32'd136314880;
      43267: inst = 32'd268468224;
      43268: inst = 32'd201345452;
      43269: inst = 32'd203423744;
      43270: inst = 32'd471859200;
      43271: inst = 32'd136314880;
      43272: inst = 32'd268468224;
      43273: inst = 32'd201345453;
      43274: inst = 32'd203423744;
      43275: inst = 32'd471859200;
      43276: inst = 32'd136314880;
      43277: inst = 32'd268468224;
      43278: inst = 32'd201345454;
      43279: inst = 32'd203423744;
      43280: inst = 32'd471859200;
      43281: inst = 32'd136314880;
      43282: inst = 32'd268468224;
      43283: inst = 32'd201345455;
      43284: inst = 32'd203423744;
      43285: inst = 32'd471859200;
      43286: inst = 32'd136314880;
      43287: inst = 32'd268468224;
      43288: inst = 32'd201345456;
      43289: inst = 32'd203423744;
      43290: inst = 32'd471859200;
      43291: inst = 32'd136314880;
      43292: inst = 32'd268468224;
      43293: inst = 32'd201345457;
      43294: inst = 32'd203423744;
      43295: inst = 32'd471859200;
      43296: inst = 32'd136314880;
      43297: inst = 32'd268468224;
      43298: inst = 32'd201345458;
      43299: inst = 32'd203423744;
      43300: inst = 32'd471859200;
      43301: inst = 32'd136314880;
      43302: inst = 32'd268468224;
      43303: inst = 32'd201345459;
      43304: inst = 32'd203423744;
      43305: inst = 32'd471859200;
      43306: inst = 32'd136314880;
      43307: inst = 32'd268468224;
      43308: inst = 32'd201345460;
      43309: inst = 32'd203423744;
      43310: inst = 32'd471859200;
      43311: inst = 32'd136314880;
      43312: inst = 32'd268468224;
      43313: inst = 32'd201345461;
      43314: inst = 32'd203423744;
      43315: inst = 32'd471859200;
      43316: inst = 32'd136314880;
      43317: inst = 32'd268468224;
      43318: inst = 32'd201345462;
      43319: inst = 32'd203423744;
      43320: inst = 32'd471859200;
      43321: inst = 32'd136314880;
      43322: inst = 32'd268468224;
      43323: inst = 32'd201345463;
      43324: inst = 32'd203423744;
      43325: inst = 32'd471859200;
      43326: inst = 32'd136314880;
      43327: inst = 32'd268468224;
      43328: inst = 32'd201345464;
      43329: inst = 32'd203423744;
      43330: inst = 32'd471859200;
      43331: inst = 32'd136314880;
      43332: inst = 32'd268468224;
      43333: inst = 32'd201345465;
      43334: inst = 32'd203423744;
      43335: inst = 32'd471859200;
      43336: inst = 32'd136314880;
      43337: inst = 32'd268468224;
      43338: inst = 32'd201345466;
      43339: inst = 32'd203423744;
      43340: inst = 32'd471859200;
      43341: inst = 32'd136314880;
      43342: inst = 32'd268468224;
      43343: inst = 32'd201345467;
      43344: inst = 32'd203423744;
      43345: inst = 32'd471859200;
      43346: inst = 32'd136314880;
      43347: inst = 32'd268468224;
      43348: inst = 32'd201345468;
      43349: inst = 32'd203423744;
      43350: inst = 32'd471859200;
      43351: inst = 32'd136314880;
      43352: inst = 32'd268468224;
      43353: inst = 32'd201345469;
      43354: inst = 32'd203423744;
      43355: inst = 32'd471859200;
      43356: inst = 32'd136314880;
      43357: inst = 32'd268468224;
      43358: inst = 32'd201345470;
      43359: inst = 32'd203423744;
      43360: inst = 32'd471859200;
      43361: inst = 32'd136314880;
      43362: inst = 32'd268468224;
      43363: inst = 32'd201345471;
      43364: inst = 32'd203423744;
      43365: inst = 32'd471859200;
      43366: inst = 32'd136314880;
      43367: inst = 32'd268468224;
      43368: inst = 32'd201345472;
      43369: inst = 32'd203423744;
      43370: inst = 32'd471859200;
      43371: inst = 32'd136314880;
      43372: inst = 32'd268468224;
      43373: inst = 32'd201345473;
      43374: inst = 32'd203423744;
      43375: inst = 32'd471859200;
      43376: inst = 32'd136314880;
      43377: inst = 32'd268468224;
      43378: inst = 32'd201345474;
      43379: inst = 32'd203423744;
      43380: inst = 32'd471859200;
      43381: inst = 32'd136314880;
      43382: inst = 32'd268468224;
      43383: inst = 32'd201345475;
      43384: inst = 32'd203423744;
      43385: inst = 32'd471859200;
      43386: inst = 32'd136314880;
      43387: inst = 32'd268468224;
      43388: inst = 32'd201345476;
      43389: inst = 32'd203423744;
      43390: inst = 32'd471859200;
      43391: inst = 32'd136314880;
      43392: inst = 32'd268468224;
      43393: inst = 32'd201345477;
      43394: inst = 32'd203423744;
      43395: inst = 32'd471859200;
      43396: inst = 32'd136314880;
      43397: inst = 32'd268468224;
      43398: inst = 32'd201345478;
      43399: inst = 32'd203423744;
      43400: inst = 32'd471859200;
      43401: inst = 32'd136314880;
      43402: inst = 32'd268468224;
      43403: inst = 32'd201345479;
      43404: inst = 32'd203423744;
      43405: inst = 32'd471859200;
      43406: inst = 32'd136314880;
      43407: inst = 32'd268468224;
      43408: inst = 32'd201345480;
      43409: inst = 32'd203423744;
      43410: inst = 32'd471859200;
      43411: inst = 32'd136314880;
      43412: inst = 32'd268468224;
      43413: inst = 32'd201345481;
      43414: inst = 32'd203423744;
      43415: inst = 32'd471859200;
      43416: inst = 32'd136314880;
      43417: inst = 32'd268468224;
      43418: inst = 32'd201345482;
      43419: inst = 32'd203423744;
      43420: inst = 32'd471859200;
      43421: inst = 32'd136314880;
      43422: inst = 32'd268468224;
      43423: inst = 32'd201345483;
      43424: inst = 32'd203423744;
      43425: inst = 32'd471859200;
      43426: inst = 32'd136314880;
      43427: inst = 32'd268468224;
      43428: inst = 32'd201345484;
      43429: inst = 32'd203423744;
      43430: inst = 32'd471859200;
      43431: inst = 32'd136314880;
      43432: inst = 32'd268468224;
      43433: inst = 32'd201345485;
      43434: inst = 32'd203423744;
      43435: inst = 32'd471859200;
      43436: inst = 32'd136314880;
      43437: inst = 32'd268468224;
      43438: inst = 32'd201345486;
      43439: inst = 32'd203423744;
      43440: inst = 32'd471859200;
      43441: inst = 32'd136314880;
      43442: inst = 32'd268468224;
      43443: inst = 32'd201345487;
      43444: inst = 32'd203423744;
      43445: inst = 32'd471859200;
      43446: inst = 32'd136314880;
      43447: inst = 32'd268468224;
      43448: inst = 32'd201345488;
      43449: inst = 32'd203423744;
      43450: inst = 32'd471859200;
      43451: inst = 32'd136314880;
      43452: inst = 32'd268468224;
      43453: inst = 32'd201345489;
      43454: inst = 32'd203423744;
      43455: inst = 32'd471859200;
      43456: inst = 32'd136314880;
      43457: inst = 32'd268468224;
      43458: inst = 32'd201345490;
      43459: inst = 32'd203423744;
      43460: inst = 32'd471859200;
      43461: inst = 32'd136314880;
      43462: inst = 32'd268468224;
      43463: inst = 32'd201345491;
      43464: inst = 32'd203423744;
      43465: inst = 32'd471859200;
      43466: inst = 32'd136314880;
      43467: inst = 32'd268468224;
      43468: inst = 32'd201345492;
      43469: inst = 32'd203423744;
      43470: inst = 32'd471859200;
      43471: inst = 32'd136314880;
      43472: inst = 32'd268468224;
      43473: inst = 32'd201345493;
      43474: inst = 32'd203423744;
      43475: inst = 32'd471859200;
      43476: inst = 32'd136314880;
      43477: inst = 32'd268468224;
      43478: inst = 32'd201345494;
      43479: inst = 32'd203423744;
      43480: inst = 32'd471859200;
      43481: inst = 32'd136314880;
      43482: inst = 32'd268468224;
      43483: inst = 32'd201345495;
      43484: inst = 32'd203423744;
      43485: inst = 32'd471859200;
      43486: inst = 32'd136314880;
      43487: inst = 32'd268468224;
      43488: inst = 32'd201345496;
      43489: inst = 32'd203423744;
      43490: inst = 32'd471859200;
      43491: inst = 32'd136314880;
      43492: inst = 32'd268468224;
      43493: inst = 32'd201345497;
      43494: inst = 32'd203423744;
      43495: inst = 32'd471859200;
      43496: inst = 32'd136314880;
      43497: inst = 32'd268468224;
      43498: inst = 32'd201345498;
      43499: inst = 32'd203423744;
      43500: inst = 32'd471859200;
      43501: inst = 32'd136314880;
      43502: inst = 32'd268468224;
      43503: inst = 32'd201345499;
      43504: inst = 32'd203423744;
      43505: inst = 32'd471859200;
      43506: inst = 32'd136314880;
      43507: inst = 32'd268468224;
      43508: inst = 32'd201345500;
      43509: inst = 32'd203423744;
      43510: inst = 32'd471859200;
      43511: inst = 32'd136314880;
      43512: inst = 32'd268468224;
      43513: inst = 32'd201345501;
      43514: inst = 32'd203423744;
      43515: inst = 32'd471859200;
      43516: inst = 32'd136314880;
      43517: inst = 32'd268468224;
      43518: inst = 32'd201345502;
      43519: inst = 32'd203423744;
      43520: inst = 32'd471859200;
      43521: inst = 32'd136314880;
      43522: inst = 32'd268468224;
      43523: inst = 32'd201345503;
      43524: inst = 32'd203423744;
      43525: inst = 32'd471859200;
      43526: inst = 32'd136314880;
      43527: inst = 32'd268468224;
      43528: inst = 32'd201345504;
      43529: inst = 32'd203423744;
      43530: inst = 32'd471859200;
      43531: inst = 32'd136314880;
      43532: inst = 32'd268468224;
      43533: inst = 32'd201345505;
      43534: inst = 32'd203423744;
      43535: inst = 32'd471859200;
      43536: inst = 32'd136314880;
      43537: inst = 32'd268468224;
      43538: inst = 32'd201345506;
      43539: inst = 32'd203423744;
      43540: inst = 32'd471859200;
      43541: inst = 32'd136314880;
      43542: inst = 32'd268468224;
      43543: inst = 32'd201345507;
      43544: inst = 32'd203423744;
      43545: inst = 32'd471859200;
      43546: inst = 32'd136314880;
      43547: inst = 32'd268468224;
      43548: inst = 32'd201345508;
      43549: inst = 32'd203423744;
      43550: inst = 32'd471859200;
      43551: inst = 32'd136314880;
      43552: inst = 32'd268468224;
      43553: inst = 32'd201345509;
      43554: inst = 32'd203423744;
      43555: inst = 32'd471859200;
      43556: inst = 32'd136314880;
      43557: inst = 32'd268468224;
      43558: inst = 32'd201345510;
      43559: inst = 32'd203423744;
      43560: inst = 32'd471859200;
      43561: inst = 32'd136314880;
      43562: inst = 32'd268468224;
      43563: inst = 32'd201345511;
      43564: inst = 32'd203423744;
      43565: inst = 32'd471859200;
      43566: inst = 32'd136314880;
      43567: inst = 32'd268468224;
      43568: inst = 32'd201345512;
      43569: inst = 32'd203423744;
      43570: inst = 32'd471859200;
      43571: inst = 32'd136314880;
      43572: inst = 32'd268468224;
      43573: inst = 32'd201345513;
      43574: inst = 32'd203423744;
      43575: inst = 32'd471859200;
      43576: inst = 32'd136314880;
      43577: inst = 32'd268468224;
      43578: inst = 32'd201345514;
      43579: inst = 32'd203423744;
      43580: inst = 32'd471859200;
      43581: inst = 32'd136314880;
      43582: inst = 32'd268468224;
      43583: inst = 32'd201345515;
      43584: inst = 32'd203423744;
      43585: inst = 32'd471859200;
      43586: inst = 32'd136314880;
      43587: inst = 32'd268468224;
      43588: inst = 32'd201345516;
      43589: inst = 32'd203423744;
      43590: inst = 32'd471859200;
      43591: inst = 32'd136314880;
      43592: inst = 32'd268468224;
      43593: inst = 32'd201345517;
      43594: inst = 32'd203423744;
      43595: inst = 32'd471859200;
      43596: inst = 32'd136314880;
      43597: inst = 32'd268468224;
      43598: inst = 32'd201345518;
      43599: inst = 32'd203423744;
      43600: inst = 32'd471859200;
      43601: inst = 32'd136314880;
      43602: inst = 32'd268468224;
      43603: inst = 32'd201345519;
      43604: inst = 32'd203423744;
      43605: inst = 32'd471859200;
      43606: inst = 32'd136314880;
      43607: inst = 32'd268468224;
      43608: inst = 32'd201345520;
      43609: inst = 32'd203423744;
      43610: inst = 32'd471859200;
      43611: inst = 32'd136314880;
      43612: inst = 32'd268468224;
      43613: inst = 32'd201345521;
      43614: inst = 32'd203423744;
      43615: inst = 32'd471859200;
      43616: inst = 32'd136314880;
      43617: inst = 32'd268468224;
      43618: inst = 32'd201345522;
      43619: inst = 32'd203423744;
      43620: inst = 32'd471859200;
      43621: inst = 32'd136314880;
      43622: inst = 32'd268468224;
      43623: inst = 32'd201345523;
      43624: inst = 32'd203423744;
      43625: inst = 32'd471859200;
      43626: inst = 32'd136314880;
      43627: inst = 32'd268468224;
      43628: inst = 32'd201345524;
      43629: inst = 32'd203423744;
      43630: inst = 32'd471859200;
      43631: inst = 32'd136314880;
      43632: inst = 32'd268468224;
      43633: inst = 32'd201345525;
      43634: inst = 32'd203423744;
      43635: inst = 32'd471859200;
      43636: inst = 32'd136314880;
      43637: inst = 32'd268468224;
      43638: inst = 32'd201345526;
      43639: inst = 32'd203423744;
      43640: inst = 32'd471859200;
      43641: inst = 32'd136314880;
      43642: inst = 32'd268468224;
      43643: inst = 32'd201345527;
      43644: inst = 32'd203423744;
      43645: inst = 32'd471859200;
      43646: inst = 32'd136314880;
      43647: inst = 32'd268468224;
      43648: inst = 32'd201345528;
      43649: inst = 32'd203423744;
      43650: inst = 32'd471859200;
      43651: inst = 32'd136314880;
      43652: inst = 32'd268468224;
      43653: inst = 32'd201345529;
      43654: inst = 32'd203423744;
      43655: inst = 32'd471859200;
      43656: inst = 32'd136314880;
      43657: inst = 32'd268468224;
      43658: inst = 32'd201345530;
      43659: inst = 32'd203423744;
      43660: inst = 32'd471859200;
      43661: inst = 32'd136314880;
      43662: inst = 32'd268468224;
      43663: inst = 32'd201345531;
      43664: inst = 32'd203423744;
      43665: inst = 32'd471859200;
      43666: inst = 32'd136314880;
      43667: inst = 32'd268468224;
      43668: inst = 32'd201345532;
      43669: inst = 32'd203423744;
      43670: inst = 32'd471859200;
      43671: inst = 32'd136314880;
      43672: inst = 32'd268468224;
      43673: inst = 32'd201345533;
      43674: inst = 32'd203423744;
      43675: inst = 32'd471859200;
      43676: inst = 32'd136314880;
      43677: inst = 32'd268468224;
      43678: inst = 32'd201345534;
      43679: inst = 32'd203423744;
      43680: inst = 32'd471859200;
      43681: inst = 32'd136314880;
      43682: inst = 32'd268468224;
      43683: inst = 32'd201345535;
      43684: inst = 32'd203423744;
      43685: inst = 32'd471859200;
      43686: inst = 32'd136314880;
      43687: inst = 32'd268468224;
      43688: inst = 32'd201345536;
      43689: inst = 32'd203423744;
      43690: inst = 32'd471859200;
      43691: inst = 32'd136314880;
      43692: inst = 32'd268468224;
      43693: inst = 32'd201345537;
      43694: inst = 32'd203423744;
      43695: inst = 32'd471859200;
      43696: inst = 32'd136314880;
      43697: inst = 32'd268468224;
      43698: inst = 32'd201345538;
      43699: inst = 32'd203423744;
      43700: inst = 32'd471859200;
      43701: inst = 32'd136314880;
      43702: inst = 32'd268468224;
      43703: inst = 32'd201345539;
      43704: inst = 32'd203423744;
      43705: inst = 32'd471859200;
      43706: inst = 32'd136314880;
      43707: inst = 32'd268468224;
      43708: inst = 32'd201345540;
      43709: inst = 32'd203423744;
      43710: inst = 32'd471859200;
      43711: inst = 32'd136314880;
      43712: inst = 32'd268468224;
      43713: inst = 32'd201345541;
      43714: inst = 32'd203423744;
      43715: inst = 32'd471859200;
      43716: inst = 32'd136314880;
      43717: inst = 32'd268468224;
      43718: inst = 32'd201345542;
      43719: inst = 32'd203423744;
      43720: inst = 32'd471859200;
      43721: inst = 32'd136314880;
      43722: inst = 32'd268468224;
      43723: inst = 32'd201345543;
      43724: inst = 32'd203423744;
      43725: inst = 32'd471859200;
      43726: inst = 32'd136314880;
      43727: inst = 32'd268468224;
      43728: inst = 32'd201345544;
      43729: inst = 32'd203423744;
      43730: inst = 32'd471859200;
      43731: inst = 32'd136314880;
      43732: inst = 32'd268468224;
      43733: inst = 32'd201345545;
      43734: inst = 32'd203423744;
      43735: inst = 32'd471859200;
      43736: inst = 32'd136314880;
      43737: inst = 32'd268468224;
      43738: inst = 32'd201345546;
      43739: inst = 32'd203423744;
      43740: inst = 32'd471859200;
      43741: inst = 32'd136314880;
      43742: inst = 32'd268468224;
      43743: inst = 32'd201345547;
      43744: inst = 32'd203423744;
      43745: inst = 32'd471859200;
      43746: inst = 32'd136314880;
      43747: inst = 32'd268468224;
      43748: inst = 32'd201345548;
      43749: inst = 32'd203423744;
      43750: inst = 32'd471859200;
      43751: inst = 32'd136314880;
      43752: inst = 32'd268468224;
      43753: inst = 32'd201345549;
      43754: inst = 32'd203423744;
      43755: inst = 32'd471859200;
      43756: inst = 32'd136314880;
      43757: inst = 32'd268468224;
      43758: inst = 32'd201345550;
      43759: inst = 32'd203423744;
      43760: inst = 32'd471859200;
      43761: inst = 32'd136314880;
      43762: inst = 32'd268468224;
      43763: inst = 32'd201345551;
      43764: inst = 32'd203423744;
      43765: inst = 32'd471859200;
      43766: inst = 32'd136314880;
      43767: inst = 32'd268468224;
      43768: inst = 32'd201345552;
      43769: inst = 32'd203423744;
      43770: inst = 32'd471859200;
      43771: inst = 32'd136314880;
      43772: inst = 32'd268468224;
      43773: inst = 32'd201345553;
      43774: inst = 32'd203423744;
      43775: inst = 32'd471859200;
      43776: inst = 32'd136314880;
      43777: inst = 32'd268468224;
      43778: inst = 32'd201345554;
      43779: inst = 32'd203423744;
      43780: inst = 32'd471859200;
      43781: inst = 32'd136314880;
      43782: inst = 32'd268468224;
      43783: inst = 32'd201345555;
      43784: inst = 32'd203423744;
      43785: inst = 32'd471859200;
      43786: inst = 32'd136314880;
      43787: inst = 32'd268468224;
      43788: inst = 32'd201345556;
      43789: inst = 32'd203423744;
      43790: inst = 32'd471859200;
      43791: inst = 32'd136314880;
      43792: inst = 32'd268468224;
      43793: inst = 32'd201345557;
      43794: inst = 32'd203423744;
      43795: inst = 32'd471859200;
      43796: inst = 32'd136314880;
      43797: inst = 32'd268468224;
      43798: inst = 32'd201345558;
      43799: inst = 32'd203423744;
      43800: inst = 32'd471859200;
      43801: inst = 32'd136314880;
      43802: inst = 32'd268468224;
      43803: inst = 32'd201345559;
      43804: inst = 32'd203423744;
      43805: inst = 32'd471859200;
      43806: inst = 32'd136314880;
      43807: inst = 32'd268468224;
      43808: inst = 32'd201345560;
      43809: inst = 32'd203423744;
      43810: inst = 32'd471859200;
      43811: inst = 32'd136314880;
      43812: inst = 32'd268468224;
      43813: inst = 32'd201345561;
      43814: inst = 32'd203423744;
      43815: inst = 32'd471859200;
      43816: inst = 32'd136314880;
      43817: inst = 32'd268468224;
      43818: inst = 32'd201345562;
      43819: inst = 32'd203423744;
      43820: inst = 32'd471859200;
      43821: inst = 32'd136314880;
      43822: inst = 32'd268468224;
      43823: inst = 32'd201345563;
      43824: inst = 32'd203423744;
      43825: inst = 32'd471859200;
      43826: inst = 32'd136314880;
      43827: inst = 32'd268468224;
      43828: inst = 32'd201345564;
      43829: inst = 32'd203423744;
      43830: inst = 32'd471859200;
      43831: inst = 32'd136314880;
      43832: inst = 32'd268468224;
      43833: inst = 32'd201345565;
      43834: inst = 32'd203423744;
      43835: inst = 32'd471859200;
      43836: inst = 32'd136314880;
      43837: inst = 32'd268468224;
      43838: inst = 32'd201345566;
      43839: inst = 32'd203423744;
      43840: inst = 32'd471859200;
      43841: inst = 32'd136314880;
      43842: inst = 32'd268468224;
      43843: inst = 32'd201345567;
      43844: inst = 32'd203423744;
      43845: inst = 32'd471859200;
      43846: inst = 32'd136314880;
      43847: inst = 32'd268468224;
      43848: inst = 32'd201345568;
      43849: inst = 32'd203423744;
      43850: inst = 32'd471859200;
      43851: inst = 32'd136314880;
      43852: inst = 32'd268468224;
      43853: inst = 32'd201345569;
      43854: inst = 32'd203423744;
      43855: inst = 32'd471859200;
      43856: inst = 32'd136314880;
      43857: inst = 32'd268468224;
      43858: inst = 32'd201345570;
      43859: inst = 32'd203423744;
      43860: inst = 32'd471859200;
      43861: inst = 32'd136314880;
      43862: inst = 32'd268468224;
      43863: inst = 32'd201345571;
      43864: inst = 32'd203423744;
      43865: inst = 32'd471859200;
      43866: inst = 32'd136314880;
      43867: inst = 32'd268468224;
      43868: inst = 32'd201345572;
      43869: inst = 32'd203423744;
      43870: inst = 32'd471859200;
      43871: inst = 32'd136314880;
      43872: inst = 32'd268468224;
      43873: inst = 32'd201345573;
      43874: inst = 32'd203423744;
      43875: inst = 32'd471859200;
      43876: inst = 32'd136314880;
      43877: inst = 32'd268468224;
      43878: inst = 32'd201345574;
      43879: inst = 32'd203423744;
      43880: inst = 32'd471859200;
      43881: inst = 32'd136314880;
      43882: inst = 32'd268468224;
      43883: inst = 32'd201345575;
      43884: inst = 32'd203423744;
      43885: inst = 32'd471859200;
      43886: inst = 32'd136314880;
      43887: inst = 32'd268468224;
      43888: inst = 32'd201345576;
      43889: inst = 32'd203423744;
      43890: inst = 32'd471859200;
      43891: inst = 32'd136314880;
      43892: inst = 32'd268468224;
      43893: inst = 32'd201345577;
      43894: inst = 32'd203423744;
      43895: inst = 32'd471859200;
      43896: inst = 32'd136314880;
      43897: inst = 32'd268468224;
      43898: inst = 32'd201345578;
      43899: inst = 32'd203423744;
      43900: inst = 32'd471859200;
      43901: inst = 32'd136314880;
      43902: inst = 32'd268468224;
      43903: inst = 32'd201345579;
      43904: inst = 32'd203423744;
      43905: inst = 32'd471859200;
      43906: inst = 32'd136314880;
      43907: inst = 32'd268468224;
      43908: inst = 32'd201345580;
      43909: inst = 32'd203423744;
      43910: inst = 32'd471859200;
      43911: inst = 32'd136314880;
      43912: inst = 32'd268468224;
      43913: inst = 32'd201345581;
      43914: inst = 32'd203423744;
      43915: inst = 32'd471859200;
      43916: inst = 32'd136314880;
      43917: inst = 32'd268468224;
      43918: inst = 32'd201345582;
      43919: inst = 32'd203423744;
      43920: inst = 32'd471859200;
      43921: inst = 32'd136314880;
      43922: inst = 32'd268468224;
      43923: inst = 32'd201345583;
      43924: inst = 32'd203423744;
      43925: inst = 32'd471859200;
      43926: inst = 32'd136314880;
      43927: inst = 32'd268468224;
      43928: inst = 32'd201345584;
      43929: inst = 32'd203423744;
      43930: inst = 32'd471859200;
      43931: inst = 32'd136314880;
      43932: inst = 32'd268468224;
      43933: inst = 32'd201345585;
      43934: inst = 32'd203423744;
      43935: inst = 32'd471859200;
      43936: inst = 32'd136314880;
      43937: inst = 32'd268468224;
      43938: inst = 32'd201345586;
      43939: inst = 32'd203423744;
      43940: inst = 32'd471859200;
      43941: inst = 32'd136314880;
      43942: inst = 32'd268468224;
      43943: inst = 32'd201345587;
      43944: inst = 32'd203423744;
      43945: inst = 32'd471859200;
      43946: inst = 32'd136314880;
      43947: inst = 32'd268468224;
      43948: inst = 32'd201345588;
      43949: inst = 32'd203423744;
      43950: inst = 32'd471859200;
      43951: inst = 32'd136314880;
      43952: inst = 32'd268468224;
      43953: inst = 32'd201345589;
      43954: inst = 32'd203423744;
      43955: inst = 32'd471859200;
      43956: inst = 32'd136314880;
      43957: inst = 32'd268468224;
      43958: inst = 32'd201345590;
      43959: inst = 32'd203423744;
      43960: inst = 32'd471859200;
      43961: inst = 32'd136314880;
      43962: inst = 32'd268468224;
      43963: inst = 32'd201345591;
      43964: inst = 32'd203423744;
      43965: inst = 32'd471859200;
      43966: inst = 32'd136314880;
      43967: inst = 32'd268468224;
      43968: inst = 32'd201345592;
      43969: inst = 32'd203423744;
      43970: inst = 32'd471859200;
      43971: inst = 32'd136314880;
      43972: inst = 32'd268468224;
      43973: inst = 32'd201345593;
      43974: inst = 32'd203423744;
      43975: inst = 32'd471859200;
      43976: inst = 32'd136314880;
      43977: inst = 32'd268468224;
      43978: inst = 32'd201345594;
      43979: inst = 32'd203423744;
      43980: inst = 32'd471859200;
      43981: inst = 32'd136314880;
      43982: inst = 32'd268468224;
      43983: inst = 32'd201345595;
      43984: inst = 32'd203423744;
      43985: inst = 32'd471859200;
      43986: inst = 32'd136314880;
      43987: inst = 32'd268468224;
      43988: inst = 32'd201345596;
      43989: inst = 32'd203423744;
      43990: inst = 32'd471859200;
      43991: inst = 32'd136314880;
      43992: inst = 32'd268468224;
      43993: inst = 32'd201345597;
      43994: inst = 32'd203423744;
      43995: inst = 32'd471859200;
      43996: inst = 32'd136314880;
      43997: inst = 32'd268468224;
      43998: inst = 32'd201345598;
      43999: inst = 32'd203423744;
      44000: inst = 32'd471859200;
      44001: inst = 32'd136314880;
      44002: inst = 32'd268468224;
      44003: inst = 32'd201345599;
      44004: inst = 32'd203423744;
      44005: inst = 32'd471859200;
      44006: inst = 32'd136314880;
      44007: inst = 32'd268468224;
      44008: inst = 32'd201345600;
      44009: inst = 32'd203423744;
      44010: inst = 32'd471859200;
      44011: inst = 32'd136314880;
      44012: inst = 32'd268468224;
      44013: inst = 32'd201345601;
      44014: inst = 32'd203423744;
      44015: inst = 32'd471859200;
      44016: inst = 32'd136314880;
      44017: inst = 32'd268468224;
      44018: inst = 32'd201345602;
      44019: inst = 32'd203423744;
      44020: inst = 32'd471859200;
      44021: inst = 32'd136314880;
      44022: inst = 32'd268468224;
      44023: inst = 32'd201345603;
      44024: inst = 32'd203423744;
      44025: inst = 32'd471859200;
      44026: inst = 32'd136314880;
      44027: inst = 32'd268468224;
      44028: inst = 32'd201345604;
      44029: inst = 32'd203423744;
      44030: inst = 32'd471859200;
      44031: inst = 32'd136314880;
      44032: inst = 32'd268468224;
      44033: inst = 32'd201345605;
      44034: inst = 32'd203423744;
      44035: inst = 32'd471859200;
      44036: inst = 32'd136314880;
      44037: inst = 32'd268468224;
      44038: inst = 32'd201345606;
      44039: inst = 32'd203423744;
      44040: inst = 32'd471859200;
      44041: inst = 32'd136314880;
      44042: inst = 32'd268468224;
      44043: inst = 32'd201345607;
      44044: inst = 32'd203423744;
      44045: inst = 32'd471859200;
      44046: inst = 32'd136314880;
      44047: inst = 32'd268468224;
      44048: inst = 32'd201345608;
      44049: inst = 32'd203423744;
      44050: inst = 32'd471859200;
      44051: inst = 32'd136314880;
      44052: inst = 32'd268468224;
      44053: inst = 32'd201345609;
      44054: inst = 32'd203423744;
      44055: inst = 32'd471859200;
      44056: inst = 32'd136314880;
      44057: inst = 32'd268468224;
      44058: inst = 32'd201345610;
      44059: inst = 32'd203423744;
      44060: inst = 32'd471859200;
      44061: inst = 32'd136314880;
      44062: inst = 32'd268468224;
      44063: inst = 32'd201345611;
      44064: inst = 32'd203423744;
      44065: inst = 32'd471859200;
      44066: inst = 32'd136314880;
      44067: inst = 32'd268468224;
      44068: inst = 32'd201345612;
      44069: inst = 32'd203423744;
      44070: inst = 32'd471859200;
      44071: inst = 32'd136314880;
      44072: inst = 32'd268468224;
      44073: inst = 32'd201345613;
      44074: inst = 32'd203423744;
      44075: inst = 32'd471859200;
      44076: inst = 32'd136314880;
      44077: inst = 32'd268468224;
      44078: inst = 32'd201345614;
      44079: inst = 32'd203423744;
      44080: inst = 32'd471859200;
      44081: inst = 32'd136314880;
      44082: inst = 32'd268468224;
      44083: inst = 32'd201345615;
      44084: inst = 32'd203423744;
      44085: inst = 32'd471859200;
      44086: inst = 32'd136314880;
      44087: inst = 32'd268468224;
      44088: inst = 32'd201345616;
      44089: inst = 32'd203423744;
      44090: inst = 32'd471859200;
      44091: inst = 32'd136314880;
      44092: inst = 32'd268468224;
      44093: inst = 32'd201345617;
      44094: inst = 32'd203423744;
      44095: inst = 32'd471859200;
      44096: inst = 32'd136314880;
      44097: inst = 32'd268468224;
      44098: inst = 32'd201345618;
      44099: inst = 32'd203423744;
      44100: inst = 32'd471859200;
      44101: inst = 32'd136314880;
      44102: inst = 32'd268468224;
      44103: inst = 32'd201345619;
      44104: inst = 32'd203423744;
      44105: inst = 32'd471859200;
      44106: inst = 32'd136314880;
      44107: inst = 32'd268468224;
      44108: inst = 32'd201345620;
      44109: inst = 32'd203423744;
      44110: inst = 32'd471859200;
      44111: inst = 32'd136314880;
      44112: inst = 32'd268468224;
      44113: inst = 32'd201345621;
      44114: inst = 32'd203423744;
      44115: inst = 32'd471859200;
      44116: inst = 32'd136314880;
      44117: inst = 32'd268468224;
      44118: inst = 32'd201345622;
      44119: inst = 32'd203423744;
      44120: inst = 32'd471859200;
      44121: inst = 32'd136314880;
      44122: inst = 32'd268468224;
      44123: inst = 32'd201345623;
      44124: inst = 32'd203423744;
      44125: inst = 32'd471859200;
      44126: inst = 32'd136314880;
      44127: inst = 32'd268468224;
      44128: inst = 32'd201345624;
      44129: inst = 32'd203423744;
      44130: inst = 32'd471859200;
      44131: inst = 32'd136314880;
      44132: inst = 32'd268468224;
      44133: inst = 32'd201345625;
      44134: inst = 32'd203423744;
      44135: inst = 32'd471859200;
      44136: inst = 32'd136314880;
      44137: inst = 32'd268468224;
      44138: inst = 32'd201345626;
      44139: inst = 32'd203423744;
      44140: inst = 32'd471859200;
      44141: inst = 32'd136314880;
      44142: inst = 32'd268468224;
      44143: inst = 32'd201345627;
      44144: inst = 32'd203423744;
      44145: inst = 32'd471859200;
      44146: inst = 32'd136314880;
      44147: inst = 32'd268468224;
      44148: inst = 32'd201345628;
      44149: inst = 32'd203423744;
      44150: inst = 32'd471859200;
      44151: inst = 32'd136314880;
      44152: inst = 32'd268468224;
      44153: inst = 32'd201345629;
      44154: inst = 32'd203423744;
      44155: inst = 32'd471859200;
      44156: inst = 32'd136314880;
      44157: inst = 32'd268468224;
      44158: inst = 32'd201345630;
      44159: inst = 32'd203423744;
      44160: inst = 32'd471859200;
      44161: inst = 32'd136314880;
      44162: inst = 32'd268468224;
      44163: inst = 32'd201345631;
      44164: inst = 32'd203423744;
      44165: inst = 32'd471859200;
      44166: inst = 32'd136314880;
      44167: inst = 32'd268468224;
      44168: inst = 32'd201345632;
      44169: inst = 32'd203423744;
      44170: inst = 32'd471859200;
      44171: inst = 32'd136314880;
      44172: inst = 32'd268468224;
      44173: inst = 32'd201345633;
      44174: inst = 32'd203423744;
      44175: inst = 32'd471859200;
      44176: inst = 32'd136314880;
      44177: inst = 32'd268468224;
      44178: inst = 32'd201345634;
      44179: inst = 32'd203423744;
      44180: inst = 32'd471859200;
      44181: inst = 32'd136314880;
      44182: inst = 32'd268468224;
      44183: inst = 32'd201345635;
      44184: inst = 32'd203423744;
      44185: inst = 32'd471859200;
      44186: inst = 32'd136314880;
      44187: inst = 32'd268468224;
      44188: inst = 32'd201345636;
      44189: inst = 32'd203423744;
      44190: inst = 32'd471859200;
      44191: inst = 32'd136314880;
      44192: inst = 32'd268468224;
      44193: inst = 32'd201345637;
      44194: inst = 32'd203423744;
      44195: inst = 32'd471859200;
      44196: inst = 32'd136314880;
      44197: inst = 32'd268468224;
      44198: inst = 32'd201345638;
      44199: inst = 32'd203423744;
      44200: inst = 32'd471859200;
      44201: inst = 32'd136314880;
      44202: inst = 32'd268468224;
      44203: inst = 32'd201345639;
      44204: inst = 32'd203423744;
      44205: inst = 32'd471859200;
      44206: inst = 32'd136314880;
      44207: inst = 32'd268468224;
      44208: inst = 32'd201345640;
      44209: inst = 32'd203423744;
      44210: inst = 32'd471859200;
      44211: inst = 32'd136314880;
      44212: inst = 32'd268468224;
      44213: inst = 32'd201345641;
      44214: inst = 32'd203423744;
      44215: inst = 32'd471859200;
      44216: inst = 32'd136314880;
      44217: inst = 32'd268468224;
      44218: inst = 32'd201345642;
      44219: inst = 32'd203423744;
      44220: inst = 32'd471859200;
      44221: inst = 32'd136314880;
      44222: inst = 32'd268468224;
      44223: inst = 32'd201345643;
      44224: inst = 32'd203423744;
      44225: inst = 32'd471859200;
      44226: inst = 32'd136314880;
      44227: inst = 32'd268468224;
      44228: inst = 32'd201345644;
      44229: inst = 32'd203423744;
      44230: inst = 32'd471859200;
      44231: inst = 32'd136314880;
      44232: inst = 32'd268468224;
      44233: inst = 32'd201345645;
      44234: inst = 32'd203423744;
      44235: inst = 32'd471859200;
      44236: inst = 32'd136314880;
      44237: inst = 32'd268468224;
      44238: inst = 32'd201345646;
      44239: inst = 32'd203423744;
      44240: inst = 32'd471859200;
      44241: inst = 32'd136314880;
      44242: inst = 32'd268468224;
      44243: inst = 32'd201345647;
      44244: inst = 32'd203423744;
      44245: inst = 32'd471859200;
      44246: inst = 32'd136314880;
      44247: inst = 32'd268468224;
      44248: inst = 32'd201345648;
      44249: inst = 32'd203423744;
      44250: inst = 32'd471859200;
      44251: inst = 32'd136314880;
      44252: inst = 32'd268468224;
      44253: inst = 32'd201345649;
      44254: inst = 32'd203423744;
      44255: inst = 32'd471859200;
      44256: inst = 32'd136314880;
      44257: inst = 32'd268468224;
      44258: inst = 32'd201345650;
      44259: inst = 32'd203423744;
      44260: inst = 32'd471859200;
      44261: inst = 32'd136314880;
      44262: inst = 32'd268468224;
      44263: inst = 32'd201345651;
      44264: inst = 32'd203423744;
      44265: inst = 32'd471859200;
      44266: inst = 32'd136314880;
      44267: inst = 32'd268468224;
      44268: inst = 32'd201345652;
      44269: inst = 32'd203423744;
      44270: inst = 32'd471859200;
      44271: inst = 32'd136314880;
      44272: inst = 32'd268468224;
      44273: inst = 32'd201345653;
      44274: inst = 32'd203423744;
      44275: inst = 32'd471859200;
      44276: inst = 32'd136314880;
      44277: inst = 32'd268468224;
      44278: inst = 32'd201345654;
      44279: inst = 32'd203423744;
      44280: inst = 32'd471859200;
      44281: inst = 32'd136314880;
      44282: inst = 32'd268468224;
      44283: inst = 32'd201345655;
      44284: inst = 32'd203423744;
      44285: inst = 32'd471859200;
      44286: inst = 32'd136314880;
      44287: inst = 32'd268468224;
      44288: inst = 32'd201345656;
      44289: inst = 32'd203423744;
      44290: inst = 32'd471859200;
      44291: inst = 32'd136314880;
      44292: inst = 32'd268468224;
      44293: inst = 32'd201345657;
      44294: inst = 32'd203423744;
      44295: inst = 32'd471859200;
      44296: inst = 32'd136314880;
      44297: inst = 32'd268468224;
      44298: inst = 32'd201345658;
      44299: inst = 32'd203423744;
      44300: inst = 32'd471859200;
      44301: inst = 32'd136314880;
      44302: inst = 32'd268468224;
      44303: inst = 32'd201345659;
      44304: inst = 32'd203423744;
      44305: inst = 32'd471859200;
      44306: inst = 32'd136314880;
      44307: inst = 32'd268468224;
      44308: inst = 32'd201345660;
      44309: inst = 32'd203423744;
      44310: inst = 32'd471859200;
      44311: inst = 32'd136314880;
      44312: inst = 32'd268468224;
      44313: inst = 32'd201345661;
      44314: inst = 32'd203423744;
      44315: inst = 32'd471859200;
      44316: inst = 32'd136314880;
      44317: inst = 32'd268468224;
      44318: inst = 32'd201345662;
      44319: inst = 32'd203423744;
      44320: inst = 32'd471859200;
      44321: inst = 32'd136314880;
      44322: inst = 32'd268468224;
      44323: inst = 32'd201345663;
      44324: inst = 32'd203423744;
      44325: inst = 32'd471859200;
      44326: inst = 32'd136314880;
      44327: inst = 32'd268468224;
      44328: inst = 32'd201345664;
      44329: inst = 32'd203423744;
      44330: inst = 32'd471859200;
      44331: inst = 32'd136314880;
      44332: inst = 32'd268468224;
      44333: inst = 32'd201345665;
      44334: inst = 32'd203423744;
      44335: inst = 32'd471859200;
      44336: inst = 32'd136314880;
      44337: inst = 32'd268468224;
      44338: inst = 32'd201345666;
      44339: inst = 32'd203423744;
      44340: inst = 32'd471859200;
      44341: inst = 32'd136314880;
      44342: inst = 32'd268468224;
      44343: inst = 32'd201345667;
      44344: inst = 32'd203423744;
      44345: inst = 32'd471859200;
      44346: inst = 32'd136314880;
      44347: inst = 32'd268468224;
      44348: inst = 32'd201345668;
      44349: inst = 32'd203423744;
      44350: inst = 32'd471859200;
      44351: inst = 32'd136314880;
      44352: inst = 32'd268468224;
      44353: inst = 32'd201345669;
      44354: inst = 32'd203423744;
      44355: inst = 32'd471859200;
      44356: inst = 32'd136314880;
      44357: inst = 32'd268468224;
      44358: inst = 32'd201345670;
      44359: inst = 32'd203423744;
      44360: inst = 32'd471859200;
      44361: inst = 32'd136314880;
      44362: inst = 32'd268468224;
      44363: inst = 32'd201345671;
      44364: inst = 32'd203423744;
      44365: inst = 32'd471859200;
      44366: inst = 32'd136314880;
      44367: inst = 32'd268468224;
      44368: inst = 32'd201345672;
      44369: inst = 32'd203423744;
      44370: inst = 32'd471859200;
      44371: inst = 32'd136314880;
      44372: inst = 32'd268468224;
      44373: inst = 32'd201345673;
      44374: inst = 32'd203423744;
      44375: inst = 32'd471859200;
      44376: inst = 32'd136314880;
      44377: inst = 32'd268468224;
      44378: inst = 32'd201345674;
      44379: inst = 32'd203423744;
      44380: inst = 32'd471859200;
      44381: inst = 32'd136314880;
      44382: inst = 32'd268468224;
      44383: inst = 32'd201345675;
      44384: inst = 32'd203423744;
      44385: inst = 32'd471859200;
      44386: inst = 32'd136314880;
      44387: inst = 32'd268468224;
      44388: inst = 32'd201345676;
      44389: inst = 32'd203423744;
      44390: inst = 32'd471859200;
      44391: inst = 32'd136314880;
      44392: inst = 32'd268468224;
      44393: inst = 32'd201345677;
      44394: inst = 32'd203423744;
      44395: inst = 32'd471859200;
      44396: inst = 32'd136314880;
      44397: inst = 32'd268468224;
      44398: inst = 32'd201345678;
      44399: inst = 32'd203423744;
      44400: inst = 32'd471859200;
      44401: inst = 32'd136314880;
      44402: inst = 32'd268468224;
      44403: inst = 32'd201345679;
      44404: inst = 32'd203423744;
      44405: inst = 32'd471859200;
      44406: inst = 32'd136314880;
      44407: inst = 32'd268468224;
      44408: inst = 32'd201345680;
      44409: inst = 32'd203423744;
      44410: inst = 32'd471859200;
      44411: inst = 32'd136314880;
      44412: inst = 32'd268468224;
      44413: inst = 32'd201345681;
      44414: inst = 32'd203423744;
      44415: inst = 32'd471859200;
      44416: inst = 32'd136314880;
      44417: inst = 32'd268468224;
      44418: inst = 32'd201345682;
      44419: inst = 32'd203423744;
      44420: inst = 32'd471859200;
      44421: inst = 32'd136314880;
      44422: inst = 32'd268468224;
      44423: inst = 32'd201345683;
      44424: inst = 32'd203423744;
      44425: inst = 32'd471859200;
      44426: inst = 32'd136314880;
      44427: inst = 32'd268468224;
      44428: inst = 32'd201345684;
      44429: inst = 32'd203423744;
      44430: inst = 32'd471859200;
      44431: inst = 32'd136314880;
      44432: inst = 32'd268468224;
      44433: inst = 32'd201345685;
      44434: inst = 32'd203423744;
      44435: inst = 32'd471859200;
      44436: inst = 32'd136314880;
      44437: inst = 32'd268468224;
      44438: inst = 32'd201345686;
      44439: inst = 32'd203423744;
      44440: inst = 32'd471859200;
      44441: inst = 32'd136314880;
      44442: inst = 32'd268468224;
      44443: inst = 32'd201345687;
      44444: inst = 32'd203423744;
      44445: inst = 32'd471859200;
      44446: inst = 32'd136314880;
      44447: inst = 32'd268468224;
      44448: inst = 32'd201345688;
      44449: inst = 32'd203423744;
      44450: inst = 32'd471859200;
      44451: inst = 32'd136314880;
      44452: inst = 32'd268468224;
      44453: inst = 32'd201345689;
      44454: inst = 32'd203423744;
      44455: inst = 32'd471859200;
      44456: inst = 32'd136314880;
      44457: inst = 32'd268468224;
      44458: inst = 32'd201345690;
      44459: inst = 32'd203423744;
      44460: inst = 32'd471859200;
      44461: inst = 32'd136314880;
      44462: inst = 32'd268468224;
      44463: inst = 32'd201345691;
      44464: inst = 32'd203423744;
      44465: inst = 32'd471859200;
      44466: inst = 32'd136314880;
      44467: inst = 32'd268468224;
      44468: inst = 32'd201345692;
      44469: inst = 32'd203423744;
      44470: inst = 32'd471859200;
      44471: inst = 32'd136314880;
      44472: inst = 32'd268468224;
      44473: inst = 32'd201345693;
      44474: inst = 32'd203423744;
      44475: inst = 32'd471859200;
      44476: inst = 32'd136314880;
      44477: inst = 32'd268468224;
      44478: inst = 32'd201345694;
      44479: inst = 32'd203423744;
      44480: inst = 32'd471859200;
      44481: inst = 32'd136314880;
      44482: inst = 32'd268468224;
      44483: inst = 32'd201345695;
      44484: inst = 32'd203423744;
      44485: inst = 32'd471859200;
      44486: inst = 32'd136314880;
      44487: inst = 32'd268468224;
      44488: inst = 32'd201345696;
      44489: inst = 32'd203423744;
      44490: inst = 32'd471859200;
      44491: inst = 32'd136314880;
      44492: inst = 32'd268468224;
      44493: inst = 32'd201345697;
      44494: inst = 32'd203423744;
      44495: inst = 32'd471859200;
      44496: inst = 32'd136314880;
      44497: inst = 32'd268468224;
      44498: inst = 32'd201345698;
      44499: inst = 32'd203423744;
      44500: inst = 32'd471859200;
      44501: inst = 32'd136314880;
      44502: inst = 32'd268468224;
      44503: inst = 32'd201345699;
      44504: inst = 32'd203423744;
      44505: inst = 32'd471859200;
      44506: inst = 32'd136314880;
      44507: inst = 32'd268468224;
      44508: inst = 32'd201345700;
      44509: inst = 32'd203423744;
      44510: inst = 32'd471859200;
      44511: inst = 32'd136314880;
      44512: inst = 32'd268468224;
      44513: inst = 32'd201345701;
      44514: inst = 32'd203423744;
      44515: inst = 32'd471859200;
      44516: inst = 32'd136314880;
      44517: inst = 32'd268468224;
      44518: inst = 32'd201345702;
      44519: inst = 32'd203423744;
      44520: inst = 32'd471859200;
      44521: inst = 32'd136314880;
      44522: inst = 32'd268468224;
      44523: inst = 32'd201345703;
      44524: inst = 32'd203423744;
      44525: inst = 32'd471859200;
      44526: inst = 32'd136314880;
      44527: inst = 32'd268468224;
      44528: inst = 32'd201345704;
      44529: inst = 32'd203423744;
      44530: inst = 32'd471859200;
      44531: inst = 32'd136314880;
      44532: inst = 32'd268468224;
      44533: inst = 32'd201345705;
      44534: inst = 32'd203423744;
      44535: inst = 32'd471859200;
      44536: inst = 32'd136314880;
      44537: inst = 32'd268468224;
      44538: inst = 32'd201345706;
      44539: inst = 32'd203423744;
      44540: inst = 32'd471859200;
      44541: inst = 32'd136314880;
      44542: inst = 32'd268468224;
      44543: inst = 32'd201345707;
      44544: inst = 32'd203423744;
      44545: inst = 32'd471859200;
      44546: inst = 32'd136314880;
      44547: inst = 32'd268468224;
      44548: inst = 32'd201345708;
      44549: inst = 32'd203423744;
      44550: inst = 32'd471859200;
      44551: inst = 32'd136314880;
      44552: inst = 32'd268468224;
      44553: inst = 32'd201345709;
      44554: inst = 32'd203423744;
      44555: inst = 32'd471859200;
      44556: inst = 32'd136314880;
      44557: inst = 32'd268468224;
      44558: inst = 32'd201345710;
      44559: inst = 32'd203423744;
      44560: inst = 32'd471859200;
      44561: inst = 32'd136314880;
      44562: inst = 32'd268468224;
      44563: inst = 32'd201345711;
      44564: inst = 32'd203423744;
      44565: inst = 32'd471859200;
      44566: inst = 32'd136314880;
      44567: inst = 32'd268468224;
      44568: inst = 32'd201345712;
      44569: inst = 32'd203423744;
      44570: inst = 32'd471859200;
      44571: inst = 32'd136314880;
      44572: inst = 32'd268468224;
      44573: inst = 32'd201345713;
      44574: inst = 32'd203423744;
      44575: inst = 32'd471859200;
      44576: inst = 32'd136314880;
      44577: inst = 32'd268468224;
      44578: inst = 32'd201345714;
      44579: inst = 32'd203423744;
      44580: inst = 32'd471859200;
      44581: inst = 32'd136314880;
      44582: inst = 32'd268468224;
      44583: inst = 32'd201345715;
      44584: inst = 32'd203423744;
      44585: inst = 32'd471859200;
      44586: inst = 32'd136314880;
      44587: inst = 32'd268468224;
      44588: inst = 32'd201345716;
      44589: inst = 32'd203423744;
      44590: inst = 32'd471859200;
      44591: inst = 32'd136314880;
      44592: inst = 32'd268468224;
      44593: inst = 32'd201345717;
      44594: inst = 32'd203423744;
      44595: inst = 32'd471859200;
      44596: inst = 32'd136314880;
      44597: inst = 32'd268468224;
      44598: inst = 32'd201345718;
      44599: inst = 32'd203423744;
      44600: inst = 32'd471859200;
      44601: inst = 32'd136314880;
      44602: inst = 32'd268468224;
      44603: inst = 32'd201345719;
      44604: inst = 32'd203423744;
      44605: inst = 32'd471859200;
      44606: inst = 32'd136314880;
      44607: inst = 32'd268468224;
      44608: inst = 32'd201345720;
      44609: inst = 32'd203423744;
      44610: inst = 32'd471859200;
      44611: inst = 32'd136314880;
      44612: inst = 32'd268468224;
      44613: inst = 32'd201345721;
      44614: inst = 32'd203423744;
      44615: inst = 32'd471859200;
      44616: inst = 32'd136314880;
      44617: inst = 32'd268468224;
      44618: inst = 32'd201345722;
      44619: inst = 32'd203423744;
      44620: inst = 32'd471859200;
      44621: inst = 32'd136314880;
      44622: inst = 32'd268468224;
      44623: inst = 32'd201345723;
      44624: inst = 32'd203423744;
      44625: inst = 32'd471859200;
      44626: inst = 32'd136314880;
      44627: inst = 32'd268468224;
      44628: inst = 32'd201345724;
      44629: inst = 32'd203423744;
      44630: inst = 32'd471859200;
      44631: inst = 32'd136314880;
      44632: inst = 32'd268468224;
      44633: inst = 32'd201345725;
      44634: inst = 32'd203423744;
      44635: inst = 32'd471859200;
      44636: inst = 32'd136314880;
      44637: inst = 32'd268468224;
      44638: inst = 32'd201345726;
      44639: inst = 32'd203423744;
      44640: inst = 32'd471859200;
      44641: inst = 32'd136314880;
      44642: inst = 32'd268468224;
      44643: inst = 32'd201345727;
      44644: inst = 32'd203423744;
      44645: inst = 32'd471859200;
      44646: inst = 32'd136314880;
      44647: inst = 32'd268468224;
      44648: inst = 32'd201345728;
      44649: inst = 32'd203423744;
      44650: inst = 32'd471859200;
      44651: inst = 32'd136314880;
      44652: inst = 32'd268468224;
      44653: inst = 32'd201345729;
      44654: inst = 32'd203423744;
      44655: inst = 32'd471859200;
      44656: inst = 32'd136314880;
      44657: inst = 32'd268468224;
      44658: inst = 32'd201345730;
      44659: inst = 32'd203423744;
      44660: inst = 32'd471859200;
      44661: inst = 32'd136314880;
      44662: inst = 32'd268468224;
      44663: inst = 32'd201345731;
      44664: inst = 32'd203423744;
      44665: inst = 32'd471859200;
      44666: inst = 32'd136314880;
      44667: inst = 32'd268468224;
      44668: inst = 32'd201345732;
      44669: inst = 32'd203423744;
      44670: inst = 32'd471859200;
      44671: inst = 32'd136314880;
      44672: inst = 32'd268468224;
      44673: inst = 32'd201345733;
      44674: inst = 32'd203423744;
      44675: inst = 32'd471859200;
      44676: inst = 32'd136314880;
      44677: inst = 32'd268468224;
      44678: inst = 32'd201345734;
      44679: inst = 32'd203423744;
      44680: inst = 32'd471859200;
      44681: inst = 32'd136314880;
      44682: inst = 32'd268468224;
      44683: inst = 32'd201345735;
      44684: inst = 32'd203423744;
      44685: inst = 32'd471859200;
      44686: inst = 32'd136314880;
      44687: inst = 32'd268468224;
      44688: inst = 32'd201345736;
      44689: inst = 32'd203423744;
      44690: inst = 32'd471859200;
      44691: inst = 32'd136314880;
      44692: inst = 32'd268468224;
      44693: inst = 32'd201345737;
      44694: inst = 32'd203423744;
      44695: inst = 32'd471859200;
      44696: inst = 32'd136314880;
      44697: inst = 32'd268468224;
      44698: inst = 32'd201345738;
      44699: inst = 32'd203423744;
      44700: inst = 32'd471859200;
      44701: inst = 32'd136314880;
      44702: inst = 32'd268468224;
      44703: inst = 32'd201345739;
      44704: inst = 32'd203423744;
      44705: inst = 32'd471859200;
      44706: inst = 32'd136314880;
      44707: inst = 32'd268468224;
      44708: inst = 32'd201345740;
      44709: inst = 32'd203423744;
      44710: inst = 32'd471859200;
      44711: inst = 32'd136314880;
      44712: inst = 32'd268468224;
      44713: inst = 32'd201345741;
      44714: inst = 32'd203423744;
      44715: inst = 32'd471859200;
      44716: inst = 32'd136314880;
      44717: inst = 32'd268468224;
      44718: inst = 32'd201345742;
      44719: inst = 32'd203423744;
      44720: inst = 32'd471859200;
      44721: inst = 32'd136314880;
      44722: inst = 32'd268468224;
      44723: inst = 32'd201345743;
      44724: inst = 32'd203423744;
      44725: inst = 32'd471859200;
      44726: inst = 32'd136314880;
      44727: inst = 32'd268468224;
      44728: inst = 32'd201345744;
      44729: inst = 32'd203423744;
      44730: inst = 32'd471859200;
      44731: inst = 32'd136314880;
      44732: inst = 32'd268468224;
      44733: inst = 32'd201345745;
      44734: inst = 32'd203423744;
      44735: inst = 32'd471859200;
      44736: inst = 32'd136314880;
      44737: inst = 32'd268468224;
      44738: inst = 32'd201345746;
      44739: inst = 32'd203423744;
      44740: inst = 32'd471859200;
      44741: inst = 32'd136314880;
      44742: inst = 32'd268468224;
      44743: inst = 32'd201345747;
      44744: inst = 32'd203423744;
      44745: inst = 32'd471859200;
      44746: inst = 32'd136314880;
      44747: inst = 32'd268468224;
      44748: inst = 32'd201345748;
      44749: inst = 32'd203423744;
      44750: inst = 32'd471859200;
      44751: inst = 32'd136314880;
      44752: inst = 32'd268468224;
      44753: inst = 32'd201345749;
      44754: inst = 32'd203423744;
      44755: inst = 32'd471859200;
      44756: inst = 32'd136314880;
      44757: inst = 32'd268468224;
      44758: inst = 32'd201345750;
      44759: inst = 32'd203423744;
      44760: inst = 32'd471859200;
      44761: inst = 32'd136314880;
      44762: inst = 32'd268468224;
      44763: inst = 32'd201345751;
      44764: inst = 32'd203423744;
      44765: inst = 32'd471859200;
      44766: inst = 32'd136314880;
      44767: inst = 32'd268468224;
      44768: inst = 32'd201345752;
      44769: inst = 32'd203423744;
      44770: inst = 32'd471859200;
      44771: inst = 32'd136314880;
      44772: inst = 32'd268468224;
      44773: inst = 32'd201345753;
      44774: inst = 32'd203423744;
      44775: inst = 32'd471859200;
      44776: inst = 32'd136314880;
      44777: inst = 32'd268468224;
      44778: inst = 32'd201345754;
      44779: inst = 32'd203423744;
      44780: inst = 32'd471859200;
      44781: inst = 32'd136314880;
      44782: inst = 32'd268468224;
      44783: inst = 32'd201345755;
      44784: inst = 32'd203423744;
      44785: inst = 32'd471859200;
      44786: inst = 32'd136314880;
      44787: inst = 32'd268468224;
      44788: inst = 32'd201345756;
      44789: inst = 32'd203423744;
      44790: inst = 32'd471859200;
      44791: inst = 32'd136314880;
      44792: inst = 32'd268468224;
      44793: inst = 32'd201345757;
      44794: inst = 32'd203423744;
      44795: inst = 32'd471859200;
      44796: inst = 32'd136314880;
      44797: inst = 32'd268468224;
      44798: inst = 32'd201345758;
      44799: inst = 32'd203423744;
      44800: inst = 32'd471859200;
      44801: inst = 32'd136314880;
      44802: inst = 32'd268468224;
      44803: inst = 32'd201345759;
      44804: inst = 32'd203423744;
      44805: inst = 32'd471859200;
      44806: inst = 32'd136314880;
      44807: inst = 32'd268468224;
      44808: inst = 32'd201345760;
      44809: inst = 32'd203423744;
      44810: inst = 32'd471859200;
      44811: inst = 32'd136314880;
      44812: inst = 32'd268468224;
      44813: inst = 32'd201345761;
      44814: inst = 32'd203423744;
      44815: inst = 32'd471859200;
      44816: inst = 32'd136314880;
      44817: inst = 32'd268468224;
      44818: inst = 32'd201345762;
      44819: inst = 32'd203423744;
      44820: inst = 32'd471859200;
      44821: inst = 32'd136314880;
      44822: inst = 32'd268468224;
      44823: inst = 32'd201345763;
      44824: inst = 32'd203423744;
      44825: inst = 32'd471859200;
      44826: inst = 32'd136314880;
      44827: inst = 32'd268468224;
      44828: inst = 32'd201345764;
      44829: inst = 32'd203423744;
      44830: inst = 32'd471859200;
      44831: inst = 32'd136314880;
      44832: inst = 32'd268468224;
      44833: inst = 32'd201345765;
      44834: inst = 32'd203423744;
      44835: inst = 32'd471859200;
      44836: inst = 32'd136314880;
      44837: inst = 32'd268468224;
      44838: inst = 32'd201345766;
      44839: inst = 32'd203423744;
      44840: inst = 32'd471859200;
      44841: inst = 32'd136314880;
      44842: inst = 32'd268468224;
      44843: inst = 32'd201345767;
      44844: inst = 32'd203423744;
      44845: inst = 32'd471859200;
      44846: inst = 32'd136314880;
      44847: inst = 32'd268468224;
      44848: inst = 32'd201345768;
      44849: inst = 32'd203423744;
      44850: inst = 32'd471859200;
      44851: inst = 32'd136314880;
      44852: inst = 32'd268468224;
      44853: inst = 32'd201345769;
      44854: inst = 32'd203423744;
      44855: inst = 32'd471859200;
      44856: inst = 32'd136314880;
      44857: inst = 32'd268468224;
      44858: inst = 32'd201345770;
      44859: inst = 32'd203423744;
      44860: inst = 32'd471859200;
      44861: inst = 32'd136314880;
      44862: inst = 32'd268468224;
      44863: inst = 32'd201345771;
      44864: inst = 32'd203423744;
      44865: inst = 32'd471859200;
      44866: inst = 32'd136314880;
      44867: inst = 32'd268468224;
      44868: inst = 32'd201345772;
      44869: inst = 32'd203423744;
      44870: inst = 32'd471859200;
      44871: inst = 32'd136314880;
      44872: inst = 32'd268468224;
      44873: inst = 32'd201345773;
      44874: inst = 32'd203423744;
      44875: inst = 32'd471859200;
      44876: inst = 32'd136314880;
      44877: inst = 32'd268468224;
      44878: inst = 32'd201345774;
      44879: inst = 32'd203423744;
      44880: inst = 32'd471859200;
      44881: inst = 32'd136314880;
      44882: inst = 32'd268468224;
      44883: inst = 32'd201345775;
      44884: inst = 32'd203423744;
      44885: inst = 32'd471859200;
      44886: inst = 32'd136314880;
      44887: inst = 32'd268468224;
      44888: inst = 32'd201345776;
      44889: inst = 32'd203423744;
      44890: inst = 32'd471859200;
      44891: inst = 32'd136314880;
      44892: inst = 32'd268468224;
      44893: inst = 32'd201345777;
      44894: inst = 32'd203423744;
      44895: inst = 32'd471859200;
      44896: inst = 32'd136314880;
      44897: inst = 32'd268468224;
      44898: inst = 32'd201345778;
      44899: inst = 32'd203423744;
      44900: inst = 32'd471859200;
      44901: inst = 32'd136314880;
      44902: inst = 32'd268468224;
      44903: inst = 32'd201345779;
      44904: inst = 32'd203423744;
      44905: inst = 32'd471859200;
      44906: inst = 32'd136314880;
      44907: inst = 32'd268468224;
      44908: inst = 32'd201345780;
      44909: inst = 32'd203423744;
      44910: inst = 32'd471859200;
      44911: inst = 32'd136314880;
      44912: inst = 32'd268468224;
      44913: inst = 32'd201345781;
      44914: inst = 32'd203423744;
      44915: inst = 32'd471859200;
      44916: inst = 32'd136314880;
      44917: inst = 32'd268468224;
      44918: inst = 32'd201345782;
      44919: inst = 32'd203423744;
      44920: inst = 32'd471859200;
      44921: inst = 32'd136314880;
      44922: inst = 32'd268468224;
      44923: inst = 32'd201345783;
      44924: inst = 32'd203423744;
      44925: inst = 32'd471859200;
      44926: inst = 32'd136314880;
      44927: inst = 32'd268468224;
      44928: inst = 32'd201345784;
      44929: inst = 32'd203423744;
      44930: inst = 32'd471859200;
      44931: inst = 32'd136314880;
      44932: inst = 32'd268468224;
      44933: inst = 32'd201345785;
      44934: inst = 32'd203423744;
      44935: inst = 32'd471859200;
      44936: inst = 32'd136314880;
      44937: inst = 32'd268468224;
      44938: inst = 32'd201345786;
      44939: inst = 32'd203423744;
      44940: inst = 32'd471859200;
      44941: inst = 32'd136314880;
      44942: inst = 32'd268468224;
      44943: inst = 32'd201345787;
      44944: inst = 32'd203423744;
      44945: inst = 32'd471859200;
      44946: inst = 32'd136314880;
      44947: inst = 32'd268468224;
      44948: inst = 32'd201345788;
      44949: inst = 32'd203423744;
      44950: inst = 32'd471859200;
      44951: inst = 32'd136314880;
      44952: inst = 32'd268468224;
      44953: inst = 32'd201345789;
      44954: inst = 32'd203423744;
      44955: inst = 32'd471859200;
      44956: inst = 32'd136314880;
      44957: inst = 32'd268468224;
      44958: inst = 32'd201345790;
      44959: inst = 32'd203423744;
      44960: inst = 32'd471859200;
      44961: inst = 32'd136314880;
      44962: inst = 32'd268468224;
      44963: inst = 32'd201345791;
      44964: inst = 32'd203423744;
      44965: inst = 32'd471859200;
      44966: inst = 32'd136314880;
      44967: inst = 32'd268468224;
      44968: inst = 32'd201345792;
      44969: inst = 32'd203423744;
      44970: inst = 32'd471859200;
      44971: inst = 32'd136314880;
      44972: inst = 32'd268468224;
      44973: inst = 32'd201345793;
      44974: inst = 32'd203423744;
      44975: inst = 32'd471859200;
      44976: inst = 32'd136314880;
      44977: inst = 32'd268468224;
      44978: inst = 32'd201345794;
      44979: inst = 32'd203423744;
      44980: inst = 32'd471859200;
      44981: inst = 32'd136314880;
      44982: inst = 32'd268468224;
      44983: inst = 32'd201345795;
      44984: inst = 32'd203423744;
      44985: inst = 32'd471859200;
      44986: inst = 32'd136314880;
      44987: inst = 32'd268468224;
      44988: inst = 32'd201345796;
      44989: inst = 32'd203423744;
      44990: inst = 32'd471859200;
      44991: inst = 32'd136314880;
      44992: inst = 32'd268468224;
      44993: inst = 32'd201345797;
      44994: inst = 32'd203423744;
      44995: inst = 32'd471859200;
      44996: inst = 32'd136314880;
      44997: inst = 32'd268468224;
      44998: inst = 32'd201345798;
      44999: inst = 32'd203423744;
      45000: inst = 32'd471859200;
      45001: inst = 32'd136314880;
      45002: inst = 32'd268468224;
      45003: inst = 32'd201345799;
      45004: inst = 32'd203423744;
      45005: inst = 32'd471859200;
      45006: inst = 32'd136314880;
      45007: inst = 32'd268468224;
      45008: inst = 32'd201345800;
      45009: inst = 32'd203423744;
      45010: inst = 32'd471859200;
      45011: inst = 32'd136314880;
      45012: inst = 32'd268468224;
      45013: inst = 32'd201345801;
      45014: inst = 32'd203423744;
      45015: inst = 32'd471859200;
      45016: inst = 32'd136314880;
      45017: inst = 32'd268468224;
      45018: inst = 32'd201345802;
      45019: inst = 32'd203423744;
      45020: inst = 32'd471859200;
      45021: inst = 32'd136314880;
      45022: inst = 32'd268468224;
      45023: inst = 32'd201345803;
      45024: inst = 32'd203423744;
      45025: inst = 32'd471859200;
      45026: inst = 32'd136314880;
      45027: inst = 32'd268468224;
      45028: inst = 32'd201345804;
      45029: inst = 32'd203423744;
      45030: inst = 32'd471859200;
      45031: inst = 32'd136314880;
      45032: inst = 32'd268468224;
      45033: inst = 32'd201345805;
      45034: inst = 32'd203423744;
      45035: inst = 32'd471859200;
      45036: inst = 32'd136314880;
      45037: inst = 32'd268468224;
      45038: inst = 32'd201345806;
      45039: inst = 32'd203423744;
      45040: inst = 32'd471859200;
      45041: inst = 32'd136314880;
      45042: inst = 32'd268468224;
      45043: inst = 32'd201345807;
      45044: inst = 32'd203423744;
      45045: inst = 32'd471859200;
      45046: inst = 32'd136314880;
      45047: inst = 32'd268468224;
      45048: inst = 32'd201345808;
      45049: inst = 32'd203423744;
      45050: inst = 32'd471859200;
      45051: inst = 32'd136314880;
      45052: inst = 32'd268468224;
      45053: inst = 32'd201345809;
      45054: inst = 32'd203423744;
      45055: inst = 32'd471859200;
      45056: inst = 32'd136314880;
      45057: inst = 32'd268468224;
      45058: inst = 32'd201345810;
      45059: inst = 32'd203423744;
      45060: inst = 32'd471859200;
      45061: inst = 32'd136314880;
      45062: inst = 32'd268468224;
      45063: inst = 32'd201345811;
      45064: inst = 32'd203423744;
      45065: inst = 32'd471859200;
      45066: inst = 32'd136314880;
      45067: inst = 32'd268468224;
      45068: inst = 32'd201345812;
      45069: inst = 32'd203423744;
      45070: inst = 32'd471859200;
      45071: inst = 32'd136314880;
      45072: inst = 32'd268468224;
      45073: inst = 32'd201345813;
      45074: inst = 32'd203423744;
      45075: inst = 32'd471859200;
      45076: inst = 32'd136314880;
      45077: inst = 32'd268468224;
      45078: inst = 32'd201345814;
      45079: inst = 32'd203423744;
      45080: inst = 32'd471859200;
      45081: inst = 32'd136314880;
      45082: inst = 32'd268468224;
      45083: inst = 32'd201345815;
      45084: inst = 32'd203423744;
      45085: inst = 32'd471859200;
      45086: inst = 32'd136314880;
      45087: inst = 32'd268468224;
      45088: inst = 32'd201345816;
      45089: inst = 32'd203423744;
      45090: inst = 32'd471859200;
      45091: inst = 32'd136314880;
      45092: inst = 32'd268468224;
      45093: inst = 32'd201345817;
      45094: inst = 32'd203423744;
      45095: inst = 32'd471859200;
      45096: inst = 32'd136314880;
      45097: inst = 32'd268468224;
      45098: inst = 32'd201345818;
      45099: inst = 32'd203423744;
      45100: inst = 32'd471859200;
      45101: inst = 32'd136314880;
      45102: inst = 32'd268468224;
      45103: inst = 32'd201345819;
      45104: inst = 32'd203423744;
      45105: inst = 32'd471859200;
      45106: inst = 32'd136314880;
      45107: inst = 32'd268468224;
      45108: inst = 32'd201345820;
      45109: inst = 32'd203423744;
      45110: inst = 32'd471859200;
      45111: inst = 32'd136314880;
      45112: inst = 32'd268468224;
      45113: inst = 32'd201345821;
      45114: inst = 32'd203423744;
      45115: inst = 32'd471859200;
      45116: inst = 32'd136314880;
      45117: inst = 32'd268468224;
      45118: inst = 32'd201345822;
      45119: inst = 32'd203423744;
      45120: inst = 32'd471859200;
      45121: inst = 32'd136314880;
      45122: inst = 32'd268468224;
      45123: inst = 32'd201345823;
      45124: inst = 32'd203423744;
      45125: inst = 32'd471859200;
      45126: inst = 32'd136314880;
      45127: inst = 32'd268468224;
      45128: inst = 32'd201345824;
      45129: inst = 32'd203423744;
      45130: inst = 32'd471859200;
      45131: inst = 32'd136314880;
      45132: inst = 32'd268468224;
      45133: inst = 32'd201345825;
      45134: inst = 32'd203423744;
      45135: inst = 32'd471859200;
      45136: inst = 32'd136314880;
      45137: inst = 32'd268468224;
      45138: inst = 32'd201345826;
      45139: inst = 32'd203423744;
      45140: inst = 32'd471859200;
      45141: inst = 32'd136314880;
      45142: inst = 32'd268468224;
      45143: inst = 32'd201345827;
      45144: inst = 32'd203423744;
      45145: inst = 32'd471859200;
      45146: inst = 32'd136314880;
      45147: inst = 32'd268468224;
      45148: inst = 32'd201345828;
      45149: inst = 32'd203423744;
      45150: inst = 32'd471859200;
      45151: inst = 32'd136314880;
      45152: inst = 32'd268468224;
      45153: inst = 32'd201345829;
      45154: inst = 32'd203423744;
      45155: inst = 32'd471859200;
      45156: inst = 32'd136314880;
      45157: inst = 32'd268468224;
      45158: inst = 32'd201345830;
      45159: inst = 32'd203423744;
      45160: inst = 32'd471859200;
      45161: inst = 32'd136314880;
      45162: inst = 32'd268468224;
      45163: inst = 32'd201345831;
      45164: inst = 32'd203423744;
      45165: inst = 32'd471859200;
      45166: inst = 32'd136314880;
      45167: inst = 32'd268468224;
      45168: inst = 32'd201345832;
      45169: inst = 32'd203423744;
      45170: inst = 32'd471859200;
      45171: inst = 32'd136314880;
      45172: inst = 32'd268468224;
      45173: inst = 32'd201345833;
      45174: inst = 32'd203423744;
      45175: inst = 32'd471859200;
      45176: inst = 32'd136314880;
      45177: inst = 32'd268468224;
      45178: inst = 32'd201345834;
      45179: inst = 32'd203423744;
      45180: inst = 32'd471859200;
      45181: inst = 32'd136314880;
      45182: inst = 32'd268468224;
      45183: inst = 32'd201345835;
      45184: inst = 32'd203423744;
      45185: inst = 32'd471859200;
      45186: inst = 32'd136314880;
      45187: inst = 32'd268468224;
      45188: inst = 32'd201345836;
      45189: inst = 32'd203423744;
      45190: inst = 32'd471859200;
      45191: inst = 32'd136314880;
      45192: inst = 32'd268468224;
      45193: inst = 32'd201345837;
      45194: inst = 32'd203423744;
      45195: inst = 32'd471859200;
      45196: inst = 32'd136314880;
      45197: inst = 32'd268468224;
      45198: inst = 32'd201345838;
      45199: inst = 32'd203423744;
      45200: inst = 32'd471859200;
      45201: inst = 32'd136314880;
      45202: inst = 32'd268468224;
      45203: inst = 32'd201345839;
      45204: inst = 32'd203423744;
      45205: inst = 32'd471859200;
      45206: inst = 32'd136314880;
      45207: inst = 32'd268468224;
      45208: inst = 32'd201345840;
      45209: inst = 32'd203423744;
      45210: inst = 32'd471859200;
      45211: inst = 32'd136314880;
      45212: inst = 32'd268468224;
      45213: inst = 32'd201345841;
      45214: inst = 32'd203423744;
      45215: inst = 32'd471859200;
      45216: inst = 32'd136314880;
      45217: inst = 32'd268468224;
      45218: inst = 32'd201345842;
      45219: inst = 32'd203423744;
      45220: inst = 32'd471859200;
      45221: inst = 32'd136314880;
      45222: inst = 32'd268468224;
      45223: inst = 32'd201345843;
      45224: inst = 32'd203423744;
      45225: inst = 32'd471859200;
      45226: inst = 32'd136314880;
      45227: inst = 32'd268468224;
      45228: inst = 32'd201345844;
      45229: inst = 32'd203423744;
      45230: inst = 32'd471859200;
      45231: inst = 32'd136314880;
      45232: inst = 32'd268468224;
      45233: inst = 32'd201345845;
      45234: inst = 32'd203423744;
      45235: inst = 32'd471859200;
      45236: inst = 32'd136314880;
      45237: inst = 32'd268468224;
      45238: inst = 32'd201345846;
      45239: inst = 32'd203423744;
      45240: inst = 32'd471859200;
      45241: inst = 32'd136314880;
      45242: inst = 32'd268468224;
      45243: inst = 32'd201345847;
      45244: inst = 32'd203423744;
      45245: inst = 32'd471859200;
      45246: inst = 32'd136314880;
      45247: inst = 32'd268468224;
      45248: inst = 32'd201345848;
      45249: inst = 32'd203423744;
      45250: inst = 32'd471859200;
      45251: inst = 32'd136314880;
      45252: inst = 32'd268468224;
      45253: inst = 32'd201345849;
      45254: inst = 32'd203423744;
      45255: inst = 32'd471859200;
      45256: inst = 32'd136314880;
      45257: inst = 32'd268468224;
      45258: inst = 32'd201345850;
      45259: inst = 32'd203423744;
      45260: inst = 32'd471859200;
      45261: inst = 32'd136314880;
      45262: inst = 32'd268468224;
      45263: inst = 32'd201345851;
      45264: inst = 32'd203423744;
      45265: inst = 32'd471859200;
      45266: inst = 32'd136314880;
      45267: inst = 32'd268468224;
      45268: inst = 32'd201345852;
      45269: inst = 32'd203423744;
      45270: inst = 32'd471859200;
      45271: inst = 32'd136314880;
      45272: inst = 32'd268468224;
      45273: inst = 32'd201345853;
      45274: inst = 32'd203423744;
      45275: inst = 32'd471859200;
      45276: inst = 32'd136314880;
      45277: inst = 32'd268468224;
      45278: inst = 32'd201345854;
      45279: inst = 32'd203423744;
      45280: inst = 32'd471859200;
      45281: inst = 32'd136314880;
      45282: inst = 32'd268468224;
      45283: inst = 32'd201345855;
      45284: inst = 32'd203423744;
      45285: inst = 32'd471859200;
      45286: inst = 32'd136314880;
      45287: inst = 32'd268468224;
      45288: inst = 32'd201345856;
      45289: inst = 32'd203423744;
      45290: inst = 32'd471859200;
      45291: inst = 32'd136314880;
      45292: inst = 32'd268468224;
      45293: inst = 32'd201345857;
      45294: inst = 32'd203423744;
      45295: inst = 32'd471859200;
      45296: inst = 32'd136314880;
      45297: inst = 32'd268468224;
      45298: inst = 32'd201345858;
      45299: inst = 32'd203423744;
      45300: inst = 32'd471859200;
      45301: inst = 32'd136314880;
      45302: inst = 32'd268468224;
      45303: inst = 32'd201345859;
      45304: inst = 32'd203423744;
      45305: inst = 32'd471859200;
      45306: inst = 32'd136314880;
      45307: inst = 32'd268468224;
      45308: inst = 32'd201345860;
      45309: inst = 32'd203423744;
      45310: inst = 32'd471859200;
      45311: inst = 32'd136314880;
      45312: inst = 32'd268468224;
      45313: inst = 32'd201345861;
      45314: inst = 32'd203423744;
      45315: inst = 32'd471859200;
      45316: inst = 32'd136314880;
      45317: inst = 32'd268468224;
      45318: inst = 32'd201345862;
      45319: inst = 32'd203423744;
      45320: inst = 32'd471859200;
      45321: inst = 32'd136314880;
      45322: inst = 32'd268468224;
      45323: inst = 32'd201345863;
      45324: inst = 32'd203423744;
      45325: inst = 32'd471859200;
      45326: inst = 32'd136314880;
      45327: inst = 32'd268468224;
      45328: inst = 32'd201345864;
      45329: inst = 32'd203423744;
      45330: inst = 32'd471859200;
      45331: inst = 32'd136314880;
      45332: inst = 32'd268468224;
      45333: inst = 32'd201345865;
      45334: inst = 32'd203423744;
      45335: inst = 32'd471859200;
      45336: inst = 32'd136314880;
      45337: inst = 32'd268468224;
      45338: inst = 32'd201345866;
      45339: inst = 32'd203423744;
      45340: inst = 32'd471859200;
      45341: inst = 32'd136314880;
      45342: inst = 32'd268468224;
      45343: inst = 32'd201345867;
      45344: inst = 32'd203423744;
      45345: inst = 32'd471859200;
      45346: inst = 32'd136314880;
      45347: inst = 32'd268468224;
      45348: inst = 32'd201345868;
      45349: inst = 32'd203423744;
      45350: inst = 32'd471859200;
      45351: inst = 32'd136314880;
      45352: inst = 32'd268468224;
      45353: inst = 32'd201345869;
      45354: inst = 32'd203423744;
      45355: inst = 32'd471859200;
      45356: inst = 32'd136314880;
      45357: inst = 32'd268468224;
      45358: inst = 32'd201345870;
      45359: inst = 32'd203423744;
      45360: inst = 32'd471859200;
      45361: inst = 32'd136314880;
      45362: inst = 32'd268468224;
      45363: inst = 32'd201345871;
      45364: inst = 32'd203423744;
      45365: inst = 32'd471859200;
      45366: inst = 32'd136314880;
      45367: inst = 32'd268468224;
      45368: inst = 32'd201345872;
      45369: inst = 32'd203423744;
      45370: inst = 32'd471859200;
      45371: inst = 32'd136314880;
      45372: inst = 32'd268468224;
      45373: inst = 32'd201345873;
      45374: inst = 32'd203423744;
      45375: inst = 32'd471859200;
      45376: inst = 32'd136314880;
      45377: inst = 32'd268468224;
      45378: inst = 32'd201345874;
      45379: inst = 32'd203423744;
      45380: inst = 32'd471859200;
      45381: inst = 32'd136314880;
      45382: inst = 32'd268468224;
      45383: inst = 32'd201345875;
      45384: inst = 32'd203423744;
      45385: inst = 32'd471859200;
      45386: inst = 32'd136314880;
      45387: inst = 32'd268468224;
      45388: inst = 32'd201345876;
      45389: inst = 32'd203423744;
      45390: inst = 32'd471859200;
      45391: inst = 32'd136314880;
      45392: inst = 32'd268468224;
      45393: inst = 32'd201345877;
      45394: inst = 32'd203423744;
      45395: inst = 32'd471859200;
      45396: inst = 32'd136314880;
      45397: inst = 32'd268468224;
      45398: inst = 32'd201345878;
      45399: inst = 32'd203423744;
      45400: inst = 32'd471859200;
      45401: inst = 32'd136314880;
      45402: inst = 32'd268468224;
      45403: inst = 32'd201345879;
      45404: inst = 32'd203423744;
      45405: inst = 32'd471859200;
      45406: inst = 32'd136314880;
      45407: inst = 32'd268468224;
      45408: inst = 32'd201345880;
      45409: inst = 32'd203423744;
      45410: inst = 32'd471859200;
      45411: inst = 32'd136314880;
      45412: inst = 32'd268468224;
      45413: inst = 32'd201345881;
      45414: inst = 32'd203423744;
      45415: inst = 32'd471859200;
      45416: inst = 32'd136314880;
      45417: inst = 32'd268468224;
      45418: inst = 32'd201345882;
      45419: inst = 32'd203423744;
      45420: inst = 32'd471859200;
      45421: inst = 32'd136314880;
      45422: inst = 32'd268468224;
      45423: inst = 32'd201345883;
      45424: inst = 32'd203423744;
      45425: inst = 32'd471859200;
      45426: inst = 32'd136314880;
      45427: inst = 32'd268468224;
      45428: inst = 32'd201345884;
      45429: inst = 32'd203423744;
      45430: inst = 32'd471859200;
      45431: inst = 32'd136314880;
      45432: inst = 32'd268468224;
      45433: inst = 32'd201345885;
      45434: inst = 32'd203423744;
      45435: inst = 32'd471859200;
      45436: inst = 32'd136314880;
      45437: inst = 32'd268468224;
      45438: inst = 32'd201345886;
      45439: inst = 32'd203423744;
      45440: inst = 32'd471859200;
      45441: inst = 32'd136314880;
      45442: inst = 32'd268468224;
      45443: inst = 32'd201345887;
      45444: inst = 32'd203423744;
      45445: inst = 32'd471859200;
      45446: inst = 32'd136314880;
      45447: inst = 32'd268468224;
      45448: inst = 32'd201345888;
      45449: inst = 32'd203423744;
      45450: inst = 32'd471859200;
      45451: inst = 32'd136314880;
      45452: inst = 32'd268468224;
      45453: inst = 32'd201345889;
      45454: inst = 32'd203423744;
      45455: inst = 32'd471859200;
      45456: inst = 32'd136314880;
      45457: inst = 32'd268468224;
      45458: inst = 32'd201345890;
      45459: inst = 32'd203423744;
      45460: inst = 32'd471859200;
      45461: inst = 32'd136314880;
      45462: inst = 32'd268468224;
      45463: inst = 32'd201345891;
      45464: inst = 32'd203423744;
      45465: inst = 32'd471859200;
      45466: inst = 32'd136314880;
      45467: inst = 32'd268468224;
      45468: inst = 32'd201345892;
      45469: inst = 32'd203423744;
      45470: inst = 32'd471859200;
      45471: inst = 32'd136314880;
      45472: inst = 32'd268468224;
      45473: inst = 32'd201345893;
      45474: inst = 32'd203423744;
      45475: inst = 32'd471859200;
      45476: inst = 32'd136314880;
      45477: inst = 32'd268468224;
      45478: inst = 32'd201345894;
      45479: inst = 32'd203423744;
      45480: inst = 32'd471859200;
      45481: inst = 32'd136314880;
      45482: inst = 32'd268468224;
      45483: inst = 32'd201345895;
      45484: inst = 32'd203423744;
      45485: inst = 32'd471859200;
      45486: inst = 32'd136314880;
      45487: inst = 32'd268468224;
      45488: inst = 32'd201345896;
      45489: inst = 32'd203423744;
      45490: inst = 32'd471859200;
      45491: inst = 32'd136314880;
      45492: inst = 32'd268468224;
      45493: inst = 32'd201345897;
      45494: inst = 32'd203423744;
      45495: inst = 32'd471859200;
      45496: inst = 32'd136314880;
      45497: inst = 32'd268468224;
      45498: inst = 32'd201345898;
      45499: inst = 32'd203423744;
      45500: inst = 32'd471859200;
      45501: inst = 32'd136314880;
      45502: inst = 32'd268468224;
      45503: inst = 32'd201345899;
      45504: inst = 32'd203423744;
      45505: inst = 32'd471859200;
      45506: inst = 32'd136314880;
      45507: inst = 32'd268468224;
      45508: inst = 32'd201345900;
      45509: inst = 32'd203423744;
      45510: inst = 32'd471859200;
      45511: inst = 32'd136314880;
      45512: inst = 32'd268468224;
      45513: inst = 32'd201345901;
      45514: inst = 32'd203423744;
      45515: inst = 32'd471859200;
      45516: inst = 32'd136314880;
      45517: inst = 32'd268468224;
      45518: inst = 32'd201345902;
      45519: inst = 32'd203423744;
      45520: inst = 32'd471859200;
      45521: inst = 32'd136314880;
      45522: inst = 32'd268468224;
      45523: inst = 32'd201345903;
      45524: inst = 32'd203423744;
      45525: inst = 32'd471859200;
      45526: inst = 32'd136314880;
      45527: inst = 32'd268468224;
      45528: inst = 32'd201345904;
      45529: inst = 32'd203423744;
      45530: inst = 32'd471859200;
      45531: inst = 32'd136314880;
      45532: inst = 32'd268468224;
      45533: inst = 32'd201345905;
      45534: inst = 32'd203423744;
      45535: inst = 32'd471859200;
      45536: inst = 32'd136314880;
      45537: inst = 32'd268468224;
      45538: inst = 32'd201345906;
      45539: inst = 32'd203423744;
      45540: inst = 32'd471859200;
      45541: inst = 32'd136314880;
      45542: inst = 32'd268468224;
      45543: inst = 32'd201345907;
      45544: inst = 32'd203423744;
      45545: inst = 32'd471859200;
      45546: inst = 32'd136314880;
      45547: inst = 32'd268468224;
      45548: inst = 32'd201345908;
      45549: inst = 32'd203423744;
      45550: inst = 32'd471859200;
      45551: inst = 32'd136314880;
      45552: inst = 32'd268468224;
      45553: inst = 32'd201345909;
      45554: inst = 32'd203423744;
      45555: inst = 32'd471859200;
      45556: inst = 32'd136314880;
      45557: inst = 32'd268468224;
      45558: inst = 32'd201345910;
      45559: inst = 32'd203423744;
      45560: inst = 32'd471859200;
      45561: inst = 32'd136314880;
      45562: inst = 32'd268468224;
      45563: inst = 32'd201345911;
      45564: inst = 32'd203423744;
      45565: inst = 32'd471859200;
      45566: inst = 32'd136314880;
      45567: inst = 32'd268468224;
      45568: inst = 32'd201345912;
      45569: inst = 32'd203423744;
      45570: inst = 32'd471859200;
      45571: inst = 32'd136314880;
      45572: inst = 32'd268468224;
      45573: inst = 32'd201345913;
      45574: inst = 32'd203423744;
      45575: inst = 32'd471859200;
      45576: inst = 32'd136314880;
      45577: inst = 32'd268468224;
      45578: inst = 32'd201345914;
      45579: inst = 32'd203423744;
      45580: inst = 32'd471859200;
      45581: inst = 32'd136314880;
      45582: inst = 32'd268468224;
      45583: inst = 32'd201345915;
      45584: inst = 32'd203423744;
      45585: inst = 32'd471859200;
      45586: inst = 32'd136314880;
      45587: inst = 32'd268468224;
      45588: inst = 32'd201345916;
      45589: inst = 32'd203423744;
      45590: inst = 32'd471859200;
      45591: inst = 32'd136314880;
      45592: inst = 32'd268468224;
      45593: inst = 32'd201345917;
      45594: inst = 32'd203423744;
      45595: inst = 32'd471859200;
      45596: inst = 32'd136314880;
      45597: inst = 32'd268468224;
      45598: inst = 32'd201345918;
      45599: inst = 32'd203423744;
      45600: inst = 32'd471859200;
      45601: inst = 32'd136314880;
      45602: inst = 32'd268468224;
      45603: inst = 32'd201345919;
      45604: inst = 32'd203423744;
      45605: inst = 32'd471859200;
      45606: inst = 32'd136314880;
      45607: inst = 32'd268468224;
      45608: inst = 32'd201345920;
      45609: inst = 32'd203423744;
      45610: inst = 32'd471859200;
      45611: inst = 32'd136314880;
      45612: inst = 32'd268468224;
      45613: inst = 32'd201345921;
      45614: inst = 32'd203423744;
      45615: inst = 32'd471859200;
      45616: inst = 32'd136314880;
      45617: inst = 32'd268468224;
      45618: inst = 32'd201345922;
      45619: inst = 32'd203423744;
      45620: inst = 32'd471859200;
      45621: inst = 32'd136314880;
      45622: inst = 32'd268468224;
      45623: inst = 32'd201345923;
      45624: inst = 32'd203423744;
      45625: inst = 32'd471859200;
      45626: inst = 32'd136314880;
      45627: inst = 32'd268468224;
      45628: inst = 32'd201345924;
      45629: inst = 32'd203423744;
      45630: inst = 32'd471859200;
      45631: inst = 32'd136314880;
      45632: inst = 32'd268468224;
      45633: inst = 32'd201345925;
      45634: inst = 32'd203423744;
      45635: inst = 32'd471859200;
      45636: inst = 32'd136314880;
      45637: inst = 32'd268468224;
      45638: inst = 32'd201345926;
      45639: inst = 32'd203423744;
      45640: inst = 32'd471859200;
      45641: inst = 32'd136314880;
      45642: inst = 32'd268468224;
      45643: inst = 32'd201345927;
      45644: inst = 32'd203423744;
      45645: inst = 32'd471859200;
      45646: inst = 32'd136314880;
      45647: inst = 32'd268468224;
      45648: inst = 32'd201345928;
      45649: inst = 32'd203423744;
      45650: inst = 32'd471859200;
      45651: inst = 32'd136314880;
      45652: inst = 32'd268468224;
      45653: inst = 32'd201345929;
      45654: inst = 32'd203423744;
      45655: inst = 32'd471859200;
      45656: inst = 32'd136314880;
      45657: inst = 32'd268468224;
      45658: inst = 32'd201345930;
      45659: inst = 32'd203423744;
      45660: inst = 32'd471859200;
      45661: inst = 32'd136314880;
      45662: inst = 32'd268468224;
      45663: inst = 32'd201345931;
      45664: inst = 32'd203423744;
      45665: inst = 32'd471859200;
      45666: inst = 32'd136314880;
      45667: inst = 32'd268468224;
      45668: inst = 32'd201345932;
      45669: inst = 32'd203423744;
      45670: inst = 32'd471859200;
      45671: inst = 32'd136314880;
      45672: inst = 32'd268468224;
      45673: inst = 32'd201345933;
      45674: inst = 32'd203423744;
      45675: inst = 32'd471859200;
      45676: inst = 32'd136314880;
      45677: inst = 32'd268468224;
      45678: inst = 32'd201345934;
      45679: inst = 32'd203423744;
      45680: inst = 32'd471859200;
      45681: inst = 32'd136314880;
      45682: inst = 32'd268468224;
      45683: inst = 32'd201345935;
      45684: inst = 32'd203423744;
      45685: inst = 32'd471859200;
      45686: inst = 32'd136314880;
      45687: inst = 32'd268468224;
      45688: inst = 32'd201345936;
      45689: inst = 32'd203423744;
      45690: inst = 32'd471859200;
      45691: inst = 32'd136314880;
      45692: inst = 32'd268468224;
      45693: inst = 32'd201345937;
      45694: inst = 32'd203423744;
      45695: inst = 32'd471859200;
      45696: inst = 32'd136314880;
      45697: inst = 32'd268468224;
      45698: inst = 32'd201345938;
      45699: inst = 32'd203423744;
      45700: inst = 32'd471859200;
      45701: inst = 32'd136314880;
      45702: inst = 32'd268468224;
      45703: inst = 32'd201345939;
      45704: inst = 32'd203423744;
      45705: inst = 32'd471859200;
      45706: inst = 32'd136314880;
      45707: inst = 32'd268468224;
      45708: inst = 32'd201345940;
      45709: inst = 32'd203423744;
      45710: inst = 32'd471859200;
      45711: inst = 32'd136314880;
      45712: inst = 32'd268468224;
      45713: inst = 32'd201345941;
      45714: inst = 32'd203423744;
      45715: inst = 32'd471859200;
      45716: inst = 32'd136314880;
      45717: inst = 32'd268468224;
      45718: inst = 32'd201345942;
      45719: inst = 32'd203423744;
      45720: inst = 32'd471859200;
      45721: inst = 32'd136314880;
      45722: inst = 32'd268468224;
      45723: inst = 32'd201345943;
      45724: inst = 32'd203423744;
      45725: inst = 32'd471859200;
      45726: inst = 32'd136314880;
      45727: inst = 32'd268468224;
      45728: inst = 32'd201345944;
      45729: inst = 32'd203423744;
      45730: inst = 32'd471859200;
      45731: inst = 32'd136314880;
      45732: inst = 32'd268468224;
      45733: inst = 32'd201345945;
      45734: inst = 32'd203423744;
      45735: inst = 32'd471859200;
      45736: inst = 32'd136314880;
      45737: inst = 32'd268468224;
      45738: inst = 32'd201345946;
      45739: inst = 32'd203423744;
      45740: inst = 32'd471859200;
      45741: inst = 32'd136314880;
      45742: inst = 32'd268468224;
      45743: inst = 32'd201345947;
      45744: inst = 32'd203423744;
      45745: inst = 32'd471859200;
      45746: inst = 32'd136314880;
      45747: inst = 32'd268468224;
      45748: inst = 32'd201345948;
      45749: inst = 32'd203423744;
      45750: inst = 32'd471859200;
      45751: inst = 32'd136314880;
      45752: inst = 32'd268468224;
      45753: inst = 32'd201345949;
      45754: inst = 32'd203423744;
      45755: inst = 32'd471859200;
      45756: inst = 32'd136314880;
      45757: inst = 32'd268468224;
      45758: inst = 32'd201345950;
      45759: inst = 32'd203423744;
      45760: inst = 32'd471859200;
      45761: inst = 32'd136314880;
      45762: inst = 32'd268468224;
      45763: inst = 32'd201345951;
      45764: inst = 32'd203423744;
      45765: inst = 32'd471859200;
      45766: inst = 32'd136314880;
      45767: inst = 32'd268468224;
      45768: inst = 32'd201345952;
      45769: inst = 32'd203423744;
      45770: inst = 32'd471859200;
      45771: inst = 32'd136314880;
      45772: inst = 32'd268468224;
      45773: inst = 32'd201345953;
      45774: inst = 32'd203423744;
      45775: inst = 32'd471859200;
      45776: inst = 32'd136314880;
      45777: inst = 32'd268468224;
      45778: inst = 32'd201345954;
      45779: inst = 32'd203423744;
      45780: inst = 32'd471859200;
      45781: inst = 32'd136314880;
      45782: inst = 32'd268468224;
      45783: inst = 32'd201345955;
      45784: inst = 32'd203423744;
      45785: inst = 32'd471859200;
      45786: inst = 32'd136314880;
      45787: inst = 32'd268468224;
      45788: inst = 32'd201345956;
      45789: inst = 32'd203423744;
      45790: inst = 32'd471859200;
      45791: inst = 32'd136314880;
      45792: inst = 32'd268468224;
      45793: inst = 32'd201345957;
      45794: inst = 32'd203423744;
      45795: inst = 32'd471859200;
      45796: inst = 32'd136314880;
      45797: inst = 32'd268468224;
      45798: inst = 32'd201345958;
      45799: inst = 32'd203423744;
      45800: inst = 32'd471859200;
      45801: inst = 32'd136314880;
      45802: inst = 32'd268468224;
      45803: inst = 32'd201345959;
      45804: inst = 32'd203423744;
      45805: inst = 32'd471859200;
      45806: inst = 32'd136314880;
      45807: inst = 32'd268468224;
      45808: inst = 32'd201345960;
      45809: inst = 32'd203423744;
      45810: inst = 32'd471859200;
      45811: inst = 32'd136314880;
      45812: inst = 32'd268468224;
      45813: inst = 32'd201345961;
      45814: inst = 32'd203423744;
      45815: inst = 32'd471859200;
      45816: inst = 32'd136314880;
      45817: inst = 32'd268468224;
      45818: inst = 32'd201345962;
      45819: inst = 32'd203423744;
      45820: inst = 32'd471859200;
      45821: inst = 32'd136314880;
      45822: inst = 32'd268468224;
      45823: inst = 32'd201345963;
      45824: inst = 32'd203423744;
      45825: inst = 32'd471859200;
      45826: inst = 32'd136314880;
      45827: inst = 32'd268468224;
      45828: inst = 32'd201345964;
      45829: inst = 32'd203423744;
      45830: inst = 32'd471859200;
      45831: inst = 32'd136314880;
      45832: inst = 32'd268468224;
      45833: inst = 32'd201345965;
      45834: inst = 32'd203423744;
      45835: inst = 32'd471859200;
      45836: inst = 32'd136314880;
      45837: inst = 32'd268468224;
      45838: inst = 32'd201345966;
      45839: inst = 32'd203423744;
      45840: inst = 32'd471859200;
      45841: inst = 32'd136314880;
      45842: inst = 32'd268468224;
      45843: inst = 32'd201345967;
      45844: inst = 32'd203423744;
      45845: inst = 32'd471859200;
      45846: inst = 32'd136314880;
      45847: inst = 32'd268468224;
      45848: inst = 32'd201345968;
      45849: inst = 32'd203423744;
      45850: inst = 32'd471859200;
      45851: inst = 32'd136314880;
      45852: inst = 32'd268468224;
      45853: inst = 32'd201345969;
      45854: inst = 32'd203423744;
      45855: inst = 32'd471859200;
      45856: inst = 32'd136314880;
      45857: inst = 32'd268468224;
      45858: inst = 32'd201345970;
      45859: inst = 32'd203423744;
      45860: inst = 32'd471859200;
      45861: inst = 32'd136314880;
      45862: inst = 32'd268468224;
      45863: inst = 32'd201345971;
      45864: inst = 32'd203423744;
      45865: inst = 32'd471859200;
      45866: inst = 32'd136314880;
      45867: inst = 32'd268468224;
      45868: inst = 32'd201345972;
      45869: inst = 32'd203423744;
      45870: inst = 32'd471859200;
      45871: inst = 32'd136314880;
      45872: inst = 32'd268468224;
      45873: inst = 32'd201345973;
      45874: inst = 32'd203423744;
      45875: inst = 32'd471859200;
      45876: inst = 32'd136314880;
      45877: inst = 32'd268468224;
      45878: inst = 32'd201345974;
      45879: inst = 32'd203423744;
      45880: inst = 32'd471859200;
      45881: inst = 32'd136314880;
      45882: inst = 32'd268468224;
      45883: inst = 32'd201345975;
      45884: inst = 32'd203423744;
      45885: inst = 32'd471859200;
      45886: inst = 32'd136314880;
      45887: inst = 32'd268468224;
      45888: inst = 32'd201345976;
      45889: inst = 32'd203423744;
      45890: inst = 32'd471859200;
      45891: inst = 32'd136314880;
      45892: inst = 32'd268468224;
      45893: inst = 32'd201345977;
      45894: inst = 32'd203423744;
      45895: inst = 32'd471859200;
      45896: inst = 32'd136314880;
      45897: inst = 32'd268468224;
      45898: inst = 32'd201345978;
      45899: inst = 32'd203423744;
      45900: inst = 32'd471859200;
      45901: inst = 32'd136314880;
      45902: inst = 32'd268468224;
      45903: inst = 32'd201345979;
      45904: inst = 32'd203423744;
      45905: inst = 32'd471859200;
      45906: inst = 32'd136314880;
      45907: inst = 32'd268468224;
      45908: inst = 32'd201345980;
      45909: inst = 32'd203423744;
      45910: inst = 32'd471859200;
      45911: inst = 32'd136314880;
      45912: inst = 32'd268468224;
      45913: inst = 32'd201345981;
      45914: inst = 32'd203423744;
      45915: inst = 32'd471859200;
      45916: inst = 32'd136314880;
      45917: inst = 32'd268468224;
      45918: inst = 32'd201345982;
      45919: inst = 32'd203423744;
      45920: inst = 32'd471859200;
      45921: inst = 32'd136314880;
      45922: inst = 32'd268468224;
      45923: inst = 32'd201345983;
      45924: inst = 32'd203423744;
      45925: inst = 32'd471859200;
      45926: inst = 32'd136314880;
      45927: inst = 32'd268468224;
      45928: inst = 32'd201345984;
      45929: inst = 32'd203423744;
      45930: inst = 32'd471859200;
      45931: inst = 32'd136314880;
      45932: inst = 32'd268468224;
      45933: inst = 32'd201345985;
      45934: inst = 32'd203423744;
      45935: inst = 32'd471859200;
      45936: inst = 32'd136314880;
      45937: inst = 32'd268468224;
      45938: inst = 32'd201345986;
      45939: inst = 32'd203423744;
      45940: inst = 32'd471859200;
      45941: inst = 32'd136314880;
      45942: inst = 32'd268468224;
      45943: inst = 32'd201345987;
      45944: inst = 32'd203423744;
      45945: inst = 32'd471859200;
      45946: inst = 32'd136314880;
      45947: inst = 32'd268468224;
      45948: inst = 32'd201345988;
      45949: inst = 32'd203423744;
      45950: inst = 32'd471859200;
      45951: inst = 32'd136314880;
      45952: inst = 32'd268468224;
      45953: inst = 32'd201345989;
      45954: inst = 32'd203423744;
      45955: inst = 32'd471859200;
      45956: inst = 32'd136314880;
      45957: inst = 32'd268468224;
      45958: inst = 32'd201345990;
      45959: inst = 32'd203423744;
      45960: inst = 32'd471859200;
      45961: inst = 32'd136314880;
      45962: inst = 32'd268468224;
      45963: inst = 32'd201345991;
      45964: inst = 32'd203423744;
      45965: inst = 32'd471859200;
      45966: inst = 32'd136314880;
      45967: inst = 32'd268468224;
      45968: inst = 32'd201345992;
      45969: inst = 32'd203423744;
      45970: inst = 32'd471859200;
      45971: inst = 32'd136314880;
      45972: inst = 32'd268468224;
      45973: inst = 32'd201345993;
      45974: inst = 32'd203423744;
      45975: inst = 32'd471859200;
      45976: inst = 32'd136314880;
      45977: inst = 32'd268468224;
      45978: inst = 32'd201345994;
      45979: inst = 32'd203423744;
      45980: inst = 32'd471859200;
      45981: inst = 32'd136314880;
      45982: inst = 32'd268468224;
      45983: inst = 32'd201345995;
      45984: inst = 32'd203423744;
      45985: inst = 32'd471859200;
      45986: inst = 32'd136314880;
      45987: inst = 32'd268468224;
      45988: inst = 32'd201345996;
      45989: inst = 32'd203423744;
      45990: inst = 32'd471859200;
      45991: inst = 32'd136314880;
      45992: inst = 32'd268468224;
      45993: inst = 32'd201345997;
      45994: inst = 32'd203423744;
      45995: inst = 32'd471859200;
      45996: inst = 32'd136314880;
      45997: inst = 32'd268468224;
      45998: inst = 32'd201345998;
      45999: inst = 32'd203423744;
      46000: inst = 32'd471859200;
      46001: inst = 32'd136314880;
      46002: inst = 32'd268468224;
      46003: inst = 32'd201345999;
      46004: inst = 32'd203423744;
      46005: inst = 32'd471859200;
      46006: inst = 32'd136314880;
      46007: inst = 32'd268468224;
      46008: inst = 32'd201346000;
      46009: inst = 32'd203423744;
      46010: inst = 32'd471859200;
      46011: inst = 32'd136314880;
      46012: inst = 32'd268468224;
      46013: inst = 32'd201346001;
      46014: inst = 32'd203423744;
      46015: inst = 32'd471859200;
      46016: inst = 32'd136314880;
      46017: inst = 32'd268468224;
      46018: inst = 32'd201346002;
      46019: inst = 32'd203423744;
      46020: inst = 32'd471859200;
      46021: inst = 32'd136314880;
      46022: inst = 32'd268468224;
      46023: inst = 32'd201346003;
      46024: inst = 32'd203423744;
      46025: inst = 32'd471859200;
      46026: inst = 32'd136314880;
      46027: inst = 32'd268468224;
      46028: inst = 32'd201346004;
      46029: inst = 32'd203423744;
      46030: inst = 32'd471859200;
      46031: inst = 32'd136314880;
      46032: inst = 32'd268468224;
      46033: inst = 32'd201346005;
      46034: inst = 32'd203423744;
      46035: inst = 32'd471859200;
      46036: inst = 32'd136314880;
      46037: inst = 32'd268468224;
      46038: inst = 32'd201346006;
      46039: inst = 32'd203423744;
      46040: inst = 32'd471859200;
      46041: inst = 32'd136314880;
      46042: inst = 32'd268468224;
      46043: inst = 32'd201346007;
      46044: inst = 32'd203423744;
      46045: inst = 32'd471859200;
      46046: inst = 32'd136314880;
      46047: inst = 32'd268468224;
      46048: inst = 32'd201346008;
      46049: inst = 32'd203423744;
      46050: inst = 32'd471859200;
      46051: inst = 32'd136314880;
      46052: inst = 32'd268468224;
      46053: inst = 32'd201346009;
      46054: inst = 32'd203423744;
      46055: inst = 32'd471859200;
      46056: inst = 32'd136314880;
      46057: inst = 32'd268468224;
      46058: inst = 32'd201346010;
      46059: inst = 32'd203423744;
      46060: inst = 32'd471859200;
      46061: inst = 32'd136314880;
      46062: inst = 32'd268468224;
      46063: inst = 32'd201346011;
      46064: inst = 32'd203423744;
      46065: inst = 32'd471859200;
      46066: inst = 32'd136314880;
      46067: inst = 32'd268468224;
      46068: inst = 32'd201346012;
      46069: inst = 32'd203423744;
      46070: inst = 32'd471859200;
      46071: inst = 32'd136314880;
      46072: inst = 32'd268468224;
      46073: inst = 32'd201346013;
      46074: inst = 32'd203423744;
      46075: inst = 32'd471859200;
      46076: inst = 32'd136314880;
      46077: inst = 32'd268468224;
      46078: inst = 32'd201346014;
      46079: inst = 32'd203423744;
      46080: inst = 32'd471859200;
      46081: inst = 32'd136314880;
      46082: inst = 32'd268468224;
      46083: inst = 32'd201346015;
      46084: inst = 32'd203423744;
      46085: inst = 32'd471859200;
      46086: inst = 32'd136314880;
      46087: inst = 32'd268468224;
      46088: inst = 32'd201346016;
      46089: inst = 32'd203423744;
      46090: inst = 32'd471859200;
      46091: inst = 32'd136314880;
      46092: inst = 32'd268468224;
      46093: inst = 32'd201346017;
      46094: inst = 32'd203423744;
      46095: inst = 32'd471859200;
      46096: inst = 32'd136314880;
      46097: inst = 32'd268468224;
      46098: inst = 32'd201346018;
      46099: inst = 32'd203423744;
      46100: inst = 32'd471859200;
      46101: inst = 32'd136314880;
      46102: inst = 32'd268468224;
      46103: inst = 32'd201346019;
      46104: inst = 32'd203423744;
      46105: inst = 32'd471859200;
      46106: inst = 32'd136314880;
      46107: inst = 32'd268468224;
      46108: inst = 32'd201346020;
      46109: inst = 32'd203423744;
      46110: inst = 32'd471859200;
      46111: inst = 32'd136314880;
      46112: inst = 32'd268468224;
      46113: inst = 32'd201346021;
      46114: inst = 32'd203423744;
      46115: inst = 32'd471859200;
      46116: inst = 32'd136314880;
      46117: inst = 32'd268468224;
      46118: inst = 32'd201346022;
      46119: inst = 32'd203423744;
      46120: inst = 32'd471859200;
      46121: inst = 32'd136314880;
      46122: inst = 32'd268468224;
      46123: inst = 32'd201346023;
      46124: inst = 32'd203423744;
      46125: inst = 32'd471859200;
      46126: inst = 32'd136314880;
      46127: inst = 32'd268468224;
      46128: inst = 32'd201346024;
      46129: inst = 32'd203423744;
      46130: inst = 32'd471859200;
      46131: inst = 32'd136314880;
      46132: inst = 32'd268468224;
      46133: inst = 32'd201346025;
      46134: inst = 32'd203423744;
      46135: inst = 32'd471859200;
      46136: inst = 32'd136314880;
      46137: inst = 32'd268468224;
      46138: inst = 32'd201346026;
      46139: inst = 32'd203423744;
      46140: inst = 32'd471859200;
      46141: inst = 32'd136314880;
      46142: inst = 32'd268468224;
      46143: inst = 32'd201346027;
      46144: inst = 32'd203423744;
      46145: inst = 32'd471859200;
      46146: inst = 32'd136314880;
      46147: inst = 32'd268468224;
      46148: inst = 32'd201346028;
      46149: inst = 32'd203423744;
      46150: inst = 32'd471859200;
      46151: inst = 32'd136314880;
      46152: inst = 32'd268468224;
      46153: inst = 32'd201346029;
      46154: inst = 32'd203423744;
      46155: inst = 32'd471859200;
      46156: inst = 32'd136314880;
      46157: inst = 32'd268468224;
      46158: inst = 32'd201346030;
      46159: inst = 32'd203483685;
      46160: inst = 32'd471859200;
      46161: inst = 32'd136314880;
      46162: inst = 32'd268468224;
      46163: inst = 32'd201346031;
      46164: inst = 32'd203483685;
      46165: inst = 32'd471859200;
      46166: inst = 32'd136314880;
      46167: inst = 32'd268468224;
      46168: inst = 32'd201346032;
      46169: inst = 32'd203483685;
      46170: inst = 32'd471859200;
      46171: inst = 32'd136314880;
      46172: inst = 32'd268468224;
      46173: inst = 32'd201346033;
      46174: inst = 32'd203483685;
      46175: inst = 32'd471859200;
      46176: inst = 32'd136314880;
      46177: inst = 32'd268468224;
      46178: inst = 32'd201346034;
      46179: inst = 32'd203483685;
      46180: inst = 32'd471859200;
      46181: inst = 32'd136314880;
      46182: inst = 32'd268468224;
      46183: inst = 32'd201346035;
      46184: inst = 32'd203483685;
      46185: inst = 32'd471859200;
      46186: inst = 32'd136314880;
      46187: inst = 32'd268468224;
      46188: inst = 32'd201346036;
      46189: inst = 32'd203483685;
      46190: inst = 32'd471859200;
      46191: inst = 32'd136314880;
      46192: inst = 32'd268468224;
      46193: inst = 32'd201346037;
      46194: inst = 32'd203483685;
      46195: inst = 32'd471859200;
      46196: inst = 32'd136314880;
      46197: inst = 32'd268468224;
      46198: inst = 32'd201346038;
      46199: inst = 32'd203483685;
      46200: inst = 32'd471859200;
      46201: inst = 32'd136314880;
      46202: inst = 32'd268468224;
      46203: inst = 32'd201346039;
      46204: inst = 32'd203483685;
      46205: inst = 32'd471859200;
      46206: inst = 32'd136314880;
      46207: inst = 32'd268468224;
      46208: inst = 32'd201346040;
      46209: inst = 32'd203483685;
      46210: inst = 32'd471859200;
      46211: inst = 32'd136314880;
      46212: inst = 32'd268468224;
      46213: inst = 32'd201346041;
      46214: inst = 32'd203483685;
      46215: inst = 32'd471859200;
      46216: inst = 32'd136314880;
      46217: inst = 32'd268468224;
      46218: inst = 32'd201346042;
      46219: inst = 32'd203483685;
      46220: inst = 32'd471859200;
      46221: inst = 32'd136314880;
      46222: inst = 32'd268468224;
      46223: inst = 32'd201346043;
      46224: inst = 32'd203483685;
      46225: inst = 32'd471859200;
      46226: inst = 32'd136314880;
      46227: inst = 32'd268468224;
      46228: inst = 32'd201346044;
      46229: inst = 32'd203483685;
      46230: inst = 32'd471859200;
      46231: inst = 32'd136314880;
      46232: inst = 32'd268468224;
      46233: inst = 32'd201346045;
      46234: inst = 32'd203483685;
      46235: inst = 32'd471859200;
      46236: inst = 32'd136314880;
      46237: inst = 32'd268468224;
      46238: inst = 32'd201346046;
      46239: inst = 32'd203483685;
      46240: inst = 32'd471859200;
      46241: inst = 32'd136314880;
      46242: inst = 32'd268468224;
      46243: inst = 32'd201346047;
      46244: inst = 32'd203483685;
      46245: inst = 32'd471859200;
      46246: inst = 32'd136314880;
      46247: inst = 32'd268468224;
      46248: inst = 32'd201346048;
      46249: inst = 32'd203483685;
      46250: inst = 32'd471859200;
      46251: inst = 32'd136314880;
      46252: inst = 32'd268468224;
      46253: inst = 32'd201346049;
      46254: inst = 32'd203483685;
      46255: inst = 32'd471859200;
      46256: inst = 32'd136314880;
      46257: inst = 32'd268468224;
      46258: inst = 32'd201346050;
      46259: inst = 32'd203483685;
      46260: inst = 32'd471859200;
      46261: inst = 32'd136314880;
      46262: inst = 32'd268468224;
      46263: inst = 32'd201346051;
      46264: inst = 32'd203483685;
      46265: inst = 32'd471859200;
      46266: inst = 32'd136314880;
      46267: inst = 32'd268468224;
      46268: inst = 32'd201346052;
      46269: inst = 32'd203483685;
      46270: inst = 32'd471859200;
      46271: inst = 32'd136314880;
      46272: inst = 32'd268468224;
      46273: inst = 32'd201346053;
      46274: inst = 32'd203483685;
      46275: inst = 32'd471859200;
      46276: inst = 32'd136314880;
      46277: inst = 32'd268468224;
      46278: inst = 32'd201346054;
      46279: inst = 32'd203483685;
      46280: inst = 32'd471859200;
      46281: inst = 32'd136314880;
      46282: inst = 32'd268468224;
      46283: inst = 32'd201346055;
      46284: inst = 32'd203483685;
      46285: inst = 32'd471859200;
      46286: inst = 32'd136314880;
      46287: inst = 32'd268468224;
      46288: inst = 32'd201346056;
      46289: inst = 32'd203483685;
      46290: inst = 32'd471859200;
      46291: inst = 32'd136314880;
      46292: inst = 32'd268468224;
      46293: inst = 32'd201346057;
      46294: inst = 32'd203483685;
      46295: inst = 32'd471859200;
      46296: inst = 32'd136314880;
      46297: inst = 32'd268468224;
      46298: inst = 32'd201346058;
      46299: inst = 32'd203483685;
      46300: inst = 32'd471859200;
      46301: inst = 32'd136314880;
      46302: inst = 32'd268468224;
      46303: inst = 32'd201346059;
      46304: inst = 32'd203483685;
      46305: inst = 32'd471859200;
      46306: inst = 32'd136314880;
      46307: inst = 32'd268468224;
      46308: inst = 32'd201346060;
      46309: inst = 32'd203483685;
      46310: inst = 32'd471859200;
      46311: inst = 32'd136314880;
      46312: inst = 32'd268468224;
      46313: inst = 32'd201346061;
      46314: inst = 32'd203483685;
      46315: inst = 32'd471859200;
      46316: inst = 32'd136314880;
      46317: inst = 32'd268468224;
      46318: inst = 32'd201346062;
      46319: inst = 32'd203483685;
      46320: inst = 32'd471859200;
      46321: inst = 32'd136314880;
      46322: inst = 32'd268468224;
      46323: inst = 32'd201346063;
      46324: inst = 32'd203483685;
      46325: inst = 32'd471859200;
      46326: inst = 32'd136314880;
      46327: inst = 32'd268468224;
      46328: inst = 32'd201346064;
      46329: inst = 32'd203483685;
      46330: inst = 32'd471859200;
      46331: inst = 32'd136314880;
      46332: inst = 32'd268468224;
      46333: inst = 32'd201346065;
      46334: inst = 32'd203483685;
      46335: inst = 32'd471859200;
      46336: inst = 32'd136314880;
      46337: inst = 32'd268468224;
      46338: inst = 32'd201346066;
      46339: inst = 32'd203483685;
      46340: inst = 32'd471859200;
      46341: inst = 32'd136314880;
      46342: inst = 32'd268468224;
      46343: inst = 32'd201346067;
      46344: inst = 32'd203483685;
      46345: inst = 32'd471859200;
      46346: inst = 32'd136314880;
      46347: inst = 32'd268468224;
      46348: inst = 32'd201346068;
      46349: inst = 32'd203483685;
      46350: inst = 32'd471859200;
      46351: inst = 32'd136314880;
      46352: inst = 32'd268468224;
      46353: inst = 32'd201346069;
      46354: inst = 32'd203483685;
      46355: inst = 32'd471859200;
      46356: inst = 32'd136314880;
      46357: inst = 32'd268468224;
      46358: inst = 32'd201346070;
      46359: inst = 32'd203423744;
      46360: inst = 32'd471859200;
      46361: inst = 32'd136314880;
      46362: inst = 32'd268468224;
      46363: inst = 32'd201346071;
      46364: inst = 32'd203423744;
      46365: inst = 32'd471859200;
      46366: inst = 32'd136314880;
      46367: inst = 32'd268468224;
      46368: inst = 32'd201346072;
      46369: inst = 32'd203423744;
      46370: inst = 32'd471859200;
      46371: inst = 32'd136314880;
      46372: inst = 32'd268468224;
      46373: inst = 32'd201346073;
      46374: inst = 32'd203423744;
      46375: inst = 32'd471859200;
      46376: inst = 32'd136314880;
      46377: inst = 32'd268468224;
      46378: inst = 32'd201346074;
      46379: inst = 32'd203423744;
      46380: inst = 32'd471859200;
      46381: inst = 32'd136314880;
      46382: inst = 32'd268468224;
      46383: inst = 32'd201346075;
      46384: inst = 32'd203423744;
      46385: inst = 32'd471859200;
      46386: inst = 32'd136314880;
      46387: inst = 32'd268468224;
      46388: inst = 32'd201346076;
      46389: inst = 32'd203423744;
      46390: inst = 32'd471859200;
      46391: inst = 32'd136314880;
      46392: inst = 32'd268468224;
      46393: inst = 32'd201346077;
      46394: inst = 32'd203423744;
      46395: inst = 32'd471859200;
      46396: inst = 32'd136314880;
      46397: inst = 32'd268468224;
      46398: inst = 32'd201346078;
      46399: inst = 32'd203483685;
      46400: inst = 32'd471859200;
      46401: inst = 32'd136314880;
      46402: inst = 32'd268468224;
      46403: inst = 32'd201346079;
      46404: inst = 32'd203483685;
      46405: inst = 32'd471859200;
      46406: inst = 32'd136314880;
      46407: inst = 32'd268468224;
      46408: inst = 32'd201346080;
      46409: inst = 32'd203483685;
      46410: inst = 32'd471859200;
      46411: inst = 32'd136314880;
      46412: inst = 32'd268468224;
      46413: inst = 32'd201346081;
      46414: inst = 32'd203483685;
      46415: inst = 32'd471859200;
      46416: inst = 32'd136314880;
      46417: inst = 32'd268468224;
      46418: inst = 32'd201346082;
      46419: inst = 32'd203483685;
      46420: inst = 32'd471859200;
      46421: inst = 32'd136314880;
      46422: inst = 32'd268468224;
      46423: inst = 32'd201346083;
      46424: inst = 32'd203483685;
      46425: inst = 32'd471859200;
      46426: inst = 32'd136314880;
      46427: inst = 32'd268468224;
      46428: inst = 32'd201346084;
      46429: inst = 32'd203483685;
      46430: inst = 32'd471859200;
      46431: inst = 32'd136314880;
      46432: inst = 32'd268468224;
      46433: inst = 32'd201346085;
      46434: inst = 32'd203483685;
      46435: inst = 32'd471859200;
      46436: inst = 32'd136314880;
      46437: inst = 32'd268468224;
      46438: inst = 32'd201346086;
      46439: inst = 32'd203483685;
      46440: inst = 32'd471859200;
      46441: inst = 32'd136314880;
      46442: inst = 32'd268468224;
      46443: inst = 32'd201346087;
      46444: inst = 32'd203483685;
      46445: inst = 32'd471859200;
      46446: inst = 32'd136314880;
      46447: inst = 32'd268468224;
      46448: inst = 32'd201346088;
      46449: inst = 32'd203483685;
      46450: inst = 32'd471859200;
      46451: inst = 32'd136314880;
      46452: inst = 32'd268468224;
      46453: inst = 32'd201346089;
      46454: inst = 32'd203483685;
      46455: inst = 32'd471859200;
      46456: inst = 32'd136314880;
      46457: inst = 32'd268468224;
      46458: inst = 32'd201346090;
      46459: inst = 32'd203483685;
      46460: inst = 32'd471859200;
      46461: inst = 32'd136314880;
      46462: inst = 32'd268468224;
      46463: inst = 32'd201346091;
      46464: inst = 32'd203423744;
      46465: inst = 32'd471859200;
      46466: inst = 32'd136314880;
      46467: inst = 32'd268468224;
      46468: inst = 32'd201346092;
      46469: inst = 32'd203483685;
      46470: inst = 32'd471859200;
      46471: inst = 32'd136314880;
      46472: inst = 32'd268468224;
      46473: inst = 32'd201346093;
      46474: inst = 32'd203483685;
      46475: inst = 32'd471859200;
      46476: inst = 32'd136314880;
      46477: inst = 32'd268468224;
      46478: inst = 32'd201346094;
      46479: inst = 32'd203483685;
      46480: inst = 32'd471859200;
      46481: inst = 32'd136314880;
      46482: inst = 32'd268468224;
      46483: inst = 32'd201346095;
      46484: inst = 32'd203483685;
      46485: inst = 32'd471859200;
      46486: inst = 32'd136314880;
      46487: inst = 32'd268468224;
      46488: inst = 32'd201346096;
      46489: inst = 32'd203483685;
      46490: inst = 32'd471859200;
      46491: inst = 32'd136314880;
      46492: inst = 32'd268468224;
      46493: inst = 32'd201346097;
      46494: inst = 32'd203483685;
      46495: inst = 32'd471859200;
      46496: inst = 32'd136314880;
      46497: inst = 32'd268468224;
      46498: inst = 32'd201346098;
      46499: inst = 32'd203483685;
      46500: inst = 32'd471859200;
      46501: inst = 32'd136314880;
      46502: inst = 32'd268468224;
      46503: inst = 32'd201346099;
      46504: inst = 32'd203483685;
      46505: inst = 32'd471859200;
      46506: inst = 32'd136314880;
      46507: inst = 32'd268468224;
      46508: inst = 32'd201346100;
      46509: inst = 32'd203483685;
      46510: inst = 32'd471859200;
      46511: inst = 32'd136314880;
      46512: inst = 32'd268468224;
      46513: inst = 32'd201346101;
      46514: inst = 32'd203483685;
      46515: inst = 32'd471859200;
      46516: inst = 32'd136314880;
      46517: inst = 32'd268468224;
      46518: inst = 32'd201346102;
      46519: inst = 32'd203423744;
      46520: inst = 32'd471859200;
      46521: inst = 32'd136314880;
      46522: inst = 32'd268468224;
      46523: inst = 32'd201346103;
      46524: inst = 32'd203423744;
      46525: inst = 32'd471859200;
      46526: inst = 32'd136314880;
      46527: inst = 32'd268468224;
      46528: inst = 32'd201346104;
      46529: inst = 32'd203423744;
      46530: inst = 32'd471859200;
      46531: inst = 32'd136314880;
      46532: inst = 32'd268468224;
      46533: inst = 32'd201346105;
      46534: inst = 32'd203423744;
      46535: inst = 32'd471859200;
      46536: inst = 32'd136314880;
      46537: inst = 32'd268468224;
      46538: inst = 32'd201346106;
      46539: inst = 32'd203423744;
      46540: inst = 32'd471859200;
      46541: inst = 32'd136314880;
      46542: inst = 32'd268468224;
      46543: inst = 32'd201346107;
      46544: inst = 32'd203423744;
      46545: inst = 32'd471859200;
      46546: inst = 32'd136314880;
      46547: inst = 32'd268468224;
      46548: inst = 32'd201346108;
      46549: inst = 32'd203423744;
      46550: inst = 32'd471859200;
      46551: inst = 32'd136314880;
      46552: inst = 32'd268468224;
      46553: inst = 32'd201346109;
      46554: inst = 32'd203423744;
      46555: inst = 32'd471859200;
      46556: inst = 32'd136314880;
      46557: inst = 32'd268468224;
      46558: inst = 32'd201346110;
      46559: inst = 32'd203423744;
      46560: inst = 32'd471859200;
      46561: inst = 32'd136314880;
      46562: inst = 32'd268468224;
      46563: inst = 32'd201346111;
      46564: inst = 32'd203423744;
      46565: inst = 32'd471859200;
      46566: inst = 32'd136314880;
      46567: inst = 32'd268468224;
      46568: inst = 32'd201346112;
      46569: inst = 32'd203423744;
      46570: inst = 32'd471859200;
      46571: inst = 32'd136314880;
      46572: inst = 32'd268468224;
      46573: inst = 32'd201346113;
      46574: inst = 32'd203423744;
      46575: inst = 32'd471859200;
      46576: inst = 32'd136314880;
      46577: inst = 32'd268468224;
      46578: inst = 32'd201346114;
      46579: inst = 32'd203423744;
      46580: inst = 32'd471859200;
      46581: inst = 32'd136314880;
      46582: inst = 32'd268468224;
      46583: inst = 32'd201346115;
      46584: inst = 32'd203423744;
      46585: inst = 32'd471859200;
      46586: inst = 32'd136314880;
      46587: inst = 32'd268468224;
      46588: inst = 32'd201346116;
      46589: inst = 32'd203423744;
      46590: inst = 32'd471859200;
      46591: inst = 32'd136314880;
      46592: inst = 32'd268468224;
      46593: inst = 32'd201346117;
      46594: inst = 32'd203423744;
      46595: inst = 32'd471859200;
      46596: inst = 32'd136314880;
      46597: inst = 32'd268468224;
      46598: inst = 32'd201346118;
      46599: inst = 32'd203423744;
      46600: inst = 32'd471859200;
      46601: inst = 32'd136314880;
      46602: inst = 32'd268468224;
      46603: inst = 32'd201346119;
      46604: inst = 32'd203423744;
      46605: inst = 32'd471859200;
      46606: inst = 32'd136314880;
      46607: inst = 32'd268468224;
      46608: inst = 32'd201346120;
      46609: inst = 32'd203423744;
      46610: inst = 32'd471859200;
      46611: inst = 32'd136314880;
      46612: inst = 32'd268468224;
      46613: inst = 32'd201346121;
      46614: inst = 32'd203423744;
      46615: inst = 32'd471859200;
      46616: inst = 32'd136314880;
      46617: inst = 32'd268468224;
      46618: inst = 32'd201346122;
      46619: inst = 32'd203423744;
      46620: inst = 32'd471859200;
      46621: inst = 32'd136314880;
      46622: inst = 32'd268468224;
      46623: inst = 32'd201346123;
      46624: inst = 32'd203423744;
      46625: inst = 32'd471859200;
      46626: inst = 32'd136314880;
      46627: inst = 32'd268468224;
      46628: inst = 32'd201346124;
      46629: inst = 32'd203423744;
      46630: inst = 32'd471859200;
      46631: inst = 32'd136314880;
      46632: inst = 32'd268468224;
      46633: inst = 32'd201346125;
      46634: inst = 32'd203483685;
      46635: inst = 32'd471859200;
      46636: inst = 32'd136314880;
      46637: inst = 32'd268468224;
      46638: inst = 32'd201346126;
      46639: inst = 32'd203483685;
      46640: inst = 32'd471859200;
      46641: inst = 32'd136314880;
      46642: inst = 32'd268468224;
      46643: inst = 32'd201346127;
      46644: inst = 32'd203483685;
      46645: inst = 32'd471859200;
      46646: inst = 32'd136314880;
      46647: inst = 32'd268468224;
      46648: inst = 32'd201346128;
      46649: inst = 32'd203483685;
      46650: inst = 32'd471859200;
      46651: inst = 32'd136314880;
      46652: inst = 32'd268468224;
      46653: inst = 32'd201346129;
      46654: inst = 32'd203483685;
      46655: inst = 32'd471859200;
      46656: inst = 32'd136314880;
      46657: inst = 32'd268468224;
      46658: inst = 32'd201346130;
      46659: inst = 32'd203483685;
      46660: inst = 32'd471859200;
      46661: inst = 32'd136314880;
      46662: inst = 32'd268468224;
      46663: inst = 32'd201346131;
      46664: inst = 32'd203483685;
      46665: inst = 32'd471859200;
      46666: inst = 32'd136314880;
      46667: inst = 32'd268468224;
      46668: inst = 32'd201346132;
      46669: inst = 32'd203483685;
      46670: inst = 32'd471859200;
      46671: inst = 32'd136314880;
      46672: inst = 32'd268468224;
      46673: inst = 32'd201346133;
      46674: inst = 32'd203483685;
      46675: inst = 32'd471859200;
      46676: inst = 32'd136314880;
      46677: inst = 32'd268468224;
      46678: inst = 32'd201346134;
      46679: inst = 32'd203483685;
      46680: inst = 32'd471859200;
      46681: inst = 32'd136314880;
      46682: inst = 32'd268468224;
      46683: inst = 32'd201346135;
      46684: inst = 32'd203483685;
      46685: inst = 32'd471859200;
      46686: inst = 32'd136314880;
      46687: inst = 32'd268468224;
      46688: inst = 32'd201346136;
      46689: inst = 32'd203483685;
      46690: inst = 32'd471859200;
      46691: inst = 32'd136314880;
      46692: inst = 32'd268468224;
      46693: inst = 32'd201346137;
      46694: inst = 32'd203483685;
      46695: inst = 32'd471859200;
      46696: inst = 32'd136314880;
      46697: inst = 32'd268468224;
      46698: inst = 32'd201346138;
      46699: inst = 32'd203483685;
      46700: inst = 32'd471859200;
      46701: inst = 32'd136314880;
      46702: inst = 32'd268468224;
      46703: inst = 32'd201346139;
      46704: inst = 32'd203483685;
      46705: inst = 32'd471859200;
      46706: inst = 32'd136314880;
      46707: inst = 32'd268468224;
      46708: inst = 32'd201346140;
      46709: inst = 32'd203483685;
      46710: inst = 32'd471859200;
      46711: inst = 32'd136314880;
      46712: inst = 32'd268468224;
      46713: inst = 32'd201346141;
      46714: inst = 32'd203483685;
      46715: inst = 32'd471859200;
      46716: inst = 32'd136314880;
      46717: inst = 32'd268468224;
      46718: inst = 32'd201346142;
      46719: inst = 32'd203483685;
      46720: inst = 32'd471859200;
      46721: inst = 32'd136314880;
      46722: inst = 32'd268468224;
      46723: inst = 32'd201346143;
      46724: inst = 32'd203483685;
      46725: inst = 32'd471859200;
      46726: inst = 32'd136314880;
      46727: inst = 32'd268468224;
      46728: inst = 32'd201346144;
      46729: inst = 32'd203483685;
      46730: inst = 32'd471859200;
      46731: inst = 32'd136314880;
      46732: inst = 32'd268468224;
      46733: inst = 32'd201346145;
      46734: inst = 32'd203483685;
      46735: inst = 32'd471859200;
      46736: inst = 32'd136314880;
      46737: inst = 32'd268468224;
      46738: inst = 32'd201346146;
      46739: inst = 32'd203483685;
      46740: inst = 32'd471859200;
      46741: inst = 32'd136314880;
      46742: inst = 32'd268468224;
      46743: inst = 32'd201346147;
      46744: inst = 32'd203483685;
      46745: inst = 32'd471859200;
      46746: inst = 32'd136314880;
      46747: inst = 32'd268468224;
      46748: inst = 32'd201346148;
      46749: inst = 32'd203483685;
      46750: inst = 32'd471859200;
      46751: inst = 32'd136314880;
      46752: inst = 32'd268468224;
      46753: inst = 32'd201346149;
      46754: inst = 32'd203483685;
      46755: inst = 32'd471859200;
      46756: inst = 32'd136314880;
      46757: inst = 32'd268468224;
      46758: inst = 32'd201346150;
      46759: inst = 32'd203483685;
      46760: inst = 32'd471859200;
      46761: inst = 32'd136314880;
      46762: inst = 32'd268468224;
      46763: inst = 32'd201346151;
      46764: inst = 32'd203483685;
      46765: inst = 32'd471859200;
      46766: inst = 32'd136314880;
      46767: inst = 32'd268468224;
      46768: inst = 32'd201346152;
      46769: inst = 32'd203483685;
      46770: inst = 32'd471859200;
      46771: inst = 32'd136314880;
      46772: inst = 32'd268468224;
      46773: inst = 32'd201346153;
      46774: inst = 32'd203483685;
      46775: inst = 32'd471859200;
      46776: inst = 32'd136314880;
      46777: inst = 32'd268468224;
      46778: inst = 32'd201346154;
      46779: inst = 32'd203483685;
      46780: inst = 32'd471859200;
      46781: inst = 32'd136314880;
      46782: inst = 32'd268468224;
      46783: inst = 32'd201346155;
      46784: inst = 32'd203483685;
      46785: inst = 32'd471859200;
      46786: inst = 32'd136314880;
      46787: inst = 32'd268468224;
      46788: inst = 32'd201346156;
      46789: inst = 32'd203483685;
      46790: inst = 32'd471859200;
      46791: inst = 32'd136314880;
      46792: inst = 32'd268468224;
      46793: inst = 32'd201346157;
      46794: inst = 32'd203483685;
      46795: inst = 32'd471859200;
      46796: inst = 32'd136314880;
      46797: inst = 32'd268468224;
      46798: inst = 32'd201346158;
      46799: inst = 32'd203483685;
      46800: inst = 32'd471859200;
      46801: inst = 32'd136314880;
      46802: inst = 32'd268468224;
      46803: inst = 32'd201346159;
      46804: inst = 32'd203483685;
      46805: inst = 32'd471859200;
      46806: inst = 32'd136314880;
      46807: inst = 32'd268468224;
      46808: inst = 32'd201346160;
      46809: inst = 32'd203483685;
      46810: inst = 32'd471859200;
      46811: inst = 32'd136314880;
      46812: inst = 32'd268468224;
      46813: inst = 32'd201346161;
      46814: inst = 32'd203483685;
      46815: inst = 32'd471859200;
      46816: inst = 32'd136314880;
      46817: inst = 32'd268468224;
      46818: inst = 32'd201346162;
      46819: inst = 32'd203483685;
      46820: inst = 32'd471859200;
      46821: inst = 32'd136314880;
      46822: inst = 32'd268468224;
      46823: inst = 32'd201346163;
      46824: inst = 32'd203483685;
      46825: inst = 32'd471859200;
      46826: inst = 32'd136314880;
      46827: inst = 32'd268468224;
      46828: inst = 32'd201346164;
      46829: inst = 32'd203483685;
      46830: inst = 32'd471859200;
      46831: inst = 32'd136314880;
      46832: inst = 32'd268468224;
      46833: inst = 32'd201346165;
      46834: inst = 32'd203483685;
      46835: inst = 32'd471859200;
      46836: inst = 32'd136314880;
      46837: inst = 32'd268468224;
      46838: inst = 32'd201346166;
      46839: inst = 32'd203483685;
      46840: inst = 32'd471859200;
      46841: inst = 32'd136314880;
      46842: inst = 32'd268468224;
      46843: inst = 32'd201346167;
      46844: inst = 32'd203423744;
      46845: inst = 32'd471859200;
      46846: inst = 32'd136314880;
      46847: inst = 32'd268468224;
      46848: inst = 32'd201346168;
      46849: inst = 32'd203423744;
      46850: inst = 32'd471859200;
      46851: inst = 32'd136314880;
      46852: inst = 32'd268468224;
      46853: inst = 32'd201346169;
      46854: inst = 32'd203423744;
      46855: inst = 32'd471859200;
      46856: inst = 32'd136314880;
      46857: inst = 32'd268468224;
      46858: inst = 32'd201346170;
      46859: inst = 32'd203423744;
      46860: inst = 32'd471859200;
      46861: inst = 32'd136314880;
      46862: inst = 32'd268468224;
      46863: inst = 32'd201346171;
      46864: inst = 32'd203423744;
      46865: inst = 32'd471859200;
      46866: inst = 32'd136314880;
      46867: inst = 32'd268468224;
      46868: inst = 32'd201346172;
      46869: inst = 32'd203423744;
      46870: inst = 32'd471859200;
      46871: inst = 32'd136314880;
      46872: inst = 32'd268468224;
      46873: inst = 32'd201346173;
      46874: inst = 32'd203423744;
      46875: inst = 32'd471859200;
      46876: inst = 32'd136314880;
      46877: inst = 32'd268468224;
      46878: inst = 32'd201346174;
      46879: inst = 32'd203483685;
      46880: inst = 32'd471859200;
      46881: inst = 32'd136314880;
      46882: inst = 32'd268468224;
      46883: inst = 32'd201346175;
      46884: inst = 32'd203483685;
      46885: inst = 32'd471859200;
      46886: inst = 32'd136314880;
      46887: inst = 32'd268468224;
      46888: inst = 32'd201346176;
      46889: inst = 32'd203483685;
      46890: inst = 32'd471859200;
      46891: inst = 32'd136314880;
      46892: inst = 32'd268468224;
      46893: inst = 32'd201346177;
      46894: inst = 32'd203483685;
      46895: inst = 32'd471859200;
      46896: inst = 32'd136314880;
      46897: inst = 32'd268468224;
      46898: inst = 32'd201346178;
      46899: inst = 32'd203483685;
      46900: inst = 32'd471859200;
      46901: inst = 32'd136314880;
      46902: inst = 32'd268468224;
      46903: inst = 32'd201346179;
      46904: inst = 32'd203483685;
      46905: inst = 32'd471859200;
      46906: inst = 32'd136314880;
      46907: inst = 32'd268468224;
      46908: inst = 32'd201346180;
      46909: inst = 32'd203483685;
      46910: inst = 32'd471859200;
      46911: inst = 32'd136314880;
      46912: inst = 32'd268468224;
      46913: inst = 32'd201346181;
      46914: inst = 32'd203483685;
      46915: inst = 32'd471859200;
      46916: inst = 32'd136314880;
      46917: inst = 32'd268468224;
      46918: inst = 32'd201346182;
      46919: inst = 32'd203483685;
      46920: inst = 32'd471859200;
      46921: inst = 32'd136314880;
      46922: inst = 32'd268468224;
      46923: inst = 32'd201346183;
      46924: inst = 32'd203483685;
      46925: inst = 32'd471859200;
      46926: inst = 32'd136314880;
      46927: inst = 32'd268468224;
      46928: inst = 32'd201346184;
      46929: inst = 32'd203483685;
      46930: inst = 32'd471859200;
      46931: inst = 32'd136314880;
      46932: inst = 32'd268468224;
      46933: inst = 32'd201346185;
      46934: inst = 32'd203483685;
      46935: inst = 32'd471859200;
      46936: inst = 32'd136314880;
      46937: inst = 32'd268468224;
      46938: inst = 32'd201346186;
      46939: inst = 32'd203423744;
      46940: inst = 32'd471859200;
      46941: inst = 32'd136314880;
      46942: inst = 32'd268468224;
      46943: inst = 32'd201346187;
      46944: inst = 32'd203483685;
      46945: inst = 32'd471859200;
      46946: inst = 32'd136314880;
      46947: inst = 32'd268468224;
      46948: inst = 32'd201346188;
      46949: inst = 32'd203483685;
      46950: inst = 32'd471859200;
      46951: inst = 32'd136314880;
      46952: inst = 32'd268468224;
      46953: inst = 32'd201346189;
      46954: inst = 32'd203483685;
      46955: inst = 32'd471859200;
      46956: inst = 32'd136314880;
      46957: inst = 32'd268468224;
      46958: inst = 32'd201346190;
      46959: inst = 32'd203483685;
      46960: inst = 32'd471859200;
      46961: inst = 32'd136314880;
      46962: inst = 32'd268468224;
      46963: inst = 32'd201346191;
      46964: inst = 32'd203483685;
      46965: inst = 32'd471859200;
      46966: inst = 32'd136314880;
      46967: inst = 32'd268468224;
      46968: inst = 32'd201346192;
      46969: inst = 32'd203483685;
      46970: inst = 32'd471859200;
      46971: inst = 32'd136314880;
      46972: inst = 32'd268468224;
      46973: inst = 32'd201346193;
      46974: inst = 32'd203483685;
      46975: inst = 32'd471859200;
      46976: inst = 32'd136314880;
      46977: inst = 32'd268468224;
      46978: inst = 32'd201346194;
      46979: inst = 32'd203483685;
      46980: inst = 32'd471859200;
      46981: inst = 32'd136314880;
      46982: inst = 32'd268468224;
      46983: inst = 32'd201346195;
      46984: inst = 32'd203483685;
      46985: inst = 32'd471859200;
      46986: inst = 32'd136314880;
      46987: inst = 32'd268468224;
      46988: inst = 32'd201346196;
      46989: inst = 32'd203483685;
      46990: inst = 32'd471859200;
      46991: inst = 32'd136314880;
      46992: inst = 32'd268468224;
      46993: inst = 32'd201346197;
      46994: inst = 32'd203483685;
      46995: inst = 32'd471859200;
      46996: inst = 32'd136314880;
      46997: inst = 32'd268468224;
      46998: inst = 32'd201346198;
      46999: inst = 32'd203423744;
      47000: inst = 32'd471859200;
      47001: inst = 32'd136314880;
      47002: inst = 32'd268468224;
      47003: inst = 32'd201346199;
      47004: inst = 32'd203423744;
      47005: inst = 32'd471859200;
      47006: inst = 32'd136314880;
      47007: inst = 32'd268468224;
      47008: inst = 32'd201346200;
      47009: inst = 32'd203423744;
      47010: inst = 32'd471859200;
      47011: inst = 32'd136314880;
      47012: inst = 32'd268468224;
      47013: inst = 32'd201346201;
      47014: inst = 32'd203423744;
      47015: inst = 32'd471859200;
      47016: inst = 32'd136314880;
      47017: inst = 32'd268468224;
      47018: inst = 32'd201346202;
      47019: inst = 32'd203423744;
      47020: inst = 32'd471859200;
      47021: inst = 32'd136314880;
      47022: inst = 32'd268468224;
      47023: inst = 32'd201346203;
      47024: inst = 32'd203423744;
      47025: inst = 32'd471859200;
      47026: inst = 32'd136314880;
      47027: inst = 32'd268468224;
      47028: inst = 32'd201346204;
      47029: inst = 32'd203423744;
      47030: inst = 32'd471859200;
      47031: inst = 32'd136314880;
      47032: inst = 32'd268468224;
      47033: inst = 32'd201346205;
      47034: inst = 32'd203423744;
      47035: inst = 32'd471859200;
      47036: inst = 32'd136314880;
      47037: inst = 32'd268468224;
      47038: inst = 32'd201346206;
      47039: inst = 32'd203423744;
      47040: inst = 32'd471859200;
      47041: inst = 32'd136314880;
      47042: inst = 32'd268468224;
      47043: inst = 32'd201346207;
      47044: inst = 32'd203423744;
      47045: inst = 32'd471859200;
      47046: inst = 32'd136314880;
      47047: inst = 32'd268468224;
      47048: inst = 32'd201346208;
      47049: inst = 32'd203423744;
      47050: inst = 32'd471859200;
      47051: inst = 32'd136314880;
      47052: inst = 32'd268468224;
      47053: inst = 32'd201346209;
      47054: inst = 32'd203423744;
      47055: inst = 32'd471859200;
      47056: inst = 32'd136314880;
      47057: inst = 32'd268468224;
      47058: inst = 32'd201346210;
      47059: inst = 32'd203423744;
      47060: inst = 32'd471859200;
      47061: inst = 32'd136314880;
      47062: inst = 32'd268468224;
      47063: inst = 32'd201346211;
      47064: inst = 32'd203423744;
      47065: inst = 32'd471859200;
      47066: inst = 32'd136314880;
      47067: inst = 32'd268468224;
      47068: inst = 32'd201346212;
      47069: inst = 32'd203423744;
      47070: inst = 32'd471859200;
      47071: inst = 32'd136314880;
      47072: inst = 32'd268468224;
      47073: inst = 32'd201346213;
      47074: inst = 32'd203423744;
      47075: inst = 32'd471859200;
      47076: inst = 32'd136314880;
      47077: inst = 32'd268468224;
      47078: inst = 32'd201346214;
      47079: inst = 32'd203423744;
      47080: inst = 32'd471859200;
      47081: inst = 32'd136314880;
      47082: inst = 32'd268468224;
      47083: inst = 32'd201346215;
      47084: inst = 32'd203423744;
      47085: inst = 32'd471859200;
      47086: inst = 32'd136314880;
      47087: inst = 32'd268468224;
      47088: inst = 32'd201346216;
      47089: inst = 32'd203423744;
      47090: inst = 32'd471859200;
      47091: inst = 32'd136314880;
      47092: inst = 32'd268468224;
      47093: inst = 32'd201346217;
      47094: inst = 32'd203423744;
      47095: inst = 32'd471859200;
      47096: inst = 32'd136314880;
      47097: inst = 32'd268468224;
      47098: inst = 32'd201346218;
      47099: inst = 32'd203423744;
      47100: inst = 32'd471859200;
      47101: inst = 32'd136314880;
      47102: inst = 32'd268468224;
      47103: inst = 32'd201346219;
      47104: inst = 32'd203423744;
      47105: inst = 32'd471859200;
      47106: inst = 32'd136314880;
      47107: inst = 32'd268468224;
      47108: inst = 32'd201346220;
      47109: inst = 32'd203423744;
      47110: inst = 32'd471859200;
      47111: inst = 32'd136314880;
      47112: inst = 32'd268468224;
      47113: inst = 32'd201346221;
      47114: inst = 32'd203483685;
      47115: inst = 32'd471859200;
      47116: inst = 32'd136314880;
      47117: inst = 32'd268468224;
      47118: inst = 32'd201346222;
      47119: inst = 32'd203483685;
      47120: inst = 32'd471859200;
      47121: inst = 32'd136314880;
      47122: inst = 32'd268468224;
      47123: inst = 32'd201346223;
      47124: inst = 32'd203483685;
      47125: inst = 32'd471859200;
      47126: inst = 32'd136314880;
      47127: inst = 32'd268468224;
      47128: inst = 32'd201346224;
      47129: inst = 32'd203483685;
      47130: inst = 32'd471859200;
      47131: inst = 32'd136314880;
      47132: inst = 32'd268468224;
      47133: inst = 32'd201346225;
      47134: inst = 32'd203483685;
      47135: inst = 32'd471859200;
      47136: inst = 32'd136314880;
      47137: inst = 32'd268468224;
      47138: inst = 32'd201346226;
      47139: inst = 32'd203483685;
      47140: inst = 32'd471859200;
      47141: inst = 32'd136314880;
      47142: inst = 32'd268468224;
      47143: inst = 32'd201346227;
      47144: inst = 32'd203483685;
      47145: inst = 32'd471859200;
      47146: inst = 32'd136314880;
      47147: inst = 32'd268468224;
      47148: inst = 32'd201346228;
      47149: inst = 32'd203483685;
      47150: inst = 32'd471859200;
      47151: inst = 32'd136314880;
      47152: inst = 32'd268468224;
      47153: inst = 32'd201346229;
      47154: inst = 32'd203483685;
      47155: inst = 32'd471859200;
      47156: inst = 32'd136314880;
      47157: inst = 32'd268468224;
      47158: inst = 32'd201346230;
      47159: inst = 32'd203483685;
      47160: inst = 32'd471859200;
      47161: inst = 32'd136314880;
      47162: inst = 32'd268468224;
      47163: inst = 32'd201346231;
      47164: inst = 32'd203483685;
      47165: inst = 32'd471859200;
      47166: inst = 32'd136314880;
      47167: inst = 32'd268468224;
      47168: inst = 32'd201346232;
      47169: inst = 32'd203483685;
      47170: inst = 32'd471859200;
      47171: inst = 32'd136314880;
      47172: inst = 32'd268468224;
      47173: inst = 32'd201346233;
      47174: inst = 32'd203423744;
      47175: inst = 32'd471859200;
      47176: inst = 32'd136314880;
      47177: inst = 32'd268468224;
      47178: inst = 32'd201346234;
      47179: inst = 32'd203483685;
      47180: inst = 32'd471859200;
      47181: inst = 32'd136314880;
      47182: inst = 32'd268468224;
      47183: inst = 32'd201346235;
      47184: inst = 32'd203483685;
      47185: inst = 32'd471859200;
      47186: inst = 32'd136314880;
      47187: inst = 32'd268468224;
      47188: inst = 32'd201346236;
      47189: inst = 32'd203483685;
      47190: inst = 32'd471859200;
      47191: inst = 32'd136314880;
      47192: inst = 32'd268468224;
      47193: inst = 32'd201346237;
      47194: inst = 32'd203483685;
      47195: inst = 32'd471859200;
      47196: inst = 32'd136314880;
      47197: inst = 32'd268468224;
      47198: inst = 32'd201346238;
      47199: inst = 32'd203483685;
      47200: inst = 32'd471859200;
      47201: inst = 32'd136314880;
      47202: inst = 32'd268468224;
      47203: inst = 32'd201346239;
      47204: inst = 32'd203483685;
      47205: inst = 32'd471859200;
      47206: inst = 32'd136314880;
      47207: inst = 32'd268468224;
      47208: inst = 32'd201346240;
      47209: inst = 32'd203483685;
      47210: inst = 32'd471859200;
      47211: inst = 32'd136314880;
      47212: inst = 32'd268468224;
      47213: inst = 32'd201346241;
      47214: inst = 32'd203483685;
      47215: inst = 32'd471859200;
      47216: inst = 32'd136314880;
      47217: inst = 32'd268468224;
      47218: inst = 32'd201346242;
      47219: inst = 32'd203483685;
      47220: inst = 32'd471859200;
      47221: inst = 32'd136314880;
      47222: inst = 32'd268468224;
      47223: inst = 32'd201346243;
      47224: inst = 32'd203483685;
      47225: inst = 32'd471859200;
      47226: inst = 32'd136314880;
      47227: inst = 32'd268468224;
      47228: inst = 32'd201346244;
      47229: inst = 32'd203483685;
      47230: inst = 32'd471859200;
      47231: inst = 32'd136314880;
      47232: inst = 32'd268468224;
      47233: inst = 32'd201346245;
      47234: inst = 32'd203483685;
      47235: inst = 32'd471859200;
      47236: inst = 32'd136314880;
      47237: inst = 32'd268468224;
      47238: inst = 32'd201346246;
      47239: inst = 32'd203483685;
      47240: inst = 32'd471859200;
      47241: inst = 32'd136314880;
      47242: inst = 32'd268468224;
      47243: inst = 32'd201346247;
      47244: inst = 32'd203483685;
      47245: inst = 32'd471859200;
      47246: inst = 32'd136314880;
      47247: inst = 32'd268468224;
      47248: inst = 32'd201346248;
      47249: inst = 32'd203483685;
      47250: inst = 32'd471859200;
      47251: inst = 32'd136314880;
      47252: inst = 32'd268468224;
      47253: inst = 32'd201346249;
      47254: inst = 32'd203483685;
      47255: inst = 32'd471859200;
      47256: inst = 32'd136314880;
      47257: inst = 32'd268468224;
      47258: inst = 32'd201346250;
      47259: inst = 32'd203483685;
      47260: inst = 32'd471859200;
      47261: inst = 32'd136314880;
      47262: inst = 32'd268468224;
      47263: inst = 32'd201346251;
      47264: inst = 32'd203483685;
      47265: inst = 32'd471859200;
      47266: inst = 32'd136314880;
      47267: inst = 32'd268468224;
      47268: inst = 32'd201346252;
      47269: inst = 32'd203483685;
      47270: inst = 32'd471859200;
      47271: inst = 32'd136314880;
      47272: inst = 32'd268468224;
      47273: inst = 32'd201346253;
      47274: inst = 32'd203483685;
      47275: inst = 32'd471859200;
      47276: inst = 32'd136314880;
      47277: inst = 32'd268468224;
      47278: inst = 32'd201346254;
      47279: inst = 32'd203483685;
      47280: inst = 32'd471859200;
      47281: inst = 32'd136314880;
      47282: inst = 32'd268468224;
      47283: inst = 32'd201346255;
      47284: inst = 32'd203483685;
      47285: inst = 32'd471859200;
      47286: inst = 32'd136314880;
      47287: inst = 32'd268468224;
      47288: inst = 32'd201346256;
      47289: inst = 32'd203483685;
      47290: inst = 32'd471859200;
      47291: inst = 32'd136314880;
      47292: inst = 32'd268468224;
      47293: inst = 32'd201346257;
      47294: inst = 32'd203483685;
      47295: inst = 32'd471859200;
      47296: inst = 32'd136314880;
      47297: inst = 32'd268468224;
      47298: inst = 32'd201346258;
      47299: inst = 32'd203483685;
      47300: inst = 32'd471859200;
      47301: inst = 32'd136314880;
      47302: inst = 32'd268468224;
      47303: inst = 32'd201346259;
      47304: inst = 32'd203483685;
      47305: inst = 32'd471859200;
      47306: inst = 32'd136314880;
      47307: inst = 32'd268468224;
      47308: inst = 32'd201346260;
      47309: inst = 32'd203483685;
      47310: inst = 32'd471859200;
      47311: inst = 32'd136314880;
      47312: inst = 32'd268468224;
      47313: inst = 32'd201346261;
      47314: inst = 32'd203483685;
      47315: inst = 32'd471859200;
      47316: inst = 32'd136314880;
      47317: inst = 32'd268468224;
      47318: inst = 32'd201346262;
      47319: inst = 32'd203483685;
      47320: inst = 32'd471859200;
      47321: inst = 32'd136314880;
      47322: inst = 32'd268468224;
      47323: inst = 32'd201346263;
      47324: inst = 32'd203483685;
      47325: inst = 32'd471859200;
      47326: inst = 32'd136314880;
      47327: inst = 32'd268468224;
      47328: inst = 32'd201346264;
      47329: inst = 32'd203423744;
      47330: inst = 32'd471859200;
      47331: inst = 32'd136314880;
      47332: inst = 32'd268468224;
      47333: inst = 32'd201346265;
      47334: inst = 32'd203423744;
      47335: inst = 32'd471859200;
      47336: inst = 32'd136314880;
      47337: inst = 32'd268468224;
      47338: inst = 32'd201346266;
      47339: inst = 32'd203423744;
      47340: inst = 32'd471859200;
      47341: inst = 32'd136314880;
      47342: inst = 32'd268468224;
      47343: inst = 32'd201346267;
      47344: inst = 32'd203423744;
      47345: inst = 32'd471859200;
      47346: inst = 32'd136314880;
      47347: inst = 32'd268468224;
      47348: inst = 32'd201346268;
      47349: inst = 32'd203423744;
      47350: inst = 32'd471859200;
      47351: inst = 32'd136314880;
      47352: inst = 32'd268468224;
      47353: inst = 32'd201346269;
      47354: inst = 32'd203423744;
      47355: inst = 32'd471859200;
      47356: inst = 32'd136314880;
      47357: inst = 32'd268468224;
      47358: inst = 32'd201346270;
      47359: inst = 32'd203483685;
      47360: inst = 32'd471859200;
      47361: inst = 32'd136314880;
      47362: inst = 32'd268468224;
      47363: inst = 32'd201346271;
      47364: inst = 32'd203483685;
      47365: inst = 32'd471859200;
      47366: inst = 32'd136314880;
      47367: inst = 32'd268468224;
      47368: inst = 32'd201346272;
      47369: inst = 32'd203483685;
      47370: inst = 32'd471859200;
      47371: inst = 32'd136314880;
      47372: inst = 32'd268468224;
      47373: inst = 32'd201346273;
      47374: inst = 32'd203483685;
      47375: inst = 32'd471859200;
      47376: inst = 32'd136314880;
      47377: inst = 32'd268468224;
      47378: inst = 32'd201346274;
      47379: inst = 32'd203483685;
      47380: inst = 32'd471859200;
      47381: inst = 32'd136314880;
      47382: inst = 32'd268468224;
      47383: inst = 32'd201346275;
      47384: inst = 32'd203483685;
      47385: inst = 32'd471859200;
      47386: inst = 32'd136314880;
      47387: inst = 32'd268468224;
      47388: inst = 32'd201346276;
      47389: inst = 32'd203483685;
      47390: inst = 32'd471859200;
      47391: inst = 32'd136314880;
      47392: inst = 32'd268468224;
      47393: inst = 32'd201346277;
      47394: inst = 32'd203483685;
      47395: inst = 32'd471859200;
      47396: inst = 32'd136314880;
      47397: inst = 32'd268468224;
      47398: inst = 32'd201346278;
      47399: inst = 32'd203483685;
      47400: inst = 32'd471859200;
      47401: inst = 32'd136314880;
      47402: inst = 32'd268468224;
      47403: inst = 32'd201346279;
      47404: inst = 32'd203483685;
      47405: inst = 32'd471859200;
      47406: inst = 32'd136314880;
      47407: inst = 32'd268468224;
      47408: inst = 32'd201346280;
      47409: inst = 32'd203483685;
      47410: inst = 32'd471859200;
      47411: inst = 32'd136314880;
      47412: inst = 32'd268468224;
      47413: inst = 32'd201346281;
      47414: inst = 32'd203423744;
      47415: inst = 32'd471859200;
      47416: inst = 32'd136314880;
      47417: inst = 32'd268468224;
      47418: inst = 32'd201346282;
      47419: inst = 32'd203483685;
      47420: inst = 32'd471859200;
      47421: inst = 32'd136314880;
      47422: inst = 32'd268468224;
      47423: inst = 32'd201346283;
      47424: inst = 32'd203483685;
      47425: inst = 32'd471859200;
      47426: inst = 32'd136314880;
      47427: inst = 32'd268468224;
      47428: inst = 32'd201346284;
      47429: inst = 32'd203483685;
      47430: inst = 32'd471859200;
      47431: inst = 32'd136314880;
      47432: inst = 32'd268468224;
      47433: inst = 32'd201346285;
      47434: inst = 32'd203483685;
      47435: inst = 32'd471859200;
      47436: inst = 32'd136314880;
      47437: inst = 32'd268468224;
      47438: inst = 32'd201346286;
      47439: inst = 32'd203483685;
      47440: inst = 32'd471859200;
      47441: inst = 32'd136314880;
      47442: inst = 32'd268468224;
      47443: inst = 32'd201346287;
      47444: inst = 32'd203483685;
      47445: inst = 32'd471859200;
      47446: inst = 32'd136314880;
      47447: inst = 32'd268468224;
      47448: inst = 32'd201346288;
      47449: inst = 32'd203483685;
      47450: inst = 32'd471859200;
      47451: inst = 32'd136314880;
      47452: inst = 32'd268468224;
      47453: inst = 32'd201346289;
      47454: inst = 32'd203483685;
      47455: inst = 32'd471859200;
      47456: inst = 32'd136314880;
      47457: inst = 32'd268468224;
      47458: inst = 32'd201346290;
      47459: inst = 32'd203483685;
      47460: inst = 32'd471859200;
      47461: inst = 32'd136314880;
      47462: inst = 32'd268468224;
      47463: inst = 32'd201346291;
      47464: inst = 32'd203483685;
      47465: inst = 32'd471859200;
      47466: inst = 32'd136314880;
      47467: inst = 32'd268468224;
      47468: inst = 32'd201346292;
      47469: inst = 32'd203483685;
      47470: inst = 32'd471859200;
      47471: inst = 32'd136314880;
      47472: inst = 32'd268468224;
      47473: inst = 32'd201346293;
      47474: inst = 32'd203483685;
      47475: inst = 32'd471859200;
      47476: inst = 32'd136314880;
      47477: inst = 32'd268468224;
      47478: inst = 32'd201346294;
      47479: inst = 32'd203423744;
      47480: inst = 32'd471859200;
      47481: inst = 32'd136314880;
      47482: inst = 32'd268468224;
      47483: inst = 32'd201346295;
      47484: inst = 32'd203423744;
      47485: inst = 32'd471859200;
      47486: inst = 32'd136314880;
      47487: inst = 32'd268468224;
      47488: inst = 32'd201346296;
      47489: inst = 32'd203423744;
      47490: inst = 32'd471859200;
      47491: inst = 32'd136314880;
      47492: inst = 32'd268468224;
      47493: inst = 32'd201346297;
      47494: inst = 32'd203423744;
      47495: inst = 32'd471859200;
      47496: inst = 32'd136314880;
      47497: inst = 32'd268468224;
      47498: inst = 32'd201346298;
      47499: inst = 32'd203423744;
      47500: inst = 32'd471859200;
      47501: inst = 32'd136314880;
      47502: inst = 32'd268468224;
      47503: inst = 32'd201346299;
      47504: inst = 32'd203423744;
      47505: inst = 32'd471859200;
      47506: inst = 32'd136314880;
      47507: inst = 32'd268468224;
      47508: inst = 32'd201346300;
      47509: inst = 32'd203423744;
      47510: inst = 32'd471859200;
      47511: inst = 32'd136314880;
      47512: inst = 32'd268468224;
      47513: inst = 32'd201346301;
      47514: inst = 32'd203423744;
      47515: inst = 32'd471859200;
      47516: inst = 32'd136314880;
      47517: inst = 32'd268468224;
      47518: inst = 32'd201346302;
      47519: inst = 32'd203423744;
      47520: inst = 32'd471859200;
      47521: inst = 32'd136314880;
      47522: inst = 32'd268468224;
      47523: inst = 32'd201346303;
      47524: inst = 32'd203423744;
      47525: inst = 32'd471859200;
      47526: inst = 32'd136314880;
      47527: inst = 32'd268468224;
      47528: inst = 32'd201346304;
      47529: inst = 32'd203423744;
      47530: inst = 32'd471859200;
      47531: inst = 32'd136314880;
      47532: inst = 32'd268468224;
      47533: inst = 32'd201346305;
      47534: inst = 32'd203423744;
      47535: inst = 32'd471859200;
      47536: inst = 32'd136314880;
      47537: inst = 32'd268468224;
      47538: inst = 32'd201346306;
      47539: inst = 32'd203423744;
      47540: inst = 32'd471859200;
      47541: inst = 32'd136314880;
      47542: inst = 32'd268468224;
      47543: inst = 32'd201346307;
      47544: inst = 32'd203423744;
      47545: inst = 32'd471859200;
      47546: inst = 32'd136314880;
      47547: inst = 32'd268468224;
      47548: inst = 32'd201346308;
      47549: inst = 32'd203423744;
      47550: inst = 32'd471859200;
      47551: inst = 32'd136314880;
      47552: inst = 32'd268468224;
      47553: inst = 32'd201346309;
      47554: inst = 32'd203423744;
      47555: inst = 32'd471859200;
      47556: inst = 32'd136314880;
      47557: inst = 32'd268468224;
      47558: inst = 32'd201346310;
      47559: inst = 32'd203423744;
      47560: inst = 32'd471859200;
      47561: inst = 32'd136314880;
      47562: inst = 32'd268468224;
      47563: inst = 32'd201346311;
      47564: inst = 32'd203423744;
      47565: inst = 32'd471859200;
      47566: inst = 32'd136314880;
      47567: inst = 32'd268468224;
      47568: inst = 32'd201346312;
      47569: inst = 32'd203423744;
      47570: inst = 32'd471859200;
      47571: inst = 32'd136314880;
      47572: inst = 32'd268468224;
      47573: inst = 32'd201346313;
      47574: inst = 32'd203423744;
      47575: inst = 32'd471859200;
      47576: inst = 32'd136314880;
      47577: inst = 32'd268468224;
      47578: inst = 32'd201346314;
      47579: inst = 32'd203423744;
      47580: inst = 32'd471859200;
      47581: inst = 32'd136314880;
      47582: inst = 32'd268468224;
      47583: inst = 32'd201346315;
      47584: inst = 32'd203423744;
      47585: inst = 32'd471859200;
      47586: inst = 32'd136314880;
      47587: inst = 32'd268468224;
      47588: inst = 32'd201346316;
      47589: inst = 32'd203423744;
      47590: inst = 32'd471859200;
      47591: inst = 32'd136314880;
      47592: inst = 32'd268468224;
      47593: inst = 32'd201346317;
      47594: inst = 32'd203483685;
      47595: inst = 32'd471859200;
      47596: inst = 32'd136314880;
      47597: inst = 32'd268468224;
      47598: inst = 32'd201346318;
      47599: inst = 32'd203483685;
      47600: inst = 32'd471859200;
      47601: inst = 32'd136314880;
      47602: inst = 32'd268468224;
      47603: inst = 32'd201346319;
      47604: inst = 32'd203483685;
      47605: inst = 32'd471859200;
      47606: inst = 32'd136314880;
      47607: inst = 32'd268468224;
      47608: inst = 32'd201346320;
      47609: inst = 32'd203423744;
      47610: inst = 32'd471859200;
      47611: inst = 32'd136314880;
      47612: inst = 32'd268468224;
      47613: inst = 32'd201346321;
      47614: inst = 32'd203423744;
      47615: inst = 32'd471859200;
      47616: inst = 32'd136314880;
      47617: inst = 32'd268468224;
      47618: inst = 32'd201346322;
      47619: inst = 32'd203423744;
      47620: inst = 32'd471859200;
      47621: inst = 32'd136314880;
      47622: inst = 32'd268468224;
      47623: inst = 32'd201346323;
      47624: inst = 32'd203423744;
      47625: inst = 32'd471859200;
      47626: inst = 32'd136314880;
      47627: inst = 32'd268468224;
      47628: inst = 32'd201346324;
      47629: inst = 32'd203423744;
      47630: inst = 32'd471859200;
      47631: inst = 32'd136314880;
      47632: inst = 32'd268468224;
      47633: inst = 32'd201346325;
      47634: inst = 32'd203423744;
      47635: inst = 32'd471859200;
      47636: inst = 32'd136314880;
      47637: inst = 32'd268468224;
      47638: inst = 32'd201346326;
      47639: inst = 32'd203423744;
      47640: inst = 32'd471859200;
      47641: inst = 32'd136314880;
      47642: inst = 32'd268468224;
      47643: inst = 32'd201346327;
      47644: inst = 32'd203423744;
      47645: inst = 32'd471859200;
      47646: inst = 32'd136314880;
      47647: inst = 32'd268468224;
      47648: inst = 32'd201346328;
      47649: inst = 32'd203423744;
      47650: inst = 32'd471859200;
      47651: inst = 32'd136314880;
      47652: inst = 32'd268468224;
      47653: inst = 32'd201346329;
      47654: inst = 32'd203423744;
      47655: inst = 32'd471859200;
      47656: inst = 32'd136314880;
      47657: inst = 32'd268468224;
      47658: inst = 32'd201346330;
      47659: inst = 32'd203423744;
      47660: inst = 32'd471859200;
      47661: inst = 32'd136314880;
      47662: inst = 32'd268468224;
      47663: inst = 32'd201346331;
      47664: inst = 32'd203483685;
      47665: inst = 32'd471859200;
      47666: inst = 32'd136314880;
      47667: inst = 32'd268468224;
      47668: inst = 32'd201346332;
      47669: inst = 32'd203483685;
      47670: inst = 32'd471859200;
      47671: inst = 32'd136314880;
      47672: inst = 32'd268468224;
      47673: inst = 32'd201346333;
      47674: inst = 32'd203483685;
      47675: inst = 32'd471859200;
      47676: inst = 32'd136314880;
      47677: inst = 32'd268468224;
      47678: inst = 32'd201346334;
      47679: inst = 32'd203483685;
      47680: inst = 32'd471859200;
      47681: inst = 32'd136314880;
      47682: inst = 32'd268468224;
      47683: inst = 32'd201346335;
      47684: inst = 32'd203483685;
      47685: inst = 32'd471859200;
      47686: inst = 32'd136314880;
      47687: inst = 32'd268468224;
      47688: inst = 32'd201346336;
      47689: inst = 32'd203423744;
      47690: inst = 32'd471859200;
      47691: inst = 32'd136314880;
      47692: inst = 32'd268468224;
      47693: inst = 32'd201346337;
      47694: inst = 32'd203423744;
      47695: inst = 32'd471859200;
      47696: inst = 32'd136314880;
      47697: inst = 32'd268468224;
      47698: inst = 32'd201346338;
      47699: inst = 32'd203423744;
      47700: inst = 32'd471859200;
      47701: inst = 32'd136314880;
      47702: inst = 32'd268468224;
      47703: inst = 32'd201346339;
      47704: inst = 32'd203423744;
      47705: inst = 32'd471859200;
      47706: inst = 32'd136314880;
      47707: inst = 32'd268468224;
      47708: inst = 32'd201346340;
      47709: inst = 32'd203423744;
      47710: inst = 32'd471859200;
      47711: inst = 32'd136314880;
      47712: inst = 32'd268468224;
      47713: inst = 32'd201346341;
      47714: inst = 32'd203483685;
      47715: inst = 32'd471859200;
      47716: inst = 32'd136314880;
      47717: inst = 32'd268468224;
      47718: inst = 32'd201346342;
      47719: inst = 32'd203483685;
      47720: inst = 32'd471859200;
      47721: inst = 32'd136314880;
      47722: inst = 32'd268468224;
      47723: inst = 32'd201346343;
      47724: inst = 32'd203483685;
      47725: inst = 32'd471859200;
      47726: inst = 32'd136314880;
      47727: inst = 32'd268468224;
      47728: inst = 32'd201346344;
      47729: inst = 32'd203483685;
      47730: inst = 32'd471859200;
      47731: inst = 32'd136314880;
      47732: inst = 32'd268468224;
      47733: inst = 32'd201346345;
      47734: inst = 32'd203423744;
      47735: inst = 32'd471859200;
      47736: inst = 32'd136314880;
      47737: inst = 32'd268468224;
      47738: inst = 32'd201346346;
      47739: inst = 32'd203423744;
      47740: inst = 32'd471859200;
      47741: inst = 32'd136314880;
      47742: inst = 32'd268468224;
      47743: inst = 32'd201346347;
      47744: inst = 32'd203423744;
      47745: inst = 32'd471859200;
      47746: inst = 32'd136314880;
      47747: inst = 32'd268468224;
      47748: inst = 32'd201346348;
      47749: inst = 32'd203423744;
      47750: inst = 32'd471859200;
      47751: inst = 32'd136314880;
      47752: inst = 32'd268468224;
      47753: inst = 32'd201346349;
      47754: inst = 32'd203423744;
      47755: inst = 32'd471859200;
      47756: inst = 32'd136314880;
      47757: inst = 32'd268468224;
      47758: inst = 32'd201346350;
      47759: inst = 32'd203483685;
      47760: inst = 32'd471859200;
      47761: inst = 32'd136314880;
      47762: inst = 32'd268468224;
      47763: inst = 32'd201346351;
      47764: inst = 32'd203483685;
      47765: inst = 32'd471859200;
      47766: inst = 32'd136314880;
      47767: inst = 32'd268468224;
      47768: inst = 32'd201346352;
      47769: inst = 32'd203423744;
      47770: inst = 32'd471859200;
      47771: inst = 32'd136314880;
      47772: inst = 32'd268468224;
      47773: inst = 32'd201346353;
      47774: inst = 32'd203483685;
      47775: inst = 32'd471859200;
      47776: inst = 32'd136314880;
      47777: inst = 32'd268468224;
      47778: inst = 32'd201346354;
      47779: inst = 32'd203483685;
      47780: inst = 32'd471859200;
      47781: inst = 32'd136314880;
      47782: inst = 32'd268468224;
      47783: inst = 32'd201346355;
      47784: inst = 32'd203483685;
      47785: inst = 32'd471859200;
      47786: inst = 32'd136314880;
      47787: inst = 32'd268468224;
      47788: inst = 32'd201346356;
      47789: inst = 32'd203483685;
      47790: inst = 32'd471859200;
      47791: inst = 32'd136314880;
      47792: inst = 32'd268468224;
      47793: inst = 32'd201346357;
      47794: inst = 32'd203483685;
      47795: inst = 32'd471859200;
      47796: inst = 32'd136314880;
      47797: inst = 32'd268468224;
      47798: inst = 32'd201346358;
      47799: inst = 32'd203483685;
      47800: inst = 32'd471859200;
      47801: inst = 32'd136314880;
      47802: inst = 32'd268468224;
      47803: inst = 32'd201346359;
      47804: inst = 32'd203483685;
      47805: inst = 32'd471859200;
      47806: inst = 32'd136314880;
      47807: inst = 32'd268468224;
      47808: inst = 32'd201346360;
      47809: inst = 32'd203483685;
      47810: inst = 32'd471859200;
      47811: inst = 32'd136314880;
      47812: inst = 32'd268468224;
      47813: inst = 32'd201346361;
      47814: inst = 32'd203423744;
      47815: inst = 32'd471859200;
      47816: inst = 32'd136314880;
      47817: inst = 32'd268468224;
      47818: inst = 32'd201346362;
      47819: inst = 32'd203423744;
      47820: inst = 32'd471859200;
      47821: inst = 32'd136314880;
      47822: inst = 32'd268468224;
      47823: inst = 32'd201346363;
      47824: inst = 32'd203423744;
      47825: inst = 32'd471859200;
      47826: inst = 32'd136314880;
      47827: inst = 32'd268468224;
      47828: inst = 32'd201346364;
      47829: inst = 32'd203423744;
      47830: inst = 32'd471859200;
      47831: inst = 32'd136314880;
      47832: inst = 32'd268468224;
      47833: inst = 32'd201346365;
      47834: inst = 32'd203423744;
      47835: inst = 32'd471859200;
      47836: inst = 32'd136314880;
      47837: inst = 32'd268468224;
      47838: inst = 32'd201346366;
      47839: inst = 32'd203483685;
      47840: inst = 32'd471859200;
      47841: inst = 32'd136314880;
      47842: inst = 32'd268468224;
      47843: inst = 32'd201346367;
      47844: inst = 32'd203483685;
      47845: inst = 32'd471859200;
      47846: inst = 32'd136314880;
      47847: inst = 32'd268468224;
      47848: inst = 32'd201346368;
      47849: inst = 32'd203483685;
      47850: inst = 32'd471859200;
      47851: inst = 32'd136314880;
      47852: inst = 32'd268468224;
      47853: inst = 32'd201346369;
      47854: inst = 32'd203423744;
      47855: inst = 32'd471859200;
      47856: inst = 32'd136314880;
      47857: inst = 32'd268468224;
      47858: inst = 32'd201346370;
      47859: inst = 32'd203423744;
      47860: inst = 32'd471859200;
      47861: inst = 32'd136314880;
      47862: inst = 32'd268468224;
      47863: inst = 32'd201346371;
      47864: inst = 32'd203483685;
      47865: inst = 32'd471859200;
      47866: inst = 32'd136314880;
      47867: inst = 32'd268468224;
      47868: inst = 32'd201346372;
      47869: inst = 32'd203483685;
      47870: inst = 32'd471859200;
      47871: inst = 32'd136314880;
      47872: inst = 32'd268468224;
      47873: inst = 32'd201346373;
      47874: inst = 32'd203483685;
      47875: inst = 32'd471859200;
      47876: inst = 32'd136314880;
      47877: inst = 32'd268468224;
      47878: inst = 32'd201346374;
      47879: inst = 32'd203483685;
      47880: inst = 32'd471859200;
      47881: inst = 32'd136314880;
      47882: inst = 32'd268468224;
      47883: inst = 32'd201346375;
      47884: inst = 32'd203483685;
      47885: inst = 32'd471859200;
      47886: inst = 32'd136314880;
      47887: inst = 32'd268468224;
      47888: inst = 32'd201346376;
      47889: inst = 32'd203423744;
      47890: inst = 32'd471859200;
      47891: inst = 32'd136314880;
      47892: inst = 32'd268468224;
      47893: inst = 32'd201346377;
      47894: inst = 32'd203423744;
      47895: inst = 32'd471859200;
      47896: inst = 32'd136314880;
      47897: inst = 32'd268468224;
      47898: inst = 32'd201346378;
      47899: inst = 32'd203483685;
      47900: inst = 32'd471859200;
      47901: inst = 32'd136314880;
      47902: inst = 32'd268468224;
      47903: inst = 32'd201346379;
      47904: inst = 32'd203483685;
      47905: inst = 32'd471859200;
      47906: inst = 32'd136314880;
      47907: inst = 32'd268468224;
      47908: inst = 32'd201346380;
      47909: inst = 32'd203483685;
      47910: inst = 32'd471859200;
      47911: inst = 32'd136314880;
      47912: inst = 32'd268468224;
      47913: inst = 32'd201346381;
      47914: inst = 32'd203483685;
      47915: inst = 32'd471859200;
      47916: inst = 32'd136314880;
      47917: inst = 32'd268468224;
      47918: inst = 32'd201346382;
      47919: inst = 32'd203423744;
      47920: inst = 32'd471859200;
      47921: inst = 32'd136314880;
      47922: inst = 32'd268468224;
      47923: inst = 32'd201346383;
      47924: inst = 32'd203423744;
      47925: inst = 32'd471859200;
      47926: inst = 32'd136314880;
      47927: inst = 32'd268468224;
      47928: inst = 32'd201346384;
      47929: inst = 32'd203423744;
      47930: inst = 32'd471859200;
      47931: inst = 32'd136314880;
      47932: inst = 32'd268468224;
      47933: inst = 32'd201346385;
      47934: inst = 32'd203423744;
      47935: inst = 32'd471859200;
      47936: inst = 32'd136314880;
      47937: inst = 32'd268468224;
      47938: inst = 32'd201346386;
      47939: inst = 32'd203423744;
      47940: inst = 32'd471859200;
      47941: inst = 32'd136314880;
      47942: inst = 32'd268468224;
      47943: inst = 32'd201346387;
      47944: inst = 32'd203423744;
      47945: inst = 32'd471859200;
      47946: inst = 32'd136314880;
      47947: inst = 32'd268468224;
      47948: inst = 32'd201346388;
      47949: inst = 32'd203423744;
      47950: inst = 32'd471859200;
      47951: inst = 32'd136314880;
      47952: inst = 32'd268468224;
      47953: inst = 32'd201346389;
      47954: inst = 32'd203423744;
      47955: inst = 32'd471859200;
      47956: inst = 32'd136314880;
      47957: inst = 32'd268468224;
      47958: inst = 32'd201346390;
      47959: inst = 32'd203423744;
      47960: inst = 32'd471859200;
      47961: inst = 32'd136314880;
      47962: inst = 32'd268468224;
      47963: inst = 32'd201346391;
      47964: inst = 32'd203423744;
      47965: inst = 32'd471859200;
      47966: inst = 32'd136314880;
      47967: inst = 32'd268468224;
      47968: inst = 32'd201346392;
      47969: inst = 32'd203423744;
      47970: inst = 32'd471859200;
      47971: inst = 32'd136314880;
      47972: inst = 32'd268468224;
      47973: inst = 32'd201346393;
      47974: inst = 32'd203423744;
      47975: inst = 32'd471859200;
      47976: inst = 32'd136314880;
      47977: inst = 32'd268468224;
      47978: inst = 32'd201346394;
      47979: inst = 32'd203423744;
      47980: inst = 32'd471859200;
      47981: inst = 32'd136314880;
      47982: inst = 32'd268468224;
      47983: inst = 32'd201346395;
      47984: inst = 32'd203423744;
      47985: inst = 32'd471859200;
      47986: inst = 32'd136314880;
      47987: inst = 32'd268468224;
      47988: inst = 32'd201346396;
      47989: inst = 32'd203423744;
      47990: inst = 32'd471859200;
      47991: inst = 32'd136314880;
      47992: inst = 32'd268468224;
      47993: inst = 32'd201346397;
      47994: inst = 32'd203423744;
      47995: inst = 32'd471859200;
      47996: inst = 32'd136314880;
      47997: inst = 32'd268468224;
      47998: inst = 32'd201346398;
      47999: inst = 32'd203423744;
      48000: inst = 32'd471859200;
      48001: inst = 32'd136314880;
      48002: inst = 32'd268468224;
      48003: inst = 32'd201346399;
      48004: inst = 32'd203423744;
      48005: inst = 32'd471859200;
      48006: inst = 32'd136314880;
      48007: inst = 32'd268468224;
      48008: inst = 32'd201346400;
      48009: inst = 32'd203423744;
      48010: inst = 32'd471859200;
      48011: inst = 32'd136314880;
      48012: inst = 32'd268468224;
      48013: inst = 32'd201346401;
      48014: inst = 32'd203423744;
      48015: inst = 32'd471859200;
      48016: inst = 32'd136314880;
      48017: inst = 32'd268468224;
      48018: inst = 32'd201346402;
      48019: inst = 32'd203423744;
      48020: inst = 32'd471859200;
      48021: inst = 32'd136314880;
      48022: inst = 32'd268468224;
      48023: inst = 32'd201346403;
      48024: inst = 32'd203423744;
      48025: inst = 32'd471859200;
      48026: inst = 32'd136314880;
      48027: inst = 32'd268468224;
      48028: inst = 32'd201346404;
      48029: inst = 32'd203423744;
      48030: inst = 32'd471859200;
      48031: inst = 32'd136314880;
      48032: inst = 32'd268468224;
      48033: inst = 32'd201346405;
      48034: inst = 32'd203423744;
      48035: inst = 32'd471859200;
      48036: inst = 32'd136314880;
      48037: inst = 32'd268468224;
      48038: inst = 32'd201346406;
      48039: inst = 32'd203423744;
      48040: inst = 32'd471859200;
      48041: inst = 32'd136314880;
      48042: inst = 32'd268468224;
      48043: inst = 32'd201346407;
      48044: inst = 32'd203423744;
      48045: inst = 32'd471859200;
      48046: inst = 32'd136314880;
      48047: inst = 32'd268468224;
      48048: inst = 32'd201346408;
      48049: inst = 32'd203423744;
      48050: inst = 32'd471859200;
      48051: inst = 32'd136314880;
      48052: inst = 32'd268468224;
      48053: inst = 32'd201346409;
      48054: inst = 32'd203423744;
      48055: inst = 32'd471859200;
      48056: inst = 32'd136314880;
      48057: inst = 32'd268468224;
      48058: inst = 32'd201346410;
      48059: inst = 32'd203423744;
      48060: inst = 32'd471859200;
      48061: inst = 32'd136314880;
      48062: inst = 32'd268468224;
      48063: inst = 32'd201346411;
      48064: inst = 32'd203423744;
      48065: inst = 32'd471859200;
      48066: inst = 32'd136314880;
      48067: inst = 32'd268468224;
      48068: inst = 32'd201346412;
      48069: inst = 32'd203423744;
      48070: inst = 32'd471859200;
      48071: inst = 32'd136314880;
      48072: inst = 32'd268468224;
      48073: inst = 32'd201346413;
      48074: inst = 32'd203483685;
      48075: inst = 32'd471859200;
      48076: inst = 32'd136314880;
      48077: inst = 32'd268468224;
      48078: inst = 32'd201346414;
      48079: inst = 32'd203483685;
      48080: inst = 32'd471859200;
      48081: inst = 32'd136314880;
      48082: inst = 32'd268468224;
      48083: inst = 32'd201346415;
      48084: inst = 32'd203483685;
      48085: inst = 32'd471859200;
      48086: inst = 32'd136314880;
      48087: inst = 32'd268468224;
      48088: inst = 32'd201346416;
      48089: inst = 32'd203483685;
      48090: inst = 32'd471859200;
      48091: inst = 32'd136314880;
      48092: inst = 32'd268468224;
      48093: inst = 32'd201346417;
      48094: inst = 32'd203483685;
      48095: inst = 32'd471859200;
      48096: inst = 32'd136314880;
      48097: inst = 32'd268468224;
      48098: inst = 32'd201346418;
      48099: inst = 32'd203483685;
      48100: inst = 32'd471859200;
      48101: inst = 32'd136314880;
      48102: inst = 32'd268468224;
      48103: inst = 32'd201346419;
      48104: inst = 32'd203483685;
      48105: inst = 32'd471859200;
      48106: inst = 32'd136314880;
      48107: inst = 32'd268468224;
      48108: inst = 32'd201346420;
      48109: inst = 32'd203483685;
      48110: inst = 32'd471859200;
      48111: inst = 32'd136314880;
      48112: inst = 32'd268468224;
      48113: inst = 32'd201346421;
      48114: inst = 32'd203423744;
      48115: inst = 32'd471859200;
      48116: inst = 32'd136314880;
      48117: inst = 32'd268468224;
      48118: inst = 32'd201346422;
      48119: inst = 32'd203423744;
      48120: inst = 32'd471859200;
      48121: inst = 32'd136314880;
      48122: inst = 32'd268468224;
      48123: inst = 32'd201346423;
      48124: inst = 32'd203423744;
      48125: inst = 32'd471859200;
      48126: inst = 32'd136314880;
      48127: inst = 32'd268468224;
      48128: inst = 32'd201346424;
      48129: inst = 32'd203423744;
      48130: inst = 32'd471859200;
      48131: inst = 32'd136314880;
      48132: inst = 32'd268468224;
      48133: inst = 32'd201346425;
      48134: inst = 32'd203423744;
      48135: inst = 32'd471859200;
      48136: inst = 32'd136314880;
      48137: inst = 32'd268468224;
      48138: inst = 32'd201346426;
      48139: inst = 32'd203423744;
      48140: inst = 32'd471859200;
      48141: inst = 32'd136314880;
      48142: inst = 32'd268468224;
      48143: inst = 32'd201346427;
      48144: inst = 32'd203423744;
      48145: inst = 32'd471859200;
      48146: inst = 32'd136314880;
      48147: inst = 32'd268468224;
      48148: inst = 32'd201346428;
      48149: inst = 32'd203483685;
      48150: inst = 32'd471859200;
      48151: inst = 32'd136314880;
      48152: inst = 32'd268468224;
      48153: inst = 32'd201346429;
      48154: inst = 32'd203483685;
      48155: inst = 32'd471859200;
      48156: inst = 32'd136314880;
      48157: inst = 32'd268468224;
      48158: inst = 32'd201346430;
      48159: inst = 32'd203483685;
      48160: inst = 32'd471859200;
      48161: inst = 32'd136314880;
      48162: inst = 32'd268468224;
      48163: inst = 32'd201346431;
      48164: inst = 32'd203483685;
      48165: inst = 32'd471859200;
      48166: inst = 32'd136314880;
      48167: inst = 32'd268468224;
      48168: inst = 32'd201346432;
      48169: inst = 32'd203483685;
      48170: inst = 32'd471859200;
      48171: inst = 32'd136314880;
      48172: inst = 32'd268468224;
      48173: inst = 32'd201346433;
      48174: inst = 32'd203423744;
      48175: inst = 32'd471859200;
      48176: inst = 32'd136314880;
      48177: inst = 32'd268468224;
      48178: inst = 32'd201346434;
      48179: inst = 32'd203423744;
      48180: inst = 32'd471859200;
      48181: inst = 32'd136314880;
      48182: inst = 32'd268468224;
      48183: inst = 32'd201346435;
      48184: inst = 32'd203423744;
      48185: inst = 32'd471859200;
      48186: inst = 32'd136314880;
      48187: inst = 32'd268468224;
      48188: inst = 32'd201346436;
      48189: inst = 32'd203423744;
      48190: inst = 32'd471859200;
      48191: inst = 32'd136314880;
      48192: inst = 32'd268468224;
      48193: inst = 32'd201346437;
      48194: inst = 32'd203483685;
      48195: inst = 32'd471859200;
      48196: inst = 32'd136314880;
      48197: inst = 32'd268468224;
      48198: inst = 32'd201346438;
      48199: inst = 32'd203483685;
      48200: inst = 32'd471859200;
      48201: inst = 32'd136314880;
      48202: inst = 32'd268468224;
      48203: inst = 32'd201346439;
      48204: inst = 32'd203483685;
      48205: inst = 32'd471859200;
      48206: inst = 32'd136314880;
      48207: inst = 32'd268468224;
      48208: inst = 32'd201346440;
      48209: inst = 32'd203483685;
      48210: inst = 32'd471859200;
      48211: inst = 32'd136314880;
      48212: inst = 32'd268468224;
      48213: inst = 32'd201346441;
      48214: inst = 32'd203423744;
      48215: inst = 32'd471859200;
      48216: inst = 32'd136314880;
      48217: inst = 32'd268468224;
      48218: inst = 32'd201346442;
      48219: inst = 32'd203423744;
      48220: inst = 32'd471859200;
      48221: inst = 32'd136314880;
      48222: inst = 32'd268468224;
      48223: inst = 32'd201346443;
      48224: inst = 32'd203423744;
      48225: inst = 32'd471859200;
      48226: inst = 32'd136314880;
      48227: inst = 32'd268468224;
      48228: inst = 32'd201346444;
      48229: inst = 32'd203423744;
      48230: inst = 32'd471859200;
      48231: inst = 32'd136314880;
      48232: inst = 32'd268468224;
      48233: inst = 32'd201346445;
      48234: inst = 32'd203483685;
      48235: inst = 32'd471859200;
      48236: inst = 32'd136314880;
      48237: inst = 32'd268468224;
      48238: inst = 32'd201346446;
      48239: inst = 32'd203483685;
      48240: inst = 32'd471859200;
      48241: inst = 32'd136314880;
      48242: inst = 32'd268468224;
      48243: inst = 32'd201346447;
      48244: inst = 32'd203423744;
      48245: inst = 32'd471859200;
      48246: inst = 32'd136314880;
      48247: inst = 32'd268468224;
      48248: inst = 32'd201346448;
      48249: inst = 32'd203423744;
      48250: inst = 32'd471859200;
      48251: inst = 32'd136314880;
      48252: inst = 32'd268468224;
      48253: inst = 32'd201346449;
      48254: inst = 32'd203483685;
      48255: inst = 32'd471859200;
      48256: inst = 32'd136314880;
      48257: inst = 32'd268468224;
      48258: inst = 32'd201346450;
      48259: inst = 32'd203483685;
      48260: inst = 32'd471859200;
      48261: inst = 32'd136314880;
      48262: inst = 32'd268468224;
      48263: inst = 32'd201346451;
      48264: inst = 32'd203483685;
      48265: inst = 32'd471859200;
      48266: inst = 32'd136314880;
      48267: inst = 32'd268468224;
      48268: inst = 32'd201346452;
      48269: inst = 32'd203483685;
      48270: inst = 32'd471859200;
      48271: inst = 32'd136314880;
      48272: inst = 32'd268468224;
      48273: inst = 32'd201346453;
      48274: inst = 32'd203483685;
      48275: inst = 32'd471859200;
      48276: inst = 32'd136314880;
      48277: inst = 32'd268468224;
      48278: inst = 32'd201346454;
      48279: inst = 32'd203483685;
      48280: inst = 32'd471859200;
      48281: inst = 32'd136314880;
      48282: inst = 32'd268468224;
      48283: inst = 32'd201346455;
      48284: inst = 32'd203483685;
      48285: inst = 32'd471859200;
      48286: inst = 32'd136314880;
      48287: inst = 32'd268468224;
      48288: inst = 32'd201346456;
      48289: inst = 32'd203483685;
      48290: inst = 32'd471859200;
      48291: inst = 32'd136314880;
      48292: inst = 32'd268468224;
      48293: inst = 32'd201346457;
      48294: inst = 32'd203483685;
      48295: inst = 32'd471859200;
      48296: inst = 32'd136314880;
      48297: inst = 32'd268468224;
      48298: inst = 32'd201346458;
      48299: inst = 32'd203423744;
      48300: inst = 32'd471859200;
      48301: inst = 32'd136314880;
      48302: inst = 32'd268468224;
      48303: inst = 32'd201346459;
      48304: inst = 32'd203423744;
      48305: inst = 32'd471859200;
      48306: inst = 32'd136314880;
      48307: inst = 32'd268468224;
      48308: inst = 32'd201346460;
      48309: inst = 32'd203423744;
      48310: inst = 32'd471859200;
      48311: inst = 32'd136314880;
      48312: inst = 32'd268468224;
      48313: inst = 32'd201346461;
      48314: inst = 32'd203423744;
      48315: inst = 32'd471859200;
      48316: inst = 32'd136314880;
      48317: inst = 32'd268468224;
      48318: inst = 32'd201346462;
      48319: inst = 32'd203483685;
      48320: inst = 32'd471859200;
      48321: inst = 32'd136314880;
      48322: inst = 32'd268468224;
      48323: inst = 32'd201346463;
      48324: inst = 32'd203483685;
      48325: inst = 32'd471859200;
      48326: inst = 32'd136314880;
      48327: inst = 32'd268468224;
      48328: inst = 32'd201346464;
      48329: inst = 32'd203483685;
      48330: inst = 32'd471859200;
      48331: inst = 32'd136314880;
      48332: inst = 32'd268468224;
      48333: inst = 32'd201346465;
      48334: inst = 32'd203483685;
      48335: inst = 32'd471859200;
      48336: inst = 32'd136314880;
      48337: inst = 32'd268468224;
      48338: inst = 32'd201346466;
      48339: inst = 32'd203483685;
      48340: inst = 32'd471859200;
      48341: inst = 32'd136314880;
      48342: inst = 32'd268468224;
      48343: inst = 32'd201346467;
      48344: inst = 32'd203483685;
      48345: inst = 32'd471859200;
      48346: inst = 32'd136314880;
      48347: inst = 32'd268468224;
      48348: inst = 32'd201346468;
      48349: inst = 32'd203483685;
      48350: inst = 32'd471859200;
      48351: inst = 32'd136314880;
      48352: inst = 32'd268468224;
      48353: inst = 32'd201346469;
      48354: inst = 32'd203483685;
      48355: inst = 32'd471859200;
      48356: inst = 32'd136314880;
      48357: inst = 32'd268468224;
      48358: inst = 32'd201346470;
      48359: inst = 32'd203483685;
      48360: inst = 32'd471859200;
      48361: inst = 32'd136314880;
      48362: inst = 32'd268468224;
      48363: inst = 32'd201346471;
      48364: inst = 32'd203423744;
      48365: inst = 32'd471859200;
      48366: inst = 32'd136314880;
      48367: inst = 32'd268468224;
      48368: inst = 32'd201346472;
      48369: inst = 32'd203423744;
      48370: inst = 32'd471859200;
      48371: inst = 32'd136314880;
      48372: inst = 32'd268468224;
      48373: inst = 32'd201346473;
      48374: inst = 32'd203423744;
      48375: inst = 32'd471859200;
      48376: inst = 32'd136314880;
      48377: inst = 32'd268468224;
      48378: inst = 32'd201346474;
      48379: inst = 32'd203483685;
      48380: inst = 32'd471859200;
      48381: inst = 32'd136314880;
      48382: inst = 32'd268468224;
      48383: inst = 32'd201346475;
      48384: inst = 32'd203483685;
      48385: inst = 32'd471859200;
      48386: inst = 32'd136314880;
      48387: inst = 32'd268468224;
      48388: inst = 32'd201346476;
      48389: inst = 32'd203483685;
      48390: inst = 32'd471859200;
      48391: inst = 32'd136314880;
      48392: inst = 32'd268468224;
      48393: inst = 32'd201346477;
      48394: inst = 32'd203483685;
      48395: inst = 32'd471859200;
      48396: inst = 32'd136314880;
      48397: inst = 32'd268468224;
      48398: inst = 32'd201346478;
      48399: inst = 32'd203483685;
      48400: inst = 32'd471859200;
      48401: inst = 32'd136314880;
      48402: inst = 32'd268468224;
      48403: inst = 32'd201346479;
      48404: inst = 32'd203483685;
      48405: inst = 32'd471859200;
      48406: inst = 32'd136314880;
      48407: inst = 32'd268468224;
      48408: inst = 32'd201346480;
      48409: inst = 32'd203483685;
      48410: inst = 32'd471859200;
      48411: inst = 32'd136314880;
      48412: inst = 32'd268468224;
      48413: inst = 32'd201346481;
      48414: inst = 32'd203483685;
      48415: inst = 32'd471859200;
      48416: inst = 32'd136314880;
      48417: inst = 32'd268468224;
      48418: inst = 32'd201346482;
      48419: inst = 32'd203483685;
      48420: inst = 32'd471859200;
      48421: inst = 32'd136314880;
      48422: inst = 32'd268468224;
      48423: inst = 32'd201346483;
      48424: inst = 32'd203423744;
      48425: inst = 32'd471859200;
      48426: inst = 32'd136314880;
      48427: inst = 32'd268468224;
      48428: inst = 32'd201346484;
      48429: inst = 32'd203423744;
      48430: inst = 32'd471859200;
      48431: inst = 32'd136314880;
      48432: inst = 32'd268468224;
      48433: inst = 32'd201346485;
      48434: inst = 32'd203423744;
      48435: inst = 32'd471859200;
      48436: inst = 32'd136314880;
      48437: inst = 32'd268468224;
      48438: inst = 32'd201346486;
      48439: inst = 32'd203423744;
      48440: inst = 32'd471859200;
      48441: inst = 32'd136314880;
      48442: inst = 32'd268468224;
      48443: inst = 32'd201346487;
      48444: inst = 32'd203423744;
      48445: inst = 32'd471859200;
      48446: inst = 32'd136314880;
      48447: inst = 32'd268468224;
      48448: inst = 32'd201346488;
      48449: inst = 32'd203423744;
      48450: inst = 32'd471859200;
      48451: inst = 32'd136314880;
      48452: inst = 32'd268468224;
      48453: inst = 32'd201346489;
      48454: inst = 32'd203423744;
      48455: inst = 32'd471859200;
      48456: inst = 32'd136314880;
      48457: inst = 32'd268468224;
      48458: inst = 32'd201346490;
      48459: inst = 32'd203423744;
      48460: inst = 32'd471859200;
      48461: inst = 32'd136314880;
      48462: inst = 32'd268468224;
      48463: inst = 32'd201346491;
      48464: inst = 32'd203423744;
      48465: inst = 32'd471859200;
      48466: inst = 32'd136314880;
      48467: inst = 32'd268468224;
      48468: inst = 32'd201346492;
      48469: inst = 32'd203423744;
      48470: inst = 32'd471859200;
      48471: inst = 32'd136314880;
      48472: inst = 32'd268468224;
      48473: inst = 32'd201346493;
      48474: inst = 32'd203423744;
      48475: inst = 32'd471859200;
      48476: inst = 32'd136314880;
      48477: inst = 32'd268468224;
      48478: inst = 32'd201346494;
      48479: inst = 32'd203423744;
      48480: inst = 32'd471859200;
      48481: inst = 32'd136314880;
      48482: inst = 32'd268468224;
      48483: inst = 32'd201346495;
      48484: inst = 32'd203423744;
      48485: inst = 32'd471859200;
      48486: inst = 32'd136314880;
      48487: inst = 32'd268468224;
      48488: inst = 32'd201346496;
      48489: inst = 32'd203423744;
      48490: inst = 32'd471859200;
      48491: inst = 32'd136314880;
      48492: inst = 32'd268468224;
      48493: inst = 32'd201346497;
      48494: inst = 32'd203423744;
      48495: inst = 32'd471859200;
      48496: inst = 32'd136314880;
      48497: inst = 32'd268468224;
      48498: inst = 32'd201346498;
      48499: inst = 32'd203423744;
      48500: inst = 32'd471859200;
      48501: inst = 32'd136314880;
      48502: inst = 32'd268468224;
      48503: inst = 32'd201346499;
      48504: inst = 32'd203423744;
      48505: inst = 32'd471859200;
      48506: inst = 32'd136314880;
      48507: inst = 32'd268468224;
      48508: inst = 32'd201346500;
      48509: inst = 32'd203423744;
      48510: inst = 32'd471859200;
      48511: inst = 32'd136314880;
      48512: inst = 32'd268468224;
      48513: inst = 32'd201346501;
      48514: inst = 32'd203423744;
      48515: inst = 32'd471859200;
      48516: inst = 32'd136314880;
      48517: inst = 32'd268468224;
      48518: inst = 32'd201346502;
      48519: inst = 32'd203423744;
      48520: inst = 32'd471859200;
      48521: inst = 32'd136314880;
      48522: inst = 32'd268468224;
      48523: inst = 32'd201346503;
      48524: inst = 32'd203423744;
      48525: inst = 32'd471859200;
      48526: inst = 32'd136314880;
      48527: inst = 32'd268468224;
      48528: inst = 32'd201346504;
      48529: inst = 32'd203423744;
      48530: inst = 32'd471859200;
      48531: inst = 32'd136314880;
      48532: inst = 32'd268468224;
      48533: inst = 32'd201346505;
      48534: inst = 32'd203423744;
      48535: inst = 32'd471859200;
      48536: inst = 32'd136314880;
      48537: inst = 32'd268468224;
      48538: inst = 32'd201346506;
      48539: inst = 32'd203423744;
      48540: inst = 32'd471859200;
      48541: inst = 32'd136314880;
      48542: inst = 32'd268468224;
      48543: inst = 32'd201346507;
      48544: inst = 32'd203423744;
      48545: inst = 32'd471859200;
      48546: inst = 32'd136314880;
      48547: inst = 32'd268468224;
      48548: inst = 32'd201346508;
      48549: inst = 32'd203423744;
      48550: inst = 32'd471859200;
      48551: inst = 32'd136314880;
      48552: inst = 32'd268468224;
      48553: inst = 32'd201346509;
      48554: inst = 32'd203483685;
      48555: inst = 32'd471859200;
      48556: inst = 32'd136314880;
      48557: inst = 32'd268468224;
      48558: inst = 32'd201346510;
      48559: inst = 32'd203483685;
      48560: inst = 32'd471859200;
      48561: inst = 32'd136314880;
      48562: inst = 32'd268468224;
      48563: inst = 32'd201346511;
      48564: inst = 32'd203483685;
      48565: inst = 32'd471859200;
      48566: inst = 32'd136314880;
      48567: inst = 32'd268468224;
      48568: inst = 32'd201346512;
      48569: inst = 32'd203483685;
      48570: inst = 32'd471859200;
      48571: inst = 32'd136314880;
      48572: inst = 32'd268468224;
      48573: inst = 32'd201346513;
      48574: inst = 32'd203483685;
      48575: inst = 32'd471859200;
      48576: inst = 32'd136314880;
      48577: inst = 32'd268468224;
      48578: inst = 32'd201346514;
      48579: inst = 32'd203483685;
      48580: inst = 32'd471859200;
      48581: inst = 32'd136314880;
      48582: inst = 32'd268468224;
      48583: inst = 32'd201346515;
      48584: inst = 32'd203483685;
      48585: inst = 32'd471859200;
      48586: inst = 32'd136314880;
      48587: inst = 32'd268468224;
      48588: inst = 32'd201346516;
      48589: inst = 32'd203483685;
      48590: inst = 32'd471859200;
      48591: inst = 32'd136314880;
      48592: inst = 32'd268468224;
      48593: inst = 32'd201346517;
      48594: inst = 32'd203423744;
      48595: inst = 32'd471859200;
      48596: inst = 32'd136314880;
      48597: inst = 32'd268468224;
      48598: inst = 32'd201346518;
      48599: inst = 32'd203423744;
      48600: inst = 32'd471859200;
      48601: inst = 32'd136314880;
      48602: inst = 32'd268468224;
      48603: inst = 32'd201346519;
      48604: inst = 32'd203423744;
      48605: inst = 32'd471859200;
      48606: inst = 32'd136314880;
      48607: inst = 32'd268468224;
      48608: inst = 32'd201346520;
      48609: inst = 32'd203423744;
      48610: inst = 32'd471859200;
      48611: inst = 32'd136314880;
      48612: inst = 32'd268468224;
      48613: inst = 32'd201346521;
      48614: inst = 32'd203423744;
      48615: inst = 32'd471859200;
      48616: inst = 32'd136314880;
      48617: inst = 32'd268468224;
      48618: inst = 32'd201346522;
      48619: inst = 32'd203423744;
      48620: inst = 32'd471859200;
      48621: inst = 32'd136314880;
      48622: inst = 32'd268468224;
      48623: inst = 32'd201346523;
      48624: inst = 32'd203423744;
      48625: inst = 32'd471859200;
      48626: inst = 32'd136314880;
      48627: inst = 32'd268468224;
      48628: inst = 32'd201346524;
      48629: inst = 32'd203423744;
      48630: inst = 32'd471859200;
      48631: inst = 32'd136314880;
      48632: inst = 32'd268468224;
      48633: inst = 32'd201346525;
      48634: inst = 32'd203483685;
      48635: inst = 32'd471859200;
      48636: inst = 32'd136314880;
      48637: inst = 32'd268468224;
      48638: inst = 32'd201346526;
      48639: inst = 32'd203483685;
      48640: inst = 32'd471859200;
      48641: inst = 32'd136314880;
      48642: inst = 32'd268468224;
      48643: inst = 32'd201346527;
      48644: inst = 32'd203483685;
      48645: inst = 32'd471859200;
      48646: inst = 32'd136314880;
      48647: inst = 32'd268468224;
      48648: inst = 32'd201346528;
      48649: inst = 32'd203483685;
      48650: inst = 32'd471859200;
      48651: inst = 32'd136314880;
      48652: inst = 32'd268468224;
      48653: inst = 32'd201346529;
      48654: inst = 32'd203483685;
      48655: inst = 32'd471859200;
      48656: inst = 32'd136314880;
      48657: inst = 32'd268468224;
      48658: inst = 32'd201346530;
      48659: inst = 32'd203423744;
      48660: inst = 32'd471859200;
      48661: inst = 32'd136314880;
      48662: inst = 32'd268468224;
      48663: inst = 32'd201346531;
      48664: inst = 32'd203423744;
      48665: inst = 32'd471859200;
      48666: inst = 32'd136314880;
      48667: inst = 32'd268468224;
      48668: inst = 32'd201346532;
      48669: inst = 32'd203423744;
      48670: inst = 32'd471859200;
      48671: inst = 32'd136314880;
      48672: inst = 32'd268468224;
      48673: inst = 32'd201346533;
      48674: inst = 32'd203483685;
      48675: inst = 32'd471859200;
      48676: inst = 32'd136314880;
      48677: inst = 32'd268468224;
      48678: inst = 32'd201346534;
      48679: inst = 32'd203483685;
      48680: inst = 32'd471859200;
      48681: inst = 32'd136314880;
      48682: inst = 32'd268468224;
      48683: inst = 32'd201346535;
      48684: inst = 32'd203483685;
      48685: inst = 32'd471859200;
      48686: inst = 32'd136314880;
      48687: inst = 32'd268468224;
      48688: inst = 32'd201346536;
      48689: inst = 32'd203483685;
      48690: inst = 32'd471859200;
      48691: inst = 32'd136314880;
      48692: inst = 32'd268468224;
      48693: inst = 32'd201346537;
      48694: inst = 32'd203423744;
      48695: inst = 32'd471859200;
      48696: inst = 32'd136314880;
      48697: inst = 32'd268468224;
      48698: inst = 32'd201346538;
      48699: inst = 32'd203423744;
      48700: inst = 32'd471859200;
      48701: inst = 32'd136314880;
      48702: inst = 32'd268468224;
      48703: inst = 32'd201346539;
      48704: inst = 32'd203423744;
      48705: inst = 32'd471859200;
      48706: inst = 32'd136314880;
      48707: inst = 32'd268468224;
      48708: inst = 32'd201346540;
      48709: inst = 32'd203423744;
      48710: inst = 32'd471859200;
      48711: inst = 32'd136314880;
      48712: inst = 32'd268468224;
      48713: inst = 32'd201346541;
      48714: inst = 32'd203423744;
      48715: inst = 32'd471859200;
      48716: inst = 32'd136314880;
      48717: inst = 32'd268468224;
      48718: inst = 32'd201346542;
      48719: inst = 32'd203423744;
      48720: inst = 32'd471859200;
      48721: inst = 32'd136314880;
      48722: inst = 32'd268468224;
      48723: inst = 32'd201346543;
      48724: inst = 32'd203423744;
      48725: inst = 32'd471859200;
      48726: inst = 32'd136314880;
      48727: inst = 32'd268468224;
      48728: inst = 32'd201346544;
      48729: inst = 32'd203423744;
      48730: inst = 32'd471859200;
      48731: inst = 32'd136314880;
      48732: inst = 32'd268468224;
      48733: inst = 32'd201346545;
      48734: inst = 32'd203483685;
      48735: inst = 32'd471859200;
      48736: inst = 32'd136314880;
      48737: inst = 32'd268468224;
      48738: inst = 32'd201346546;
      48739: inst = 32'd203483685;
      48740: inst = 32'd471859200;
      48741: inst = 32'd136314880;
      48742: inst = 32'd268468224;
      48743: inst = 32'd201346547;
      48744: inst = 32'd203483685;
      48745: inst = 32'd471859200;
      48746: inst = 32'd136314880;
      48747: inst = 32'd268468224;
      48748: inst = 32'd201346548;
      48749: inst = 32'd203483685;
      48750: inst = 32'd471859200;
      48751: inst = 32'd136314880;
      48752: inst = 32'd268468224;
      48753: inst = 32'd201346549;
      48754: inst = 32'd203483685;
      48755: inst = 32'd471859200;
      48756: inst = 32'd136314880;
      48757: inst = 32'd268468224;
      48758: inst = 32'd201346550;
      48759: inst = 32'd203483685;
      48760: inst = 32'd471859200;
      48761: inst = 32'd136314880;
      48762: inst = 32'd268468224;
      48763: inst = 32'd201346551;
      48764: inst = 32'd203483685;
      48765: inst = 32'd471859200;
      48766: inst = 32'd136314880;
      48767: inst = 32'd268468224;
      48768: inst = 32'd201346552;
      48769: inst = 32'd203483685;
      48770: inst = 32'd471859200;
      48771: inst = 32'd136314880;
      48772: inst = 32'd268468224;
      48773: inst = 32'd201346553;
      48774: inst = 32'd203483685;
      48775: inst = 32'd471859200;
      48776: inst = 32'd136314880;
      48777: inst = 32'd268468224;
      48778: inst = 32'd201346554;
      48779: inst = 32'd203483685;
      48780: inst = 32'd471859200;
      48781: inst = 32'd136314880;
      48782: inst = 32'd268468224;
      48783: inst = 32'd201346555;
      48784: inst = 32'd203423744;
      48785: inst = 32'd471859200;
      48786: inst = 32'd136314880;
      48787: inst = 32'd268468224;
      48788: inst = 32'd201346556;
      48789: inst = 32'd203423744;
      48790: inst = 32'd471859200;
      48791: inst = 32'd136314880;
      48792: inst = 32'd268468224;
      48793: inst = 32'd201346557;
      48794: inst = 32'd203423744;
      48795: inst = 32'd471859200;
      48796: inst = 32'd136314880;
      48797: inst = 32'd268468224;
      48798: inst = 32'd201346558;
      48799: inst = 32'd203483685;
      48800: inst = 32'd471859200;
      48801: inst = 32'd136314880;
      48802: inst = 32'd268468224;
      48803: inst = 32'd201346559;
      48804: inst = 32'd203483685;
      48805: inst = 32'd471859200;
      48806: inst = 32'd136314880;
      48807: inst = 32'd268468224;
      48808: inst = 32'd201346560;
      48809: inst = 32'd203483685;
      48810: inst = 32'd471859200;
      48811: inst = 32'd136314880;
      48812: inst = 32'd268468224;
      48813: inst = 32'd201346561;
      48814: inst = 32'd203483685;
      48815: inst = 32'd471859200;
      48816: inst = 32'd136314880;
      48817: inst = 32'd268468224;
      48818: inst = 32'd201346562;
      48819: inst = 32'd203483685;
      48820: inst = 32'd471859200;
      48821: inst = 32'd136314880;
      48822: inst = 32'd268468224;
      48823: inst = 32'd201346563;
      48824: inst = 32'd203483685;
      48825: inst = 32'd471859200;
      48826: inst = 32'd136314880;
      48827: inst = 32'd268468224;
      48828: inst = 32'd201346564;
      48829: inst = 32'd203483685;
      48830: inst = 32'd471859200;
      48831: inst = 32'd136314880;
      48832: inst = 32'd268468224;
      48833: inst = 32'd201346565;
      48834: inst = 32'd203483685;
      48835: inst = 32'd471859200;
      48836: inst = 32'd136314880;
      48837: inst = 32'd268468224;
      48838: inst = 32'd201346566;
      48839: inst = 32'd203423744;
      48840: inst = 32'd471859200;
      48841: inst = 32'd136314880;
      48842: inst = 32'd268468224;
      48843: inst = 32'd201346567;
      48844: inst = 32'd203423744;
      48845: inst = 32'd471859200;
      48846: inst = 32'd136314880;
      48847: inst = 32'd268468224;
      48848: inst = 32'd201346568;
      48849: inst = 32'd203423744;
      48850: inst = 32'd471859200;
      48851: inst = 32'd136314880;
      48852: inst = 32'd268468224;
      48853: inst = 32'd201346569;
      48854: inst = 32'd203423744;
      48855: inst = 32'd471859200;
      48856: inst = 32'd136314880;
      48857: inst = 32'd268468224;
      48858: inst = 32'd201346570;
      48859: inst = 32'd203483685;
      48860: inst = 32'd471859200;
      48861: inst = 32'd136314880;
      48862: inst = 32'd268468224;
      48863: inst = 32'd201346571;
      48864: inst = 32'd203483685;
      48865: inst = 32'd471859200;
      48866: inst = 32'd136314880;
      48867: inst = 32'd268468224;
      48868: inst = 32'd201346572;
      48869: inst = 32'd203483685;
      48870: inst = 32'd471859200;
      48871: inst = 32'd136314880;
      48872: inst = 32'd268468224;
      48873: inst = 32'd201346573;
      48874: inst = 32'd203483685;
      48875: inst = 32'd471859200;
      48876: inst = 32'd136314880;
      48877: inst = 32'd268468224;
      48878: inst = 32'd201346574;
      48879: inst = 32'd203483685;
      48880: inst = 32'd471859200;
      48881: inst = 32'd136314880;
      48882: inst = 32'd268468224;
      48883: inst = 32'd201346575;
      48884: inst = 32'd203483685;
      48885: inst = 32'd471859200;
      48886: inst = 32'd136314880;
      48887: inst = 32'd268468224;
      48888: inst = 32'd201346576;
      48889: inst = 32'd203483685;
      48890: inst = 32'd471859200;
      48891: inst = 32'd136314880;
      48892: inst = 32'd268468224;
      48893: inst = 32'd201346577;
      48894: inst = 32'd203483685;
      48895: inst = 32'd471859200;
      48896: inst = 32'd136314880;
      48897: inst = 32'd268468224;
      48898: inst = 32'd201346578;
      48899: inst = 32'd203483685;
      48900: inst = 32'd471859200;
      48901: inst = 32'd136314880;
      48902: inst = 32'd268468224;
      48903: inst = 32'd201346579;
      48904: inst = 32'd203423744;
      48905: inst = 32'd471859200;
      48906: inst = 32'd136314880;
      48907: inst = 32'd268468224;
      48908: inst = 32'd201346580;
      48909: inst = 32'd203423744;
      48910: inst = 32'd471859200;
      48911: inst = 32'd136314880;
      48912: inst = 32'd268468224;
      48913: inst = 32'd201346581;
      48914: inst = 32'd203423744;
      48915: inst = 32'd471859200;
      48916: inst = 32'd136314880;
      48917: inst = 32'd268468224;
      48918: inst = 32'd201346582;
      48919: inst = 32'd203423744;
      48920: inst = 32'd471859200;
      48921: inst = 32'd136314880;
      48922: inst = 32'd268468224;
      48923: inst = 32'd201346583;
      48924: inst = 32'd203423744;
      48925: inst = 32'd471859200;
      48926: inst = 32'd136314880;
      48927: inst = 32'd268468224;
      48928: inst = 32'd201346584;
      48929: inst = 32'd203423744;
      48930: inst = 32'd471859200;
      48931: inst = 32'd136314880;
      48932: inst = 32'd268468224;
      48933: inst = 32'd201346585;
      48934: inst = 32'd203423744;
      48935: inst = 32'd471859200;
      48936: inst = 32'd136314880;
      48937: inst = 32'd268468224;
      48938: inst = 32'd201346586;
      48939: inst = 32'd203423744;
      48940: inst = 32'd471859200;
      48941: inst = 32'd136314880;
      48942: inst = 32'd268468224;
      48943: inst = 32'd201346587;
      48944: inst = 32'd203423744;
      48945: inst = 32'd471859200;
      48946: inst = 32'd136314880;
      48947: inst = 32'd268468224;
      48948: inst = 32'd201346588;
      48949: inst = 32'd203423744;
      48950: inst = 32'd471859200;
      48951: inst = 32'd136314880;
      48952: inst = 32'd268468224;
      48953: inst = 32'd201346589;
      48954: inst = 32'd203423744;
      48955: inst = 32'd471859200;
      48956: inst = 32'd136314880;
      48957: inst = 32'd268468224;
      48958: inst = 32'd201346590;
      48959: inst = 32'd203423744;
      48960: inst = 32'd471859200;
      48961: inst = 32'd136314880;
      48962: inst = 32'd268468224;
      48963: inst = 32'd201346591;
      48964: inst = 32'd203423744;
      48965: inst = 32'd471859200;
      48966: inst = 32'd136314880;
      48967: inst = 32'd268468224;
      48968: inst = 32'd201346592;
      48969: inst = 32'd203423744;
      48970: inst = 32'd471859200;
      48971: inst = 32'd136314880;
      48972: inst = 32'd268468224;
      48973: inst = 32'd201346593;
      48974: inst = 32'd203423744;
      48975: inst = 32'd471859200;
      48976: inst = 32'd136314880;
      48977: inst = 32'd268468224;
      48978: inst = 32'd201346594;
      48979: inst = 32'd203423744;
      48980: inst = 32'd471859200;
      48981: inst = 32'd136314880;
      48982: inst = 32'd268468224;
      48983: inst = 32'd201346595;
      48984: inst = 32'd203423744;
      48985: inst = 32'd471859200;
      48986: inst = 32'd136314880;
      48987: inst = 32'd268468224;
      48988: inst = 32'd201346596;
      48989: inst = 32'd203423744;
      48990: inst = 32'd471859200;
      48991: inst = 32'd136314880;
      48992: inst = 32'd268468224;
      48993: inst = 32'd201346597;
      48994: inst = 32'd203423744;
      48995: inst = 32'd471859200;
      48996: inst = 32'd136314880;
      48997: inst = 32'd268468224;
      48998: inst = 32'd201346598;
      48999: inst = 32'd203423744;
      49000: inst = 32'd471859200;
      49001: inst = 32'd136314880;
      49002: inst = 32'd268468224;
      49003: inst = 32'd201346599;
      49004: inst = 32'd203423744;
      49005: inst = 32'd471859200;
      49006: inst = 32'd136314880;
      49007: inst = 32'd268468224;
      49008: inst = 32'd201346600;
      49009: inst = 32'd203423744;
      49010: inst = 32'd471859200;
      49011: inst = 32'd136314880;
      49012: inst = 32'd268468224;
      49013: inst = 32'd201346601;
      49014: inst = 32'd203423744;
      49015: inst = 32'd471859200;
      49016: inst = 32'd136314880;
      49017: inst = 32'd268468224;
      49018: inst = 32'd201346602;
      49019: inst = 32'd203423744;
      49020: inst = 32'd471859200;
      49021: inst = 32'd136314880;
      49022: inst = 32'd268468224;
      49023: inst = 32'd201346603;
      49024: inst = 32'd203423744;
      49025: inst = 32'd471859200;
      49026: inst = 32'd136314880;
      49027: inst = 32'd268468224;
      49028: inst = 32'd201346604;
      49029: inst = 32'd203423744;
      49030: inst = 32'd471859200;
      49031: inst = 32'd136314880;
      49032: inst = 32'd268468224;
      49033: inst = 32'd201346605;
      49034: inst = 32'd203483685;
      49035: inst = 32'd471859200;
      49036: inst = 32'd136314880;
      49037: inst = 32'd268468224;
      49038: inst = 32'd201346606;
      49039: inst = 32'd203483685;
      49040: inst = 32'd471859200;
      49041: inst = 32'd136314880;
      49042: inst = 32'd268468224;
      49043: inst = 32'd201346607;
      49044: inst = 32'd203483685;
      49045: inst = 32'd471859200;
      49046: inst = 32'd136314880;
      49047: inst = 32'd268468224;
      49048: inst = 32'd201346608;
      49049: inst = 32'd203483685;
      49050: inst = 32'd471859200;
      49051: inst = 32'd136314880;
      49052: inst = 32'd268468224;
      49053: inst = 32'd201346609;
      49054: inst = 32'd203483685;
      49055: inst = 32'd471859200;
      49056: inst = 32'd136314880;
      49057: inst = 32'd268468224;
      49058: inst = 32'd201346610;
      49059: inst = 32'd203483685;
      49060: inst = 32'd471859200;
      49061: inst = 32'd136314880;
      49062: inst = 32'd268468224;
      49063: inst = 32'd201346611;
      49064: inst = 32'd203483685;
      49065: inst = 32'd471859200;
      49066: inst = 32'd136314880;
      49067: inst = 32'd268468224;
      49068: inst = 32'd201346612;
      49069: inst = 32'd203483685;
      49070: inst = 32'd471859200;
      49071: inst = 32'd136314880;
      49072: inst = 32'd268468224;
      49073: inst = 32'd201346613;
      49074: inst = 32'd203423744;
      49075: inst = 32'd471859200;
      49076: inst = 32'd136314880;
      49077: inst = 32'd268468224;
      49078: inst = 32'd201346614;
      49079: inst = 32'd203423744;
      49080: inst = 32'd471859200;
      49081: inst = 32'd136314880;
      49082: inst = 32'd268468224;
      49083: inst = 32'd201346615;
      49084: inst = 32'd203423744;
      49085: inst = 32'd471859200;
      49086: inst = 32'd136314880;
      49087: inst = 32'd268468224;
      49088: inst = 32'd201346616;
      49089: inst = 32'd203423744;
      49090: inst = 32'd471859200;
      49091: inst = 32'd136314880;
      49092: inst = 32'd268468224;
      49093: inst = 32'd201346617;
      49094: inst = 32'd203423744;
      49095: inst = 32'd471859200;
      49096: inst = 32'd136314880;
      49097: inst = 32'd268468224;
      49098: inst = 32'd201346618;
      49099: inst = 32'd203423744;
      49100: inst = 32'd471859200;
      49101: inst = 32'd136314880;
      49102: inst = 32'd268468224;
      49103: inst = 32'd201346619;
      49104: inst = 32'd203423744;
      49105: inst = 32'd471859200;
      49106: inst = 32'd136314880;
      49107: inst = 32'd268468224;
      49108: inst = 32'd201346620;
      49109: inst = 32'd203423744;
      49110: inst = 32'd471859200;
      49111: inst = 32'd136314880;
      49112: inst = 32'd268468224;
      49113: inst = 32'd201346621;
      49114: inst = 32'd203423744;
      49115: inst = 32'd471859200;
      49116: inst = 32'd136314880;
      49117: inst = 32'd268468224;
      49118: inst = 32'd201346622;
      49119: inst = 32'd203483685;
      49120: inst = 32'd471859200;
      49121: inst = 32'd136314880;
      49122: inst = 32'd268468224;
      49123: inst = 32'd201346623;
      49124: inst = 32'd203483685;
      49125: inst = 32'd471859200;
      49126: inst = 32'd136314880;
      49127: inst = 32'd268468224;
      49128: inst = 32'd201346624;
      49129: inst = 32'd203483685;
      49130: inst = 32'd471859200;
      49131: inst = 32'd136314880;
      49132: inst = 32'd268468224;
      49133: inst = 32'd201346625;
      49134: inst = 32'd203483685;
      49135: inst = 32'd471859200;
      49136: inst = 32'd136314880;
      49137: inst = 32'd268468224;
      49138: inst = 32'd201346626;
      49139: inst = 32'd203483685;
      49140: inst = 32'd471859200;
      49141: inst = 32'd136314880;
      49142: inst = 32'd268468224;
      49143: inst = 32'd201346627;
      49144: inst = 32'd203423744;
      49145: inst = 32'd471859200;
      49146: inst = 32'd136314880;
      49147: inst = 32'd268468224;
      49148: inst = 32'd201346628;
      49149: inst = 32'd203423744;
      49150: inst = 32'd471859200;
      49151: inst = 32'd136314880;
      49152: inst = 32'd268468224;
      49153: inst = 32'd201346629;
      49154: inst = 32'd203483685;
      49155: inst = 32'd471859200;
      49156: inst = 32'd136314880;
      49157: inst = 32'd268468224;
      49158: inst = 32'd201346630;
      49159: inst = 32'd203483685;
      49160: inst = 32'd471859200;
      49161: inst = 32'd136314880;
      49162: inst = 32'd268468224;
      49163: inst = 32'd201346631;
      49164: inst = 32'd203483685;
      49165: inst = 32'd471859200;
      49166: inst = 32'd136314880;
      49167: inst = 32'd268468224;
      49168: inst = 32'd201346632;
      49169: inst = 32'd203483685;
      49170: inst = 32'd471859200;
      49171: inst = 32'd136314880;
      49172: inst = 32'd268468224;
      49173: inst = 32'd201346633;
      49174: inst = 32'd203423744;
      49175: inst = 32'd471859200;
      49176: inst = 32'd136314880;
      49177: inst = 32'd268468224;
      49178: inst = 32'd201346634;
      49179: inst = 32'd203423744;
      49180: inst = 32'd471859200;
      49181: inst = 32'd136314880;
      49182: inst = 32'd268468224;
      49183: inst = 32'd201346635;
      49184: inst = 32'd203423744;
      49185: inst = 32'd471859200;
      49186: inst = 32'd136314880;
      49187: inst = 32'd268468224;
      49188: inst = 32'd201346636;
      49189: inst = 32'd203423744;
      49190: inst = 32'd471859200;
      49191: inst = 32'd136314880;
      49192: inst = 32'd268468224;
      49193: inst = 32'd201346637;
      49194: inst = 32'd203423744;
      49195: inst = 32'd471859200;
      49196: inst = 32'd136314880;
      49197: inst = 32'd268468224;
      49198: inst = 32'd201346638;
      49199: inst = 32'd203423744;
      49200: inst = 32'd471859200;
      49201: inst = 32'd136314880;
      49202: inst = 32'd268468224;
      49203: inst = 32'd201346639;
      49204: inst = 32'd203423744;
      49205: inst = 32'd471859200;
      49206: inst = 32'd136314880;
      49207: inst = 32'd268468224;
      49208: inst = 32'd201346640;
      49209: inst = 32'd203423744;
      49210: inst = 32'd471859200;
      49211: inst = 32'd136314880;
      49212: inst = 32'd268468224;
      49213: inst = 32'd201346641;
      49214: inst = 32'd203483685;
      49215: inst = 32'd471859200;
      49216: inst = 32'd136314880;
      49217: inst = 32'd268468224;
      49218: inst = 32'd201346642;
      49219: inst = 32'd203483685;
      49220: inst = 32'd471859200;
      49221: inst = 32'd136314880;
      49222: inst = 32'd268468224;
      49223: inst = 32'd201346643;
      49224: inst = 32'd203483685;
      49225: inst = 32'd471859200;
      49226: inst = 32'd136314880;
      49227: inst = 32'd268468224;
      49228: inst = 32'd201346644;
      49229: inst = 32'd203483685;
      49230: inst = 32'd471859200;
      49231: inst = 32'd136314880;
      49232: inst = 32'd268468224;
      49233: inst = 32'd201346645;
      49234: inst = 32'd203483685;
      49235: inst = 32'd471859200;
      49236: inst = 32'd136314880;
      49237: inst = 32'd268468224;
      49238: inst = 32'd201346646;
      49239: inst = 32'd203483685;
      49240: inst = 32'd471859200;
      49241: inst = 32'd136314880;
      49242: inst = 32'd268468224;
      49243: inst = 32'd201346647;
      49244: inst = 32'd203483685;
      49245: inst = 32'd471859200;
      49246: inst = 32'd136314880;
      49247: inst = 32'd268468224;
      49248: inst = 32'd201346648;
      49249: inst = 32'd203483685;
      49250: inst = 32'd471859200;
      49251: inst = 32'd136314880;
      49252: inst = 32'd268468224;
      49253: inst = 32'd201346649;
      49254: inst = 32'd203483685;
      49255: inst = 32'd471859200;
      49256: inst = 32'd136314880;
      49257: inst = 32'd268468224;
      49258: inst = 32'd201346650;
      49259: inst = 32'd203483685;
      49260: inst = 32'd471859200;
      49261: inst = 32'd136314880;
      49262: inst = 32'd268468224;
      49263: inst = 32'd201346651;
      49264: inst = 32'd203483685;
      49265: inst = 32'd471859200;
      49266: inst = 32'd136314880;
      49267: inst = 32'd268468224;
      49268: inst = 32'd201346652;
      49269: inst = 32'd203423744;
      49270: inst = 32'd471859200;
      49271: inst = 32'd136314880;
      49272: inst = 32'd268468224;
      49273: inst = 32'd201346653;
      49274: inst = 32'd203423744;
      49275: inst = 32'd471859200;
      49276: inst = 32'd136314880;
      49277: inst = 32'd268468224;
      49278: inst = 32'd201346654;
      49279: inst = 32'd203483685;
      49280: inst = 32'd471859200;
      49281: inst = 32'd136314880;
      49282: inst = 32'd268468224;
      49283: inst = 32'd201346655;
      49284: inst = 32'd203483685;
      49285: inst = 32'd471859200;
      49286: inst = 32'd136314880;
      49287: inst = 32'd268468224;
      49288: inst = 32'd201346656;
      49289: inst = 32'd203483685;
      49290: inst = 32'd471859200;
      49291: inst = 32'd136314880;
      49292: inst = 32'd268468224;
      49293: inst = 32'd201346657;
      49294: inst = 32'd203483685;
      49295: inst = 32'd471859200;
      49296: inst = 32'd136314880;
      49297: inst = 32'd268468224;
      49298: inst = 32'd201346658;
      49299: inst = 32'd203483685;
      49300: inst = 32'd471859200;
      49301: inst = 32'd136314880;
      49302: inst = 32'd268468224;
      49303: inst = 32'd201346659;
      49304: inst = 32'd203483685;
      49305: inst = 32'd471859200;
      49306: inst = 32'd136314880;
      49307: inst = 32'd268468224;
      49308: inst = 32'd201346660;
      49309: inst = 32'd203483685;
      49310: inst = 32'd471859200;
      49311: inst = 32'd136314880;
      49312: inst = 32'd268468224;
      49313: inst = 32'd201346661;
      49314: inst = 32'd203483685;
      49315: inst = 32'd471859200;
      49316: inst = 32'd136314880;
      49317: inst = 32'd268468224;
      49318: inst = 32'd201346662;
      49319: inst = 32'd203423744;
      49320: inst = 32'd471859200;
      49321: inst = 32'd136314880;
      49322: inst = 32'd268468224;
      49323: inst = 32'd201346663;
      49324: inst = 32'd203423744;
      49325: inst = 32'd471859200;
      49326: inst = 32'd136314880;
      49327: inst = 32'd268468224;
      49328: inst = 32'd201346664;
      49329: inst = 32'd203423744;
      49330: inst = 32'd471859200;
      49331: inst = 32'd136314880;
      49332: inst = 32'd268468224;
      49333: inst = 32'd201346665;
      49334: inst = 32'd203423744;
      49335: inst = 32'd471859200;
      49336: inst = 32'd136314880;
      49337: inst = 32'd268468224;
      49338: inst = 32'd201346666;
      49339: inst = 32'd203483685;
      49340: inst = 32'd471859200;
      49341: inst = 32'd136314880;
      49342: inst = 32'd268468224;
      49343: inst = 32'd201346667;
      49344: inst = 32'd203483685;
      49345: inst = 32'd471859200;
      49346: inst = 32'd136314880;
      49347: inst = 32'd268468224;
      49348: inst = 32'd201346668;
      49349: inst = 32'd203483685;
      49350: inst = 32'd471859200;
      49351: inst = 32'd136314880;
      49352: inst = 32'd268468224;
      49353: inst = 32'd201346669;
      49354: inst = 32'd203483685;
      49355: inst = 32'd471859200;
      49356: inst = 32'd136314880;
      49357: inst = 32'd268468224;
      49358: inst = 32'd201346670;
      49359: inst = 32'd203483685;
      49360: inst = 32'd471859200;
      49361: inst = 32'd136314880;
      49362: inst = 32'd268468224;
      49363: inst = 32'd201346671;
      49364: inst = 32'd203483685;
      49365: inst = 32'd471859200;
      49366: inst = 32'd136314880;
      49367: inst = 32'd268468224;
      49368: inst = 32'd201346672;
      49369: inst = 32'd203483685;
      49370: inst = 32'd471859200;
      49371: inst = 32'd136314880;
      49372: inst = 32'd268468224;
      49373: inst = 32'd201346673;
      49374: inst = 32'd203483685;
      49375: inst = 32'd471859200;
      49376: inst = 32'd136314880;
      49377: inst = 32'd268468224;
      49378: inst = 32'd201346674;
      49379: inst = 32'd203483685;
      49380: inst = 32'd471859200;
      49381: inst = 32'd136314880;
      49382: inst = 32'd268468224;
      49383: inst = 32'd201346675;
      49384: inst = 32'd203423744;
      49385: inst = 32'd471859200;
      49386: inst = 32'd136314880;
      49387: inst = 32'd268468224;
      49388: inst = 32'd201346676;
      49389: inst = 32'd203423744;
      49390: inst = 32'd471859200;
      49391: inst = 32'd136314880;
      49392: inst = 32'd268468224;
      49393: inst = 32'd201346677;
      49394: inst = 32'd203423744;
      49395: inst = 32'd471859200;
      49396: inst = 32'd136314880;
      49397: inst = 32'd268468224;
      49398: inst = 32'd201346678;
      49399: inst = 32'd203423744;
      49400: inst = 32'd471859200;
      49401: inst = 32'd136314880;
      49402: inst = 32'd268468224;
      49403: inst = 32'd201346679;
      49404: inst = 32'd203423744;
      49405: inst = 32'd471859200;
      49406: inst = 32'd136314880;
      49407: inst = 32'd268468224;
      49408: inst = 32'd201346680;
      49409: inst = 32'd203423744;
      49410: inst = 32'd471859200;
      49411: inst = 32'd136314880;
      49412: inst = 32'd268468224;
      49413: inst = 32'd201346681;
      49414: inst = 32'd203423744;
      49415: inst = 32'd471859200;
      49416: inst = 32'd136314880;
      49417: inst = 32'd268468224;
      49418: inst = 32'd201346682;
      49419: inst = 32'd203423744;
      49420: inst = 32'd471859200;
      49421: inst = 32'd136314880;
      49422: inst = 32'd268468224;
      49423: inst = 32'd201346683;
      49424: inst = 32'd203423744;
      49425: inst = 32'd471859200;
      49426: inst = 32'd136314880;
      49427: inst = 32'd268468224;
      49428: inst = 32'd201346684;
      49429: inst = 32'd203423744;
      49430: inst = 32'd471859200;
      49431: inst = 32'd136314880;
      49432: inst = 32'd268468224;
      49433: inst = 32'd201346685;
      49434: inst = 32'd203423744;
      49435: inst = 32'd471859200;
      49436: inst = 32'd136314880;
      49437: inst = 32'd268468224;
      49438: inst = 32'd201346686;
      49439: inst = 32'd203423744;
      49440: inst = 32'd471859200;
      49441: inst = 32'd136314880;
      49442: inst = 32'd268468224;
      49443: inst = 32'd201346687;
      49444: inst = 32'd203423744;
      49445: inst = 32'd471859200;
      49446: inst = 32'd136314880;
      49447: inst = 32'd268468224;
      49448: inst = 32'd201346688;
      49449: inst = 32'd203423744;
      49450: inst = 32'd471859200;
      49451: inst = 32'd136314880;
      49452: inst = 32'd268468224;
      49453: inst = 32'd201346689;
      49454: inst = 32'd203423744;
      49455: inst = 32'd471859200;
      49456: inst = 32'd136314880;
      49457: inst = 32'd268468224;
      49458: inst = 32'd201346690;
      49459: inst = 32'd203423744;
      49460: inst = 32'd471859200;
      49461: inst = 32'd136314880;
      49462: inst = 32'd268468224;
      49463: inst = 32'd201346691;
      49464: inst = 32'd203423744;
      49465: inst = 32'd471859200;
      49466: inst = 32'd136314880;
      49467: inst = 32'd268468224;
      49468: inst = 32'd201346692;
      49469: inst = 32'd203423744;
      49470: inst = 32'd471859200;
      49471: inst = 32'd136314880;
      49472: inst = 32'd268468224;
      49473: inst = 32'd201346693;
      49474: inst = 32'd203423744;
      49475: inst = 32'd471859200;
      49476: inst = 32'd136314880;
      49477: inst = 32'd268468224;
      49478: inst = 32'd201346694;
      49479: inst = 32'd203423744;
      49480: inst = 32'd471859200;
      49481: inst = 32'd136314880;
      49482: inst = 32'd268468224;
      49483: inst = 32'd201346695;
      49484: inst = 32'd203423744;
      49485: inst = 32'd471859200;
      49486: inst = 32'd136314880;
      49487: inst = 32'd268468224;
      49488: inst = 32'd201346696;
      49489: inst = 32'd203423744;
      49490: inst = 32'd471859200;
      49491: inst = 32'd136314880;
      49492: inst = 32'd268468224;
      49493: inst = 32'd201346697;
      49494: inst = 32'd203423744;
      49495: inst = 32'd471859200;
      49496: inst = 32'd136314880;
      49497: inst = 32'd268468224;
      49498: inst = 32'd201346698;
      49499: inst = 32'd203423744;
      49500: inst = 32'd471859200;
      49501: inst = 32'd136314880;
      49502: inst = 32'd268468224;
      49503: inst = 32'd201346699;
      49504: inst = 32'd203423744;
      49505: inst = 32'd471859200;
      49506: inst = 32'd136314880;
      49507: inst = 32'd268468224;
      49508: inst = 32'd201346700;
      49509: inst = 32'd203423744;
      49510: inst = 32'd471859200;
      49511: inst = 32'd136314880;
      49512: inst = 32'd268468224;
      49513: inst = 32'd201346701;
      49514: inst = 32'd203483685;
      49515: inst = 32'd471859200;
      49516: inst = 32'd136314880;
      49517: inst = 32'd268468224;
      49518: inst = 32'd201346702;
      49519: inst = 32'd203483685;
      49520: inst = 32'd471859200;
      49521: inst = 32'd136314880;
      49522: inst = 32'd268468224;
      49523: inst = 32'd201346703;
      49524: inst = 32'd203483685;
      49525: inst = 32'd471859200;
      49526: inst = 32'd136314880;
      49527: inst = 32'd268468224;
      49528: inst = 32'd201346704;
      49529: inst = 32'd203483685;
      49530: inst = 32'd471859200;
      49531: inst = 32'd136314880;
      49532: inst = 32'd268468224;
      49533: inst = 32'd201346705;
      49534: inst = 32'd203483685;
      49535: inst = 32'd471859200;
      49536: inst = 32'd136314880;
      49537: inst = 32'd268468224;
      49538: inst = 32'd201346706;
      49539: inst = 32'd203483685;
      49540: inst = 32'd471859200;
      49541: inst = 32'd136314880;
      49542: inst = 32'd268468224;
      49543: inst = 32'd201346707;
      49544: inst = 32'd203483685;
      49545: inst = 32'd471859200;
      49546: inst = 32'd136314880;
      49547: inst = 32'd268468224;
      49548: inst = 32'd201346708;
      49549: inst = 32'd203483685;
      49550: inst = 32'd471859200;
      49551: inst = 32'd136314880;
      49552: inst = 32'd268468224;
      49553: inst = 32'd201346709;
      49554: inst = 32'd203483685;
      49555: inst = 32'd471859200;
      49556: inst = 32'd136314880;
      49557: inst = 32'd268468224;
      49558: inst = 32'd201346710;
      49559: inst = 32'd203483685;
      49560: inst = 32'd471859200;
      49561: inst = 32'd136314880;
      49562: inst = 32'd268468224;
      49563: inst = 32'd201346711;
      49564: inst = 32'd203483685;
      49565: inst = 32'd471859200;
      49566: inst = 32'd136314880;
      49567: inst = 32'd268468224;
      49568: inst = 32'd201346712;
      49569: inst = 32'd203483685;
      49570: inst = 32'd471859200;
      49571: inst = 32'd136314880;
      49572: inst = 32'd268468224;
      49573: inst = 32'd201346713;
      49574: inst = 32'd203483685;
      49575: inst = 32'd471859200;
      49576: inst = 32'd136314880;
      49577: inst = 32'd268468224;
      49578: inst = 32'd201346714;
      49579: inst = 32'd203483685;
      49580: inst = 32'd471859200;
      49581: inst = 32'd136314880;
      49582: inst = 32'd268468224;
      49583: inst = 32'd201346715;
      49584: inst = 32'd203483685;
      49585: inst = 32'd471859200;
      49586: inst = 32'd136314880;
      49587: inst = 32'd268468224;
      49588: inst = 32'd201346716;
      49589: inst = 32'd203483685;
      49590: inst = 32'd471859200;
      49591: inst = 32'd136314880;
      49592: inst = 32'd268468224;
      49593: inst = 32'd201346717;
      49594: inst = 32'd203483685;
      49595: inst = 32'd471859200;
      49596: inst = 32'd136314880;
      49597: inst = 32'd268468224;
      49598: inst = 32'd201346718;
      49599: inst = 32'd203483685;
      49600: inst = 32'd471859200;
      49601: inst = 32'd136314880;
      49602: inst = 32'd268468224;
      49603: inst = 32'd201346719;
      49604: inst = 32'd203483685;
      49605: inst = 32'd471859200;
      49606: inst = 32'd136314880;
      49607: inst = 32'd268468224;
      49608: inst = 32'd201346720;
      49609: inst = 32'd203483685;
      49610: inst = 32'd471859200;
      49611: inst = 32'd136314880;
      49612: inst = 32'd268468224;
      49613: inst = 32'd201346721;
      49614: inst = 32'd203483685;
      49615: inst = 32'd471859200;
      49616: inst = 32'd136314880;
      49617: inst = 32'd268468224;
      49618: inst = 32'd201346722;
      49619: inst = 32'd203483685;
      49620: inst = 32'd471859200;
      49621: inst = 32'd136314880;
      49622: inst = 32'd268468224;
      49623: inst = 32'd201346723;
      49624: inst = 32'd203483685;
      49625: inst = 32'd471859200;
      49626: inst = 32'd136314880;
      49627: inst = 32'd268468224;
      49628: inst = 32'd201346724;
      49629: inst = 32'd203423744;
      49630: inst = 32'd471859200;
      49631: inst = 32'd136314880;
      49632: inst = 32'd268468224;
      49633: inst = 32'd201346725;
      49634: inst = 32'd203483685;
      49635: inst = 32'd471859200;
      49636: inst = 32'd136314880;
      49637: inst = 32'd268468224;
      49638: inst = 32'd201346726;
      49639: inst = 32'd203483685;
      49640: inst = 32'd471859200;
      49641: inst = 32'd136314880;
      49642: inst = 32'd268468224;
      49643: inst = 32'd201346727;
      49644: inst = 32'd203483685;
      49645: inst = 32'd471859200;
      49646: inst = 32'd136314880;
      49647: inst = 32'd268468224;
      49648: inst = 32'd201346728;
      49649: inst = 32'd203483685;
      49650: inst = 32'd471859200;
      49651: inst = 32'd136314880;
      49652: inst = 32'd268468224;
      49653: inst = 32'd201346729;
      49654: inst = 32'd203483685;
      49655: inst = 32'd471859200;
      49656: inst = 32'd136314880;
      49657: inst = 32'd268468224;
      49658: inst = 32'd201346730;
      49659: inst = 32'd203483685;
      49660: inst = 32'd471859200;
      49661: inst = 32'd136314880;
      49662: inst = 32'd268468224;
      49663: inst = 32'd201346731;
      49664: inst = 32'd203483685;
      49665: inst = 32'd471859200;
      49666: inst = 32'd136314880;
      49667: inst = 32'd268468224;
      49668: inst = 32'd201346732;
      49669: inst = 32'd203483685;
      49670: inst = 32'd471859200;
      49671: inst = 32'd136314880;
      49672: inst = 32'd268468224;
      49673: inst = 32'd201346733;
      49674: inst = 32'd203483685;
      49675: inst = 32'd471859200;
      49676: inst = 32'd136314880;
      49677: inst = 32'd268468224;
      49678: inst = 32'd201346734;
      49679: inst = 32'd203483685;
      49680: inst = 32'd471859200;
      49681: inst = 32'd136314880;
      49682: inst = 32'd268468224;
      49683: inst = 32'd201346735;
      49684: inst = 32'd203483685;
      49685: inst = 32'd471859200;
      49686: inst = 32'd136314880;
      49687: inst = 32'd268468224;
      49688: inst = 32'd201346736;
      49689: inst = 32'd203483685;
      49690: inst = 32'd471859200;
      49691: inst = 32'd136314880;
      49692: inst = 32'd268468224;
      49693: inst = 32'd201346737;
      49694: inst = 32'd203483685;
      49695: inst = 32'd471859200;
      49696: inst = 32'd136314880;
      49697: inst = 32'd268468224;
      49698: inst = 32'd201346738;
      49699: inst = 32'd203483685;
      49700: inst = 32'd471859200;
      49701: inst = 32'd136314880;
      49702: inst = 32'd268468224;
      49703: inst = 32'd201346739;
      49704: inst = 32'd203483685;
      49705: inst = 32'd471859200;
      49706: inst = 32'd136314880;
      49707: inst = 32'd268468224;
      49708: inst = 32'd201346740;
      49709: inst = 32'd203483685;
      49710: inst = 32'd471859200;
      49711: inst = 32'd136314880;
      49712: inst = 32'd268468224;
      49713: inst = 32'd201346741;
      49714: inst = 32'd203483685;
      49715: inst = 32'd471859200;
      49716: inst = 32'd136314880;
      49717: inst = 32'd268468224;
      49718: inst = 32'd201346742;
      49719: inst = 32'd203483685;
      49720: inst = 32'd471859200;
      49721: inst = 32'd136314880;
      49722: inst = 32'd268468224;
      49723: inst = 32'd201346743;
      49724: inst = 32'd203483685;
      49725: inst = 32'd471859200;
      49726: inst = 32'd136314880;
      49727: inst = 32'd268468224;
      49728: inst = 32'd201346744;
      49729: inst = 32'd203483685;
      49730: inst = 32'd471859200;
      49731: inst = 32'd136314880;
      49732: inst = 32'd268468224;
      49733: inst = 32'd201346745;
      49734: inst = 32'd203483685;
      49735: inst = 32'd471859200;
      49736: inst = 32'd136314880;
      49737: inst = 32'd268468224;
      49738: inst = 32'd201346746;
      49739: inst = 32'd203483685;
      49740: inst = 32'd471859200;
      49741: inst = 32'd136314880;
      49742: inst = 32'd268468224;
      49743: inst = 32'd201346747;
      49744: inst = 32'd203483685;
      49745: inst = 32'd471859200;
      49746: inst = 32'd136314880;
      49747: inst = 32'd268468224;
      49748: inst = 32'd201346748;
      49749: inst = 32'd203483685;
      49750: inst = 32'd471859200;
      49751: inst = 32'd136314880;
      49752: inst = 32'd268468224;
      49753: inst = 32'd201346749;
      49754: inst = 32'd203423744;
      49755: inst = 32'd471859200;
      49756: inst = 32'd136314880;
      49757: inst = 32'd268468224;
      49758: inst = 32'd201346750;
      49759: inst = 32'd203483685;
      49760: inst = 32'd471859200;
      49761: inst = 32'd136314880;
      49762: inst = 32'd268468224;
      49763: inst = 32'd201346751;
      49764: inst = 32'd203483685;
      49765: inst = 32'd471859200;
      49766: inst = 32'd136314880;
      49767: inst = 32'd268468224;
      49768: inst = 32'd201346752;
      49769: inst = 32'd203483685;
      49770: inst = 32'd471859200;
      49771: inst = 32'd136314880;
      49772: inst = 32'd268468224;
      49773: inst = 32'd201346753;
      49774: inst = 32'd203423744;
      49775: inst = 32'd471859200;
      49776: inst = 32'd136314880;
      49777: inst = 32'd268468224;
      49778: inst = 32'd201346754;
      49779: inst = 32'd203423744;
      49780: inst = 32'd471859200;
      49781: inst = 32'd136314880;
      49782: inst = 32'd268468224;
      49783: inst = 32'd201346755;
      49784: inst = 32'd203423744;
      49785: inst = 32'd471859200;
      49786: inst = 32'd136314880;
      49787: inst = 32'd268468224;
      49788: inst = 32'd201346756;
      49789: inst = 32'd203423744;
      49790: inst = 32'd471859200;
      49791: inst = 32'd136314880;
      49792: inst = 32'd268468224;
      49793: inst = 32'd201346757;
      49794: inst = 32'd203423744;
      49795: inst = 32'd471859200;
      49796: inst = 32'd136314880;
      49797: inst = 32'd268468224;
      49798: inst = 32'd201346758;
      49799: inst = 32'd203423744;
      49800: inst = 32'd471859200;
      49801: inst = 32'd136314880;
      49802: inst = 32'd268468224;
      49803: inst = 32'd201346759;
      49804: inst = 32'd203423744;
      49805: inst = 32'd471859200;
      49806: inst = 32'd136314880;
      49807: inst = 32'd268468224;
      49808: inst = 32'd201346760;
      49809: inst = 32'd203423744;
      49810: inst = 32'd471859200;
      49811: inst = 32'd136314880;
      49812: inst = 32'd268468224;
      49813: inst = 32'd201346761;
      49814: inst = 32'd203423744;
      49815: inst = 32'd471859200;
      49816: inst = 32'd136314880;
      49817: inst = 32'd268468224;
      49818: inst = 32'd201346762;
      49819: inst = 32'd203483685;
      49820: inst = 32'd471859200;
      49821: inst = 32'd136314880;
      49822: inst = 32'd268468224;
      49823: inst = 32'd201346763;
      49824: inst = 32'd203483685;
      49825: inst = 32'd471859200;
      49826: inst = 32'd136314880;
      49827: inst = 32'd268468224;
      49828: inst = 32'd201346764;
      49829: inst = 32'd203483685;
      49830: inst = 32'd471859200;
      49831: inst = 32'd136314880;
      49832: inst = 32'd268468224;
      49833: inst = 32'd201346765;
      49834: inst = 32'd203483685;
      49835: inst = 32'd471859200;
      49836: inst = 32'd136314880;
      49837: inst = 32'd268468224;
      49838: inst = 32'd201346766;
      49839: inst = 32'd203483685;
      49840: inst = 32'd471859200;
      49841: inst = 32'd136314880;
      49842: inst = 32'd268468224;
      49843: inst = 32'd201346767;
      49844: inst = 32'd203483685;
      49845: inst = 32'd471859200;
      49846: inst = 32'd136314880;
      49847: inst = 32'd268468224;
      49848: inst = 32'd201346768;
      49849: inst = 32'd203483685;
      49850: inst = 32'd471859200;
      49851: inst = 32'd136314880;
      49852: inst = 32'd268468224;
      49853: inst = 32'd201346769;
      49854: inst = 32'd203483685;
      49855: inst = 32'd471859200;
      49856: inst = 32'd136314880;
      49857: inst = 32'd268468224;
      49858: inst = 32'd201346770;
      49859: inst = 32'd203483685;
      49860: inst = 32'd471859200;
      49861: inst = 32'd136314880;
      49862: inst = 32'd268468224;
      49863: inst = 32'd201346771;
      49864: inst = 32'd203483685;
      49865: inst = 32'd471859200;
      49866: inst = 32'd136314880;
      49867: inst = 32'd268468224;
      49868: inst = 32'd201346772;
      49869: inst = 32'd203483685;
      49870: inst = 32'd471859200;
      49871: inst = 32'd136314880;
      49872: inst = 32'd268468224;
      49873: inst = 32'd201346773;
      49874: inst = 32'd203483685;
      49875: inst = 32'd471859200;
      49876: inst = 32'd136314880;
      49877: inst = 32'd268468224;
      49878: inst = 32'd201346774;
      49879: inst = 32'd203423744;
      49880: inst = 32'd471859200;
      49881: inst = 32'd136314880;
      49882: inst = 32'd268468224;
      49883: inst = 32'd201346775;
      49884: inst = 32'd203423744;
      49885: inst = 32'd471859200;
      49886: inst = 32'd136314880;
      49887: inst = 32'd268468224;
      49888: inst = 32'd201346776;
      49889: inst = 32'd203423744;
      49890: inst = 32'd471859200;
      49891: inst = 32'd136314880;
      49892: inst = 32'd268468224;
      49893: inst = 32'd201346777;
      49894: inst = 32'd203423744;
      49895: inst = 32'd471859200;
      49896: inst = 32'd136314880;
      49897: inst = 32'd268468224;
      49898: inst = 32'd201346778;
      49899: inst = 32'd203423744;
      49900: inst = 32'd471859200;
      49901: inst = 32'd136314880;
      49902: inst = 32'd268468224;
      49903: inst = 32'd201346779;
      49904: inst = 32'd203423744;
      49905: inst = 32'd471859200;
      49906: inst = 32'd136314880;
      49907: inst = 32'd268468224;
      49908: inst = 32'd201346780;
      49909: inst = 32'd203423744;
      49910: inst = 32'd471859200;
      49911: inst = 32'd136314880;
      49912: inst = 32'd268468224;
      49913: inst = 32'd201346781;
      49914: inst = 32'd203423744;
      49915: inst = 32'd471859200;
      49916: inst = 32'd136314880;
      49917: inst = 32'd268468224;
      49918: inst = 32'd201346782;
      49919: inst = 32'd203423744;
      49920: inst = 32'd471859200;
      49921: inst = 32'd136314880;
      49922: inst = 32'd268468224;
      49923: inst = 32'd201346783;
      49924: inst = 32'd203423744;
      49925: inst = 32'd471859200;
      49926: inst = 32'd136314880;
      49927: inst = 32'd268468224;
      49928: inst = 32'd201346784;
      49929: inst = 32'd203423744;
      49930: inst = 32'd471859200;
      49931: inst = 32'd136314880;
      49932: inst = 32'd268468224;
      49933: inst = 32'd201346785;
      49934: inst = 32'd203423744;
      49935: inst = 32'd471859200;
      49936: inst = 32'd136314880;
      49937: inst = 32'd268468224;
      49938: inst = 32'd201346786;
      49939: inst = 32'd203423744;
      49940: inst = 32'd471859200;
      49941: inst = 32'd136314880;
      49942: inst = 32'd268468224;
      49943: inst = 32'd201346787;
      49944: inst = 32'd203423744;
      49945: inst = 32'd471859200;
      49946: inst = 32'd136314880;
      49947: inst = 32'd268468224;
      49948: inst = 32'd201346788;
      49949: inst = 32'd203423744;
      49950: inst = 32'd471859200;
      49951: inst = 32'd136314880;
      49952: inst = 32'd268468224;
      49953: inst = 32'd201346789;
      49954: inst = 32'd203423744;
      49955: inst = 32'd471859200;
      49956: inst = 32'd136314880;
      49957: inst = 32'd268468224;
      49958: inst = 32'd201346790;
      49959: inst = 32'd203423744;
      49960: inst = 32'd471859200;
      49961: inst = 32'd136314880;
      49962: inst = 32'd268468224;
      49963: inst = 32'd201346791;
      49964: inst = 32'd203423744;
      49965: inst = 32'd471859200;
      49966: inst = 32'd136314880;
      49967: inst = 32'd268468224;
      49968: inst = 32'd201346792;
      49969: inst = 32'd203423744;
      49970: inst = 32'd471859200;
      49971: inst = 32'd136314880;
      49972: inst = 32'd268468224;
      49973: inst = 32'd201346793;
      49974: inst = 32'd203423744;
      49975: inst = 32'd471859200;
      49976: inst = 32'd136314880;
      49977: inst = 32'd268468224;
      49978: inst = 32'd201346794;
      49979: inst = 32'd203423744;
      49980: inst = 32'd471859200;
      49981: inst = 32'd136314880;
      49982: inst = 32'd268468224;
      49983: inst = 32'd201346795;
      49984: inst = 32'd203423744;
      49985: inst = 32'd471859200;
      49986: inst = 32'd136314880;
      49987: inst = 32'd268468224;
      49988: inst = 32'd201346796;
      49989: inst = 32'd203423744;
      49990: inst = 32'd471859200;
      49991: inst = 32'd136314880;
      49992: inst = 32'd268468224;
      49993: inst = 32'd201346797;
      49994: inst = 32'd203483685;
      49995: inst = 32'd471859200;
      49996: inst = 32'd136314880;
      49997: inst = 32'd268468224;
      49998: inst = 32'd201346798;
      49999: inst = 32'd203483685;
      50000: inst = 32'd471859200;
      50001: inst = 32'd136314880;
      50002: inst = 32'd268468224;
      50003: inst = 32'd201346799;
      50004: inst = 32'd203483685;
      50005: inst = 32'd471859200;
      50006: inst = 32'd136314880;
      50007: inst = 32'd268468224;
      50008: inst = 32'd201346800;
      50009: inst = 32'd203483685;
      50010: inst = 32'd471859200;
      50011: inst = 32'd136314880;
      50012: inst = 32'd268468224;
      50013: inst = 32'd201346801;
      50014: inst = 32'd203483685;
      50015: inst = 32'd471859200;
      50016: inst = 32'd136314880;
      50017: inst = 32'd268468224;
      50018: inst = 32'd201346802;
      50019: inst = 32'd203483685;
      50020: inst = 32'd471859200;
      50021: inst = 32'd136314880;
      50022: inst = 32'd268468224;
      50023: inst = 32'd201346803;
      50024: inst = 32'd203483685;
      50025: inst = 32'd471859200;
      50026: inst = 32'd136314880;
      50027: inst = 32'd268468224;
      50028: inst = 32'd201346804;
      50029: inst = 32'd203483685;
      50030: inst = 32'd471859200;
      50031: inst = 32'd136314880;
      50032: inst = 32'd268468224;
      50033: inst = 32'd201346805;
      50034: inst = 32'd203483685;
      50035: inst = 32'd471859200;
      50036: inst = 32'd136314880;
      50037: inst = 32'd268468224;
      50038: inst = 32'd201346806;
      50039: inst = 32'd203483685;
      50040: inst = 32'd471859200;
      50041: inst = 32'd136314880;
      50042: inst = 32'd268468224;
      50043: inst = 32'd201346807;
      50044: inst = 32'd203483685;
      50045: inst = 32'd471859200;
      50046: inst = 32'd136314880;
      50047: inst = 32'd268468224;
      50048: inst = 32'd201346808;
      50049: inst = 32'd203483685;
      50050: inst = 32'd471859200;
      50051: inst = 32'd136314880;
      50052: inst = 32'd268468224;
      50053: inst = 32'd201346809;
      50054: inst = 32'd203483685;
      50055: inst = 32'd471859200;
      50056: inst = 32'd136314880;
      50057: inst = 32'd268468224;
      50058: inst = 32'd201346810;
      50059: inst = 32'd203483685;
      50060: inst = 32'd471859200;
      50061: inst = 32'd136314880;
      50062: inst = 32'd268468224;
      50063: inst = 32'd201346811;
      50064: inst = 32'd203483685;
      50065: inst = 32'd471859200;
      50066: inst = 32'd136314880;
      50067: inst = 32'd268468224;
      50068: inst = 32'd201346812;
      50069: inst = 32'd203483685;
      50070: inst = 32'd471859200;
      50071: inst = 32'd136314880;
      50072: inst = 32'd268468224;
      50073: inst = 32'd201346813;
      50074: inst = 32'd203483685;
      50075: inst = 32'd471859200;
      50076: inst = 32'd136314880;
      50077: inst = 32'd268468224;
      50078: inst = 32'd201346814;
      50079: inst = 32'd203483685;
      50080: inst = 32'd471859200;
      50081: inst = 32'd136314880;
      50082: inst = 32'd268468224;
      50083: inst = 32'd201346815;
      50084: inst = 32'd203483685;
      50085: inst = 32'd471859200;
      50086: inst = 32'd136314880;
      50087: inst = 32'd268468224;
      50088: inst = 32'd201346816;
      50089: inst = 32'd203483685;
      50090: inst = 32'd471859200;
      50091: inst = 32'd136314880;
      50092: inst = 32'd268468224;
      50093: inst = 32'd201346817;
      50094: inst = 32'd203483685;
      50095: inst = 32'd471859200;
      50096: inst = 32'd136314880;
      50097: inst = 32'd268468224;
      50098: inst = 32'd201346818;
      50099: inst = 32'd203483685;
      50100: inst = 32'd471859200;
      50101: inst = 32'd136314880;
      50102: inst = 32'd268468224;
      50103: inst = 32'd201346819;
      50104: inst = 32'd203483685;
      50105: inst = 32'd471859200;
      50106: inst = 32'd136314880;
      50107: inst = 32'd268468224;
      50108: inst = 32'd201346820;
      50109: inst = 32'd203483685;
      50110: inst = 32'd471859200;
      50111: inst = 32'd136314880;
      50112: inst = 32'd268468224;
      50113: inst = 32'd201346821;
      50114: inst = 32'd203423744;
      50115: inst = 32'd471859200;
      50116: inst = 32'd136314880;
      50117: inst = 32'd268468224;
      50118: inst = 32'd201346822;
      50119: inst = 32'd203483685;
      50120: inst = 32'd471859200;
      50121: inst = 32'd136314880;
      50122: inst = 32'd268468224;
      50123: inst = 32'd201346823;
      50124: inst = 32'd203483685;
      50125: inst = 32'd471859200;
      50126: inst = 32'd136314880;
      50127: inst = 32'd268468224;
      50128: inst = 32'd201346824;
      50129: inst = 32'd203483685;
      50130: inst = 32'd471859200;
      50131: inst = 32'd136314880;
      50132: inst = 32'd268468224;
      50133: inst = 32'd201346825;
      50134: inst = 32'd203483685;
      50135: inst = 32'd471859200;
      50136: inst = 32'd136314880;
      50137: inst = 32'd268468224;
      50138: inst = 32'd201346826;
      50139: inst = 32'd203483685;
      50140: inst = 32'd471859200;
      50141: inst = 32'd136314880;
      50142: inst = 32'd268468224;
      50143: inst = 32'd201346827;
      50144: inst = 32'd203483685;
      50145: inst = 32'd471859200;
      50146: inst = 32'd136314880;
      50147: inst = 32'd268468224;
      50148: inst = 32'd201346828;
      50149: inst = 32'd203483685;
      50150: inst = 32'd471859200;
      50151: inst = 32'd136314880;
      50152: inst = 32'd268468224;
      50153: inst = 32'd201346829;
      50154: inst = 32'd203483685;
      50155: inst = 32'd471859200;
      50156: inst = 32'd136314880;
      50157: inst = 32'd268468224;
      50158: inst = 32'd201346830;
      50159: inst = 32'd203483685;
      50160: inst = 32'd471859200;
      50161: inst = 32'd136314880;
      50162: inst = 32'd268468224;
      50163: inst = 32'd201346831;
      50164: inst = 32'd203483685;
      50165: inst = 32'd471859200;
      50166: inst = 32'd136314880;
      50167: inst = 32'd268468224;
      50168: inst = 32'd201346832;
      50169: inst = 32'd203483685;
      50170: inst = 32'd471859200;
      50171: inst = 32'd136314880;
      50172: inst = 32'd268468224;
      50173: inst = 32'd201346833;
      50174: inst = 32'd203483685;
      50175: inst = 32'd471859200;
      50176: inst = 32'd136314880;
      50177: inst = 32'd268468224;
      50178: inst = 32'd201346834;
      50179: inst = 32'd203483685;
      50180: inst = 32'd471859200;
      50181: inst = 32'd136314880;
      50182: inst = 32'd268468224;
      50183: inst = 32'd201346835;
      50184: inst = 32'd203483685;
      50185: inst = 32'd471859200;
      50186: inst = 32'd136314880;
      50187: inst = 32'd268468224;
      50188: inst = 32'd201346836;
      50189: inst = 32'd203423744;
      50190: inst = 32'd471859200;
      50191: inst = 32'd136314880;
      50192: inst = 32'd268468224;
      50193: inst = 32'd201346837;
      50194: inst = 32'd203423744;
      50195: inst = 32'd471859200;
      50196: inst = 32'd136314880;
      50197: inst = 32'd268468224;
      50198: inst = 32'd201346838;
      50199: inst = 32'd203423744;
      50200: inst = 32'd471859200;
      50201: inst = 32'd136314880;
      50202: inst = 32'd268468224;
      50203: inst = 32'd201346839;
      50204: inst = 32'd203423744;
      50205: inst = 32'd471859200;
      50206: inst = 32'd136314880;
      50207: inst = 32'd268468224;
      50208: inst = 32'd201346840;
      50209: inst = 32'd203483685;
      50210: inst = 32'd471859200;
      50211: inst = 32'd136314880;
      50212: inst = 32'd268468224;
      50213: inst = 32'd201346841;
      50214: inst = 32'd203483685;
      50215: inst = 32'd471859200;
      50216: inst = 32'd136314880;
      50217: inst = 32'd268468224;
      50218: inst = 32'd201346842;
      50219: inst = 32'd203483685;
      50220: inst = 32'd471859200;
      50221: inst = 32'd136314880;
      50222: inst = 32'd268468224;
      50223: inst = 32'd201346843;
      50224: inst = 32'd203483685;
      50225: inst = 32'd471859200;
      50226: inst = 32'd136314880;
      50227: inst = 32'd268468224;
      50228: inst = 32'd201346844;
      50229: inst = 32'd203483685;
      50230: inst = 32'd471859200;
      50231: inst = 32'd136314880;
      50232: inst = 32'd268468224;
      50233: inst = 32'd201346845;
      50234: inst = 32'd203483685;
      50235: inst = 32'd471859200;
      50236: inst = 32'd136314880;
      50237: inst = 32'd268468224;
      50238: inst = 32'd201346846;
      50239: inst = 32'd203483685;
      50240: inst = 32'd471859200;
      50241: inst = 32'd136314880;
      50242: inst = 32'd268468224;
      50243: inst = 32'd201346847;
      50244: inst = 32'd203483685;
      50245: inst = 32'd471859200;
      50246: inst = 32'd136314880;
      50247: inst = 32'd268468224;
      50248: inst = 32'd201346848;
      50249: inst = 32'd203483685;
      50250: inst = 32'd471859200;
      50251: inst = 32'd136314880;
      50252: inst = 32'd268468224;
      50253: inst = 32'd201346849;
      50254: inst = 32'd203423744;
      50255: inst = 32'd471859200;
      50256: inst = 32'd136314880;
      50257: inst = 32'd268468224;
      50258: inst = 32'd201346850;
      50259: inst = 32'd203423744;
      50260: inst = 32'd471859200;
      50261: inst = 32'd136314880;
      50262: inst = 32'd268468224;
      50263: inst = 32'd201346851;
      50264: inst = 32'd203423744;
      50265: inst = 32'd471859200;
      50266: inst = 32'd136314880;
      50267: inst = 32'd268468224;
      50268: inst = 32'd201346852;
      50269: inst = 32'd203423744;
      50270: inst = 32'd471859200;
      50271: inst = 32'd136314880;
      50272: inst = 32'd268468224;
      50273: inst = 32'd201346853;
      50274: inst = 32'd203423744;
      50275: inst = 32'd471859200;
      50276: inst = 32'd136314880;
      50277: inst = 32'd268468224;
      50278: inst = 32'd201346854;
      50279: inst = 32'd203423744;
      50280: inst = 32'd471859200;
      50281: inst = 32'd136314880;
      50282: inst = 32'd268468224;
      50283: inst = 32'd201346855;
      50284: inst = 32'd203423744;
      50285: inst = 32'd471859200;
      50286: inst = 32'd136314880;
      50287: inst = 32'd268468224;
      50288: inst = 32'd201346856;
      50289: inst = 32'd203423744;
      50290: inst = 32'd471859200;
      50291: inst = 32'd136314880;
      50292: inst = 32'd268468224;
      50293: inst = 32'd201346857;
      50294: inst = 32'd203423744;
      50295: inst = 32'd471859200;
      50296: inst = 32'd136314880;
      50297: inst = 32'd268468224;
      50298: inst = 32'd201346858;
      50299: inst = 32'd203483685;
      50300: inst = 32'd471859200;
      50301: inst = 32'd136314880;
      50302: inst = 32'd268468224;
      50303: inst = 32'd201346859;
      50304: inst = 32'd203483685;
      50305: inst = 32'd471859200;
      50306: inst = 32'd136314880;
      50307: inst = 32'd268468224;
      50308: inst = 32'd201346860;
      50309: inst = 32'd203483685;
      50310: inst = 32'd471859200;
      50311: inst = 32'd136314880;
      50312: inst = 32'd268468224;
      50313: inst = 32'd201346861;
      50314: inst = 32'd203483685;
      50315: inst = 32'd471859200;
      50316: inst = 32'd136314880;
      50317: inst = 32'd268468224;
      50318: inst = 32'd201346862;
      50319: inst = 32'd203483685;
      50320: inst = 32'd471859200;
      50321: inst = 32'd136314880;
      50322: inst = 32'd268468224;
      50323: inst = 32'd201346863;
      50324: inst = 32'd203483685;
      50325: inst = 32'd471859200;
      50326: inst = 32'd136314880;
      50327: inst = 32'd268468224;
      50328: inst = 32'd201346864;
      50329: inst = 32'd203483685;
      50330: inst = 32'd471859200;
      50331: inst = 32'd136314880;
      50332: inst = 32'd268468224;
      50333: inst = 32'd201346865;
      50334: inst = 32'd203483685;
      50335: inst = 32'd471859200;
      50336: inst = 32'd136314880;
      50337: inst = 32'd268468224;
      50338: inst = 32'd201346866;
      50339: inst = 32'd203483685;
      50340: inst = 32'd471859200;
      50341: inst = 32'd136314880;
      50342: inst = 32'd268468224;
      50343: inst = 32'd201346867;
      50344: inst = 32'd203483685;
      50345: inst = 32'd471859200;
      50346: inst = 32'd136314880;
      50347: inst = 32'd268468224;
      50348: inst = 32'd201346868;
      50349: inst = 32'd203483685;
      50350: inst = 32'd471859200;
      50351: inst = 32'd136314880;
      50352: inst = 32'd268468224;
      50353: inst = 32'd201346869;
      50354: inst = 32'd203483685;
      50355: inst = 32'd471859200;
      50356: inst = 32'd136314880;
      50357: inst = 32'd268468224;
      50358: inst = 32'd201346870;
      50359: inst = 32'd203423744;
      50360: inst = 32'd471859200;
      50361: inst = 32'd136314880;
      50362: inst = 32'd268468224;
      50363: inst = 32'd201346871;
      50364: inst = 32'd203423744;
      50365: inst = 32'd471859200;
      50366: inst = 32'd136314880;
      50367: inst = 32'd268468224;
      50368: inst = 32'd201346872;
      50369: inst = 32'd203423744;
      50370: inst = 32'd471859200;
      50371: inst = 32'd136314880;
      50372: inst = 32'd268468224;
      50373: inst = 32'd201346873;
      50374: inst = 32'd203423744;
      50375: inst = 32'd471859200;
      50376: inst = 32'd136314880;
      50377: inst = 32'd268468224;
      50378: inst = 32'd201346874;
      50379: inst = 32'd203423744;
      50380: inst = 32'd471859200;
      50381: inst = 32'd136314880;
      50382: inst = 32'd268468224;
      50383: inst = 32'd201346875;
      50384: inst = 32'd203423744;
      50385: inst = 32'd471859200;
      50386: inst = 32'd136314880;
      50387: inst = 32'd268468224;
      50388: inst = 32'd201346876;
      50389: inst = 32'd203423744;
      50390: inst = 32'd471859200;
      50391: inst = 32'd136314880;
      50392: inst = 32'd268468224;
      50393: inst = 32'd201346877;
      50394: inst = 32'd203423744;
      50395: inst = 32'd471859200;
      50396: inst = 32'd136314880;
      50397: inst = 32'd268468224;
      50398: inst = 32'd201346878;
      50399: inst = 32'd203423744;
      50400: inst = 32'd471859200;
      50401: inst = 32'd136314880;
      50402: inst = 32'd268468224;
      50403: inst = 32'd201346879;
      50404: inst = 32'd203423744;
      50405: inst = 32'd471859200;
      50406: inst = 32'd136314880;
      50407: inst = 32'd268468224;
      50408: inst = 32'd201346880;
      50409: inst = 32'd203423744;
      50410: inst = 32'd471859200;
      50411: inst = 32'd136314880;
      50412: inst = 32'd268468224;
      50413: inst = 32'd201346881;
      50414: inst = 32'd203423744;
      50415: inst = 32'd471859200;
      50416: inst = 32'd136314880;
      50417: inst = 32'd268468224;
      50418: inst = 32'd201346882;
      50419: inst = 32'd203423744;
      50420: inst = 32'd471859200;
      50421: inst = 32'd136314880;
      50422: inst = 32'd268468224;
      50423: inst = 32'd201346883;
      50424: inst = 32'd203423744;
      50425: inst = 32'd471859200;
      50426: inst = 32'd136314880;
      50427: inst = 32'd268468224;
      50428: inst = 32'd201346884;
      50429: inst = 32'd203423744;
      50430: inst = 32'd471859200;
      50431: inst = 32'd136314880;
      50432: inst = 32'd268468224;
      50433: inst = 32'd201346885;
      50434: inst = 32'd203423744;
      50435: inst = 32'd471859200;
      50436: inst = 32'd136314880;
      50437: inst = 32'd268468224;
      50438: inst = 32'd201346886;
      50439: inst = 32'd203423744;
      50440: inst = 32'd471859200;
      50441: inst = 32'd136314880;
      50442: inst = 32'd268468224;
      50443: inst = 32'd201346887;
      50444: inst = 32'd203423744;
      50445: inst = 32'd471859200;
      50446: inst = 32'd136314880;
      50447: inst = 32'd268468224;
      50448: inst = 32'd201346888;
      50449: inst = 32'd203423744;
      50450: inst = 32'd471859200;
      50451: inst = 32'd136314880;
      50452: inst = 32'd268468224;
      50453: inst = 32'd201346889;
      50454: inst = 32'd203423744;
      50455: inst = 32'd471859200;
      50456: inst = 32'd136314880;
      50457: inst = 32'd268468224;
      50458: inst = 32'd201346890;
      50459: inst = 32'd203423744;
      50460: inst = 32'd471859200;
      50461: inst = 32'd136314880;
      50462: inst = 32'd268468224;
      50463: inst = 32'd201346891;
      50464: inst = 32'd203423744;
      50465: inst = 32'd471859200;
      50466: inst = 32'd136314880;
      50467: inst = 32'd268468224;
      50468: inst = 32'd201346892;
      50469: inst = 32'd203423744;
      50470: inst = 32'd471859200;
      50471: inst = 32'd136314880;
      50472: inst = 32'd268468224;
      50473: inst = 32'd201346893;
      50474: inst = 32'd203483685;
      50475: inst = 32'd471859200;
      50476: inst = 32'd136314880;
      50477: inst = 32'd268468224;
      50478: inst = 32'd201346894;
      50479: inst = 32'd203483685;
      50480: inst = 32'd471859200;
      50481: inst = 32'd136314880;
      50482: inst = 32'd268468224;
      50483: inst = 32'd201346895;
      50484: inst = 32'd203483685;
      50485: inst = 32'd471859200;
      50486: inst = 32'd136314880;
      50487: inst = 32'd268468224;
      50488: inst = 32'd201346896;
      50489: inst = 32'd203483685;
      50490: inst = 32'd471859200;
      50491: inst = 32'd136314880;
      50492: inst = 32'd268468224;
      50493: inst = 32'd201346897;
      50494: inst = 32'd203483685;
      50495: inst = 32'd471859200;
      50496: inst = 32'd136314880;
      50497: inst = 32'd268468224;
      50498: inst = 32'd201346898;
      50499: inst = 32'd203483685;
      50500: inst = 32'd471859200;
      50501: inst = 32'd136314880;
      50502: inst = 32'd268468224;
      50503: inst = 32'd201346899;
      50504: inst = 32'd203483685;
      50505: inst = 32'd471859200;
      50506: inst = 32'd136314880;
      50507: inst = 32'd268468224;
      50508: inst = 32'd201346900;
      50509: inst = 32'd203483685;
      50510: inst = 32'd471859200;
      50511: inst = 32'd136314880;
      50512: inst = 32'd268468224;
      50513: inst = 32'd201346901;
      50514: inst = 32'd203483685;
      50515: inst = 32'd471859200;
      50516: inst = 32'd136314880;
      50517: inst = 32'd268468224;
      50518: inst = 32'd201346902;
      50519: inst = 32'd203483685;
      50520: inst = 32'd471859200;
      50521: inst = 32'd136314880;
      50522: inst = 32'd268468224;
      50523: inst = 32'd201346903;
      50524: inst = 32'd203423744;
      50525: inst = 32'd471859200;
      50526: inst = 32'd136314880;
      50527: inst = 32'd268468224;
      50528: inst = 32'd201346904;
      50529: inst = 32'd203483685;
      50530: inst = 32'd471859200;
      50531: inst = 32'd136314880;
      50532: inst = 32'd268468224;
      50533: inst = 32'd201346905;
      50534: inst = 32'd203483685;
      50535: inst = 32'd471859200;
      50536: inst = 32'd136314880;
      50537: inst = 32'd268468224;
      50538: inst = 32'd201346906;
      50539: inst = 32'd203483685;
      50540: inst = 32'd471859200;
      50541: inst = 32'd136314880;
      50542: inst = 32'd268468224;
      50543: inst = 32'd201346907;
      50544: inst = 32'd203483685;
      50545: inst = 32'd471859200;
      50546: inst = 32'd136314880;
      50547: inst = 32'd268468224;
      50548: inst = 32'd201346908;
      50549: inst = 32'd203483685;
      50550: inst = 32'd471859200;
      50551: inst = 32'd136314880;
      50552: inst = 32'd268468224;
      50553: inst = 32'd201346909;
      50554: inst = 32'd203483685;
      50555: inst = 32'd471859200;
      50556: inst = 32'd136314880;
      50557: inst = 32'd268468224;
      50558: inst = 32'd201346910;
      50559: inst = 32'd203483685;
      50560: inst = 32'd471859200;
      50561: inst = 32'd136314880;
      50562: inst = 32'd268468224;
      50563: inst = 32'd201346911;
      50564: inst = 32'd203483685;
      50565: inst = 32'd471859200;
      50566: inst = 32'd136314880;
      50567: inst = 32'd268468224;
      50568: inst = 32'd201346912;
      50569: inst = 32'd203483685;
      50570: inst = 32'd471859200;
      50571: inst = 32'd136314880;
      50572: inst = 32'd268468224;
      50573: inst = 32'd201346913;
      50574: inst = 32'd203483685;
      50575: inst = 32'd471859200;
      50576: inst = 32'd136314880;
      50577: inst = 32'd268468224;
      50578: inst = 32'd201346914;
      50579: inst = 32'd203483685;
      50580: inst = 32'd471859200;
      50581: inst = 32'd136314880;
      50582: inst = 32'd268468224;
      50583: inst = 32'd201346915;
      50584: inst = 32'd203483685;
      50585: inst = 32'd471859200;
      50586: inst = 32'd136314880;
      50587: inst = 32'd268468224;
      50588: inst = 32'd201346916;
      50589: inst = 32'd203483685;
      50590: inst = 32'd471859200;
      50591: inst = 32'd136314880;
      50592: inst = 32'd268468224;
      50593: inst = 32'd201346917;
      50594: inst = 32'd203423744;
      50595: inst = 32'd471859200;
      50596: inst = 32'd136314880;
      50597: inst = 32'd268468224;
      50598: inst = 32'd201346918;
      50599: inst = 32'd203423744;
      50600: inst = 32'd471859200;
      50601: inst = 32'd136314880;
      50602: inst = 32'd268468224;
      50603: inst = 32'd201346919;
      50604: inst = 32'd203483685;
      50605: inst = 32'd471859200;
      50606: inst = 32'd136314880;
      50607: inst = 32'd268468224;
      50608: inst = 32'd201346920;
      50609: inst = 32'd203483685;
      50610: inst = 32'd471859200;
      50611: inst = 32'd136314880;
      50612: inst = 32'd268468224;
      50613: inst = 32'd201346921;
      50614: inst = 32'd203483685;
      50615: inst = 32'd471859200;
      50616: inst = 32'd136314880;
      50617: inst = 32'd268468224;
      50618: inst = 32'd201346922;
      50619: inst = 32'd203483685;
      50620: inst = 32'd471859200;
      50621: inst = 32'd136314880;
      50622: inst = 32'd268468224;
      50623: inst = 32'd201346923;
      50624: inst = 32'd203483685;
      50625: inst = 32'd471859200;
      50626: inst = 32'd136314880;
      50627: inst = 32'd268468224;
      50628: inst = 32'd201346924;
      50629: inst = 32'd203483685;
      50630: inst = 32'd471859200;
      50631: inst = 32'd136314880;
      50632: inst = 32'd268468224;
      50633: inst = 32'd201346925;
      50634: inst = 32'd203483685;
      50635: inst = 32'd471859200;
      50636: inst = 32'd136314880;
      50637: inst = 32'd268468224;
      50638: inst = 32'd201346926;
      50639: inst = 32'd203483685;
      50640: inst = 32'd471859200;
      50641: inst = 32'd136314880;
      50642: inst = 32'd268468224;
      50643: inst = 32'd201346927;
      50644: inst = 32'd203483685;
      50645: inst = 32'd471859200;
      50646: inst = 32'd136314880;
      50647: inst = 32'd268468224;
      50648: inst = 32'd201346928;
      50649: inst = 32'd203483685;
      50650: inst = 32'd471859200;
      50651: inst = 32'd136314880;
      50652: inst = 32'd268468224;
      50653: inst = 32'd201346929;
      50654: inst = 32'd203483685;
      50655: inst = 32'd471859200;
      50656: inst = 32'd136314880;
      50657: inst = 32'd268468224;
      50658: inst = 32'd201346930;
      50659: inst = 32'd203483685;
      50660: inst = 32'd471859200;
      50661: inst = 32'd136314880;
      50662: inst = 32'd268468224;
      50663: inst = 32'd201346931;
      50664: inst = 32'd203483685;
      50665: inst = 32'd471859200;
      50666: inst = 32'd136314880;
      50667: inst = 32'd268468224;
      50668: inst = 32'd201346932;
      50669: inst = 32'd203423744;
      50670: inst = 32'd471859200;
      50671: inst = 32'd136314880;
      50672: inst = 32'd268468224;
      50673: inst = 32'd201346933;
      50674: inst = 32'd203423744;
      50675: inst = 32'd471859200;
      50676: inst = 32'd136314880;
      50677: inst = 32'd268468224;
      50678: inst = 32'd201346934;
      50679: inst = 32'd203423744;
      50680: inst = 32'd471859200;
      50681: inst = 32'd136314880;
      50682: inst = 32'd268468224;
      50683: inst = 32'd201346935;
      50684: inst = 32'd203423744;
      50685: inst = 32'd471859200;
      50686: inst = 32'd136314880;
      50687: inst = 32'd268468224;
      50688: inst = 32'd201346936;
      50689: inst = 32'd203423744;
      50690: inst = 32'd471859200;
      50691: inst = 32'd136314880;
      50692: inst = 32'd268468224;
      50693: inst = 32'd201346937;
      50694: inst = 32'd203483685;
      50695: inst = 32'd471859200;
      50696: inst = 32'd136314880;
      50697: inst = 32'd268468224;
      50698: inst = 32'd201346938;
      50699: inst = 32'd203483685;
      50700: inst = 32'd471859200;
      50701: inst = 32'd136314880;
      50702: inst = 32'd268468224;
      50703: inst = 32'd201346939;
      50704: inst = 32'd203483685;
      50705: inst = 32'd471859200;
      50706: inst = 32'd136314880;
      50707: inst = 32'd268468224;
      50708: inst = 32'd201346940;
      50709: inst = 32'd203483685;
      50710: inst = 32'd471859200;
      50711: inst = 32'd136314880;
      50712: inst = 32'd268468224;
      50713: inst = 32'd201346941;
      50714: inst = 32'd203483685;
      50715: inst = 32'd471859200;
      50716: inst = 32'd136314880;
      50717: inst = 32'd268468224;
      50718: inst = 32'd201346942;
      50719: inst = 32'd203483685;
      50720: inst = 32'd471859200;
      50721: inst = 32'd136314880;
      50722: inst = 32'd268468224;
      50723: inst = 32'd201346943;
      50724: inst = 32'd203483685;
      50725: inst = 32'd471859200;
      50726: inst = 32'd136314880;
      50727: inst = 32'd268468224;
      50728: inst = 32'd201346944;
      50729: inst = 32'd203483685;
      50730: inst = 32'd471859200;
      50731: inst = 32'd136314880;
      50732: inst = 32'd268468224;
      50733: inst = 32'd201346945;
      50734: inst = 32'd203423744;
      50735: inst = 32'd471859200;
      50736: inst = 32'd136314880;
      50737: inst = 32'd268468224;
      50738: inst = 32'd201346946;
      50739: inst = 32'd203423744;
      50740: inst = 32'd471859200;
      50741: inst = 32'd136314880;
      50742: inst = 32'd268468224;
      50743: inst = 32'd201346947;
      50744: inst = 32'd203423744;
      50745: inst = 32'd471859200;
      50746: inst = 32'd136314880;
      50747: inst = 32'd268468224;
      50748: inst = 32'd201346948;
      50749: inst = 32'd203423744;
      50750: inst = 32'd471859200;
      50751: inst = 32'd136314880;
      50752: inst = 32'd268468224;
      50753: inst = 32'd201346949;
      50754: inst = 32'd203423744;
      50755: inst = 32'd471859200;
      50756: inst = 32'd136314880;
      50757: inst = 32'd268468224;
      50758: inst = 32'd201346950;
      50759: inst = 32'd203423744;
      50760: inst = 32'd471859200;
      50761: inst = 32'd136314880;
      50762: inst = 32'd268468224;
      50763: inst = 32'd201346951;
      50764: inst = 32'd203423744;
      50765: inst = 32'd471859200;
      50766: inst = 32'd136314880;
      50767: inst = 32'd268468224;
      50768: inst = 32'd201346952;
      50769: inst = 32'd203423744;
      50770: inst = 32'd471859200;
      50771: inst = 32'd136314880;
      50772: inst = 32'd268468224;
      50773: inst = 32'd201346953;
      50774: inst = 32'd203423744;
      50775: inst = 32'd471859200;
      50776: inst = 32'd136314880;
      50777: inst = 32'd268468224;
      50778: inst = 32'd201346954;
      50779: inst = 32'd203483685;
      50780: inst = 32'd471859200;
      50781: inst = 32'd136314880;
      50782: inst = 32'd268468224;
      50783: inst = 32'd201346955;
      50784: inst = 32'd203483685;
      50785: inst = 32'd471859200;
      50786: inst = 32'd136314880;
      50787: inst = 32'd268468224;
      50788: inst = 32'd201346956;
      50789: inst = 32'd203483685;
      50790: inst = 32'd471859200;
      50791: inst = 32'd136314880;
      50792: inst = 32'd268468224;
      50793: inst = 32'd201346957;
      50794: inst = 32'd203483685;
      50795: inst = 32'd471859200;
      50796: inst = 32'd136314880;
      50797: inst = 32'd268468224;
      50798: inst = 32'd201346958;
      50799: inst = 32'd203483685;
      50800: inst = 32'd471859200;
      50801: inst = 32'd136314880;
      50802: inst = 32'd268468224;
      50803: inst = 32'd201346959;
      50804: inst = 32'd203483685;
      50805: inst = 32'd471859200;
      50806: inst = 32'd136314880;
      50807: inst = 32'd268468224;
      50808: inst = 32'd201346960;
      50809: inst = 32'd203483685;
      50810: inst = 32'd471859200;
      50811: inst = 32'd136314880;
      50812: inst = 32'd268468224;
      50813: inst = 32'd201346961;
      50814: inst = 32'd203483685;
      50815: inst = 32'd471859200;
      50816: inst = 32'd136314880;
      50817: inst = 32'd268468224;
      50818: inst = 32'd201346962;
      50819: inst = 32'd203483685;
      50820: inst = 32'd471859200;
      50821: inst = 32'd136314880;
      50822: inst = 32'd268468224;
      50823: inst = 32'd201346963;
      50824: inst = 32'd203483685;
      50825: inst = 32'd471859200;
      50826: inst = 32'd136314880;
      50827: inst = 32'd268468224;
      50828: inst = 32'd201346964;
      50829: inst = 32'd203423744;
      50830: inst = 32'd471859200;
      50831: inst = 32'd136314880;
      50832: inst = 32'd268468224;
      50833: inst = 32'd201346965;
      50834: inst = 32'd203423744;
      50835: inst = 32'd471859200;
      50836: inst = 32'd136314880;
      50837: inst = 32'd268468224;
      50838: inst = 32'd201346966;
      50839: inst = 32'd203423744;
      50840: inst = 32'd471859200;
      50841: inst = 32'd136314880;
      50842: inst = 32'd268468224;
      50843: inst = 32'd201346967;
      50844: inst = 32'd203423744;
      50845: inst = 32'd471859200;
      50846: inst = 32'd136314880;
      50847: inst = 32'd268468224;
      50848: inst = 32'd201346968;
      50849: inst = 32'd203423744;
      50850: inst = 32'd471859200;
      50851: inst = 32'd136314880;
      50852: inst = 32'd268468224;
      50853: inst = 32'd201346969;
      50854: inst = 32'd203423744;
      50855: inst = 32'd471859200;
      50856: inst = 32'd136314880;
      50857: inst = 32'd268468224;
      50858: inst = 32'd201346970;
      50859: inst = 32'd203423744;
      50860: inst = 32'd471859200;
      50861: inst = 32'd136314880;
      50862: inst = 32'd268468224;
      50863: inst = 32'd201346971;
      50864: inst = 32'd203423744;
      50865: inst = 32'd471859200;
      50866: inst = 32'd136314880;
      50867: inst = 32'd268468224;
      50868: inst = 32'd201346972;
      50869: inst = 32'd203423744;
      50870: inst = 32'd471859200;
      50871: inst = 32'd136314880;
      50872: inst = 32'd268468224;
      50873: inst = 32'd201346973;
      50874: inst = 32'd203423744;
      50875: inst = 32'd471859200;
      50876: inst = 32'd136314880;
      50877: inst = 32'd268468224;
      50878: inst = 32'd201346974;
      50879: inst = 32'd203423744;
      50880: inst = 32'd471859200;
      50881: inst = 32'd136314880;
      50882: inst = 32'd268468224;
      50883: inst = 32'd201346975;
      50884: inst = 32'd203423744;
      50885: inst = 32'd471859200;
      50886: inst = 32'd136314880;
      50887: inst = 32'd268468224;
      50888: inst = 32'd201346976;
      50889: inst = 32'd203423744;
      50890: inst = 32'd471859200;
      50891: inst = 32'd136314880;
      50892: inst = 32'd268468224;
      50893: inst = 32'd201346977;
      50894: inst = 32'd203423744;
      50895: inst = 32'd471859200;
      50896: inst = 32'd136314880;
      50897: inst = 32'd268468224;
      50898: inst = 32'd201346978;
      50899: inst = 32'd203423744;
      50900: inst = 32'd471859200;
      50901: inst = 32'd136314880;
      50902: inst = 32'd268468224;
      50903: inst = 32'd201346979;
      50904: inst = 32'd203423744;
      50905: inst = 32'd471859200;
      50906: inst = 32'd136314880;
      50907: inst = 32'd268468224;
      50908: inst = 32'd201346980;
      50909: inst = 32'd203423744;
      50910: inst = 32'd471859200;
      50911: inst = 32'd136314880;
      50912: inst = 32'd268468224;
      50913: inst = 32'd201346981;
      50914: inst = 32'd203423744;
      50915: inst = 32'd471859200;
      50916: inst = 32'd136314880;
      50917: inst = 32'd268468224;
      50918: inst = 32'd201346982;
      50919: inst = 32'd203423744;
      50920: inst = 32'd471859200;
      50921: inst = 32'd136314880;
      50922: inst = 32'd268468224;
      50923: inst = 32'd201346983;
      50924: inst = 32'd203423744;
      50925: inst = 32'd471859200;
      50926: inst = 32'd136314880;
      50927: inst = 32'd268468224;
      50928: inst = 32'd201346984;
      50929: inst = 32'd203423744;
      50930: inst = 32'd471859200;
      50931: inst = 32'd136314880;
      50932: inst = 32'd268468224;
      50933: inst = 32'd201346985;
      50934: inst = 32'd203423744;
      50935: inst = 32'd471859200;
      50936: inst = 32'd136314880;
      50937: inst = 32'd268468224;
      50938: inst = 32'd201346986;
      50939: inst = 32'd203423744;
      50940: inst = 32'd471859200;
      50941: inst = 32'd136314880;
      50942: inst = 32'd268468224;
      50943: inst = 32'd201346987;
      50944: inst = 32'd203423744;
      50945: inst = 32'd471859200;
      50946: inst = 32'd136314880;
      50947: inst = 32'd268468224;
      50948: inst = 32'd201346988;
      50949: inst = 32'd203423744;
      50950: inst = 32'd471859200;
      50951: inst = 32'd136314880;
      50952: inst = 32'd268468224;
      50953: inst = 32'd201346989;
      50954: inst = 32'd203423744;
      50955: inst = 32'd471859200;
      50956: inst = 32'd136314880;
      50957: inst = 32'd268468224;
      50958: inst = 32'd201346990;
      50959: inst = 32'd203423744;
      50960: inst = 32'd471859200;
      50961: inst = 32'd136314880;
      50962: inst = 32'd268468224;
      50963: inst = 32'd201346991;
      50964: inst = 32'd203423744;
      50965: inst = 32'd471859200;
      50966: inst = 32'd136314880;
      50967: inst = 32'd268468224;
      50968: inst = 32'd201346992;
      50969: inst = 32'd203423744;
      50970: inst = 32'd471859200;
      50971: inst = 32'd136314880;
      50972: inst = 32'd268468224;
      50973: inst = 32'd201346993;
      50974: inst = 32'd203423744;
      50975: inst = 32'd471859200;
      50976: inst = 32'd136314880;
      50977: inst = 32'd268468224;
      50978: inst = 32'd201346994;
      50979: inst = 32'd203423744;
      50980: inst = 32'd471859200;
      50981: inst = 32'd136314880;
      50982: inst = 32'd268468224;
      50983: inst = 32'd201346995;
      50984: inst = 32'd203423744;
      50985: inst = 32'd471859200;
      50986: inst = 32'd136314880;
      50987: inst = 32'd268468224;
      50988: inst = 32'd201346996;
      50989: inst = 32'd203423744;
      50990: inst = 32'd471859200;
      50991: inst = 32'd136314880;
      50992: inst = 32'd268468224;
      50993: inst = 32'd201346997;
      50994: inst = 32'd203423744;
      50995: inst = 32'd471859200;
      50996: inst = 32'd136314880;
      50997: inst = 32'd268468224;
      50998: inst = 32'd201346998;
      50999: inst = 32'd203423744;
      51000: inst = 32'd471859200;
      51001: inst = 32'd136314880;
      51002: inst = 32'd268468224;
      51003: inst = 32'd201346999;
      51004: inst = 32'd203423744;
      51005: inst = 32'd471859200;
      51006: inst = 32'd136314880;
      51007: inst = 32'd268468224;
      51008: inst = 32'd201347000;
      51009: inst = 32'd203423744;
      51010: inst = 32'd471859200;
      51011: inst = 32'd136314880;
      51012: inst = 32'd268468224;
      51013: inst = 32'd201347001;
      51014: inst = 32'd203423744;
      51015: inst = 32'd471859200;
      51016: inst = 32'd136314880;
      51017: inst = 32'd268468224;
      51018: inst = 32'd201347002;
      51019: inst = 32'd203423744;
      51020: inst = 32'd471859200;
      51021: inst = 32'd136314880;
      51022: inst = 32'd268468224;
      51023: inst = 32'd201347003;
      51024: inst = 32'd203423744;
      51025: inst = 32'd471859200;
      51026: inst = 32'd136314880;
      51027: inst = 32'd268468224;
      51028: inst = 32'd201347004;
      51029: inst = 32'd203423744;
      51030: inst = 32'd471859200;
      51031: inst = 32'd136314880;
      51032: inst = 32'd268468224;
      51033: inst = 32'd201347005;
      51034: inst = 32'd203423744;
      51035: inst = 32'd471859200;
      51036: inst = 32'd136314880;
      51037: inst = 32'd268468224;
      51038: inst = 32'd201347006;
      51039: inst = 32'd203423744;
      51040: inst = 32'd471859200;
      51041: inst = 32'd136314880;
      51042: inst = 32'd268468224;
      51043: inst = 32'd201347007;
      51044: inst = 32'd203423744;
      51045: inst = 32'd471859200;
      51046: inst = 32'd136314880;
      51047: inst = 32'd268468224;
      51048: inst = 32'd201347008;
      51049: inst = 32'd203423744;
      51050: inst = 32'd471859200;
      51051: inst = 32'd136314880;
      51052: inst = 32'd268468224;
      51053: inst = 32'd201347009;
      51054: inst = 32'd203423744;
      51055: inst = 32'd471859200;
      51056: inst = 32'd136314880;
      51057: inst = 32'd268468224;
      51058: inst = 32'd201347010;
      51059: inst = 32'd203423744;
      51060: inst = 32'd471859200;
      51061: inst = 32'd136314880;
      51062: inst = 32'd268468224;
      51063: inst = 32'd201347011;
      51064: inst = 32'd203423744;
      51065: inst = 32'd471859200;
      51066: inst = 32'd136314880;
      51067: inst = 32'd268468224;
      51068: inst = 32'd201347012;
      51069: inst = 32'd203423744;
      51070: inst = 32'd471859200;
      51071: inst = 32'd136314880;
      51072: inst = 32'd268468224;
      51073: inst = 32'd201347013;
      51074: inst = 32'd203423744;
      51075: inst = 32'd471859200;
      51076: inst = 32'd136314880;
      51077: inst = 32'd268468224;
      51078: inst = 32'd201347014;
      51079: inst = 32'd203423744;
      51080: inst = 32'd471859200;
      51081: inst = 32'd136314880;
      51082: inst = 32'd268468224;
      51083: inst = 32'd201347015;
      51084: inst = 32'd203423744;
      51085: inst = 32'd471859200;
      51086: inst = 32'd136314880;
      51087: inst = 32'd268468224;
      51088: inst = 32'd201347016;
      51089: inst = 32'd203423744;
      51090: inst = 32'd471859200;
      51091: inst = 32'd136314880;
      51092: inst = 32'd268468224;
      51093: inst = 32'd201347017;
      51094: inst = 32'd203423744;
      51095: inst = 32'd471859200;
      51096: inst = 32'd136314880;
      51097: inst = 32'd268468224;
      51098: inst = 32'd201347018;
      51099: inst = 32'd203423744;
      51100: inst = 32'd471859200;
      51101: inst = 32'd136314880;
      51102: inst = 32'd268468224;
      51103: inst = 32'd201347019;
      51104: inst = 32'd203423744;
      51105: inst = 32'd471859200;
      51106: inst = 32'd136314880;
      51107: inst = 32'd268468224;
      51108: inst = 32'd201347020;
      51109: inst = 32'd203423744;
      51110: inst = 32'd471859200;
      51111: inst = 32'd136314880;
      51112: inst = 32'd268468224;
      51113: inst = 32'd201347021;
      51114: inst = 32'd203423744;
      51115: inst = 32'd471859200;
      51116: inst = 32'd136314880;
      51117: inst = 32'd268468224;
      51118: inst = 32'd201347022;
      51119: inst = 32'd203423744;
      51120: inst = 32'd471859200;
      51121: inst = 32'd136314880;
      51122: inst = 32'd268468224;
      51123: inst = 32'd201347023;
      51124: inst = 32'd203423744;
      51125: inst = 32'd471859200;
      51126: inst = 32'd136314880;
      51127: inst = 32'd268468224;
      51128: inst = 32'd201347024;
      51129: inst = 32'd203423744;
      51130: inst = 32'd471859200;
      51131: inst = 32'd136314880;
      51132: inst = 32'd268468224;
      51133: inst = 32'd201347025;
      51134: inst = 32'd203423744;
      51135: inst = 32'd471859200;
      51136: inst = 32'd136314880;
      51137: inst = 32'd268468224;
      51138: inst = 32'd201347026;
      51139: inst = 32'd203423744;
      51140: inst = 32'd471859200;
      51141: inst = 32'd136314880;
      51142: inst = 32'd268468224;
      51143: inst = 32'd201347027;
      51144: inst = 32'd203423744;
      51145: inst = 32'd471859200;
      51146: inst = 32'd136314880;
      51147: inst = 32'd268468224;
      51148: inst = 32'd201347028;
      51149: inst = 32'd203423744;
      51150: inst = 32'd471859200;
      51151: inst = 32'd136314880;
      51152: inst = 32'd268468224;
      51153: inst = 32'd201347029;
      51154: inst = 32'd203423744;
      51155: inst = 32'd471859200;
      51156: inst = 32'd136314880;
      51157: inst = 32'd268468224;
      51158: inst = 32'd201347030;
      51159: inst = 32'd203423744;
      51160: inst = 32'd471859200;
      51161: inst = 32'd136314880;
      51162: inst = 32'd268468224;
      51163: inst = 32'd201347031;
      51164: inst = 32'd203423744;
      51165: inst = 32'd471859200;
      51166: inst = 32'd136314880;
      51167: inst = 32'd268468224;
      51168: inst = 32'd201347032;
      51169: inst = 32'd203423744;
      51170: inst = 32'd471859200;
      51171: inst = 32'd136314880;
      51172: inst = 32'd268468224;
      51173: inst = 32'd201347033;
      51174: inst = 32'd203423744;
      51175: inst = 32'd471859200;
      51176: inst = 32'd136314880;
      51177: inst = 32'd268468224;
      51178: inst = 32'd201347034;
      51179: inst = 32'd203423744;
      51180: inst = 32'd471859200;
      51181: inst = 32'd136314880;
      51182: inst = 32'd268468224;
      51183: inst = 32'd201347035;
      51184: inst = 32'd203423744;
      51185: inst = 32'd471859200;
      51186: inst = 32'd136314880;
      51187: inst = 32'd268468224;
      51188: inst = 32'd201347036;
      51189: inst = 32'd203423744;
      51190: inst = 32'd471859200;
      51191: inst = 32'd136314880;
      51192: inst = 32'd268468224;
      51193: inst = 32'd201347037;
      51194: inst = 32'd203423744;
      51195: inst = 32'd471859200;
      51196: inst = 32'd136314880;
      51197: inst = 32'd268468224;
      51198: inst = 32'd201347038;
      51199: inst = 32'd203423744;
      51200: inst = 32'd471859200;
      51201: inst = 32'd136314880;
      51202: inst = 32'd268468224;
      51203: inst = 32'd201347039;
      51204: inst = 32'd203423744;
      51205: inst = 32'd471859200;
      51206: inst = 32'd136314880;
      51207: inst = 32'd268468224;
      51208: inst = 32'd201347040;
      51209: inst = 32'd203423744;
      51210: inst = 32'd471859200;
      51211: inst = 32'd136314880;
      51212: inst = 32'd268468224;
      51213: inst = 32'd201347041;
      51214: inst = 32'd203423744;
      51215: inst = 32'd471859200;
      51216: inst = 32'd136314880;
      51217: inst = 32'd268468224;
      51218: inst = 32'd201347042;
      51219: inst = 32'd203423744;
      51220: inst = 32'd471859200;
      51221: inst = 32'd136314880;
      51222: inst = 32'd268468224;
      51223: inst = 32'd201347043;
      51224: inst = 32'd203423744;
      51225: inst = 32'd471859200;
      51226: inst = 32'd136314880;
      51227: inst = 32'd268468224;
      51228: inst = 32'd201347044;
      51229: inst = 32'd203423744;
      51230: inst = 32'd471859200;
      51231: inst = 32'd136314880;
      51232: inst = 32'd268468224;
      51233: inst = 32'd201347045;
      51234: inst = 32'd203423744;
      51235: inst = 32'd471859200;
      51236: inst = 32'd136314880;
      51237: inst = 32'd268468224;
      51238: inst = 32'd201347046;
      51239: inst = 32'd203423744;
      51240: inst = 32'd471859200;
      51241: inst = 32'd136314880;
      51242: inst = 32'd268468224;
      51243: inst = 32'd201347047;
      51244: inst = 32'd203423744;
      51245: inst = 32'd471859200;
      51246: inst = 32'd136314880;
      51247: inst = 32'd268468224;
      51248: inst = 32'd201347048;
      51249: inst = 32'd203423744;
      51250: inst = 32'd471859200;
      51251: inst = 32'd136314880;
      51252: inst = 32'd268468224;
      51253: inst = 32'd201347049;
      51254: inst = 32'd203423744;
      51255: inst = 32'd471859200;
      51256: inst = 32'd136314880;
      51257: inst = 32'd268468224;
      51258: inst = 32'd201347050;
      51259: inst = 32'd203423744;
      51260: inst = 32'd471859200;
      51261: inst = 32'd136314880;
      51262: inst = 32'd268468224;
      51263: inst = 32'd201347051;
      51264: inst = 32'd203423744;
      51265: inst = 32'd471859200;
      51266: inst = 32'd136314880;
      51267: inst = 32'd268468224;
      51268: inst = 32'd201347052;
      51269: inst = 32'd203423744;
      51270: inst = 32'd471859200;
      51271: inst = 32'd136314880;
      51272: inst = 32'd268468224;
      51273: inst = 32'd201347053;
      51274: inst = 32'd203423744;
      51275: inst = 32'd471859200;
      51276: inst = 32'd136314880;
      51277: inst = 32'd268468224;
      51278: inst = 32'd201347054;
      51279: inst = 32'd203423744;
      51280: inst = 32'd471859200;
      51281: inst = 32'd136314880;
      51282: inst = 32'd268468224;
      51283: inst = 32'd201347055;
      51284: inst = 32'd203423744;
      51285: inst = 32'd471859200;
      51286: inst = 32'd136314880;
      51287: inst = 32'd268468224;
      51288: inst = 32'd201347056;
      51289: inst = 32'd203423744;
      51290: inst = 32'd471859200;
      51291: inst = 32'd136314880;
      51292: inst = 32'd268468224;
      51293: inst = 32'd201347057;
      51294: inst = 32'd203423744;
      51295: inst = 32'd471859200;
      51296: inst = 32'd136314880;
      51297: inst = 32'd268468224;
      51298: inst = 32'd201347058;
      51299: inst = 32'd203423744;
      51300: inst = 32'd471859200;
      51301: inst = 32'd136314880;
      51302: inst = 32'd268468224;
      51303: inst = 32'd201347059;
      51304: inst = 32'd203423744;
      51305: inst = 32'd471859200;
      51306: inst = 32'd136314880;
      51307: inst = 32'd268468224;
      51308: inst = 32'd201347060;
      51309: inst = 32'd203423744;
      51310: inst = 32'd471859200;
      51311: inst = 32'd136314880;
      51312: inst = 32'd268468224;
      51313: inst = 32'd201347061;
      51314: inst = 32'd203423744;
      51315: inst = 32'd471859200;
      51316: inst = 32'd136314880;
      51317: inst = 32'd268468224;
      51318: inst = 32'd201347062;
      51319: inst = 32'd203423744;
      51320: inst = 32'd471859200;
      51321: inst = 32'd136314880;
      51322: inst = 32'd268468224;
      51323: inst = 32'd201347063;
      51324: inst = 32'd203423744;
      51325: inst = 32'd471859200;
      51326: inst = 32'd136314880;
      51327: inst = 32'd268468224;
      51328: inst = 32'd201347064;
      51329: inst = 32'd203423744;
      51330: inst = 32'd471859200;
      51331: inst = 32'd136314880;
      51332: inst = 32'd268468224;
      51333: inst = 32'd201347065;
      51334: inst = 32'd203423744;
      51335: inst = 32'd471859200;
      51336: inst = 32'd136314880;
      51337: inst = 32'd268468224;
      51338: inst = 32'd201347066;
      51339: inst = 32'd203423744;
      51340: inst = 32'd471859200;
      51341: inst = 32'd136314880;
      51342: inst = 32'd268468224;
      51343: inst = 32'd201347067;
      51344: inst = 32'd203423744;
      51345: inst = 32'd471859200;
      51346: inst = 32'd136314880;
      51347: inst = 32'd268468224;
      51348: inst = 32'd201347068;
      51349: inst = 32'd203423744;
      51350: inst = 32'd471859200;
      51351: inst = 32'd136314880;
      51352: inst = 32'd268468224;
      51353: inst = 32'd201347069;
      51354: inst = 32'd203423744;
      51355: inst = 32'd471859200;
      51356: inst = 32'd136314880;
      51357: inst = 32'd268468224;
      51358: inst = 32'd201347070;
      51359: inst = 32'd203423744;
      51360: inst = 32'd471859200;
      51361: inst = 32'd136314880;
      51362: inst = 32'd268468224;
      51363: inst = 32'd201347071;
      51364: inst = 32'd203423744;
      51365: inst = 32'd471859200;
      51366: inst = 32'd136314880;
      51367: inst = 32'd268468224;
      51368: inst = 32'd201347072;
      51369: inst = 32'd203423744;
      51370: inst = 32'd471859200;
      51371: inst = 32'd136314880;
      51372: inst = 32'd268468224;
      51373: inst = 32'd201347073;
      51374: inst = 32'd203423744;
      51375: inst = 32'd471859200;
      51376: inst = 32'd136314880;
      51377: inst = 32'd268468224;
      51378: inst = 32'd201347074;
      51379: inst = 32'd203423744;
      51380: inst = 32'd471859200;
      51381: inst = 32'd136314880;
      51382: inst = 32'd268468224;
      51383: inst = 32'd201347075;
      51384: inst = 32'd203423744;
      51385: inst = 32'd471859200;
      51386: inst = 32'd136314880;
      51387: inst = 32'd268468224;
      51388: inst = 32'd201347076;
      51389: inst = 32'd203423744;
      51390: inst = 32'd471859200;
      51391: inst = 32'd136314880;
      51392: inst = 32'd268468224;
      51393: inst = 32'd201347077;
      51394: inst = 32'd203423744;
      51395: inst = 32'd471859200;
      51396: inst = 32'd136314880;
      51397: inst = 32'd268468224;
      51398: inst = 32'd201347078;
      51399: inst = 32'd203423744;
      51400: inst = 32'd471859200;
      51401: inst = 32'd136314880;
      51402: inst = 32'd268468224;
      51403: inst = 32'd201347079;
      51404: inst = 32'd203423744;
      51405: inst = 32'd471859200;
      51406: inst = 32'd136314880;
      51407: inst = 32'd268468224;
      51408: inst = 32'd201347080;
      51409: inst = 32'd203423744;
      51410: inst = 32'd471859200;
      51411: inst = 32'd136314880;
      51412: inst = 32'd268468224;
      51413: inst = 32'd201347081;
      51414: inst = 32'd203423744;
      51415: inst = 32'd471859200;
      51416: inst = 32'd136314880;
      51417: inst = 32'd268468224;
      51418: inst = 32'd201347082;
      51419: inst = 32'd203423744;
      51420: inst = 32'd471859200;
      51421: inst = 32'd136314880;
      51422: inst = 32'd268468224;
      51423: inst = 32'd201347083;
      51424: inst = 32'd203423744;
      51425: inst = 32'd471859200;
      51426: inst = 32'd136314880;
      51427: inst = 32'd268468224;
      51428: inst = 32'd201347084;
      51429: inst = 32'd203423744;
      51430: inst = 32'd471859200;
      51431: inst = 32'd136314880;
      51432: inst = 32'd268468224;
      51433: inst = 32'd201347085;
      51434: inst = 32'd203423744;
      51435: inst = 32'd471859200;
      51436: inst = 32'd136314880;
      51437: inst = 32'd268468224;
      51438: inst = 32'd201347086;
      51439: inst = 32'd203423744;
      51440: inst = 32'd471859200;
      51441: inst = 32'd136314880;
      51442: inst = 32'd268468224;
      51443: inst = 32'd201347087;
      51444: inst = 32'd203423744;
      51445: inst = 32'd471859200;
      51446: inst = 32'd136314880;
      51447: inst = 32'd268468224;
      51448: inst = 32'd201347088;
      51449: inst = 32'd203423744;
      51450: inst = 32'd471859200;
      51451: inst = 32'd136314880;
      51452: inst = 32'd268468224;
      51453: inst = 32'd201347089;
      51454: inst = 32'd203423744;
      51455: inst = 32'd471859200;
      51456: inst = 32'd136314880;
      51457: inst = 32'd268468224;
      51458: inst = 32'd201347090;
      51459: inst = 32'd203423744;
      51460: inst = 32'd471859200;
      51461: inst = 32'd136314880;
      51462: inst = 32'd268468224;
      51463: inst = 32'd201347091;
      51464: inst = 32'd203423744;
      51465: inst = 32'd471859200;
      51466: inst = 32'd136314880;
      51467: inst = 32'd268468224;
      51468: inst = 32'd201347092;
      51469: inst = 32'd203423744;
      51470: inst = 32'd471859200;
      51471: inst = 32'd136314880;
      51472: inst = 32'd268468224;
      51473: inst = 32'd201347093;
      51474: inst = 32'd203423744;
      51475: inst = 32'd471859200;
      51476: inst = 32'd136314880;
      51477: inst = 32'd268468224;
      51478: inst = 32'd201347094;
      51479: inst = 32'd203423744;
      51480: inst = 32'd471859200;
      51481: inst = 32'd136314880;
      51482: inst = 32'd268468224;
      51483: inst = 32'd201347095;
      51484: inst = 32'd203423744;
      51485: inst = 32'd471859200;
      51486: inst = 32'd136314880;
      51487: inst = 32'd268468224;
      51488: inst = 32'd201347096;
      51489: inst = 32'd203423744;
      51490: inst = 32'd471859200;
      51491: inst = 32'd136314880;
      51492: inst = 32'd268468224;
      51493: inst = 32'd201347097;
      51494: inst = 32'd203423744;
      51495: inst = 32'd471859200;
      51496: inst = 32'd136314880;
      51497: inst = 32'd268468224;
      51498: inst = 32'd201347098;
      51499: inst = 32'd203423744;
      51500: inst = 32'd471859200;
      51501: inst = 32'd136314880;
      51502: inst = 32'd268468224;
      51503: inst = 32'd201347099;
      51504: inst = 32'd203423744;
      51505: inst = 32'd471859200;
      51506: inst = 32'd136314880;
      51507: inst = 32'd268468224;
      51508: inst = 32'd201347100;
      51509: inst = 32'd203423744;
      51510: inst = 32'd471859200;
      51511: inst = 32'd136314880;
      51512: inst = 32'd268468224;
      51513: inst = 32'd201347101;
      51514: inst = 32'd203423744;
      51515: inst = 32'd471859200;
      51516: inst = 32'd136314880;
      51517: inst = 32'd268468224;
      51518: inst = 32'd201347102;
      51519: inst = 32'd203423744;
      51520: inst = 32'd471859200;
      51521: inst = 32'd136314880;
      51522: inst = 32'd268468224;
      51523: inst = 32'd201347103;
      51524: inst = 32'd203423744;
      51525: inst = 32'd471859200;
      51526: inst = 32'd136314880;
      51527: inst = 32'd268468224;
      51528: inst = 32'd201347104;
      51529: inst = 32'd203423744;
      51530: inst = 32'd471859200;
      51531: inst = 32'd136314880;
      51532: inst = 32'd268468224;
      51533: inst = 32'd201347105;
      51534: inst = 32'd203423744;
      51535: inst = 32'd471859200;
      51536: inst = 32'd136314880;
      51537: inst = 32'd268468224;
      51538: inst = 32'd201347106;
      51539: inst = 32'd203423744;
      51540: inst = 32'd471859200;
      51541: inst = 32'd136314880;
      51542: inst = 32'd268468224;
      51543: inst = 32'd201347107;
      51544: inst = 32'd203423744;
      51545: inst = 32'd471859200;
      51546: inst = 32'd136314880;
      51547: inst = 32'd268468224;
      51548: inst = 32'd201347108;
      51549: inst = 32'd203423744;
      51550: inst = 32'd471859200;
      51551: inst = 32'd136314880;
      51552: inst = 32'd268468224;
      51553: inst = 32'd201347109;
      51554: inst = 32'd203423744;
      51555: inst = 32'd471859200;
      51556: inst = 32'd136314880;
      51557: inst = 32'd268468224;
      51558: inst = 32'd201347110;
      51559: inst = 32'd203423744;
      51560: inst = 32'd471859200;
      51561: inst = 32'd136314880;
      51562: inst = 32'd268468224;
      51563: inst = 32'd201347111;
      51564: inst = 32'd203423744;
      51565: inst = 32'd471859200;
      51566: inst = 32'd136314880;
      51567: inst = 32'd268468224;
      51568: inst = 32'd201347112;
      51569: inst = 32'd203423744;
      51570: inst = 32'd471859200;
      51571: inst = 32'd136314880;
      51572: inst = 32'd268468224;
      51573: inst = 32'd201347113;
      51574: inst = 32'd203423744;
      51575: inst = 32'd471859200;
      51576: inst = 32'd136314880;
      51577: inst = 32'd268468224;
      51578: inst = 32'd201347114;
      51579: inst = 32'd203423744;
      51580: inst = 32'd471859200;
      51581: inst = 32'd136314880;
      51582: inst = 32'd268468224;
      51583: inst = 32'd201347115;
      51584: inst = 32'd203423744;
      51585: inst = 32'd471859200;
      51586: inst = 32'd136314880;
      51587: inst = 32'd268468224;
      51588: inst = 32'd201347116;
      51589: inst = 32'd203423744;
      51590: inst = 32'd471859200;
      51591: inst = 32'd136314880;
      51592: inst = 32'd268468224;
      51593: inst = 32'd201347117;
      51594: inst = 32'd203423744;
      51595: inst = 32'd471859200;
      51596: inst = 32'd136314880;
      51597: inst = 32'd268468224;
      51598: inst = 32'd201347118;
      51599: inst = 32'd203423744;
      51600: inst = 32'd471859200;
      51601: inst = 32'd136314880;
      51602: inst = 32'd268468224;
      51603: inst = 32'd201347119;
      51604: inst = 32'd203423744;
      51605: inst = 32'd471859200;
      51606: inst = 32'd136314880;
      51607: inst = 32'd268468224;
      51608: inst = 32'd201347120;
      51609: inst = 32'd203423744;
      51610: inst = 32'd471859200;
      51611: inst = 32'd136314880;
      51612: inst = 32'd268468224;
      51613: inst = 32'd201347121;
      51614: inst = 32'd203423744;
      51615: inst = 32'd471859200;
      51616: inst = 32'd136314880;
      51617: inst = 32'd268468224;
      51618: inst = 32'd201347122;
      51619: inst = 32'd203423744;
      51620: inst = 32'd471859200;
      51621: inst = 32'd136314880;
      51622: inst = 32'd268468224;
      51623: inst = 32'd201347123;
      51624: inst = 32'd203423744;
      51625: inst = 32'd471859200;
      51626: inst = 32'd136314880;
      51627: inst = 32'd268468224;
      51628: inst = 32'd201347124;
      51629: inst = 32'd203423744;
      51630: inst = 32'd471859200;
      51631: inst = 32'd136314880;
      51632: inst = 32'd268468224;
      51633: inst = 32'd201347125;
      51634: inst = 32'd203423744;
      51635: inst = 32'd471859200;
      51636: inst = 32'd136314880;
      51637: inst = 32'd268468224;
      51638: inst = 32'd201347126;
      51639: inst = 32'd203423744;
      51640: inst = 32'd471859200;
      51641: inst = 32'd136314880;
      51642: inst = 32'd268468224;
      51643: inst = 32'd201347127;
      51644: inst = 32'd203423744;
      51645: inst = 32'd471859200;
      51646: inst = 32'd136314880;
      51647: inst = 32'd268468224;
      51648: inst = 32'd201347128;
      51649: inst = 32'd203423744;
      51650: inst = 32'd471859200;
      51651: inst = 32'd136314880;
      51652: inst = 32'd268468224;
      51653: inst = 32'd201347129;
      51654: inst = 32'd203423744;
      51655: inst = 32'd471859200;
      51656: inst = 32'd136314880;
      51657: inst = 32'd268468224;
      51658: inst = 32'd201347130;
      51659: inst = 32'd203423744;
      51660: inst = 32'd471859200;
      51661: inst = 32'd136314880;
      51662: inst = 32'd268468224;
      51663: inst = 32'd201347131;
      51664: inst = 32'd203423744;
      51665: inst = 32'd471859200;
      51666: inst = 32'd136314880;
      51667: inst = 32'd268468224;
      51668: inst = 32'd201347132;
      51669: inst = 32'd203423744;
      51670: inst = 32'd471859200;
      51671: inst = 32'd136314880;
      51672: inst = 32'd268468224;
      51673: inst = 32'd201347133;
      51674: inst = 32'd203423744;
      51675: inst = 32'd471859200;
      51676: inst = 32'd136314880;
      51677: inst = 32'd268468224;
      51678: inst = 32'd201347134;
      51679: inst = 32'd203423744;
      51680: inst = 32'd471859200;
      51681: inst = 32'd136314880;
      51682: inst = 32'd268468224;
      51683: inst = 32'd201347135;
      51684: inst = 32'd203423744;
      51685: inst = 32'd471859200;
      51686: inst = 32'd136314880;
      51687: inst = 32'd268468224;
      51688: inst = 32'd201347136;
      51689: inst = 32'd203423744;
      51690: inst = 32'd471859200;
      51691: inst = 32'd136314880;
      51692: inst = 32'd268468224;
      51693: inst = 32'd201347137;
      51694: inst = 32'd203423744;
      51695: inst = 32'd471859200;
      51696: inst = 32'd136314880;
      51697: inst = 32'd268468224;
      51698: inst = 32'd201347138;
      51699: inst = 32'd203423744;
      51700: inst = 32'd471859200;
      51701: inst = 32'd136314880;
      51702: inst = 32'd268468224;
      51703: inst = 32'd201347139;
      51704: inst = 32'd203423744;
      51705: inst = 32'd471859200;
      51706: inst = 32'd136314880;
      51707: inst = 32'd268468224;
      51708: inst = 32'd201347140;
      51709: inst = 32'd203423744;
      51710: inst = 32'd471859200;
      51711: inst = 32'd136314880;
      51712: inst = 32'd268468224;
      51713: inst = 32'd201347141;
      51714: inst = 32'd203423744;
      51715: inst = 32'd471859200;
      51716: inst = 32'd136314880;
      51717: inst = 32'd268468224;
      51718: inst = 32'd201347142;
      51719: inst = 32'd203423744;
      51720: inst = 32'd471859200;
      51721: inst = 32'd136314880;
      51722: inst = 32'd268468224;
      51723: inst = 32'd201347143;
      51724: inst = 32'd203423744;
      51725: inst = 32'd471859200;
      51726: inst = 32'd136314880;
      51727: inst = 32'd268468224;
      51728: inst = 32'd201347144;
      51729: inst = 32'd203423744;
      51730: inst = 32'd471859200;
      51731: inst = 32'd136314880;
      51732: inst = 32'd268468224;
      51733: inst = 32'd201347145;
      51734: inst = 32'd203423744;
      51735: inst = 32'd471859200;
      51736: inst = 32'd136314880;
      51737: inst = 32'd268468224;
      51738: inst = 32'd201347146;
      51739: inst = 32'd203423744;
      51740: inst = 32'd471859200;
      51741: inst = 32'd136314880;
      51742: inst = 32'd268468224;
      51743: inst = 32'd201347147;
      51744: inst = 32'd203423744;
      51745: inst = 32'd471859200;
      51746: inst = 32'd136314880;
      51747: inst = 32'd268468224;
      51748: inst = 32'd201347148;
      51749: inst = 32'd203423744;
      51750: inst = 32'd471859200;
      51751: inst = 32'd136314880;
      51752: inst = 32'd268468224;
      51753: inst = 32'd201347149;
      51754: inst = 32'd203423744;
      51755: inst = 32'd471859200;
      51756: inst = 32'd136314880;
      51757: inst = 32'd268468224;
      51758: inst = 32'd201347150;
      51759: inst = 32'd203423744;
      51760: inst = 32'd471859200;
      51761: inst = 32'd136314880;
      51762: inst = 32'd268468224;
      51763: inst = 32'd201347151;
      51764: inst = 32'd203423744;
      51765: inst = 32'd471859200;
      51766: inst = 32'd136314880;
      51767: inst = 32'd268468224;
      51768: inst = 32'd201347152;
      51769: inst = 32'd203423744;
      51770: inst = 32'd471859200;
      51771: inst = 32'd136314880;
      51772: inst = 32'd268468224;
      51773: inst = 32'd201347153;
      51774: inst = 32'd203423744;
      51775: inst = 32'd471859200;
      51776: inst = 32'd136314880;
      51777: inst = 32'd268468224;
      51778: inst = 32'd201347154;
      51779: inst = 32'd203423744;
      51780: inst = 32'd471859200;
      51781: inst = 32'd136314880;
      51782: inst = 32'd268468224;
      51783: inst = 32'd201347155;
      51784: inst = 32'd203423744;
      51785: inst = 32'd471859200;
      51786: inst = 32'd136314880;
      51787: inst = 32'd268468224;
      51788: inst = 32'd201347156;
      51789: inst = 32'd203423744;
      51790: inst = 32'd471859200;
      51791: inst = 32'd136314880;
      51792: inst = 32'd268468224;
      51793: inst = 32'd201347157;
      51794: inst = 32'd203423744;
      51795: inst = 32'd471859200;
      51796: inst = 32'd136314880;
      51797: inst = 32'd268468224;
      51798: inst = 32'd201347158;
      51799: inst = 32'd203423744;
      51800: inst = 32'd471859200;
      51801: inst = 32'd136314880;
      51802: inst = 32'd268468224;
      51803: inst = 32'd201347159;
      51804: inst = 32'd203423744;
      51805: inst = 32'd471859200;
      51806: inst = 32'd136314880;
      51807: inst = 32'd268468224;
      51808: inst = 32'd201347160;
      51809: inst = 32'd203423744;
      51810: inst = 32'd471859200;
      51811: inst = 32'd136314880;
      51812: inst = 32'd268468224;
      51813: inst = 32'd201347161;
      51814: inst = 32'd203423744;
      51815: inst = 32'd471859200;
      51816: inst = 32'd136314880;
      51817: inst = 32'd268468224;
      51818: inst = 32'd201347162;
      51819: inst = 32'd203423744;
      51820: inst = 32'd471859200;
      51821: inst = 32'd136314880;
      51822: inst = 32'd268468224;
      51823: inst = 32'd201347163;
      51824: inst = 32'd203423744;
      51825: inst = 32'd471859200;
      51826: inst = 32'd136314880;
      51827: inst = 32'd268468224;
      51828: inst = 32'd201347164;
      51829: inst = 32'd203423744;
      51830: inst = 32'd471859200;
      51831: inst = 32'd136314880;
      51832: inst = 32'd268468224;
      51833: inst = 32'd201347165;
      51834: inst = 32'd203423744;
      51835: inst = 32'd471859200;
      51836: inst = 32'd136314880;
      51837: inst = 32'd268468224;
      51838: inst = 32'd201347166;
      51839: inst = 32'd203423744;
      51840: inst = 32'd471859200;
      51841: inst = 32'd136314880;
      51842: inst = 32'd268468224;
      51843: inst = 32'd201347167;
      51844: inst = 32'd203423744;
      51845: inst = 32'd471859200;
      51846: inst = 32'd136314880;
      51847: inst = 32'd268468224;
      51848: inst = 32'd201347168;
      51849: inst = 32'd203423744;
      51850: inst = 32'd471859200;
      51851: inst = 32'd136314880;
      51852: inst = 32'd268468224;
      51853: inst = 32'd201347169;
      51854: inst = 32'd203423744;
      51855: inst = 32'd471859200;
      51856: inst = 32'd136314880;
      51857: inst = 32'd268468224;
      51858: inst = 32'd201347170;
      51859: inst = 32'd203423744;
      51860: inst = 32'd471859200;
      51861: inst = 32'd136314880;
      51862: inst = 32'd268468224;
      51863: inst = 32'd201347171;
      51864: inst = 32'd203423744;
      51865: inst = 32'd471859200;
      51866: inst = 32'd136314880;
      51867: inst = 32'd268468224;
      51868: inst = 32'd201347172;
      51869: inst = 32'd203423744;
      51870: inst = 32'd471859200;
      51871: inst = 32'd136314880;
      51872: inst = 32'd268468224;
      51873: inst = 32'd201347173;
      51874: inst = 32'd203423744;
      51875: inst = 32'd471859200;
      51876: inst = 32'd136314880;
      51877: inst = 32'd268468224;
      51878: inst = 32'd201347174;
      51879: inst = 32'd203423744;
      51880: inst = 32'd471859200;
      51881: inst = 32'd136314880;
      51882: inst = 32'd268468224;
      51883: inst = 32'd201347175;
      51884: inst = 32'd203423744;
      51885: inst = 32'd471859200;
      51886: inst = 32'd136314880;
      51887: inst = 32'd268468224;
      51888: inst = 32'd201347176;
      51889: inst = 32'd203423744;
      51890: inst = 32'd471859200;
      51891: inst = 32'd136314880;
      51892: inst = 32'd268468224;
      51893: inst = 32'd201347177;
      51894: inst = 32'd203423744;
      51895: inst = 32'd471859200;
      51896: inst = 32'd136314880;
      51897: inst = 32'd268468224;
      51898: inst = 32'd201347178;
      51899: inst = 32'd203423744;
      51900: inst = 32'd471859200;
      51901: inst = 32'd136314880;
      51902: inst = 32'd268468224;
      51903: inst = 32'd201347179;
      51904: inst = 32'd203423744;
      51905: inst = 32'd471859200;
      51906: inst = 32'd136314880;
      51907: inst = 32'd268468224;
      51908: inst = 32'd201347180;
      51909: inst = 32'd203423744;
      51910: inst = 32'd471859200;
      51911: inst = 32'd136314880;
      51912: inst = 32'd268468224;
      51913: inst = 32'd201347181;
      51914: inst = 32'd203423744;
      51915: inst = 32'd471859200;
      51916: inst = 32'd136314880;
      51917: inst = 32'd268468224;
      51918: inst = 32'd201347182;
      51919: inst = 32'd203423744;
      51920: inst = 32'd471859200;
      51921: inst = 32'd136314880;
      51922: inst = 32'd268468224;
      51923: inst = 32'd201347183;
      51924: inst = 32'd203423744;
      51925: inst = 32'd471859200;
      51926: inst = 32'd136314880;
      51927: inst = 32'd268468224;
      51928: inst = 32'd201347184;
      51929: inst = 32'd203423744;
      51930: inst = 32'd471859200;
      51931: inst = 32'd136314880;
      51932: inst = 32'd268468224;
      51933: inst = 32'd201347185;
      51934: inst = 32'd203423744;
      51935: inst = 32'd471859200;
      51936: inst = 32'd136314880;
      51937: inst = 32'd268468224;
      51938: inst = 32'd201347186;
      51939: inst = 32'd203423744;
      51940: inst = 32'd471859200;
      51941: inst = 32'd136314880;
      51942: inst = 32'd268468224;
      51943: inst = 32'd201347187;
      51944: inst = 32'd203423744;
      51945: inst = 32'd471859200;
      51946: inst = 32'd136314880;
      51947: inst = 32'd268468224;
      51948: inst = 32'd201347188;
      51949: inst = 32'd203423744;
      51950: inst = 32'd471859200;
      51951: inst = 32'd136314880;
      51952: inst = 32'd268468224;
      51953: inst = 32'd201347189;
      51954: inst = 32'd203423744;
      51955: inst = 32'd471859200;
      51956: inst = 32'd136314880;
      51957: inst = 32'd268468224;
      51958: inst = 32'd201347190;
      51959: inst = 32'd203423744;
      51960: inst = 32'd471859200;
      51961: inst = 32'd136314880;
      51962: inst = 32'd268468224;
      51963: inst = 32'd201347191;
      51964: inst = 32'd203423744;
      51965: inst = 32'd471859200;
      51966: inst = 32'd136314880;
      51967: inst = 32'd268468224;
      51968: inst = 32'd201347192;
      51969: inst = 32'd203423744;
      51970: inst = 32'd471859200;
      51971: inst = 32'd136314880;
      51972: inst = 32'd268468224;
      51973: inst = 32'd201347193;
      51974: inst = 32'd203423744;
      51975: inst = 32'd471859200;
      51976: inst = 32'd136314880;
      51977: inst = 32'd268468224;
      51978: inst = 32'd201347194;
      51979: inst = 32'd203423744;
      51980: inst = 32'd471859200;
      51981: inst = 32'd136314880;
      51982: inst = 32'd268468224;
      51983: inst = 32'd201347195;
      51984: inst = 32'd203423744;
      51985: inst = 32'd471859200;
      51986: inst = 32'd136314880;
      51987: inst = 32'd268468224;
      51988: inst = 32'd201347196;
      51989: inst = 32'd203423744;
      51990: inst = 32'd471859200;
      51991: inst = 32'd136314880;
      51992: inst = 32'd268468224;
      51993: inst = 32'd201347197;
      51994: inst = 32'd203423744;
      51995: inst = 32'd471859200;
      51996: inst = 32'd136314880;
      51997: inst = 32'd268468224;
      51998: inst = 32'd201347198;
      51999: inst = 32'd203423744;
      52000: inst = 32'd471859200;
      52001: inst = 32'd136314880;
      52002: inst = 32'd268468224;
      52003: inst = 32'd201347199;
      52004: inst = 32'd203423744;
      52005: inst = 32'd471859200;
      52006: inst = 32'd136314880;
      52007: inst = 32'd268468224;
      52008: inst = 32'd201347200;
      52009: inst = 32'd203423744;
      52010: inst = 32'd471859200;
      52011: inst = 32'd136314880;
      52012: inst = 32'd268468224;
      52013: inst = 32'd201347201;
      52014: inst = 32'd203423744;
      52015: inst = 32'd471859200;
      52016: inst = 32'd136314880;
      52017: inst = 32'd268468224;
      52018: inst = 32'd201347202;
      52019: inst = 32'd203423744;
      52020: inst = 32'd471859200;
      52021: inst = 32'd136314880;
      52022: inst = 32'd268468224;
      52023: inst = 32'd201347203;
      52024: inst = 32'd203423744;
      52025: inst = 32'd471859200;
      52026: inst = 32'd136314880;
      52027: inst = 32'd268468224;
      52028: inst = 32'd201347204;
      52029: inst = 32'd203423744;
      52030: inst = 32'd471859200;
      52031: inst = 32'd136314880;
      52032: inst = 32'd268468224;
      52033: inst = 32'd201347205;
      52034: inst = 32'd203423744;
      52035: inst = 32'd471859200;
      52036: inst = 32'd136314880;
      52037: inst = 32'd268468224;
      52038: inst = 32'd201347206;
      52039: inst = 32'd203423744;
      52040: inst = 32'd471859200;
      52041: inst = 32'd136314880;
      52042: inst = 32'd268468224;
      52043: inst = 32'd201347207;
      52044: inst = 32'd203423744;
      52045: inst = 32'd471859200;
      52046: inst = 32'd136314880;
      52047: inst = 32'd268468224;
      52048: inst = 32'd201347208;
      52049: inst = 32'd203423744;
      52050: inst = 32'd471859200;
      52051: inst = 32'd136314880;
      52052: inst = 32'd268468224;
      52053: inst = 32'd201347209;
      52054: inst = 32'd203423744;
      52055: inst = 32'd471859200;
      52056: inst = 32'd136314880;
      52057: inst = 32'd268468224;
      52058: inst = 32'd201347210;
      52059: inst = 32'd203423744;
      52060: inst = 32'd471859200;
      52061: inst = 32'd136314880;
      52062: inst = 32'd268468224;
      52063: inst = 32'd201347211;
      52064: inst = 32'd203423744;
      52065: inst = 32'd471859200;
      52066: inst = 32'd136314880;
      52067: inst = 32'd268468224;
      52068: inst = 32'd201347212;
      52069: inst = 32'd203423744;
      52070: inst = 32'd471859200;
      52071: inst = 32'd136314880;
      52072: inst = 32'd268468224;
      52073: inst = 32'd201347213;
      52074: inst = 32'd203423744;
      52075: inst = 32'd471859200;
      52076: inst = 32'd136314880;
      52077: inst = 32'd268468224;
      52078: inst = 32'd201347214;
      52079: inst = 32'd203423744;
      52080: inst = 32'd471859200;
      52081: inst = 32'd136314880;
      52082: inst = 32'd268468224;
      52083: inst = 32'd201347215;
      52084: inst = 32'd203423744;
      52085: inst = 32'd471859200;
      52086: inst = 32'd136314880;
      52087: inst = 32'd268468224;
      52088: inst = 32'd201347216;
      52089: inst = 32'd203423744;
      52090: inst = 32'd471859200;
      52091: inst = 32'd136314880;
      52092: inst = 32'd268468224;
      52093: inst = 32'd201347217;
      52094: inst = 32'd203423744;
      52095: inst = 32'd471859200;
      52096: inst = 32'd136314880;
      52097: inst = 32'd268468224;
      52098: inst = 32'd201347218;
      52099: inst = 32'd203423744;
      52100: inst = 32'd471859200;
      52101: inst = 32'd136314880;
      52102: inst = 32'd268468224;
      52103: inst = 32'd201347219;
      52104: inst = 32'd203423744;
      52105: inst = 32'd471859200;
      52106: inst = 32'd136314880;
      52107: inst = 32'd268468224;
      52108: inst = 32'd201347220;
      52109: inst = 32'd203423744;
      52110: inst = 32'd471859200;
      52111: inst = 32'd136314880;
      52112: inst = 32'd268468224;
      52113: inst = 32'd201347221;
      52114: inst = 32'd203423744;
      52115: inst = 32'd471859200;
      52116: inst = 32'd136314880;
      52117: inst = 32'd268468224;
      52118: inst = 32'd201347222;
      52119: inst = 32'd203423744;
      52120: inst = 32'd471859200;
      52121: inst = 32'd136314880;
      52122: inst = 32'd268468224;
      52123: inst = 32'd201347223;
      52124: inst = 32'd203423744;
      52125: inst = 32'd471859200;
      52126: inst = 32'd136314880;
      52127: inst = 32'd268468224;
      52128: inst = 32'd201347224;
      52129: inst = 32'd203423744;
      52130: inst = 32'd471859200;
      52131: inst = 32'd136314880;
      52132: inst = 32'd268468224;
      52133: inst = 32'd201347225;
      52134: inst = 32'd203423744;
      52135: inst = 32'd471859200;
      52136: inst = 32'd136314880;
      52137: inst = 32'd268468224;
      52138: inst = 32'd201347226;
      52139: inst = 32'd203423744;
      52140: inst = 32'd471859200;
      52141: inst = 32'd136314880;
      52142: inst = 32'd268468224;
      52143: inst = 32'd201347227;
      52144: inst = 32'd203423744;
      52145: inst = 32'd471859200;
      52146: inst = 32'd136314880;
      52147: inst = 32'd268468224;
      52148: inst = 32'd201347228;
      52149: inst = 32'd203423744;
      52150: inst = 32'd471859200;
      52151: inst = 32'd136314880;
      52152: inst = 32'd268468224;
      52153: inst = 32'd201347229;
      52154: inst = 32'd203423744;
      52155: inst = 32'd471859200;
      52156: inst = 32'd136314880;
      52157: inst = 32'd268468224;
      52158: inst = 32'd201347230;
      52159: inst = 32'd203423744;
      52160: inst = 32'd471859200;
      52161: inst = 32'd136314880;
      52162: inst = 32'd268468224;
      52163: inst = 32'd201347231;
      52164: inst = 32'd203423744;
      52165: inst = 32'd471859200;
      52166: inst = 32'd136314880;
      52167: inst = 32'd268468224;
      52168: inst = 32'd201347232;
      52169: inst = 32'd203423744;
      52170: inst = 32'd471859200;
      52171: inst = 32'd136314880;
      52172: inst = 32'd268468224;
      52173: inst = 32'd201347233;
      52174: inst = 32'd203423744;
      52175: inst = 32'd471859200;
      52176: inst = 32'd136314880;
      52177: inst = 32'd268468224;
      52178: inst = 32'd201347234;
      52179: inst = 32'd203423744;
      52180: inst = 32'd471859200;
      52181: inst = 32'd136314880;
      52182: inst = 32'd268468224;
      52183: inst = 32'd201347235;
      52184: inst = 32'd203423744;
      52185: inst = 32'd471859200;
      52186: inst = 32'd136314880;
      52187: inst = 32'd268468224;
      52188: inst = 32'd201347236;
      52189: inst = 32'd203423744;
      52190: inst = 32'd471859200;
      52191: inst = 32'd136314880;
      52192: inst = 32'd268468224;
      52193: inst = 32'd201347237;
      52194: inst = 32'd203423744;
      52195: inst = 32'd471859200;
      52196: inst = 32'd136314880;
      52197: inst = 32'd268468224;
      52198: inst = 32'd201347238;
      52199: inst = 32'd203423744;
      52200: inst = 32'd471859200;
      52201: inst = 32'd136314880;
      52202: inst = 32'd268468224;
      52203: inst = 32'd201347239;
      52204: inst = 32'd203423744;
      52205: inst = 32'd471859200;
      52206: inst = 32'd136314880;
      52207: inst = 32'd268468224;
      52208: inst = 32'd201347240;
      52209: inst = 32'd203423744;
      52210: inst = 32'd471859200;
      52211: inst = 32'd136314880;
      52212: inst = 32'd268468224;
      52213: inst = 32'd201347241;
      52214: inst = 32'd203423744;
      52215: inst = 32'd471859200;
      52216: inst = 32'd136314880;
      52217: inst = 32'd268468224;
      52218: inst = 32'd201347242;
      52219: inst = 32'd203423744;
      52220: inst = 32'd471859200;
      52221: inst = 32'd136314880;
      52222: inst = 32'd268468224;
      52223: inst = 32'd201347243;
      52224: inst = 32'd203423744;
      52225: inst = 32'd471859200;
      52226: inst = 32'd136314880;
      52227: inst = 32'd268468224;
      52228: inst = 32'd201347244;
      52229: inst = 32'd203423744;
      52230: inst = 32'd471859200;
      52231: inst = 32'd136314880;
      52232: inst = 32'd268468224;
      52233: inst = 32'd201347245;
      52234: inst = 32'd203423744;
      52235: inst = 32'd471859200;
      52236: inst = 32'd136314880;
      52237: inst = 32'd268468224;
      52238: inst = 32'd201347246;
      52239: inst = 32'd203423744;
      52240: inst = 32'd471859200;
      52241: inst = 32'd136314880;
      52242: inst = 32'd268468224;
      52243: inst = 32'd201347247;
      52244: inst = 32'd203423744;
      52245: inst = 32'd471859200;
      52246: inst = 32'd136314880;
      52247: inst = 32'd268468224;
      52248: inst = 32'd201347248;
      52249: inst = 32'd203423744;
      52250: inst = 32'd471859200;
      52251: inst = 32'd136314880;
      52252: inst = 32'd268468224;
      52253: inst = 32'd201347249;
      52254: inst = 32'd203423744;
      52255: inst = 32'd471859200;
      52256: inst = 32'd136314880;
      52257: inst = 32'd268468224;
      52258: inst = 32'd201347250;
      52259: inst = 32'd203423744;
      52260: inst = 32'd471859200;
      52261: inst = 32'd136314880;
      52262: inst = 32'd268468224;
      52263: inst = 32'd201347251;
      52264: inst = 32'd203423744;
      52265: inst = 32'd471859200;
      52266: inst = 32'd136314880;
      52267: inst = 32'd268468224;
      52268: inst = 32'd201347252;
      52269: inst = 32'd203423744;
      52270: inst = 32'd471859200;
      52271: inst = 32'd136314880;
      52272: inst = 32'd268468224;
      52273: inst = 32'd201347253;
      52274: inst = 32'd203423744;
      52275: inst = 32'd471859200;
      52276: inst = 32'd136314880;
      52277: inst = 32'd268468224;
      52278: inst = 32'd201347254;
      52279: inst = 32'd203423744;
      52280: inst = 32'd471859200;
      52281: inst = 32'd136314880;
      52282: inst = 32'd268468224;
      52283: inst = 32'd201347255;
      52284: inst = 32'd203423744;
      52285: inst = 32'd471859200;
      52286: inst = 32'd136314880;
      52287: inst = 32'd268468224;
      52288: inst = 32'd201347256;
      52289: inst = 32'd203423744;
      52290: inst = 32'd471859200;
      52291: inst = 32'd136314880;
      52292: inst = 32'd268468224;
      52293: inst = 32'd201347257;
      52294: inst = 32'd203423744;
      52295: inst = 32'd471859200;
      52296: inst = 32'd136314880;
      52297: inst = 32'd268468224;
      52298: inst = 32'd201347258;
      52299: inst = 32'd203423744;
      52300: inst = 32'd471859200;
      52301: inst = 32'd136314880;
      52302: inst = 32'd268468224;
      52303: inst = 32'd201347259;
      52304: inst = 32'd203423744;
      52305: inst = 32'd471859200;
      52306: inst = 32'd136314880;
      52307: inst = 32'd268468224;
      52308: inst = 32'd201347260;
      52309: inst = 32'd203423744;
      52310: inst = 32'd471859200;
      52311: inst = 32'd136314880;
      52312: inst = 32'd268468224;
      52313: inst = 32'd201347261;
      52314: inst = 32'd203423744;
      52315: inst = 32'd471859200;
      52316: inst = 32'd136314880;
      52317: inst = 32'd268468224;
      52318: inst = 32'd201347262;
      52319: inst = 32'd203423744;
      52320: inst = 32'd471859200;
      52321: inst = 32'd136314880;
      52322: inst = 32'd268468224;
      52323: inst = 32'd201347263;
      52324: inst = 32'd203423744;
      52325: inst = 32'd471859200;
      52326: inst = 32'd136314880;
      52327: inst = 32'd268468224;
      52328: inst = 32'd201347264;
      52329: inst = 32'd203423744;
      52330: inst = 32'd471859200;
      52331: inst = 32'd136314880;
      52332: inst = 32'd268468224;
      52333: inst = 32'd201347265;
      52334: inst = 32'd203423744;
      52335: inst = 32'd471859200;
      52336: inst = 32'd136314880;
      52337: inst = 32'd268468224;
      52338: inst = 32'd201347266;
      52339: inst = 32'd203423744;
      52340: inst = 32'd471859200;
      52341: inst = 32'd136314880;
      52342: inst = 32'd268468224;
      52343: inst = 32'd201347267;
      52344: inst = 32'd203423744;
      52345: inst = 32'd471859200;
      52346: inst = 32'd136314880;
      52347: inst = 32'd268468224;
      52348: inst = 32'd201347268;
      52349: inst = 32'd203423744;
      52350: inst = 32'd471859200;
      52351: inst = 32'd136314880;
      52352: inst = 32'd268468224;
      52353: inst = 32'd201347269;
      52354: inst = 32'd203423744;
      52355: inst = 32'd471859200;
      52356: inst = 32'd136314880;
      52357: inst = 32'd268468224;
      52358: inst = 32'd201347270;
      52359: inst = 32'd203423744;
      52360: inst = 32'd471859200;
      52361: inst = 32'd136314880;
      52362: inst = 32'd268468224;
      52363: inst = 32'd201347271;
      52364: inst = 32'd203423744;
      52365: inst = 32'd471859200;
      52366: inst = 32'd136314880;
      52367: inst = 32'd268468224;
      52368: inst = 32'd201347272;
      52369: inst = 32'd203423744;
      52370: inst = 32'd471859200;
      52371: inst = 32'd136314880;
      52372: inst = 32'd268468224;
      52373: inst = 32'd201347273;
      52374: inst = 32'd203423744;
      52375: inst = 32'd471859200;
      52376: inst = 32'd136314880;
      52377: inst = 32'd268468224;
      52378: inst = 32'd201347274;
      52379: inst = 32'd203423744;
      52380: inst = 32'd471859200;
      52381: inst = 32'd136314880;
      52382: inst = 32'd268468224;
      52383: inst = 32'd201347275;
      52384: inst = 32'd203423744;
      52385: inst = 32'd471859200;
      52386: inst = 32'd136314880;
      52387: inst = 32'd268468224;
      52388: inst = 32'd201347276;
      52389: inst = 32'd203423744;
      52390: inst = 32'd471859200;
      52391: inst = 32'd136314880;
      52392: inst = 32'd268468224;
      52393: inst = 32'd201347277;
      52394: inst = 32'd203423744;
      52395: inst = 32'd471859200;
      52396: inst = 32'd136314880;
      52397: inst = 32'd268468224;
      52398: inst = 32'd201347278;
      52399: inst = 32'd203423744;
      52400: inst = 32'd471859200;
      52401: inst = 32'd136314880;
      52402: inst = 32'd268468224;
      52403: inst = 32'd201347279;
      52404: inst = 32'd203423744;
      52405: inst = 32'd471859200;
      52406: inst = 32'd136314880;
      52407: inst = 32'd268468224;
      52408: inst = 32'd201347280;
      52409: inst = 32'd203423744;
      52410: inst = 32'd471859200;
      52411: inst = 32'd136314880;
      52412: inst = 32'd268468224;
      52413: inst = 32'd201347281;
      52414: inst = 32'd203423744;
      52415: inst = 32'd471859200;
      52416: inst = 32'd136314880;
      52417: inst = 32'd268468224;
      52418: inst = 32'd201347282;
      52419: inst = 32'd203423744;
      52420: inst = 32'd471859200;
      52421: inst = 32'd136314880;
      52422: inst = 32'd268468224;
      52423: inst = 32'd201347283;
      52424: inst = 32'd203423744;
      52425: inst = 32'd471859200;
      52426: inst = 32'd136314880;
      52427: inst = 32'd268468224;
      52428: inst = 32'd201347284;
      52429: inst = 32'd203423744;
      52430: inst = 32'd471859200;
      52431: inst = 32'd136314880;
      52432: inst = 32'd268468224;
      52433: inst = 32'd201347285;
      52434: inst = 32'd203423744;
      52435: inst = 32'd471859200;
      52436: inst = 32'd136314880;
      52437: inst = 32'd268468224;
      52438: inst = 32'd201347286;
      52439: inst = 32'd203423744;
      52440: inst = 32'd471859200;
      52441: inst = 32'd136314880;
      52442: inst = 32'd268468224;
      52443: inst = 32'd201347287;
      52444: inst = 32'd203423744;
      52445: inst = 32'd471859200;
      52446: inst = 32'd136314880;
      52447: inst = 32'd268468224;
      52448: inst = 32'd201347288;
      52449: inst = 32'd203423744;
      52450: inst = 32'd471859200;
      52451: inst = 32'd136314880;
      52452: inst = 32'd268468224;
      52453: inst = 32'd201347289;
      52454: inst = 32'd203423744;
      52455: inst = 32'd471859200;
      52456: inst = 32'd136314880;
      52457: inst = 32'd268468224;
      52458: inst = 32'd201347290;
      52459: inst = 32'd203423744;
      52460: inst = 32'd471859200;
      52461: inst = 32'd136314880;
      52462: inst = 32'd268468224;
      52463: inst = 32'd201347291;
      52464: inst = 32'd203423744;
      52465: inst = 32'd471859200;
      52466: inst = 32'd136314880;
      52467: inst = 32'd268468224;
      52468: inst = 32'd201347292;
      52469: inst = 32'd203423744;
      52470: inst = 32'd471859200;
      52471: inst = 32'd136314880;
      52472: inst = 32'd268468224;
      52473: inst = 32'd201347293;
      52474: inst = 32'd203423744;
      52475: inst = 32'd471859200;
      52476: inst = 32'd136314880;
      52477: inst = 32'd268468224;
      52478: inst = 32'd201347294;
      52479: inst = 32'd203423744;
      52480: inst = 32'd471859200;
      52481: inst = 32'd136314880;
      52482: inst = 32'd268468224;
      52483: inst = 32'd201347295;
      52484: inst = 32'd203423744;
      52485: inst = 32'd471859200;
      52486: inst = 32'd136314880;
      52487: inst = 32'd268468224;
      52488: inst = 32'd201347296;
      52489: inst = 32'd203423744;
      52490: inst = 32'd471859200;
      52491: inst = 32'd136314880;
      52492: inst = 32'd268468224;
      52493: inst = 32'd201347297;
      52494: inst = 32'd203423744;
      52495: inst = 32'd471859200;
      52496: inst = 32'd136314880;
      52497: inst = 32'd268468224;
      52498: inst = 32'd201347298;
      52499: inst = 32'd203423744;
      52500: inst = 32'd471859200;
      52501: inst = 32'd136314880;
      52502: inst = 32'd268468224;
      52503: inst = 32'd201347299;
      52504: inst = 32'd203423744;
      52505: inst = 32'd471859200;
      52506: inst = 32'd136314880;
      52507: inst = 32'd268468224;
      52508: inst = 32'd201347300;
      52509: inst = 32'd203423744;
      52510: inst = 32'd471859200;
      52511: inst = 32'd136314880;
      52512: inst = 32'd268468224;
      52513: inst = 32'd201347301;
      52514: inst = 32'd203423744;
      52515: inst = 32'd471859200;
      52516: inst = 32'd136314880;
      52517: inst = 32'd268468224;
      52518: inst = 32'd201347302;
      52519: inst = 32'd203423744;
      52520: inst = 32'd471859200;
      52521: inst = 32'd136314880;
      52522: inst = 32'd268468224;
      52523: inst = 32'd201347303;
      52524: inst = 32'd203423744;
      52525: inst = 32'd471859200;
      52526: inst = 32'd136314880;
      52527: inst = 32'd268468224;
      52528: inst = 32'd201347304;
      52529: inst = 32'd203423744;
      52530: inst = 32'd471859200;
      52531: inst = 32'd136314880;
      52532: inst = 32'd268468224;
      52533: inst = 32'd201347305;
      52534: inst = 32'd203423744;
      52535: inst = 32'd471859200;
      52536: inst = 32'd136314880;
      52537: inst = 32'd268468224;
      52538: inst = 32'd201347306;
      52539: inst = 32'd203423744;
      52540: inst = 32'd471859200;
      52541: inst = 32'd136314880;
      52542: inst = 32'd268468224;
      52543: inst = 32'd201347307;
      52544: inst = 32'd203423744;
      52545: inst = 32'd471859200;
      52546: inst = 32'd136314880;
      52547: inst = 32'd268468224;
      52548: inst = 32'd201347308;
      52549: inst = 32'd203423744;
      52550: inst = 32'd471859200;
      52551: inst = 32'd136314880;
      52552: inst = 32'd268468224;
      52553: inst = 32'd201347309;
      52554: inst = 32'd203423744;
      52555: inst = 32'd471859200;
      52556: inst = 32'd136314880;
      52557: inst = 32'd268468224;
      52558: inst = 32'd201347310;
      52559: inst = 32'd203423744;
      52560: inst = 32'd471859200;
      52561: inst = 32'd136314880;
      52562: inst = 32'd268468224;
      52563: inst = 32'd201347311;
      52564: inst = 32'd203423744;
      52565: inst = 32'd471859200;
      52566: inst = 32'd136314880;
      52567: inst = 32'd268468224;
      52568: inst = 32'd201347312;
      52569: inst = 32'd203423744;
      52570: inst = 32'd471859200;
      52571: inst = 32'd136314880;
      52572: inst = 32'd268468224;
      52573: inst = 32'd201347313;
      52574: inst = 32'd203423744;
      52575: inst = 32'd471859200;
      52576: inst = 32'd136314880;
      52577: inst = 32'd268468224;
      52578: inst = 32'd201347314;
      52579: inst = 32'd203423744;
      52580: inst = 32'd471859200;
      52581: inst = 32'd136314880;
      52582: inst = 32'd268468224;
      52583: inst = 32'd201347315;
      52584: inst = 32'd203423744;
      52585: inst = 32'd471859200;
      52586: inst = 32'd136314880;
      52587: inst = 32'd268468224;
      52588: inst = 32'd201347316;
      52589: inst = 32'd203423744;
      52590: inst = 32'd471859200;
      52591: inst = 32'd136314880;
      52592: inst = 32'd268468224;
      52593: inst = 32'd201347317;
      52594: inst = 32'd203423744;
      52595: inst = 32'd471859200;
      52596: inst = 32'd136314880;
      52597: inst = 32'd268468224;
      52598: inst = 32'd201347318;
      52599: inst = 32'd203423744;
      52600: inst = 32'd471859200;
      52601: inst = 32'd136314880;
      52602: inst = 32'd268468224;
      52603: inst = 32'd201347319;
      52604: inst = 32'd203423744;
      52605: inst = 32'd471859200;
      52606: inst = 32'd136314880;
      52607: inst = 32'd268468224;
      52608: inst = 32'd201347320;
      52609: inst = 32'd203423744;
      52610: inst = 32'd471859200;
      52611: inst = 32'd136314880;
      52612: inst = 32'd268468224;
      52613: inst = 32'd201347321;
      52614: inst = 32'd203423744;
      52615: inst = 32'd471859200;
      52616: inst = 32'd136314880;
      52617: inst = 32'd268468224;
      52618: inst = 32'd201347322;
      52619: inst = 32'd203423744;
      52620: inst = 32'd471859200;
      52621: inst = 32'd136314880;
      52622: inst = 32'd268468224;
      52623: inst = 32'd201347323;
      52624: inst = 32'd203423744;
      52625: inst = 32'd471859200;
      52626: inst = 32'd136314880;
      52627: inst = 32'd268468224;
      52628: inst = 32'd201347324;
      52629: inst = 32'd203423744;
      52630: inst = 32'd471859200;
      52631: inst = 32'd136314880;
      52632: inst = 32'd268468224;
      52633: inst = 32'd201347325;
      52634: inst = 32'd203423744;
      52635: inst = 32'd471859200;
      52636: inst = 32'd136314880;
      52637: inst = 32'd268468224;
      52638: inst = 32'd201347326;
      52639: inst = 32'd203423744;
      52640: inst = 32'd471859200;
      52641: inst = 32'd136314880;
      52642: inst = 32'd268468224;
      52643: inst = 32'd201347327;
      52644: inst = 32'd203423744;
      52645: inst = 32'd471859200;
      52646: inst = 32'd136314880;
      52647: inst = 32'd268468224;
      52648: inst = 32'd201347328;
      52649: inst = 32'd203423744;
      52650: inst = 32'd471859200;
      52651: inst = 32'd136314880;
      52652: inst = 32'd268468224;
      52653: inst = 32'd201347329;
      52654: inst = 32'd203423744;
      52655: inst = 32'd471859200;
      52656: inst = 32'd136314880;
      52657: inst = 32'd268468224;
      52658: inst = 32'd201347330;
      52659: inst = 32'd203423744;
      52660: inst = 32'd471859200;
      52661: inst = 32'd136314880;
      52662: inst = 32'd268468224;
      52663: inst = 32'd201347331;
      52664: inst = 32'd203423744;
      52665: inst = 32'd471859200;
      52666: inst = 32'd136314880;
      52667: inst = 32'd268468224;
      52668: inst = 32'd201347332;
      52669: inst = 32'd203423744;
      52670: inst = 32'd471859200;
      52671: inst = 32'd136314880;
      52672: inst = 32'd268468224;
      52673: inst = 32'd201347333;
      52674: inst = 32'd203423744;
      52675: inst = 32'd471859200;
      52676: inst = 32'd136314880;
      52677: inst = 32'd268468224;
      52678: inst = 32'd201347334;
      52679: inst = 32'd203423744;
      52680: inst = 32'd471859200;
      52681: inst = 32'd136314880;
      52682: inst = 32'd268468224;
      52683: inst = 32'd201347335;
      52684: inst = 32'd203423744;
      52685: inst = 32'd471859200;
      52686: inst = 32'd136314880;
      52687: inst = 32'd268468224;
      52688: inst = 32'd201347336;
      52689: inst = 32'd203423744;
      52690: inst = 32'd471859200;
      52691: inst = 32'd136314880;
      52692: inst = 32'd268468224;
      52693: inst = 32'd201347337;
      52694: inst = 32'd203423744;
      52695: inst = 32'd471859200;
      52696: inst = 32'd136314880;
      52697: inst = 32'd268468224;
      52698: inst = 32'd201347338;
      52699: inst = 32'd203423744;
      52700: inst = 32'd471859200;
      52701: inst = 32'd136314880;
      52702: inst = 32'd268468224;
      52703: inst = 32'd201347339;
      52704: inst = 32'd203423744;
      52705: inst = 32'd471859200;
      52706: inst = 32'd136314880;
      52707: inst = 32'd268468224;
      52708: inst = 32'd201347340;
      52709: inst = 32'd203423744;
      52710: inst = 32'd471859200;
      52711: inst = 32'd136314880;
      52712: inst = 32'd268468224;
      52713: inst = 32'd201347341;
      52714: inst = 32'd203423744;
      52715: inst = 32'd471859200;
      52716: inst = 32'd136314880;
      52717: inst = 32'd268468224;
      52718: inst = 32'd201347342;
      52719: inst = 32'd203423744;
      52720: inst = 32'd471859200;
      52721: inst = 32'd136314880;
      52722: inst = 32'd268468224;
      52723: inst = 32'd201347343;
      52724: inst = 32'd203423744;
      52725: inst = 32'd471859200;
      52726: inst = 32'd136314880;
      52727: inst = 32'd268468224;
      52728: inst = 32'd201347344;
      52729: inst = 32'd203423744;
      52730: inst = 32'd471859200;
      52731: inst = 32'd136314880;
      52732: inst = 32'd268468224;
      52733: inst = 32'd201347345;
      52734: inst = 32'd203423744;
      52735: inst = 32'd471859200;
      52736: inst = 32'd136314880;
      52737: inst = 32'd268468224;
      52738: inst = 32'd201347346;
      52739: inst = 32'd203423744;
      52740: inst = 32'd471859200;
      52741: inst = 32'd136314880;
      52742: inst = 32'd268468224;
      52743: inst = 32'd201347347;
      52744: inst = 32'd203423744;
      52745: inst = 32'd471859200;
      52746: inst = 32'd136314880;
      52747: inst = 32'd268468224;
      52748: inst = 32'd201347348;
      52749: inst = 32'd203423744;
      52750: inst = 32'd471859200;
      52751: inst = 32'd136314880;
      52752: inst = 32'd268468224;
      52753: inst = 32'd201347349;
      52754: inst = 32'd203423744;
      52755: inst = 32'd471859200;
      52756: inst = 32'd136314880;
      52757: inst = 32'd268468224;
      52758: inst = 32'd201347350;
      52759: inst = 32'd203423744;
      52760: inst = 32'd471859200;
      52761: inst = 32'd136314880;
      52762: inst = 32'd268468224;
      52763: inst = 32'd201347351;
      52764: inst = 32'd203423744;
      52765: inst = 32'd471859200;
      52766: inst = 32'd136314880;
      52767: inst = 32'd268468224;
      52768: inst = 32'd201347352;
      52769: inst = 32'd203423744;
      52770: inst = 32'd471859200;
      52771: inst = 32'd136314880;
      52772: inst = 32'd268468224;
      52773: inst = 32'd201347353;
      52774: inst = 32'd203423744;
      52775: inst = 32'd471859200;
      52776: inst = 32'd136314880;
      52777: inst = 32'd268468224;
      52778: inst = 32'd201347354;
      52779: inst = 32'd203423744;
      52780: inst = 32'd471859200;
      52781: inst = 32'd136314880;
      52782: inst = 32'd268468224;
      52783: inst = 32'd201347355;
      52784: inst = 32'd203423744;
      52785: inst = 32'd471859200;
      52786: inst = 32'd136314880;
      52787: inst = 32'd268468224;
      52788: inst = 32'd201347356;
      52789: inst = 32'd203423744;
      52790: inst = 32'd471859200;
      52791: inst = 32'd136314880;
      52792: inst = 32'd268468224;
      52793: inst = 32'd201347357;
      52794: inst = 32'd203423744;
      52795: inst = 32'd471859200;
      52796: inst = 32'd136314880;
      52797: inst = 32'd268468224;
      52798: inst = 32'd201347358;
      52799: inst = 32'd203423744;
      52800: inst = 32'd471859200;
      52801: inst = 32'd136314880;
      52802: inst = 32'd268468224;
      52803: inst = 32'd201347359;
      52804: inst = 32'd203423744;
      52805: inst = 32'd471859200;
      52806: inst = 32'd136314880;
      52807: inst = 32'd268468224;
      52808: inst = 32'd201347360;
      52809: inst = 32'd203423744;
      52810: inst = 32'd471859200;
      52811: inst = 32'd136314880;
      52812: inst = 32'd268468224;
      52813: inst = 32'd201347361;
      52814: inst = 32'd203423744;
      52815: inst = 32'd471859200;
      52816: inst = 32'd136314880;
      52817: inst = 32'd268468224;
      52818: inst = 32'd201347362;
      52819: inst = 32'd203423744;
      52820: inst = 32'd471859200;
      52821: inst = 32'd136314880;
      52822: inst = 32'd268468224;
      52823: inst = 32'd201347363;
      52824: inst = 32'd203423744;
      52825: inst = 32'd471859200;
      52826: inst = 32'd136314880;
      52827: inst = 32'd268468224;
      52828: inst = 32'd201347364;
      52829: inst = 32'd203423744;
      52830: inst = 32'd471859200;
      52831: inst = 32'd136314880;
      52832: inst = 32'd268468224;
      52833: inst = 32'd201347365;
      52834: inst = 32'd203423744;
      52835: inst = 32'd471859200;
      52836: inst = 32'd136314880;
      52837: inst = 32'd268468224;
      52838: inst = 32'd201347366;
      52839: inst = 32'd203423744;
      52840: inst = 32'd471859200;
      52841: inst = 32'd136314880;
      52842: inst = 32'd268468224;
      52843: inst = 32'd201347367;
      52844: inst = 32'd203423744;
      52845: inst = 32'd471859200;
      52846: inst = 32'd136314880;
      52847: inst = 32'd268468224;
      52848: inst = 32'd201347368;
      52849: inst = 32'd203423744;
      52850: inst = 32'd471859200;
      52851: inst = 32'd136314880;
      52852: inst = 32'd268468224;
      52853: inst = 32'd201347369;
      52854: inst = 32'd203423744;
      52855: inst = 32'd471859200;
      52856: inst = 32'd136314880;
      52857: inst = 32'd268468224;
      52858: inst = 32'd201347370;
      52859: inst = 32'd203423744;
      52860: inst = 32'd471859200;
      52861: inst = 32'd136314880;
      52862: inst = 32'd268468224;
      52863: inst = 32'd201347371;
      52864: inst = 32'd203423744;
      52865: inst = 32'd471859200;
      52866: inst = 32'd136314880;
      52867: inst = 32'd268468224;
      52868: inst = 32'd201347372;
      52869: inst = 32'd203423744;
      52870: inst = 32'd471859200;
      52871: inst = 32'd136314880;
      52872: inst = 32'd268468224;
      52873: inst = 32'd201347373;
      52874: inst = 32'd203423744;
      52875: inst = 32'd471859200;
      52876: inst = 32'd136314880;
      52877: inst = 32'd268468224;
      52878: inst = 32'd201347374;
      52879: inst = 32'd203423744;
      52880: inst = 32'd471859200;
      52881: inst = 32'd136314880;
      52882: inst = 32'd268468224;
      52883: inst = 32'd201347375;
      52884: inst = 32'd203423744;
      52885: inst = 32'd471859200;
      52886: inst = 32'd136314880;
      52887: inst = 32'd268468224;
      52888: inst = 32'd201347376;
      52889: inst = 32'd203423744;
      52890: inst = 32'd471859200;
      52891: inst = 32'd136314880;
      52892: inst = 32'd268468224;
      52893: inst = 32'd201347377;
      52894: inst = 32'd203423744;
      52895: inst = 32'd471859200;
      52896: inst = 32'd136314880;
      52897: inst = 32'd268468224;
      52898: inst = 32'd201347378;
      52899: inst = 32'd203423744;
      52900: inst = 32'd471859200;
      52901: inst = 32'd136314880;
      52902: inst = 32'd268468224;
      52903: inst = 32'd201347379;
      52904: inst = 32'd203423744;
      52905: inst = 32'd471859200;
      52906: inst = 32'd136314880;
      52907: inst = 32'd268468224;
      52908: inst = 32'd201347380;
      52909: inst = 32'd203423744;
      52910: inst = 32'd471859200;
      52911: inst = 32'd136314880;
      52912: inst = 32'd268468224;
      52913: inst = 32'd201347381;
      52914: inst = 32'd203423744;
      52915: inst = 32'd471859200;
      52916: inst = 32'd136314880;
      52917: inst = 32'd268468224;
      52918: inst = 32'd201347382;
      52919: inst = 32'd203423744;
      52920: inst = 32'd471859200;
      52921: inst = 32'd136314880;
      52922: inst = 32'd268468224;
      52923: inst = 32'd201347383;
      52924: inst = 32'd203423744;
      52925: inst = 32'd471859200;
      52926: inst = 32'd136314880;
      52927: inst = 32'd268468224;
      52928: inst = 32'd201347384;
      52929: inst = 32'd203423744;
      52930: inst = 32'd471859200;
      52931: inst = 32'd136314880;
      52932: inst = 32'd268468224;
      52933: inst = 32'd201347385;
      52934: inst = 32'd203423744;
      52935: inst = 32'd471859200;
      52936: inst = 32'd136314880;
      52937: inst = 32'd268468224;
      52938: inst = 32'd201347386;
      52939: inst = 32'd203423744;
      52940: inst = 32'd471859200;
      52941: inst = 32'd136314880;
      52942: inst = 32'd268468224;
      52943: inst = 32'd201347387;
      52944: inst = 32'd203423744;
      52945: inst = 32'd471859200;
      52946: inst = 32'd136314880;
      52947: inst = 32'd268468224;
      52948: inst = 32'd201347388;
      52949: inst = 32'd203423744;
      52950: inst = 32'd471859200;
      52951: inst = 32'd136314880;
      52952: inst = 32'd268468224;
      52953: inst = 32'd201347389;
      52954: inst = 32'd203423744;
      52955: inst = 32'd471859200;
      52956: inst = 32'd136314880;
      52957: inst = 32'd268468224;
      52958: inst = 32'd201347390;
      52959: inst = 32'd203423744;
      52960: inst = 32'd471859200;
      52961: inst = 32'd136314880;
      52962: inst = 32'd268468224;
      52963: inst = 32'd201347391;
      52964: inst = 32'd203423744;
      52965: inst = 32'd471859200;
      52966: inst = 32'd136314880;
      52967: inst = 32'd268468224;
      52968: inst = 32'd201347392;
      52969: inst = 32'd203423744;
      52970: inst = 32'd471859200;
      52971: inst = 32'd136314880;
      52972: inst = 32'd268468224;
      52973: inst = 32'd201347393;
      52974: inst = 32'd203423744;
      52975: inst = 32'd471859200;
      52976: inst = 32'd136314880;
      52977: inst = 32'd268468224;
      52978: inst = 32'd201347394;
      52979: inst = 32'd203423744;
      52980: inst = 32'd471859200;
      52981: inst = 32'd136314880;
      52982: inst = 32'd268468224;
      52983: inst = 32'd201347395;
      52984: inst = 32'd203423744;
      52985: inst = 32'd471859200;
      52986: inst = 32'd136314880;
      52987: inst = 32'd268468224;
      52988: inst = 32'd201347396;
      52989: inst = 32'd203423744;
      52990: inst = 32'd471859200;
      52991: inst = 32'd136314880;
      52992: inst = 32'd268468224;
      52993: inst = 32'd201347397;
      52994: inst = 32'd203423744;
      52995: inst = 32'd471859200;
      52996: inst = 32'd136314880;
      52997: inst = 32'd268468224;
      52998: inst = 32'd201347398;
      52999: inst = 32'd203423744;
      53000: inst = 32'd471859200;
      53001: inst = 32'd136314880;
      53002: inst = 32'd268468224;
      53003: inst = 32'd201347399;
      53004: inst = 32'd203423744;
      53005: inst = 32'd471859200;
      53006: inst = 32'd136314880;
      53007: inst = 32'd268468224;
      53008: inst = 32'd201347400;
      53009: inst = 32'd203423744;
      53010: inst = 32'd471859200;
      53011: inst = 32'd136314880;
      53012: inst = 32'd268468224;
      53013: inst = 32'd201347401;
      53014: inst = 32'd203423744;
      53015: inst = 32'd471859200;
      53016: inst = 32'd136314880;
      53017: inst = 32'd268468224;
      53018: inst = 32'd201347402;
      53019: inst = 32'd203423744;
      53020: inst = 32'd471859200;
      53021: inst = 32'd136314880;
      53022: inst = 32'd268468224;
      53023: inst = 32'd201347403;
      53024: inst = 32'd203423744;
      53025: inst = 32'd471859200;
      53026: inst = 32'd136314880;
      53027: inst = 32'd268468224;
      53028: inst = 32'd201347404;
      53029: inst = 32'd203423744;
      53030: inst = 32'd471859200;
      53031: inst = 32'd136314880;
      53032: inst = 32'd268468224;
      53033: inst = 32'd201347405;
      53034: inst = 32'd203423744;
      53035: inst = 32'd471859200;
      53036: inst = 32'd136314880;
      53037: inst = 32'd268468224;
      53038: inst = 32'd201347406;
      53039: inst = 32'd203423744;
      53040: inst = 32'd471859200;
      53041: inst = 32'd136314880;
      53042: inst = 32'd268468224;
      53043: inst = 32'd201347407;
      53044: inst = 32'd203423744;
      53045: inst = 32'd471859200;
      53046: inst = 32'd136314880;
      53047: inst = 32'd268468224;
      53048: inst = 32'd201347408;
      53049: inst = 32'd203423744;
      53050: inst = 32'd471859200;
      53051: inst = 32'd136314880;
      53052: inst = 32'd268468224;
      53053: inst = 32'd201347409;
      53054: inst = 32'd203423744;
      53055: inst = 32'd471859200;
      53056: inst = 32'd136314880;
      53057: inst = 32'd268468224;
      53058: inst = 32'd201347410;
      53059: inst = 32'd203423744;
      53060: inst = 32'd471859200;
      53061: inst = 32'd136314880;
      53062: inst = 32'd268468224;
      53063: inst = 32'd201347411;
      53064: inst = 32'd203423744;
      53065: inst = 32'd471859200;
      53066: inst = 32'd136314880;
      53067: inst = 32'd268468224;
      53068: inst = 32'd201347412;
      53069: inst = 32'd203423744;
      53070: inst = 32'd471859200;
      53071: inst = 32'd136314880;
      53072: inst = 32'd268468224;
      53073: inst = 32'd201347413;
      53074: inst = 32'd203423744;
      53075: inst = 32'd471859200;
      53076: inst = 32'd136314880;
      53077: inst = 32'd268468224;
      53078: inst = 32'd201347414;
      53079: inst = 32'd203423744;
      53080: inst = 32'd471859200;
      53081: inst = 32'd136314880;
      53082: inst = 32'd268468224;
      53083: inst = 32'd201347415;
      53084: inst = 32'd203423744;
      53085: inst = 32'd471859200;
      53086: inst = 32'd136314880;
      53087: inst = 32'd268468224;
      53088: inst = 32'd201347416;
      53089: inst = 32'd203423744;
      53090: inst = 32'd471859200;
      53091: inst = 32'd136314880;
      53092: inst = 32'd268468224;
      53093: inst = 32'd201347417;
      53094: inst = 32'd203423744;
      53095: inst = 32'd471859200;
      53096: inst = 32'd136314880;
      53097: inst = 32'd268468224;
      53098: inst = 32'd201347418;
      53099: inst = 32'd203423744;
      53100: inst = 32'd471859200;
      53101: inst = 32'd136314880;
      53102: inst = 32'd268468224;
      53103: inst = 32'd201347419;
      53104: inst = 32'd203423744;
      53105: inst = 32'd471859200;
      53106: inst = 32'd136314880;
      53107: inst = 32'd268468224;
      53108: inst = 32'd201347420;
      53109: inst = 32'd203423744;
      53110: inst = 32'd471859200;
      53111: inst = 32'd136314880;
      53112: inst = 32'd268468224;
      53113: inst = 32'd201347421;
      53114: inst = 32'd203423744;
      53115: inst = 32'd471859200;
      53116: inst = 32'd136314880;
      53117: inst = 32'd268468224;
      53118: inst = 32'd201347422;
      53119: inst = 32'd203423744;
      53120: inst = 32'd471859200;
      53121: inst = 32'd136314880;
      53122: inst = 32'd268468224;
      53123: inst = 32'd201347423;
      53124: inst = 32'd203423744;
      53125: inst = 32'd471859200;
      53126: inst = 32'd136314880;
      53127: inst = 32'd268468224;
      53128: inst = 32'd201347424;
      53129: inst = 32'd203423744;
      53130: inst = 32'd471859200;
      53131: inst = 32'd136314880;
      53132: inst = 32'd268468224;
      53133: inst = 32'd201347425;
      53134: inst = 32'd203423744;
      53135: inst = 32'd471859200;
      53136: inst = 32'd136314880;
      53137: inst = 32'd268468224;
      53138: inst = 32'd201347426;
      53139: inst = 32'd203423744;
      53140: inst = 32'd471859200;
      53141: inst = 32'd136314880;
      53142: inst = 32'd268468224;
      53143: inst = 32'd201347427;
      53144: inst = 32'd203423744;
      53145: inst = 32'd471859200;
      53146: inst = 32'd136314880;
      53147: inst = 32'd268468224;
      53148: inst = 32'd201347428;
      53149: inst = 32'd203423744;
      53150: inst = 32'd471859200;
      53151: inst = 32'd136314880;
      53152: inst = 32'd268468224;
      53153: inst = 32'd201347429;
      53154: inst = 32'd203423744;
      53155: inst = 32'd471859200;
      53156: inst = 32'd136314880;
      53157: inst = 32'd268468224;
      53158: inst = 32'd201347430;
      53159: inst = 32'd203423744;
      53160: inst = 32'd471859200;
      53161: inst = 32'd136314880;
      53162: inst = 32'd268468224;
      53163: inst = 32'd201347431;
      53164: inst = 32'd203423744;
      53165: inst = 32'd471859200;
      53166: inst = 32'd136314880;
      53167: inst = 32'd268468224;
      53168: inst = 32'd201347432;
      53169: inst = 32'd203423744;
      53170: inst = 32'd471859200;
      53171: inst = 32'd136314880;
      53172: inst = 32'd268468224;
      53173: inst = 32'd201347433;
      53174: inst = 32'd203423744;
      53175: inst = 32'd471859200;
      53176: inst = 32'd136314880;
      53177: inst = 32'd268468224;
      53178: inst = 32'd201347434;
      53179: inst = 32'd203423744;
      53180: inst = 32'd471859200;
      53181: inst = 32'd136314880;
      53182: inst = 32'd268468224;
      53183: inst = 32'd201347435;
      53184: inst = 32'd203423744;
      53185: inst = 32'd471859200;
      53186: inst = 32'd136314880;
      53187: inst = 32'd268468224;
      53188: inst = 32'd201347436;
      53189: inst = 32'd203423744;
      53190: inst = 32'd471859200;
      53191: inst = 32'd136314880;
      53192: inst = 32'd268468224;
      53193: inst = 32'd201347437;
      53194: inst = 32'd203423744;
      53195: inst = 32'd471859200;
      53196: inst = 32'd136314880;
      53197: inst = 32'd268468224;
      53198: inst = 32'd201347438;
      53199: inst = 32'd203423744;
      53200: inst = 32'd471859200;
      53201: inst = 32'd136314880;
      53202: inst = 32'd268468224;
      53203: inst = 32'd201347439;
      53204: inst = 32'd203423744;
      53205: inst = 32'd471859200;
      53206: inst = 32'd136314880;
      53207: inst = 32'd268468224;
      53208: inst = 32'd201347440;
      53209: inst = 32'd203423744;
      53210: inst = 32'd471859200;
      53211: inst = 32'd136314880;
      53212: inst = 32'd268468224;
      53213: inst = 32'd201347441;
      53214: inst = 32'd203423744;
      53215: inst = 32'd471859200;
      53216: inst = 32'd136314880;
      53217: inst = 32'd268468224;
      53218: inst = 32'd201347442;
      53219: inst = 32'd203423744;
      53220: inst = 32'd471859200;
      53221: inst = 32'd136314880;
      53222: inst = 32'd268468224;
      53223: inst = 32'd201347443;
      53224: inst = 32'd203423744;
      53225: inst = 32'd471859200;
      53226: inst = 32'd136314880;
      53227: inst = 32'd268468224;
      53228: inst = 32'd201347444;
      53229: inst = 32'd203423744;
      53230: inst = 32'd471859200;
      53231: inst = 32'd136314880;
      53232: inst = 32'd268468224;
      53233: inst = 32'd201347445;
      53234: inst = 32'd203423744;
      53235: inst = 32'd471859200;
      53236: inst = 32'd136314880;
      53237: inst = 32'd268468224;
      53238: inst = 32'd201347446;
      53239: inst = 32'd203423744;
      53240: inst = 32'd471859200;
      53241: inst = 32'd136314880;
      53242: inst = 32'd268468224;
      53243: inst = 32'd201347447;
      53244: inst = 32'd203423744;
      53245: inst = 32'd471859200;
      53246: inst = 32'd136314880;
      53247: inst = 32'd268468224;
      53248: inst = 32'd201347448;
      53249: inst = 32'd203423744;
      53250: inst = 32'd471859200;
      53251: inst = 32'd136314880;
      53252: inst = 32'd268468224;
      53253: inst = 32'd201347449;
      53254: inst = 32'd203423744;
      53255: inst = 32'd471859200;
      53256: inst = 32'd136314880;
      53257: inst = 32'd268468224;
      53258: inst = 32'd201347450;
      53259: inst = 32'd203423744;
      53260: inst = 32'd471859200;
      53261: inst = 32'd136314880;
      53262: inst = 32'd268468224;
      53263: inst = 32'd201347451;
      53264: inst = 32'd203423744;
      53265: inst = 32'd471859200;
      53266: inst = 32'd136314880;
      53267: inst = 32'd268468224;
      53268: inst = 32'd201347452;
      53269: inst = 32'd203423744;
      53270: inst = 32'd471859200;
      53271: inst = 32'd136314880;
      53272: inst = 32'd268468224;
      53273: inst = 32'd201347453;
      53274: inst = 32'd203423744;
      53275: inst = 32'd471859200;
      53276: inst = 32'd136314880;
      53277: inst = 32'd268468224;
      53278: inst = 32'd201347454;
      53279: inst = 32'd203423744;
      53280: inst = 32'd471859200;
      53281: inst = 32'd136314880;
      53282: inst = 32'd268468224;
      53283: inst = 32'd201347455;
      53284: inst = 32'd203423744;
      53285: inst = 32'd471859200;
      53286: inst = 32'd136314880;
      53287: inst = 32'd268468224;
      53288: inst = 32'd201347456;
      53289: inst = 32'd203423744;
      53290: inst = 32'd471859200;
      53291: inst = 32'd136314880;
      53292: inst = 32'd268468224;
      53293: inst = 32'd201347457;
      53294: inst = 32'd203423744;
      53295: inst = 32'd471859200;
      53296: inst = 32'd136314880;
      53297: inst = 32'd268468224;
      53298: inst = 32'd201347458;
      53299: inst = 32'd203423744;
      53300: inst = 32'd471859200;
      53301: inst = 32'd136314880;
      53302: inst = 32'd268468224;
      53303: inst = 32'd201347459;
      53304: inst = 32'd203423744;
      53305: inst = 32'd471859200;
      53306: inst = 32'd136314880;
      53307: inst = 32'd268468224;
      53308: inst = 32'd201347460;
      53309: inst = 32'd203423744;
      53310: inst = 32'd471859200;
      53311: inst = 32'd136314880;
      53312: inst = 32'd268468224;
      53313: inst = 32'd201347461;
      53314: inst = 32'd203423744;
      53315: inst = 32'd471859200;
      53316: inst = 32'd136314880;
      53317: inst = 32'd268468224;
      53318: inst = 32'd201347462;
      53319: inst = 32'd203423744;
      53320: inst = 32'd471859200;
      53321: inst = 32'd136314880;
      53322: inst = 32'd268468224;
      53323: inst = 32'd201347463;
      53324: inst = 32'd203423744;
      53325: inst = 32'd471859200;
      53326: inst = 32'd136314880;
      53327: inst = 32'd268468224;
      53328: inst = 32'd201347464;
      53329: inst = 32'd203423744;
      53330: inst = 32'd471859200;
      53331: inst = 32'd136314880;
      53332: inst = 32'd268468224;
      53333: inst = 32'd201347465;
      53334: inst = 32'd203423744;
      53335: inst = 32'd471859200;
      53336: inst = 32'd136314880;
      53337: inst = 32'd268468224;
      53338: inst = 32'd201347466;
      53339: inst = 32'd203423744;
      53340: inst = 32'd471859200;
      53341: inst = 32'd136314880;
      53342: inst = 32'd268468224;
      53343: inst = 32'd201347467;
      53344: inst = 32'd203423744;
      53345: inst = 32'd471859200;
      53346: inst = 32'd136314880;
      53347: inst = 32'd268468224;
      53348: inst = 32'd201347468;
      53349: inst = 32'd203423744;
      53350: inst = 32'd471859200;
      53351: inst = 32'd136314880;
      53352: inst = 32'd268468224;
      53353: inst = 32'd201347469;
      53354: inst = 32'd203423744;
      53355: inst = 32'd471859200;
      53356: inst = 32'd136314880;
      53357: inst = 32'd268468224;
      53358: inst = 32'd201347470;
      53359: inst = 32'd203423744;
      53360: inst = 32'd471859200;
      53361: inst = 32'd136314880;
      53362: inst = 32'd268468224;
      53363: inst = 32'd201347471;
      53364: inst = 32'd203423744;
      53365: inst = 32'd471859200;
      53366: inst = 32'd136314880;
      53367: inst = 32'd268468224;
      53368: inst = 32'd201347472;
      53369: inst = 32'd203423744;
      53370: inst = 32'd471859200;
      53371: inst = 32'd136314880;
      53372: inst = 32'd268468224;
      53373: inst = 32'd201347473;
      53374: inst = 32'd203423744;
      53375: inst = 32'd471859200;
      53376: inst = 32'd136314880;
      53377: inst = 32'd268468224;
      53378: inst = 32'd201347474;
      53379: inst = 32'd203423744;
      53380: inst = 32'd471859200;
      53381: inst = 32'd136314880;
      53382: inst = 32'd268468224;
      53383: inst = 32'd201347475;
      53384: inst = 32'd203423744;
      53385: inst = 32'd471859200;
      53386: inst = 32'd136314880;
      53387: inst = 32'd268468224;
      53388: inst = 32'd201347476;
      53389: inst = 32'd203423744;
      53390: inst = 32'd471859200;
      53391: inst = 32'd136314880;
      53392: inst = 32'd268468224;
      53393: inst = 32'd201347477;
      53394: inst = 32'd203423744;
      53395: inst = 32'd471859200;
      53396: inst = 32'd136314880;
      53397: inst = 32'd268468224;
      53398: inst = 32'd201347478;
      53399: inst = 32'd203423744;
      53400: inst = 32'd471859200;
      53401: inst = 32'd136314880;
      53402: inst = 32'd268468224;
      53403: inst = 32'd201347479;
      53404: inst = 32'd203423744;
      53405: inst = 32'd471859200;
      53406: inst = 32'd136314880;
      53407: inst = 32'd268468224;
      53408: inst = 32'd201347480;
      53409: inst = 32'd203423744;
      53410: inst = 32'd471859200;
      53411: inst = 32'd136314880;
      53412: inst = 32'd268468224;
      53413: inst = 32'd201347481;
      53414: inst = 32'd203423744;
      53415: inst = 32'd471859200;
      53416: inst = 32'd136314880;
      53417: inst = 32'd268468224;
      53418: inst = 32'd201347482;
      53419: inst = 32'd203423744;
      53420: inst = 32'd471859200;
      53421: inst = 32'd136314880;
      53422: inst = 32'd268468224;
      53423: inst = 32'd201347483;
      53424: inst = 32'd203423744;
      53425: inst = 32'd471859200;
      53426: inst = 32'd136314880;
      53427: inst = 32'd268468224;
      53428: inst = 32'd201347484;
      53429: inst = 32'd203423744;
      53430: inst = 32'd471859200;
      53431: inst = 32'd136314880;
      53432: inst = 32'd268468224;
      53433: inst = 32'd201347485;
      53434: inst = 32'd203423744;
      53435: inst = 32'd471859200;
      53436: inst = 32'd136314880;
      53437: inst = 32'd268468224;
      53438: inst = 32'd201347486;
      53439: inst = 32'd203423744;
      53440: inst = 32'd471859200;
      53441: inst = 32'd136314880;
      53442: inst = 32'd268468224;
      53443: inst = 32'd201347487;
      53444: inst = 32'd203423744;
      53445: inst = 32'd471859200;
      53446: inst = 32'd136314880;
      53447: inst = 32'd268468224;
      53448: inst = 32'd201347488;
      53449: inst = 32'd203423744;
      53450: inst = 32'd471859200;
      53451: inst = 32'd136314880;
      53452: inst = 32'd268468224;
      53453: inst = 32'd201347489;
      53454: inst = 32'd203423744;
      53455: inst = 32'd471859200;
      53456: inst = 32'd136314880;
      53457: inst = 32'd268468224;
      53458: inst = 32'd201347490;
      53459: inst = 32'd203423744;
      53460: inst = 32'd471859200;
      53461: inst = 32'd136314880;
      53462: inst = 32'd268468224;
      53463: inst = 32'd201347491;
      53464: inst = 32'd203423744;
      53465: inst = 32'd471859200;
      53466: inst = 32'd136314880;
      53467: inst = 32'd268468224;
      53468: inst = 32'd201347492;
      53469: inst = 32'd203423744;
      53470: inst = 32'd471859200;
      53471: inst = 32'd136314880;
      53472: inst = 32'd268468224;
      53473: inst = 32'd201347493;
      53474: inst = 32'd203423744;
      53475: inst = 32'd471859200;
      53476: inst = 32'd136314880;
      53477: inst = 32'd268468224;
      53478: inst = 32'd201347494;
      53479: inst = 32'd203423744;
      53480: inst = 32'd471859200;
      53481: inst = 32'd136314880;
      53482: inst = 32'd268468224;
      53483: inst = 32'd201347495;
      53484: inst = 32'd203423744;
      53485: inst = 32'd471859200;
      53486: inst = 32'd136314880;
      53487: inst = 32'd268468224;
      53488: inst = 32'd201347496;
      53489: inst = 32'd203423744;
      53490: inst = 32'd471859200;
      53491: inst = 32'd136314880;
      53492: inst = 32'd268468224;
      53493: inst = 32'd201347497;
      53494: inst = 32'd203423744;
      53495: inst = 32'd471859200;
      53496: inst = 32'd136314880;
      53497: inst = 32'd268468224;
      53498: inst = 32'd201347498;
      53499: inst = 32'd203423744;
      53500: inst = 32'd471859200;
      53501: inst = 32'd136314880;
      53502: inst = 32'd268468224;
      53503: inst = 32'd201347499;
      53504: inst = 32'd203423744;
      53505: inst = 32'd471859200;
      53506: inst = 32'd136314880;
      53507: inst = 32'd268468224;
      53508: inst = 32'd201347500;
      53509: inst = 32'd203423744;
      53510: inst = 32'd471859200;
      53511: inst = 32'd136314880;
      53512: inst = 32'd268468224;
      53513: inst = 32'd201347501;
      53514: inst = 32'd203423744;
      53515: inst = 32'd471859200;
      53516: inst = 32'd136314880;
      53517: inst = 32'd268468224;
      53518: inst = 32'd201347502;
      53519: inst = 32'd203423744;
      53520: inst = 32'd471859200;
      53521: inst = 32'd136314880;
      53522: inst = 32'd268468224;
      53523: inst = 32'd201347503;
      53524: inst = 32'd203423744;
      53525: inst = 32'd471859200;
      53526: inst = 32'd136314880;
      53527: inst = 32'd268468224;
      53528: inst = 32'd201347504;
      53529: inst = 32'd203423744;
      53530: inst = 32'd471859200;
      53531: inst = 32'd136314880;
      53532: inst = 32'd268468224;
      53533: inst = 32'd201347505;
      53534: inst = 32'd203423744;
      53535: inst = 32'd471859200;
      53536: inst = 32'd136314880;
      53537: inst = 32'd268468224;
      53538: inst = 32'd201347506;
      53539: inst = 32'd203423744;
      53540: inst = 32'd471859200;
      53541: inst = 32'd136314880;
      53542: inst = 32'd268468224;
      53543: inst = 32'd201347507;
      53544: inst = 32'd203423744;
      53545: inst = 32'd471859200;
      53546: inst = 32'd136314880;
      53547: inst = 32'd268468224;
      53548: inst = 32'd201347508;
      53549: inst = 32'd203423744;
      53550: inst = 32'd471859200;
      53551: inst = 32'd136314880;
      53552: inst = 32'd268468224;
      53553: inst = 32'd201347509;
      53554: inst = 32'd203423744;
      53555: inst = 32'd471859200;
      53556: inst = 32'd136314880;
      53557: inst = 32'd268468224;
      53558: inst = 32'd201347510;
      53559: inst = 32'd203423744;
      53560: inst = 32'd471859200;
      53561: inst = 32'd136314880;
      53562: inst = 32'd268468224;
      53563: inst = 32'd201347511;
      53564: inst = 32'd203423744;
      53565: inst = 32'd471859200;
      53566: inst = 32'd136314880;
      53567: inst = 32'd268468224;
      53568: inst = 32'd201347512;
      53569: inst = 32'd203423744;
      53570: inst = 32'd471859200;
      53571: inst = 32'd136314880;
      53572: inst = 32'd268468224;
      53573: inst = 32'd201347513;
      53574: inst = 32'd203423744;
      53575: inst = 32'd471859200;
      53576: inst = 32'd136314880;
      53577: inst = 32'd268468224;
      53578: inst = 32'd201347514;
      53579: inst = 32'd203423744;
      53580: inst = 32'd471859200;
      53581: inst = 32'd136314880;
      53582: inst = 32'd268468224;
      53583: inst = 32'd201347515;
      53584: inst = 32'd203423744;
      53585: inst = 32'd471859200;
      53586: inst = 32'd136314880;
      53587: inst = 32'd268468224;
      53588: inst = 32'd201347516;
      53589: inst = 32'd203423744;
      53590: inst = 32'd471859200;
      53591: inst = 32'd136314880;
      53592: inst = 32'd268468224;
      53593: inst = 32'd201347517;
      53594: inst = 32'd203423744;
      53595: inst = 32'd471859200;
      53596: inst = 32'd136314880;
      53597: inst = 32'd268468224;
      53598: inst = 32'd201347518;
      53599: inst = 32'd203423744;
      53600: inst = 32'd471859200;
      53601: inst = 32'd136314880;
      53602: inst = 32'd268468224;
      53603: inst = 32'd201347519;
      53604: inst = 32'd203423744;
      53605: inst = 32'd471859200;
      53606: inst = 32'd136314880;
      53607: inst = 32'd268468224;
      53608: inst = 32'd201347520;
      53609: inst = 32'd203423744;
      53610: inst = 32'd471859200;
      53611: inst = 32'd136314880;
      53612: inst = 32'd268468224;
      53613: inst = 32'd201347521;
      53614: inst = 32'd203423744;
      53615: inst = 32'd471859200;
      53616: inst = 32'd136314880;
      53617: inst = 32'd268468224;
      53618: inst = 32'd201347522;
      53619: inst = 32'd203423744;
      53620: inst = 32'd471859200;
      53621: inst = 32'd136314880;
      53622: inst = 32'd268468224;
      53623: inst = 32'd201347523;
      53624: inst = 32'd203423744;
      53625: inst = 32'd471859200;
      53626: inst = 32'd136314880;
      53627: inst = 32'd268468224;
      53628: inst = 32'd201347524;
      53629: inst = 32'd203423744;
      53630: inst = 32'd471859200;
      53631: inst = 32'd136314880;
      53632: inst = 32'd268468224;
      53633: inst = 32'd201347525;
      53634: inst = 32'd203423744;
      53635: inst = 32'd471859200;
      53636: inst = 32'd136314880;
      53637: inst = 32'd268468224;
      53638: inst = 32'd201347526;
      53639: inst = 32'd203423744;
      53640: inst = 32'd471859200;
      53641: inst = 32'd136314880;
      53642: inst = 32'd268468224;
      53643: inst = 32'd201347527;
      53644: inst = 32'd203423744;
      53645: inst = 32'd471859200;
      53646: inst = 32'd136314880;
      53647: inst = 32'd268468224;
      53648: inst = 32'd201347528;
      53649: inst = 32'd203423744;
      53650: inst = 32'd471859200;
      53651: inst = 32'd136314880;
      53652: inst = 32'd268468224;
      53653: inst = 32'd201347529;
      53654: inst = 32'd203423744;
      53655: inst = 32'd471859200;
      53656: inst = 32'd136314880;
      53657: inst = 32'd268468224;
      53658: inst = 32'd201347530;
      53659: inst = 32'd203423744;
      53660: inst = 32'd471859200;
      53661: inst = 32'd136314880;
      53662: inst = 32'd268468224;
      53663: inst = 32'd201347531;
      53664: inst = 32'd203423744;
      53665: inst = 32'd471859200;
      53666: inst = 32'd136314880;
      53667: inst = 32'd268468224;
      53668: inst = 32'd201347532;
      53669: inst = 32'd203423744;
      53670: inst = 32'd471859200;
      53671: inst = 32'd136314880;
      53672: inst = 32'd268468224;
      53673: inst = 32'd201347533;
      53674: inst = 32'd203423744;
      53675: inst = 32'd471859200;
      53676: inst = 32'd136314880;
      53677: inst = 32'd268468224;
      53678: inst = 32'd201347534;
      53679: inst = 32'd203423744;
      53680: inst = 32'd471859200;
      53681: inst = 32'd136314880;
      53682: inst = 32'd268468224;
      53683: inst = 32'd201347535;
      53684: inst = 32'd203423744;
      53685: inst = 32'd471859200;
      53686: inst = 32'd136314880;
      53687: inst = 32'd268468224;
      53688: inst = 32'd201347536;
      53689: inst = 32'd203423744;
      53690: inst = 32'd471859200;
      53691: inst = 32'd136314880;
      53692: inst = 32'd268468224;
      53693: inst = 32'd201347537;
      53694: inst = 32'd203423744;
      53695: inst = 32'd471859200;
      53696: inst = 32'd136314880;
      53697: inst = 32'd268468224;
      53698: inst = 32'd201347538;
      53699: inst = 32'd203423744;
      53700: inst = 32'd471859200;
      53701: inst = 32'd136314880;
      53702: inst = 32'd268468224;
      53703: inst = 32'd201347539;
      53704: inst = 32'd203423744;
      53705: inst = 32'd471859200;
      53706: inst = 32'd136314880;
      53707: inst = 32'd268468224;
      53708: inst = 32'd201347540;
      53709: inst = 32'd203423744;
      53710: inst = 32'd471859200;
      53711: inst = 32'd136314880;
      53712: inst = 32'd268468224;
      53713: inst = 32'd201347541;
      53714: inst = 32'd203423744;
      53715: inst = 32'd471859200;
      53716: inst = 32'd136314880;
      53717: inst = 32'd268468224;
      53718: inst = 32'd201347542;
      53719: inst = 32'd203423744;
      53720: inst = 32'd471859200;
      53721: inst = 32'd136314880;
      53722: inst = 32'd268468224;
      53723: inst = 32'd201347543;
      53724: inst = 32'd203423744;
      53725: inst = 32'd471859200;
      53726: inst = 32'd136314880;
      53727: inst = 32'd268468224;
      53728: inst = 32'd201347544;
      53729: inst = 32'd203423744;
      53730: inst = 32'd471859200;
      53731: inst = 32'd136314880;
      53732: inst = 32'd268468224;
      53733: inst = 32'd201347545;
      53734: inst = 32'd203423744;
      53735: inst = 32'd471859200;
      53736: inst = 32'd136314880;
      53737: inst = 32'd268468224;
      53738: inst = 32'd201347546;
      53739: inst = 32'd203423744;
      53740: inst = 32'd471859200;
      53741: inst = 32'd136314880;
      53742: inst = 32'd268468224;
      53743: inst = 32'd201347547;
      53744: inst = 32'd203423744;
      53745: inst = 32'd471859200;
      53746: inst = 32'd136314880;
      53747: inst = 32'd268468224;
      53748: inst = 32'd201347548;
      53749: inst = 32'd203423744;
      53750: inst = 32'd471859200;
      53751: inst = 32'd136314880;
      53752: inst = 32'd268468224;
      53753: inst = 32'd201347549;
      53754: inst = 32'd203423744;
      53755: inst = 32'd471859200;
      53756: inst = 32'd136314880;
      53757: inst = 32'd268468224;
      53758: inst = 32'd201347550;
      53759: inst = 32'd203423744;
      53760: inst = 32'd471859200;
      53761: inst = 32'd136314880;
      53762: inst = 32'd268468224;
      53763: inst = 32'd201347551;
      53764: inst = 32'd203423744;
      53765: inst = 32'd471859200;
      53766: inst = 32'd136314880;
      53767: inst = 32'd268468224;
      53768: inst = 32'd201347552;
      53769: inst = 32'd203423744;
      53770: inst = 32'd471859200;
      53771: inst = 32'd136314880;
      53772: inst = 32'd268468224;
      53773: inst = 32'd201347553;
      53774: inst = 32'd203423744;
      53775: inst = 32'd471859200;
      53776: inst = 32'd136314880;
      53777: inst = 32'd268468224;
      53778: inst = 32'd201347554;
      53779: inst = 32'd203423744;
      53780: inst = 32'd471859200;
      53781: inst = 32'd136314880;
      53782: inst = 32'd268468224;
      53783: inst = 32'd201347555;
      53784: inst = 32'd203423744;
      53785: inst = 32'd471859200;
      53786: inst = 32'd136314880;
      53787: inst = 32'd268468224;
      53788: inst = 32'd201347556;
      53789: inst = 32'd203423744;
      53790: inst = 32'd471859200;
      53791: inst = 32'd136314880;
      53792: inst = 32'd268468224;
      53793: inst = 32'd201347557;
      53794: inst = 32'd203423744;
      53795: inst = 32'd471859200;
      53796: inst = 32'd136314880;
      53797: inst = 32'd268468224;
      53798: inst = 32'd201347558;
      53799: inst = 32'd203423744;
      53800: inst = 32'd471859200;
      53801: inst = 32'd136314880;
      53802: inst = 32'd268468224;
      53803: inst = 32'd201347559;
      53804: inst = 32'd203423744;
      53805: inst = 32'd471859200;
      53806: inst = 32'd136314880;
      53807: inst = 32'd268468224;
      53808: inst = 32'd201347560;
      53809: inst = 32'd203423744;
      53810: inst = 32'd471859200;
      53811: inst = 32'd136314880;
      53812: inst = 32'd268468224;
      53813: inst = 32'd201347561;
      53814: inst = 32'd203423744;
      53815: inst = 32'd471859200;
      53816: inst = 32'd136314880;
      53817: inst = 32'd268468224;
      53818: inst = 32'd201347562;
      53819: inst = 32'd203423744;
      53820: inst = 32'd471859200;
      53821: inst = 32'd136314880;
      53822: inst = 32'd268468224;
      53823: inst = 32'd201347563;
      53824: inst = 32'd203423744;
      53825: inst = 32'd471859200;
      53826: inst = 32'd136314880;
      53827: inst = 32'd268468224;
      53828: inst = 32'd201347564;
      53829: inst = 32'd203423744;
      53830: inst = 32'd471859200;
      53831: inst = 32'd136314880;
      53832: inst = 32'd268468224;
      53833: inst = 32'd201347565;
      53834: inst = 32'd203423744;
      53835: inst = 32'd471859200;
      53836: inst = 32'd136314880;
      53837: inst = 32'd268468224;
      53838: inst = 32'd201347566;
      53839: inst = 32'd203423744;
      53840: inst = 32'd471859200;
      53841: inst = 32'd136314880;
      53842: inst = 32'd268468224;
      53843: inst = 32'd201347567;
      53844: inst = 32'd203423744;
      53845: inst = 32'd471859200;
      53846: inst = 32'd136314880;
      53847: inst = 32'd268468224;
      53848: inst = 32'd201347568;
      53849: inst = 32'd203423744;
      53850: inst = 32'd471859200;
      53851: inst = 32'd136314880;
      53852: inst = 32'd268468224;
      53853: inst = 32'd201347569;
      53854: inst = 32'd203423744;
      53855: inst = 32'd471859200;
      53856: inst = 32'd136314880;
      53857: inst = 32'd268468224;
      53858: inst = 32'd201347570;
      53859: inst = 32'd203423744;
      53860: inst = 32'd471859200;
      53861: inst = 32'd136314880;
      53862: inst = 32'd268468224;
      53863: inst = 32'd201347571;
      53864: inst = 32'd203423744;
      53865: inst = 32'd471859200;
      53866: inst = 32'd136314880;
      53867: inst = 32'd268468224;
      53868: inst = 32'd201347572;
      53869: inst = 32'd203423744;
      53870: inst = 32'd471859200;
      53871: inst = 32'd136314880;
      53872: inst = 32'd268468224;
      53873: inst = 32'd201347573;
      53874: inst = 32'd203423744;
      53875: inst = 32'd471859200;
      53876: inst = 32'd136314880;
      53877: inst = 32'd268468224;
      53878: inst = 32'd201347574;
      53879: inst = 32'd203423744;
      53880: inst = 32'd471859200;
      53881: inst = 32'd136314880;
      53882: inst = 32'd268468224;
      53883: inst = 32'd201347575;
      53884: inst = 32'd203423744;
      53885: inst = 32'd471859200;
      53886: inst = 32'd136314880;
      53887: inst = 32'd268468224;
      53888: inst = 32'd201347576;
      53889: inst = 32'd203423744;
      53890: inst = 32'd471859200;
      53891: inst = 32'd136314880;
      53892: inst = 32'd268468224;
      53893: inst = 32'd201347577;
      53894: inst = 32'd203423744;
      53895: inst = 32'd471859200;
      53896: inst = 32'd136314880;
      53897: inst = 32'd268468224;
      53898: inst = 32'd201347578;
      53899: inst = 32'd203423744;
      53900: inst = 32'd471859200;
      53901: inst = 32'd136314880;
      53902: inst = 32'd268468224;
      53903: inst = 32'd201347579;
      53904: inst = 32'd203423744;
      53905: inst = 32'd471859200;
      53906: inst = 32'd136314880;
      53907: inst = 32'd268468224;
      53908: inst = 32'd201347580;
      53909: inst = 32'd203423744;
      53910: inst = 32'd471859200;
      53911: inst = 32'd136314880;
      53912: inst = 32'd268468224;
      53913: inst = 32'd201347581;
      53914: inst = 32'd203423744;
      53915: inst = 32'd471859200;
      53916: inst = 32'd136314880;
      53917: inst = 32'd268468224;
      53918: inst = 32'd201347582;
      53919: inst = 32'd203423744;
      53920: inst = 32'd471859200;
      53921: inst = 32'd136314880;
      53922: inst = 32'd268468224;
      53923: inst = 32'd201347583;
      53924: inst = 32'd203423744;
      53925: inst = 32'd471859200;
      53926: inst = 32'd136314880;
      53927: inst = 32'd268468224;
      53928: inst = 32'd201347584;
      53929: inst = 32'd203423744;
      53930: inst = 32'd471859200;
      53931: inst = 32'd136314880;
      53932: inst = 32'd268468224;
      53933: inst = 32'd201347585;
      53934: inst = 32'd203423744;
      53935: inst = 32'd471859200;
      53936: inst = 32'd136314880;
      53937: inst = 32'd268468224;
      53938: inst = 32'd201347586;
      53939: inst = 32'd203423744;
      53940: inst = 32'd471859200;
      53941: inst = 32'd136314880;
      53942: inst = 32'd268468224;
      53943: inst = 32'd201347587;
      53944: inst = 32'd203423744;
      53945: inst = 32'd471859200;
      53946: inst = 32'd136314880;
      53947: inst = 32'd268468224;
      53948: inst = 32'd201347588;
      53949: inst = 32'd203423744;
      53950: inst = 32'd471859200;
      53951: inst = 32'd136314880;
      53952: inst = 32'd268468224;
      53953: inst = 32'd201347589;
      53954: inst = 32'd203423744;
      53955: inst = 32'd471859200;
      53956: inst = 32'd136314880;
      53957: inst = 32'd268468224;
      53958: inst = 32'd201347590;
      53959: inst = 32'd203423744;
      53960: inst = 32'd471859200;
      53961: inst = 32'd136314880;
      53962: inst = 32'd268468224;
      53963: inst = 32'd201347591;
      53964: inst = 32'd203423744;
      53965: inst = 32'd471859200;
      53966: inst = 32'd136314880;
      53967: inst = 32'd268468224;
      53968: inst = 32'd201347592;
      53969: inst = 32'd203423744;
      53970: inst = 32'd471859200;
      53971: inst = 32'd136314880;
      53972: inst = 32'd268468224;
      53973: inst = 32'd201347593;
      53974: inst = 32'd203423744;
      53975: inst = 32'd471859200;
      53976: inst = 32'd136314880;
      53977: inst = 32'd268468224;
      53978: inst = 32'd201347594;
      53979: inst = 32'd203423744;
      53980: inst = 32'd471859200;
      53981: inst = 32'd136314880;
      53982: inst = 32'd268468224;
      53983: inst = 32'd201347595;
      53984: inst = 32'd203423744;
      53985: inst = 32'd471859200;
      53986: inst = 32'd136314880;
      53987: inst = 32'd268468224;
      53988: inst = 32'd201347596;
      53989: inst = 32'd203423744;
      53990: inst = 32'd471859200;
      53991: inst = 32'd136314880;
      53992: inst = 32'd268468224;
      53993: inst = 32'd201347597;
      53994: inst = 32'd203423744;
      53995: inst = 32'd471859200;
      53996: inst = 32'd136314880;
      53997: inst = 32'd268468224;
      53998: inst = 32'd201347598;
      53999: inst = 32'd203423744;
      54000: inst = 32'd471859200;
      54001: inst = 32'd136314880;
      54002: inst = 32'd268468224;
      54003: inst = 32'd201347599;
      54004: inst = 32'd203423744;
      54005: inst = 32'd471859200;
      54006: inst = 32'd136314880;
      54007: inst = 32'd268468224;
      54008: inst = 32'd201347600;
      54009: inst = 32'd203423744;
      54010: inst = 32'd471859200;
      54011: inst = 32'd136314880;
      54012: inst = 32'd268468224;
      54013: inst = 32'd201347601;
      54014: inst = 32'd203423744;
      54015: inst = 32'd471859200;
      54016: inst = 32'd136314880;
      54017: inst = 32'd268468224;
      54018: inst = 32'd201347602;
      54019: inst = 32'd203423744;
      54020: inst = 32'd471859200;
      54021: inst = 32'd136314880;
      54022: inst = 32'd268468224;
      54023: inst = 32'd201347603;
      54024: inst = 32'd203423744;
      54025: inst = 32'd471859200;
      54026: inst = 32'd136314880;
      54027: inst = 32'd268468224;
      54028: inst = 32'd201347604;
      54029: inst = 32'd203423744;
      54030: inst = 32'd471859200;
      54031: inst = 32'd136314880;
      54032: inst = 32'd268468224;
      54033: inst = 32'd201347605;
      54034: inst = 32'd203423744;
      54035: inst = 32'd471859200;
      54036: inst = 32'd136314880;
      54037: inst = 32'd268468224;
      54038: inst = 32'd201347606;
      54039: inst = 32'd203423744;
      54040: inst = 32'd471859200;
      54041: inst = 32'd136314880;
      54042: inst = 32'd268468224;
      54043: inst = 32'd201347607;
      54044: inst = 32'd203423744;
      54045: inst = 32'd471859200;
      54046: inst = 32'd136314880;
      54047: inst = 32'd268468224;
      54048: inst = 32'd201347608;
      54049: inst = 32'd203423744;
      54050: inst = 32'd471859200;
      54051: inst = 32'd136314880;
      54052: inst = 32'd268468224;
      54053: inst = 32'd201347609;
      54054: inst = 32'd203423744;
      54055: inst = 32'd471859200;
      54056: inst = 32'd136314880;
      54057: inst = 32'd268468224;
      54058: inst = 32'd201347610;
      54059: inst = 32'd203423744;
      54060: inst = 32'd471859200;
      54061: inst = 32'd136314880;
      54062: inst = 32'd268468224;
      54063: inst = 32'd201347611;
      54064: inst = 32'd203423744;
      54065: inst = 32'd471859200;
      54066: inst = 32'd136314880;
      54067: inst = 32'd268468224;
      54068: inst = 32'd201347612;
      54069: inst = 32'd203423744;
      54070: inst = 32'd471859200;
      54071: inst = 32'd136314880;
      54072: inst = 32'd268468224;
      54073: inst = 32'd201347613;
      54074: inst = 32'd203423744;
      54075: inst = 32'd471859200;
      54076: inst = 32'd136314880;
      54077: inst = 32'd268468224;
      54078: inst = 32'd201347614;
      54079: inst = 32'd203423744;
      54080: inst = 32'd471859200;
      54081: inst = 32'd136314880;
      54082: inst = 32'd268468224;
      54083: inst = 32'd201347615;
      54084: inst = 32'd203423744;
      54085: inst = 32'd471859200;
      54086: inst = 32'd136314880;
      54087: inst = 32'd268468224;
      54088: inst = 32'd201347616;
      54089: inst = 32'd203423744;
      54090: inst = 32'd471859200;
      54091: inst = 32'd136314880;
      54092: inst = 32'd268468224;
      54093: inst = 32'd201347617;
      54094: inst = 32'd203423744;
      54095: inst = 32'd471859200;
      54096: inst = 32'd136314880;
      54097: inst = 32'd268468224;
      54098: inst = 32'd201347618;
      54099: inst = 32'd203423744;
      54100: inst = 32'd471859200;
      54101: inst = 32'd136314880;
      54102: inst = 32'd268468224;
      54103: inst = 32'd201347619;
      54104: inst = 32'd203423744;
      54105: inst = 32'd471859200;
      54106: inst = 32'd136314880;
      54107: inst = 32'd268468224;
      54108: inst = 32'd201347620;
      54109: inst = 32'd203423744;
      54110: inst = 32'd471859200;
      54111: inst = 32'd136314880;
      54112: inst = 32'd268468224;
      54113: inst = 32'd201347621;
      54114: inst = 32'd203423744;
      54115: inst = 32'd471859200;
      54116: inst = 32'd136314880;
      54117: inst = 32'd268468224;
      54118: inst = 32'd201347622;
      54119: inst = 32'd203423744;
      54120: inst = 32'd471859200;
      54121: inst = 32'd136314880;
      54122: inst = 32'd268468224;
      54123: inst = 32'd201347623;
      54124: inst = 32'd203423744;
      54125: inst = 32'd471859200;
      54126: inst = 32'd136314880;
      54127: inst = 32'd268468224;
      54128: inst = 32'd201347624;
      54129: inst = 32'd203423744;
      54130: inst = 32'd471859200;
      54131: inst = 32'd136314880;
      54132: inst = 32'd268468224;
      54133: inst = 32'd201347625;
      54134: inst = 32'd203423744;
      54135: inst = 32'd471859200;
      54136: inst = 32'd136314880;
      54137: inst = 32'd268468224;
      54138: inst = 32'd201347626;
      54139: inst = 32'd203423744;
      54140: inst = 32'd471859200;
      54141: inst = 32'd136314880;
      54142: inst = 32'd268468224;
      54143: inst = 32'd201347627;
      54144: inst = 32'd203423744;
      54145: inst = 32'd471859200;
      54146: inst = 32'd136314880;
      54147: inst = 32'd268468224;
      54148: inst = 32'd201347628;
      54149: inst = 32'd203423744;
      54150: inst = 32'd471859200;
      54151: inst = 32'd136314880;
      54152: inst = 32'd268468224;
      54153: inst = 32'd201347629;
      54154: inst = 32'd203423744;
      54155: inst = 32'd471859200;
      54156: inst = 32'd136314880;
      54157: inst = 32'd268468224;
      54158: inst = 32'd201347630;
      54159: inst = 32'd203423744;
      54160: inst = 32'd471859200;
      54161: inst = 32'd136314880;
      54162: inst = 32'd268468224;
      54163: inst = 32'd201347631;
      54164: inst = 32'd203423744;
      54165: inst = 32'd471859200;
      54166: inst = 32'd136314880;
      54167: inst = 32'd268468224;
      54168: inst = 32'd201347632;
      54169: inst = 32'd203423744;
      54170: inst = 32'd471859200;
      54171: inst = 32'd136314880;
      54172: inst = 32'd268468224;
      54173: inst = 32'd201347633;
      54174: inst = 32'd203423744;
      54175: inst = 32'd471859200;
      54176: inst = 32'd136314880;
      54177: inst = 32'd268468224;
      54178: inst = 32'd201347634;
      54179: inst = 32'd203423744;
      54180: inst = 32'd471859200;
      54181: inst = 32'd136314880;
      54182: inst = 32'd268468224;
      54183: inst = 32'd201347635;
      54184: inst = 32'd203423744;
      54185: inst = 32'd471859200;
      54186: inst = 32'd136314880;
      54187: inst = 32'd268468224;
      54188: inst = 32'd201347636;
      54189: inst = 32'd203423744;
      54190: inst = 32'd471859200;
      54191: inst = 32'd136314880;
      54192: inst = 32'd268468224;
      54193: inst = 32'd201347637;
      54194: inst = 32'd203423744;
      54195: inst = 32'd471859200;
      54196: inst = 32'd136314880;
      54197: inst = 32'd268468224;
      54198: inst = 32'd201347638;
      54199: inst = 32'd203423744;
      54200: inst = 32'd471859200;
      54201: inst = 32'd136314880;
      54202: inst = 32'd268468224;
      54203: inst = 32'd201347639;
      54204: inst = 32'd203423744;
      54205: inst = 32'd471859200;
      54206: inst = 32'd136314880;
      54207: inst = 32'd268468224;
      54208: inst = 32'd201347640;
      54209: inst = 32'd203423744;
      54210: inst = 32'd471859200;
      54211: inst = 32'd136314880;
      54212: inst = 32'd268468224;
      54213: inst = 32'd201347641;
      54214: inst = 32'd203423744;
      54215: inst = 32'd471859200;
      54216: inst = 32'd136314880;
      54217: inst = 32'd268468224;
      54218: inst = 32'd201347642;
      54219: inst = 32'd203423744;
      54220: inst = 32'd471859200;
      54221: inst = 32'd136314880;
      54222: inst = 32'd268468224;
      54223: inst = 32'd201347643;
      54224: inst = 32'd203423744;
      54225: inst = 32'd471859200;
      54226: inst = 32'd136314880;
      54227: inst = 32'd268468224;
      54228: inst = 32'd201347644;
      54229: inst = 32'd203423744;
      54230: inst = 32'd471859200;
      54231: inst = 32'd136314880;
      54232: inst = 32'd268468224;
      54233: inst = 32'd201347645;
      54234: inst = 32'd203423744;
      54235: inst = 32'd471859200;
      54236: inst = 32'd136314880;
      54237: inst = 32'd268468224;
      54238: inst = 32'd201347646;
      54239: inst = 32'd203423744;
      54240: inst = 32'd471859200;
      54241: inst = 32'd136314880;
      54242: inst = 32'd268468224;
      54243: inst = 32'd201347647;
      54244: inst = 32'd203423744;
      54245: inst = 32'd471859200;
      54246: inst = 32'd136314880;
      54247: inst = 32'd268468224;
      54248: inst = 32'd201347648;
      54249: inst = 32'd203423744;
      54250: inst = 32'd471859200;
      54251: inst = 32'd136314880;
      54252: inst = 32'd268468224;
      54253: inst = 32'd201347649;
      54254: inst = 32'd203423744;
      54255: inst = 32'd471859200;
      54256: inst = 32'd136314880;
      54257: inst = 32'd268468224;
      54258: inst = 32'd201347650;
      54259: inst = 32'd203423744;
      54260: inst = 32'd471859200;
      54261: inst = 32'd136314880;
      54262: inst = 32'd268468224;
      54263: inst = 32'd201347651;
      54264: inst = 32'd203423744;
      54265: inst = 32'd471859200;
      54266: inst = 32'd136314880;
      54267: inst = 32'd268468224;
      54268: inst = 32'd201347652;
      54269: inst = 32'd203423744;
      54270: inst = 32'd471859200;
      54271: inst = 32'd136314880;
      54272: inst = 32'd268468224;
      54273: inst = 32'd201347653;
      54274: inst = 32'd203423744;
      54275: inst = 32'd471859200;
      54276: inst = 32'd136314880;
      54277: inst = 32'd268468224;
      54278: inst = 32'd201347654;
      54279: inst = 32'd203423744;
      54280: inst = 32'd471859200;
      54281: inst = 32'd136314880;
      54282: inst = 32'd268468224;
      54283: inst = 32'd201347655;
      54284: inst = 32'd203423744;
      54285: inst = 32'd471859200;
      54286: inst = 32'd136314880;
      54287: inst = 32'd268468224;
      54288: inst = 32'd201347656;
      54289: inst = 32'd203423744;
      54290: inst = 32'd471859200;
      54291: inst = 32'd136314880;
      54292: inst = 32'd268468224;
      54293: inst = 32'd201347657;
      54294: inst = 32'd203423744;
      54295: inst = 32'd471859200;
      54296: inst = 32'd136314880;
      54297: inst = 32'd268468224;
      54298: inst = 32'd201347658;
      54299: inst = 32'd203423744;
      54300: inst = 32'd471859200;
      54301: inst = 32'd136314880;
      54302: inst = 32'd268468224;
      54303: inst = 32'd201347659;
      54304: inst = 32'd203423744;
      54305: inst = 32'd471859200;
      54306: inst = 32'd136314880;
      54307: inst = 32'd268468224;
      54308: inst = 32'd201347660;
      54309: inst = 32'd203423744;
      54310: inst = 32'd471859200;
      54311: inst = 32'd136314880;
      54312: inst = 32'd268468224;
      54313: inst = 32'd201347661;
      54314: inst = 32'd203423744;
      54315: inst = 32'd471859200;
      54316: inst = 32'd136314880;
      54317: inst = 32'd268468224;
      54318: inst = 32'd201347662;
      54319: inst = 32'd203423744;
      54320: inst = 32'd471859200;
      54321: inst = 32'd136314880;
      54322: inst = 32'd268468224;
      54323: inst = 32'd201347663;
      54324: inst = 32'd203423744;
      54325: inst = 32'd471859200;
      54326: inst = 32'd136314880;
      54327: inst = 32'd268468224;
      54328: inst = 32'd201347664;
      54329: inst = 32'd203423744;
      54330: inst = 32'd471859200;
      54331: inst = 32'd136314880;
      54332: inst = 32'd268468224;
      54333: inst = 32'd201347665;
      54334: inst = 32'd203423744;
      54335: inst = 32'd471859200;
      54336: inst = 32'd136314880;
      54337: inst = 32'd268468224;
      54338: inst = 32'd201347666;
      54339: inst = 32'd203423744;
      54340: inst = 32'd471859200;
      54341: inst = 32'd136314880;
      54342: inst = 32'd268468224;
      54343: inst = 32'd201347667;
      54344: inst = 32'd203423744;
      54345: inst = 32'd471859200;
      54346: inst = 32'd136314880;
      54347: inst = 32'd268468224;
      54348: inst = 32'd201347668;
      54349: inst = 32'd203423744;
      54350: inst = 32'd471859200;
      54351: inst = 32'd136314880;
      54352: inst = 32'd268468224;
      54353: inst = 32'd201347669;
      54354: inst = 32'd203423744;
      54355: inst = 32'd471859200;
      54356: inst = 32'd136314880;
      54357: inst = 32'd268468224;
      54358: inst = 32'd201347670;
      54359: inst = 32'd203423744;
      54360: inst = 32'd471859200;
      54361: inst = 32'd136314880;
      54362: inst = 32'd268468224;
      54363: inst = 32'd201347671;
      54364: inst = 32'd203423744;
      54365: inst = 32'd471859200;
      54366: inst = 32'd136314880;
      54367: inst = 32'd268468224;
      54368: inst = 32'd201347672;
      54369: inst = 32'd203423744;
      54370: inst = 32'd471859200;
      54371: inst = 32'd136314880;
      54372: inst = 32'd268468224;
      54373: inst = 32'd201347673;
      54374: inst = 32'd203423744;
      54375: inst = 32'd471859200;
      54376: inst = 32'd136314880;
      54377: inst = 32'd268468224;
      54378: inst = 32'd201347674;
      54379: inst = 32'd203423744;
      54380: inst = 32'd471859200;
      54381: inst = 32'd136314880;
      54382: inst = 32'd268468224;
      54383: inst = 32'd201347675;
      54384: inst = 32'd203423744;
      54385: inst = 32'd471859200;
      54386: inst = 32'd136314880;
      54387: inst = 32'd268468224;
      54388: inst = 32'd201347676;
      54389: inst = 32'd203423744;
      54390: inst = 32'd471859200;
      54391: inst = 32'd136314880;
      54392: inst = 32'd268468224;
      54393: inst = 32'd201347677;
      54394: inst = 32'd203423744;
      54395: inst = 32'd471859200;
      54396: inst = 32'd136314880;
      54397: inst = 32'd268468224;
      54398: inst = 32'd201347678;
      54399: inst = 32'd203423744;
      54400: inst = 32'd471859200;
      54401: inst = 32'd136314880;
      54402: inst = 32'd268468224;
      54403: inst = 32'd201347679;
      54404: inst = 32'd203423744;
      54405: inst = 32'd471859200;
      54406: inst = 32'd136314880;
      54407: inst = 32'd268468224;
      54408: inst = 32'd201347680;
      54409: inst = 32'd203423744;
      54410: inst = 32'd471859200;
      54411: inst = 32'd136314880;
      54412: inst = 32'd268468224;
      54413: inst = 32'd201347681;
      54414: inst = 32'd203423744;
      54415: inst = 32'd471859200;
      54416: inst = 32'd136314880;
      54417: inst = 32'd268468224;
      54418: inst = 32'd201347682;
      54419: inst = 32'd203423744;
      54420: inst = 32'd471859200;
      54421: inst = 32'd136314880;
      54422: inst = 32'd268468224;
      54423: inst = 32'd201347683;
      54424: inst = 32'd203423744;
      54425: inst = 32'd471859200;
      54426: inst = 32'd136314880;
      54427: inst = 32'd268468224;
      54428: inst = 32'd201347684;
      54429: inst = 32'd203423744;
      54430: inst = 32'd471859200;
      54431: inst = 32'd136314880;
      54432: inst = 32'd268468224;
      54433: inst = 32'd201347685;
      54434: inst = 32'd203423744;
      54435: inst = 32'd471859200;
      54436: inst = 32'd136314880;
      54437: inst = 32'd268468224;
      54438: inst = 32'd201347686;
      54439: inst = 32'd203423744;
      54440: inst = 32'd471859200;
      54441: inst = 32'd136314880;
      54442: inst = 32'd268468224;
      54443: inst = 32'd201347687;
      54444: inst = 32'd203423744;
      54445: inst = 32'd471859200;
      54446: inst = 32'd136314880;
      54447: inst = 32'd268468224;
      54448: inst = 32'd201347688;
      54449: inst = 32'd203423744;
      54450: inst = 32'd471859200;
      54451: inst = 32'd136314880;
      54452: inst = 32'd268468224;
      54453: inst = 32'd201347689;
      54454: inst = 32'd203423744;
      54455: inst = 32'd471859200;
      54456: inst = 32'd136314880;
      54457: inst = 32'd268468224;
      54458: inst = 32'd201347690;
      54459: inst = 32'd203423744;
      54460: inst = 32'd471859200;
      54461: inst = 32'd136314880;
      54462: inst = 32'd268468224;
      54463: inst = 32'd201347691;
      54464: inst = 32'd203423744;
      54465: inst = 32'd471859200;
      54466: inst = 32'd136314880;
      54467: inst = 32'd268468224;
      54468: inst = 32'd201347692;
      54469: inst = 32'd203423744;
      54470: inst = 32'd471859200;
      54471: inst = 32'd136314880;
      54472: inst = 32'd268468224;
      54473: inst = 32'd201347693;
      54474: inst = 32'd203423744;
      54475: inst = 32'd471859200;
      54476: inst = 32'd136314880;
      54477: inst = 32'd268468224;
      54478: inst = 32'd201347694;
      54479: inst = 32'd203423744;
      54480: inst = 32'd471859200;
      54481: inst = 32'd136314880;
      54482: inst = 32'd268468224;
      54483: inst = 32'd201347695;
      54484: inst = 32'd203423744;
      54485: inst = 32'd471859200;
      54486: inst = 32'd136314880;
      54487: inst = 32'd268468224;
      54488: inst = 32'd201347696;
      54489: inst = 32'd203423744;
      54490: inst = 32'd471859200;
      54491: inst = 32'd136314880;
      54492: inst = 32'd268468224;
      54493: inst = 32'd201347697;
      54494: inst = 32'd203423744;
      54495: inst = 32'd471859200;
      54496: inst = 32'd136314880;
      54497: inst = 32'd268468224;
      54498: inst = 32'd201347698;
      54499: inst = 32'd203423744;
      54500: inst = 32'd471859200;
      54501: inst = 32'd136314880;
      54502: inst = 32'd268468224;
      54503: inst = 32'd201347699;
      54504: inst = 32'd203423744;
      54505: inst = 32'd471859200;
      54506: inst = 32'd136314880;
      54507: inst = 32'd268468224;
      54508: inst = 32'd201347700;
      54509: inst = 32'd203423744;
      54510: inst = 32'd471859200;
      54511: inst = 32'd136314880;
      54512: inst = 32'd268468224;
      54513: inst = 32'd201347701;
      54514: inst = 32'd203423744;
      54515: inst = 32'd471859200;
      54516: inst = 32'd136314880;
      54517: inst = 32'd268468224;
      54518: inst = 32'd201347702;
      54519: inst = 32'd203423744;
      54520: inst = 32'd471859200;
      54521: inst = 32'd136314880;
      54522: inst = 32'd268468224;
      54523: inst = 32'd201347703;
      54524: inst = 32'd203423744;
      54525: inst = 32'd471859200;
      54526: inst = 32'd136314880;
      54527: inst = 32'd268468224;
      54528: inst = 32'd201347704;
      54529: inst = 32'd203423744;
      54530: inst = 32'd471859200;
      54531: inst = 32'd136314880;
      54532: inst = 32'd268468224;
      54533: inst = 32'd201347705;
      54534: inst = 32'd203423744;
      54535: inst = 32'd471859200;
      54536: inst = 32'd136314880;
      54537: inst = 32'd268468224;
      54538: inst = 32'd201347706;
      54539: inst = 32'd203423744;
      54540: inst = 32'd471859200;
      54541: inst = 32'd136314880;
      54542: inst = 32'd268468224;
      54543: inst = 32'd201347707;
      54544: inst = 32'd203423744;
      54545: inst = 32'd471859200;
      54546: inst = 32'd136314880;
      54547: inst = 32'd268468224;
      54548: inst = 32'd201347708;
      54549: inst = 32'd203423744;
      54550: inst = 32'd471859200;
      54551: inst = 32'd136314880;
      54552: inst = 32'd268468224;
      54553: inst = 32'd201347709;
      54554: inst = 32'd203423744;
      54555: inst = 32'd471859200;
      54556: inst = 32'd136314880;
      54557: inst = 32'd268468224;
      54558: inst = 32'd201347710;
      54559: inst = 32'd203423744;
      54560: inst = 32'd471859200;
      54561: inst = 32'd136314880;
      54562: inst = 32'd268468224;
      54563: inst = 32'd201347711;
      54564: inst = 32'd203423744;
      54565: inst = 32'd471859200;
      54566: inst = 32'd136314880;
      54567: inst = 32'd268468224;
      54568: inst = 32'd201347712;
      54569: inst = 32'd203423744;
      54570: inst = 32'd471859200;
      54571: inst = 32'd136314880;
      54572: inst = 32'd268468224;
      54573: inst = 32'd201347713;
      54574: inst = 32'd203423744;
      54575: inst = 32'd471859200;
      54576: inst = 32'd136314880;
      54577: inst = 32'd268468224;
      54578: inst = 32'd201347714;
      54579: inst = 32'd203423744;
      54580: inst = 32'd471859200;
      54581: inst = 32'd136314880;
      54582: inst = 32'd268468224;
      54583: inst = 32'd201347715;
      54584: inst = 32'd203423744;
      54585: inst = 32'd471859200;
      54586: inst = 32'd136314880;
      54587: inst = 32'd268468224;
      54588: inst = 32'd201347716;
      54589: inst = 32'd203423744;
      54590: inst = 32'd471859200;
      54591: inst = 32'd136314880;
      54592: inst = 32'd268468224;
      54593: inst = 32'd201347717;
      54594: inst = 32'd203423744;
      54595: inst = 32'd471859200;
      54596: inst = 32'd136314880;
      54597: inst = 32'd268468224;
      54598: inst = 32'd201347718;
      54599: inst = 32'd203423744;
      54600: inst = 32'd471859200;
      54601: inst = 32'd136314880;
      54602: inst = 32'd268468224;
      54603: inst = 32'd201347719;
      54604: inst = 32'd203423744;
      54605: inst = 32'd471859200;
      54606: inst = 32'd136314880;
      54607: inst = 32'd268468224;
      54608: inst = 32'd201347720;
      54609: inst = 32'd203423744;
      54610: inst = 32'd471859200;
      54611: inst = 32'd136314880;
      54612: inst = 32'd268468224;
      54613: inst = 32'd201347721;
      54614: inst = 32'd203423744;
      54615: inst = 32'd471859200;
      54616: inst = 32'd136314880;
      54617: inst = 32'd268468224;
      54618: inst = 32'd201347722;
      54619: inst = 32'd203423744;
      54620: inst = 32'd471859200;
      54621: inst = 32'd136314880;
      54622: inst = 32'd268468224;
      54623: inst = 32'd201347723;
      54624: inst = 32'd203423744;
      54625: inst = 32'd471859200;
      54626: inst = 32'd136314880;
      54627: inst = 32'd268468224;
      54628: inst = 32'd201347724;
      54629: inst = 32'd203423744;
      54630: inst = 32'd471859200;
      54631: inst = 32'd136314880;
      54632: inst = 32'd268468224;
      54633: inst = 32'd201347725;
      54634: inst = 32'd203423744;
      54635: inst = 32'd471859200;
      54636: inst = 32'd136314880;
      54637: inst = 32'd268468224;
      54638: inst = 32'd201347726;
      54639: inst = 32'd203423744;
      54640: inst = 32'd471859200;
      54641: inst = 32'd136314880;
      54642: inst = 32'd268468224;
      54643: inst = 32'd201347727;
      54644: inst = 32'd203423744;
      54645: inst = 32'd471859200;
      54646: inst = 32'd136314880;
      54647: inst = 32'd268468224;
      54648: inst = 32'd201347728;
      54649: inst = 32'd203423744;
      54650: inst = 32'd471859200;
      54651: inst = 32'd136314880;
      54652: inst = 32'd268468224;
      54653: inst = 32'd201347729;
      54654: inst = 32'd203423744;
      54655: inst = 32'd471859200;
      54656: inst = 32'd136314880;
      54657: inst = 32'd268468224;
      54658: inst = 32'd201347730;
      54659: inst = 32'd203423744;
      54660: inst = 32'd471859200;
      54661: inst = 32'd136314880;
      54662: inst = 32'd268468224;
      54663: inst = 32'd201347731;
      54664: inst = 32'd203423744;
      54665: inst = 32'd471859200;
      54666: inst = 32'd136314880;
      54667: inst = 32'd268468224;
      54668: inst = 32'd201347732;
      54669: inst = 32'd203423744;
      54670: inst = 32'd471859200;
      54671: inst = 32'd136314880;
      54672: inst = 32'd268468224;
      54673: inst = 32'd201347733;
      54674: inst = 32'd203423744;
      54675: inst = 32'd471859200;
      54676: inst = 32'd136314880;
      54677: inst = 32'd268468224;
      54678: inst = 32'd201347734;
      54679: inst = 32'd203423744;
      54680: inst = 32'd471859200;
      54681: inst = 32'd136314880;
      54682: inst = 32'd268468224;
      54683: inst = 32'd201347735;
      54684: inst = 32'd203423744;
      54685: inst = 32'd471859200;
      54686: inst = 32'd136314880;
      54687: inst = 32'd268468224;
      54688: inst = 32'd201347736;
      54689: inst = 32'd203423744;
      54690: inst = 32'd471859200;
      54691: inst = 32'd136314880;
      54692: inst = 32'd268468224;
      54693: inst = 32'd201347737;
      54694: inst = 32'd203423744;
      54695: inst = 32'd471859200;
      54696: inst = 32'd136314880;
      54697: inst = 32'd268468224;
      54698: inst = 32'd201347738;
      54699: inst = 32'd203423744;
      54700: inst = 32'd471859200;
      54701: inst = 32'd136314880;
      54702: inst = 32'd268468224;
      54703: inst = 32'd201347739;
      54704: inst = 32'd203423744;
      54705: inst = 32'd471859200;
      54706: inst = 32'd136314880;
      54707: inst = 32'd268468224;
      54708: inst = 32'd201347740;
      54709: inst = 32'd203423744;
      54710: inst = 32'd471859200;
      54711: inst = 32'd136314880;
      54712: inst = 32'd268468224;
      54713: inst = 32'd201347741;
      54714: inst = 32'd203423744;
      54715: inst = 32'd471859200;
      54716: inst = 32'd136314880;
      54717: inst = 32'd268468224;
      54718: inst = 32'd201347742;
      54719: inst = 32'd203423744;
      54720: inst = 32'd471859200;
      54721: inst = 32'd136314880;
      54722: inst = 32'd268468224;
      54723: inst = 32'd201347743;
      54724: inst = 32'd203423744;
      54725: inst = 32'd471859200;
      54726: inst = 32'd136314880;
      54727: inst = 32'd268468224;
      54728: inst = 32'd201347744;
      54729: inst = 32'd203423744;
      54730: inst = 32'd471859200;
      54731: inst = 32'd136314880;
      54732: inst = 32'd268468224;
      54733: inst = 32'd201347745;
      54734: inst = 32'd203423744;
      54735: inst = 32'd471859200;
      54736: inst = 32'd136314880;
      54737: inst = 32'd268468224;
      54738: inst = 32'd201347746;
      54739: inst = 32'd203423744;
      54740: inst = 32'd471859200;
      54741: inst = 32'd136314880;
      54742: inst = 32'd268468224;
      54743: inst = 32'd201347747;
      54744: inst = 32'd203423744;
      54745: inst = 32'd471859200;
      54746: inst = 32'd136314880;
      54747: inst = 32'd268468224;
      54748: inst = 32'd201347748;
      54749: inst = 32'd203423744;
      54750: inst = 32'd471859200;
      54751: inst = 32'd136314880;
      54752: inst = 32'd268468224;
      54753: inst = 32'd201347749;
      54754: inst = 32'd203423744;
      54755: inst = 32'd471859200;
      54756: inst = 32'd136314880;
      54757: inst = 32'd268468224;
      54758: inst = 32'd201347750;
      54759: inst = 32'd203423744;
      54760: inst = 32'd471859200;
      54761: inst = 32'd136314880;
      54762: inst = 32'd268468224;
      54763: inst = 32'd201347751;
      54764: inst = 32'd203423744;
      54765: inst = 32'd471859200;
      54766: inst = 32'd136314880;
      54767: inst = 32'd268468224;
      54768: inst = 32'd201347752;
      54769: inst = 32'd203423744;
      54770: inst = 32'd471859200;
      54771: inst = 32'd136314880;
      54772: inst = 32'd268468224;
      54773: inst = 32'd201347753;
      54774: inst = 32'd203423744;
      54775: inst = 32'd471859200;
      54776: inst = 32'd136314880;
      54777: inst = 32'd268468224;
      54778: inst = 32'd201347754;
      54779: inst = 32'd203423744;
      54780: inst = 32'd471859200;
      54781: inst = 32'd136314880;
      54782: inst = 32'd268468224;
      54783: inst = 32'd201347755;
      54784: inst = 32'd203423744;
      54785: inst = 32'd471859200;
      54786: inst = 32'd136314880;
      54787: inst = 32'd268468224;
      54788: inst = 32'd201347756;
      54789: inst = 32'd203423744;
      54790: inst = 32'd471859200;
      54791: inst = 32'd136314880;
      54792: inst = 32'd268468224;
      54793: inst = 32'd201347757;
      54794: inst = 32'd203423744;
      54795: inst = 32'd471859200;
      54796: inst = 32'd136314880;
      54797: inst = 32'd268468224;
      54798: inst = 32'd201347758;
      54799: inst = 32'd203423744;
      54800: inst = 32'd471859200;
      54801: inst = 32'd136314880;
      54802: inst = 32'd268468224;
      54803: inst = 32'd201347759;
      54804: inst = 32'd203423744;
      54805: inst = 32'd471859200;
      54806: inst = 32'd136314880;
      54807: inst = 32'd268468224;
      54808: inst = 32'd201347760;
      54809: inst = 32'd203423744;
      54810: inst = 32'd471859200;
      54811: inst = 32'd136314880;
      54812: inst = 32'd268468224;
      54813: inst = 32'd201347761;
      54814: inst = 32'd203423744;
      54815: inst = 32'd471859200;
      54816: inst = 32'd136314880;
      54817: inst = 32'd268468224;
      54818: inst = 32'd201347762;
      54819: inst = 32'd203423744;
      54820: inst = 32'd471859200;
      54821: inst = 32'd136314880;
      54822: inst = 32'd268468224;
      54823: inst = 32'd201347763;
      54824: inst = 32'd203423744;
      54825: inst = 32'd471859200;
      54826: inst = 32'd136314880;
      54827: inst = 32'd268468224;
      54828: inst = 32'd201347764;
      54829: inst = 32'd203423744;
      54830: inst = 32'd471859200;
      54831: inst = 32'd136314880;
      54832: inst = 32'd268468224;
      54833: inst = 32'd201347765;
      54834: inst = 32'd203423744;
      54835: inst = 32'd471859200;
      54836: inst = 32'd136314880;
      54837: inst = 32'd268468224;
      54838: inst = 32'd201347766;
      54839: inst = 32'd203423744;
      54840: inst = 32'd471859200;
      54841: inst = 32'd136314880;
      54842: inst = 32'd268468224;
      54843: inst = 32'd201347767;
      54844: inst = 32'd203423744;
      54845: inst = 32'd471859200;
      54846: inst = 32'd136314880;
      54847: inst = 32'd268468224;
      54848: inst = 32'd201347768;
      54849: inst = 32'd203423744;
      54850: inst = 32'd471859200;
      54851: inst = 32'd136314880;
      54852: inst = 32'd268468224;
      54853: inst = 32'd201347769;
      54854: inst = 32'd203423744;
      54855: inst = 32'd471859200;
      54856: inst = 32'd136314880;
      54857: inst = 32'd268468224;
      54858: inst = 32'd201347770;
      54859: inst = 32'd203423744;
      54860: inst = 32'd471859200;
      54861: inst = 32'd136314880;
      54862: inst = 32'd268468224;
      54863: inst = 32'd201347771;
      54864: inst = 32'd203423744;
      54865: inst = 32'd471859200;
      54866: inst = 32'd136314880;
      54867: inst = 32'd268468224;
      54868: inst = 32'd201347772;
      54869: inst = 32'd203423744;
      54870: inst = 32'd471859200;
      54871: inst = 32'd136314880;
      54872: inst = 32'd268468224;
      54873: inst = 32'd201347773;
      54874: inst = 32'd203423744;
      54875: inst = 32'd471859200;
      54876: inst = 32'd136314880;
      54877: inst = 32'd268468224;
      54878: inst = 32'd201347774;
      54879: inst = 32'd203423744;
      54880: inst = 32'd471859200;
      54881: inst = 32'd136314880;
      54882: inst = 32'd268468224;
      54883: inst = 32'd201347775;
      54884: inst = 32'd203423744;
      54885: inst = 32'd471859200;
      54886: inst = 32'd136314880;
      54887: inst = 32'd268468224;
      54888: inst = 32'd201347776;
      54889: inst = 32'd203423744;
      54890: inst = 32'd471859200;
      54891: inst = 32'd136314880;
      54892: inst = 32'd268468224;
      54893: inst = 32'd201347777;
      54894: inst = 32'd203423744;
      54895: inst = 32'd471859200;
      54896: inst = 32'd136314880;
      54897: inst = 32'd268468224;
      54898: inst = 32'd201347778;
      54899: inst = 32'd203423744;
      54900: inst = 32'd471859200;
      54901: inst = 32'd136314880;
      54902: inst = 32'd268468224;
      54903: inst = 32'd201347779;
      54904: inst = 32'd203423744;
      54905: inst = 32'd471859200;
      54906: inst = 32'd136314880;
      54907: inst = 32'd268468224;
      54908: inst = 32'd201347780;
      54909: inst = 32'd203423744;
      54910: inst = 32'd471859200;
      54911: inst = 32'd136314880;
      54912: inst = 32'd268468224;
      54913: inst = 32'd201347781;
      54914: inst = 32'd203423744;
      54915: inst = 32'd471859200;
      54916: inst = 32'd136314880;
      54917: inst = 32'd268468224;
      54918: inst = 32'd201347782;
      54919: inst = 32'd203423744;
      54920: inst = 32'd471859200;
      54921: inst = 32'd136314880;
      54922: inst = 32'd268468224;
      54923: inst = 32'd201347783;
      54924: inst = 32'd203423744;
      54925: inst = 32'd471859200;
      54926: inst = 32'd136314880;
      54927: inst = 32'd268468224;
      54928: inst = 32'd201347784;
      54929: inst = 32'd203423744;
      54930: inst = 32'd471859200;
      54931: inst = 32'd136314880;
      54932: inst = 32'd268468224;
      54933: inst = 32'd201347785;
      54934: inst = 32'd203423744;
      54935: inst = 32'd471859200;
      54936: inst = 32'd136314880;
      54937: inst = 32'd268468224;
      54938: inst = 32'd201347786;
      54939: inst = 32'd203423744;
      54940: inst = 32'd471859200;
      54941: inst = 32'd136314880;
      54942: inst = 32'd268468224;
      54943: inst = 32'd201347787;
      54944: inst = 32'd203423744;
      54945: inst = 32'd471859200;
      54946: inst = 32'd136314880;
      54947: inst = 32'd268468224;
      54948: inst = 32'd201347788;
      54949: inst = 32'd203423744;
      54950: inst = 32'd471859200;
      54951: inst = 32'd136314880;
      54952: inst = 32'd268468224;
      54953: inst = 32'd201347789;
      54954: inst = 32'd203423744;
      54955: inst = 32'd471859200;
      54956: inst = 32'd136314880;
      54957: inst = 32'd268468224;
      54958: inst = 32'd201347790;
      54959: inst = 32'd203423744;
      54960: inst = 32'd471859200;
      54961: inst = 32'd136314880;
      54962: inst = 32'd268468224;
      54963: inst = 32'd201347791;
      54964: inst = 32'd203423744;
      54965: inst = 32'd471859200;
      54966: inst = 32'd136314880;
      54967: inst = 32'd268468224;
      54968: inst = 32'd201347792;
      54969: inst = 32'd203423744;
      54970: inst = 32'd471859200;
      54971: inst = 32'd136314880;
      54972: inst = 32'd268468224;
      54973: inst = 32'd201347793;
      54974: inst = 32'd203423744;
      54975: inst = 32'd471859200;
      54976: inst = 32'd136314880;
      54977: inst = 32'd268468224;
      54978: inst = 32'd201347794;
      54979: inst = 32'd203423744;
      54980: inst = 32'd471859200;
      54981: inst = 32'd136314880;
      54982: inst = 32'd268468224;
      54983: inst = 32'd201347795;
      54984: inst = 32'd203423744;
      54985: inst = 32'd471859200;
      54986: inst = 32'd136314880;
      54987: inst = 32'd268468224;
      54988: inst = 32'd201347796;
      54989: inst = 32'd203423744;
      54990: inst = 32'd471859200;
      54991: inst = 32'd136314880;
      54992: inst = 32'd268468224;
      54993: inst = 32'd201347797;
      54994: inst = 32'd203423744;
      54995: inst = 32'd471859200;
      54996: inst = 32'd136314880;
      54997: inst = 32'd268468224;
      54998: inst = 32'd201347798;
      54999: inst = 32'd203423744;
      55000: inst = 32'd471859200;
      55001: inst = 32'd136314880;
      55002: inst = 32'd268468224;
      55003: inst = 32'd201347799;
      55004: inst = 32'd203423744;
      55005: inst = 32'd471859200;
      55006: inst = 32'd136314880;
      55007: inst = 32'd268468224;
      55008: inst = 32'd201347800;
      55009: inst = 32'd203423744;
      55010: inst = 32'd471859200;
      55011: inst = 32'd136314880;
      55012: inst = 32'd268468224;
      55013: inst = 32'd201347801;
      55014: inst = 32'd203423744;
      55015: inst = 32'd471859200;
      55016: inst = 32'd136314880;
      55017: inst = 32'd268468224;
      55018: inst = 32'd201347802;
      55019: inst = 32'd203423744;
      55020: inst = 32'd471859200;
      55021: inst = 32'd136314880;
      55022: inst = 32'd268468224;
      55023: inst = 32'd201347803;
      55024: inst = 32'd203423744;
      55025: inst = 32'd471859200;
      55026: inst = 32'd136314880;
      55027: inst = 32'd268468224;
      55028: inst = 32'd201347804;
      55029: inst = 32'd203423744;
      55030: inst = 32'd471859200;
      55031: inst = 32'd136314880;
      55032: inst = 32'd268468224;
      55033: inst = 32'd201347805;
      55034: inst = 32'd203423744;
      55035: inst = 32'd471859200;
      55036: inst = 32'd136314880;
      55037: inst = 32'd268468224;
      55038: inst = 32'd201347806;
      55039: inst = 32'd203423744;
      55040: inst = 32'd471859200;
      55041: inst = 32'd136314880;
      55042: inst = 32'd268468224;
      55043: inst = 32'd201347807;
      55044: inst = 32'd203423744;
      55045: inst = 32'd471859200;
      55046: inst = 32'd136314880;
      55047: inst = 32'd268468224;
      55048: inst = 32'd201347808;
      55049: inst = 32'd203423744;
      55050: inst = 32'd471859200;
      55051: inst = 32'd136314880;
      55052: inst = 32'd268468224;
      55053: inst = 32'd201347809;
      55054: inst = 32'd203423744;
      55055: inst = 32'd471859200;
      55056: inst = 32'd136314880;
      55057: inst = 32'd268468224;
      55058: inst = 32'd201347810;
      55059: inst = 32'd203423744;
      55060: inst = 32'd471859200;
      55061: inst = 32'd136314880;
      55062: inst = 32'd268468224;
      55063: inst = 32'd201347811;
      55064: inst = 32'd203423744;
      55065: inst = 32'd471859200;
      55066: inst = 32'd136314880;
      55067: inst = 32'd268468224;
      55068: inst = 32'd201347812;
      55069: inst = 32'd203423744;
      55070: inst = 32'd471859200;
      55071: inst = 32'd136314880;
      55072: inst = 32'd268468224;
      55073: inst = 32'd201347813;
      55074: inst = 32'd203423744;
      55075: inst = 32'd471859200;
      55076: inst = 32'd136314880;
      55077: inst = 32'd268468224;
      55078: inst = 32'd201347814;
      55079: inst = 32'd203423744;
      55080: inst = 32'd471859200;
      55081: inst = 32'd136314880;
      55082: inst = 32'd268468224;
      55083: inst = 32'd201347815;
      55084: inst = 32'd203423744;
      55085: inst = 32'd471859200;
      55086: inst = 32'd136314880;
      55087: inst = 32'd268468224;
      55088: inst = 32'd201347816;
      55089: inst = 32'd203423744;
      55090: inst = 32'd471859200;
      55091: inst = 32'd136314880;
      55092: inst = 32'd268468224;
      55093: inst = 32'd201347817;
      55094: inst = 32'd203423744;
      55095: inst = 32'd471859200;
      55096: inst = 32'd136314880;
      55097: inst = 32'd268468224;
      55098: inst = 32'd201347818;
      55099: inst = 32'd203423744;
      55100: inst = 32'd471859200;
      55101: inst = 32'd136314880;
      55102: inst = 32'd268468224;
      55103: inst = 32'd201347819;
      55104: inst = 32'd203423744;
      55105: inst = 32'd471859200;
      55106: inst = 32'd136314880;
      55107: inst = 32'd268468224;
      55108: inst = 32'd201347820;
      55109: inst = 32'd203423744;
      55110: inst = 32'd471859200;
      55111: inst = 32'd136314880;
      55112: inst = 32'd268468224;
      55113: inst = 32'd201347821;
      55114: inst = 32'd203423744;
      55115: inst = 32'd471859200;
      55116: inst = 32'd136314880;
      55117: inst = 32'd268468224;
      55118: inst = 32'd201347822;
      55119: inst = 32'd203423744;
      55120: inst = 32'd471859200;
      55121: inst = 32'd136314880;
      55122: inst = 32'd268468224;
      55123: inst = 32'd201347823;
      55124: inst = 32'd203423744;
      55125: inst = 32'd471859200;
      55126: inst = 32'd136314880;
      55127: inst = 32'd268468224;
      55128: inst = 32'd201347824;
      55129: inst = 32'd203423744;
      55130: inst = 32'd471859200;
      55131: inst = 32'd136314880;
      55132: inst = 32'd268468224;
      55133: inst = 32'd201347825;
      55134: inst = 32'd203423744;
      55135: inst = 32'd471859200;
      55136: inst = 32'd136314880;
      55137: inst = 32'd268468224;
      55138: inst = 32'd201347826;
      55139: inst = 32'd203423744;
      55140: inst = 32'd471859200;
      55141: inst = 32'd136314880;
      55142: inst = 32'd268468224;
      55143: inst = 32'd201347827;
      55144: inst = 32'd203423744;
      55145: inst = 32'd471859200;
      55146: inst = 32'd136314880;
      55147: inst = 32'd268468224;
      55148: inst = 32'd201347828;
      55149: inst = 32'd203423744;
      55150: inst = 32'd471859200;
      55151: inst = 32'd136314880;
      55152: inst = 32'd268468224;
      55153: inst = 32'd201347829;
      55154: inst = 32'd203423744;
      55155: inst = 32'd471859200;
      55156: inst = 32'd136314880;
      55157: inst = 32'd268468224;
      55158: inst = 32'd201347830;
      55159: inst = 32'd203423744;
      55160: inst = 32'd471859200;
      55161: inst = 32'd136314880;
      55162: inst = 32'd268468224;
      55163: inst = 32'd201347831;
      55164: inst = 32'd203423744;
      55165: inst = 32'd471859200;
      55166: inst = 32'd136314880;
      55167: inst = 32'd268468224;
      55168: inst = 32'd201347832;
      55169: inst = 32'd203423744;
      55170: inst = 32'd471859200;
      55171: inst = 32'd136314880;
      55172: inst = 32'd268468224;
      55173: inst = 32'd201347833;
      55174: inst = 32'd203423744;
      55175: inst = 32'd471859200;
      55176: inst = 32'd136314880;
      55177: inst = 32'd268468224;
      55178: inst = 32'd201347834;
      55179: inst = 32'd203423744;
      55180: inst = 32'd471859200;
      55181: inst = 32'd136314880;
      55182: inst = 32'd268468224;
      55183: inst = 32'd201347835;
      55184: inst = 32'd203423744;
      55185: inst = 32'd471859200;
      55186: inst = 32'd136314880;
      55187: inst = 32'd268468224;
      55188: inst = 32'd201347836;
      55189: inst = 32'd203423744;
      55190: inst = 32'd471859200;
      55191: inst = 32'd136314880;
      55192: inst = 32'd268468224;
      55193: inst = 32'd201347837;
      55194: inst = 32'd203423744;
      55195: inst = 32'd471859200;
      55196: inst = 32'd136314880;
      55197: inst = 32'd268468224;
      55198: inst = 32'd201347838;
      55199: inst = 32'd203423744;
      55200: inst = 32'd471859200;
      55201: inst = 32'd136314880;
      55202: inst = 32'd268468224;
      55203: inst = 32'd201347839;
      55204: inst = 32'd203423744;
      55205: inst = 32'd471859200;
      55206: inst = 32'd136314880;
      55207: inst = 32'd268468224;
      55208: inst = 32'd201347840;
      55209: inst = 32'd203423744;
      55210: inst = 32'd471859200;
      55211: inst = 32'd136314880;
      55212: inst = 32'd268468224;
      55213: inst = 32'd201347841;
      55214: inst = 32'd203423744;
      55215: inst = 32'd471859200;
      55216: inst = 32'd136314880;
      55217: inst = 32'd268468224;
      55218: inst = 32'd201347842;
      55219: inst = 32'd203423744;
      55220: inst = 32'd471859200;
      55221: inst = 32'd136314880;
      55222: inst = 32'd268468224;
      55223: inst = 32'd201347843;
      55224: inst = 32'd203423744;
      55225: inst = 32'd471859200;
      55226: inst = 32'd136314880;
      55227: inst = 32'd268468224;
      55228: inst = 32'd201347844;
      55229: inst = 32'd203423744;
      55230: inst = 32'd471859200;
      55231: inst = 32'd136314880;
      55232: inst = 32'd268468224;
      55233: inst = 32'd201347845;
      55234: inst = 32'd203423744;
      55235: inst = 32'd471859200;
      55236: inst = 32'd136314880;
      55237: inst = 32'd268468224;
      55238: inst = 32'd201347846;
      55239: inst = 32'd203423744;
      55240: inst = 32'd471859200;
      55241: inst = 32'd136314880;
      55242: inst = 32'd268468224;
      55243: inst = 32'd201347847;
      55244: inst = 32'd203423744;
      55245: inst = 32'd471859200;
      55246: inst = 32'd136314880;
      55247: inst = 32'd268468224;
      55248: inst = 32'd201347848;
      55249: inst = 32'd203423744;
      55250: inst = 32'd471859200;
      55251: inst = 32'd136314880;
      55252: inst = 32'd268468224;
      55253: inst = 32'd201347849;
      55254: inst = 32'd203423744;
      55255: inst = 32'd471859200;
      55256: inst = 32'd136314880;
      55257: inst = 32'd268468224;
      55258: inst = 32'd201347850;
      55259: inst = 32'd203423744;
      55260: inst = 32'd471859200;
      55261: inst = 32'd136314880;
      55262: inst = 32'd268468224;
      55263: inst = 32'd201347851;
      55264: inst = 32'd203423744;
      55265: inst = 32'd471859200;
      55266: inst = 32'd136314880;
      55267: inst = 32'd268468224;
      55268: inst = 32'd201347852;
      55269: inst = 32'd203423744;
      55270: inst = 32'd471859200;
      55271: inst = 32'd136314880;
      55272: inst = 32'd268468224;
      55273: inst = 32'd201347853;
      55274: inst = 32'd203423744;
      55275: inst = 32'd471859200;
      55276: inst = 32'd136314880;
      55277: inst = 32'd268468224;
      55278: inst = 32'd201347854;
      55279: inst = 32'd203423744;
      55280: inst = 32'd471859200;
      55281: inst = 32'd136314880;
      55282: inst = 32'd268468224;
      55283: inst = 32'd201347855;
      55284: inst = 32'd203423744;
      55285: inst = 32'd471859200;
      55286: inst = 32'd136314880;
      55287: inst = 32'd268468224;
      55288: inst = 32'd201347856;
      55289: inst = 32'd203423744;
      55290: inst = 32'd471859200;
      55291: inst = 32'd136314880;
      55292: inst = 32'd268468224;
      55293: inst = 32'd201347857;
      55294: inst = 32'd203423744;
      55295: inst = 32'd471859200;
      55296: inst = 32'd136314880;
      55297: inst = 32'd268468224;
      55298: inst = 32'd201347858;
      55299: inst = 32'd203423744;
      55300: inst = 32'd471859200;
      55301: inst = 32'd136314880;
      55302: inst = 32'd268468224;
      55303: inst = 32'd201347859;
      55304: inst = 32'd203423744;
      55305: inst = 32'd471859200;
      55306: inst = 32'd136314880;
      55307: inst = 32'd268468224;
      55308: inst = 32'd201347860;
      55309: inst = 32'd203423744;
      55310: inst = 32'd471859200;
      55311: inst = 32'd136314880;
      55312: inst = 32'd268468224;
      55313: inst = 32'd201347861;
      55314: inst = 32'd203423744;
      55315: inst = 32'd471859200;
      55316: inst = 32'd136314880;
      55317: inst = 32'd268468224;
      55318: inst = 32'd201347862;
      55319: inst = 32'd203423744;
      55320: inst = 32'd471859200;
      55321: inst = 32'd136314880;
      55322: inst = 32'd268468224;
      55323: inst = 32'd201347863;
      55324: inst = 32'd203423744;
      55325: inst = 32'd471859200;
      55326: inst = 32'd136314880;
      55327: inst = 32'd268468224;
      55328: inst = 32'd201347864;
      55329: inst = 32'd203423744;
      55330: inst = 32'd471859200;
      55331: inst = 32'd136314880;
      55332: inst = 32'd268468224;
      55333: inst = 32'd201347865;
      55334: inst = 32'd203423744;
      55335: inst = 32'd471859200;
      55336: inst = 32'd136314880;
      55337: inst = 32'd268468224;
      55338: inst = 32'd201347866;
      55339: inst = 32'd203423744;
      55340: inst = 32'd471859200;
      55341: inst = 32'd136314880;
      55342: inst = 32'd268468224;
      55343: inst = 32'd201347867;
      55344: inst = 32'd203423744;
      55345: inst = 32'd471859200;
      55346: inst = 32'd136314880;
      55347: inst = 32'd268468224;
      55348: inst = 32'd201347868;
      55349: inst = 32'd203423744;
      55350: inst = 32'd471859200;
      55351: inst = 32'd136314880;
      55352: inst = 32'd268468224;
      55353: inst = 32'd201347869;
      55354: inst = 32'd203423744;
      55355: inst = 32'd471859200;
      55356: inst = 32'd136314880;
      55357: inst = 32'd268468224;
      55358: inst = 32'd201347870;
      55359: inst = 32'd203423744;
      55360: inst = 32'd471859200;
      55361: inst = 32'd136314880;
      55362: inst = 32'd268468224;
      55363: inst = 32'd201347871;
      55364: inst = 32'd203423744;
      55365: inst = 32'd471859200;
      55366: inst = 32'd136314880;
      55367: inst = 32'd268468224;
      55368: inst = 32'd201347872;
      55369: inst = 32'd203423744;
      55370: inst = 32'd471859200;
      55371: inst = 32'd136314880;
      55372: inst = 32'd268468224;
      55373: inst = 32'd201347873;
      55374: inst = 32'd203423744;
      55375: inst = 32'd471859200;
      55376: inst = 32'd136314880;
      55377: inst = 32'd268468224;
      55378: inst = 32'd201347874;
      55379: inst = 32'd203423744;
      55380: inst = 32'd471859200;
      55381: inst = 32'd136314880;
      55382: inst = 32'd268468224;
      55383: inst = 32'd201347875;
      55384: inst = 32'd203423744;
      55385: inst = 32'd471859200;
      55386: inst = 32'd136314880;
      55387: inst = 32'd268468224;
      55388: inst = 32'd201347876;
      55389: inst = 32'd203423744;
      55390: inst = 32'd471859200;
      55391: inst = 32'd136314880;
      55392: inst = 32'd268468224;
      55393: inst = 32'd201347877;
      55394: inst = 32'd203423744;
      55395: inst = 32'd471859200;
      55396: inst = 32'd136314880;
      55397: inst = 32'd268468224;
      55398: inst = 32'd201347878;
      55399: inst = 32'd203423744;
      55400: inst = 32'd471859200;
      55401: inst = 32'd136314880;
      55402: inst = 32'd268468224;
      55403: inst = 32'd201347879;
      55404: inst = 32'd203423744;
      55405: inst = 32'd471859200;
      55406: inst = 32'd136314880;
      55407: inst = 32'd268468224;
      55408: inst = 32'd201347880;
      55409: inst = 32'd203423744;
      55410: inst = 32'd471859200;
      55411: inst = 32'd136314880;
      55412: inst = 32'd268468224;
      55413: inst = 32'd201347881;
      55414: inst = 32'd203423744;
      55415: inst = 32'd471859200;
      55416: inst = 32'd136314880;
      55417: inst = 32'd268468224;
      55418: inst = 32'd201347882;
      55419: inst = 32'd203423744;
      55420: inst = 32'd471859200;
      55421: inst = 32'd136314880;
      55422: inst = 32'd268468224;
      55423: inst = 32'd201347883;
      55424: inst = 32'd203423744;
      55425: inst = 32'd471859200;
      55426: inst = 32'd136314880;
      55427: inst = 32'd268468224;
      55428: inst = 32'd201347884;
      55429: inst = 32'd203423744;
      55430: inst = 32'd471859200;
      55431: inst = 32'd136314880;
      55432: inst = 32'd268468224;
      55433: inst = 32'd201347885;
      55434: inst = 32'd203423744;
      55435: inst = 32'd471859200;
      55436: inst = 32'd136314880;
      55437: inst = 32'd268468224;
      55438: inst = 32'd201347886;
      55439: inst = 32'd203423744;
      55440: inst = 32'd471859200;
      55441: inst = 32'd136314880;
      55442: inst = 32'd268468224;
      55443: inst = 32'd201347887;
      55444: inst = 32'd203423744;
      55445: inst = 32'd471859200;
      55446: inst = 32'd136314880;
      55447: inst = 32'd268468224;
      55448: inst = 32'd201347888;
      55449: inst = 32'd203423744;
      55450: inst = 32'd471859200;
      55451: inst = 32'd136314880;
      55452: inst = 32'd268468224;
      55453: inst = 32'd201347889;
      55454: inst = 32'd203423744;
      55455: inst = 32'd471859200;
      55456: inst = 32'd136314880;
      55457: inst = 32'd268468224;
      55458: inst = 32'd201347890;
      55459: inst = 32'd203423744;
      55460: inst = 32'd471859200;
      55461: inst = 32'd136314880;
      55462: inst = 32'd268468224;
      55463: inst = 32'd201347891;
      55464: inst = 32'd203423744;
      55465: inst = 32'd471859200;
      55466: inst = 32'd136314880;
      55467: inst = 32'd268468224;
      55468: inst = 32'd201347892;
      55469: inst = 32'd203423744;
      55470: inst = 32'd471859200;
      55471: inst = 32'd136314880;
      55472: inst = 32'd268468224;
      55473: inst = 32'd201347893;
      55474: inst = 32'd203423744;
      55475: inst = 32'd471859200;
      55476: inst = 32'd136314880;
      55477: inst = 32'd268468224;
      55478: inst = 32'd201347894;
      55479: inst = 32'd203423744;
      55480: inst = 32'd471859200;
      55481: inst = 32'd136314880;
      55482: inst = 32'd268468224;
      55483: inst = 32'd201347895;
      55484: inst = 32'd203423744;
      55485: inst = 32'd471859200;
      55486: inst = 32'd136314880;
      55487: inst = 32'd268468224;
      55488: inst = 32'd201347896;
      55489: inst = 32'd203423744;
      55490: inst = 32'd471859200;
      55491: inst = 32'd136314880;
      55492: inst = 32'd268468224;
      55493: inst = 32'd201347897;
      55494: inst = 32'd203423744;
      55495: inst = 32'd471859200;
      55496: inst = 32'd136314880;
      55497: inst = 32'd268468224;
      55498: inst = 32'd201347898;
      55499: inst = 32'd203423744;
      55500: inst = 32'd471859200;
      55501: inst = 32'd136314880;
      55502: inst = 32'd268468224;
      55503: inst = 32'd201347899;
      55504: inst = 32'd203423744;
      55505: inst = 32'd471859200;
      55506: inst = 32'd136314880;
      55507: inst = 32'd268468224;
      55508: inst = 32'd201347900;
      55509: inst = 32'd203423744;
      55510: inst = 32'd471859200;
      55511: inst = 32'd136314880;
      55512: inst = 32'd268468224;
      55513: inst = 32'd201347901;
      55514: inst = 32'd203423744;
      55515: inst = 32'd471859200;
      55516: inst = 32'd136314880;
      55517: inst = 32'd268468224;
      55518: inst = 32'd201347902;
      55519: inst = 32'd203423744;
      55520: inst = 32'd471859200;
      55521: inst = 32'd136314880;
      55522: inst = 32'd268468224;
      55523: inst = 32'd201347903;
      55524: inst = 32'd203423744;
      55525: inst = 32'd471859200;
      55526: inst = 32'd136314880;
      55527: inst = 32'd268468224;
      55528: inst = 32'd201347904;
      55529: inst = 32'd203423744;
      55530: inst = 32'd471859200;
      55531: inst = 32'd136314880;
      55532: inst = 32'd268468224;
      55533: inst = 32'd201347905;
      55534: inst = 32'd203423744;
      55535: inst = 32'd471859200;
      55536: inst = 32'd136314880;
      55537: inst = 32'd268468224;
      55538: inst = 32'd201347906;
      55539: inst = 32'd203423744;
      55540: inst = 32'd471859200;
      55541: inst = 32'd136314880;
      55542: inst = 32'd268468224;
      55543: inst = 32'd201347907;
      55544: inst = 32'd203423744;
      55545: inst = 32'd471859200;
      55546: inst = 32'd136314880;
      55547: inst = 32'd268468224;
      55548: inst = 32'd201347908;
      55549: inst = 32'd203423744;
      55550: inst = 32'd471859200;
      55551: inst = 32'd136314880;
      55552: inst = 32'd268468224;
      55553: inst = 32'd201347909;
      55554: inst = 32'd203423744;
      55555: inst = 32'd471859200;
      55556: inst = 32'd136314880;
      55557: inst = 32'd268468224;
      55558: inst = 32'd201347910;
      55559: inst = 32'd203423744;
      55560: inst = 32'd471859200;
      55561: inst = 32'd136314880;
      55562: inst = 32'd268468224;
      55563: inst = 32'd201347911;
      55564: inst = 32'd203423744;
      55565: inst = 32'd471859200;
      55566: inst = 32'd136314880;
      55567: inst = 32'd268468224;
      55568: inst = 32'd201347912;
      55569: inst = 32'd203423744;
      55570: inst = 32'd471859200;
      55571: inst = 32'd136314880;
      55572: inst = 32'd268468224;
      55573: inst = 32'd201347913;
      55574: inst = 32'd203423744;
      55575: inst = 32'd471859200;
      55576: inst = 32'd136314880;
      55577: inst = 32'd268468224;
      55578: inst = 32'd201347914;
      55579: inst = 32'd203423744;
      55580: inst = 32'd471859200;
      55581: inst = 32'd136314880;
      55582: inst = 32'd268468224;
      55583: inst = 32'd201347915;
      55584: inst = 32'd203423744;
      55585: inst = 32'd471859200;
      55586: inst = 32'd136314880;
      55587: inst = 32'd268468224;
      55588: inst = 32'd201347916;
      55589: inst = 32'd203423744;
      55590: inst = 32'd471859200;
      55591: inst = 32'd136314880;
      55592: inst = 32'd268468224;
      55593: inst = 32'd201347917;
      55594: inst = 32'd203423744;
      55595: inst = 32'd471859200;
      55596: inst = 32'd136314880;
      55597: inst = 32'd268468224;
      55598: inst = 32'd201347918;
      55599: inst = 32'd203423744;
      55600: inst = 32'd471859200;
      55601: inst = 32'd136314880;
      55602: inst = 32'd268468224;
      55603: inst = 32'd201347919;
      55604: inst = 32'd203423744;
      55605: inst = 32'd471859200;
      55606: inst = 32'd136314880;
      55607: inst = 32'd268468224;
      55608: inst = 32'd201347920;
      55609: inst = 32'd203423744;
      55610: inst = 32'd471859200;
      55611: inst = 32'd136314880;
      55612: inst = 32'd268468224;
      55613: inst = 32'd201347921;
      55614: inst = 32'd203423744;
      55615: inst = 32'd471859200;
      55616: inst = 32'd136314880;
      55617: inst = 32'd268468224;
      55618: inst = 32'd201347922;
      55619: inst = 32'd203423744;
      55620: inst = 32'd471859200;
      55621: inst = 32'd136314880;
      55622: inst = 32'd268468224;
      55623: inst = 32'd201347923;
      55624: inst = 32'd203423744;
      55625: inst = 32'd471859200;
      55626: inst = 32'd136314880;
      55627: inst = 32'd268468224;
      55628: inst = 32'd201347924;
      55629: inst = 32'd203423744;
      55630: inst = 32'd471859200;
      55631: inst = 32'd136314880;
      55632: inst = 32'd268468224;
      55633: inst = 32'd201347925;
      55634: inst = 32'd203423744;
      55635: inst = 32'd471859200;
      55636: inst = 32'd136314880;
      55637: inst = 32'd268468224;
      55638: inst = 32'd201347926;
      55639: inst = 32'd203423744;
      55640: inst = 32'd471859200;
      55641: inst = 32'd136314880;
      55642: inst = 32'd268468224;
      55643: inst = 32'd201347927;
      55644: inst = 32'd203423744;
      55645: inst = 32'd471859200;
      55646: inst = 32'd136314880;
      55647: inst = 32'd268468224;
      55648: inst = 32'd201347928;
      55649: inst = 32'd203423744;
      55650: inst = 32'd471859200;
      55651: inst = 32'd136314880;
      55652: inst = 32'd268468224;
      55653: inst = 32'd201347929;
      55654: inst = 32'd203423744;
      55655: inst = 32'd471859200;
      55656: inst = 32'd136314880;
      55657: inst = 32'd268468224;
      55658: inst = 32'd201347930;
      55659: inst = 32'd203423744;
      55660: inst = 32'd471859200;
      55661: inst = 32'd136314880;
      55662: inst = 32'd268468224;
      55663: inst = 32'd201347931;
      55664: inst = 32'd203423744;
      55665: inst = 32'd471859200;
      55666: inst = 32'd136314880;
      55667: inst = 32'd268468224;
      55668: inst = 32'd201347932;
      55669: inst = 32'd203423744;
      55670: inst = 32'd471859200;
      55671: inst = 32'd136314880;
      55672: inst = 32'd268468224;
      55673: inst = 32'd201347933;
      55674: inst = 32'd203423744;
      55675: inst = 32'd471859200;
      55676: inst = 32'd136314880;
      55677: inst = 32'd268468224;
      55678: inst = 32'd201347934;
      55679: inst = 32'd203423744;
      55680: inst = 32'd471859200;
      55681: inst = 32'd136314880;
      55682: inst = 32'd268468224;
      55683: inst = 32'd201347935;
      55684: inst = 32'd203423744;
      55685: inst = 32'd471859200;
      55686: inst = 32'd136314880;
      55687: inst = 32'd268468224;
      55688: inst = 32'd201347936;
      55689: inst = 32'd203423744;
      55690: inst = 32'd471859200;
      55691: inst = 32'd136314880;
      55692: inst = 32'd268468224;
      55693: inst = 32'd201347937;
      55694: inst = 32'd203423744;
      55695: inst = 32'd471859200;
      55696: inst = 32'd136314880;
      55697: inst = 32'd268468224;
      55698: inst = 32'd201347938;
      55699: inst = 32'd203423744;
      55700: inst = 32'd471859200;
      55701: inst = 32'd136314880;
      55702: inst = 32'd268468224;
      55703: inst = 32'd201347939;
      55704: inst = 32'd203423744;
      55705: inst = 32'd471859200;
      55706: inst = 32'd136314880;
      55707: inst = 32'd268468224;
      55708: inst = 32'd201347940;
      55709: inst = 32'd203423744;
      55710: inst = 32'd471859200;
      55711: inst = 32'd136314880;
      55712: inst = 32'd268468224;
      55713: inst = 32'd201347941;
      55714: inst = 32'd203423744;
      55715: inst = 32'd471859200;
      55716: inst = 32'd136314880;
      55717: inst = 32'd268468224;
      55718: inst = 32'd201347942;
      55719: inst = 32'd203423744;
      55720: inst = 32'd471859200;
      55721: inst = 32'd136314880;
      55722: inst = 32'd268468224;
      55723: inst = 32'd201347943;
      55724: inst = 32'd203423744;
      55725: inst = 32'd471859200;
      55726: inst = 32'd136314880;
      55727: inst = 32'd268468224;
      55728: inst = 32'd201347944;
      55729: inst = 32'd203423744;
      55730: inst = 32'd471859200;
      55731: inst = 32'd136314880;
      55732: inst = 32'd268468224;
      55733: inst = 32'd201347945;
      55734: inst = 32'd203423744;
      55735: inst = 32'd471859200;
      55736: inst = 32'd136314880;
      55737: inst = 32'd268468224;
      55738: inst = 32'd201347946;
      55739: inst = 32'd203423744;
      55740: inst = 32'd471859200;
      55741: inst = 32'd136314880;
      55742: inst = 32'd268468224;
      55743: inst = 32'd201347947;
      55744: inst = 32'd203423744;
      55745: inst = 32'd471859200;
      55746: inst = 32'd136314880;
      55747: inst = 32'd268468224;
      55748: inst = 32'd201347948;
      55749: inst = 32'd203423744;
      55750: inst = 32'd471859200;
      55751: inst = 32'd136314880;
      55752: inst = 32'd268468224;
      55753: inst = 32'd201347949;
      55754: inst = 32'd203423744;
      55755: inst = 32'd471859200;
      55756: inst = 32'd136314880;
      55757: inst = 32'd268468224;
      55758: inst = 32'd201347950;
      55759: inst = 32'd203423744;
      55760: inst = 32'd471859200;
      55761: inst = 32'd136314880;
      55762: inst = 32'd268468224;
      55763: inst = 32'd201347951;
      55764: inst = 32'd203423744;
      55765: inst = 32'd471859200;
      55766: inst = 32'd136314880;
      55767: inst = 32'd268468224;
      55768: inst = 32'd201347952;
      55769: inst = 32'd203423744;
      55770: inst = 32'd471859200;
      55771: inst = 32'd136314880;
      55772: inst = 32'd268468224;
      55773: inst = 32'd201347953;
      55774: inst = 32'd203423744;
      55775: inst = 32'd471859200;
      55776: inst = 32'd136314880;
      55777: inst = 32'd268468224;
      55778: inst = 32'd201347954;
      55779: inst = 32'd203423744;
      55780: inst = 32'd471859200;
      55781: inst = 32'd136314880;
      55782: inst = 32'd268468224;
      55783: inst = 32'd201347955;
      55784: inst = 32'd203423744;
      55785: inst = 32'd471859200;
      55786: inst = 32'd136314880;
      55787: inst = 32'd268468224;
      55788: inst = 32'd201347956;
      55789: inst = 32'd203423744;
      55790: inst = 32'd471859200;
      55791: inst = 32'd136314880;
      55792: inst = 32'd268468224;
      55793: inst = 32'd201347957;
      55794: inst = 32'd203423744;
      55795: inst = 32'd471859200;
      55796: inst = 32'd136314880;
      55797: inst = 32'd268468224;
      55798: inst = 32'd201347958;
      55799: inst = 32'd203423744;
      55800: inst = 32'd471859200;
      55801: inst = 32'd136314880;
      55802: inst = 32'd268468224;
      55803: inst = 32'd201347959;
      55804: inst = 32'd203423744;
      55805: inst = 32'd471859200;
      55806: inst = 32'd136314880;
      55807: inst = 32'd268468224;
      55808: inst = 32'd201347960;
      55809: inst = 32'd203423744;
      55810: inst = 32'd471859200;
      55811: inst = 32'd136314880;
      55812: inst = 32'd268468224;
      55813: inst = 32'd201347961;
      55814: inst = 32'd203423744;
      55815: inst = 32'd471859200;
      55816: inst = 32'd136314880;
      55817: inst = 32'd268468224;
      55818: inst = 32'd201347962;
      55819: inst = 32'd203423744;
      55820: inst = 32'd471859200;
      55821: inst = 32'd136314880;
      55822: inst = 32'd268468224;
      55823: inst = 32'd201347963;
      55824: inst = 32'd203423744;
      55825: inst = 32'd471859200;
      55826: inst = 32'd136314880;
      55827: inst = 32'd268468224;
      55828: inst = 32'd201347964;
      55829: inst = 32'd203423744;
      55830: inst = 32'd471859200;
      55831: inst = 32'd136314880;
      55832: inst = 32'd268468224;
      55833: inst = 32'd201347965;
      55834: inst = 32'd203423744;
      55835: inst = 32'd471859200;
      55836: inst = 32'd136314880;
      55837: inst = 32'd268468224;
      55838: inst = 32'd201347966;
      55839: inst = 32'd203423744;
      55840: inst = 32'd471859200;
      55841: inst = 32'd136314880;
      55842: inst = 32'd268468224;
      55843: inst = 32'd201347967;
      55844: inst = 32'd203423744;
      55845: inst = 32'd471859200;
      55846: inst = 32'd136314880;
      55847: inst = 32'd268468224;
      55848: inst = 32'd201347968;
      55849: inst = 32'd203423744;
      55850: inst = 32'd471859200;
      55851: inst = 32'd136314880;
      55852: inst = 32'd268468224;
      55853: inst = 32'd201347969;
      55854: inst = 32'd203423744;
      55855: inst = 32'd471859200;
      55856: inst = 32'd136314880;
      55857: inst = 32'd268468224;
      55858: inst = 32'd201347970;
      55859: inst = 32'd203423744;
      55860: inst = 32'd471859200;
      55861: inst = 32'd136314880;
      55862: inst = 32'd268468224;
      55863: inst = 32'd201347971;
      55864: inst = 32'd203423744;
      55865: inst = 32'd471859200;
      55866: inst = 32'd136314880;
      55867: inst = 32'd268468224;
      55868: inst = 32'd201347972;
      55869: inst = 32'd203423744;
      55870: inst = 32'd471859200;
      55871: inst = 32'd136314880;
      55872: inst = 32'd268468224;
      55873: inst = 32'd201347973;
      55874: inst = 32'd203423744;
      55875: inst = 32'd471859200;
      55876: inst = 32'd136314880;
      55877: inst = 32'd268468224;
      55878: inst = 32'd201347974;
      55879: inst = 32'd203423744;
      55880: inst = 32'd471859200;
      55881: inst = 32'd136314880;
      55882: inst = 32'd268468224;
      55883: inst = 32'd201347975;
      55884: inst = 32'd203423744;
      55885: inst = 32'd471859200;
      55886: inst = 32'd136314880;
      55887: inst = 32'd268468224;
      55888: inst = 32'd201347976;
      55889: inst = 32'd203423744;
      55890: inst = 32'd471859200;
      55891: inst = 32'd136314880;
      55892: inst = 32'd268468224;
      55893: inst = 32'd201347977;
      55894: inst = 32'd203423744;
      55895: inst = 32'd471859200;
      55896: inst = 32'd136314880;
      55897: inst = 32'd268468224;
      55898: inst = 32'd201347978;
      55899: inst = 32'd203423744;
      55900: inst = 32'd471859200;
      55901: inst = 32'd136314880;
      55902: inst = 32'd268468224;
      55903: inst = 32'd201347979;
      55904: inst = 32'd203423744;
      55905: inst = 32'd471859200;
      55906: inst = 32'd136314880;
      55907: inst = 32'd268468224;
      55908: inst = 32'd201347980;
      55909: inst = 32'd203423744;
      55910: inst = 32'd471859200;
      55911: inst = 32'd136314880;
      55912: inst = 32'd268468224;
      55913: inst = 32'd201347981;
      55914: inst = 32'd203423744;
      55915: inst = 32'd471859200;
      55916: inst = 32'd136314880;
      55917: inst = 32'd268468224;
      55918: inst = 32'd201347982;
      55919: inst = 32'd203423744;
      55920: inst = 32'd471859200;
      55921: inst = 32'd136314880;
      55922: inst = 32'd268468224;
      55923: inst = 32'd201347983;
      55924: inst = 32'd203423744;
      55925: inst = 32'd471859200;
      55926: inst = 32'd136314880;
      55927: inst = 32'd268468224;
      55928: inst = 32'd201347984;
      55929: inst = 32'd203423744;
      55930: inst = 32'd471859200;
      55931: inst = 32'd136314880;
      55932: inst = 32'd268468224;
      55933: inst = 32'd201347985;
      55934: inst = 32'd203423744;
      55935: inst = 32'd471859200;
      55936: inst = 32'd136314880;
      55937: inst = 32'd268468224;
      55938: inst = 32'd201347986;
      55939: inst = 32'd203423744;
      55940: inst = 32'd471859200;
      55941: inst = 32'd136314880;
      55942: inst = 32'd268468224;
      55943: inst = 32'd201347987;
      55944: inst = 32'd203423744;
      55945: inst = 32'd471859200;
      55946: inst = 32'd136314880;
      55947: inst = 32'd268468224;
      55948: inst = 32'd201347988;
      55949: inst = 32'd203423744;
      55950: inst = 32'd471859200;
      55951: inst = 32'd136314880;
      55952: inst = 32'd268468224;
      55953: inst = 32'd201347989;
      55954: inst = 32'd203423744;
      55955: inst = 32'd471859200;
      55956: inst = 32'd136314880;
      55957: inst = 32'd268468224;
      55958: inst = 32'd201347990;
      55959: inst = 32'd203423744;
      55960: inst = 32'd471859200;
      55961: inst = 32'd136314880;
      55962: inst = 32'd268468224;
      55963: inst = 32'd201347991;
      55964: inst = 32'd203423744;
      55965: inst = 32'd471859200;
      55966: inst = 32'd136314880;
      55967: inst = 32'd268468224;
      55968: inst = 32'd201347992;
      55969: inst = 32'd203423744;
      55970: inst = 32'd471859200;
      55971: inst = 32'd136314880;
      55972: inst = 32'd268468224;
      55973: inst = 32'd201347993;
      55974: inst = 32'd203423744;
      55975: inst = 32'd471859200;
      55976: inst = 32'd136314880;
      55977: inst = 32'd268468224;
      55978: inst = 32'd201347994;
      55979: inst = 32'd203423744;
      55980: inst = 32'd471859200;
      55981: inst = 32'd136314880;
      55982: inst = 32'd268468224;
      55983: inst = 32'd201347995;
      55984: inst = 32'd203423744;
      55985: inst = 32'd471859200;
      55986: inst = 32'd136314880;
      55987: inst = 32'd268468224;
      55988: inst = 32'd201347996;
      55989: inst = 32'd203423744;
      55990: inst = 32'd471859200;
      55991: inst = 32'd136314880;
      55992: inst = 32'd268468224;
      55993: inst = 32'd201347997;
      55994: inst = 32'd203423744;
      55995: inst = 32'd471859200;
      55996: inst = 32'd136314880;
      55997: inst = 32'd268468224;
      55998: inst = 32'd201347998;
      55999: inst = 32'd203423744;
      56000: inst = 32'd471859200;
      56001: inst = 32'd136314880;
      56002: inst = 32'd268468224;
      56003: inst = 32'd201347999;
      56004: inst = 32'd203423744;
      56005: inst = 32'd471859200;
      56006: inst = 32'd136314880;
      56007: inst = 32'd268468224;
      56008: inst = 32'd201348000;
      56009: inst = 32'd203423744;
      56010: inst = 32'd471859200;
      56011: inst = 32'd136314880;
      56012: inst = 32'd268468224;
      56013: inst = 32'd201348001;
      56014: inst = 32'd203423744;
      56015: inst = 32'd471859200;
      56016: inst = 32'd136314880;
      56017: inst = 32'd268468224;
      56018: inst = 32'd201348002;
      56019: inst = 32'd203423744;
      56020: inst = 32'd471859200;
      56021: inst = 32'd136314880;
      56022: inst = 32'd268468224;
      56023: inst = 32'd201348003;
      56024: inst = 32'd203423744;
      56025: inst = 32'd471859200;
      56026: inst = 32'd136314880;
      56027: inst = 32'd268468224;
      56028: inst = 32'd201348004;
      56029: inst = 32'd203423744;
      56030: inst = 32'd471859200;
      56031: inst = 32'd136314880;
      56032: inst = 32'd268468224;
      56033: inst = 32'd201348005;
      56034: inst = 32'd203423744;
      56035: inst = 32'd471859200;
      56036: inst = 32'd136314880;
      56037: inst = 32'd268468224;
      56038: inst = 32'd201348006;
      56039: inst = 32'd203423744;
      56040: inst = 32'd471859200;
      56041: inst = 32'd136314880;
      56042: inst = 32'd268468224;
      56043: inst = 32'd201348007;
      56044: inst = 32'd203423744;
      56045: inst = 32'd471859200;
      56046: inst = 32'd136314880;
      56047: inst = 32'd268468224;
      56048: inst = 32'd201348008;
      56049: inst = 32'd203423744;
      56050: inst = 32'd471859200;
      56051: inst = 32'd136314880;
      56052: inst = 32'd268468224;
      56053: inst = 32'd201348009;
      56054: inst = 32'd203423744;
      56055: inst = 32'd471859200;
      56056: inst = 32'd136314880;
      56057: inst = 32'd268468224;
      56058: inst = 32'd201348010;
      56059: inst = 32'd203423744;
      56060: inst = 32'd471859200;
      56061: inst = 32'd136314880;
      56062: inst = 32'd268468224;
      56063: inst = 32'd201348011;
      56064: inst = 32'd203423744;
      56065: inst = 32'd471859200;
      56066: inst = 32'd136314880;
      56067: inst = 32'd268468224;
      56068: inst = 32'd201348012;
      56069: inst = 32'd203423744;
      56070: inst = 32'd471859200;
      56071: inst = 32'd136314880;
      56072: inst = 32'd268468224;
      56073: inst = 32'd201348013;
      56074: inst = 32'd203423744;
      56075: inst = 32'd471859200;
      56076: inst = 32'd136314880;
      56077: inst = 32'd268468224;
      56078: inst = 32'd201348014;
      56079: inst = 32'd203423744;
      56080: inst = 32'd471859200;
      56081: inst = 32'd136314880;
      56082: inst = 32'd268468224;
      56083: inst = 32'd201348015;
      56084: inst = 32'd203423744;
      56085: inst = 32'd471859200;
      56086: inst = 32'd136314880;
      56087: inst = 32'd268468224;
      56088: inst = 32'd201348016;
      56089: inst = 32'd203423744;
      56090: inst = 32'd471859200;
      56091: inst = 32'd136314880;
      56092: inst = 32'd268468224;
      56093: inst = 32'd201348017;
      56094: inst = 32'd203423744;
      56095: inst = 32'd471859200;
      56096: inst = 32'd136314880;
      56097: inst = 32'd268468224;
      56098: inst = 32'd201348018;
      56099: inst = 32'd203423744;
      56100: inst = 32'd471859200;
      56101: inst = 32'd136314880;
      56102: inst = 32'd268468224;
      56103: inst = 32'd201348019;
      56104: inst = 32'd203423744;
      56105: inst = 32'd471859200;
      56106: inst = 32'd136314880;
      56107: inst = 32'd268468224;
      56108: inst = 32'd201348020;
      56109: inst = 32'd203423744;
      56110: inst = 32'd471859200;
      56111: inst = 32'd136314880;
      56112: inst = 32'd268468224;
      56113: inst = 32'd201348021;
      56114: inst = 32'd203423744;
      56115: inst = 32'd471859200;
      56116: inst = 32'd136314880;
      56117: inst = 32'd268468224;
      56118: inst = 32'd201348022;
      56119: inst = 32'd203423744;
      56120: inst = 32'd471859200;
      56121: inst = 32'd136314880;
      56122: inst = 32'd268468224;
      56123: inst = 32'd201348023;
      56124: inst = 32'd203423744;
      56125: inst = 32'd471859200;
      56126: inst = 32'd136314880;
      56127: inst = 32'd268468224;
      56128: inst = 32'd201348024;
      56129: inst = 32'd203423744;
      56130: inst = 32'd471859200;
      56131: inst = 32'd136314880;
      56132: inst = 32'd268468224;
      56133: inst = 32'd201348025;
      56134: inst = 32'd203423744;
      56135: inst = 32'd471859200;
      56136: inst = 32'd136314880;
      56137: inst = 32'd268468224;
      56138: inst = 32'd201348026;
      56139: inst = 32'd203423744;
      56140: inst = 32'd471859200;
      56141: inst = 32'd136314880;
      56142: inst = 32'd268468224;
      56143: inst = 32'd201348027;
      56144: inst = 32'd203423744;
      56145: inst = 32'd471859200;
      56146: inst = 32'd136314880;
      56147: inst = 32'd268468224;
      56148: inst = 32'd201348028;
      56149: inst = 32'd203423744;
      56150: inst = 32'd471859200;
      56151: inst = 32'd136314880;
      56152: inst = 32'd268468224;
      56153: inst = 32'd201348029;
      56154: inst = 32'd203423744;
      56155: inst = 32'd471859200;
      56156: inst = 32'd136314880;
      56157: inst = 32'd268468224;
      56158: inst = 32'd201348030;
      56159: inst = 32'd203423744;
      56160: inst = 32'd471859200;
      56161: inst = 32'd136314880;
      56162: inst = 32'd268468224;
      56163: inst = 32'd201348031;
      56164: inst = 32'd203423744;
      56165: inst = 32'd471859200;
      56166: inst = 32'd136314880;
      56167: inst = 32'd268468224;
      56168: inst = 32'd201348032;
      56169: inst = 32'd203423744;
      56170: inst = 32'd471859200;
      56171: inst = 32'd136314880;
      56172: inst = 32'd268468224;
      56173: inst = 32'd201348033;
      56174: inst = 32'd203423744;
      56175: inst = 32'd471859200;
      56176: inst = 32'd136314880;
      56177: inst = 32'd268468224;
      56178: inst = 32'd201348034;
      56179: inst = 32'd203423744;
      56180: inst = 32'd471859200;
      56181: inst = 32'd136314880;
      56182: inst = 32'd268468224;
      56183: inst = 32'd201348035;
      56184: inst = 32'd203423744;
      56185: inst = 32'd471859200;
      56186: inst = 32'd136314880;
      56187: inst = 32'd268468224;
      56188: inst = 32'd201348036;
      56189: inst = 32'd203423744;
      56190: inst = 32'd471859200;
      56191: inst = 32'd136314880;
      56192: inst = 32'd268468224;
      56193: inst = 32'd201348037;
      56194: inst = 32'd203423744;
      56195: inst = 32'd471859200;
      56196: inst = 32'd136314880;
      56197: inst = 32'd268468224;
      56198: inst = 32'd201348038;
      56199: inst = 32'd203423744;
      56200: inst = 32'd471859200;
      56201: inst = 32'd136314880;
      56202: inst = 32'd268468224;
      56203: inst = 32'd201348039;
      56204: inst = 32'd203423744;
      56205: inst = 32'd471859200;
      56206: inst = 32'd136314880;
      56207: inst = 32'd268468224;
      56208: inst = 32'd201348040;
      56209: inst = 32'd203423744;
      56210: inst = 32'd471859200;
      56211: inst = 32'd136314880;
      56212: inst = 32'd268468224;
      56213: inst = 32'd201348041;
      56214: inst = 32'd203423744;
      56215: inst = 32'd471859200;
      56216: inst = 32'd136314880;
      56217: inst = 32'd268468224;
      56218: inst = 32'd201348042;
      56219: inst = 32'd203423744;
      56220: inst = 32'd471859200;
      56221: inst = 32'd136314880;
      56222: inst = 32'd268468224;
      56223: inst = 32'd201348043;
      56224: inst = 32'd203423744;
      56225: inst = 32'd471859200;
      56226: inst = 32'd136314880;
      56227: inst = 32'd268468224;
      56228: inst = 32'd201348044;
      56229: inst = 32'd203423744;
      56230: inst = 32'd471859200;
      56231: inst = 32'd136314880;
      56232: inst = 32'd268468224;
      56233: inst = 32'd201348045;
      56234: inst = 32'd203423744;
      56235: inst = 32'd471859200;
      56236: inst = 32'd136314880;
      56237: inst = 32'd268468224;
      56238: inst = 32'd201348046;
      56239: inst = 32'd203423744;
      56240: inst = 32'd471859200;
      56241: inst = 32'd136314880;
      56242: inst = 32'd268468224;
      56243: inst = 32'd201348047;
      56244: inst = 32'd203423744;
      56245: inst = 32'd471859200;
      56246: inst = 32'd136314880;
      56247: inst = 32'd268468224;
      56248: inst = 32'd201348048;
      56249: inst = 32'd203423744;
      56250: inst = 32'd471859200;
      56251: inst = 32'd136314880;
      56252: inst = 32'd268468224;
      56253: inst = 32'd201348049;
      56254: inst = 32'd203423744;
      56255: inst = 32'd471859200;
      56256: inst = 32'd136314880;
      56257: inst = 32'd268468224;
      56258: inst = 32'd201348050;
      56259: inst = 32'd203423744;
      56260: inst = 32'd471859200;
      56261: inst = 32'd136314880;
      56262: inst = 32'd268468224;
      56263: inst = 32'd201348051;
      56264: inst = 32'd203423744;
      56265: inst = 32'd471859200;
      56266: inst = 32'd136314880;
      56267: inst = 32'd268468224;
      56268: inst = 32'd201348052;
      56269: inst = 32'd203423744;
      56270: inst = 32'd471859200;
      56271: inst = 32'd136314880;
      56272: inst = 32'd268468224;
      56273: inst = 32'd201348053;
      56274: inst = 32'd203423744;
      56275: inst = 32'd471859200;
      56276: inst = 32'd136314880;
      56277: inst = 32'd268468224;
      56278: inst = 32'd201348054;
      56279: inst = 32'd203423744;
      56280: inst = 32'd471859200;
      56281: inst = 32'd136314880;
      56282: inst = 32'd268468224;
      56283: inst = 32'd201348055;
      56284: inst = 32'd203423744;
      56285: inst = 32'd471859200;
      56286: inst = 32'd136314880;
      56287: inst = 32'd268468224;
      56288: inst = 32'd201348056;
      56289: inst = 32'd203423744;
      56290: inst = 32'd471859200;
      56291: inst = 32'd136314880;
      56292: inst = 32'd268468224;
      56293: inst = 32'd201348057;
      56294: inst = 32'd203423744;
      56295: inst = 32'd471859200;
      56296: inst = 32'd136314880;
      56297: inst = 32'd268468224;
      56298: inst = 32'd201348058;
      56299: inst = 32'd203423744;
      56300: inst = 32'd471859200;
      56301: inst = 32'd136314880;
      56302: inst = 32'd268468224;
      56303: inst = 32'd201348059;
      56304: inst = 32'd203423744;
      56305: inst = 32'd471859200;
      56306: inst = 32'd136314880;
      56307: inst = 32'd268468224;
      56308: inst = 32'd201348060;
      56309: inst = 32'd203423744;
      56310: inst = 32'd471859200;
      56311: inst = 32'd136314880;
      56312: inst = 32'd268468224;
      56313: inst = 32'd201348061;
      56314: inst = 32'd203423744;
      56315: inst = 32'd471859200;
      56316: inst = 32'd136314880;
      56317: inst = 32'd268468224;
      56318: inst = 32'd201348062;
      56319: inst = 32'd203423744;
      56320: inst = 32'd471859200;
      56321: inst = 32'd136314880;
      56322: inst = 32'd268468224;
      56323: inst = 32'd201348063;
      56324: inst = 32'd203423744;
      56325: inst = 32'd471859200;
      56326: inst = 32'd136314880;
      56327: inst = 32'd268468224;
      56328: inst = 32'd201348064;
      56329: inst = 32'd203423744;
      56330: inst = 32'd471859200;
      56331: inst = 32'd136314880;
      56332: inst = 32'd268468224;
      56333: inst = 32'd201348065;
      56334: inst = 32'd203423744;
      56335: inst = 32'd471859200;
      56336: inst = 32'd136314880;
      56337: inst = 32'd268468224;
      56338: inst = 32'd201348066;
      56339: inst = 32'd203423744;
      56340: inst = 32'd471859200;
      56341: inst = 32'd136314880;
      56342: inst = 32'd268468224;
      56343: inst = 32'd201348067;
      56344: inst = 32'd203423744;
      56345: inst = 32'd471859200;
      56346: inst = 32'd136314880;
      56347: inst = 32'd268468224;
      56348: inst = 32'd201348068;
      56349: inst = 32'd203423744;
      56350: inst = 32'd471859200;
      56351: inst = 32'd136314880;
      56352: inst = 32'd268468224;
      56353: inst = 32'd201348069;
      56354: inst = 32'd203423744;
      56355: inst = 32'd471859200;
      56356: inst = 32'd136314880;
      56357: inst = 32'd268468224;
      56358: inst = 32'd201348070;
      56359: inst = 32'd203423744;
      56360: inst = 32'd471859200;
      56361: inst = 32'd136314880;
      56362: inst = 32'd268468224;
      56363: inst = 32'd201348071;
      56364: inst = 32'd203423744;
      56365: inst = 32'd471859200;
      56366: inst = 32'd136314880;
      56367: inst = 32'd268468224;
      56368: inst = 32'd201348072;
      56369: inst = 32'd203423744;
      56370: inst = 32'd471859200;
      56371: inst = 32'd136314880;
      56372: inst = 32'd268468224;
      56373: inst = 32'd201348073;
      56374: inst = 32'd203423744;
      56375: inst = 32'd471859200;
      56376: inst = 32'd136314880;
      56377: inst = 32'd268468224;
      56378: inst = 32'd201348074;
      56379: inst = 32'd203423744;
      56380: inst = 32'd471859200;
      56381: inst = 32'd136314880;
      56382: inst = 32'd268468224;
      56383: inst = 32'd201348075;
      56384: inst = 32'd203423744;
      56385: inst = 32'd471859200;
      56386: inst = 32'd136314880;
      56387: inst = 32'd268468224;
      56388: inst = 32'd201348076;
      56389: inst = 32'd203423744;
      56390: inst = 32'd471859200;
      56391: inst = 32'd136314880;
      56392: inst = 32'd268468224;
      56393: inst = 32'd201348077;
      56394: inst = 32'd203423744;
      56395: inst = 32'd471859200;
      56396: inst = 32'd136314880;
      56397: inst = 32'd268468224;
      56398: inst = 32'd201348078;
      56399: inst = 32'd203423744;
      56400: inst = 32'd471859200;
      56401: inst = 32'd136314880;
      56402: inst = 32'd268468224;
      56403: inst = 32'd201348079;
      56404: inst = 32'd203423744;
      56405: inst = 32'd471859200;
      56406: inst = 32'd136314880;
      56407: inst = 32'd268468224;
      56408: inst = 32'd201348080;
      56409: inst = 32'd203423744;
      56410: inst = 32'd471859200;
      56411: inst = 32'd136314880;
      56412: inst = 32'd268468224;
      56413: inst = 32'd201348081;
      56414: inst = 32'd203423744;
      56415: inst = 32'd471859200;
      56416: inst = 32'd136314880;
      56417: inst = 32'd268468224;
      56418: inst = 32'd201348082;
      56419: inst = 32'd203423744;
      56420: inst = 32'd471859200;
      56421: inst = 32'd136314880;
      56422: inst = 32'd268468224;
      56423: inst = 32'd201348083;
      56424: inst = 32'd203423744;
      56425: inst = 32'd471859200;
      56426: inst = 32'd136314880;
      56427: inst = 32'd268468224;
      56428: inst = 32'd201348084;
      56429: inst = 32'd203423744;
      56430: inst = 32'd471859200;
      56431: inst = 32'd136314880;
      56432: inst = 32'd268468224;
      56433: inst = 32'd201348085;
      56434: inst = 32'd203423744;
      56435: inst = 32'd471859200;
      56436: inst = 32'd136314880;
      56437: inst = 32'd268468224;
      56438: inst = 32'd201348086;
      56439: inst = 32'd203423744;
      56440: inst = 32'd471859200;
      56441: inst = 32'd136314880;
      56442: inst = 32'd268468224;
      56443: inst = 32'd201348087;
      56444: inst = 32'd203423744;
      56445: inst = 32'd471859200;
      56446: inst = 32'd136314880;
      56447: inst = 32'd268468224;
      56448: inst = 32'd201348088;
      56449: inst = 32'd203423744;
      56450: inst = 32'd471859200;
      56451: inst = 32'd136314880;
      56452: inst = 32'd268468224;
      56453: inst = 32'd201348089;
      56454: inst = 32'd203423744;
      56455: inst = 32'd471859200;
      56456: inst = 32'd136314880;
      56457: inst = 32'd268468224;
      56458: inst = 32'd201348090;
      56459: inst = 32'd203423744;
      56460: inst = 32'd471859200;
      56461: inst = 32'd136314880;
      56462: inst = 32'd268468224;
      56463: inst = 32'd201348091;
      56464: inst = 32'd203423744;
      56465: inst = 32'd471859200;
      56466: inst = 32'd136314880;
      56467: inst = 32'd268468224;
      56468: inst = 32'd201348092;
      56469: inst = 32'd203423744;
      56470: inst = 32'd471859200;
      56471: inst = 32'd136314880;
      56472: inst = 32'd268468224;
      56473: inst = 32'd201348093;
      56474: inst = 32'd203423744;
      56475: inst = 32'd471859200;
      56476: inst = 32'd136314880;
      56477: inst = 32'd268468224;
      56478: inst = 32'd201348094;
      56479: inst = 32'd203423744;
      56480: inst = 32'd471859200;
      56481: inst = 32'd136314880;
      56482: inst = 32'd268468224;
      56483: inst = 32'd201348095;
      56484: inst = 32'd203423744;
      56485: inst = 32'd471859200;
      56486: inst = 32'd136314880;
      56487: inst = 32'd268468224;
      56488: inst = 32'd201348096;
      56489: inst = 32'd203423744;
      56490: inst = 32'd471859200;
      56491: inst = 32'd136314880;
      56492: inst = 32'd268468224;
      56493: inst = 32'd201348097;
      56494: inst = 32'd203423744;
      56495: inst = 32'd471859200;
      56496: inst = 32'd136314880;
      56497: inst = 32'd268468224;
      56498: inst = 32'd201348098;
      56499: inst = 32'd203423744;
      56500: inst = 32'd471859200;
      56501: inst = 32'd136314880;
      56502: inst = 32'd268468224;
      56503: inst = 32'd201348099;
      56504: inst = 32'd203423744;
      56505: inst = 32'd471859200;
      56506: inst = 32'd136314880;
      56507: inst = 32'd268468224;
      56508: inst = 32'd201348100;
      56509: inst = 32'd203423744;
      56510: inst = 32'd471859200;
      56511: inst = 32'd136314880;
      56512: inst = 32'd268468224;
      56513: inst = 32'd201348101;
      56514: inst = 32'd203423744;
      56515: inst = 32'd471859200;
      56516: inst = 32'd136314880;
      56517: inst = 32'd268468224;
      56518: inst = 32'd201348102;
      56519: inst = 32'd203423744;
      56520: inst = 32'd471859200;
      56521: inst = 32'd136314880;
      56522: inst = 32'd268468224;
      56523: inst = 32'd201348103;
      56524: inst = 32'd203423744;
      56525: inst = 32'd471859200;
      56526: inst = 32'd136314880;
      56527: inst = 32'd268468224;
      56528: inst = 32'd201348104;
      56529: inst = 32'd203423744;
      56530: inst = 32'd471859200;
      56531: inst = 32'd136314880;
      56532: inst = 32'd268468224;
      56533: inst = 32'd201348105;
      56534: inst = 32'd203423744;
      56535: inst = 32'd471859200;
      56536: inst = 32'd136314880;
      56537: inst = 32'd268468224;
      56538: inst = 32'd201348106;
      56539: inst = 32'd203423744;
      56540: inst = 32'd471859200;
      56541: inst = 32'd136314880;
      56542: inst = 32'd268468224;
      56543: inst = 32'd201348107;
      56544: inst = 32'd203423744;
      56545: inst = 32'd471859200;
      56546: inst = 32'd136314880;
      56547: inst = 32'd268468224;
      56548: inst = 32'd201348108;
      56549: inst = 32'd203423744;
      56550: inst = 32'd471859200;
      56551: inst = 32'd136314880;
      56552: inst = 32'd268468224;
      56553: inst = 32'd201348109;
      56554: inst = 32'd203423744;
      56555: inst = 32'd471859200;
      56556: inst = 32'd136314880;
      56557: inst = 32'd268468224;
      56558: inst = 32'd201348110;
      56559: inst = 32'd203423744;
      56560: inst = 32'd471859200;
      56561: inst = 32'd136314880;
      56562: inst = 32'd268468224;
      56563: inst = 32'd201348111;
      56564: inst = 32'd203423744;
      56565: inst = 32'd471859200;
      56566: inst = 32'd136314880;
      56567: inst = 32'd268468224;
      56568: inst = 32'd201348112;
      56569: inst = 32'd203423744;
      56570: inst = 32'd471859200;
      56571: inst = 32'd136314880;
      56572: inst = 32'd268468224;
      56573: inst = 32'd201348113;
      56574: inst = 32'd203423744;
      56575: inst = 32'd471859200;
      56576: inst = 32'd136314880;
      56577: inst = 32'd268468224;
      56578: inst = 32'd201348114;
      56579: inst = 32'd203423744;
      56580: inst = 32'd471859200;
      56581: inst = 32'd136314880;
      56582: inst = 32'd268468224;
      56583: inst = 32'd201348115;
      56584: inst = 32'd203423744;
      56585: inst = 32'd471859200;
      56586: inst = 32'd136314880;
      56587: inst = 32'd268468224;
      56588: inst = 32'd201348116;
      56589: inst = 32'd203423744;
      56590: inst = 32'd471859200;
      56591: inst = 32'd136314880;
      56592: inst = 32'd268468224;
      56593: inst = 32'd201348117;
      56594: inst = 32'd203423744;
      56595: inst = 32'd471859200;
      56596: inst = 32'd136314880;
      56597: inst = 32'd268468224;
      56598: inst = 32'd201348118;
      56599: inst = 32'd203423744;
      56600: inst = 32'd471859200;
      56601: inst = 32'd136314880;
      56602: inst = 32'd268468224;
      56603: inst = 32'd201348119;
      56604: inst = 32'd203423744;
      56605: inst = 32'd471859200;
      56606: inst = 32'd136314880;
      56607: inst = 32'd268468224;
      56608: inst = 32'd201348120;
      56609: inst = 32'd203423744;
      56610: inst = 32'd471859200;
      56611: inst = 32'd136314880;
      56612: inst = 32'd268468224;
      56613: inst = 32'd201348121;
      56614: inst = 32'd203423744;
      56615: inst = 32'd471859200;
      56616: inst = 32'd136314880;
      56617: inst = 32'd268468224;
      56618: inst = 32'd201348122;
      56619: inst = 32'd203423744;
      56620: inst = 32'd471859200;
      56621: inst = 32'd136314880;
      56622: inst = 32'd268468224;
      56623: inst = 32'd201348123;
      56624: inst = 32'd203423744;
      56625: inst = 32'd471859200;
      56626: inst = 32'd136314880;
      56627: inst = 32'd268468224;
      56628: inst = 32'd201348124;
      56629: inst = 32'd203423744;
      56630: inst = 32'd471859200;
      56631: inst = 32'd136314880;
      56632: inst = 32'd268468224;
      56633: inst = 32'd201348125;
      56634: inst = 32'd203423744;
      56635: inst = 32'd471859200;
      56636: inst = 32'd136314880;
      56637: inst = 32'd268468224;
      56638: inst = 32'd201348126;
      56639: inst = 32'd203423744;
      56640: inst = 32'd471859200;
      56641: inst = 32'd136314880;
      56642: inst = 32'd268468224;
      56643: inst = 32'd201348127;
      56644: inst = 32'd203423744;
      56645: inst = 32'd471859200;
      56646: inst = 32'd136314880;
      56647: inst = 32'd268468224;
      56648: inst = 32'd201348128;
      56649: inst = 32'd203423744;
      56650: inst = 32'd471859200;
      56651: inst = 32'd136314880;
      56652: inst = 32'd268468224;
      56653: inst = 32'd201348129;
      56654: inst = 32'd203423744;
      56655: inst = 32'd471859200;
      56656: inst = 32'd136314880;
      56657: inst = 32'd268468224;
      56658: inst = 32'd201348130;
      56659: inst = 32'd203423744;
      56660: inst = 32'd471859200;
      56661: inst = 32'd136314880;
      56662: inst = 32'd268468224;
      56663: inst = 32'd201348131;
      56664: inst = 32'd203423744;
      56665: inst = 32'd471859200;
      56666: inst = 32'd136314880;
      56667: inst = 32'd268468224;
      56668: inst = 32'd201348132;
      56669: inst = 32'd203423744;
      56670: inst = 32'd471859200;
      56671: inst = 32'd136314880;
      56672: inst = 32'd268468224;
      56673: inst = 32'd201348133;
      56674: inst = 32'd203423744;
      56675: inst = 32'd471859200;
      56676: inst = 32'd136314880;
      56677: inst = 32'd268468224;
      56678: inst = 32'd201348134;
      56679: inst = 32'd203423744;
      56680: inst = 32'd471859200;
      56681: inst = 32'd136314880;
      56682: inst = 32'd268468224;
      56683: inst = 32'd201348135;
      56684: inst = 32'd203423744;
      56685: inst = 32'd471859200;
      56686: inst = 32'd136314880;
      56687: inst = 32'd268468224;
      56688: inst = 32'd201348136;
      56689: inst = 32'd203423744;
      56690: inst = 32'd471859200;
      56691: inst = 32'd136314880;
      56692: inst = 32'd268468224;
      56693: inst = 32'd201348137;
      56694: inst = 32'd203423744;
      56695: inst = 32'd471859200;
      56696: inst = 32'd136314880;
      56697: inst = 32'd268468224;
      56698: inst = 32'd201348138;
      56699: inst = 32'd203423744;
      56700: inst = 32'd471859200;
      56701: inst = 32'd136314880;
      56702: inst = 32'd268468224;
      56703: inst = 32'd201348139;
      56704: inst = 32'd203423744;
      56705: inst = 32'd471859200;
      56706: inst = 32'd136314880;
      56707: inst = 32'd268468224;
      56708: inst = 32'd201348140;
      56709: inst = 32'd203423744;
      56710: inst = 32'd471859200;
      56711: inst = 32'd136314880;
      56712: inst = 32'd268468224;
      56713: inst = 32'd201348141;
      56714: inst = 32'd203423744;
      56715: inst = 32'd471859200;
      56716: inst = 32'd136314880;
      56717: inst = 32'd268468224;
      56718: inst = 32'd201348142;
      56719: inst = 32'd203423744;
      56720: inst = 32'd471859200;
      56721: inst = 32'd136314880;
      56722: inst = 32'd268468224;
      56723: inst = 32'd201348143;
      56724: inst = 32'd203423744;
      56725: inst = 32'd471859200;
      56726: inst = 32'd136314880;
      56727: inst = 32'd268468224;
      56728: inst = 32'd201348144;
      56729: inst = 32'd203423744;
      56730: inst = 32'd471859200;
      56731: inst = 32'd136314880;
      56732: inst = 32'd268468224;
      56733: inst = 32'd201348145;
      56734: inst = 32'd203423744;
      56735: inst = 32'd471859200;
      56736: inst = 32'd136314880;
      56737: inst = 32'd268468224;
      56738: inst = 32'd201348146;
      56739: inst = 32'd203423744;
      56740: inst = 32'd471859200;
      56741: inst = 32'd136314880;
      56742: inst = 32'd268468224;
      56743: inst = 32'd201348147;
      56744: inst = 32'd203423744;
      56745: inst = 32'd471859200;
      56746: inst = 32'd136314880;
      56747: inst = 32'd268468224;
      56748: inst = 32'd201348148;
      56749: inst = 32'd203423744;
      56750: inst = 32'd471859200;
      56751: inst = 32'd136314880;
      56752: inst = 32'd268468224;
      56753: inst = 32'd201348149;
      56754: inst = 32'd203423744;
      56755: inst = 32'd471859200;
      56756: inst = 32'd136314880;
      56757: inst = 32'd268468224;
      56758: inst = 32'd201348150;
      56759: inst = 32'd203423744;
      56760: inst = 32'd471859200;
      56761: inst = 32'd136314880;
      56762: inst = 32'd268468224;
      56763: inst = 32'd201348151;
      56764: inst = 32'd203423744;
      56765: inst = 32'd471859200;
      56766: inst = 32'd136314880;
      56767: inst = 32'd268468224;
      56768: inst = 32'd201348152;
      56769: inst = 32'd203423744;
      56770: inst = 32'd471859200;
      56771: inst = 32'd136314880;
      56772: inst = 32'd268468224;
      56773: inst = 32'd201348153;
      56774: inst = 32'd203423744;
      56775: inst = 32'd471859200;
      56776: inst = 32'd136314880;
      56777: inst = 32'd268468224;
      56778: inst = 32'd201348154;
      56779: inst = 32'd203423744;
      56780: inst = 32'd471859200;
      56781: inst = 32'd136314880;
      56782: inst = 32'd268468224;
      56783: inst = 32'd201348155;
      56784: inst = 32'd203423744;
      56785: inst = 32'd471859200;
      56786: inst = 32'd136314880;
      56787: inst = 32'd268468224;
      56788: inst = 32'd201348156;
      56789: inst = 32'd203423744;
      56790: inst = 32'd471859200;
      56791: inst = 32'd136314880;
      56792: inst = 32'd268468224;
      56793: inst = 32'd201348157;
      56794: inst = 32'd203423744;
      56795: inst = 32'd471859200;
      56796: inst = 32'd136314880;
      56797: inst = 32'd268468224;
      56798: inst = 32'd201348158;
      56799: inst = 32'd203423744;
      56800: inst = 32'd471859200;
      56801: inst = 32'd136314880;
      56802: inst = 32'd268468224;
      56803: inst = 32'd201348159;
      56804: inst = 32'd203423744;
      56805: inst = 32'd471859200;
      56806: inst = 32'd136314880;
      56807: inst = 32'd268468224;
      56808: inst = 32'd201348160;
      56809: inst = 32'd203423744;
      56810: inst = 32'd471859200;
      56811: inst = 32'd136314880;
      56812: inst = 32'd268468224;
      56813: inst = 32'd201348161;
      56814: inst = 32'd203423744;
      56815: inst = 32'd471859200;
      56816: inst = 32'd136314880;
      56817: inst = 32'd268468224;
      56818: inst = 32'd201348162;
      56819: inst = 32'd203423744;
      56820: inst = 32'd471859200;
      56821: inst = 32'd136314880;
      56822: inst = 32'd268468224;
      56823: inst = 32'd201348163;
      56824: inst = 32'd203423744;
      56825: inst = 32'd471859200;
      56826: inst = 32'd136314880;
      56827: inst = 32'd268468224;
      56828: inst = 32'd201348164;
      56829: inst = 32'd203423744;
      56830: inst = 32'd471859200;
      56831: inst = 32'd136314880;
      56832: inst = 32'd268468224;
      56833: inst = 32'd201348165;
      56834: inst = 32'd203423744;
      56835: inst = 32'd471859200;
      56836: inst = 32'd136314880;
      56837: inst = 32'd268468224;
      56838: inst = 32'd201348166;
      56839: inst = 32'd203423744;
      56840: inst = 32'd471859200;
      56841: inst = 32'd136314880;
      56842: inst = 32'd268468224;
      56843: inst = 32'd201348167;
      56844: inst = 32'd203423744;
      56845: inst = 32'd471859200;
      56846: inst = 32'd136314880;
      56847: inst = 32'd268468224;
      56848: inst = 32'd201348168;
      56849: inst = 32'd203423744;
      56850: inst = 32'd471859200;
      56851: inst = 32'd136314880;
      56852: inst = 32'd268468224;
      56853: inst = 32'd201348169;
      56854: inst = 32'd203423744;
      56855: inst = 32'd471859200;
      56856: inst = 32'd136314880;
      56857: inst = 32'd268468224;
      56858: inst = 32'd201348170;
      56859: inst = 32'd203423744;
      56860: inst = 32'd471859200;
      56861: inst = 32'd136314880;
      56862: inst = 32'd268468224;
      56863: inst = 32'd201348171;
      56864: inst = 32'd203423744;
      56865: inst = 32'd471859200;
      56866: inst = 32'd136314880;
      56867: inst = 32'd268468224;
      56868: inst = 32'd201348172;
      56869: inst = 32'd203423744;
      56870: inst = 32'd471859200;
      56871: inst = 32'd136314880;
      56872: inst = 32'd268468224;
      56873: inst = 32'd201348173;
      56874: inst = 32'd203423744;
      56875: inst = 32'd471859200;
      56876: inst = 32'd136314880;
      56877: inst = 32'd268468224;
      56878: inst = 32'd201348174;
      56879: inst = 32'd203423744;
      56880: inst = 32'd471859200;
      56881: inst = 32'd136314880;
      56882: inst = 32'd268468224;
      56883: inst = 32'd201348175;
      56884: inst = 32'd203423744;
      56885: inst = 32'd471859200;
      56886: inst = 32'd136314880;
      56887: inst = 32'd268468224;
      56888: inst = 32'd201348176;
      56889: inst = 32'd203423744;
      56890: inst = 32'd471859200;
      56891: inst = 32'd136314880;
      56892: inst = 32'd268468224;
      56893: inst = 32'd201348177;
      56894: inst = 32'd203423744;
      56895: inst = 32'd471859200;
      56896: inst = 32'd136314880;
      56897: inst = 32'd268468224;
      56898: inst = 32'd201348178;
      56899: inst = 32'd203423744;
      56900: inst = 32'd471859200;
      56901: inst = 32'd136314880;
      56902: inst = 32'd268468224;
      56903: inst = 32'd201348179;
      56904: inst = 32'd203423744;
      56905: inst = 32'd471859200;
      56906: inst = 32'd136314880;
      56907: inst = 32'd268468224;
      56908: inst = 32'd201348180;
      56909: inst = 32'd203423744;
      56910: inst = 32'd471859200;
      56911: inst = 32'd136314880;
      56912: inst = 32'd268468224;
      56913: inst = 32'd201348181;
      56914: inst = 32'd203423744;
      56915: inst = 32'd471859200;
      56916: inst = 32'd136314880;
      56917: inst = 32'd268468224;
      56918: inst = 32'd201348182;
      56919: inst = 32'd203423744;
      56920: inst = 32'd471859200;
      56921: inst = 32'd136314880;
      56922: inst = 32'd268468224;
      56923: inst = 32'd201348183;
      56924: inst = 32'd203423744;
      56925: inst = 32'd471859200;
      56926: inst = 32'd136314880;
      56927: inst = 32'd268468224;
      56928: inst = 32'd201348184;
      56929: inst = 32'd203423744;
      56930: inst = 32'd471859200;
      56931: inst = 32'd136314880;
      56932: inst = 32'd268468224;
      56933: inst = 32'd201348185;
      56934: inst = 32'd203423744;
      56935: inst = 32'd471859200;
      56936: inst = 32'd136314880;
      56937: inst = 32'd268468224;
      56938: inst = 32'd201348186;
      56939: inst = 32'd203423744;
      56940: inst = 32'd471859200;
      56941: inst = 32'd136314880;
      56942: inst = 32'd268468224;
      56943: inst = 32'd201348187;
      56944: inst = 32'd203423744;
      56945: inst = 32'd471859200;
      56946: inst = 32'd136314880;
      56947: inst = 32'd268468224;
      56948: inst = 32'd201348188;
      56949: inst = 32'd203423744;
      56950: inst = 32'd471859200;
      56951: inst = 32'd136314880;
      56952: inst = 32'd268468224;
      56953: inst = 32'd201348189;
      56954: inst = 32'd203423744;
      56955: inst = 32'd471859200;
      56956: inst = 32'd136314880;
      56957: inst = 32'd268468224;
      56958: inst = 32'd201348190;
      56959: inst = 32'd203423744;
      56960: inst = 32'd471859200;
      56961: inst = 32'd136314880;
      56962: inst = 32'd268468224;
      56963: inst = 32'd201348191;
      56964: inst = 32'd203423744;
      56965: inst = 32'd471859200;
      56966: inst = 32'd136314880;
      56967: inst = 32'd268468224;
      56968: inst = 32'd201348192;
      56969: inst = 32'd203423744;
      56970: inst = 32'd471859200;
      56971: inst = 32'd136314880;
      56972: inst = 32'd268468224;
      56973: inst = 32'd201348193;
      56974: inst = 32'd203423744;
      56975: inst = 32'd471859200;
      56976: inst = 32'd136314880;
      56977: inst = 32'd268468224;
      56978: inst = 32'd201348194;
      56979: inst = 32'd203423744;
      56980: inst = 32'd471859200;
      56981: inst = 32'd136314880;
      56982: inst = 32'd268468224;
      56983: inst = 32'd201348195;
      56984: inst = 32'd203423744;
      56985: inst = 32'd471859200;
      56986: inst = 32'd136314880;
      56987: inst = 32'd268468224;
      56988: inst = 32'd201348196;
      56989: inst = 32'd203423744;
      56990: inst = 32'd471859200;
      56991: inst = 32'd136314880;
      56992: inst = 32'd268468224;
      56993: inst = 32'd201348197;
      56994: inst = 32'd203423744;
      56995: inst = 32'd471859200;
      56996: inst = 32'd136314880;
      56997: inst = 32'd268468224;
      56998: inst = 32'd201348198;
      56999: inst = 32'd203423744;
      57000: inst = 32'd471859200;
      57001: inst = 32'd136314880;
      57002: inst = 32'd268468224;
      57003: inst = 32'd201348199;
      57004: inst = 32'd203423744;
      57005: inst = 32'd471859200;
      57006: inst = 32'd136314880;
      57007: inst = 32'd268468224;
      57008: inst = 32'd201348200;
      57009: inst = 32'd203423744;
      57010: inst = 32'd471859200;
      57011: inst = 32'd136314880;
      57012: inst = 32'd268468224;
      57013: inst = 32'd201348201;
      57014: inst = 32'd203423744;
      57015: inst = 32'd471859200;
      57016: inst = 32'd136314880;
      57017: inst = 32'd268468224;
      57018: inst = 32'd201348202;
      57019: inst = 32'd203423744;
      57020: inst = 32'd471859200;
      57021: inst = 32'd136314880;
      57022: inst = 32'd268468224;
      57023: inst = 32'd201348203;
      57024: inst = 32'd203423744;
      57025: inst = 32'd471859200;
      57026: inst = 32'd136314880;
      57027: inst = 32'd268468224;
      57028: inst = 32'd201348204;
      57029: inst = 32'd203423744;
      57030: inst = 32'd471859200;
      57031: inst = 32'd136314880;
      57032: inst = 32'd268468224;
      57033: inst = 32'd201348205;
      57034: inst = 32'd203423744;
      57035: inst = 32'd471859200;
      57036: inst = 32'd136314880;
      57037: inst = 32'd268468224;
      57038: inst = 32'd201348206;
      57039: inst = 32'd203423744;
      57040: inst = 32'd471859200;
      57041: inst = 32'd136314880;
      57042: inst = 32'd268468224;
      57043: inst = 32'd201348207;
      57044: inst = 32'd203423744;
      57045: inst = 32'd471859200;
      57046: inst = 32'd136314880;
      57047: inst = 32'd268468224;
      57048: inst = 32'd201348208;
      57049: inst = 32'd203423744;
      57050: inst = 32'd471859200;
      57051: inst = 32'd136314880;
      57052: inst = 32'd268468224;
      57053: inst = 32'd201348209;
      57054: inst = 32'd203423744;
      57055: inst = 32'd471859200;
      57056: inst = 32'd136314880;
      57057: inst = 32'd268468224;
      57058: inst = 32'd201348210;
      57059: inst = 32'd203423744;
      57060: inst = 32'd471859200;
      57061: inst = 32'd136314880;
      57062: inst = 32'd268468224;
      57063: inst = 32'd201348211;
      57064: inst = 32'd203423744;
      57065: inst = 32'd471859200;
      57066: inst = 32'd136314880;
      57067: inst = 32'd268468224;
      57068: inst = 32'd201348212;
      57069: inst = 32'd203423744;
      57070: inst = 32'd471859200;
      57071: inst = 32'd136314880;
      57072: inst = 32'd268468224;
      57073: inst = 32'd201348213;
      57074: inst = 32'd203423744;
      57075: inst = 32'd471859200;
      57076: inst = 32'd136314880;
      57077: inst = 32'd268468224;
      57078: inst = 32'd201348214;
      57079: inst = 32'd203423744;
      57080: inst = 32'd471859200;
      57081: inst = 32'd136314880;
      57082: inst = 32'd268468224;
      57083: inst = 32'd201348215;
      57084: inst = 32'd203423744;
      57085: inst = 32'd471859200;
      57086: inst = 32'd136314880;
      57087: inst = 32'd268468224;
      57088: inst = 32'd201348216;
      57089: inst = 32'd203423744;
      57090: inst = 32'd471859200;
      57091: inst = 32'd136314880;
      57092: inst = 32'd268468224;
      57093: inst = 32'd201348217;
      57094: inst = 32'd203423744;
      57095: inst = 32'd471859200;
      57096: inst = 32'd136314880;
      57097: inst = 32'd268468224;
      57098: inst = 32'd201348218;
      57099: inst = 32'd203423744;
      57100: inst = 32'd471859200;
      57101: inst = 32'd136314880;
      57102: inst = 32'd268468224;
      57103: inst = 32'd201348219;
      57104: inst = 32'd203423744;
      57105: inst = 32'd471859200;
      57106: inst = 32'd136314880;
      57107: inst = 32'd268468224;
      57108: inst = 32'd201348220;
      57109: inst = 32'd203423744;
      57110: inst = 32'd471859200;
      57111: inst = 32'd136314880;
      57112: inst = 32'd268468224;
      57113: inst = 32'd201348221;
      57114: inst = 32'd203423744;
      57115: inst = 32'd471859200;
      57116: inst = 32'd136314880;
      57117: inst = 32'd268468224;
      57118: inst = 32'd201348222;
      57119: inst = 32'd203423744;
      57120: inst = 32'd471859200;
      57121: inst = 32'd136314880;
      57122: inst = 32'd268468224;
      57123: inst = 32'd201348223;
      57124: inst = 32'd203423744;
      57125: inst = 32'd471859200;
      57126: inst = 32'd136314880;
      57127: inst = 32'd268468224;
      57128: inst = 32'd201348224;
      57129: inst = 32'd203423744;
      57130: inst = 32'd471859200;
      57131: inst = 32'd136314880;
      57132: inst = 32'd268468224;
      57133: inst = 32'd201348225;
      57134: inst = 32'd203423744;
      57135: inst = 32'd471859200;
      57136: inst = 32'd136314880;
      57137: inst = 32'd268468224;
      57138: inst = 32'd201348226;
      57139: inst = 32'd203423744;
      57140: inst = 32'd471859200;
      57141: inst = 32'd136314880;
      57142: inst = 32'd268468224;
      57143: inst = 32'd201348227;
      57144: inst = 32'd203423744;
      57145: inst = 32'd471859200;
      57146: inst = 32'd136314880;
      57147: inst = 32'd268468224;
      57148: inst = 32'd201348228;
      57149: inst = 32'd203423744;
      57150: inst = 32'd471859200;
      57151: inst = 32'd136314880;
      57152: inst = 32'd268468224;
      57153: inst = 32'd201348229;
      57154: inst = 32'd203423744;
      57155: inst = 32'd471859200;
      57156: inst = 32'd136314880;
      57157: inst = 32'd268468224;
      57158: inst = 32'd201348230;
      57159: inst = 32'd203423744;
      57160: inst = 32'd471859200;
      57161: inst = 32'd136314880;
      57162: inst = 32'd268468224;
      57163: inst = 32'd201348231;
      57164: inst = 32'd203423744;
      57165: inst = 32'd471859200;
      57166: inst = 32'd136314880;
      57167: inst = 32'd268468224;
      57168: inst = 32'd201348232;
      57169: inst = 32'd203423744;
      57170: inst = 32'd471859200;
      57171: inst = 32'd136314880;
      57172: inst = 32'd268468224;
      57173: inst = 32'd201348233;
      57174: inst = 32'd203423744;
      57175: inst = 32'd471859200;
      57176: inst = 32'd136314880;
      57177: inst = 32'd268468224;
      57178: inst = 32'd201348234;
      57179: inst = 32'd203423744;
      57180: inst = 32'd471859200;
      57181: inst = 32'd136314880;
      57182: inst = 32'd268468224;
      57183: inst = 32'd201348235;
      57184: inst = 32'd203423744;
      57185: inst = 32'd471859200;
      57186: inst = 32'd136314880;
      57187: inst = 32'd268468224;
      57188: inst = 32'd201348236;
      57189: inst = 32'd203423744;
      57190: inst = 32'd471859200;
      57191: inst = 32'd136314880;
      57192: inst = 32'd268468224;
      57193: inst = 32'd201348237;
      57194: inst = 32'd203423744;
      57195: inst = 32'd471859200;
      57196: inst = 32'd136314880;
      57197: inst = 32'd268468224;
      57198: inst = 32'd201348238;
      57199: inst = 32'd203423744;
      57200: inst = 32'd471859200;
      57201: inst = 32'd136314880;
      57202: inst = 32'd268468224;
      57203: inst = 32'd201348239;
      57204: inst = 32'd203423744;
      57205: inst = 32'd471859200;
      57206: inst = 32'd136314880;
      57207: inst = 32'd268468224;
      57208: inst = 32'd201348240;
      57209: inst = 32'd203423744;
      57210: inst = 32'd471859200;
      57211: inst = 32'd136314880;
      57212: inst = 32'd268468224;
      57213: inst = 32'd201348241;
      57214: inst = 32'd203423744;
      57215: inst = 32'd471859200;
      57216: inst = 32'd136314880;
      57217: inst = 32'd268468224;
      57218: inst = 32'd201348242;
      57219: inst = 32'd203423744;
      57220: inst = 32'd471859200;
      57221: inst = 32'd136314880;
      57222: inst = 32'd268468224;
      57223: inst = 32'd201348243;
      57224: inst = 32'd203423744;
      57225: inst = 32'd471859200;
      57226: inst = 32'd136314880;
      57227: inst = 32'd268468224;
      57228: inst = 32'd201348244;
      57229: inst = 32'd203423744;
      57230: inst = 32'd471859200;
      57231: inst = 32'd136314880;
      57232: inst = 32'd268468224;
      57233: inst = 32'd201348245;
      57234: inst = 32'd203423744;
      57235: inst = 32'd471859200;
      57236: inst = 32'd136314880;
      57237: inst = 32'd268468224;
      57238: inst = 32'd201348246;
      57239: inst = 32'd203423744;
      57240: inst = 32'd471859200;
      57241: inst = 32'd136314880;
      57242: inst = 32'd268468224;
      57243: inst = 32'd201348247;
      57244: inst = 32'd203423744;
      57245: inst = 32'd471859200;
      57246: inst = 32'd136314880;
      57247: inst = 32'd268468224;
      57248: inst = 32'd201348248;
      57249: inst = 32'd203423744;
      57250: inst = 32'd471859200;
      57251: inst = 32'd136314880;
      57252: inst = 32'd268468224;
      57253: inst = 32'd201348249;
      57254: inst = 32'd203423744;
      57255: inst = 32'd471859200;
      57256: inst = 32'd136314880;
      57257: inst = 32'd268468224;
      57258: inst = 32'd201348250;
      57259: inst = 32'd203423744;
      57260: inst = 32'd471859200;
      57261: inst = 32'd136314880;
      57262: inst = 32'd268468224;
      57263: inst = 32'd201348251;
      57264: inst = 32'd203423744;
      57265: inst = 32'd471859200;
      57266: inst = 32'd136314880;
      57267: inst = 32'd268468224;
      57268: inst = 32'd201348252;
      57269: inst = 32'd203423744;
      57270: inst = 32'd471859200;
      57271: inst = 32'd136314880;
      57272: inst = 32'd268468224;
      57273: inst = 32'd201348253;
      57274: inst = 32'd203423744;
      57275: inst = 32'd471859200;
      57276: inst = 32'd136314880;
      57277: inst = 32'd268468224;
      57278: inst = 32'd201348254;
      57279: inst = 32'd203423744;
      57280: inst = 32'd471859200;
      57281: inst = 32'd136314880;
      57282: inst = 32'd268468224;
      57283: inst = 32'd201348255;
      57284: inst = 32'd203423744;
      57285: inst = 32'd471859200;
      57286: inst = 32'd136314880;
      57287: inst = 32'd268468224;
      57288: inst = 32'd201348256;
      57289: inst = 32'd203423744;
      57290: inst = 32'd471859200;
      57291: inst = 32'd136314880;
      57292: inst = 32'd268468224;
      57293: inst = 32'd201348257;
      57294: inst = 32'd203423744;
      57295: inst = 32'd471859200;
      57296: inst = 32'd136314880;
      57297: inst = 32'd268468224;
      57298: inst = 32'd201348258;
      57299: inst = 32'd203423744;
      57300: inst = 32'd471859200;
      57301: inst = 32'd136314880;
      57302: inst = 32'd268468224;
      57303: inst = 32'd201348259;
      57304: inst = 32'd203423744;
      57305: inst = 32'd471859200;
      57306: inst = 32'd136314880;
      57307: inst = 32'd268468224;
      57308: inst = 32'd201348260;
      57309: inst = 32'd203423744;
      57310: inst = 32'd471859200;
      57311: inst = 32'd136314880;
      57312: inst = 32'd268468224;
      57313: inst = 32'd201348261;
      57314: inst = 32'd203423744;
      57315: inst = 32'd471859200;
      57316: inst = 32'd136314880;
      57317: inst = 32'd268468224;
      57318: inst = 32'd201348262;
      57319: inst = 32'd203423744;
      57320: inst = 32'd471859200;
      57321: inst = 32'd136314880;
      57322: inst = 32'd268468224;
      57323: inst = 32'd201348263;
      57324: inst = 32'd203423744;
      57325: inst = 32'd471859200;
      57326: inst = 32'd136314880;
      57327: inst = 32'd268468224;
      57328: inst = 32'd201348264;
      57329: inst = 32'd203423744;
      57330: inst = 32'd471859200;
      57331: inst = 32'd136314880;
      57332: inst = 32'd268468224;
      57333: inst = 32'd201348265;
      57334: inst = 32'd203423744;
      57335: inst = 32'd471859200;
      57336: inst = 32'd136314880;
      57337: inst = 32'd268468224;
      57338: inst = 32'd201348266;
      57339: inst = 32'd203423744;
      57340: inst = 32'd471859200;
      57341: inst = 32'd136314880;
      57342: inst = 32'd268468224;
      57343: inst = 32'd201348267;
      57344: inst = 32'd203423744;
      57345: inst = 32'd471859200;
      57346: inst = 32'd136314880;
      57347: inst = 32'd268468224;
      57348: inst = 32'd201348268;
      57349: inst = 32'd203423744;
      57350: inst = 32'd471859200;
      57351: inst = 32'd136314880;
      57352: inst = 32'd268468224;
      57353: inst = 32'd201348269;
      57354: inst = 32'd203423744;
      57355: inst = 32'd471859200;
      57356: inst = 32'd136314880;
      57357: inst = 32'd268468224;
      57358: inst = 32'd201348270;
      57359: inst = 32'd203423744;
      57360: inst = 32'd471859200;
      57361: inst = 32'd136314880;
      57362: inst = 32'd268468224;
      57363: inst = 32'd201348271;
      57364: inst = 32'd203423744;
      57365: inst = 32'd471859200;
      57366: inst = 32'd136314880;
      57367: inst = 32'd268468224;
      57368: inst = 32'd201348272;
      57369: inst = 32'd203423744;
      57370: inst = 32'd471859200;
      57371: inst = 32'd136314880;
      57372: inst = 32'd268468224;
      57373: inst = 32'd201348273;
      57374: inst = 32'd203423744;
      57375: inst = 32'd471859200;
      57376: inst = 32'd136314880;
      57377: inst = 32'd268468224;
      57378: inst = 32'd201348274;
      57379: inst = 32'd203423744;
      57380: inst = 32'd471859200;
      57381: inst = 32'd136314880;
      57382: inst = 32'd268468224;
      57383: inst = 32'd201348275;
      57384: inst = 32'd203423744;
      57385: inst = 32'd471859200;
      57386: inst = 32'd136314880;
      57387: inst = 32'd268468224;
      57388: inst = 32'd201348276;
      57389: inst = 32'd203423744;
      57390: inst = 32'd471859200;
      57391: inst = 32'd136314880;
      57392: inst = 32'd268468224;
      57393: inst = 32'd201348277;
      57394: inst = 32'd203423744;
      57395: inst = 32'd471859200;
      57396: inst = 32'd136314880;
      57397: inst = 32'd268468224;
      57398: inst = 32'd201348278;
      57399: inst = 32'd203423744;
      57400: inst = 32'd471859200;
      57401: inst = 32'd136314880;
      57402: inst = 32'd268468224;
      57403: inst = 32'd201348279;
      57404: inst = 32'd203423744;
      57405: inst = 32'd471859200;
      57406: inst = 32'd136314880;
      57407: inst = 32'd268468224;
      57408: inst = 32'd201348280;
      57409: inst = 32'd203423744;
      57410: inst = 32'd471859200;
      57411: inst = 32'd136314880;
      57412: inst = 32'd268468224;
      57413: inst = 32'd201348281;
      57414: inst = 32'd203423744;
      57415: inst = 32'd471859200;
      57416: inst = 32'd136314880;
      57417: inst = 32'd268468224;
      57418: inst = 32'd201348282;
      57419: inst = 32'd203423744;
      57420: inst = 32'd471859200;
      57421: inst = 32'd136314880;
      57422: inst = 32'd268468224;
      57423: inst = 32'd201348283;
      57424: inst = 32'd203423744;
      57425: inst = 32'd471859200;
      57426: inst = 32'd136314880;
      57427: inst = 32'd268468224;
      57428: inst = 32'd201348284;
      57429: inst = 32'd203423744;
      57430: inst = 32'd471859200;
      57431: inst = 32'd136314880;
      57432: inst = 32'd268468224;
      57433: inst = 32'd201348285;
      57434: inst = 32'd203423744;
      57435: inst = 32'd471859200;
      57436: inst = 32'd136314880;
      57437: inst = 32'd268468224;
      57438: inst = 32'd201348286;
      57439: inst = 32'd203423744;
      57440: inst = 32'd471859200;
      57441: inst = 32'd136314880;
      57442: inst = 32'd268468224;
      57443: inst = 32'd201348287;
      57444: inst = 32'd203423744;
      57445: inst = 32'd471859200;
      57446: inst = 32'd136314880;
      57447: inst = 32'd268468224;
      57448: inst = 32'd201348288;
      57449: inst = 32'd203423744;
      57450: inst = 32'd471859200;
      57451: inst = 32'd136314880;
      57452: inst = 32'd268468224;
      57453: inst = 32'd201348289;
      57454: inst = 32'd203423744;
      57455: inst = 32'd471859200;
      57456: inst = 32'd136314880;
      57457: inst = 32'd268468224;
      57458: inst = 32'd201348290;
      57459: inst = 32'd203423744;
      57460: inst = 32'd471859200;
      57461: inst = 32'd136314880;
      57462: inst = 32'd268468224;
      57463: inst = 32'd201348291;
      57464: inst = 32'd203423744;
      57465: inst = 32'd471859200;
      57466: inst = 32'd136314880;
      57467: inst = 32'd268468224;
      57468: inst = 32'd201348292;
      57469: inst = 32'd203423744;
      57470: inst = 32'd471859200;
      57471: inst = 32'd136314880;
      57472: inst = 32'd268468224;
      57473: inst = 32'd201348293;
      57474: inst = 32'd203423744;
      57475: inst = 32'd471859200;
      57476: inst = 32'd136314880;
      57477: inst = 32'd268468224;
      57478: inst = 32'd201348294;
      57479: inst = 32'd203423744;
      57480: inst = 32'd471859200;
      57481: inst = 32'd136314880;
      57482: inst = 32'd268468224;
      57483: inst = 32'd201348295;
      57484: inst = 32'd203423744;
      57485: inst = 32'd471859200;
      57486: inst = 32'd136314880;
      57487: inst = 32'd268468224;
      57488: inst = 32'd201348296;
      57489: inst = 32'd203423744;
      57490: inst = 32'd471859200;
      57491: inst = 32'd136314880;
      57492: inst = 32'd268468224;
      57493: inst = 32'd201348297;
      57494: inst = 32'd203423744;
      57495: inst = 32'd471859200;
      57496: inst = 32'd136314880;
      57497: inst = 32'd268468224;
      57498: inst = 32'd201348298;
      57499: inst = 32'd203423744;
      57500: inst = 32'd471859200;
      57501: inst = 32'd136314880;
      57502: inst = 32'd268468224;
      57503: inst = 32'd201348299;
      57504: inst = 32'd203423744;
      57505: inst = 32'd471859200;
      57506: inst = 32'd136314880;
      57507: inst = 32'd268468224;
      57508: inst = 32'd201348300;
      57509: inst = 32'd203423744;
      57510: inst = 32'd471859200;
      57511: inst = 32'd136314880;
      57512: inst = 32'd268468224;
      57513: inst = 32'd201348301;
      57514: inst = 32'd203423744;
      57515: inst = 32'd471859200;
      57516: inst = 32'd136314880;
      57517: inst = 32'd268468224;
      57518: inst = 32'd201348302;
      57519: inst = 32'd203423744;
      57520: inst = 32'd471859200;
      57521: inst = 32'd136314880;
      57522: inst = 32'd268468224;
      57523: inst = 32'd201348303;
      57524: inst = 32'd203423744;
      57525: inst = 32'd471859200;
      57526: inst = 32'd136314880;
      57527: inst = 32'd268468224;
      57528: inst = 32'd201348304;
      57529: inst = 32'd203423744;
      57530: inst = 32'd471859200;
      57531: inst = 32'd136314880;
      57532: inst = 32'd268468224;
      57533: inst = 32'd201348305;
      57534: inst = 32'd203423744;
      57535: inst = 32'd471859200;
      57536: inst = 32'd136314880;
      57537: inst = 32'd268468224;
      57538: inst = 32'd201348306;
      57539: inst = 32'd203423744;
      57540: inst = 32'd471859200;
      57541: inst = 32'd136314880;
      57542: inst = 32'd268468224;
      57543: inst = 32'd201348307;
      57544: inst = 32'd203423744;
      57545: inst = 32'd471859200;
      57546: inst = 32'd136314880;
      57547: inst = 32'd268468224;
      57548: inst = 32'd201348308;
      57549: inst = 32'd203423744;
      57550: inst = 32'd471859200;
      57551: inst = 32'd136314880;
      57552: inst = 32'd268468224;
      57553: inst = 32'd201348309;
      57554: inst = 32'd203423744;
      57555: inst = 32'd471859200;
      57556: inst = 32'd136314880;
      57557: inst = 32'd268468224;
      57558: inst = 32'd201348310;
      57559: inst = 32'd203423744;
      57560: inst = 32'd471859200;
      57561: inst = 32'd136314880;
      57562: inst = 32'd268468224;
      57563: inst = 32'd201348311;
      57564: inst = 32'd203423744;
      57565: inst = 32'd471859200;
      57566: inst = 32'd136314880;
      57567: inst = 32'd268468224;
      57568: inst = 32'd201348312;
      57569: inst = 32'd203423744;
      57570: inst = 32'd471859200;
      57571: inst = 32'd136314880;
      57572: inst = 32'd268468224;
      57573: inst = 32'd201348313;
      57574: inst = 32'd203423744;
      57575: inst = 32'd471859200;
      57576: inst = 32'd136314880;
      57577: inst = 32'd268468224;
      57578: inst = 32'd201348314;
      57579: inst = 32'd203423744;
      57580: inst = 32'd471859200;
      57581: inst = 32'd136314880;
      57582: inst = 32'd268468224;
      57583: inst = 32'd201348315;
      57584: inst = 32'd203423744;
      57585: inst = 32'd471859200;
      57586: inst = 32'd136314880;
      57587: inst = 32'd268468224;
      57588: inst = 32'd201348316;
      57589: inst = 32'd203423744;
      57590: inst = 32'd471859200;
      57591: inst = 32'd136314880;
      57592: inst = 32'd268468224;
      57593: inst = 32'd201348317;
      57594: inst = 32'd203423744;
      57595: inst = 32'd471859200;
      57596: inst = 32'd136314880;
      57597: inst = 32'd268468224;
      57598: inst = 32'd201348318;
      57599: inst = 32'd203423744;
      57600: inst = 32'd471859200;
      57601: inst = 32'd136314880;
      57602: inst = 32'd268468224;
      57603: inst = 32'd201348319;
      57604: inst = 32'd203423744;
      57605: inst = 32'd471859200;
      57606: inst = 32'd136314880;
      57607: inst = 32'd268468224;
      57608: inst = 32'd201348320;
      57609: inst = 32'd203423744;
      57610: inst = 32'd471859200;
      57611: inst = 32'd136314880;
      57612: inst = 32'd268468224;
      57613: inst = 32'd201348321;
      57614: inst = 32'd203423744;
      57615: inst = 32'd471859200;
      57616: inst = 32'd136314880;
      57617: inst = 32'd268468224;
      57618: inst = 32'd201348322;
      57619: inst = 32'd203423744;
      57620: inst = 32'd471859200;
      57621: inst = 32'd136314880;
      57622: inst = 32'd268468224;
      57623: inst = 32'd201348323;
      57624: inst = 32'd203423744;
      57625: inst = 32'd471859200;
      57626: inst = 32'd136314880;
      57627: inst = 32'd268468224;
      57628: inst = 32'd201348324;
      57629: inst = 32'd203423744;
      57630: inst = 32'd471859200;
      57631: inst = 32'd136314880;
      57632: inst = 32'd268468224;
      57633: inst = 32'd201348325;
      57634: inst = 32'd203423744;
      57635: inst = 32'd471859200;
      57636: inst = 32'd136314880;
      57637: inst = 32'd268468224;
      57638: inst = 32'd201348326;
      57639: inst = 32'd203423744;
      57640: inst = 32'd471859200;
      57641: inst = 32'd136314880;
      57642: inst = 32'd268468224;
      57643: inst = 32'd201348327;
      57644: inst = 32'd203423744;
      57645: inst = 32'd471859200;
      57646: inst = 32'd136314880;
      57647: inst = 32'd268468224;
      57648: inst = 32'd201348328;
      57649: inst = 32'd203423744;
      57650: inst = 32'd471859200;
      57651: inst = 32'd136314880;
      57652: inst = 32'd268468224;
      57653: inst = 32'd201348329;
      57654: inst = 32'd203423744;
      57655: inst = 32'd471859200;
      57656: inst = 32'd136314880;
      57657: inst = 32'd268468224;
      57658: inst = 32'd201348330;
      57659: inst = 32'd203423744;
      57660: inst = 32'd471859200;
      57661: inst = 32'd136314880;
      57662: inst = 32'd268468224;
      57663: inst = 32'd201348331;
      57664: inst = 32'd203423744;
      57665: inst = 32'd471859200;
      57666: inst = 32'd136314880;
      57667: inst = 32'd268468224;
      57668: inst = 32'd201348332;
      57669: inst = 32'd203423744;
      57670: inst = 32'd471859200;
      57671: inst = 32'd136314880;
      57672: inst = 32'd268468224;
      57673: inst = 32'd201348333;
      57674: inst = 32'd203423744;
      57675: inst = 32'd471859200;
      57676: inst = 32'd136314880;
      57677: inst = 32'd268468224;
      57678: inst = 32'd201348334;
      57679: inst = 32'd203423744;
      57680: inst = 32'd471859200;
      57681: inst = 32'd136314880;
      57682: inst = 32'd268468224;
      57683: inst = 32'd201348335;
      57684: inst = 32'd203423744;
      57685: inst = 32'd471859200;
      57686: inst = 32'd136314880;
      57687: inst = 32'd268468224;
      57688: inst = 32'd201348336;
      57689: inst = 32'd203423744;
      57690: inst = 32'd471859200;
      57691: inst = 32'd136314880;
      57692: inst = 32'd268468224;
      57693: inst = 32'd201348337;
      57694: inst = 32'd203423744;
      57695: inst = 32'd471859200;
      57696: inst = 32'd136314880;
      57697: inst = 32'd268468224;
      57698: inst = 32'd201348338;
      57699: inst = 32'd203423744;
      57700: inst = 32'd471859200;
      57701: inst = 32'd136314880;
      57702: inst = 32'd268468224;
      57703: inst = 32'd201348339;
      57704: inst = 32'd203423744;
      57705: inst = 32'd471859200;
      57706: inst = 32'd136314880;
      57707: inst = 32'd268468224;
      57708: inst = 32'd201348340;
      57709: inst = 32'd203423744;
      57710: inst = 32'd471859200;
      57711: inst = 32'd136314880;
      57712: inst = 32'd268468224;
      57713: inst = 32'd201348341;
      57714: inst = 32'd203423744;
      57715: inst = 32'd471859200;
      57716: inst = 32'd136314880;
      57717: inst = 32'd268468224;
      57718: inst = 32'd201348342;
      57719: inst = 32'd203423744;
      57720: inst = 32'd471859200;
      57721: inst = 32'd136314880;
      57722: inst = 32'd268468224;
      57723: inst = 32'd201348343;
      57724: inst = 32'd203423744;
      57725: inst = 32'd471859200;
      57726: inst = 32'd136314880;
      57727: inst = 32'd268468224;
      57728: inst = 32'd201348344;
      57729: inst = 32'd203423744;
      57730: inst = 32'd471859200;
      57731: inst = 32'd136314880;
      57732: inst = 32'd268468224;
      57733: inst = 32'd201348345;
      57734: inst = 32'd203423744;
      57735: inst = 32'd471859200;
      57736: inst = 32'd136314880;
      57737: inst = 32'd268468224;
      57738: inst = 32'd201348346;
      57739: inst = 32'd203423744;
      57740: inst = 32'd471859200;
      57741: inst = 32'd136314880;
      57742: inst = 32'd268468224;
      57743: inst = 32'd201348347;
      57744: inst = 32'd203423744;
      57745: inst = 32'd471859200;
      57746: inst = 32'd136314880;
      57747: inst = 32'd268468224;
      57748: inst = 32'd201348348;
      57749: inst = 32'd203423744;
      57750: inst = 32'd471859200;
      57751: inst = 32'd136314880;
      57752: inst = 32'd268468224;
      57753: inst = 32'd201348349;
      57754: inst = 32'd203423744;
      57755: inst = 32'd471859200;
      57756: inst = 32'd136314880;
      57757: inst = 32'd268468224;
      57758: inst = 32'd201348350;
      57759: inst = 32'd203423744;
      57760: inst = 32'd471859200;
      57761: inst = 32'd136314880;
      57762: inst = 32'd268468224;
      57763: inst = 32'd201348351;
      57764: inst = 32'd203423744;
      57765: inst = 32'd471859200;
      57766: inst = 32'd136314880;
      57767: inst = 32'd268468224;
      57768: inst = 32'd201348352;
      57769: inst = 32'd203423744;
      57770: inst = 32'd471859200;
      57771: inst = 32'd136314880;
      57772: inst = 32'd268468224;
      57773: inst = 32'd201348353;
      57774: inst = 32'd203423744;
      57775: inst = 32'd471859200;
      57776: inst = 32'd136314880;
      57777: inst = 32'd268468224;
      57778: inst = 32'd201348354;
      57779: inst = 32'd203423744;
      57780: inst = 32'd471859200;
      57781: inst = 32'd136314880;
      57782: inst = 32'd268468224;
      57783: inst = 32'd201348355;
      57784: inst = 32'd203423744;
      57785: inst = 32'd471859200;
      57786: inst = 32'd136314880;
      57787: inst = 32'd268468224;
      57788: inst = 32'd201348356;
      57789: inst = 32'd203423744;
      57790: inst = 32'd471859200;
      57791: inst = 32'd136314880;
      57792: inst = 32'd268468224;
      57793: inst = 32'd201348357;
      57794: inst = 32'd203423744;
      57795: inst = 32'd471859200;
      57796: inst = 32'd136314880;
      57797: inst = 32'd268468224;
      57798: inst = 32'd201348358;
      57799: inst = 32'd203423744;
      57800: inst = 32'd471859200;
      57801: inst = 32'd136314880;
      57802: inst = 32'd268468224;
      57803: inst = 32'd201348359;
      57804: inst = 32'd203423744;
      57805: inst = 32'd471859200;
      57806: inst = 32'd136314880;
      57807: inst = 32'd268468224;
      57808: inst = 32'd201348360;
      57809: inst = 32'd203423744;
      57810: inst = 32'd471859200;
      57811: inst = 32'd136314880;
      57812: inst = 32'd268468224;
      57813: inst = 32'd201348361;
      57814: inst = 32'd203423744;
      57815: inst = 32'd471859200;
      57816: inst = 32'd136314880;
      57817: inst = 32'd268468224;
      57818: inst = 32'd201348362;
      57819: inst = 32'd203423744;
      57820: inst = 32'd471859200;
      57821: inst = 32'd136314880;
      57822: inst = 32'd268468224;
      57823: inst = 32'd201348363;
      57824: inst = 32'd203423744;
      57825: inst = 32'd471859200;
      57826: inst = 32'd136314880;
      57827: inst = 32'd268468224;
      57828: inst = 32'd201348364;
      57829: inst = 32'd203423744;
      57830: inst = 32'd471859200;
      57831: inst = 32'd136314880;
      57832: inst = 32'd268468224;
      57833: inst = 32'd201348365;
      57834: inst = 32'd203423744;
      57835: inst = 32'd471859200;
      57836: inst = 32'd136314880;
      57837: inst = 32'd268468224;
      57838: inst = 32'd201348366;
      57839: inst = 32'd203423744;
      57840: inst = 32'd471859200;
      57841: inst = 32'd136314880;
      57842: inst = 32'd268468224;
      57843: inst = 32'd201348367;
      57844: inst = 32'd203423744;
      57845: inst = 32'd471859200;
      57846: inst = 32'd136314880;
      57847: inst = 32'd268468224;
      57848: inst = 32'd201348368;
      57849: inst = 32'd203423744;
      57850: inst = 32'd471859200;
      57851: inst = 32'd136314880;
      57852: inst = 32'd268468224;
      57853: inst = 32'd201348369;
      57854: inst = 32'd203423744;
      57855: inst = 32'd471859200;
      57856: inst = 32'd136314880;
      57857: inst = 32'd268468224;
      57858: inst = 32'd201348370;
      57859: inst = 32'd203423744;
      57860: inst = 32'd471859200;
      57861: inst = 32'd136314880;
      57862: inst = 32'd268468224;
      57863: inst = 32'd201348371;
      57864: inst = 32'd203423744;
      57865: inst = 32'd471859200;
      57866: inst = 32'd136314880;
      57867: inst = 32'd268468224;
      57868: inst = 32'd201348372;
      57869: inst = 32'd203423744;
      57870: inst = 32'd471859200;
      57871: inst = 32'd136314880;
      57872: inst = 32'd268468224;
      57873: inst = 32'd201348373;
      57874: inst = 32'd203423744;
      57875: inst = 32'd471859200;
      57876: inst = 32'd136314880;
      57877: inst = 32'd268468224;
      57878: inst = 32'd201348374;
      57879: inst = 32'd203423744;
      57880: inst = 32'd471859200;
      57881: inst = 32'd136314880;
      57882: inst = 32'd268468224;
      57883: inst = 32'd201348375;
      57884: inst = 32'd203423744;
      57885: inst = 32'd471859200;
      57886: inst = 32'd136314880;
      57887: inst = 32'd268468224;
      57888: inst = 32'd201348376;
      57889: inst = 32'd203423744;
      57890: inst = 32'd471859200;
      57891: inst = 32'd136314880;
      57892: inst = 32'd268468224;
      57893: inst = 32'd201348377;
      57894: inst = 32'd203423744;
      57895: inst = 32'd471859200;
      57896: inst = 32'd136314880;
      57897: inst = 32'd268468224;
      57898: inst = 32'd201348378;
      57899: inst = 32'd203423744;
      57900: inst = 32'd471859200;
      57901: inst = 32'd136314880;
      57902: inst = 32'd268468224;
      57903: inst = 32'd201348379;
      57904: inst = 32'd203423744;
      57905: inst = 32'd471859200;
      57906: inst = 32'd136314880;
      57907: inst = 32'd268468224;
      57908: inst = 32'd201348380;
      57909: inst = 32'd203423744;
      57910: inst = 32'd471859200;
      57911: inst = 32'd136314880;
      57912: inst = 32'd268468224;
      57913: inst = 32'd201348381;
      57914: inst = 32'd203423744;
      57915: inst = 32'd471859200;
      57916: inst = 32'd136314880;
      57917: inst = 32'd268468224;
      57918: inst = 32'd201348382;
      57919: inst = 32'd203423744;
      57920: inst = 32'd471859200;
      57921: inst = 32'd136314880;
      57922: inst = 32'd268468224;
      57923: inst = 32'd201348383;
      57924: inst = 32'd203423744;
      57925: inst = 32'd471859200;
      57926: inst = 32'd136314880;
      57927: inst = 32'd268468224;
      57928: inst = 32'd201348384;
      57929: inst = 32'd203423744;
      57930: inst = 32'd471859200;
      57931: inst = 32'd136314880;
      57932: inst = 32'd268468224;
      57933: inst = 32'd201348385;
      57934: inst = 32'd203423744;
      57935: inst = 32'd471859200;
      57936: inst = 32'd136314880;
      57937: inst = 32'd268468224;
      57938: inst = 32'd201348386;
      57939: inst = 32'd203423744;
      57940: inst = 32'd471859200;
      57941: inst = 32'd136314880;
      57942: inst = 32'd268468224;
      57943: inst = 32'd201348387;
      57944: inst = 32'd203423744;
      57945: inst = 32'd471859200;
      57946: inst = 32'd136314880;
      57947: inst = 32'd268468224;
      57948: inst = 32'd201348388;
      57949: inst = 32'd203423744;
      57950: inst = 32'd471859200;
      57951: inst = 32'd136314880;
      57952: inst = 32'd268468224;
      57953: inst = 32'd201348389;
      57954: inst = 32'd203423744;
      57955: inst = 32'd471859200;
      57956: inst = 32'd136314880;
      57957: inst = 32'd268468224;
      57958: inst = 32'd201348390;
      57959: inst = 32'd203423744;
      57960: inst = 32'd471859200;
      57961: inst = 32'd136314880;
      57962: inst = 32'd268468224;
      57963: inst = 32'd201348391;
      57964: inst = 32'd203423744;
      57965: inst = 32'd471859200;
      57966: inst = 32'd136314880;
      57967: inst = 32'd268468224;
      57968: inst = 32'd201348392;
      57969: inst = 32'd203423744;
      57970: inst = 32'd471859200;
      57971: inst = 32'd136314880;
      57972: inst = 32'd268468224;
      57973: inst = 32'd201348393;
      57974: inst = 32'd203423744;
      57975: inst = 32'd471859200;
      57976: inst = 32'd136314880;
      57977: inst = 32'd268468224;
      57978: inst = 32'd201348394;
      57979: inst = 32'd203423744;
      57980: inst = 32'd471859200;
      57981: inst = 32'd136314880;
      57982: inst = 32'd268468224;
      57983: inst = 32'd201348395;
      57984: inst = 32'd203423744;
      57985: inst = 32'd471859200;
      57986: inst = 32'd136314880;
      57987: inst = 32'd268468224;
      57988: inst = 32'd201348396;
      57989: inst = 32'd203423744;
      57990: inst = 32'd471859200;
      57991: inst = 32'd136314880;
      57992: inst = 32'd268468224;
      57993: inst = 32'd201348397;
      57994: inst = 32'd203423744;
      57995: inst = 32'd471859200;
      57996: inst = 32'd136314880;
      57997: inst = 32'd268468224;
      57998: inst = 32'd201348398;
      57999: inst = 32'd203423744;
      58000: inst = 32'd471859200;
      58001: inst = 32'd136314880;
      58002: inst = 32'd268468224;
      58003: inst = 32'd201348399;
      58004: inst = 32'd203423744;
      58005: inst = 32'd471859200;
      58006: inst = 32'd136314880;
      58007: inst = 32'd268468224;
      58008: inst = 32'd201348400;
      58009: inst = 32'd203423744;
      58010: inst = 32'd471859200;
      58011: inst = 32'd136314880;
      58012: inst = 32'd268468224;
      58013: inst = 32'd201348401;
      58014: inst = 32'd203423744;
      58015: inst = 32'd471859200;
      58016: inst = 32'd136314880;
      58017: inst = 32'd268468224;
      58018: inst = 32'd201348402;
      58019: inst = 32'd203423744;
      58020: inst = 32'd471859200;
      58021: inst = 32'd136314880;
      58022: inst = 32'd268468224;
      58023: inst = 32'd201348403;
      58024: inst = 32'd203423744;
      58025: inst = 32'd471859200;
      58026: inst = 32'd136314880;
      58027: inst = 32'd268468224;
      58028: inst = 32'd201348404;
      58029: inst = 32'd203423744;
      58030: inst = 32'd471859200;
      58031: inst = 32'd136314880;
      58032: inst = 32'd268468224;
      58033: inst = 32'd201348405;
      58034: inst = 32'd203423744;
      58035: inst = 32'd471859200;
      58036: inst = 32'd136314880;
      58037: inst = 32'd268468224;
      58038: inst = 32'd201348406;
      58039: inst = 32'd203423744;
      58040: inst = 32'd471859200;
      58041: inst = 32'd136314880;
      58042: inst = 32'd268468224;
      58043: inst = 32'd201348407;
      58044: inst = 32'd203423744;
      58045: inst = 32'd471859200;
      58046: inst = 32'd136314880;
      58047: inst = 32'd268468224;
      58048: inst = 32'd201348408;
      58049: inst = 32'd203423744;
      58050: inst = 32'd471859200;
      58051: inst = 32'd136314880;
      58052: inst = 32'd268468224;
      58053: inst = 32'd201348409;
      58054: inst = 32'd203423744;
      58055: inst = 32'd471859200;
      58056: inst = 32'd136314880;
      58057: inst = 32'd268468224;
      58058: inst = 32'd201348410;
      58059: inst = 32'd203423744;
      58060: inst = 32'd471859200;
      58061: inst = 32'd136314880;
      58062: inst = 32'd268468224;
      58063: inst = 32'd201348411;
      58064: inst = 32'd203423744;
      58065: inst = 32'd471859200;
      58066: inst = 32'd136314880;
      58067: inst = 32'd268468224;
      58068: inst = 32'd201348412;
      58069: inst = 32'd203423744;
      58070: inst = 32'd471859200;
      58071: inst = 32'd136314880;
      58072: inst = 32'd268468224;
      58073: inst = 32'd201348413;
      58074: inst = 32'd203423744;
      58075: inst = 32'd471859200;
      58076: inst = 32'd136314880;
      58077: inst = 32'd268468224;
      58078: inst = 32'd201348414;
      58079: inst = 32'd203423744;
      58080: inst = 32'd471859200;
      58081: inst = 32'd136314880;
      58082: inst = 32'd268468224;
      58083: inst = 32'd201348415;
      58084: inst = 32'd203423744;
      58085: inst = 32'd471859200;
      58086: inst = 32'd136314880;
      58087: inst = 32'd268468224;
      58088: inst = 32'd201348416;
      58089: inst = 32'd203423744;
      58090: inst = 32'd471859200;
      58091: inst = 32'd136314880;
      58092: inst = 32'd268468224;
      58093: inst = 32'd201348417;
      58094: inst = 32'd203423744;
      58095: inst = 32'd471859200;
      58096: inst = 32'd136314880;
      58097: inst = 32'd268468224;
      58098: inst = 32'd201348418;
      58099: inst = 32'd203423744;
      58100: inst = 32'd471859200;
      58101: inst = 32'd136314880;
      58102: inst = 32'd268468224;
      58103: inst = 32'd201348419;
      58104: inst = 32'd203423744;
      58105: inst = 32'd471859200;
      58106: inst = 32'd136314880;
      58107: inst = 32'd268468224;
      58108: inst = 32'd201348420;
      58109: inst = 32'd203423744;
      58110: inst = 32'd471859200;
      58111: inst = 32'd136314880;
      58112: inst = 32'd268468224;
      58113: inst = 32'd201348421;
      58114: inst = 32'd203423744;
      58115: inst = 32'd471859200;
      58116: inst = 32'd136314880;
      58117: inst = 32'd268468224;
      58118: inst = 32'd201348422;
      58119: inst = 32'd203423744;
      58120: inst = 32'd471859200;
      58121: inst = 32'd136314880;
      58122: inst = 32'd268468224;
      58123: inst = 32'd201348423;
      58124: inst = 32'd203423744;
      58125: inst = 32'd471859200;
      58126: inst = 32'd136314880;
      58127: inst = 32'd268468224;
      58128: inst = 32'd201348424;
      58129: inst = 32'd203423744;
      58130: inst = 32'd471859200;
      58131: inst = 32'd136314880;
      58132: inst = 32'd268468224;
      58133: inst = 32'd201348425;
      58134: inst = 32'd203423744;
      58135: inst = 32'd471859200;
      58136: inst = 32'd136314880;
      58137: inst = 32'd268468224;
      58138: inst = 32'd201348426;
      58139: inst = 32'd203423744;
      58140: inst = 32'd471859200;
      58141: inst = 32'd136314880;
      58142: inst = 32'd268468224;
      58143: inst = 32'd201348427;
      58144: inst = 32'd203423744;
      58145: inst = 32'd471859200;
      58146: inst = 32'd136314880;
      58147: inst = 32'd268468224;
      58148: inst = 32'd201348428;
      58149: inst = 32'd203423744;
      58150: inst = 32'd471859200;
      58151: inst = 32'd136314880;
      58152: inst = 32'd268468224;
      58153: inst = 32'd201348429;
      58154: inst = 32'd203423744;
      58155: inst = 32'd471859200;
      58156: inst = 32'd136314880;
      58157: inst = 32'd268468224;
      58158: inst = 32'd201348430;
      58159: inst = 32'd203423744;
      58160: inst = 32'd471859200;
      58161: inst = 32'd136314880;
      58162: inst = 32'd268468224;
      58163: inst = 32'd201348431;
      58164: inst = 32'd203423744;
      58165: inst = 32'd471859200;
      58166: inst = 32'd136314880;
      58167: inst = 32'd268468224;
      58168: inst = 32'd201348432;
      58169: inst = 32'd203423744;
      58170: inst = 32'd471859200;
      58171: inst = 32'd136314880;
      58172: inst = 32'd268468224;
      58173: inst = 32'd201348433;
      58174: inst = 32'd203423744;
      58175: inst = 32'd471859200;
      58176: inst = 32'd136314880;
      58177: inst = 32'd268468224;
      58178: inst = 32'd201348434;
      58179: inst = 32'd203423744;
      58180: inst = 32'd471859200;
      58181: inst = 32'd136314880;
      58182: inst = 32'd268468224;
      58183: inst = 32'd201348435;
      58184: inst = 32'd203423744;
      58185: inst = 32'd471859200;
      58186: inst = 32'd136314880;
      58187: inst = 32'd268468224;
      58188: inst = 32'd201348436;
      58189: inst = 32'd203423744;
      58190: inst = 32'd471859200;
      58191: inst = 32'd136314880;
      58192: inst = 32'd268468224;
      58193: inst = 32'd201348437;
      58194: inst = 32'd203423744;
      58195: inst = 32'd471859200;
      58196: inst = 32'd136314880;
      58197: inst = 32'd268468224;
      58198: inst = 32'd201348438;
      58199: inst = 32'd203423744;
      58200: inst = 32'd471859200;
      58201: inst = 32'd136314880;
      58202: inst = 32'd268468224;
      58203: inst = 32'd201348439;
      58204: inst = 32'd203423744;
      58205: inst = 32'd471859200;
      58206: inst = 32'd136314880;
      58207: inst = 32'd268468224;
      58208: inst = 32'd201348440;
      58209: inst = 32'd203423744;
      58210: inst = 32'd471859200;
      58211: inst = 32'd136314880;
      58212: inst = 32'd268468224;
      58213: inst = 32'd201348441;
      58214: inst = 32'd203423744;
      58215: inst = 32'd471859200;
      58216: inst = 32'd136314880;
      58217: inst = 32'd268468224;
      58218: inst = 32'd201348442;
      58219: inst = 32'd203423744;
      58220: inst = 32'd471859200;
      58221: inst = 32'd136314880;
      58222: inst = 32'd268468224;
      58223: inst = 32'd201348443;
      58224: inst = 32'd203423744;
      58225: inst = 32'd471859200;
      58226: inst = 32'd136314880;
      58227: inst = 32'd268468224;
      58228: inst = 32'd201348444;
      58229: inst = 32'd203423744;
      58230: inst = 32'd471859200;
      58231: inst = 32'd136314880;
      58232: inst = 32'd268468224;
      58233: inst = 32'd201348445;
      58234: inst = 32'd203423744;
      58235: inst = 32'd471859200;
      58236: inst = 32'd136314880;
      58237: inst = 32'd268468224;
      58238: inst = 32'd201348446;
      58239: inst = 32'd203423744;
      58240: inst = 32'd471859200;
      58241: inst = 32'd136314880;
      58242: inst = 32'd268468224;
      58243: inst = 32'd201348447;
      58244: inst = 32'd203423744;
      58245: inst = 32'd471859200;
      58246: inst = 32'd136314880;
      58247: inst = 32'd268468224;
      58248: inst = 32'd201348448;
      58249: inst = 32'd203423744;
      58250: inst = 32'd471859200;
      58251: inst = 32'd136314880;
      58252: inst = 32'd268468224;
      58253: inst = 32'd201348449;
      58254: inst = 32'd203423744;
      58255: inst = 32'd471859200;
      58256: inst = 32'd136314880;
      58257: inst = 32'd268468224;
      58258: inst = 32'd201348450;
      58259: inst = 32'd203423744;
      58260: inst = 32'd471859200;
      58261: inst = 32'd136314880;
      58262: inst = 32'd268468224;
      58263: inst = 32'd201348451;
      58264: inst = 32'd203423744;
      58265: inst = 32'd471859200;
      58266: inst = 32'd136314880;
      58267: inst = 32'd268468224;
      58268: inst = 32'd201348452;
      58269: inst = 32'd203423744;
      58270: inst = 32'd471859200;
      58271: inst = 32'd136314880;
      58272: inst = 32'd268468224;
      58273: inst = 32'd201348453;
      58274: inst = 32'd203423744;
      58275: inst = 32'd471859200;
      58276: inst = 32'd136314880;
      58277: inst = 32'd268468224;
      58278: inst = 32'd201348454;
      58279: inst = 32'd203423744;
      58280: inst = 32'd471859200;
      58281: inst = 32'd136314880;
      58282: inst = 32'd268468224;
      58283: inst = 32'd201348455;
      58284: inst = 32'd203423744;
      58285: inst = 32'd471859200;
      58286: inst = 32'd136314880;
      58287: inst = 32'd268468224;
      58288: inst = 32'd201348456;
      58289: inst = 32'd203423744;
      58290: inst = 32'd471859200;
      58291: inst = 32'd136314880;
      58292: inst = 32'd268468224;
      58293: inst = 32'd201348457;
      58294: inst = 32'd203423744;
      58295: inst = 32'd471859200;
      58296: inst = 32'd136314880;
      58297: inst = 32'd268468224;
      58298: inst = 32'd201348458;
      58299: inst = 32'd203423744;
      58300: inst = 32'd471859200;
      58301: inst = 32'd136314880;
      58302: inst = 32'd268468224;
      58303: inst = 32'd201348459;
      58304: inst = 32'd203423744;
      58305: inst = 32'd471859200;
      58306: inst = 32'd136314880;
      58307: inst = 32'd268468224;
      58308: inst = 32'd201348460;
      58309: inst = 32'd203423744;
      58310: inst = 32'd471859200;
      58311: inst = 32'd136314880;
      58312: inst = 32'd268468224;
      58313: inst = 32'd201348461;
      58314: inst = 32'd203423744;
      58315: inst = 32'd471859200;
      58316: inst = 32'd136314880;
      58317: inst = 32'd268468224;
      58318: inst = 32'd201348462;
      58319: inst = 32'd203423744;
      58320: inst = 32'd471859200;
      58321: inst = 32'd136314880;
      58322: inst = 32'd268468224;
      58323: inst = 32'd201348463;
      58324: inst = 32'd203423744;
      58325: inst = 32'd471859200;
      58326: inst = 32'd136314880;
      58327: inst = 32'd268468224;
      58328: inst = 32'd201348464;
      58329: inst = 32'd203423744;
      58330: inst = 32'd471859200;
      58331: inst = 32'd136314880;
      58332: inst = 32'd268468224;
      58333: inst = 32'd201348465;
      58334: inst = 32'd203423744;
      58335: inst = 32'd471859200;
      58336: inst = 32'd136314880;
      58337: inst = 32'd268468224;
      58338: inst = 32'd201348466;
      58339: inst = 32'd203423744;
      58340: inst = 32'd471859200;
      58341: inst = 32'd136314880;
      58342: inst = 32'd268468224;
      58343: inst = 32'd201348467;
      58344: inst = 32'd203423744;
      58345: inst = 32'd471859200;
      58346: inst = 32'd136314880;
      58347: inst = 32'd268468224;
      58348: inst = 32'd201348468;
      58349: inst = 32'd203423744;
      58350: inst = 32'd471859200;
      58351: inst = 32'd136314880;
      58352: inst = 32'd268468224;
      58353: inst = 32'd201348469;
      58354: inst = 32'd203423744;
      58355: inst = 32'd471859200;
      58356: inst = 32'd136314880;
      58357: inst = 32'd268468224;
      58358: inst = 32'd201348470;
      58359: inst = 32'd203423744;
      58360: inst = 32'd471859200;
      58361: inst = 32'd136314880;
      58362: inst = 32'd268468224;
      58363: inst = 32'd201348471;
      58364: inst = 32'd203423744;
      58365: inst = 32'd471859200;
      58366: inst = 32'd136314880;
      58367: inst = 32'd268468224;
      58368: inst = 32'd201348472;
      58369: inst = 32'd203423744;
      58370: inst = 32'd471859200;
      58371: inst = 32'd136314880;
      58372: inst = 32'd268468224;
      58373: inst = 32'd201348473;
      58374: inst = 32'd203423744;
      58375: inst = 32'd471859200;
      58376: inst = 32'd136314880;
      58377: inst = 32'd268468224;
      58378: inst = 32'd201348474;
      58379: inst = 32'd203423744;
      58380: inst = 32'd471859200;
      58381: inst = 32'd136314880;
      58382: inst = 32'd268468224;
      58383: inst = 32'd201348475;
      58384: inst = 32'd203423744;
      58385: inst = 32'd471859200;
      58386: inst = 32'd136314880;
      58387: inst = 32'd268468224;
      58388: inst = 32'd201348476;
      58389: inst = 32'd203423744;
      58390: inst = 32'd471859200;
      58391: inst = 32'd136314880;
      58392: inst = 32'd268468224;
      58393: inst = 32'd201348477;
      58394: inst = 32'd203423744;
      58395: inst = 32'd471859200;
      58396: inst = 32'd136314880;
      58397: inst = 32'd268468224;
      58398: inst = 32'd201348478;
      58399: inst = 32'd203423744;
      58400: inst = 32'd471859200;
      58401: inst = 32'd136314880;
      58402: inst = 32'd268468224;
      58403: inst = 32'd201348479;
      58404: inst = 32'd203423744;
      58405: inst = 32'd471859200;
      58406: inst = 32'd136314880;
      58407: inst = 32'd268468224;
      58408: inst = 32'd201348480;
      58409: inst = 32'd203423744;
      58410: inst = 32'd471859200;
      58411: inst = 32'd136314880;
      58412: inst = 32'd268468224;
      58413: inst = 32'd201348481;
      58414: inst = 32'd203423744;
      58415: inst = 32'd471859200;
      58416: inst = 32'd136314880;
      58417: inst = 32'd268468224;
      58418: inst = 32'd201348482;
      58419: inst = 32'd203423744;
      58420: inst = 32'd471859200;
      58421: inst = 32'd136314880;
      58422: inst = 32'd268468224;
      58423: inst = 32'd201348483;
      58424: inst = 32'd203423744;
      58425: inst = 32'd471859200;
      58426: inst = 32'd136314880;
      58427: inst = 32'd268468224;
      58428: inst = 32'd201348484;
      58429: inst = 32'd203423744;
      58430: inst = 32'd471859200;
      58431: inst = 32'd136314880;
      58432: inst = 32'd268468224;
      58433: inst = 32'd201348485;
      58434: inst = 32'd203423744;
      58435: inst = 32'd471859200;
      58436: inst = 32'd136314880;
      58437: inst = 32'd268468224;
      58438: inst = 32'd201348486;
      58439: inst = 32'd203423744;
      58440: inst = 32'd471859200;
      58441: inst = 32'd136314880;
      58442: inst = 32'd268468224;
      58443: inst = 32'd201348487;
      58444: inst = 32'd203423744;
      58445: inst = 32'd471859200;
      58446: inst = 32'd136314880;
      58447: inst = 32'd268468224;
      58448: inst = 32'd201348488;
      58449: inst = 32'd203423744;
      58450: inst = 32'd471859200;
      58451: inst = 32'd136314880;
      58452: inst = 32'd268468224;
      58453: inst = 32'd201348489;
      58454: inst = 32'd203423744;
      58455: inst = 32'd471859200;
      58456: inst = 32'd136314880;
      58457: inst = 32'd268468224;
      58458: inst = 32'd201348490;
      58459: inst = 32'd203423744;
      58460: inst = 32'd471859200;
      58461: inst = 32'd136314880;
      58462: inst = 32'd268468224;
      58463: inst = 32'd201348491;
      58464: inst = 32'd203423744;
      58465: inst = 32'd471859200;
      58466: inst = 32'd136314880;
      58467: inst = 32'd268468224;
      58468: inst = 32'd201348492;
      58469: inst = 32'd203423744;
      58470: inst = 32'd471859200;
      58471: inst = 32'd136314880;
      58472: inst = 32'd268468224;
      58473: inst = 32'd201348493;
      58474: inst = 32'd203423744;
      58475: inst = 32'd471859200;
      58476: inst = 32'd136314880;
      58477: inst = 32'd268468224;
      58478: inst = 32'd201348494;
      58479: inst = 32'd203423744;
      58480: inst = 32'd471859200;
      58481: inst = 32'd136314880;
      58482: inst = 32'd268468224;
      58483: inst = 32'd201348495;
      58484: inst = 32'd203423744;
      58485: inst = 32'd471859200;
      58486: inst = 32'd136314880;
      58487: inst = 32'd268468224;
      58488: inst = 32'd201348496;
      58489: inst = 32'd203423744;
      58490: inst = 32'd471859200;
      58491: inst = 32'd136314880;
      58492: inst = 32'd268468224;
      58493: inst = 32'd201348497;
      58494: inst = 32'd203423744;
      58495: inst = 32'd471859200;
      58496: inst = 32'd136314880;
      58497: inst = 32'd268468224;
      58498: inst = 32'd201348498;
      58499: inst = 32'd203423744;
      58500: inst = 32'd471859200;
      58501: inst = 32'd136314880;
      58502: inst = 32'd268468224;
      58503: inst = 32'd201348499;
      58504: inst = 32'd203423744;
      58505: inst = 32'd471859200;
      58506: inst = 32'd136314880;
      58507: inst = 32'd268468224;
      58508: inst = 32'd201348500;
      58509: inst = 32'd203423744;
      58510: inst = 32'd471859200;
      58511: inst = 32'd136314880;
      58512: inst = 32'd268468224;
      58513: inst = 32'd201348501;
      58514: inst = 32'd203423744;
      58515: inst = 32'd471859200;
      58516: inst = 32'd136314880;
      58517: inst = 32'd268468224;
      58518: inst = 32'd201348502;
      58519: inst = 32'd203423744;
      58520: inst = 32'd471859200;
      58521: inst = 32'd136314880;
      58522: inst = 32'd268468224;
      58523: inst = 32'd201348503;
      58524: inst = 32'd203423744;
      58525: inst = 32'd471859200;
      58526: inst = 32'd136314880;
      58527: inst = 32'd268468224;
      58528: inst = 32'd201348504;
      58529: inst = 32'd203423744;
      58530: inst = 32'd471859200;
      58531: inst = 32'd136314880;
      58532: inst = 32'd268468224;
      58533: inst = 32'd201348505;
      58534: inst = 32'd203423744;
      58535: inst = 32'd471859200;
      58536: inst = 32'd136314880;
      58537: inst = 32'd268468224;
      58538: inst = 32'd201348506;
      58539: inst = 32'd203423744;
      58540: inst = 32'd471859200;
      58541: inst = 32'd136314880;
      58542: inst = 32'd268468224;
      58543: inst = 32'd201348507;
      58544: inst = 32'd203423744;
      58545: inst = 32'd471859200;
      58546: inst = 32'd136314880;
      58547: inst = 32'd268468224;
      58548: inst = 32'd201348508;
      58549: inst = 32'd203423744;
      58550: inst = 32'd471859200;
      58551: inst = 32'd136314880;
      58552: inst = 32'd268468224;
      58553: inst = 32'd201348509;
      58554: inst = 32'd203423744;
      58555: inst = 32'd471859200;
      58556: inst = 32'd136314880;
      58557: inst = 32'd268468224;
      58558: inst = 32'd201348510;
      58559: inst = 32'd203423744;
      58560: inst = 32'd471859200;
      58561: inst = 32'd136314880;
      58562: inst = 32'd268468224;
      58563: inst = 32'd201348511;
      58564: inst = 32'd203423744;
      58565: inst = 32'd471859200;
      58566: inst = 32'd136314880;
      58567: inst = 32'd268468224;
      58568: inst = 32'd201348512;
      58569: inst = 32'd203423744;
      58570: inst = 32'd471859200;
      58571: inst = 32'd136314880;
      58572: inst = 32'd268468224;
      58573: inst = 32'd201348513;
      58574: inst = 32'd203423744;
      58575: inst = 32'd471859200;
      58576: inst = 32'd136314880;
      58577: inst = 32'd268468224;
      58578: inst = 32'd201348514;
      58579: inst = 32'd203423744;
      58580: inst = 32'd471859200;
      58581: inst = 32'd136314880;
      58582: inst = 32'd268468224;
      58583: inst = 32'd201348515;
      58584: inst = 32'd203423744;
      58585: inst = 32'd471859200;
      58586: inst = 32'd136314880;
      58587: inst = 32'd268468224;
      58588: inst = 32'd201348516;
      58589: inst = 32'd203423744;
      58590: inst = 32'd471859200;
      58591: inst = 32'd136314880;
      58592: inst = 32'd268468224;
      58593: inst = 32'd201348517;
      58594: inst = 32'd203423744;
      58595: inst = 32'd471859200;
      58596: inst = 32'd136314880;
      58597: inst = 32'd268468224;
      58598: inst = 32'd201348518;
      58599: inst = 32'd203423744;
      58600: inst = 32'd471859200;
      58601: inst = 32'd136314880;
      58602: inst = 32'd268468224;
      58603: inst = 32'd201348519;
      58604: inst = 32'd203423744;
      58605: inst = 32'd471859200;
      58606: inst = 32'd136314880;
      58607: inst = 32'd268468224;
      58608: inst = 32'd201348520;
      58609: inst = 32'd203423744;
      58610: inst = 32'd471859200;
      58611: inst = 32'd136314880;
      58612: inst = 32'd268468224;
      58613: inst = 32'd201348521;
      58614: inst = 32'd203423744;
      58615: inst = 32'd471859200;
      58616: inst = 32'd136314880;
      58617: inst = 32'd268468224;
      58618: inst = 32'd201348522;
      58619: inst = 32'd203423744;
      58620: inst = 32'd471859200;
      58621: inst = 32'd136314880;
      58622: inst = 32'd268468224;
      58623: inst = 32'd201348523;
      58624: inst = 32'd203423744;
      58625: inst = 32'd471859200;
      58626: inst = 32'd136314880;
      58627: inst = 32'd268468224;
      58628: inst = 32'd201348524;
      58629: inst = 32'd203423744;
      58630: inst = 32'd471859200;
      58631: inst = 32'd136314880;
      58632: inst = 32'd268468224;
      58633: inst = 32'd201348525;
      58634: inst = 32'd203423744;
      58635: inst = 32'd471859200;
      58636: inst = 32'd136314880;
      58637: inst = 32'd268468224;
      58638: inst = 32'd201348526;
      58639: inst = 32'd203423744;
      58640: inst = 32'd471859200;
      58641: inst = 32'd136314880;
      58642: inst = 32'd268468224;
      58643: inst = 32'd201348527;
      58644: inst = 32'd203423744;
      58645: inst = 32'd471859200;
      58646: inst = 32'd136314880;
      58647: inst = 32'd268468224;
      58648: inst = 32'd201348528;
      58649: inst = 32'd203423744;
      58650: inst = 32'd471859200;
      58651: inst = 32'd136314880;
      58652: inst = 32'd268468224;
      58653: inst = 32'd201348529;
      58654: inst = 32'd203423744;
      58655: inst = 32'd471859200;
      58656: inst = 32'd136314880;
      58657: inst = 32'd268468224;
      58658: inst = 32'd201348530;
      58659: inst = 32'd203423744;
      58660: inst = 32'd471859200;
      58661: inst = 32'd136314880;
      58662: inst = 32'd268468224;
      58663: inst = 32'd201348531;
      58664: inst = 32'd203423744;
      58665: inst = 32'd471859200;
      58666: inst = 32'd136314880;
      58667: inst = 32'd268468224;
      58668: inst = 32'd201348532;
      58669: inst = 32'd203423744;
      58670: inst = 32'd471859200;
      58671: inst = 32'd136314880;
      58672: inst = 32'd268468224;
      58673: inst = 32'd201348533;
      58674: inst = 32'd203423744;
      58675: inst = 32'd471859200;
      58676: inst = 32'd136314880;
      58677: inst = 32'd268468224;
      58678: inst = 32'd201348534;
      58679: inst = 32'd203423744;
      58680: inst = 32'd471859200;
      58681: inst = 32'd136314880;
      58682: inst = 32'd268468224;
      58683: inst = 32'd201348535;
      58684: inst = 32'd203423744;
      58685: inst = 32'd471859200;
      58686: inst = 32'd136314880;
      58687: inst = 32'd268468224;
      58688: inst = 32'd201348536;
      58689: inst = 32'd203423744;
      58690: inst = 32'd471859200;
      58691: inst = 32'd136314880;
      58692: inst = 32'd268468224;
      58693: inst = 32'd201348537;
      58694: inst = 32'd203423744;
      58695: inst = 32'd471859200;
      58696: inst = 32'd136314880;
      58697: inst = 32'd268468224;
      58698: inst = 32'd201348538;
      58699: inst = 32'd203423744;
      58700: inst = 32'd471859200;
      58701: inst = 32'd136314880;
      58702: inst = 32'd268468224;
      58703: inst = 32'd201348539;
      58704: inst = 32'd203423744;
      58705: inst = 32'd471859200;
      58706: inst = 32'd136314880;
      58707: inst = 32'd268468224;
      58708: inst = 32'd201348540;
      58709: inst = 32'd203423744;
      58710: inst = 32'd471859200;
      58711: inst = 32'd136314880;
      58712: inst = 32'd268468224;
      58713: inst = 32'd201348541;
      58714: inst = 32'd203423744;
      58715: inst = 32'd471859200;
      58716: inst = 32'd136314880;
      58717: inst = 32'd268468224;
      58718: inst = 32'd201348542;
      58719: inst = 32'd203423744;
      58720: inst = 32'd471859200;
      58721: inst = 32'd136314880;
      58722: inst = 32'd268468224;
      58723: inst = 32'd201348543;
      58724: inst = 32'd203423744;
      58725: inst = 32'd471859200;
      58726: inst = 32'd136314880;
      58727: inst = 32'd268468224;
      58728: inst = 32'd201348544;
      58729: inst = 32'd203423744;
      58730: inst = 32'd471859200;
      58731: inst = 32'd136314880;
      58732: inst = 32'd268468224;
      58733: inst = 32'd201348545;
      58734: inst = 32'd203423744;
      58735: inst = 32'd471859200;
      58736: inst = 32'd136314880;
      58737: inst = 32'd268468224;
      58738: inst = 32'd201348546;
      58739: inst = 32'd203423744;
      58740: inst = 32'd471859200;
      58741: inst = 32'd136314880;
      58742: inst = 32'd268468224;
      58743: inst = 32'd201348547;
      58744: inst = 32'd203423744;
      58745: inst = 32'd471859200;
      58746: inst = 32'd136314880;
      58747: inst = 32'd268468224;
      58748: inst = 32'd201348548;
      58749: inst = 32'd203423744;
      58750: inst = 32'd471859200;
      58751: inst = 32'd136314880;
      58752: inst = 32'd268468224;
      58753: inst = 32'd201348549;
      58754: inst = 32'd203423744;
      58755: inst = 32'd471859200;
      58756: inst = 32'd136314880;
      58757: inst = 32'd268468224;
      58758: inst = 32'd201348550;
      58759: inst = 32'd203423744;
      58760: inst = 32'd471859200;
      58761: inst = 32'd136314880;
      58762: inst = 32'd268468224;
      58763: inst = 32'd201348551;
      58764: inst = 32'd203423744;
      58765: inst = 32'd471859200;
      58766: inst = 32'd136314880;
      58767: inst = 32'd268468224;
      58768: inst = 32'd201348552;
      58769: inst = 32'd203423744;
      58770: inst = 32'd471859200;
      58771: inst = 32'd136314880;
      58772: inst = 32'd268468224;
      58773: inst = 32'd201348553;
      58774: inst = 32'd203423744;
      58775: inst = 32'd471859200;
      58776: inst = 32'd136314880;
      58777: inst = 32'd268468224;
      58778: inst = 32'd201348554;
      58779: inst = 32'd203423744;
      58780: inst = 32'd471859200;
      58781: inst = 32'd136314880;
      58782: inst = 32'd268468224;
      58783: inst = 32'd201348555;
      58784: inst = 32'd203423744;
      58785: inst = 32'd471859200;
      58786: inst = 32'd136314880;
      58787: inst = 32'd268468224;
      58788: inst = 32'd201348556;
      58789: inst = 32'd203423744;
      58790: inst = 32'd471859200;
      58791: inst = 32'd136314880;
      58792: inst = 32'd268468224;
      58793: inst = 32'd201348557;
      58794: inst = 32'd203423744;
      58795: inst = 32'd471859200;
      58796: inst = 32'd136314880;
      58797: inst = 32'd268468224;
      58798: inst = 32'd201348558;
      58799: inst = 32'd203423744;
      58800: inst = 32'd471859200;
      58801: inst = 32'd136314880;
      58802: inst = 32'd268468224;
      58803: inst = 32'd201348559;
      58804: inst = 32'd203423744;
      58805: inst = 32'd471859200;
      58806: inst = 32'd136314880;
      58807: inst = 32'd268468224;
      58808: inst = 32'd201348560;
      58809: inst = 32'd203423744;
      58810: inst = 32'd471859200;
      58811: inst = 32'd136314880;
      58812: inst = 32'd268468224;
      58813: inst = 32'd201348561;
      58814: inst = 32'd203423744;
      58815: inst = 32'd471859200;
      58816: inst = 32'd136314880;
      58817: inst = 32'd268468224;
      58818: inst = 32'd201348562;
      58819: inst = 32'd203423744;
      58820: inst = 32'd471859200;
      58821: inst = 32'd136314880;
      58822: inst = 32'd268468224;
      58823: inst = 32'd201348563;
      58824: inst = 32'd203423744;
      58825: inst = 32'd471859200;
      58826: inst = 32'd136314880;
      58827: inst = 32'd268468224;
      58828: inst = 32'd201348564;
      58829: inst = 32'd203423744;
      58830: inst = 32'd471859200;
      58831: inst = 32'd136314880;
      58832: inst = 32'd268468224;
      58833: inst = 32'd201348565;
      58834: inst = 32'd203423744;
      58835: inst = 32'd471859200;
      58836: inst = 32'd136314880;
      58837: inst = 32'd268468224;
      58838: inst = 32'd201348566;
      58839: inst = 32'd203423744;
      58840: inst = 32'd471859200;
      58841: inst = 32'd136314880;
      58842: inst = 32'd268468224;
      58843: inst = 32'd201348567;
      58844: inst = 32'd203423744;
      58845: inst = 32'd471859200;
      58846: inst = 32'd136314880;
      58847: inst = 32'd268468224;
      58848: inst = 32'd201348568;
      58849: inst = 32'd203423744;
      58850: inst = 32'd471859200;
      58851: inst = 32'd136314880;
      58852: inst = 32'd268468224;
      58853: inst = 32'd201348569;
      58854: inst = 32'd203423744;
      58855: inst = 32'd471859200;
      58856: inst = 32'd136314880;
      58857: inst = 32'd268468224;
      58858: inst = 32'd201348570;
      58859: inst = 32'd203423744;
      58860: inst = 32'd471859200;
      58861: inst = 32'd136314880;
      58862: inst = 32'd268468224;
      58863: inst = 32'd201348571;
      58864: inst = 32'd203423744;
      58865: inst = 32'd471859200;
      58866: inst = 32'd136314880;
      58867: inst = 32'd268468224;
      58868: inst = 32'd201348572;
      58869: inst = 32'd203423744;
      58870: inst = 32'd471859200;
      58871: inst = 32'd136314880;
      58872: inst = 32'd268468224;
      58873: inst = 32'd201348573;
      58874: inst = 32'd203423744;
      58875: inst = 32'd471859200;
      58876: inst = 32'd136314880;
      58877: inst = 32'd268468224;
      58878: inst = 32'd201348574;
      58879: inst = 32'd203423744;
      58880: inst = 32'd471859200;
      58881: inst = 32'd136314880;
      58882: inst = 32'd268468224;
      58883: inst = 32'd201348575;
      58884: inst = 32'd203423744;
      58885: inst = 32'd471859200;
      58886: inst = 32'd136314880;
      58887: inst = 32'd268468224;
      58888: inst = 32'd201348576;
      58889: inst = 32'd203423744;
      58890: inst = 32'd471859200;
      58891: inst = 32'd136314880;
      58892: inst = 32'd268468224;
      58893: inst = 32'd201348577;
      58894: inst = 32'd203423744;
      58895: inst = 32'd471859200;
      58896: inst = 32'd136314880;
      58897: inst = 32'd268468224;
      58898: inst = 32'd201348578;
      58899: inst = 32'd203423744;
      58900: inst = 32'd471859200;
      58901: inst = 32'd136314880;
      58902: inst = 32'd268468224;
      58903: inst = 32'd201348579;
      58904: inst = 32'd203423744;
      58905: inst = 32'd471859200;
      58906: inst = 32'd136314880;
      58907: inst = 32'd268468224;
      58908: inst = 32'd201348580;
      58909: inst = 32'd203423744;
      58910: inst = 32'd471859200;
      58911: inst = 32'd136314880;
      58912: inst = 32'd268468224;
      58913: inst = 32'd201348581;
      58914: inst = 32'd203423744;
      58915: inst = 32'd471859200;
      58916: inst = 32'd136314880;
      58917: inst = 32'd268468224;
      58918: inst = 32'd201348582;
      58919: inst = 32'd203423744;
      58920: inst = 32'd471859200;
      58921: inst = 32'd136314880;
      58922: inst = 32'd268468224;
      58923: inst = 32'd201348583;
      58924: inst = 32'd203423744;
      58925: inst = 32'd471859200;
      58926: inst = 32'd136314880;
      58927: inst = 32'd268468224;
      58928: inst = 32'd201348584;
      58929: inst = 32'd203423744;
      58930: inst = 32'd471859200;
      58931: inst = 32'd136314880;
      58932: inst = 32'd268468224;
      58933: inst = 32'd201348585;
      58934: inst = 32'd203423744;
      58935: inst = 32'd471859200;
      58936: inst = 32'd136314880;
      58937: inst = 32'd268468224;
      58938: inst = 32'd201348586;
      58939: inst = 32'd203423744;
      58940: inst = 32'd471859200;
      58941: inst = 32'd136314880;
      58942: inst = 32'd268468224;
      58943: inst = 32'd201348587;
      58944: inst = 32'd203423744;
      58945: inst = 32'd471859200;
      58946: inst = 32'd136314880;
      58947: inst = 32'd268468224;
      58948: inst = 32'd201348588;
      58949: inst = 32'd203423744;
      58950: inst = 32'd471859200;
      58951: inst = 32'd136314880;
      58952: inst = 32'd268468224;
      58953: inst = 32'd201348589;
      58954: inst = 32'd203423744;
      58955: inst = 32'd471859200;
      58956: inst = 32'd136314880;
      58957: inst = 32'd268468224;
      58958: inst = 32'd201348590;
      58959: inst = 32'd203423744;
      58960: inst = 32'd471859200;
      58961: inst = 32'd136314880;
      58962: inst = 32'd268468224;
      58963: inst = 32'd201348591;
      58964: inst = 32'd203423744;
      58965: inst = 32'd471859200;
      58966: inst = 32'd136314880;
      58967: inst = 32'd268468224;
      58968: inst = 32'd201348592;
      58969: inst = 32'd203423744;
      58970: inst = 32'd471859200;
      58971: inst = 32'd136314880;
      58972: inst = 32'd268468224;
      58973: inst = 32'd201348593;
      58974: inst = 32'd203423744;
      58975: inst = 32'd471859200;
      58976: inst = 32'd136314880;
      58977: inst = 32'd268468224;
      58978: inst = 32'd201348594;
      58979: inst = 32'd203423744;
      58980: inst = 32'd471859200;
      58981: inst = 32'd136314880;
      58982: inst = 32'd268468224;
      58983: inst = 32'd201348595;
      58984: inst = 32'd203423744;
      58985: inst = 32'd471859200;
      58986: inst = 32'd136314880;
      58987: inst = 32'd268468224;
      58988: inst = 32'd201348596;
      58989: inst = 32'd203423744;
      58990: inst = 32'd471859200;
      58991: inst = 32'd136314880;
      58992: inst = 32'd268468224;
      58993: inst = 32'd201348597;
      58994: inst = 32'd203423744;
      58995: inst = 32'd471859200;
      58996: inst = 32'd136314880;
      58997: inst = 32'd268468224;
      58998: inst = 32'd201348598;
      58999: inst = 32'd203423744;
      59000: inst = 32'd471859200;
      59001: inst = 32'd136314880;
      59002: inst = 32'd268468224;
      59003: inst = 32'd201348599;
      59004: inst = 32'd203423744;
      59005: inst = 32'd471859200;
      59006: inst = 32'd136314880;
      59007: inst = 32'd268468224;
      59008: inst = 32'd201348600;
      59009: inst = 32'd203423744;
      59010: inst = 32'd471859200;
      59011: inst = 32'd136314880;
      59012: inst = 32'd268468224;
      59013: inst = 32'd201348601;
      59014: inst = 32'd203423744;
      59015: inst = 32'd471859200;
      59016: inst = 32'd136314880;
      59017: inst = 32'd268468224;
      59018: inst = 32'd201348602;
      59019: inst = 32'd203423744;
      59020: inst = 32'd471859200;
      59021: inst = 32'd136314880;
      59022: inst = 32'd268468224;
      59023: inst = 32'd201348603;
      59024: inst = 32'd203423744;
      59025: inst = 32'd471859200;
      59026: inst = 32'd136314880;
      59027: inst = 32'd268468224;
      59028: inst = 32'd201348604;
      59029: inst = 32'd203423744;
      59030: inst = 32'd471859200;
      59031: inst = 32'd136314880;
      59032: inst = 32'd268468224;
      59033: inst = 32'd201348605;
      59034: inst = 32'd203423744;
      59035: inst = 32'd471859200;
      59036: inst = 32'd136314880;
      59037: inst = 32'd268468224;
      59038: inst = 32'd201348606;
      59039: inst = 32'd203423744;
      59040: inst = 32'd471859200;
      59041: inst = 32'd136314880;
      59042: inst = 32'd268468224;
      59043: inst = 32'd201348607;
      59044: inst = 32'd203423744;
      59045: inst = 32'd471859200;
      59046: inst = 32'd136314880;
      59047: inst = 32'd268468224;
      59048: inst = 32'd201348608;
      59049: inst = 32'd203423744;
      59050: inst = 32'd471859200;
      59051: inst = 32'd136314880;
      59052: inst = 32'd268468224;
      59053: inst = 32'd201348609;
      59054: inst = 32'd203423744;
      59055: inst = 32'd471859200;
      59056: inst = 32'd136314880;
      59057: inst = 32'd268468224;
      59058: inst = 32'd201348610;
      59059: inst = 32'd203423744;
      59060: inst = 32'd471859200;
      59061: inst = 32'd136314880;
      59062: inst = 32'd268468224;
      59063: inst = 32'd201348611;
      59064: inst = 32'd203423744;
      59065: inst = 32'd471859200;
      59066: inst = 32'd136314880;
      59067: inst = 32'd268468224;
      59068: inst = 32'd201348612;
      59069: inst = 32'd203423744;
      59070: inst = 32'd471859200;
      59071: inst = 32'd136314880;
      59072: inst = 32'd268468224;
      59073: inst = 32'd201348613;
      59074: inst = 32'd203423744;
      59075: inst = 32'd471859200;
      59076: inst = 32'd136314880;
      59077: inst = 32'd268468224;
      59078: inst = 32'd201348614;
      59079: inst = 32'd203423744;
      59080: inst = 32'd471859200;
      59081: inst = 32'd136314880;
      59082: inst = 32'd268468224;
      59083: inst = 32'd201348615;
      59084: inst = 32'd203423744;
      59085: inst = 32'd471859200;
      59086: inst = 32'd136314880;
      59087: inst = 32'd268468224;
      59088: inst = 32'd201348616;
      59089: inst = 32'd203423744;
      59090: inst = 32'd471859200;
      59091: inst = 32'd136314880;
      59092: inst = 32'd268468224;
      59093: inst = 32'd201348617;
      59094: inst = 32'd203423744;
      59095: inst = 32'd471859200;
      59096: inst = 32'd136314880;
      59097: inst = 32'd268468224;
      59098: inst = 32'd201348618;
      59099: inst = 32'd203423744;
      59100: inst = 32'd471859200;
      59101: inst = 32'd136314880;
      59102: inst = 32'd268468224;
      59103: inst = 32'd201348619;
      59104: inst = 32'd203423744;
      59105: inst = 32'd471859200;
      59106: inst = 32'd136314880;
      59107: inst = 32'd268468224;
      59108: inst = 32'd201348620;
      59109: inst = 32'd203423744;
      59110: inst = 32'd471859200;
      59111: inst = 32'd136314880;
      59112: inst = 32'd268468224;
      59113: inst = 32'd201348621;
      59114: inst = 32'd203423744;
      59115: inst = 32'd471859200;
      59116: inst = 32'd136314880;
      59117: inst = 32'd268468224;
      59118: inst = 32'd201348622;
      59119: inst = 32'd203423744;
      59120: inst = 32'd471859200;
      59121: inst = 32'd136314880;
      59122: inst = 32'd268468224;
      59123: inst = 32'd201348623;
      59124: inst = 32'd203423744;
      59125: inst = 32'd471859200;
      59126: inst = 32'd136314880;
      59127: inst = 32'd268468224;
      59128: inst = 32'd201348624;
      59129: inst = 32'd203423744;
      59130: inst = 32'd471859200;
      59131: inst = 32'd136314880;
      59132: inst = 32'd268468224;
      59133: inst = 32'd201348625;
      59134: inst = 32'd203423744;
      59135: inst = 32'd471859200;
      59136: inst = 32'd136314880;
      59137: inst = 32'd268468224;
      59138: inst = 32'd201348626;
      59139: inst = 32'd203423744;
      59140: inst = 32'd471859200;
      59141: inst = 32'd136314880;
      59142: inst = 32'd268468224;
      59143: inst = 32'd201348627;
      59144: inst = 32'd203423744;
      59145: inst = 32'd471859200;
      59146: inst = 32'd136314880;
      59147: inst = 32'd268468224;
      59148: inst = 32'd201348628;
      59149: inst = 32'd203423744;
      59150: inst = 32'd471859200;
      59151: inst = 32'd136314880;
      59152: inst = 32'd268468224;
      59153: inst = 32'd201348629;
      59154: inst = 32'd203423744;
      59155: inst = 32'd471859200;
      59156: inst = 32'd136314880;
      59157: inst = 32'd268468224;
      59158: inst = 32'd201348630;
      59159: inst = 32'd203423744;
      59160: inst = 32'd471859200;
      59161: inst = 32'd136314880;
      59162: inst = 32'd268468224;
      59163: inst = 32'd201348631;
      59164: inst = 32'd203423744;
      59165: inst = 32'd471859200;
      59166: inst = 32'd136314880;
      59167: inst = 32'd268468224;
      59168: inst = 32'd201348632;
      59169: inst = 32'd203423744;
      59170: inst = 32'd471859200;
      59171: inst = 32'd136314880;
      59172: inst = 32'd268468224;
      59173: inst = 32'd201348633;
      59174: inst = 32'd203423744;
      59175: inst = 32'd471859200;
      59176: inst = 32'd136314880;
      59177: inst = 32'd268468224;
      59178: inst = 32'd201348634;
      59179: inst = 32'd203423744;
      59180: inst = 32'd471859200;
      59181: inst = 32'd136314880;
      59182: inst = 32'd268468224;
      59183: inst = 32'd201348635;
      59184: inst = 32'd203423744;
      59185: inst = 32'd471859200;
      59186: inst = 32'd136314880;
      59187: inst = 32'd268468224;
      59188: inst = 32'd201348636;
      59189: inst = 32'd203423744;
      59190: inst = 32'd471859200;
      59191: inst = 32'd136314880;
      59192: inst = 32'd268468224;
      59193: inst = 32'd201348637;
      59194: inst = 32'd203423744;
      59195: inst = 32'd471859200;
      59196: inst = 32'd136314880;
      59197: inst = 32'd268468224;
      59198: inst = 32'd201348638;
      59199: inst = 32'd203423744;
      59200: inst = 32'd471859200;
      59201: inst = 32'd136314880;
      59202: inst = 32'd268468224;
      59203: inst = 32'd201348639;
      59204: inst = 32'd203423744;
      59205: inst = 32'd471859200;
      59206: inst = 32'd136314880;
      59207: inst = 32'd268468224;
      59208: inst = 32'd201348640;
      59209: inst = 32'd203423744;
      59210: inst = 32'd471859200;
      59211: inst = 32'd136314880;
      59212: inst = 32'd268468224;
      59213: inst = 32'd201348641;
      59214: inst = 32'd203423744;
      59215: inst = 32'd471859200;
      59216: inst = 32'd136314880;
      59217: inst = 32'd268468224;
      59218: inst = 32'd201348642;
      59219: inst = 32'd203423744;
      59220: inst = 32'd471859200;
      59221: inst = 32'd136314880;
      59222: inst = 32'd268468224;
      59223: inst = 32'd201348643;
      59224: inst = 32'd203423744;
      59225: inst = 32'd471859200;
      59226: inst = 32'd136314880;
      59227: inst = 32'd268468224;
      59228: inst = 32'd201348644;
      59229: inst = 32'd203423744;
      59230: inst = 32'd471859200;
      59231: inst = 32'd136314880;
      59232: inst = 32'd268468224;
      59233: inst = 32'd201348645;
      59234: inst = 32'd203423744;
      59235: inst = 32'd471859200;
      59236: inst = 32'd136314880;
      59237: inst = 32'd268468224;
      59238: inst = 32'd201348646;
      59239: inst = 32'd203423744;
      59240: inst = 32'd471859200;
      59241: inst = 32'd136314880;
      59242: inst = 32'd268468224;
      59243: inst = 32'd201348647;
      59244: inst = 32'd203423744;
      59245: inst = 32'd471859200;
      59246: inst = 32'd136314880;
      59247: inst = 32'd268468224;
      59248: inst = 32'd201348648;
      59249: inst = 32'd203423744;
      59250: inst = 32'd471859200;
      59251: inst = 32'd136314880;
      59252: inst = 32'd268468224;
      59253: inst = 32'd201348649;
      59254: inst = 32'd203423744;
      59255: inst = 32'd471859200;
      59256: inst = 32'd136314880;
      59257: inst = 32'd268468224;
      59258: inst = 32'd201348650;
      59259: inst = 32'd203423744;
      59260: inst = 32'd471859200;
      59261: inst = 32'd136314880;
      59262: inst = 32'd268468224;
      59263: inst = 32'd201348651;
      59264: inst = 32'd203423744;
      59265: inst = 32'd471859200;
      59266: inst = 32'd136314880;
      59267: inst = 32'd268468224;
      59268: inst = 32'd201348652;
      59269: inst = 32'd203423744;
      59270: inst = 32'd471859200;
      59271: inst = 32'd136314880;
      59272: inst = 32'd268468224;
      59273: inst = 32'd201348653;
      59274: inst = 32'd203423744;
      59275: inst = 32'd471859200;
      59276: inst = 32'd136314880;
      59277: inst = 32'd268468224;
      59278: inst = 32'd201348654;
      59279: inst = 32'd203423744;
      59280: inst = 32'd471859200;
      59281: inst = 32'd136314880;
      59282: inst = 32'd268468224;
      59283: inst = 32'd201348655;
      59284: inst = 32'd203423744;
      59285: inst = 32'd471859200;
      59286: inst = 32'd136314880;
      59287: inst = 32'd268468224;
      59288: inst = 32'd201348656;
      59289: inst = 32'd203423744;
      59290: inst = 32'd471859200;
      59291: inst = 32'd136314880;
      59292: inst = 32'd268468224;
      59293: inst = 32'd201348657;
      59294: inst = 32'd203423744;
      59295: inst = 32'd471859200;
      59296: inst = 32'd136314880;
      59297: inst = 32'd268468224;
      59298: inst = 32'd201348658;
      59299: inst = 32'd203423744;
      59300: inst = 32'd471859200;
      59301: inst = 32'd136314880;
      59302: inst = 32'd268468224;
      59303: inst = 32'd201348659;
      59304: inst = 32'd203423744;
      59305: inst = 32'd471859200;
      59306: inst = 32'd136314880;
      59307: inst = 32'd268468224;
      59308: inst = 32'd201348660;
      59309: inst = 32'd203423744;
      59310: inst = 32'd471859200;
      59311: inst = 32'd136314880;
      59312: inst = 32'd268468224;
      59313: inst = 32'd201348661;
      59314: inst = 32'd203423744;
      59315: inst = 32'd471859200;
      59316: inst = 32'd136314880;
      59317: inst = 32'd268468224;
      59318: inst = 32'd201348662;
      59319: inst = 32'd203423744;
      59320: inst = 32'd471859200;
      59321: inst = 32'd136314880;
      59322: inst = 32'd268468224;
      59323: inst = 32'd201348663;
      59324: inst = 32'd203423744;
      59325: inst = 32'd471859200;
      59326: inst = 32'd136314880;
      59327: inst = 32'd268468224;
      59328: inst = 32'd201348664;
      59329: inst = 32'd203423744;
      59330: inst = 32'd471859200;
      59331: inst = 32'd136314880;
      59332: inst = 32'd268468224;
      59333: inst = 32'd201348665;
      59334: inst = 32'd203423744;
      59335: inst = 32'd471859200;
      59336: inst = 32'd136314880;
      59337: inst = 32'd268468224;
      59338: inst = 32'd201348666;
      59339: inst = 32'd203423744;
      59340: inst = 32'd471859200;
      59341: inst = 32'd136314880;
      59342: inst = 32'd268468224;
      59343: inst = 32'd201348667;
      59344: inst = 32'd203423744;
      59345: inst = 32'd471859200;
      59346: inst = 32'd136314880;
      59347: inst = 32'd268468224;
      59348: inst = 32'd201348668;
      59349: inst = 32'd203423744;
      59350: inst = 32'd471859200;
      59351: inst = 32'd136314880;
      59352: inst = 32'd268468224;
      59353: inst = 32'd201348669;
      59354: inst = 32'd203423744;
      59355: inst = 32'd471859200;
      59356: inst = 32'd136314880;
      59357: inst = 32'd268468224;
      59358: inst = 32'd201348670;
      59359: inst = 32'd203423744;
      59360: inst = 32'd471859200;
      59361: inst = 32'd136314880;
      59362: inst = 32'd268468224;
      59363: inst = 32'd201348671;
      59364: inst = 32'd203423744;
      59365: inst = 32'd471859200;
      59366: inst = 32'd136314880;
      59367: inst = 32'd268468224;
      59368: inst = 32'd201348672;
      59369: inst = 32'd203423744;
      59370: inst = 32'd471859200;
      59371: inst = 32'd136314880;
      59372: inst = 32'd268468224;
      59373: inst = 32'd201348673;
      59374: inst = 32'd203423744;
      59375: inst = 32'd471859200;
      59376: inst = 32'd136314880;
      59377: inst = 32'd268468224;
      59378: inst = 32'd201348674;
      59379: inst = 32'd203423744;
      59380: inst = 32'd471859200;
      59381: inst = 32'd136314880;
      59382: inst = 32'd268468224;
      59383: inst = 32'd201348675;
      59384: inst = 32'd203423744;
      59385: inst = 32'd471859200;
      59386: inst = 32'd136314880;
      59387: inst = 32'd268468224;
      59388: inst = 32'd201348676;
      59389: inst = 32'd203423744;
      59390: inst = 32'd471859200;
      59391: inst = 32'd136314880;
      59392: inst = 32'd268468224;
      59393: inst = 32'd201348677;
      59394: inst = 32'd203423744;
      59395: inst = 32'd471859200;
      59396: inst = 32'd136314880;
      59397: inst = 32'd268468224;
      59398: inst = 32'd201348678;
      59399: inst = 32'd203423744;
      59400: inst = 32'd471859200;
      59401: inst = 32'd136314880;
      59402: inst = 32'd268468224;
      59403: inst = 32'd201348679;
      59404: inst = 32'd203423744;
      59405: inst = 32'd471859200;
      59406: inst = 32'd136314880;
      59407: inst = 32'd268468224;
      59408: inst = 32'd201348680;
      59409: inst = 32'd203423744;
      59410: inst = 32'd471859200;
      59411: inst = 32'd136314880;
      59412: inst = 32'd268468224;
      59413: inst = 32'd201348681;
      59414: inst = 32'd203423744;
      59415: inst = 32'd471859200;
      59416: inst = 32'd136314880;
      59417: inst = 32'd268468224;
      59418: inst = 32'd201348682;
      59419: inst = 32'd203423744;
      59420: inst = 32'd471859200;
      59421: inst = 32'd136314880;
      59422: inst = 32'd268468224;
      59423: inst = 32'd201348683;
      59424: inst = 32'd203423744;
      59425: inst = 32'd471859200;
      59426: inst = 32'd136314880;
      59427: inst = 32'd268468224;
      59428: inst = 32'd201348684;
      59429: inst = 32'd203423744;
      59430: inst = 32'd471859200;
      59431: inst = 32'd136314880;
      59432: inst = 32'd268468224;
      59433: inst = 32'd201348685;
      59434: inst = 32'd203423744;
      59435: inst = 32'd471859200;
      59436: inst = 32'd136314880;
      59437: inst = 32'd268468224;
      59438: inst = 32'd201348686;
      59439: inst = 32'd203423744;
      59440: inst = 32'd471859200;
      59441: inst = 32'd136314880;
      59442: inst = 32'd268468224;
      59443: inst = 32'd201348687;
      59444: inst = 32'd203423744;
      59445: inst = 32'd471859200;
      59446: inst = 32'd136314880;
      59447: inst = 32'd268468224;
      59448: inst = 32'd201348688;
      59449: inst = 32'd203423744;
      59450: inst = 32'd471859200;
      59451: inst = 32'd136314880;
      59452: inst = 32'd268468224;
      59453: inst = 32'd201348689;
      59454: inst = 32'd203423744;
      59455: inst = 32'd471859200;
      59456: inst = 32'd136314880;
      59457: inst = 32'd268468224;
      59458: inst = 32'd201348690;
      59459: inst = 32'd203423744;
      59460: inst = 32'd471859200;
      59461: inst = 32'd136314880;
      59462: inst = 32'd268468224;
      59463: inst = 32'd201348691;
      59464: inst = 32'd203423744;
      59465: inst = 32'd471859200;
      59466: inst = 32'd136314880;
      59467: inst = 32'd268468224;
      59468: inst = 32'd201348692;
      59469: inst = 32'd203423744;
      59470: inst = 32'd471859200;
      59471: inst = 32'd136314880;
      59472: inst = 32'd268468224;
      59473: inst = 32'd201348693;
      59474: inst = 32'd203423744;
      59475: inst = 32'd471859200;
      59476: inst = 32'd136314880;
      59477: inst = 32'd268468224;
      59478: inst = 32'd201348694;
      59479: inst = 32'd203423744;
      59480: inst = 32'd471859200;
      59481: inst = 32'd136314880;
      59482: inst = 32'd268468224;
      59483: inst = 32'd201348695;
      59484: inst = 32'd203423744;
      59485: inst = 32'd471859200;
      59486: inst = 32'd136314880;
      59487: inst = 32'd268468224;
      59488: inst = 32'd201348696;
      59489: inst = 32'd203423744;
      59490: inst = 32'd471859200;
      59491: inst = 32'd136314880;
      59492: inst = 32'd268468224;
      59493: inst = 32'd201348697;
      59494: inst = 32'd203423744;
      59495: inst = 32'd471859200;
      59496: inst = 32'd136314880;
      59497: inst = 32'd268468224;
      59498: inst = 32'd201348698;
      59499: inst = 32'd203423744;
      59500: inst = 32'd471859200;
      59501: inst = 32'd136314880;
      59502: inst = 32'd268468224;
      59503: inst = 32'd201348699;
      59504: inst = 32'd203423744;
      59505: inst = 32'd471859200;
      59506: inst = 32'd136314880;
      59507: inst = 32'd268468224;
      59508: inst = 32'd201348700;
      59509: inst = 32'd203423744;
      59510: inst = 32'd471859200;
      59511: inst = 32'd136314880;
      59512: inst = 32'd268468224;
      59513: inst = 32'd201348701;
      59514: inst = 32'd203423744;
      59515: inst = 32'd471859200;
      59516: inst = 32'd136314880;
      59517: inst = 32'd268468224;
      59518: inst = 32'd201348702;
      59519: inst = 32'd203423744;
      59520: inst = 32'd471859200;
      59521: inst = 32'd136314880;
      59522: inst = 32'd268468224;
      59523: inst = 32'd201348703;
      59524: inst = 32'd203423744;
      59525: inst = 32'd471859200;
      59526: inst = 32'd136314880;
      59527: inst = 32'd268468224;
      59528: inst = 32'd201348704;
      59529: inst = 32'd203423744;
      59530: inst = 32'd471859200;
      59531: inst = 32'd136314880;
      59532: inst = 32'd268468224;
      59533: inst = 32'd201348705;
      59534: inst = 32'd203423744;
      59535: inst = 32'd471859200;
      59536: inst = 32'd136314880;
      59537: inst = 32'd268468224;
      59538: inst = 32'd201348706;
      59539: inst = 32'd203423744;
      59540: inst = 32'd471859200;
      59541: inst = 32'd136314880;
      59542: inst = 32'd268468224;
      59543: inst = 32'd201348707;
      59544: inst = 32'd203423744;
      59545: inst = 32'd471859200;
      59546: inst = 32'd136314880;
      59547: inst = 32'd268468224;
      59548: inst = 32'd201348708;
      59549: inst = 32'd203423744;
      59550: inst = 32'd471859200;
      59551: inst = 32'd136314880;
      59552: inst = 32'd268468224;
      59553: inst = 32'd201348709;
      59554: inst = 32'd203423744;
      59555: inst = 32'd471859200;
      59556: inst = 32'd136314880;
      59557: inst = 32'd268468224;
      59558: inst = 32'd201348710;
      59559: inst = 32'd203423744;
      59560: inst = 32'd471859200;
      59561: inst = 32'd136314880;
      59562: inst = 32'd268468224;
      59563: inst = 32'd201348711;
      59564: inst = 32'd203423744;
      59565: inst = 32'd471859200;
      59566: inst = 32'd136314880;
      59567: inst = 32'd268468224;
      59568: inst = 32'd201348712;
      59569: inst = 32'd203423744;
      59570: inst = 32'd471859200;
      59571: inst = 32'd136314880;
      59572: inst = 32'd268468224;
      59573: inst = 32'd201348713;
      59574: inst = 32'd203423744;
      59575: inst = 32'd471859200;
      59576: inst = 32'd136314880;
      59577: inst = 32'd268468224;
      59578: inst = 32'd201348714;
      59579: inst = 32'd203423744;
      59580: inst = 32'd471859200;
      59581: inst = 32'd136314880;
      59582: inst = 32'd268468224;
      59583: inst = 32'd201348715;
      59584: inst = 32'd203423744;
      59585: inst = 32'd471859200;
      59586: inst = 32'd136314880;
      59587: inst = 32'd268468224;
      59588: inst = 32'd201348716;
      59589: inst = 32'd203423744;
      59590: inst = 32'd471859200;
      59591: inst = 32'd136314880;
      59592: inst = 32'd268468224;
      59593: inst = 32'd201348717;
      59594: inst = 32'd203423744;
      59595: inst = 32'd471859200;
      59596: inst = 32'd136314880;
      59597: inst = 32'd268468224;
      59598: inst = 32'd201348718;
      59599: inst = 32'd203423744;
      59600: inst = 32'd471859200;
      59601: inst = 32'd136314880;
      59602: inst = 32'd268468224;
      59603: inst = 32'd201348719;
      59604: inst = 32'd203423744;
      59605: inst = 32'd471859200;
      59606: inst = 32'd136314880;
      59607: inst = 32'd268468224;
      59608: inst = 32'd201348720;
      59609: inst = 32'd203423744;
      59610: inst = 32'd471859200;
      59611: inst = 32'd136314880;
      59612: inst = 32'd268468224;
      59613: inst = 32'd201348721;
      59614: inst = 32'd203423744;
      59615: inst = 32'd471859200;
      59616: inst = 32'd136314880;
      59617: inst = 32'd268468224;
      59618: inst = 32'd201348722;
      59619: inst = 32'd203423744;
      59620: inst = 32'd471859200;
      59621: inst = 32'd136314880;
      59622: inst = 32'd268468224;
      59623: inst = 32'd201348723;
      59624: inst = 32'd203423744;
      59625: inst = 32'd471859200;
      59626: inst = 32'd136314880;
      59627: inst = 32'd268468224;
      59628: inst = 32'd201348724;
      59629: inst = 32'd203423744;
      59630: inst = 32'd471859200;
      59631: inst = 32'd136314880;
      59632: inst = 32'd268468224;
      59633: inst = 32'd201348725;
      59634: inst = 32'd203423744;
      59635: inst = 32'd471859200;
      59636: inst = 32'd136314880;
      59637: inst = 32'd268468224;
      59638: inst = 32'd201348726;
      59639: inst = 32'd203423744;
      59640: inst = 32'd471859200;
      59641: inst = 32'd136314880;
      59642: inst = 32'd268468224;
      59643: inst = 32'd201348727;
      59644: inst = 32'd203423744;
      59645: inst = 32'd471859200;
      59646: inst = 32'd136314880;
      59647: inst = 32'd268468224;
      59648: inst = 32'd201348728;
      59649: inst = 32'd203423744;
      59650: inst = 32'd471859200;
      59651: inst = 32'd136314880;
      59652: inst = 32'd268468224;
      59653: inst = 32'd201348729;
      59654: inst = 32'd203423744;
      59655: inst = 32'd471859200;
      59656: inst = 32'd136314880;
      59657: inst = 32'd268468224;
      59658: inst = 32'd201348730;
      59659: inst = 32'd203423744;
      59660: inst = 32'd471859200;
      59661: inst = 32'd136314880;
      59662: inst = 32'd268468224;
      59663: inst = 32'd201348731;
      59664: inst = 32'd203423744;
      59665: inst = 32'd471859200;
      59666: inst = 32'd136314880;
      59667: inst = 32'd268468224;
      59668: inst = 32'd201348732;
      59669: inst = 32'd203423744;
      59670: inst = 32'd471859200;
      59671: inst = 32'd136314880;
      59672: inst = 32'd268468224;
      59673: inst = 32'd201348733;
      59674: inst = 32'd203423744;
      59675: inst = 32'd471859200;
      59676: inst = 32'd136314880;
      59677: inst = 32'd268468224;
      59678: inst = 32'd201348734;
      59679: inst = 32'd203423744;
      59680: inst = 32'd471859200;
      59681: inst = 32'd136314880;
      59682: inst = 32'd268468224;
      59683: inst = 32'd201348735;
      59684: inst = 32'd203423744;
      59685: inst = 32'd471859200;
      59686: inst = 32'd136314880;
      59687: inst = 32'd268468224;
      59688: inst = 32'd201348736;
      59689: inst = 32'd203423744;
      59690: inst = 32'd471859200;
      59691: inst = 32'd136314880;
      59692: inst = 32'd268468224;
      59693: inst = 32'd201348737;
      59694: inst = 32'd203423744;
      59695: inst = 32'd471859200;
      59696: inst = 32'd136314880;
      59697: inst = 32'd268468224;
      59698: inst = 32'd201348738;
      59699: inst = 32'd203423744;
      59700: inst = 32'd471859200;
      59701: inst = 32'd136314880;
      59702: inst = 32'd268468224;
      59703: inst = 32'd201348739;
      59704: inst = 32'd203423744;
      59705: inst = 32'd471859200;
      59706: inst = 32'd136314880;
      59707: inst = 32'd268468224;
      59708: inst = 32'd201348740;
      59709: inst = 32'd203423744;
      59710: inst = 32'd471859200;
      59711: inst = 32'd136314880;
      59712: inst = 32'd268468224;
      59713: inst = 32'd201348741;
      59714: inst = 32'd203423744;
      59715: inst = 32'd471859200;
      59716: inst = 32'd136314880;
      59717: inst = 32'd268468224;
      59718: inst = 32'd201348742;
      59719: inst = 32'd203423744;
      59720: inst = 32'd471859200;
      59721: inst = 32'd136314880;
      59722: inst = 32'd268468224;
      59723: inst = 32'd201348743;
      59724: inst = 32'd203423744;
      59725: inst = 32'd471859200;
      59726: inst = 32'd136314880;
      59727: inst = 32'd268468224;
      59728: inst = 32'd201348744;
      59729: inst = 32'd203423744;
      59730: inst = 32'd471859200;
      59731: inst = 32'd136314880;
      59732: inst = 32'd268468224;
      59733: inst = 32'd201348745;
      59734: inst = 32'd203423744;
      59735: inst = 32'd471859200;
      59736: inst = 32'd136314880;
      59737: inst = 32'd268468224;
      59738: inst = 32'd201348746;
      59739: inst = 32'd203423744;
      59740: inst = 32'd471859200;
      59741: inst = 32'd136314880;
      59742: inst = 32'd268468224;
      59743: inst = 32'd201348747;
      59744: inst = 32'd203423744;
      59745: inst = 32'd471859200;
      59746: inst = 32'd136314880;
      59747: inst = 32'd268468224;
      59748: inst = 32'd201348748;
      59749: inst = 32'd203423744;
      59750: inst = 32'd471859200;
      59751: inst = 32'd136314880;
      59752: inst = 32'd268468224;
      59753: inst = 32'd201348749;
      59754: inst = 32'd203423744;
      59755: inst = 32'd471859200;
      59756: inst = 32'd136314880;
      59757: inst = 32'd268468224;
      59758: inst = 32'd201348750;
      59759: inst = 32'd203423744;
      59760: inst = 32'd471859200;
      59761: inst = 32'd136314880;
      59762: inst = 32'd268468224;
      59763: inst = 32'd201348751;
      59764: inst = 32'd203423744;
      59765: inst = 32'd471859200;
      59766: inst = 32'd136314880;
      59767: inst = 32'd268468224;
      59768: inst = 32'd201348752;
      59769: inst = 32'd203423744;
      59770: inst = 32'd471859200;
      59771: inst = 32'd136314880;
      59772: inst = 32'd268468224;
      59773: inst = 32'd201348753;
      59774: inst = 32'd203423744;
      59775: inst = 32'd471859200;
      59776: inst = 32'd136314880;
      59777: inst = 32'd268468224;
      59778: inst = 32'd201348754;
      59779: inst = 32'd203423744;
      59780: inst = 32'd471859200;
      59781: inst = 32'd136314880;
      59782: inst = 32'd268468224;
      59783: inst = 32'd201348755;
      59784: inst = 32'd203423744;
      59785: inst = 32'd471859200;
      59786: inst = 32'd136314880;
      59787: inst = 32'd268468224;
      59788: inst = 32'd201348756;
      59789: inst = 32'd203423744;
      59790: inst = 32'd471859200;
      59791: inst = 32'd136314880;
      59792: inst = 32'd268468224;
      59793: inst = 32'd201348757;
      59794: inst = 32'd203423744;
      59795: inst = 32'd471859200;
      59796: inst = 32'd136314880;
      59797: inst = 32'd268468224;
      59798: inst = 32'd201348758;
      59799: inst = 32'd203423744;
      59800: inst = 32'd471859200;
      59801: inst = 32'd136314880;
      59802: inst = 32'd268468224;
      59803: inst = 32'd201348759;
      59804: inst = 32'd203423744;
      59805: inst = 32'd471859200;
      59806: inst = 32'd136314880;
      59807: inst = 32'd268468224;
      59808: inst = 32'd201348760;
      59809: inst = 32'd203423744;
      59810: inst = 32'd471859200;
      59811: inst = 32'd136314880;
      59812: inst = 32'd268468224;
      59813: inst = 32'd201348761;
      59814: inst = 32'd203423744;
      59815: inst = 32'd471859200;
      59816: inst = 32'd136314880;
      59817: inst = 32'd268468224;
      59818: inst = 32'd201348762;
      59819: inst = 32'd203423744;
      59820: inst = 32'd471859200;
      59821: inst = 32'd136314880;
      59822: inst = 32'd268468224;
      59823: inst = 32'd201348763;
      59824: inst = 32'd203423744;
      59825: inst = 32'd471859200;
      59826: inst = 32'd136314880;
      59827: inst = 32'd268468224;
      59828: inst = 32'd201348764;
      59829: inst = 32'd203423744;
      59830: inst = 32'd471859200;
      59831: inst = 32'd136314880;
      59832: inst = 32'd268468224;
      59833: inst = 32'd201348765;
      59834: inst = 32'd203423744;
      59835: inst = 32'd471859200;
      59836: inst = 32'd136314880;
      59837: inst = 32'd268468224;
      59838: inst = 32'd201348766;
      59839: inst = 32'd203423744;
      59840: inst = 32'd471859200;
      59841: inst = 32'd136314880;
      59842: inst = 32'd268468224;
      59843: inst = 32'd201348767;
      59844: inst = 32'd203423744;
      59845: inst = 32'd471859200;
      59846: inst = 32'd136314880;
      59847: inst = 32'd268468224;
      59848: inst = 32'd201348768;
      59849: inst = 32'd203423744;
      59850: inst = 32'd471859200;
      59851: inst = 32'd136314880;
      59852: inst = 32'd268468224;
      59853: inst = 32'd201348769;
      59854: inst = 32'd203423744;
      59855: inst = 32'd471859200;
      59856: inst = 32'd136314880;
      59857: inst = 32'd268468224;
      59858: inst = 32'd201348770;
      59859: inst = 32'd203423744;
      59860: inst = 32'd471859200;
      59861: inst = 32'd136314880;
      59862: inst = 32'd268468224;
      59863: inst = 32'd201348771;
      59864: inst = 32'd203423744;
      59865: inst = 32'd471859200;
      59866: inst = 32'd136314880;
      59867: inst = 32'd268468224;
      59868: inst = 32'd201348772;
      59869: inst = 32'd203423744;
      59870: inst = 32'd471859200;
      59871: inst = 32'd136314880;
      59872: inst = 32'd268468224;
      59873: inst = 32'd201348773;
      59874: inst = 32'd203423744;
      59875: inst = 32'd471859200;
      59876: inst = 32'd136314880;
      59877: inst = 32'd268468224;
      59878: inst = 32'd201348774;
      59879: inst = 32'd203423744;
      59880: inst = 32'd471859200;
      59881: inst = 32'd136314880;
      59882: inst = 32'd268468224;
      59883: inst = 32'd201348775;
      59884: inst = 32'd203423744;
      59885: inst = 32'd471859200;
      59886: inst = 32'd136314880;
      59887: inst = 32'd268468224;
      59888: inst = 32'd201348776;
      59889: inst = 32'd203423744;
      59890: inst = 32'd471859200;
      59891: inst = 32'd136314880;
      59892: inst = 32'd268468224;
      59893: inst = 32'd201348777;
      59894: inst = 32'd203423744;
      59895: inst = 32'd471859200;
      59896: inst = 32'd136314880;
      59897: inst = 32'd268468224;
      59898: inst = 32'd201348778;
      59899: inst = 32'd203423744;
      59900: inst = 32'd471859200;
      59901: inst = 32'd136314880;
      59902: inst = 32'd268468224;
      59903: inst = 32'd201348779;
      59904: inst = 32'd203423744;
      59905: inst = 32'd471859200;
      59906: inst = 32'd136314880;
      59907: inst = 32'd268468224;
      59908: inst = 32'd201348780;
      59909: inst = 32'd203423744;
      59910: inst = 32'd471859200;
      59911: inst = 32'd136314880;
      59912: inst = 32'd268468224;
      59913: inst = 32'd201348781;
      59914: inst = 32'd203423744;
      59915: inst = 32'd471859200;
      59916: inst = 32'd136314880;
      59917: inst = 32'd268468224;
      59918: inst = 32'd201348782;
      59919: inst = 32'd203423744;
      59920: inst = 32'd471859200;
      59921: inst = 32'd136314880;
      59922: inst = 32'd268468224;
      59923: inst = 32'd201348783;
      59924: inst = 32'd203423744;
      59925: inst = 32'd471859200;
      59926: inst = 32'd136314880;
      59927: inst = 32'd268468224;
      59928: inst = 32'd201348784;
      59929: inst = 32'd203423744;
      59930: inst = 32'd471859200;
      59931: inst = 32'd136314880;
      59932: inst = 32'd268468224;
      59933: inst = 32'd201348785;
      59934: inst = 32'd203423744;
      59935: inst = 32'd471859200;
      59936: inst = 32'd136314880;
      59937: inst = 32'd268468224;
      59938: inst = 32'd201348786;
      59939: inst = 32'd203423744;
      59940: inst = 32'd471859200;
      59941: inst = 32'd136314880;
      59942: inst = 32'd268468224;
      59943: inst = 32'd201348787;
      59944: inst = 32'd203423744;
      59945: inst = 32'd471859200;
      59946: inst = 32'd136314880;
      59947: inst = 32'd268468224;
      59948: inst = 32'd201348788;
      59949: inst = 32'd203423744;
      59950: inst = 32'd471859200;
      59951: inst = 32'd136314880;
      59952: inst = 32'd268468224;
      59953: inst = 32'd201348789;
      59954: inst = 32'd203423744;
      59955: inst = 32'd471859200;
      59956: inst = 32'd136314880;
      59957: inst = 32'd268468224;
      59958: inst = 32'd201348790;
      59959: inst = 32'd203423744;
      59960: inst = 32'd471859200;
      59961: inst = 32'd136314880;
      59962: inst = 32'd268468224;
      59963: inst = 32'd201348791;
      59964: inst = 32'd203423744;
      59965: inst = 32'd471859200;
      59966: inst = 32'd136314880;
      59967: inst = 32'd268468224;
      59968: inst = 32'd201348792;
      59969: inst = 32'd203423744;
      59970: inst = 32'd471859200;
      59971: inst = 32'd136314880;
      59972: inst = 32'd268468224;
      59973: inst = 32'd201348793;
      59974: inst = 32'd203423744;
      59975: inst = 32'd471859200;
      59976: inst = 32'd136314880;
      59977: inst = 32'd268468224;
      59978: inst = 32'd201348794;
      59979: inst = 32'd203423744;
      59980: inst = 32'd471859200;
      59981: inst = 32'd136314880;
      59982: inst = 32'd268468224;
      59983: inst = 32'd201348795;
      59984: inst = 32'd203423744;
      59985: inst = 32'd471859200;
      59986: inst = 32'd136314880;
      59987: inst = 32'd268468224;
      59988: inst = 32'd201348796;
      59989: inst = 32'd203423744;
      59990: inst = 32'd471859200;
      59991: inst = 32'd136314880;
      59992: inst = 32'd268468224;
      59993: inst = 32'd201348797;
      59994: inst = 32'd203423744;
      59995: inst = 32'd471859200;
      59996: inst = 32'd136314880;
      59997: inst = 32'd268468224;
      59998: inst = 32'd201348798;
      59999: inst = 32'd203423744;
      60000: inst = 32'd471859200;
      60001: inst = 32'd136314880;
      60002: inst = 32'd268468224;
      60003: inst = 32'd201348799;
      60004: inst = 32'd203423744;
      60005: inst = 32'd471859200;
      60006: inst = 32'd136314880;
      60007: inst = 32'd268468224;
      60008: inst = 32'd201348800;
      60009: inst = 32'd203423744;
      60010: inst = 32'd471859200;
      60011: inst = 32'd136314880;
      60012: inst = 32'd268468224;
      60013: inst = 32'd201348801;
      60014: inst = 32'd203423744;
      60015: inst = 32'd471859200;
      60016: inst = 32'd136314880;
      60017: inst = 32'd268468224;
      60018: inst = 32'd201348802;
      60019: inst = 32'd203423744;
      60020: inst = 32'd471859200;
      60021: inst = 32'd136314880;
      60022: inst = 32'd268468224;
      60023: inst = 32'd201348803;
      60024: inst = 32'd203423744;
      60025: inst = 32'd471859200;
      60026: inst = 32'd136314880;
      60027: inst = 32'd268468224;
      60028: inst = 32'd201348804;
      60029: inst = 32'd203423744;
      60030: inst = 32'd471859200;
      60031: inst = 32'd136314880;
      60032: inst = 32'd268468224;
      60033: inst = 32'd201348805;
      60034: inst = 32'd203423744;
      60035: inst = 32'd471859200;
      60036: inst = 32'd136314880;
      60037: inst = 32'd268468224;
      60038: inst = 32'd201348806;
      60039: inst = 32'd203423744;
      60040: inst = 32'd471859200;
      60041: inst = 32'd136314880;
      60042: inst = 32'd268468224;
      60043: inst = 32'd201348807;
      60044: inst = 32'd203423744;
      60045: inst = 32'd471859200;
      60046: inst = 32'd136314880;
      60047: inst = 32'd268468224;
      60048: inst = 32'd201348808;
      60049: inst = 32'd203423744;
      60050: inst = 32'd471859200;
      60051: inst = 32'd136314880;
      60052: inst = 32'd268468224;
      60053: inst = 32'd201348809;
      60054: inst = 32'd203423744;
      60055: inst = 32'd471859200;
      60056: inst = 32'd136314880;
      60057: inst = 32'd268468224;
      60058: inst = 32'd201348810;
      60059: inst = 32'd203423744;
      60060: inst = 32'd471859200;
      60061: inst = 32'd136314880;
      60062: inst = 32'd268468224;
      60063: inst = 32'd201348811;
      60064: inst = 32'd203423744;
      60065: inst = 32'd471859200;
      60066: inst = 32'd136314880;
      60067: inst = 32'd268468224;
      60068: inst = 32'd201348812;
      60069: inst = 32'd203423744;
      60070: inst = 32'd471859200;
      60071: inst = 32'd136314880;
      60072: inst = 32'd268468224;
      60073: inst = 32'd201348813;
      60074: inst = 32'd203423744;
      60075: inst = 32'd471859200;
      60076: inst = 32'd136314880;
      60077: inst = 32'd268468224;
      60078: inst = 32'd201348814;
      60079: inst = 32'd203423744;
      60080: inst = 32'd471859200;
      60081: inst = 32'd136314880;
      60082: inst = 32'd268468224;
      60083: inst = 32'd201348815;
      60084: inst = 32'd203423744;
      60085: inst = 32'd471859200;
      60086: inst = 32'd136314880;
      60087: inst = 32'd268468224;
      60088: inst = 32'd201348816;
      60089: inst = 32'd203423744;
      60090: inst = 32'd471859200;
      60091: inst = 32'd136314880;
      60092: inst = 32'd268468224;
      60093: inst = 32'd201348817;
      60094: inst = 32'd203423744;
      60095: inst = 32'd471859200;
      60096: inst = 32'd136314880;
      60097: inst = 32'd268468224;
      60098: inst = 32'd201348818;
      60099: inst = 32'd203423744;
      60100: inst = 32'd471859200;
      60101: inst = 32'd136314880;
      60102: inst = 32'd268468224;
      60103: inst = 32'd201348819;
      60104: inst = 32'd203423744;
      60105: inst = 32'd471859200;
      60106: inst = 32'd136314880;
      60107: inst = 32'd268468224;
      60108: inst = 32'd201348820;
      60109: inst = 32'd203423744;
      60110: inst = 32'd471859200;
      60111: inst = 32'd136314880;
      60112: inst = 32'd268468224;
      60113: inst = 32'd201348821;
      60114: inst = 32'd203423744;
      60115: inst = 32'd471859200;
      60116: inst = 32'd136314880;
      60117: inst = 32'd268468224;
      60118: inst = 32'd201348822;
      60119: inst = 32'd203423744;
      60120: inst = 32'd471859200;
      60121: inst = 32'd136314880;
      60122: inst = 32'd268468224;
      60123: inst = 32'd201348823;
      60124: inst = 32'd203423744;
      60125: inst = 32'd471859200;
      60126: inst = 32'd136314880;
      60127: inst = 32'd268468224;
      60128: inst = 32'd201348824;
      60129: inst = 32'd203423744;
      60130: inst = 32'd471859200;
      60131: inst = 32'd136314880;
      60132: inst = 32'd268468224;
      60133: inst = 32'd201348825;
      60134: inst = 32'd203423744;
      60135: inst = 32'd471859200;
      60136: inst = 32'd136314880;
      60137: inst = 32'd268468224;
      60138: inst = 32'd201348826;
      60139: inst = 32'd203423744;
      60140: inst = 32'd471859200;
      60141: inst = 32'd136314880;
      60142: inst = 32'd268468224;
      60143: inst = 32'd201348827;
      60144: inst = 32'd203423744;
      60145: inst = 32'd471859200;
      60146: inst = 32'd136314880;
      60147: inst = 32'd268468224;
      60148: inst = 32'd201348828;
      60149: inst = 32'd203423744;
      60150: inst = 32'd471859200;
      60151: inst = 32'd136314880;
      60152: inst = 32'd268468224;
      60153: inst = 32'd201348829;
      60154: inst = 32'd203423744;
      60155: inst = 32'd471859200;
      60156: inst = 32'd136314880;
      60157: inst = 32'd268468224;
      60158: inst = 32'd201348830;
      60159: inst = 32'd203423744;
      60160: inst = 32'd471859200;
      60161: inst = 32'd136314880;
      60162: inst = 32'd268468224;
      60163: inst = 32'd201348831;
      60164: inst = 32'd203423744;
      60165: inst = 32'd471859200;
      60166: inst = 32'd136314880;
      60167: inst = 32'd268468224;
      60168: inst = 32'd201348832;
      60169: inst = 32'd203423744;
      60170: inst = 32'd471859200;
      60171: inst = 32'd136314880;
      60172: inst = 32'd268468224;
      60173: inst = 32'd201348833;
      60174: inst = 32'd203423744;
      60175: inst = 32'd471859200;
      60176: inst = 32'd136314880;
      60177: inst = 32'd268468224;
      60178: inst = 32'd201348834;
      60179: inst = 32'd203423744;
      60180: inst = 32'd471859200;
      60181: inst = 32'd136314880;
      60182: inst = 32'd268468224;
      60183: inst = 32'd201348835;
      60184: inst = 32'd203423744;
      60185: inst = 32'd471859200;
      60186: inst = 32'd136314880;
      60187: inst = 32'd268468224;
      60188: inst = 32'd201348836;
      60189: inst = 32'd203423744;
      60190: inst = 32'd471859200;
      60191: inst = 32'd136314880;
      60192: inst = 32'd268468224;
      60193: inst = 32'd201348837;
      60194: inst = 32'd203423744;
      60195: inst = 32'd471859200;
      60196: inst = 32'd136314880;
      60197: inst = 32'd268468224;
      60198: inst = 32'd201348838;
      60199: inst = 32'd203423744;
      60200: inst = 32'd471859200;
      60201: inst = 32'd136314880;
      60202: inst = 32'd268468224;
      60203: inst = 32'd201348839;
      60204: inst = 32'd203423744;
      60205: inst = 32'd471859200;
      60206: inst = 32'd136314880;
      60207: inst = 32'd268468224;
      60208: inst = 32'd201348840;
      60209: inst = 32'd203423744;
      60210: inst = 32'd471859200;
      60211: inst = 32'd136314880;
      60212: inst = 32'd268468224;
      60213: inst = 32'd201348841;
      60214: inst = 32'd203423744;
      60215: inst = 32'd471859200;
      60216: inst = 32'd136314880;
      60217: inst = 32'd268468224;
      60218: inst = 32'd201348842;
      60219: inst = 32'd203423744;
      60220: inst = 32'd471859200;
      60221: inst = 32'd136314880;
      60222: inst = 32'd268468224;
      60223: inst = 32'd201348843;
      60224: inst = 32'd203423744;
      60225: inst = 32'd471859200;
      60226: inst = 32'd136314880;
      60227: inst = 32'd268468224;
      60228: inst = 32'd201348844;
      60229: inst = 32'd203423744;
      60230: inst = 32'd471859200;
      60231: inst = 32'd136314880;
      60232: inst = 32'd268468224;
      60233: inst = 32'd201348845;
      60234: inst = 32'd203423744;
      60235: inst = 32'd471859200;
      60236: inst = 32'd136314880;
      60237: inst = 32'd268468224;
      60238: inst = 32'd201348846;
      60239: inst = 32'd203423744;
      60240: inst = 32'd471859200;
      60241: inst = 32'd136314880;
      60242: inst = 32'd268468224;
      60243: inst = 32'd201348847;
      60244: inst = 32'd203423744;
      60245: inst = 32'd471859200;
      60246: inst = 32'd136314880;
      60247: inst = 32'd268468224;
      60248: inst = 32'd201348848;
      60249: inst = 32'd203423744;
      60250: inst = 32'd471859200;
      60251: inst = 32'd136314880;
      60252: inst = 32'd268468224;
      60253: inst = 32'd201348849;
      60254: inst = 32'd203423744;
      60255: inst = 32'd471859200;
      60256: inst = 32'd136314880;
      60257: inst = 32'd268468224;
      60258: inst = 32'd201348850;
      60259: inst = 32'd203423744;
      60260: inst = 32'd471859200;
      60261: inst = 32'd136314880;
      60262: inst = 32'd268468224;
      60263: inst = 32'd201348851;
      60264: inst = 32'd203423744;
      60265: inst = 32'd471859200;
      60266: inst = 32'd136314880;
      60267: inst = 32'd268468224;
      60268: inst = 32'd201348852;
      60269: inst = 32'd203423744;
      60270: inst = 32'd471859200;
      60271: inst = 32'd136314880;
      60272: inst = 32'd268468224;
      60273: inst = 32'd201348853;
      60274: inst = 32'd203423744;
      60275: inst = 32'd471859200;
      60276: inst = 32'd136314880;
      60277: inst = 32'd268468224;
      60278: inst = 32'd201348854;
      60279: inst = 32'd203423744;
      60280: inst = 32'd471859200;
      60281: inst = 32'd136314880;
      60282: inst = 32'd268468224;
      60283: inst = 32'd201348855;
      60284: inst = 32'd203423744;
      60285: inst = 32'd471859200;
      60286: inst = 32'd136314880;
      60287: inst = 32'd268468224;
      60288: inst = 32'd201348856;
      60289: inst = 32'd203423744;
      60290: inst = 32'd471859200;
      60291: inst = 32'd136314880;
      60292: inst = 32'd268468224;
      60293: inst = 32'd201348857;
      60294: inst = 32'd203423744;
      60295: inst = 32'd471859200;
      60296: inst = 32'd136314880;
      60297: inst = 32'd268468224;
      60298: inst = 32'd201348858;
      60299: inst = 32'd203423744;
      60300: inst = 32'd471859200;
      60301: inst = 32'd136314880;
      60302: inst = 32'd268468224;
      60303: inst = 32'd201348859;
      60304: inst = 32'd203423744;
      60305: inst = 32'd471859200;
      60306: inst = 32'd136314880;
      60307: inst = 32'd268468224;
      60308: inst = 32'd201348860;
      60309: inst = 32'd203423744;
      60310: inst = 32'd471859200;
      60311: inst = 32'd136314880;
      60312: inst = 32'd268468224;
      60313: inst = 32'd201348861;
      60314: inst = 32'd203423744;
      60315: inst = 32'd471859200;
      60316: inst = 32'd136314880;
      60317: inst = 32'd268468224;
      60318: inst = 32'd201348862;
      60319: inst = 32'd203423744;
      60320: inst = 32'd471859200;
      60321: inst = 32'd136314880;
      60322: inst = 32'd268468224;
      60323: inst = 32'd201348863;
      60324: inst = 32'd203423744;
      60325: inst = 32'd471859200;
      60326: inst = 32'd136314880;
      60327: inst = 32'd268468224;
      60328: inst = 32'd201348864;
      60329: inst = 32'd203423744;
      60330: inst = 32'd471859200;
      60331: inst = 32'd136314880;
      60332: inst = 32'd268468224;
      60333: inst = 32'd201348865;
      60334: inst = 32'd203423744;
      60335: inst = 32'd471859200;
      60336: inst = 32'd136314880;
      60337: inst = 32'd268468224;
      60338: inst = 32'd201348866;
      60339: inst = 32'd203423744;
      60340: inst = 32'd471859200;
      60341: inst = 32'd136314880;
      60342: inst = 32'd268468224;
      60343: inst = 32'd201348867;
      60344: inst = 32'd203423744;
      60345: inst = 32'd471859200;
      60346: inst = 32'd136314880;
      60347: inst = 32'd268468224;
      60348: inst = 32'd201348868;
      60349: inst = 32'd203423744;
      60350: inst = 32'd471859200;
      60351: inst = 32'd136314880;
      60352: inst = 32'd268468224;
      60353: inst = 32'd201348869;
      60354: inst = 32'd203423744;
      60355: inst = 32'd471859200;
      60356: inst = 32'd136314880;
      60357: inst = 32'd268468224;
      60358: inst = 32'd201348870;
      60359: inst = 32'd203423744;
      60360: inst = 32'd471859200;
      60361: inst = 32'd136314880;
      60362: inst = 32'd268468224;
      60363: inst = 32'd201348871;
      60364: inst = 32'd203423744;
      60365: inst = 32'd471859200;
      60366: inst = 32'd136314880;
      60367: inst = 32'd268468224;
      60368: inst = 32'd201348872;
      60369: inst = 32'd203423744;
      60370: inst = 32'd471859200;
      60371: inst = 32'd136314880;
      60372: inst = 32'd268468224;
      60373: inst = 32'd201348873;
      60374: inst = 32'd203423744;
      60375: inst = 32'd471859200;
      60376: inst = 32'd136314880;
      60377: inst = 32'd268468224;
      60378: inst = 32'd201348874;
      60379: inst = 32'd203423744;
      60380: inst = 32'd471859200;
      60381: inst = 32'd136314880;
      60382: inst = 32'd268468224;
      60383: inst = 32'd201348875;
      60384: inst = 32'd203423744;
      60385: inst = 32'd471859200;
      60386: inst = 32'd136314880;
      60387: inst = 32'd268468224;
      60388: inst = 32'd201348876;
      60389: inst = 32'd203423744;
      60390: inst = 32'd471859200;
      60391: inst = 32'd136314880;
      60392: inst = 32'd268468224;
      60393: inst = 32'd201348877;
      60394: inst = 32'd203423744;
      60395: inst = 32'd471859200;
      60396: inst = 32'd136314880;
      60397: inst = 32'd268468224;
      60398: inst = 32'd201348878;
      60399: inst = 32'd203423744;
      60400: inst = 32'd471859200;
      60401: inst = 32'd136314880;
      60402: inst = 32'd268468224;
      60403: inst = 32'd201348879;
      60404: inst = 32'd203423744;
      60405: inst = 32'd471859200;
      60406: inst = 32'd136314880;
      60407: inst = 32'd268468224;
      60408: inst = 32'd201348880;
      60409: inst = 32'd203423744;
      60410: inst = 32'd471859200;
      60411: inst = 32'd136314880;
      60412: inst = 32'd268468224;
      60413: inst = 32'd201348881;
      60414: inst = 32'd203423744;
      60415: inst = 32'd471859200;
      60416: inst = 32'd136314880;
      60417: inst = 32'd268468224;
      60418: inst = 32'd201348882;
      60419: inst = 32'd203423744;
      60420: inst = 32'd471859200;
      60421: inst = 32'd136314880;
      60422: inst = 32'd268468224;
      60423: inst = 32'd201348883;
      60424: inst = 32'd203423744;
      60425: inst = 32'd471859200;
      60426: inst = 32'd136314880;
      60427: inst = 32'd268468224;
      60428: inst = 32'd201348884;
      60429: inst = 32'd203423744;
      60430: inst = 32'd471859200;
      60431: inst = 32'd136314880;
      60432: inst = 32'd268468224;
      60433: inst = 32'd201348885;
      60434: inst = 32'd203423744;
      60435: inst = 32'd471859200;
      60436: inst = 32'd136314880;
      60437: inst = 32'd268468224;
      60438: inst = 32'd201348886;
      60439: inst = 32'd203423744;
      60440: inst = 32'd471859200;
      60441: inst = 32'd136314880;
      60442: inst = 32'd268468224;
      60443: inst = 32'd201348887;
      60444: inst = 32'd203423744;
      60445: inst = 32'd471859200;
      60446: inst = 32'd136314880;
      60447: inst = 32'd268468224;
      60448: inst = 32'd201348888;
      60449: inst = 32'd203423744;
      60450: inst = 32'd471859200;
      60451: inst = 32'd136314880;
      60452: inst = 32'd268468224;
      60453: inst = 32'd201348889;
      60454: inst = 32'd203423744;
      60455: inst = 32'd471859200;
      60456: inst = 32'd136314880;
      60457: inst = 32'd268468224;
      60458: inst = 32'd201348890;
      60459: inst = 32'd203423744;
      60460: inst = 32'd471859200;
      60461: inst = 32'd136314880;
      60462: inst = 32'd268468224;
      60463: inst = 32'd201348891;
      60464: inst = 32'd203423744;
      60465: inst = 32'd471859200;
      60466: inst = 32'd136314880;
      60467: inst = 32'd268468224;
      60468: inst = 32'd201348892;
      60469: inst = 32'd203423744;
      60470: inst = 32'd471859200;
      60471: inst = 32'd136314880;
      60472: inst = 32'd268468224;
      60473: inst = 32'd201348893;
      60474: inst = 32'd203423744;
      60475: inst = 32'd471859200;
      60476: inst = 32'd136314880;
      60477: inst = 32'd268468224;
      60478: inst = 32'd201348894;
      60479: inst = 32'd203423744;
      60480: inst = 32'd471859200;
      60481: inst = 32'd136314880;
      60482: inst = 32'd268468224;
      60483: inst = 32'd201348895;
      60484: inst = 32'd203423744;
      60485: inst = 32'd471859200;
      60486: inst = 32'd136314880;
      60487: inst = 32'd268468224;
      60488: inst = 32'd201348896;
      60489: inst = 32'd203423744;
      60490: inst = 32'd471859200;
      60491: inst = 32'd136314880;
      60492: inst = 32'd268468224;
      60493: inst = 32'd201348897;
      60494: inst = 32'd203423744;
      60495: inst = 32'd471859200;
      60496: inst = 32'd136314880;
      60497: inst = 32'd268468224;
      60498: inst = 32'd201348898;
      60499: inst = 32'd203423744;
      60500: inst = 32'd471859200;
      60501: inst = 32'd136314880;
      60502: inst = 32'd268468224;
      60503: inst = 32'd201348899;
      60504: inst = 32'd203423744;
      60505: inst = 32'd471859200;
      60506: inst = 32'd136314880;
      60507: inst = 32'd268468224;
      60508: inst = 32'd201348900;
      60509: inst = 32'd203423744;
      60510: inst = 32'd471859200;
      60511: inst = 32'd136314880;
      60512: inst = 32'd268468224;
      60513: inst = 32'd201348901;
      60514: inst = 32'd203423744;
      60515: inst = 32'd471859200;
      60516: inst = 32'd136314880;
      60517: inst = 32'd268468224;
      60518: inst = 32'd201348902;
      60519: inst = 32'd203423744;
      60520: inst = 32'd471859200;
      60521: inst = 32'd136314880;
      60522: inst = 32'd268468224;
      60523: inst = 32'd201348903;
      60524: inst = 32'd203423744;
      60525: inst = 32'd471859200;
      60526: inst = 32'd136314880;
      60527: inst = 32'd268468224;
      60528: inst = 32'd201348904;
      60529: inst = 32'd203423744;
      60530: inst = 32'd471859200;
      60531: inst = 32'd136314880;
      60532: inst = 32'd268468224;
      60533: inst = 32'd201348905;
      60534: inst = 32'd203423744;
      60535: inst = 32'd471859200;
      60536: inst = 32'd136314880;
      60537: inst = 32'd268468224;
      60538: inst = 32'd201348906;
      60539: inst = 32'd203423744;
      60540: inst = 32'd471859200;
      60541: inst = 32'd136314880;
      60542: inst = 32'd268468224;
      60543: inst = 32'd201348907;
      60544: inst = 32'd203423744;
      60545: inst = 32'd471859200;
      60546: inst = 32'd136314880;
      60547: inst = 32'd268468224;
      60548: inst = 32'd201348908;
      60549: inst = 32'd203423744;
      60550: inst = 32'd471859200;
      60551: inst = 32'd136314880;
      60552: inst = 32'd268468224;
      60553: inst = 32'd201348909;
      60554: inst = 32'd203423744;
      60555: inst = 32'd471859200;
      60556: inst = 32'd136314880;
      60557: inst = 32'd268468224;
      60558: inst = 32'd201348910;
      60559: inst = 32'd203423744;
      60560: inst = 32'd471859200;
      60561: inst = 32'd136314880;
      60562: inst = 32'd268468224;
      60563: inst = 32'd201348911;
      60564: inst = 32'd203423744;
      60565: inst = 32'd471859200;
      60566: inst = 32'd136314880;
      60567: inst = 32'd268468224;
      60568: inst = 32'd201348912;
      60569: inst = 32'd203423744;
      60570: inst = 32'd471859200;
      60571: inst = 32'd136314880;
      60572: inst = 32'd268468224;
      60573: inst = 32'd201348913;
      60574: inst = 32'd203423744;
      60575: inst = 32'd471859200;
      60576: inst = 32'd136314880;
      60577: inst = 32'd268468224;
      60578: inst = 32'd201348914;
      60579: inst = 32'd203423744;
      60580: inst = 32'd471859200;
      60581: inst = 32'd136314880;
      60582: inst = 32'd268468224;
      60583: inst = 32'd201348915;
      60584: inst = 32'd203423744;
      60585: inst = 32'd471859200;
      60586: inst = 32'd136314880;
      60587: inst = 32'd268468224;
      60588: inst = 32'd201348916;
      60589: inst = 32'd203423744;
      60590: inst = 32'd471859200;
      60591: inst = 32'd136314880;
      60592: inst = 32'd268468224;
      60593: inst = 32'd201348917;
      60594: inst = 32'd203423744;
      60595: inst = 32'd471859200;
      60596: inst = 32'd136314880;
      60597: inst = 32'd268468224;
      60598: inst = 32'd201348918;
      60599: inst = 32'd203423744;
      60600: inst = 32'd471859200;
      60601: inst = 32'd136314880;
      60602: inst = 32'd268468224;
      60603: inst = 32'd201348919;
      60604: inst = 32'd203423744;
      60605: inst = 32'd471859200;
      60606: inst = 32'd136314880;
      60607: inst = 32'd268468224;
      60608: inst = 32'd201348920;
      60609: inst = 32'd203423744;
      60610: inst = 32'd471859200;
      60611: inst = 32'd136314880;
      60612: inst = 32'd268468224;
      60613: inst = 32'd201348921;
      60614: inst = 32'd203423744;
      60615: inst = 32'd471859200;
      60616: inst = 32'd136314880;
      60617: inst = 32'd268468224;
      60618: inst = 32'd201348922;
      60619: inst = 32'd203423744;
      60620: inst = 32'd471859200;
      60621: inst = 32'd136314880;
      60622: inst = 32'd268468224;
      60623: inst = 32'd201348923;
      60624: inst = 32'd203423744;
      60625: inst = 32'd471859200;
      60626: inst = 32'd136314880;
      60627: inst = 32'd268468224;
      60628: inst = 32'd201348924;
      60629: inst = 32'd203423744;
      60630: inst = 32'd471859200;
      60631: inst = 32'd136314880;
      60632: inst = 32'd268468224;
      60633: inst = 32'd201348925;
      60634: inst = 32'd203423744;
      60635: inst = 32'd471859200;
      60636: inst = 32'd136314880;
      60637: inst = 32'd268468224;
      60638: inst = 32'd201348926;
      60639: inst = 32'd203423744;
      60640: inst = 32'd471859200;
      60641: inst = 32'd136314880;
      60642: inst = 32'd268468224;
      60643: inst = 32'd201348927;
      60644: inst = 32'd203423744;
      60645: inst = 32'd471859200;
      60646: inst = 32'd136314880;
      60647: inst = 32'd268468224;
      60648: inst = 32'd201348928;
      60649: inst = 32'd203423744;
      60650: inst = 32'd471859200;
      60651: inst = 32'd136314880;
      60652: inst = 32'd268468224;
      60653: inst = 32'd201348929;
      60654: inst = 32'd203423744;
      60655: inst = 32'd471859200;
      60656: inst = 32'd136314880;
      60657: inst = 32'd268468224;
      60658: inst = 32'd201348930;
      60659: inst = 32'd203423744;
      60660: inst = 32'd471859200;
      60661: inst = 32'd136314880;
      60662: inst = 32'd268468224;
      60663: inst = 32'd201348931;
      60664: inst = 32'd203423744;
      60665: inst = 32'd471859200;
      60666: inst = 32'd136314880;
      60667: inst = 32'd268468224;
      60668: inst = 32'd201348932;
      60669: inst = 32'd203423744;
      60670: inst = 32'd471859200;
      60671: inst = 32'd136314880;
      60672: inst = 32'd268468224;
      60673: inst = 32'd201348933;
      60674: inst = 32'd203423744;
      60675: inst = 32'd471859200;
      60676: inst = 32'd136314880;
      60677: inst = 32'd268468224;
      60678: inst = 32'd201348934;
      60679: inst = 32'd203423744;
      60680: inst = 32'd471859200;
      60681: inst = 32'd136314880;
      60682: inst = 32'd268468224;
      60683: inst = 32'd201348935;
      60684: inst = 32'd203423744;
      60685: inst = 32'd471859200;
      60686: inst = 32'd136314880;
      60687: inst = 32'd268468224;
      60688: inst = 32'd201348936;
      60689: inst = 32'd203423744;
      60690: inst = 32'd471859200;
      60691: inst = 32'd136314880;
      60692: inst = 32'd268468224;
      60693: inst = 32'd201348937;
      60694: inst = 32'd203423744;
      60695: inst = 32'd471859200;
      60696: inst = 32'd136314880;
      60697: inst = 32'd268468224;
      60698: inst = 32'd201348938;
      60699: inst = 32'd203423744;
      60700: inst = 32'd471859200;
      60701: inst = 32'd136314880;
      60702: inst = 32'd268468224;
      60703: inst = 32'd201348939;
      60704: inst = 32'd203423744;
      60705: inst = 32'd471859200;
      60706: inst = 32'd136314880;
      60707: inst = 32'd268468224;
      60708: inst = 32'd201348940;
      60709: inst = 32'd203423744;
      60710: inst = 32'd471859200;
      60711: inst = 32'd136314880;
      60712: inst = 32'd268468224;
      60713: inst = 32'd201348941;
      60714: inst = 32'd203423744;
      60715: inst = 32'd471859200;
      60716: inst = 32'd136314880;
      60717: inst = 32'd268468224;
      60718: inst = 32'd201348942;
      60719: inst = 32'd203423744;
      60720: inst = 32'd471859200;
      60721: inst = 32'd136314880;
      60722: inst = 32'd268468224;
      60723: inst = 32'd201348943;
      60724: inst = 32'd203423744;
      60725: inst = 32'd471859200;
      60726: inst = 32'd136314880;
      60727: inst = 32'd268468224;
      60728: inst = 32'd201348944;
      60729: inst = 32'd203423744;
      60730: inst = 32'd471859200;
      60731: inst = 32'd136314880;
      60732: inst = 32'd268468224;
      60733: inst = 32'd201348945;
      60734: inst = 32'd203423744;
      60735: inst = 32'd471859200;
      60736: inst = 32'd136314880;
      60737: inst = 32'd268468224;
      60738: inst = 32'd201348946;
      60739: inst = 32'd203423744;
      60740: inst = 32'd471859200;
      60741: inst = 32'd136314880;
      60742: inst = 32'd268468224;
      60743: inst = 32'd201348947;
      60744: inst = 32'd203423744;
      60745: inst = 32'd471859200;
      60746: inst = 32'd136314880;
      60747: inst = 32'd268468224;
      60748: inst = 32'd201348948;
      60749: inst = 32'd203423744;
      60750: inst = 32'd471859200;
      60751: inst = 32'd136314880;
      60752: inst = 32'd268468224;
      60753: inst = 32'd201348949;
      60754: inst = 32'd203423744;
      60755: inst = 32'd471859200;
      60756: inst = 32'd136314880;
      60757: inst = 32'd268468224;
      60758: inst = 32'd201348950;
      60759: inst = 32'd203423744;
      60760: inst = 32'd471859200;
      60761: inst = 32'd136314880;
      60762: inst = 32'd268468224;
      60763: inst = 32'd201348951;
      60764: inst = 32'd203423744;
      60765: inst = 32'd471859200;
      60766: inst = 32'd136314880;
      60767: inst = 32'd268468224;
      60768: inst = 32'd201348952;
      60769: inst = 32'd203423744;
      60770: inst = 32'd471859200;
      60771: inst = 32'd136314880;
      60772: inst = 32'd268468224;
      60773: inst = 32'd201348953;
      60774: inst = 32'd203423744;
      60775: inst = 32'd471859200;
      60776: inst = 32'd136314880;
      60777: inst = 32'd268468224;
      60778: inst = 32'd201348954;
      60779: inst = 32'd203423744;
      60780: inst = 32'd471859200;
      60781: inst = 32'd136314880;
      60782: inst = 32'd268468224;
      60783: inst = 32'd201348955;
      60784: inst = 32'd203423744;
      60785: inst = 32'd471859200;
      60786: inst = 32'd136314880;
      60787: inst = 32'd268468224;
      60788: inst = 32'd201348956;
      60789: inst = 32'd203423744;
      60790: inst = 32'd471859200;
      60791: inst = 32'd136314880;
      60792: inst = 32'd268468224;
      60793: inst = 32'd201348957;
      60794: inst = 32'd203423744;
      60795: inst = 32'd471859200;
      60796: inst = 32'd136314880;
      60797: inst = 32'd268468224;
      60798: inst = 32'd201348958;
      60799: inst = 32'd203423744;
      60800: inst = 32'd471859200;
      60801: inst = 32'd136314880;
      60802: inst = 32'd268468224;
      60803: inst = 32'd201348959;
      60804: inst = 32'd203423744;
      60805: inst = 32'd471859200;
      60806: inst = 32'd136314880;
      60807: inst = 32'd268468224;
      60808: inst = 32'd201348960;
      60809: inst = 32'd203423744;
      60810: inst = 32'd471859200;
      60811: inst = 32'd136314880;
      60812: inst = 32'd268468224;
      60813: inst = 32'd201348961;
      60814: inst = 32'd203423744;
      60815: inst = 32'd471859200;
      60816: inst = 32'd136314880;
      60817: inst = 32'd268468224;
      60818: inst = 32'd201348962;
      60819: inst = 32'd203423744;
      60820: inst = 32'd471859200;
      60821: inst = 32'd136314880;
      60822: inst = 32'd268468224;
      60823: inst = 32'd201348963;
      60824: inst = 32'd203423744;
      60825: inst = 32'd471859200;
      60826: inst = 32'd136314880;
      60827: inst = 32'd268468224;
      60828: inst = 32'd201348964;
      60829: inst = 32'd203423744;
      60830: inst = 32'd471859200;
      60831: inst = 32'd136314880;
      60832: inst = 32'd268468224;
      60833: inst = 32'd201348965;
      60834: inst = 32'd203423744;
      60835: inst = 32'd471859200;
      60836: inst = 32'd136314880;
      60837: inst = 32'd268468224;
      60838: inst = 32'd201348966;
      60839: inst = 32'd203423744;
      60840: inst = 32'd471859200;
      60841: inst = 32'd136314880;
      60842: inst = 32'd268468224;
      60843: inst = 32'd201348967;
      60844: inst = 32'd203423744;
      60845: inst = 32'd471859200;
      60846: inst = 32'd136314880;
      60847: inst = 32'd268468224;
      60848: inst = 32'd201348968;
      60849: inst = 32'd203423744;
      60850: inst = 32'd471859200;
      60851: inst = 32'd136314880;
      60852: inst = 32'd268468224;
      60853: inst = 32'd201348969;
      60854: inst = 32'd203423744;
      60855: inst = 32'd471859200;
      60856: inst = 32'd136314880;
      60857: inst = 32'd268468224;
      60858: inst = 32'd201348970;
      60859: inst = 32'd203423744;
      60860: inst = 32'd471859200;
      60861: inst = 32'd136314880;
      60862: inst = 32'd268468224;
      60863: inst = 32'd201348971;
      60864: inst = 32'd203423744;
      60865: inst = 32'd471859200;
      60866: inst = 32'd136314880;
      60867: inst = 32'd268468224;
      60868: inst = 32'd201348972;
      60869: inst = 32'd203423744;
      60870: inst = 32'd471859200;
      60871: inst = 32'd136314880;
      60872: inst = 32'd268468224;
      60873: inst = 32'd201348973;
      60874: inst = 32'd203423744;
      60875: inst = 32'd471859200;
      60876: inst = 32'd136314880;
      60877: inst = 32'd268468224;
      60878: inst = 32'd201348974;
      60879: inst = 32'd203423744;
      60880: inst = 32'd471859200;
      60881: inst = 32'd136314880;
      60882: inst = 32'd268468224;
      60883: inst = 32'd201348975;
      60884: inst = 32'd203423744;
      60885: inst = 32'd471859200;
      60886: inst = 32'd136314880;
      60887: inst = 32'd268468224;
      60888: inst = 32'd201348976;
      60889: inst = 32'd203423744;
      60890: inst = 32'd471859200;
      60891: inst = 32'd136314880;
      60892: inst = 32'd268468224;
      60893: inst = 32'd201348977;
      60894: inst = 32'd203423744;
      60895: inst = 32'd471859200;
      60896: inst = 32'd136314880;
      60897: inst = 32'd268468224;
      60898: inst = 32'd201348978;
      60899: inst = 32'd203423744;
      60900: inst = 32'd471859200;
      60901: inst = 32'd136314880;
      60902: inst = 32'd268468224;
      60903: inst = 32'd201348979;
      60904: inst = 32'd203423744;
      60905: inst = 32'd471859200;
      60906: inst = 32'd136314880;
      60907: inst = 32'd268468224;
      60908: inst = 32'd201348980;
      60909: inst = 32'd203423744;
      60910: inst = 32'd471859200;
      60911: inst = 32'd136314880;
      60912: inst = 32'd268468224;
      60913: inst = 32'd201348981;
      60914: inst = 32'd203423744;
      60915: inst = 32'd471859200;
      60916: inst = 32'd136314880;
      60917: inst = 32'd268468224;
      60918: inst = 32'd201348982;
      60919: inst = 32'd203423744;
      60920: inst = 32'd471859200;
      60921: inst = 32'd136314880;
      60922: inst = 32'd268468224;
      60923: inst = 32'd201348983;
      60924: inst = 32'd203423744;
      60925: inst = 32'd471859200;
      60926: inst = 32'd136314880;
      60927: inst = 32'd268468224;
      60928: inst = 32'd201348984;
      60929: inst = 32'd203423744;
      60930: inst = 32'd471859200;
      60931: inst = 32'd136314880;
      60932: inst = 32'd268468224;
      60933: inst = 32'd201348985;
      60934: inst = 32'd203423744;
      60935: inst = 32'd471859200;
      60936: inst = 32'd136314880;
      60937: inst = 32'd268468224;
      60938: inst = 32'd201348986;
      60939: inst = 32'd203423744;
      60940: inst = 32'd471859200;
      60941: inst = 32'd136314880;
      60942: inst = 32'd268468224;
      60943: inst = 32'd201348987;
      60944: inst = 32'd203423744;
      60945: inst = 32'd471859200;
      60946: inst = 32'd136314880;
      60947: inst = 32'd268468224;
      60948: inst = 32'd201348988;
      60949: inst = 32'd203423744;
      60950: inst = 32'd471859200;
      60951: inst = 32'd136314880;
      60952: inst = 32'd268468224;
      60953: inst = 32'd201348989;
      60954: inst = 32'd203423744;
      60955: inst = 32'd471859200;
      60956: inst = 32'd136314880;
      60957: inst = 32'd268468224;
      60958: inst = 32'd201348990;
      60959: inst = 32'd203423744;
      60960: inst = 32'd471859200;
      60961: inst = 32'd136314880;
      60962: inst = 32'd268468224;
      60963: inst = 32'd201348991;
      60964: inst = 32'd203423744;
      60965: inst = 32'd471859200;
      60966: inst = 32'd136314880;
      60967: inst = 32'd268468224;
      60968: inst = 32'd201348992;
      60969: inst = 32'd203423744;
      60970: inst = 32'd471859200;
      60971: inst = 32'd136314880;
      60972: inst = 32'd268468224;
      60973: inst = 32'd201348993;
      60974: inst = 32'd203423744;
      60975: inst = 32'd471859200;
      60976: inst = 32'd136314880;
      60977: inst = 32'd268468224;
      60978: inst = 32'd201348994;
      60979: inst = 32'd203423744;
      60980: inst = 32'd471859200;
      60981: inst = 32'd136314880;
      60982: inst = 32'd268468224;
      60983: inst = 32'd201348995;
      60984: inst = 32'd203423744;
      60985: inst = 32'd471859200;
      60986: inst = 32'd136314880;
      60987: inst = 32'd268468224;
      60988: inst = 32'd201348996;
      60989: inst = 32'd203423744;
      60990: inst = 32'd471859200;
      60991: inst = 32'd136314880;
      60992: inst = 32'd268468224;
      60993: inst = 32'd201348997;
      60994: inst = 32'd203423744;
      60995: inst = 32'd471859200;
      60996: inst = 32'd136314880;
      60997: inst = 32'd268468224;
      60998: inst = 32'd201348998;
      60999: inst = 32'd203423744;
      61000: inst = 32'd471859200;
      61001: inst = 32'd136314880;
      61002: inst = 32'd268468224;
      61003: inst = 32'd201348999;
      61004: inst = 32'd203423744;
      61005: inst = 32'd471859200;
      61006: inst = 32'd136314880;
      61007: inst = 32'd268468224;
      61008: inst = 32'd201349000;
      61009: inst = 32'd203423744;
      61010: inst = 32'd471859200;
      61011: inst = 32'd136314880;
      61012: inst = 32'd268468224;
      61013: inst = 32'd201349001;
      61014: inst = 32'd203423744;
      61015: inst = 32'd471859200;
      61016: inst = 32'd136314880;
      61017: inst = 32'd268468224;
      61018: inst = 32'd201349002;
      61019: inst = 32'd203423744;
      61020: inst = 32'd471859200;
      61021: inst = 32'd136314880;
      61022: inst = 32'd268468224;
      61023: inst = 32'd201349003;
      61024: inst = 32'd203423744;
      61025: inst = 32'd471859200;
      61026: inst = 32'd136314880;
      61027: inst = 32'd268468224;
      61028: inst = 32'd201349004;
      61029: inst = 32'd203423744;
      61030: inst = 32'd471859200;
      61031: inst = 32'd136314880;
      61032: inst = 32'd268468224;
      61033: inst = 32'd201349005;
      61034: inst = 32'd203423744;
      61035: inst = 32'd471859200;
      61036: inst = 32'd136314880;
      61037: inst = 32'd268468224;
      61038: inst = 32'd201349006;
      61039: inst = 32'd203423744;
      61040: inst = 32'd471859200;
      61041: inst = 32'd136314880;
      61042: inst = 32'd268468224;
      61043: inst = 32'd201349007;
      61044: inst = 32'd203423744;
      61045: inst = 32'd471859200;
      61046: inst = 32'd136314880;
      61047: inst = 32'd268468224;
      61048: inst = 32'd201349008;
      61049: inst = 32'd203423744;
      61050: inst = 32'd471859200;
      61051: inst = 32'd136314880;
      61052: inst = 32'd268468224;
      61053: inst = 32'd201349009;
      61054: inst = 32'd203423744;
      61055: inst = 32'd471859200;
      61056: inst = 32'd136314880;
      61057: inst = 32'd268468224;
      61058: inst = 32'd201349010;
      61059: inst = 32'd203423744;
      61060: inst = 32'd471859200;
      61061: inst = 32'd136314880;
      61062: inst = 32'd268468224;
      61063: inst = 32'd201349011;
      61064: inst = 32'd203423744;
      61065: inst = 32'd471859200;
      61066: inst = 32'd136314880;
      61067: inst = 32'd268468224;
      61068: inst = 32'd201349012;
      61069: inst = 32'd203423744;
      61070: inst = 32'd471859200;
      61071: inst = 32'd136314880;
      61072: inst = 32'd268468224;
      61073: inst = 32'd201349013;
      61074: inst = 32'd203423744;
      61075: inst = 32'd471859200;
      61076: inst = 32'd136314880;
      61077: inst = 32'd268468224;
      61078: inst = 32'd201349014;
      61079: inst = 32'd203423744;
      61080: inst = 32'd471859200;
      61081: inst = 32'd136314880;
      61082: inst = 32'd268468224;
      61083: inst = 32'd201349015;
      61084: inst = 32'd203423744;
      61085: inst = 32'd471859200;
      61086: inst = 32'd136314880;
      61087: inst = 32'd268468224;
      61088: inst = 32'd201349016;
      61089: inst = 32'd203423744;
      61090: inst = 32'd471859200;
      61091: inst = 32'd136314880;
      61092: inst = 32'd268468224;
      61093: inst = 32'd201349017;
      61094: inst = 32'd203423744;
      61095: inst = 32'd471859200;
      61096: inst = 32'd136314880;
      61097: inst = 32'd268468224;
      61098: inst = 32'd201349018;
      61099: inst = 32'd203423744;
      61100: inst = 32'd471859200;
      61101: inst = 32'd136314880;
      61102: inst = 32'd268468224;
      61103: inst = 32'd201349019;
      61104: inst = 32'd203423744;
      61105: inst = 32'd471859200;
      61106: inst = 32'd136314880;
      61107: inst = 32'd268468224;
      61108: inst = 32'd201349020;
      61109: inst = 32'd203423744;
      61110: inst = 32'd471859200;
      61111: inst = 32'd136314880;
      61112: inst = 32'd268468224;
      61113: inst = 32'd201349021;
      61114: inst = 32'd203423744;
      61115: inst = 32'd471859200;
      61116: inst = 32'd136314880;
      61117: inst = 32'd268468224;
      61118: inst = 32'd201349022;
      61119: inst = 32'd203423744;
      61120: inst = 32'd471859200;
      61121: inst = 32'd136314880;
      61122: inst = 32'd268468224;
      61123: inst = 32'd201349023;
      61124: inst = 32'd203423744;
      61125: inst = 32'd471859200;
      61126: inst = 32'd136314880;
      61127: inst = 32'd268468224;
      61128: inst = 32'd201349024;
      61129: inst = 32'd203423744;
      61130: inst = 32'd471859200;
      61131: inst = 32'd136314880;
      61132: inst = 32'd268468224;
      61133: inst = 32'd201349025;
      61134: inst = 32'd203423744;
      61135: inst = 32'd471859200;
      61136: inst = 32'd136314880;
      61137: inst = 32'd268468224;
      61138: inst = 32'd201349026;
      61139: inst = 32'd203423744;
      61140: inst = 32'd471859200;
      61141: inst = 32'd136314880;
      61142: inst = 32'd268468224;
      61143: inst = 32'd201349027;
      61144: inst = 32'd203423744;
      61145: inst = 32'd471859200;
      61146: inst = 32'd136314880;
      61147: inst = 32'd268468224;
      61148: inst = 32'd201349028;
      61149: inst = 32'd203423744;
      61150: inst = 32'd471859200;
      61151: inst = 32'd136314880;
      61152: inst = 32'd268468224;
      61153: inst = 32'd201349029;
      61154: inst = 32'd203423744;
      61155: inst = 32'd471859200;
      61156: inst = 32'd136314880;
      61157: inst = 32'd268468224;
      61158: inst = 32'd201349030;
      61159: inst = 32'd203423744;
      61160: inst = 32'd471859200;
      61161: inst = 32'd136314880;
      61162: inst = 32'd268468224;
      61163: inst = 32'd201349031;
      61164: inst = 32'd203423744;
      61165: inst = 32'd471859200;
      61166: inst = 32'd136314880;
      61167: inst = 32'd268468224;
      61168: inst = 32'd201349032;
      61169: inst = 32'd203423744;
      61170: inst = 32'd471859200;
      61171: inst = 32'd136314880;
      61172: inst = 32'd268468224;
      61173: inst = 32'd201349033;
      61174: inst = 32'd203423744;
      61175: inst = 32'd471859200;
      61176: inst = 32'd136314880;
      61177: inst = 32'd268468224;
      61178: inst = 32'd201349034;
      61179: inst = 32'd203423744;
      61180: inst = 32'd471859200;
      61181: inst = 32'd136314880;
      61182: inst = 32'd268468224;
      61183: inst = 32'd201349035;
      61184: inst = 32'd203423744;
      61185: inst = 32'd471859200;
      61186: inst = 32'd136314880;
      61187: inst = 32'd268468224;
      61188: inst = 32'd201349036;
      61189: inst = 32'd203423744;
      61190: inst = 32'd471859200;
      61191: inst = 32'd136314880;
      61192: inst = 32'd268468224;
      61193: inst = 32'd201349037;
      61194: inst = 32'd203423744;
      61195: inst = 32'd471859200;
      61196: inst = 32'd136314880;
      61197: inst = 32'd268468224;
      61198: inst = 32'd201349038;
      61199: inst = 32'd203423744;
      61200: inst = 32'd471859200;
      61201: inst = 32'd136314880;
      61202: inst = 32'd268468224;
      61203: inst = 32'd201349039;
      61204: inst = 32'd203423744;
      61205: inst = 32'd471859200;
      61206: inst = 32'd136314880;
      61207: inst = 32'd268468224;
      61208: inst = 32'd201349040;
      61209: inst = 32'd203423744;
      61210: inst = 32'd471859200;
      61211: inst = 32'd136314880;
      61212: inst = 32'd268468224;
      61213: inst = 32'd201349041;
      61214: inst = 32'd203423744;
      61215: inst = 32'd471859200;
      61216: inst = 32'd136314880;
      61217: inst = 32'd268468224;
      61218: inst = 32'd201349042;
      61219: inst = 32'd203423744;
      61220: inst = 32'd471859200;
      61221: inst = 32'd136314880;
      61222: inst = 32'd268468224;
      61223: inst = 32'd201349043;
      61224: inst = 32'd203423744;
      61225: inst = 32'd471859200;
      61226: inst = 32'd136314880;
      61227: inst = 32'd268468224;
      61228: inst = 32'd201349044;
      61229: inst = 32'd203423744;
      61230: inst = 32'd471859200;
      61231: inst = 32'd136314880;
      61232: inst = 32'd268468224;
      61233: inst = 32'd201349045;
      61234: inst = 32'd203423744;
      61235: inst = 32'd471859200;
      61236: inst = 32'd136314880;
      61237: inst = 32'd268468224;
      61238: inst = 32'd201349046;
      61239: inst = 32'd203423744;
      61240: inst = 32'd471859200;
      61241: inst = 32'd136314880;
      61242: inst = 32'd268468224;
      61243: inst = 32'd201349047;
      61244: inst = 32'd203423744;
      61245: inst = 32'd471859200;
      61246: inst = 32'd136314880;
      61247: inst = 32'd268468224;
      61248: inst = 32'd201349048;
      61249: inst = 32'd203423744;
      61250: inst = 32'd471859200;
      61251: inst = 32'd136314880;
      61252: inst = 32'd268468224;
      61253: inst = 32'd201349049;
      61254: inst = 32'd203423744;
      61255: inst = 32'd471859200;
      61256: inst = 32'd136314880;
      61257: inst = 32'd268468224;
      61258: inst = 32'd201349050;
      61259: inst = 32'd203423744;
      61260: inst = 32'd471859200;
      61261: inst = 32'd136314880;
      61262: inst = 32'd268468224;
      61263: inst = 32'd201349051;
      61264: inst = 32'd203423744;
      61265: inst = 32'd471859200;
      61266: inst = 32'd136314880;
      61267: inst = 32'd268468224;
      61268: inst = 32'd201349052;
      61269: inst = 32'd203423744;
      61270: inst = 32'd471859200;
      61271: inst = 32'd136314880;
      61272: inst = 32'd268468224;
      61273: inst = 32'd201349053;
      61274: inst = 32'd203423744;
      61275: inst = 32'd471859200;
      61276: inst = 32'd136314880;
      61277: inst = 32'd268468224;
      61278: inst = 32'd201349054;
      61279: inst = 32'd203423744;
      61280: inst = 32'd471859200;
      61281: inst = 32'd136314880;
      61282: inst = 32'd268468224;
      61283: inst = 32'd201349055;
      61284: inst = 32'd203423744;
      61285: inst = 32'd471859200;
      61286: inst = 32'd136314880;
      61287: inst = 32'd268468224;
      61288: inst = 32'd201349056;
      61289: inst = 32'd203423744;
      61290: inst = 32'd471859200;
      61291: inst = 32'd136314880;
      61292: inst = 32'd268468224;
      61293: inst = 32'd201349057;
      61294: inst = 32'd203423744;
      61295: inst = 32'd471859200;
      61296: inst = 32'd136314880;
      61297: inst = 32'd268468224;
      61298: inst = 32'd201349058;
      61299: inst = 32'd203423744;
      61300: inst = 32'd471859200;
      61301: inst = 32'd136314880;
      61302: inst = 32'd268468224;
      61303: inst = 32'd201349059;
      61304: inst = 32'd203423744;
      61305: inst = 32'd471859200;
      61306: inst = 32'd136314880;
      61307: inst = 32'd268468224;
      61308: inst = 32'd201349060;
      61309: inst = 32'd203423744;
      61310: inst = 32'd471859200;
      61311: inst = 32'd136314880;
      61312: inst = 32'd268468224;
      61313: inst = 32'd201349061;
      61314: inst = 32'd203423744;
      61315: inst = 32'd471859200;
      61316: inst = 32'd136314880;
      61317: inst = 32'd268468224;
      61318: inst = 32'd201349062;
      61319: inst = 32'd203423744;
      61320: inst = 32'd471859200;
      61321: inst = 32'd136314880;
      61322: inst = 32'd268468224;
      61323: inst = 32'd201349063;
      61324: inst = 32'd203423744;
      61325: inst = 32'd471859200;
      61326: inst = 32'd136314880;
      61327: inst = 32'd268468224;
      61328: inst = 32'd201349064;
      61329: inst = 32'd203423744;
      61330: inst = 32'd471859200;
      61331: inst = 32'd136314880;
      61332: inst = 32'd268468224;
      61333: inst = 32'd201349065;
      61334: inst = 32'd203423744;
      61335: inst = 32'd471859200;
      61336: inst = 32'd136314880;
      61337: inst = 32'd268468224;
      61338: inst = 32'd201349066;
      61339: inst = 32'd203423744;
      61340: inst = 32'd471859200;
      61341: inst = 32'd136314880;
      61342: inst = 32'd268468224;
      61343: inst = 32'd201349067;
      61344: inst = 32'd203423744;
      61345: inst = 32'd471859200;
      61346: inst = 32'd136314880;
      61347: inst = 32'd268468224;
      61348: inst = 32'd201349068;
      61349: inst = 32'd203423744;
      61350: inst = 32'd471859200;
      61351: inst = 32'd136314880;
      61352: inst = 32'd268468224;
      61353: inst = 32'd201349069;
      61354: inst = 32'd203423744;
      61355: inst = 32'd471859200;
      61356: inst = 32'd136314880;
      61357: inst = 32'd268468224;
      61358: inst = 32'd201349070;
      61359: inst = 32'd203423744;
      61360: inst = 32'd471859200;
      61361: inst = 32'd136314880;
      61362: inst = 32'd268468224;
      61363: inst = 32'd201349071;
      61364: inst = 32'd203423744;
      61365: inst = 32'd471859200;
      61366: inst = 32'd136314880;
      61367: inst = 32'd268468224;
      61368: inst = 32'd201349072;
      61369: inst = 32'd203423744;
      61370: inst = 32'd471859200;
      61371: inst = 32'd136314880;
      61372: inst = 32'd268468224;
      61373: inst = 32'd201349073;
      61374: inst = 32'd203423744;
      61375: inst = 32'd471859200;
      61376: inst = 32'd136314880;
      61377: inst = 32'd268468224;
      61378: inst = 32'd201349074;
      61379: inst = 32'd203423744;
      61380: inst = 32'd471859200;
      61381: inst = 32'd136314880;
      61382: inst = 32'd268468224;
      61383: inst = 32'd201349075;
      61384: inst = 32'd203423744;
      61385: inst = 32'd471859200;
      61386: inst = 32'd136314880;
      61387: inst = 32'd268468224;
      61388: inst = 32'd201349076;
      61389: inst = 32'd203423744;
      61390: inst = 32'd471859200;
      61391: inst = 32'd136314880;
      61392: inst = 32'd268468224;
      61393: inst = 32'd201349077;
      61394: inst = 32'd203423744;
      61395: inst = 32'd471859200;
      61396: inst = 32'd136314880;
      61397: inst = 32'd268468224;
      61398: inst = 32'd201349078;
      61399: inst = 32'd203423744;
      61400: inst = 32'd471859200;
      61401: inst = 32'd136314880;
      61402: inst = 32'd268468224;
      61403: inst = 32'd201349079;
      61404: inst = 32'd203423744;
      61405: inst = 32'd471859200;
      61406: inst = 32'd136314880;
      61407: inst = 32'd268468224;
      61408: inst = 32'd201349080;
      61409: inst = 32'd203423744;
      61410: inst = 32'd471859200;
      61411: inst = 32'd136314880;
      61412: inst = 32'd268468224;
      61413: inst = 32'd201349081;
      61414: inst = 32'd203423744;
      61415: inst = 32'd471859200;
      61416: inst = 32'd136314880;
      61417: inst = 32'd268468224;
      61418: inst = 32'd201349082;
      61419: inst = 32'd203423744;
      61420: inst = 32'd471859200;
      61421: inst = 32'd136314880;
      61422: inst = 32'd268468224;
      61423: inst = 32'd201349083;
      61424: inst = 32'd203423744;
      61425: inst = 32'd471859200;
      61426: inst = 32'd136314880;
      61427: inst = 32'd268468224;
      61428: inst = 32'd201349084;
      61429: inst = 32'd203423744;
      61430: inst = 32'd471859200;
      61431: inst = 32'd136314880;
      61432: inst = 32'd268468224;
      61433: inst = 32'd201349085;
      61434: inst = 32'd203423744;
      61435: inst = 32'd471859200;
      61436: inst = 32'd136314880;
      61437: inst = 32'd268468224;
      61438: inst = 32'd201349086;
      61439: inst = 32'd203423744;
      61440: inst = 32'd471859200;
      61441: inst = 32'd136314880;
      61442: inst = 32'd268468224;
      61443: inst = 32'd201349087;
      61444: inst = 32'd203423744;
      61445: inst = 32'd471859200;
      61446: inst = 32'd136314880;
      61447: inst = 32'd272629792;
      61448: inst = 32'd205520896;
      61449: inst = 32'd809631745;
      61450: inst = 32'd333447168;
      61451: inst = 32'd266399753;
      61452: inst = 32'd473956352;
      61453: inst = 32'd1541406720;
      61454: inst = 32'd333447168;
      61455: inst = 32'd266338304;
      61456: inst = 32'd1541406720;
    endcase
  end
endmodule
