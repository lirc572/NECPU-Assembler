`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: lirc572
// Engineer: lirc572
// 
// Create Date: 
// Design Name: NECPU
// Module Name: InstMem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module instMem (
    input  [31:0]  address,
    output reg [31:0] inst
  );
  always @ (address) begin
    inst = 32'd0;
    case (address)
      0: inst = 32'h10000000;
      1: inst = 32'hc000005;
      2: inst = 32'h13e00000;
      3: inst = 32'hfe00055;
      4: inst = 32'h5be00000;
      5: inst = 32'h13c0007f;
      6: inst = 32'hfc02815;
      7: inst = 32'h33de0001;
      8: inst = 32'h13e00000;
      9: inst = 32'hfe00007;
      10: inst = 32'h1fc00000;
      11: inst = 32'h5be00000;
      12: inst = 32'h10000000;
      13: inst = 32'hc000011;
      14: inst = 32'h13e00000;
      15: inst = 32'hfe048ad;
      16: inst = 32'h5be00000;
      17: inst = 32'h13c0007f;
      18: inst = 32'hfc02815;
      19: inst = 32'h33de0001;
      20: inst = 32'h13e00000;
      21: inst = 32'hfe00013;
      22: inst = 32'h1fc00000;
      23: inst = 32'h5be00000;
      24: inst = 32'h10000000;
      25: inst = 32'hc000000;
      26: inst = 32'h10200000;
      27: inst = 32'hc20001f;
      28: inst = 32'h13e00000;
      29: inst = 32'hfe08960;
      30: inst = 32'h5be00000;
      31: inst = 32'h10000000;
      32: inst = 32'hc000024;
      33: inst = 32'h13e00000;
      34: inst = 32'hfe050fe;
      35: inst = 32'h5be00000;
      36: inst = 32'h13c001fc;
      37: inst = 32'hfc0a055;
      38: inst = 32'h33de0001;
      39: inst = 32'h13e00000;
      40: inst = 32'hfe00026;
      41: inst = 32'h1fc00000;
      42: inst = 32'h5be00000;
      43: inst = 32'h10000000;
      44: inst = 32'hc00002b;
      45: inst = 32'h10200000;
      46: inst = 32'hc200032;
      47: inst = 32'h13e00000;
      48: inst = 32'hfe08960;
      49: inst = 32'h5be00000;
      50: inst = 32'h10200000;
      51: inst = 32'hc20000c;
      52: inst = 32'h10400000;
      53: inst = 32'hc400009;
      54: inst = 32'h10000000;
      55: inst = 32'hc00003b;
      56: inst = 32'h13e00000;
      57: inst = 32'hfe0896a;
      58: inst = 32'h5be00000;
      59: inst = 32'h10200000;
      60: inst = 32'hc200000;
      61: inst = 32'h10000000;
      62: inst = 32'hc000042;
      63: inst = 32'h13e00000;
      64: inst = 32'hfe085ad;
      65: inst = 32'h5be00000;
      66: inst = 32'h13e00000;
      67: inst = 32'hfe00045;
      68: inst = 32'h5be00000;
      69: inst = 32'h10608000;
      70: inst = 32'hc600000;
      71: inst = 32'h10200000;
      72: inst = 32'hc20aaaa;
      73: inst = 32'h4c210000;
      74: inst = 32'h8230000;
      75: inst = 32'h104000fe;
      76: inst = 32'hc40502a;
      77: inst = 32'h30420001;
      78: inst = 32'h13e00000;
      79: inst = 32'hfe0004d;
      80: inst = 32'h1c400000;
      81: inst = 32'h5be00000;
      82: inst = 32'h13e00000;
      83: inst = 32'hfe00049;
      84: inst = 32'h5be00000;
      85: inst = 32'hc20eeb6;
      86: inst = 32'h10408000;
      87: inst = 32'hc403fe0;
      88: inst = 32'h8220000;
      89: inst = 32'h10408000;
      90: inst = 32'hc403fe1;
      91: inst = 32'h8220000;
      92: inst = 32'h10408000;
      93: inst = 32'hc403fe2;
      94: inst = 32'h8220000;
      95: inst = 32'h10408000;
      96: inst = 32'hc403fe3;
      97: inst = 32'h8220000;
      98: inst = 32'h10408000;
      99: inst = 32'hc403fe4;
      100: inst = 32'h8220000;
      101: inst = 32'h10408000;
      102: inst = 32'hc403fe5;
      103: inst = 32'h8220000;
      104: inst = 32'h10408000;
      105: inst = 32'hc403fe6;
      106: inst = 32'h8220000;
      107: inst = 32'h10408000;
      108: inst = 32'hc403fe7;
      109: inst = 32'h8220000;
      110: inst = 32'h10408000;
      111: inst = 32'hc403fe8;
      112: inst = 32'h8220000;
      113: inst = 32'h10408000;
      114: inst = 32'hc403fe9;
      115: inst = 32'h8220000;
      116: inst = 32'h10408000;
      117: inst = 32'hc403fea;
      118: inst = 32'h8220000;
      119: inst = 32'h10408000;
      120: inst = 32'hc403fec;
      121: inst = 32'h8220000;
      122: inst = 32'h10408000;
      123: inst = 32'hc403fed;
      124: inst = 32'h8220000;
      125: inst = 32'h10408000;
      126: inst = 32'hc403fee;
      127: inst = 32'h8220000;
      128: inst = 32'h10408000;
      129: inst = 32'hc403fef;
      130: inst = 32'h8220000;
      131: inst = 32'h10408000;
      132: inst = 32'hc403ff0;
      133: inst = 32'h8220000;
      134: inst = 32'h10408000;
      135: inst = 32'hc403ff1;
      136: inst = 32'h8220000;
      137: inst = 32'h10408000;
      138: inst = 32'hc403ff2;
      139: inst = 32'h8220000;
      140: inst = 32'h10408000;
      141: inst = 32'hc403ff3;
      142: inst = 32'h8220000;
      143: inst = 32'h10408000;
      144: inst = 32'hc403ff4;
      145: inst = 32'h8220000;
      146: inst = 32'h10408000;
      147: inst = 32'hc403ff5;
      148: inst = 32'h8220000;
      149: inst = 32'h10408000;
      150: inst = 32'hc403ff6;
      151: inst = 32'h8220000;
      152: inst = 32'h10408000;
      153: inst = 32'hc403ff7;
      154: inst = 32'h8220000;
      155: inst = 32'h10408000;
      156: inst = 32'hc403ff8;
      157: inst = 32'h8220000;
      158: inst = 32'h10408000;
      159: inst = 32'hc403ff9;
      160: inst = 32'h8220000;
      161: inst = 32'h10408000;
      162: inst = 32'hc403ffa;
      163: inst = 32'h8220000;
      164: inst = 32'h10408000;
      165: inst = 32'hc403ffb;
      166: inst = 32'h8220000;
      167: inst = 32'h10408000;
      168: inst = 32'hc403ffc;
      169: inst = 32'h8220000;
      170: inst = 32'h10408000;
      171: inst = 32'hc403ffd;
      172: inst = 32'h8220000;
      173: inst = 32'h10408000;
      174: inst = 32'hc403ffe;
      175: inst = 32'h8220000;
      176: inst = 32'h10408000;
      177: inst = 32'hc403fff;
      178: inst = 32'h8220000;
      179: inst = 32'h10408000;
      180: inst = 32'hc404000;
      181: inst = 32'h8220000;
      182: inst = 32'h10408000;
      183: inst = 32'hc404001;
      184: inst = 32'h8220000;
      185: inst = 32'h10408000;
      186: inst = 32'hc404002;
      187: inst = 32'h8220000;
      188: inst = 32'h10408000;
      189: inst = 32'hc404003;
      190: inst = 32'h8220000;
      191: inst = 32'h10408000;
      192: inst = 32'hc404004;
      193: inst = 32'h8220000;
      194: inst = 32'h10408000;
      195: inst = 32'hc404005;
      196: inst = 32'h8220000;
      197: inst = 32'h10408000;
      198: inst = 32'hc404006;
      199: inst = 32'h8220000;
      200: inst = 32'h10408000;
      201: inst = 32'hc404007;
      202: inst = 32'h8220000;
      203: inst = 32'h10408000;
      204: inst = 32'hc404008;
      205: inst = 32'h8220000;
      206: inst = 32'h10408000;
      207: inst = 32'hc404009;
      208: inst = 32'h8220000;
      209: inst = 32'h10408000;
      210: inst = 32'hc40400a;
      211: inst = 32'h8220000;
      212: inst = 32'h10408000;
      213: inst = 32'hc40400b;
      214: inst = 32'h8220000;
      215: inst = 32'h10408000;
      216: inst = 32'hc40400c;
      217: inst = 32'h8220000;
      218: inst = 32'h10408000;
      219: inst = 32'hc40400d;
      220: inst = 32'h8220000;
      221: inst = 32'h10408000;
      222: inst = 32'hc40400e;
      223: inst = 32'h8220000;
      224: inst = 32'h10408000;
      225: inst = 32'hc40400f;
      226: inst = 32'h8220000;
      227: inst = 32'h10408000;
      228: inst = 32'hc404010;
      229: inst = 32'h8220000;
      230: inst = 32'h10408000;
      231: inst = 32'hc404011;
      232: inst = 32'h8220000;
      233: inst = 32'h10408000;
      234: inst = 32'hc404012;
      235: inst = 32'h8220000;
      236: inst = 32'h10408000;
      237: inst = 32'hc404013;
      238: inst = 32'h8220000;
      239: inst = 32'h10408000;
      240: inst = 32'hc404014;
      241: inst = 32'h8220000;
      242: inst = 32'h10408000;
      243: inst = 32'hc404015;
      244: inst = 32'h8220000;
      245: inst = 32'h10408000;
      246: inst = 32'hc404016;
      247: inst = 32'h8220000;
      248: inst = 32'h10408000;
      249: inst = 32'hc404017;
      250: inst = 32'h8220000;
      251: inst = 32'h10408000;
      252: inst = 32'hc404018;
      253: inst = 32'h8220000;
      254: inst = 32'h10408000;
      255: inst = 32'hc404019;
      256: inst = 32'h8220000;
      257: inst = 32'h10408000;
      258: inst = 32'hc40401a;
      259: inst = 32'h8220000;
      260: inst = 32'h10408000;
      261: inst = 32'hc40401b;
      262: inst = 32'h8220000;
      263: inst = 32'h10408000;
      264: inst = 32'hc40401c;
      265: inst = 32'h8220000;
      266: inst = 32'h10408000;
      267: inst = 32'hc40401d;
      268: inst = 32'h8220000;
      269: inst = 32'h10408000;
      270: inst = 32'hc40401e;
      271: inst = 32'h8220000;
      272: inst = 32'h10408000;
      273: inst = 32'hc40401f;
      274: inst = 32'h8220000;
      275: inst = 32'h10408000;
      276: inst = 32'hc404020;
      277: inst = 32'h8220000;
      278: inst = 32'h10408000;
      279: inst = 32'hc404021;
      280: inst = 32'h8220000;
      281: inst = 32'h10408000;
      282: inst = 32'hc404022;
      283: inst = 32'h8220000;
      284: inst = 32'h10408000;
      285: inst = 32'hc404023;
      286: inst = 32'h8220000;
      287: inst = 32'h10408000;
      288: inst = 32'hc404024;
      289: inst = 32'h8220000;
      290: inst = 32'h10408000;
      291: inst = 32'hc404025;
      292: inst = 32'h8220000;
      293: inst = 32'h10408000;
      294: inst = 32'hc404026;
      295: inst = 32'h8220000;
      296: inst = 32'h10408000;
      297: inst = 32'hc404027;
      298: inst = 32'h8220000;
      299: inst = 32'h10408000;
      300: inst = 32'hc404028;
      301: inst = 32'h8220000;
      302: inst = 32'h10408000;
      303: inst = 32'hc404029;
      304: inst = 32'h8220000;
      305: inst = 32'h10408000;
      306: inst = 32'hc40402a;
      307: inst = 32'h8220000;
      308: inst = 32'h10408000;
      309: inst = 32'hc40402b;
      310: inst = 32'h8220000;
      311: inst = 32'h10408000;
      312: inst = 32'hc40402c;
      313: inst = 32'h8220000;
      314: inst = 32'h10408000;
      315: inst = 32'hc40402d;
      316: inst = 32'h8220000;
      317: inst = 32'h10408000;
      318: inst = 32'hc40402e;
      319: inst = 32'h8220000;
      320: inst = 32'h10408000;
      321: inst = 32'hc40402f;
      322: inst = 32'h8220000;
      323: inst = 32'h10408000;
      324: inst = 32'hc404030;
      325: inst = 32'h8220000;
      326: inst = 32'h10408000;
      327: inst = 32'hc404031;
      328: inst = 32'h8220000;
      329: inst = 32'h10408000;
      330: inst = 32'hc404032;
      331: inst = 32'h8220000;
      332: inst = 32'h10408000;
      333: inst = 32'hc404033;
      334: inst = 32'h8220000;
      335: inst = 32'h10408000;
      336: inst = 32'hc404034;
      337: inst = 32'h8220000;
      338: inst = 32'h10408000;
      339: inst = 32'hc404035;
      340: inst = 32'h8220000;
      341: inst = 32'h10408000;
      342: inst = 32'hc404036;
      343: inst = 32'h8220000;
      344: inst = 32'h10408000;
      345: inst = 32'hc404037;
      346: inst = 32'h8220000;
      347: inst = 32'h10408000;
      348: inst = 32'hc404038;
      349: inst = 32'h8220000;
      350: inst = 32'h10408000;
      351: inst = 32'hc404039;
      352: inst = 32'h8220000;
      353: inst = 32'h10408000;
      354: inst = 32'hc40403a;
      355: inst = 32'h8220000;
      356: inst = 32'h10408000;
      357: inst = 32'hc40403b;
      358: inst = 32'h8220000;
      359: inst = 32'h10408000;
      360: inst = 32'hc40403c;
      361: inst = 32'h8220000;
      362: inst = 32'h10408000;
      363: inst = 32'hc40403d;
      364: inst = 32'h8220000;
      365: inst = 32'h10408000;
      366: inst = 32'hc40403e;
      367: inst = 32'h8220000;
      368: inst = 32'h10408000;
      369: inst = 32'hc40403f;
      370: inst = 32'h8220000;
      371: inst = 32'h10408000;
      372: inst = 32'hc404040;
      373: inst = 32'h8220000;
      374: inst = 32'h10408000;
      375: inst = 32'hc404041;
      376: inst = 32'h8220000;
      377: inst = 32'h10408000;
      378: inst = 32'hc404042;
      379: inst = 32'h8220000;
      380: inst = 32'h10408000;
      381: inst = 32'hc404043;
      382: inst = 32'h8220000;
      383: inst = 32'h10408000;
      384: inst = 32'hc404044;
      385: inst = 32'h8220000;
      386: inst = 32'h10408000;
      387: inst = 32'hc404045;
      388: inst = 32'h8220000;
      389: inst = 32'h10408000;
      390: inst = 32'hc404046;
      391: inst = 32'h8220000;
      392: inst = 32'h10408000;
      393: inst = 32'hc404047;
      394: inst = 32'h8220000;
      395: inst = 32'h10408000;
      396: inst = 32'hc404048;
      397: inst = 32'h8220000;
      398: inst = 32'h10408000;
      399: inst = 32'hc404049;
      400: inst = 32'h8220000;
      401: inst = 32'h10408000;
      402: inst = 32'hc40404a;
      403: inst = 32'h8220000;
      404: inst = 32'h10408000;
      405: inst = 32'hc40404c;
      406: inst = 32'h8220000;
      407: inst = 32'h10408000;
      408: inst = 32'hc40404d;
      409: inst = 32'h8220000;
      410: inst = 32'h10408000;
      411: inst = 32'hc40404e;
      412: inst = 32'h8220000;
      413: inst = 32'h10408000;
      414: inst = 32'hc40404f;
      415: inst = 32'h8220000;
      416: inst = 32'h10408000;
      417: inst = 32'hc404050;
      418: inst = 32'h8220000;
      419: inst = 32'h10408000;
      420: inst = 32'hc404051;
      421: inst = 32'h8220000;
      422: inst = 32'h10408000;
      423: inst = 32'hc404052;
      424: inst = 32'h8220000;
      425: inst = 32'h10408000;
      426: inst = 32'hc404053;
      427: inst = 32'h8220000;
      428: inst = 32'h10408000;
      429: inst = 32'hc404054;
      430: inst = 32'h8220000;
      431: inst = 32'h10408000;
      432: inst = 32'hc404055;
      433: inst = 32'h8220000;
      434: inst = 32'h10408000;
      435: inst = 32'hc404056;
      436: inst = 32'h8220000;
      437: inst = 32'h10408000;
      438: inst = 32'hc404057;
      439: inst = 32'h8220000;
      440: inst = 32'h10408000;
      441: inst = 32'hc404058;
      442: inst = 32'h8220000;
      443: inst = 32'h10408000;
      444: inst = 32'hc404059;
      445: inst = 32'h8220000;
      446: inst = 32'h10408000;
      447: inst = 32'hc40405a;
      448: inst = 32'h8220000;
      449: inst = 32'h10408000;
      450: inst = 32'hc40405b;
      451: inst = 32'h8220000;
      452: inst = 32'h10408000;
      453: inst = 32'hc40405c;
      454: inst = 32'h8220000;
      455: inst = 32'h10408000;
      456: inst = 32'hc40405d;
      457: inst = 32'h8220000;
      458: inst = 32'h10408000;
      459: inst = 32'hc40405e;
      460: inst = 32'h8220000;
      461: inst = 32'h10408000;
      462: inst = 32'hc40405f;
      463: inst = 32'h8220000;
      464: inst = 32'h10408000;
      465: inst = 32'hc404060;
      466: inst = 32'h8220000;
      467: inst = 32'h10408000;
      468: inst = 32'hc404061;
      469: inst = 32'h8220000;
      470: inst = 32'h10408000;
      471: inst = 32'hc404062;
      472: inst = 32'h8220000;
      473: inst = 32'h10408000;
      474: inst = 32'hc404063;
      475: inst = 32'h8220000;
      476: inst = 32'h10408000;
      477: inst = 32'hc404064;
      478: inst = 32'h8220000;
      479: inst = 32'h10408000;
      480: inst = 32'hc404065;
      481: inst = 32'h8220000;
      482: inst = 32'h10408000;
      483: inst = 32'hc404066;
      484: inst = 32'h8220000;
      485: inst = 32'h10408000;
      486: inst = 32'hc404067;
      487: inst = 32'h8220000;
      488: inst = 32'h10408000;
      489: inst = 32'hc404068;
      490: inst = 32'h8220000;
      491: inst = 32'h10408000;
      492: inst = 32'hc404069;
      493: inst = 32'h8220000;
      494: inst = 32'h10408000;
      495: inst = 32'hc40406a;
      496: inst = 32'h8220000;
      497: inst = 32'h10408000;
      498: inst = 32'hc40406b;
      499: inst = 32'h8220000;
      500: inst = 32'h10408000;
      501: inst = 32'hc40406c;
      502: inst = 32'h8220000;
      503: inst = 32'h10408000;
      504: inst = 32'hc40406d;
      505: inst = 32'h8220000;
      506: inst = 32'h10408000;
      507: inst = 32'hc40406e;
      508: inst = 32'h8220000;
      509: inst = 32'h10408000;
      510: inst = 32'hc40406f;
      511: inst = 32'h8220000;
      512: inst = 32'h10408000;
      513: inst = 32'hc404070;
      514: inst = 32'h8220000;
      515: inst = 32'h10408000;
      516: inst = 32'hc404071;
      517: inst = 32'h8220000;
      518: inst = 32'h10408000;
      519: inst = 32'hc404072;
      520: inst = 32'h8220000;
      521: inst = 32'h10408000;
      522: inst = 32'hc404073;
      523: inst = 32'h8220000;
      524: inst = 32'h10408000;
      525: inst = 32'hc404074;
      526: inst = 32'h8220000;
      527: inst = 32'h10408000;
      528: inst = 32'hc404075;
      529: inst = 32'h8220000;
      530: inst = 32'h10408000;
      531: inst = 32'hc404076;
      532: inst = 32'h8220000;
      533: inst = 32'h10408000;
      534: inst = 32'hc404077;
      535: inst = 32'h8220000;
      536: inst = 32'h10408000;
      537: inst = 32'hc404078;
      538: inst = 32'h8220000;
      539: inst = 32'h10408000;
      540: inst = 32'hc404079;
      541: inst = 32'h8220000;
      542: inst = 32'h10408000;
      543: inst = 32'hc40407a;
      544: inst = 32'h8220000;
      545: inst = 32'h10408000;
      546: inst = 32'hc40407b;
      547: inst = 32'h8220000;
      548: inst = 32'h10408000;
      549: inst = 32'hc40407c;
      550: inst = 32'h8220000;
      551: inst = 32'h10408000;
      552: inst = 32'hc40407d;
      553: inst = 32'h8220000;
      554: inst = 32'h10408000;
      555: inst = 32'hc40407e;
      556: inst = 32'h8220000;
      557: inst = 32'h10408000;
      558: inst = 32'hc40407f;
      559: inst = 32'h8220000;
      560: inst = 32'h10408000;
      561: inst = 32'hc404080;
      562: inst = 32'h8220000;
      563: inst = 32'h10408000;
      564: inst = 32'hc404081;
      565: inst = 32'h8220000;
      566: inst = 32'h10408000;
      567: inst = 32'hc404082;
      568: inst = 32'h8220000;
      569: inst = 32'h10408000;
      570: inst = 32'hc404083;
      571: inst = 32'h8220000;
      572: inst = 32'h10408000;
      573: inst = 32'hc404084;
      574: inst = 32'h8220000;
      575: inst = 32'h10408000;
      576: inst = 32'hc404085;
      577: inst = 32'h8220000;
      578: inst = 32'h10408000;
      579: inst = 32'hc404086;
      580: inst = 32'h8220000;
      581: inst = 32'h10408000;
      582: inst = 32'hc404087;
      583: inst = 32'h8220000;
      584: inst = 32'h10408000;
      585: inst = 32'hc404088;
      586: inst = 32'h8220000;
      587: inst = 32'h10408000;
      588: inst = 32'hc404089;
      589: inst = 32'h8220000;
      590: inst = 32'h10408000;
      591: inst = 32'hc40408a;
      592: inst = 32'h8220000;
      593: inst = 32'h10408000;
      594: inst = 32'hc40408b;
      595: inst = 32'h8220000;
      596: inst = 32'h10408000;
      597: inst = 32'hc40408c;
      598: inst = 32'h8220000;
      599: inst = 32'h10408000;
      600: inst = 32'hc40408d;
      601: inst = 32'h8220000;
      602: inst = 32'h10408000;
      603: inst = 32'hc40408e;
      604: inst = 32'h8220000;
      605: inst = 32'h10408000;
      606: inst = 32'hc40408f;
      607: inst = 32'h8220000;
      608: inst = 32'h10408000;
      609: inst = 32'hc404090;
      610: inst = 32'h8220000;
      611: inst = 32'h10408000;
      612: inst = 32'hc404091;
      613: inst = 32'h8220000;
      614: inst = 32'h10408000;
      615: inst = 32'hc404092;
      616: inst = 32'h8220000;
      617: inst = 32'h10408000;
      618: inst = 32'hc404093;
      619: inst = 32'h8220000;
      620: inst = 32'h10408000;
      621: inst = 32'hc404094;
      622: inst = 32'h8220000;
      623: inst = 32'h10408000;
      624: inst = 32'hc404095;
      625: inst = 32'h8220000;
      626: inst = 32'h10408000;
      627: inst = 32'hc404096;
      628: inst = 32'h8220000;
      629: inst = 32'h10408000;
      630: inst = 32'hc404097;
      631: inst = 32'h8220000;
      632: inst = 32'h10408000;
      633: inst = 32'hc404098;
      634: inst = 32'h8220000;
      635: inst = 32'h10408000;
      636: inst = 32'hc404099;
      637: inst = 32'h8220000;
      638: inst = 32'h10408000;
      639: inst = 32'hc40409a;
      640: inst = 32'h8220000;
      641: inst = 32'h10408000;
      642: inst = 32'hc40409b;
      643: inst = 32'h8220000;
      644: inst = 32'h10408000;
      645: inst = 32'hc40409c;
      646: inst = 32'h8220000;
      647: inst = 32'h10408000;
      648: inst = 32'hc40409d;
      649: inst = 32'h8220000;
      650: inst = 32'h10408000;
      651: inst = 32'hc40409e;
      652: inst = 32'h8220000;
      653: inst = 32'h10408000;
      654: inst = 32'hc40409f;
      655: inst = 32'h8220000;
      656: inst = 32'h10408000;
      657: inst = 32'hc4040a0;
      658: inst = 32'h8220000;
      659: inst = 32'h10408000;
      660: inst = 32'hc4040a1;
      661: inst = 32'h8220000;
      662: inst = 32'h10408000;
      663: inst = 32'hc4040a2;
      664: inst = 32'h8220000;
      665: inst = 32'h10408000;
      666: inst = 32'hc4040a3;
      667: inst = 32'h8220000;
      668: inst = 32'h10408000;
      669: inst = 32'hc4040a4;
      670: inst = 32'h8220000;
      671: inst = 32'h10408000;
      672: inst = 32'hc4040a5;
      673: inst = 32'h8220000;
      674: inst = 32'h10408000;
      675: inst = 32'hc4040a6;
      676: inst = 32'h8220000;
      677: inst = 32'h10408000;
      678: inst = 32'hc4040a7;
      679: inst = 32'h8220000;
      680: inst = 32'h10408000;
      681: inst = 32'hc4040a8;
      682: inst = 32'h8220000;
      683: inst = 32'h10408000;
      684: inst = 32'hc4040a9;
      685: inst = 32'h8220000;
      686: inst = 32'h10408000;
      687: inst = 32'hc4040aa;
      688: inst = 32'h8220000;
      689: inst = 32'h10408000;
      690: inst = 32'hc4040ac;
      691: inst = 32'h8220000;
      692: inst = 32'h10408000;
      693: inst = 32'hc4040ad;
      694: inst = 32'h8220000;
      695: inst = 32'h10408000;
      696: inst = 32'hc4040ae;
      697: inst = 32'h8220000;
      698: inst = 32'h10408000;
      699: inst = 32'hc4040af;
      700: inst = 32'h8220000;
      701: inst = 32'h10408000;
      702: inst = 32'hc4040b0;
      703: inst = 32'h8220000;
      704: inst = 32'h10408000;
      705: inst = 32'hc4040b1;
      706: inst = 32'h8220000;
      707: inst = 32'h10408000;
      708: inst = 32'hc4040b2;
      709: inst = 32'h8220000;
      710: inst = 32'h10408000;
      711: inst = 32'hc4040b3;
      712: inst = 32'h8220000;
      713: inst = 32'h10408000;
      714: inst = 32'hc4040b4;
      715: inst = 32'h8220000;
      716: inst = 32'h10408000;
      717: inst = 32'hc4040b5;
      718: inst = 32'h8220000;
      719: inst = 32'h10408000;
      720: inst = 32'hc4040b6;
      721: inst = 32'h8220000;
      722: inst = 32'h10408000;
      723: inst = 32'hc4040b7;
      724: inst = 32'h8220000;
      725: inst = 32'h10408000;
      726: inst = 32'hc4040b8;
      727: inst = 32'h8220000;
      728: inst = 32'h10408000;
      729: inst = 32'hc4040b9;
      730: inst = 32'h8220000;
      731: inst = 32'h10408000;
      732: inst = 32'hc4040ba;
      733: inst = 32'h8220000;
      734: inst = 32'h10408000;
      735: inst = 32'hc4040bb;
      736: inst = 32'h8220000;
      737: inst = 32'h10408000;
      738: inst = 32'hc4040bc;
      739: inst = 32'h8220000;
      740: inst = 32'h10408000;
      741: inst = 32'hc4040bd;
      742: inst = 32'h8220000;
      743: inst = 32'h10408000;
      744: inst = 32'hc4040be;
      745: inst = 32'h8220000;
      746: inst = 32'h10408000;
      747: inst = 32'hc4040bf;
      748: inst = 32'h8220000;
      749: inst = 32'h10408000;
      750: inst = 32'hc4040c0;
      751: inst = 32'h8220000;
      752: inst = 32'h10408000;
      753: inst = 32'hc4040c1;
      754: inst = 32'h8220000;
      755: inst = 32'h10408000;
      756: inst = 32'hc4040c2;
      757: inst = 32'h8220000;
      758: inst = 32'h10408000;
      759: inst = 32'hc4040c3;
      760: inst = 32'h8220000;
      761: inst = 32'h10408000;
      762: inst = 32'hc4040c4;
      763: inst = 32'h8220000;
      764: inst = 32'h10408000;
      765: inst = 32'hc4040c5;
      766: inst = 32'h8220000;
      767: inst = 32'h10408000;
      768: inst = 32'hc4040c6;
      769: inst = 32'h8220000;
      770: inst = 32'h10408000;
      771: inst = 32'hc4040c7;
      772: inst = 32'h8220000;
      773: inst = 32'h10408000;
      774: inst = 32'hc4040c8;
      775: inst = 32'h8220000;
      776: inst = 32'h10408000;
      777: inst = 32'hc4040c9;
      778: inst = 32'h8220000;
      779: inst = 32'h10408000;
      780: inst = 32'hc4040ca;
      781: inst = 32'h8220000;
      782: inst = 32'h10408000;
      783: inst = 32'hc4040cb;
      784: inst = 32'h8220000;
      785: inst = 32'h10408000;
      786: inst = 32'hc4040cc;
      787: inst = 32'h8220000;
      788: inst = 32'h10408000;
      789: inst = 32'hc4040cd;
      790: inst = 32'h8220000;
      791: inst = 32'h10408000;
      792: inst = 32'hc4040ce;
      793: inst = 32'h8220000;
      794: inst = 32'h10408000;
      795: inst = 32'hc4040cf;
      796: inst = 32'h8220000;
      797: inst = 32'h10408000;
      798: inst = 32'hc4040d0;
      799: inst = 32'h8220000;
      800: inst = 32'h10408000;
      801: inst = 32'hc4040d1;
      802: inst = 32'h8220000;
      803: inst = 32'h10408000;
      804: inst = 32'hc4040d2;
      805: inst = 32'h8220000;
      806: inst = 32'h10408000;
      807: inst = 32'hc4040d3;
      808: inst = 32'h8220000;
      809: inst = 32'h10408000;
      810: inst = 32'hc4040d4;
      811: inst = 32'h8220000;
      812: inst = 32'h10408000;
      813: inst = 32'hc4040d5;
      814: inst = 32'h8220000;
      815: inst = 32'h10408000;
      816: inst = 32'hc4040d6;
      817: inst = 32'h8220000;
      818: inst = 32'h10408000;
      819: inst = 32'hc4040d7;
      820: inst = 32'h8220000;
      821: inst = 32'h10408000;
      822: inst = 32'hc4040d8;
      823: inst = 32'h8220000;
      824: inst = 32'h10408000;
      825: inst = 32'hc4040d9;
      826: inst = 32'h8220000;
      827: inst = 32'h10408000;
      828: inst = 32'hc4040da;
      829: inst = 32'h8220000;
      830: inst = 32'h10408000;
      831: inst = 32'hc4040db;
      832: inst = 32'h8220000;
      833: inst = 32'h10408000;
      834: inst = 32'hc4040dc;
      835: inst = 32'h8220000;
      836: inst = 32'h10408000;
      837: inst = 32'hc4040dd;
      838: inst = 32'h8220000;
      839: inst = 32'h10408000;
      840: inst = 32'hc4040de;
      841: inst = 32'h8220000;
      842: inst = 32'h10408000;
      843: inst = 32'hc4040df;
      844: inst = 32'h8220000;
      845: inst = 32'h10408000;
      846: inst = 32'hc4040e0;
      847: inst = 32'h8220000;
      848: inst = 32'h10408000;
      849: inst = 32'hc4040e1;
      850: inst = 32'h8220000;
      851: inst = 32'h10408000;
      852: inst = 32'hc4040e2;
      853: inst = 32'h8220000;
      854: inst = 32'h10408000;
      855: inst = 32'hc4040e3;
      856: inst = 32'h8220000;
      857: inst = 32'h10408000;
      858: inst = 32'hc4040e4;
      859: inst = 32'h8220000;
      860: inst = 32'h10408000;
      861: inst = 32'hc4040e5;
      862: inst = 32'h8220000;
      863: inst = 32'h10408000;
      864: inst = 32'hc4040e6;
      865: inst = 32'h8220000;
      866: inst = 32'h10408000;
      867: inst = 32'hc4040e7;
      868: inst = 32'h8220000;
      869: inst = 32'h10408000;
      870: inst = 32'hc4040e8;
      871: inst = 32'h8220000;
      872: inst = 32'h10408000;
      873: inst = 32'hc4040e9;
      874: inst = 32'h8220000;
      875: inst = 32'h10408000;
      876: inst = 32'hc4040ea;
      877: inst = 32'h8220000;
      878: inst = 32'h10408000;
      879: inst = 32'hc4040eb;
      880: inst = 32'h8220000;
      881: inst = 32'h10408000;
      882: inst = 32'hc4040ec;
      883: inst = 32'h8220000;
      884: inst = 32'h10408000;
      885: inst = 32'hc4040ed;
      886: inst = 32'h8220000;
      887: inst = 32'h10408000;
      888: inst = 32'hc4040ee;
      889: inst = 32'h8220000;
      890: inst = 32'h10408000;
      891: inst = 32'hc4040ef;
      892: inst = 32'h8220000;
      893: inst = 32'h10408000;
      894: inst = 32'hc4040f0;
      895: inst = 32'h8220000;
      896: inst = 32'h10408000;
      897: inst = 32'hc4040f1;
      898: inst = 32'h8220000;
      899: inst = 32'h10408000;
      900: inst = 32'hc4040f2;
      901: inst = 32'h8220000;
      902: inst = 32'h10408000;
      903: inst = 32'hc4040f3;
      904: inst = 32'h8220000;
      905: inst = 32'h10408000;
      906: inst = 32'hc4040f4;
      907: inst = 32'h8220000;
      908: inst = 32'h10408000;
      909: inst = 32'hc4040f5;
      910: inst = 32'h8220000;
      911: inst = 32'h10408000;
      912: inst = 32'hc4040f6;
      913: inst = 32'h8220000;
      914: inst = 32'h10408000;
      915: inst = 32'hc4040f7;
      916: inst = 32'h8220000;
      917: inst = 32'h10408000;
      918: inst = 32'hc4040f8;
      919: inst = 32'h8220000;
      920: inst = 32'h10408000;
      921: inst = 32'hc4040f9;
      922: inst = 32'h8220000;
      923: inst = 32'h10408000;
      924: inst = 32'hc4040fa;
      925: inst = 32'h8220000;
      926: inst = 32'h10408000;
      927: inst = 32'hc4040fb;
      928: inst = 32'h8220000;
      929: inst = 32'h10408000;
      930: inst = 32'hc4040fc;
      931: inst = 32'h8220000;
      932: inst = 32'h10408000;
      933: inst = 32'hc4040fd;
      934: inst = 32'h8220000;
      935: inst = 32'h10408000;
      936: inst = 32'hc4040fe;
      937: inst = 32'h8220000;
      938: inst = 32'h10408000;
      939: inst = 32'hc4040ff;
      940: inst = 32'h8220000;
      941: inst = 32'h10408000;
      942: inst = 32'hc404100;
      943: inst = 32'h8220000;
      944: inst = 32'h10408000;
      945: inst = 32'hc404101;
      946: inst = 32'h8220000;
      947: inst = 32'h10408000;
      948: inst = 32'hc404102;
      949: inst = 32'h8220000;
      950: inst = 32'h10408000;
      951: inst = 32'hc404103;
      952: inst = 32'h8220000;
      953: inst = 32'h10408000;
      954: inst = 32'hc404104;
      955: inst = 32'h8220000;
      956: inst = 32'h10408000;
      957: inst = 32'hc404105;
      958: inst = 32'h8220000;
      959: inst = 32'h10408000;
      960: inst = 32'hc404106;
      961: inst = 32'h8220000;
      962: inst = 32'h10408000;
      963: inst = 32'hc404107;
      964: inst = 32'h8220000;
      965: inst = 32'h10408000;
      966: inst = 32'hc404108;
      967: inst = 32'h8220000;
      968: inst = 32'h10408000;
      969: inst = 32'hc404109;
      970: inst = 32'h8220000;
      971: inst = 32'h10408000;
      972: inst = 32'hc40410a;
      973: inst = 32'h8220000;
      974: inst = 32'h10408000;
      975: inst = 32'hc40410c;
      976: inst = 32'h8220000;
      977: inst = 32'h10408000;
      978: inst = 32'hc40410d;
      979: inst = 32'h8220000;
      980: inst = 32'h10408000;
      981: inst = 32'hc40410e;
      982: inst = 32'h8220000;
      983: inst = 32'h10408000;
      984: inst = 32'hc40410f;
      985: inst = 32'h8220000;
      986: inst = 32'h10408000;
      987: inst = 32'hc404110;
      988: inst = 32'h8220000;
      989: inst = 32'h10408000;
      990: inst = 32'hc404111;
      991: inst = 32'h8220000;
      992: inst = 32'h10408000;
      993: inst = 32'hc404112;
      994: inst = 32'h8220000;
      995: inst = 32'h10408000;
      996: inst = 32'hc404113;
      997: inst = 32'h8220000;
      998: inst = 32'h10408000;
      999: inst = 32'hc404114;
      1000: inst = 32'h8220000;
      1001: inst = 32'h10408000;
      1002: inst = 32'hc404115;
      1003: inst = 32'h8220000;
      1004: inst = 32'h10408000;
      1005: inst = 32'hc404116;
      1006: inst = 32'h8220000;
      1007: inst = 32'h10408000;
      1008: inst = 32'hc404117;
      1009: inst = 32'h8220000;
      1010: inst = 32'h10408000;
      1011: inst = 32'hc404118;
      1012: inst = 32'h8220000;
      1013: inst = 32'h10408000;
      1014: inst = 32'hc404119;
      1015: inst = 32'h8220000;
      1016: inst = 32'h10408000;
      1017: inst = 32'hc40411a;
      1018: inst = 32'h8220000;
      1019: inst = 32'h10408000;
      1020: inst = 32'hc40411b;
      1021: inst = 32'h8220000;
      1022: inst = 32'h10408000;
      1023: inst = 32'hc40411c;
      1024: inst = 32'h8220000;
      1025: inst = 32'h10408000;
      1026: inst = 32'hc40411d;
      1027: inst = 32'h8220000;
      1028: inst = 32'h10408000;
      1029: inst = 32'hc40411e;
      1030: inst = 32'h8220000;
      1031: inst = 32'h10408000;
      1032: inst = 32'hc40411f;
      1033: inst = 32'h8220000;
      1034: inst = 32'h10408000;
      1035: inst = 32'hc404120;
      1036: inst = 32'h8220000;
      1037: inst = 32'h10408000;
      1038: inst = 32'hc404121;
      1039: inst = 32'h8220000;
      1040: inst = 32'h10408000;
      1041: inst = 32'hc404122;
      1042: inst = 32'h8220000;
      1043: inst = 32'h10408000;
      1044: inst = 32'hc404123;
      1045: inst = 32'h8220000;
      1046: inst = 32'h10408000;
      1047: inst = 32'hc404124;
      1048: inst = 32'h8220000;
      1049: inst = 32'h10408000;
      1050: inst = 32'hc404125;
      1051: inst = 32'h8220000;
      1052: inst = 32'h10408000;
      1053: inst = 32'hc404126;
      1054: inst = 32'h8220000;
      1055: inst = 32'h10408000;
      1056: inst = 32'hc404127;
      1057: inst = 32'h8220000;
      1058: inst = 32'h10408000;
      1059: inst = 32'hc404128;
      1060: inst = 32'h8220000;
      1061: inst = 32'h10408000;
      1062: inst = 32'hc404129;
      1063: inst = 32'h8220000;
      1064: inst = 32'h10408000;
      1065: inst = 32'hc40412a;
      1066: inst = 32'h8220000;
      1067: inst = 32'h10408000;
      1068: inst = 32'hc40412b;
      1069: inst = 32'h8220000;
      1070: inst = 32'h10408000;
      1071: inst = 32'hc40412c;
      1072: inst = 32'h8220000;
      1073: inst = 32'h10408000;
      1074: inst = 32'hc40412d;
      1075: inst = 32'h8220000;
      1076: inst = 32'h10408000;
      1077: inst = 32'hc40412e;
      1078: inst = 32'h8220000;
      1079: inst = 32'h10408000;
      1080: inst = 32'hc40412f;
      1081: inst = 32'h8220000;
      1082: inst = 32'h10408000;
      1083: inst = 32'hc404130;
      1084: inst = 32'h8220000;
      1085: inst = 32'h10408000;
      1086: inst = 32'hc404131;
      1087: inst = 32'h8220000;
      1088: inst = 32'h10408000;
      1089: inst = 32'hc404132;
      1090: inst = 32'h8220000;
      1091: inst = 32'h10408000;
      1092: inst = 32'hc404133;
      1093: inst = 32'h8220000;
      1094: inst = 32'h10408000;
      1095: inst = 32'hc404134;
      1096: inst = 32'h8220000;
      1097: inst = 32'h10408000;
      1098: inst = 32'hc404135;
      1099: inst = 32'h8220000;
      1100: inst = 32'h10408000;
      1101: inst = 32'hc404136;
      1102: inst = 32'h8220000;
      1103: inst = 32'h10408000;
      1104: inst = 32'hc404137;
      1105: inst = 32'h8220000;
      1106: inst = 32'h10408000;
      1107: inst = 32'hc404138;
      1108: inst = 32'h8220000;
      1109: inst = 32'h10408000;
      1110: inst = 32'hc404139;
      1111: inst = 32'h8220000;
      1112: inst = 32'h10408000;
      1113: inst = 32'hc40413a;
      1114: inst = 32'h8220000;
      1115: inst = 32'h10408000;
      1116: inst = 32'hc40413b;
      1117: inst = 32'h8220000;
      1118: inst = 32'h10408000;
      1119: inst = 32'hc40413c;
      1120: inst = 32'h8220000;
      1121: inst = 32'h10408000;
      1122: inst = 32'hc40413d;
      1123: inst = 32'h8220000;
      1124: inst = 32'h10408000;
      1125: inst = 32'hc40413e;
      1126: inst = 32'h8220000;
      1127: inst = 32'h10408000;
      1128: inst = 32'hc40413f;
      1129: inst = 32'h8220000;
      1130: inst = 32'h10408000;
      1131: inst = 32'hc404140;
      1132: inst = 32'h8220000;
      1133: inst = 32'h10408000;
      1134: inst = 32'hc404141;
      1135: inst = 32'h8220000;
      1136: inst = 32'h10408000;
      1137: inst = 32'hc404142;
      1138: inst = 32'h8220000;
      1139: inst = 32'h10408000;
      1140: inst = 32'hc404143;
      1141: inst = 32'h8220000;
      1142: inst = 32'h10408000;
      1143: inst = 32'hc404144;
      1144: inst = 32'h8220000;
      1145: inst = 32'h10408000;
      1146: inst = 32'hc404145;
      1147: inst = 32'h8220000;
      1148: inst = 32'h10408000;
      1149: inst = 32'hc404146;
      1150: inst = 32'h8220000;
      1151: inst = 32'h10408000;
      1152: inst = 32'hc404147;
      1153: inst = 32'h8220000;
      1154: inst = 32'h10408000;
      1155: inst = 32'hc404148;
      1156: inst = 32'h8220000;
      1157: inst = 32'h10408000;
      1158: inst = 32'hc404149;
      1159: inst = 32'h8220000;
      1160: inst = 32'h10408000;
      1161: inst = 32'hc40414a;
      1162: inst = 32'h8220000;
      1163: inst = 32'h10408000;
      1164: inst = 32'hc40414b;
      1165: inst = 32'h8220000;
      1166: inst = 32'h10408000;
      1167: inst = 32'hc40414c;
      1168: inst = 32'h8220000;
      1169: inst = 32'h10408000;
      1170: inst = 32'hc40414d;
      1171: inst = 32'h8220000;
      1172: inst = 32'h10408000;
      1173: inst = 32'hc40414e;
      1174: inst = 32'h8220000;
      1175: inst = 32'h10408000;
      1176: inst = 32'hc40414f;
      1177: inst = 32'h8220000;
      1178: inst = 32'h10408000;
      1179: inst = 32'hc404150;
      1180: inst = 32'h8220000;
      1181: inst = 32'h10408000;
      1182: inst = 32'hc404151;
      1183: inst = 32'h8220000;
      1184: inst = 32'h10408000;
      1185: inst = 32'hc404152;
      1186: inst = 32'h8220000;
      1187: inst = 32'h10408000;
      1188: inst = 32'hc404153;
      1189: inst = 32'h8220000;
      1190: inst = 32'h10408000;
      1191: inst = 32'hc404154;
      1192: inst = 32'h8220000;
      1193: inst = 32'h10408000;
      1194: inst = 32'hc404155;
      1195: inst = 32'h8220000;
      1196: inst = 32'h10408000;
      1197: inst = 32'hc404156;
      1198: inst = 32'h8220000;
      1199: inst = 32'h10408000;
      1200: inst = 32'hc404157;
      1201: inst = 32'h8220000;
      1202: inst = 32'h10408000;
      1203: inst = 32'hc404158;
      1204: inst = 32'h8220000;
      1205: inst = 32'h10408000;
      1206: inst = 32'hc404159;
      1207: inst = 32'h8220000;
      1208: inst = 32'h10408000;
      1209: inst = 32'hc40415a;
      1210: inst = 32'h8220000;
      1211: inst = 32'h10408000;
      1212: inst = 32'hc40415b;
      1213: inst = 32'h8220000;
      1214: inst = 32'h10408000;
      1215: inst = 32'hc40415c;
      1216: inst = 32'h8220000;
      1217: inst = 32'h10408000;
      1218: inst = 32'hc40415d;
      1219: inst = 32'h8220000;
      1220: inst = 32'h10408000;
      1221: inst = 32'hc40415e;
      1222: inst = 32'h8220000;
      1223: inst = 32'h10408000;
      1224: inst = 32'hc40415f;
      1225: inst = 32'h8220000;
      1226: inst = 32'h10408000;
      1227: inst = 32'hc404160;
      1228: inst = 32'h8220000;
      1229: inst = 32'h10408000;
      1230: inst = 32'hc404161;
      1231: inst = 32'h8220000;
      1232: inst = 32'h10408000;
      1233: inst = 32'hc404162;
      1234: inst = 32'h8220000;
      1235: inst = 32'h10408000;
      1236: inst = 32'hc404163;
      1237: inst = 32'h8220000;
      1238: inst = 32'h10408000;
      1239: inst = 32'hc404164;
      1240: inst = 32'h8220000;
      1241: inst = 32'h10408000;
      1242: inst = 32'hc404165;
      1243: inst = 32'h8220000;
      1244: inst = 32'h10408000;
      1245: inst = 32'hc404166;
      1246: inst = 32'h8220000;
      1247: inst = 32'h10408000;
      1248: inst = 32'hc404167;
      1249: inst = 32'h8220000;
      1250: inst = 32'h10408000;
      1251: inst = 32'hc404168;
      1252: inst = 32'h8220000;
      1253: inst = 32'h10408000;
      1254: inst = 32'hc404169;
      1255: inst = 32'h8220000;
      1256: inst = 32'h10408000;
      1257: inst = 32'hc40416a;
      1258: inst = 32'h8220000;
      1259: inst = 32'h10408000;
      1260: inst = 32'hc40416c;
      1261: inst = 32'h8220000;
      1262: inst = 32'h10408000;
      1263: inst = 32'hc40416d;
      1264: inst = 32'h8220000;
      1265: inst = 32'h10408000;
      1266: inst = 32'hc40416e;
      1267: inst = 32'h8220000;
      1268: inst = 32'h10408000;
      1269: inst = 32'hc40416f;
      1270: inst = 32'h8220000;
      1271: inst = 32'h10408000;
      1272: inst = 32'hc404170;
      1273: inst = 32'h8220000;
      1274: inst = 32'h10408000;
      1275: inst = 32'hc404171;
      1276: inst = 32'h8220000;
      1277: inst = 32'h10408000;
      1278: inst = 32'hc404172;
      1279: inst = 32'h8220000;
      1280: inst = 32'h10408000;
      1281: inst = 32'hc404173;
      1282: inst = 32'h8220000;
      1283: inst = 32'h10408000;
      1284: inst = 32'hc404174;
      1285: inst = 32'h8220000;
      1286: inst = 32'h10408000;
      1287: inst = 32'hc404175;
      1288: inst = 32'h8220000;
      1289: inst = 32'h10408000;
      1290: inst = 32'hc404176;
      1291: inst = 32'h8220000;
      1292: inst = 32'h10408000;
      1293: inst = 32'hc404177;
      1294: inst = 32'h8220000;
      1295: inst = 32'h10408000;
      1296: inst = 32'hc404178;
      1297: inst = 32'h8220000;
      1298: inst = 32'h10408000;
      1299: inst = 32'hc404179;
      1300: inst = 32'h8220000;
      1301: inst = 32'h10408000;
      1302: inst = 32'hc40417a;
      1303: inst = 32'h8220000;
      1304: inst = 32'h10408000;
      1305: inst = 32'hc40417b;
      1306: inst = 32'h8220000;
      1307: inst = 32'h10408000;
      1308: inst = 32'hc40417c;
      1309: inst = 32'h8220000;
      1310: inst = 32'h10408000;
      1311: inst = 32'hc40417d;
      1312: inst = 32'h8220000;
      1313: inst = 32'h10408000;
      1314: inst = 32'hc40417e;
      1315: inst = 32'h8220000;
      1316: inst = 32'h10408000;
      1317: inst = 32'hc40417f;
      1318: inst = 32'h8220000;
      1319: inst = 32'h10408000;
      1320: inst = 32'hc404180;
      1321: inst = 32'h8220000;
      1322: inst = 32'h10408000;
      1323: inst = 32'hc404181;
      1324: inst = 32'h8220000;
      1325: inst = 32'h10408000;
      1326: inst = 32'hc404182;
      1327: inst = 32'h8220000;
      1328: inst = 32'h10408000;
      1329: inst = 32'hc404183;
      1330: inst = 32'h8220000;
      1331: inst = 32'h10408000;
      1332: inst = 32'hc404184;
      1333: inst = 32'h8220000;
      1334: inst = 32'h10408000;
      1335: inst = 32'hc404185;
      1336: inst = 32'h8220000;
      1337: inst = 32'h10408000;
      1338: inst = 32'hc404186;
      1339: inst = 32'h8220000;
      1340: inst = 32'h10408000;
      1341: inst = 32'hc404187;
      1342: inst = 32'h8220000;
      1343: inst = 32'h10408000;
      1344: inst = 32'hc404188;
      1345: inst = 32'h8220000;
      1346: inst = 32'h10408000;
      1347: inst = 32'hc404189;
      1348: inst = 32'h8220000;
      1349: inst = 32'h10408000;
      1350: inst = 32'hc40418a;
      1351: inst = 32'h8220000;
      1352: inst = 32'h10408000;
      1353: inst = 32'hc40418b;
      1354: inst = 32'h8220000;
      1355: inst = 32'h10408000;
      1356: inst = 32'hc40418c;
      1357: inst = 32'h8220000;
      1358: inst = 32'h10408000;
      1359: inst = 32'hc40418d;
      1360: inst = 32'h8220000;
      1361: inst = 32'h10408000;
      1362: inst = 32'hc40418e;
      1363: inst = 32'h8220000;
      1364: inst = 32'h10408000;
      1365: inst = 32'hc40418f;
      1366: inst = 32'h8220000;
      1367: inst = 32'h10408000;
      1368: inst = 32'hc404190;
      1369: inst = 32'h8220000;
      1370: inst = 32'h10408000;
      1371: inst = 32'hc404191;
      1372: inst = 32'h8220000;
      1373: inst = 32'h10408000;
      1374: inst = 32'hc404192;
      1375: inst = 32'h8220000;
      1376: inst = 32'h10408000;
      1377: inst = 32'hc404193;
      1378: inst = 32'h8220000;
      1379: inst = 32'h10408000;
      1380: inst = 32'hc404194;
      1381: inst = 32'h8220000;
      1382: inst = 32'h10408000;
      1383: inst = 32'hc404195;
      1384: inst = 32'h8220000;
      1385: inst = 32'h10408000;
      1386: inst = 32'hc404196;
      1387: inst = 32'h8220000;
      1388: inst = 32'h10408000;
      1389: inst = 32'hc404197;
      1390: inst = 32'h8220000;
      1391: inst = 32'h10408000;
      1392: inst = 32'hc404198;
      1393: inst = 32'h8220000;
      1394: inst = 32'h10408000;
      1395: inst = 32'hc404199;
      1396: inst = 32'h8220000;
      1397: inst = 32'h10408000;
      1398: inst = 32'hc40419a;
      1399: inst = 32'h8220000;
      1400: inst = 32'h10408000;
      1401: inst = 32'hc40419b;
      1402: inst = 32'h8220000;
      1403: inst = 32'h10408000;
      1404: inst = 32'hc40419c;
      1405: inst = 32'h8220000;
      1406: inst = 32'h10408000;
      1407: inst = 32'hc40419d;
      1408: inst = 32'h8220000;
      1409: inst = 32'h10408000;
      1410: inst = 32'hc40419e;
      1411: inst = 32'h8220000;
      1412: inst = 32'h10408000;
      1413: inst = 32'hc40419f;
      1414: inst = 32'h8220000;
      1415: inst = 32'h10408000;
      1416: inst = 32'hc4041a0;
      1417: inst = 32'h8220000;
      1418: inst = 32'h10408000;
      1419: inst = 32'hc4041a1;
      1420: inst = 32'h8220000;
      1421: inst = 32'h10408000;
      1422: inst = 32'hc4041a2;
      1423: inst = 32'h8220000;
      1424: inst = 32'h10408000;
      1425: inst = 32'hc4041a3;
      1426: inst = 32'h8220000;
      1427: inst = 32'h10408000;
      1428: inst = 32'hc4041a4;
      1429: inst = 32'h8220000;
      1430: inst = 32'h10408000;
      1431: inst = 32'hc4041a5;
      1432: inst = 32'h8220000;
      1433: inst = 32'h10408000;
      1434: inst = 32'hc4041a6;
      1435: inst = 32'h8220000;
      1436: inst = 32'h10408000;
      1437: inst = 32'hc4041a7;
      1438: inst = 32'h8220000;
      1439: inst = 32'h10408000;
      1440: inst = 32'hc4041a8;
      1441: inst = 32'h8220000;
      1442: inst = 32'h10408000;
      1443: inst = 32'hc4041a9;
      1444: inst = 32'h8220000;
      1445: inst = 32'h10408000;
      1446: inst = 32'hc4041aa;
      1447: inst = 32'h8220000;
      1448: inst = 32'h10408000;
      1449: inst = 32'hc4041ab;
      1450: inst = 32'h8220000;
      1451: inst = 32'h10408000;
      1452: inst = 32'hc4041ac;
      1453: inst = 32'h8220000;
      1454: inst = 32'h10408000;
      1455: inst = 32'hc4041ad;
      1456: inst = 32'h8220000;
      1457: inst = 32'h10408000;
      1458: inst = 32'hc4041ae;
      1459: inst = 32'h8220000;
      1460: inst = 32'h10408000;
      1461: inst = 32'hc4041af;
      1462: inst = 32'h8220000;
      1463: inst = 32'h10408000;
      1464: inst = 32'hc4041b0;
      1465: inst = 32'h8220000;
      1466: inst = 32'h10408000;
      1467: inst = 32'hc4041b1;
      1468: inst = 32'h8220000;
      1469: inst = 32'h10408000;
      1470: inst = 32'hc4041b2;
      1471: inst = 32'h8220000;
      1472: inst = 32'h10408000;
      1473: inst = 32'hc4041b3;
      1474: inst = 32'h8220000;
      1475: inst = 32'h10408000;
      1476: inst = 32'hc4041b4;
      1477: inst = 32'h8220000;
      1478: inst = 32'h10408000;
      1479: inst = 32'hc4041b5;
      1480: inst = 32'h8220000;
      1481: inst = 32'h10408000;
      1482: inst = 32'hc4041b6;
      1483: inst = 32'h8220000;
      1484: inst = 32'h10408000;
      1485: inst = 32'hc4041b7;
      1486: inst = 32'h8220000;
      1487: inst = 32'h10408000;
      1488: inst = 32'hc4041b8;
      1489: inst = 32'h8220000;
      1490: inst = 32'h10408000;
      1491: inst = 32'hc4041b9;
      1492: inst = 32'h8220000;
      1493: inst = 32'h10408000;
      1494: inst = 32'hc4041ba;
      1495: inst = 32'h8220000;
      1496: inst = 32'h10408000;
      1497: inst = 32'hc4041bb;
      1498: inst = 32'h8220000;
      1499: inst = 32'h10408000;
      1500: inst = 32'hc4041bc;
      1501: inst = 32'h8220000;
      1502: inst = 32'h10408000;
      1503: inst = 32'hc4041bd;
      1504: inst = 32'h8220000;
      1505: inst = 32'h10408000;
      1506: inst = 32'hc4041be;
      1507: inst = 32'h8220000;
      1508: inst = 32'h10408000;
      1509: inst = 32'hc4041bf;
      1510: inst = 32'h8220000;
      1511: inst = 32'h10408000;
      1512: inst = 32'hc4041c0;
      1513: inst = 32'h8220000;
      1514: inst = 32'h10408000;
      1515: inst = 32'hc4041c1;
      1516: inst = 32'h8220000;
      1517: inst = 32'h10408000;
      1518: inst = 32'hc4041c2;
      1519: inst = 32'h8220000;
      1520: inst = 32'h10408000;
      1521: inst = 32'hc4041c3;
      1522: inst = 32'h8220000;
      1523: inst = 32'h10408000;
      1524: inst = 32'hc4041c4;
      1525: inst = 32'h8220000;
      1526: inst = 32'h10408000;
      1527: inst = 32'hc4041c5;
      1528: inst = 32'h8220000;
      1529: inst = 32'h10408000;
      1530: inst = 32'hc4041c6;
      1531: inst = 32'h8220000;
      1532: inst = 32'h10408000;
      1533: inst = 32'hc4041c7;
      1534: inst = 32'h8220000;
      1535: inst = 32'h10408000;
      1536: inst = 32'hc4041c8;
      1537: inst = 32'h8220000;
      1538: inst = 32'h10408000;
      1539: inst = 32'hc4041c9;
      1540: inst = 32'h8220000;
      1541: inst = 32'h10408000;
      1542: inst = 32'hc4041ca;
      1543: inst = 32'h8220000;
      1544: inst = 32'h10408000;
      1545: inst = 32'hc4041cc;
      1546: inst = 32'h8220000;
      1547: inst = 32'h10408000;
      1548: inst = 32'hc4041cd;
      1549: inst = 32'h8220000;
      1550: inst = 32'h10408000;
      1551: inst = 32'hc4041ce;
      1552: inst = 32'h8220000;
      1553: inst = 32'h10408000;
      1554: inst = 32'hc4041cf;
      1555: inst = 32'h8220000;
      1556: inst = 32'h10408000;
      1557: inst = 32'hc4041d0;
      1558: inst = 32'h8220000;
      1559: inst = 32'h10408000;
      1560: inst = 32'hc4041d1;
      1561: inst = 32'h8220000;
      1562: inst = 32'h10408000;
      1563: inst = 32'hc4041d2;
      1564: inst = 32'h8220000;
      1565: inst = 32'h10408000;
      1566: inst = 32'hc4041d3;
      1567: inst = 32'h8220000;
      1568: inst = 32'h10408000;
      1569: inst = 32'hc4041d4;
      1570: inst = 32'h8220000;
      1571: inst = 32'h10408000;
      1572: inst = 32'hc4041d5;
      1573: inst = 32'h8220000;
      1574: inst = 32'h10408000;
      1575: inst = 32'hc4041d6;
      1576: inst = 32'h8220000;
      1577: inst = 32'h10408000;
      1578: inst = 32'hc4041d7;
      1579: inst = 32'h8220000;
      1580: inst = 32'h10408000;
      1581: inst = 32'hc4041d8;
      1582: inst = 32'h8220000;
      1583: inst = 32'h10408000;
      1584: inst = 32'hc4041d9;
      1585: inst = 32'h8220000;
      1586: inst = 32'h10408000;
      1587: inst = 32'hc404206;
      1588: inst = 32'h8220000;
      1589: inst = 32'h10408000;
      1590: inst = 32'hc404207;
      1591: inst = 32'h8220000;
      1592: inst = 32'h10408000;
      1593: inst = 32'hc404208;
      1594: inst = 32'h8220000;
      1595: inst = 32'h10408000;
      1596: inst = 32'hc404209;
      1597: inst = 32'h8220000;
      1598: inst = 32'h10408000;
      1599: inst = 32'hc40420a;
      1600: inst = 32'h8220000;
      1601: inst = 32'h10408000;
      1602: inst = 32'hc40420b;
      1603: inst = 32'h8220000;
      1604: inst = 32'h10408000;
      1605: inst = 32'hc40420c;
      1606: inst = 32'h8220000;
      1607: inst = 32'h10408000;
      1608: inst = 32'hc40420d;
      1609: inst = 32'h8220000;
      1610: inst = 32'h10408000;
      1611: inst = 32'hc40420e;
      1612: inst = 32'h8220000;
      1613: inst = 32'h10408000;
      1614: inst = 32'hc40420f;
      1615: inst = 32'h8220000;
      1616: inst = 32'h10408000;
      1617: inst = 32'hc404210;
      1618: inst = 32'h8220000;
      1619: inst = 32'h10408000;
      1620: inst = 32'hc404211;
      1621: inst = 32'h8220000;
      1622: inst = 32'h10408000;
      1623: inst = 32'hc404212;
      1624: inst = 32'h8220000;
      1625: inst = 32'h10408000;
      1626: inst = 32'hc404213;
      1627: inst = 32'h8220000;
      1628: inst = 32'h10408000;
      1629: inst = 32'hc404214;
      1630: inst = 32'h8220000;
      1631: inst = 32'h10408000;
      1632: inst = 32'hc404215;
      1633: inst = 32'h8220000;
      1634: inst = 32'h10408000;
      1635: inst = 32'hc404216;
      1636: inst = 32'h8220000;
      1637: inst = 32'h10408000;
      1638: inst = 32'hc404217;
      1639: inst = 32'h8220000;
      1640: inst = 32'h10408000;
      1641: inst = 32'hc404218;
      1642: inst = 32'h8220000;
      1643: inst = 32'h10408000;
      1644: inst = 32'hc404219;
      1645: inst = 32'h8220000;
      1646: inst = 32'h10408000;
      1647: inst = 32'hc40421a;
      1648: inst = 32'h8220000;
      1649: inst = 32'h10408000;
      1650: inst = 32'hc40421b;
      1651: inst = 32'h8220000;
      1652: inst = 32'h10408000;
      1653: inst = 32'hc40421c;
      1654: inst = 32'h8220000;
      1655: inst = 32'h10408000;
      1656: inst = 32'hc40421d;
      1657: inst = 32'h8220000;
      1658: inst = 32'h10408000;
      1659: inst = 32'hc40421e;
      1660: inst = 32'h8220000;
      1661: inst = 32'h10408000;
      1662: inst = 32'hc40421f;
      1663: inst = 32'h8220000;
      1664: inst = 32'h10408000;
      1665: inst = 32'hc404220;
      1666: inst = 32'h8220000;
      1667: inst = 32'h10408000;
      1668: inst = 32'hc404221;
      1669: inst = 32'h8220000;
      1670: inst = 32'h10408000;
      1671: inst = 32'hc404222;
      1672: inst = 32'h8220000;
      1673: inst = 32'h10408000;
      1674: inst = 32'hc404223;
      1675: inst = 32'h8220000;
      1676: inst = 32'h10408000;
      1677: inst = 32'hc404224;
      1678: inst = 32'h8220000;
      1679: inst = 32'h10408000;
      1680: inst = 32'hc404225;
      1681: inst = 32'h8220000;
      1682: inst = 32'h10408000;
      1683: inst = 32'hc404226;
      1684: inst = 32'h8220000;
      1685: inst = 32'h10408000;
      1686: inst = 32'hc404227;
      1687: inst = 32'h8220000;
      1688: inst = 32'h10408000;
      1689: inst = 32'hc404228;
      1690: inst = 32'h8220000;
      1691: inst = 32'h10408000;
      1692: inst = 32'hc404229;
      1693: inst = 32'h8220000;
      1694: inst = 32'h10408000;
      1695: inst = 32'hc40422a;
      1696: inst = 32'h8220000;
      1697: inst = 32'h10408000;
      1698: inst = 32'hc40422c;
      1699: inst = 32'h8220000;
      1700: inst = 32'h10408000;
      1701: inst = 32'hc40422d;
      1702: inst = 32'h8220000;
      1703: inst = 32'h10408000;
      1704: inst = 32'hc40422e;
      1705: inst = 32'h8220000;
      1706: inst = 32'h10408000;
      1707: inst = 32'hc40422f;
      1708: inst = 32'h8220000;
      1709: inst = 32'h10408000;
      1710: inst = 32'hc404230;
      1711: inst = 32'h8220000;
      1712: inst = 32'h10408000;
      1713: inst = 32'hc404231;
      1714: inst = 32'h8220000;
      1715: inst = 32'h10408000;
      1716: inst = 32'hc404232;
      1717: inst = 32'h8220000;
      1718: inst = 32'h10408000;
      1719: inst = 32'hc404233;
      1720: inst = 32'h8220000;
      1721: inst = 32'h10408000;
      1722: inst = 32'hc404234;
      1723: inst = 32'h8220000;
      1724: inst = 32'h10408000;
      1725: inst = 32'hc404235;
      1726: inst = 32'h8220000;
      1727: inst = 32'h10408000;
      1728: inst = 32'hc404236;
      1729: inst = 32'h8220000;
      1730: inst = 32'h10408000;
      1731: inst = 32'hc404237;
      1732: inst = 32'h8220000;
      1733: inst = 32'h10408000;
      1734: inst = 32'hc404238;
      1735: inst = 32'h8220000;
      1736: inst = 32'h10408000;
      1737: inst = 32'hc404239;
      1738: inst = 32'h8220000;
      1739: inst = 32'h10408000;
      1740: inst = 32'hc40423a;
      1741: inst = 32'h8220000;
      1742: inst = 32'h10408000;
      1743: inst = 32'hc40423b;
      1744: inst = 32'h8220000;
      1745: inst = 32'h10408000;
      1746: inst = 32'hc404264;
      1747: inst = 32'h8220000;
      1748: inst = 32'h10408000;
      1749: inst = 32'hc404265;
      1750: inst = 32'h8220000;
      1751: inst = 32'h10408000;
      1752: inst = 32'hc404266;
      1753: inst = 32'h8220000;
      1754: inst = 32'h10408000;
      1755: inst = 32'hc404267;
      1756: inst = 32'h8220000;
      1757: inst = 32'h10408000;
      1758: inst = 32'hc404268;
      1759: inst = 32'h8220000;
      1760: inst = 32'h10408000;
      1761: inst = 32'hc404269;
      1762: inst = 32'h8220000;
      1763: inst = 32'h10408000;
      1764: inst = 32'hc40426a;
      1765: inst = 32'h8220000;
      1766: inst = 32'h10408000;
      1767: inst = 32'hc40426b;
      1768: inst = 32'h8220000;
      1769: inst = 32'h10408000;
      1770: inst = 32'hc40426c;
      1771: inst = 32'h8220000;
      1772: inst = 32'h10408000;
      1773: inst = 32'hc40426d;
      1774: inst = 32'h8220000;
      1775: inst = 32'h10408000;
      1776: inst = 32'hc40426e;
      1777: inst = 32'h8220000;
      1778: inst = 32'h10408000;
      1779: inst = 32'hc40426f;
      1780: inst = 32'h8220000;
      1781: inst = 32'h10408000;
      1782: inst = 32'hc404270;
      1783: inst = 32'h8220000;
      1784: inst = 32'h10408000;
      1785: inst = 32'hc404271;
      1786: inst = 32'h8220000;
      1787: inst = 32'h10408000;
      1788: inst = 32'hc404272;
      1789: inst = 32'h8220000;
      1790: inst = 32'h10408000;
      1791: inst = 32'hc404273;
      1792: inst = 32'h8220000;
      1793: inst = 32'h10408000;
      1794: inst = 32'hc404274;
      1795: inst = 32'h8220000;
      1796: inst = 32'h10408000;
      1797: inst = 32'hc404275;
      1798: inst = 32'h8220000;
      1799: inst = 32'h10408000;
      1800: inst = 32'hc404276;
      1801: inst = 32'h8220000;
      1802: inst = 32'h10408000;
      1803: inst = 32'hc404277;
      1804: inst = 32'h8220000;
      1805: inst = 32'h10408000;
      1806: inst = 32'hc404278;
      1807: inst = 32'h8220000;
      1808: inst = 32'h10408000;
      1809: inst = 32'hc404279;
      1810: inst = 32'h8220000;
      1811: inst = 32'h10408000;
      1812: inst = 32'hc40427a;
      1813: inst = 32'h8220000;
      1814: inst = 32'h10408000;
      1815: inst = 32'hc40427b;
      1816: inst = 32'h8220000;
      1817: inst = 32'h10408000;
      1818: inst = 32'hc40427c;
      1819: inst = 32'h8220000;
      1820: inst = 32'h10408000;
      1821: inst = 32'hc40427d;
      1822: inst = 32'h8220000;
      1823: inst = 32'h10408000;
      1824: inst = 32'hc40427e;
      1825: inst = 32'h8220000;
      1826: inst = 32'h10408000;
      1827: inst = 32'hc40427f;
      1828: inst = 32'h8220000;
      1829: inst = 32'h10408000;
      1830: inst = 32'hc404280;
      1831: inst = 32'h8220000;
      1832: inst = 32'h10408000;
      1833: inst = 32'hc404281;
      1834: inst = 32'h8220000;
      1835: inst = 32'h10408000;
      1836: inst = 32'hc404282;
      1837: inst = 32'h8220000;
      1838: inst = 32'h10408000;
      1839: inst = 32'hc404283;
      1840: inst = 32'h8220000;
      1841: inst = 32'h10408000;
      1842: inst = 32'hc404284;
      1843: inst = 32'h8220000;
      1844: inst = 32'h10408000;
      1845: inst = 32'hc404285;
      1846: inst = 32'h8220000;
      1847: inst = 32'h10408000;
      1848: inst = 32'hc404286;
      1849: inst = 32'h8220000;
      1850: inst = 32'h10408000;
      1851: inst = 32'hc404287;
      1852: inst = 32'h8220000;
      1853: inst = 32'h10408000;
      1854: inst = 32'hc404288;
      1855: inst = 32'h8220000;
      1856: inst = 32'h10408000;
      1857: inst = 32'hc404289;
      1858: inst = 32'h8220000;
      1859: inst = 32'h10408000;
      1860: inst = 32'hc40428a;
      1861: inst = 32'h8220000;
      1862: inst = 32'h10408000;
      1863: inst = 32'hc40428c;
      1864: inst = 32'h8220000;
      1865: inst = 32'h10408000;
      1866: inst = 32'hc40428d;
      1867: inst = 32'h8220000;
      1868: inst = 32'h10408000;
      1869: inst = 32'hc40428e;
      1870: inst = 32'h8220000;
      1871: inst = 32'h10408000;
      1872: inst = 32'hc40428f;
      1873: inst = 32'h8220000;
      1874: inst = 32'h10408000;
      1875: inst = 32'hc404290;
      1876: inst = 32'h8220000;
      1877: inst = 32'h10408000;
      1878: inst = 32'hc404291;
      1879: inst = 32'h8220000;
      1880: inst = 32'h10408000;
      1881: inst = 32'hc404292;
      1882: inst = 32'h8220000;
      1883: inst = 32'h10408000;
      1884: inst = 32'hc404293;
      1885: inst = 32'h8220000;
      1886: inst = 32'h10408000;
      1887: inst = 32'hc404294;
      1888: inst = 32'h8220000;
      1889: inst = 32'h10408000;
      1890: inst = 32'hc404295;
      1891: inst = 32'h8220000;
      1892: inst = 32'h10408000;
      1893: inst = 32'hc404296;
      1894: inst = 32'h8220000;
      1895: inst = 32'h10408000;
      1896: inst = 32'hc404297;
      1897: inst = 32'h8220000;
      1898: inst = 32'h10408000;
      1899: inst = 32'hc404298;
      1900: inst = 32'h8220000;
      1901: inst = 32'h10408000;
      1902: inst = 32'hc404299;
      1903: inst = 32'h8220000;
      1904: inst = 32'h10408000;
      1905: inst = 32'hc40429a;
      1906: inst = 32'h8220000;
      1907: inst = 32'h10408000;
      1908: inst = 32'hc40429b;
      1909: inst = 32'h8220000;
      1910: inst = 32'h10408000;
      1911: inst = 32'hc4042c4;
      1912: inst = 32'h8220000;
      1913: inst = 32'h10408000;
      1914: inst = 32'hc4042c5;
      1915: inst = 32'h8220000;
      1916: inst = 32'h10408000;
      1917: inst = 32'hc4042c6;
      1918: inst = 32'h8220000;
      1919: inst = 32'h10408000;
      1920: inst = 32'hc4042c7;
      1921: inst = 32'h8220000;
      1922: inst = 32'h10408000;
      1923: inst = 32'hc4042c8;
      1924: inst = 32'h8220000;
      1925: inst = 32'h10408000;
      1926: inst = 32'hc4042c9;
      1927: inst = 32'h8220000;
      1928: inst = 32'h10408000;
      1929: inst = 32'hc4042ca;
      1930: inst = 32'h8220000;
      1931: inst = 32'h10408000;
      1932: inst = 32'hc4042cb;
      1933: inst = 32'h8220000;
      1934: inst = 32'h10408000;
      1935: inst = 32'hc4042cc;
      1936: inst = 32'h8220000;
      1937: inst = 32'h10408000;
      1938: inst = 32'hc4042cd;
      1939: inst = 32'h8220000;
      1940: inst = 32'h10408000;
      1941: inst = 32'hc4042ce;
      1942: inst = 32'h8220000;
      1943: inst = 32'h10408000;
      1944: inst = 32'hc4042cf;
      1945: inst = 32'h8220000;
      1946: inst = 32'h10408000;
      1947: inst = 32'hc4042d0;
      1948: inst = 32'h8220000;
      1949: inst = 32'h10408000;
      1950: inst = 32'hc4042d1;
      1951: inst = 32'h8220000;
      1952: inst = 32'h10408000;
      1953: inst = 32'hc4042d2;
      1954: inst = 32'h8220000;
      1955: inst = 32'h10408000;
      1956: inst = 32'hc4042d3;
      1957: inst = 32'h8220000;
      1958: inst = 32'h10408000;
      1959: inst = 32'hc4042d4;
      1960: inst = 32'h8220000;
      1961: inst = 32'h10408000;
      1962: inst = 32'hc4042d5;
      1963: inst = 32'h8220000;
      1964: inst = 32'h10408000;
      1965: inst = 32'hc4042d6;
      1966: inst = 32'h8220000;
      1967: inst = 32'h10408000;
      1968: inst = 32'hc4042d7;
      1969: inst = 32'h8220000;
      1970: inst = 32'h10408000;
      1971: inst = 32'hc4042d8;
      1972: inst = 32'h8220000;
      1973: inst = 32'h10408000;
      1974: inst = 32'hc4042d9;
      1975: inst = 32'h8220000;
      1976: inst = 32'h10408000;
      1977: inst = 32'hc4042da;
      1978: inst = 32'h8220000;
      1979: inst = 32'h10408000;
      1980: inst = 32'hc4042db;
      1981: inst = 32'h8220000;
      1982: inst = 32'h10408000;
      1983: inst = 32'hc4042dc;
      1984: inst = 32'h8220000;
      1985: inst = 32'h10408000;
      1986: inst = 32'hc4042dd;
      1987: inst = 32'h8220000;
      1988: inst = 32'h10408000;
      1989: inst = 32'hc4042de;
      1990: inst = 32'h8220000;
      1991: inst = 32'h10408000;
      1992: inst = 32'hc4042df;
      1993: inst = 32'h8220000;
      1994: inst = 32'h10408000;
      1995: inst = 32'hc4042e0;
      1996: inst = 32'h8220000;
      1997: inst = 32'h10408000;
      1998: inst = 32'hc4042e1;
      1999: inst = 32'h8220000;
      2000: inst = 32'h10408000;
      2001: inst = 32'hc4042e2;
      2002: inst = 32'h8220000;
      2003: inst = 32'h10408000;
      2004: inst = 32'hc4042e3;
      2005: inst = 32'h8220000;
      2006: inst = 32'h10408000;
      2007: inst = 32'hc4042e4;
      2008: inst = 32'h8220000;
      2009: inst = 32'h10408000;
      2010: inst = 32'hc4042e5;
      2011: inst = 32'h8220000;
      2012: inst = 32'h10408000;
      2013: inst = 32'hc4042e6;
      2014: inst = 32'h8220000;
      2015: inst = 32'h10408000;
      2016: inst = 32'hc4042e7;
      2017: inst = 32'h8220000;
      2018: inst = 32'h10408000;
      2019: inst = 32'hc4042e8;
      2020: inst = 32'h8220000;
      2021: inst = 32'h10408000;
      2022: inst = 32'hc4042e9;
      2023: inst = 32'h8220000;
      2024: inst = 32'h10408000;
      2025: inst = 32'hc4042ee;
      2026: inst = 32'h8220000;
      2027: inst = 32'h10408000;
      2028: inst = 32'hc4042ef;
      2029: inst = 32'h8220000;
      2030: inst = 32'h10408000;
      2031: inst = 32'hc4042f0;
      2032: inst = 32'h8220000;
      2033: inst = 32'h10408000;
      2034: inst = 32'hc4042f1;
      2035: inst = 32'h8220000;
      2036: inst = 32'h10408000;
      2037: inst = 32'hc4042f2;
      2038: inst = 32'h8220000;
      2039: inst = 32'h10408000;
      2040: inst = 32'hc4042f3;
      2041: inst = 32'h8220000;
      2042: inst = 32'h10408000;
      2043: inst = 32'hc4042f4;
      2044: inst = 32'h8220000;
      2045: inst = 32'h10408000;
      2046: inst = 32'hc4042f5;
      2047: inst = 32'h8220000;
      2048: inst = 32'h10408000;
      2049: inst = 32'hc4042f6;
      2050: inst = 32'h8220000;
      2051: inst = 32'h10408000;
      2052: inst = 32'hc4042f7;
      2053: inst = 32'h8220000;
      2054: inst = 32'h10408000;
      2055: inst = 32'hc4042f8;
      2056: inst = 32'h8220000;
      2057: inst = 32'h10408000;
      2058: inst = 32'hc4042f9;
      2059: inst = 32'h8220000;
      2060: inst = 32'h10408000;
      2061: inst = 32'hc4042fa;
      2062: inst = 32'h8220000;
      2063: inst = 32'h10408000;
      2064: inst = 32'hc4042fb;
      2065: inst = 32'h8220000;
      2066: inst = 32'h10408000;
      2067: inst = 32'hc404324;
      2068: inst = 32'h8220000;
      2069: inst = 32'h10408000;
      2070: inst = 32'hc404325;
      2071: inst = 32'h8220000;
      2072: inst = 32'h10408000;
      2073: inst = 32'hc404326;
      2074: inst = 32'h8220000;
      2075: inst = 32'h10408000;
      2076: inst = 32'hc404327;
      2077: inst = 32'h8220000;
      2078: inst = 32'h10408000;
      2079: inst = 32'hc404328;
      2080: inst = 32'h8220000;
      2081: inst = 32'h10408000;
      2082: inst = 32'hc404329;
      2083: inst = 32'h8220000;
      2084: inst = 32'h10408000;
      2085: inst = 32'hc40432a;
      2086: inst = 32'h8220000;
      2087: inst = 32'h10408000;
      2088: inst = 32'hc40432b;
      2089: inst = 32'h8220000;
      2090: inst = 32'h10408000;
      2091: inst = 32'hc40432c;
      2092: inst = 32'h8220000;
      2093: inst = 32'h10408000;
      2094: inst = 32'hc40432d;
      2095: inst = 32'h8220000;
      2096: inst = 32'h10408000;
      2097: inst = 32'hc40432e;
      2098: inst = 32'h8220000;
      2099: inst = 32'h10408000;
      2100: inst = 32'hc40432f;
      2101: inst = 32'h8220000;
      2102: inst = 32'h10408000;
      2103: inst = 32'hc404330;
      2104: inst = 32'h8220000;
      2105: inst = 32'h10408000;
      2106: inst = 32'hc404331;
      2107: inst = 32'h8220000;
      2108: inst = 32'h10408000;
      2109: inst = 32'hc404332;
      2110: inst = 32'h8220000;
      2111: inst = 32'h10408000;
      2112: inst = 32'hc404333;
      2113: inst = 32'h8220000;
      2114: inst = 32'h10408000;
      2115: inst = 32'hc404334;
      2116: inst = 32'h8220000;
      2117: inst = 32'h10408000;
      2118: inst = 32'hc404335;
      2119: inst = 32'h8220000;
      2120: inst = 32'h10408000;
      2121: inst = 32'hc404336;
      2122: inst = 32'h8220000;
      2123: inst = 32'h10408000;
      2124: inst = 32'hc404337;
      2125: inst = 32'h8220000;
      2126: inst = 32'h10408000;
      2127: inst = 32'hc404338;
      2128: inst = 32'h8220000;
      2129: inst = 32'h10408000;
      2130: inst = 32'hc404339;
      2131: inst = 32'h8220000;
      2132: inst = 32'h10408000;
      2133: inst = 32'hc40433a;
      2134: inst = 32'h8220000;
      2135: inst = 32'h10408000;
      2136: inst = 32'hc40433b;
      2137: inst = 32'h8220000;
      2138: inst = 32'h10408000;
      2139: inst = 32'hc40433c;
      2140: inst = 32'h8220000;
      2141: inst = 32'h10408000;
      2142: inst = 32'hc40433d;
      2143: inst = 32'h8220000;
      2144: inst = 32'h10408000;
      2145: inst = 32'hc40433e;
      2146: inst = 32'h8220000;
      2147: inst = 32'h10408000;
      2148: inst = 32'hc40433f;
      2149: inst = 32'h8220000;
      2150: inst = 32'h10408000;
      2151: inst = 32'hc404340;
      2152: inst = 32'h8220000;
      2153: inst = 32'h10408000;
      2154: inst = 32'hc404341;
      2155: inst = 32'h8220000;
      2156: inst = 32'h10408000;
      2157: inst = 32'hc404342;
      2158: inst = 32'h8220000;
      2159: inst = 32'h10408000;
      2160: inst = 32'hc404343;
      2161: inst = 32'h8220000;
      2162: inst = 32'h10408000;
      2163: inst = 32'hc404344;
      2164: inst = 32'h8220000;
      2165: inst = 32'h10408000;
      2166: inst = 32'hc404345;
      2167: inst = 32'h8220000;
      2168: inst = 32'h10408000;
      2169: inst = 32'hc404346;
      2170: inst = 32'h8220000;
      2171: inst = 32'h10408000;
      2172: inst = 32'hc404347;
      2173: inst = 32'h8220000;
      2174: inst = 32'h10408000;
      2175: inst = 32'hc404348;
      2176: inst = 32'h8220000;
      2177: inst = 32'h10408000;
      2178: inst = 32'hc40434f;
      2179: inst = 32'h8220000;
      2180: inst = 32'h10408000;
      2181: inst = 32'hc404350;
      2182: inst = 32'h8220000;
      2183: inst = 32'h10408000;
      2184: inst = 32'hc404351;
      2185: inst = 32'h8220000;
      2186: inst = 32'h10408000;
      2187: inst = 32'hc404352;
      2188: inst = 32'h8220000;
      2189: inst = 32'h10408000;
      2190: inst = 32'hc404353;
      2191: inst = 32'h8220000;
      2192: inst = 32'h10408000;
      2193: inst = 32'hc404354;
      2194: inst = 32'h8220000;
      2195: inst = 32'h10408000;
      2196: inst = 32'hc404355;
      2197: inst = 32'h8220000;
      2198: inst = 32'h10408000;
      2199: inst = 32'hc404356;
      2200: inst = 32'h8220000;
      2201: inst = 32'h10408000;
      2202: inst = 32'hc404357;
      2203: inst = 32'h8220000;
      2204: inst = 32'h10408000;
      2205: inst = 32'hc404358;
      2206: inst = 32'h8220000;
      2207: inst = 32'h10408000;
      2208: inst = 32'hc404359;
      2209: inst = 32'h8220000;
      2210: inst = 32'h10408000;
      2211: inst = 32'hc40435a;
      2212: inst = 32'h8220000;
      2213: inst = 32'h10408000;
      2214: inst = 32'hc40435b;
      2215: inst = 32'h8220000;
      2216: inst = 32'h10408000;
      2217: inst = 32'hc404384;
      2218: inst = 32'h8220000;
      2219: inst = 32'h10408000;
      2220: inst = 32'hc404385;
      2221: inst = 32'h8220000;
      2222: inst = 32'h10408000;
      2223: inst = 32'hc404386;
      2224: inst = 32'h8220000;
      2225: inst = 32'h10408000;
      2226: inst = 32'hc404387;
      2227: inst = 32'h8220000;
      2228: inst = 32'h10408000;
      2229: inst = 32'hc404388;
      2230: inst = 32'h8220000;
      2231: inst = 32'h10408000;
      2232: inst = 32'hc404389;
      2233: inst = 32'h8220000;
      2234: inst = 32'h10408000;
      2235: inst = 32'hc40438a;
      2236: inst = 32'h8220000;
      2237: inst = 32'h10408000;
      2238: inst = 32'hc40438b;
      2239: inst = 32'h8220000;
      2240: inst = 32'h10408000;
      2241: inst = 32'hc40438c;
      2242: inst = 32'h8220000;
      2243: inst = 32'h10408000;
      2244: inst = 32'hc40438d;
      2245: inst = 32'h8220000;
      2246: inst = 32'h10408000;
      2247: inst = 32'hc40438e;
      2248: inst = 32'h8220000;
      2249: inst = 32'h10408000;
      2250: inst = 32'hc40438f;
      2251: inst = 32'h8220000;
      2252: inst = 32'h10408000;
      2253: inst = 32'hc404390;
      2254: inst = 32'h8220000;
      2255: inst = 32'h10408000;
      2256: inst = 32'hc404391;
      2257: inst = 32'h8220000;
      2258: inst = 32'h10408000;
      2259: inst = 32'hc404392;
      2260: inst = 32'h8220000;
      2261: inst = 32'h10408000;
      2262: inst = 32'hc404393;
      2263: inst = 32'h8220000;
      2264: inst = 32'h10408000;
      2265: inst = 32'hc404394;
      2266: inst = 32'h8220000;
      2267: inst = 32'h10408000;
      2268: inst = 32'hc404395;
      2269: inst = 32'h8220000;
      2270: inst = 32'h10408000;
      2271: inst = 32'hc404396;
      2272: inst = 32'h8220000;
      2273: inst = 32'h10408000;
      2274: inst = 32'hc404397;
      2275: inst = 32'h8220000;
      2276: inst = 32'h10408000;
      2277: inst = 32'hc404398;
      2278: inst = 32'h8220000;
      2279: inst = 32'h10408000;
      2280: inst = 32'hc404399;
      2281: inst = 32'h8220000;
      2282: inst = 32'h10408000;
      2283: inst = 32'hc40439a;
      2284: inst = 32'h8220000;
      2285: inst = 32'h10408000;
      2286: inst = 32'hc40439b;
      2287: inst = 32'h8220000;
      2288: inst = 32'h10408000;
      2289: inst = 32'hc40439c;
      2290: inst = 32'h8220000;
      2291: inst = 32'h10408000;
      2292: inst = 32'hc40439d;
      2293: inst = 32'h8220000;
      2294: inst = 32'h10408000;
      2295: inst = 32'hc40439e;
      2296: inst = 32'h8220000;
      2297: inst = 32'h10408000;
      2298: inst = 32'hc40439f;
      2299: inst = 32'h8220000;
      2300: inst = 32'h10408000;
      2301: inst = 32'hc4043a0;
      2302: inst = 32'h8220000;
      2303: inst = 32'h10408000;
      2304: inst = 32'hc4043a1;
      2305: inst = 32'h8220000;
      2306: inst = 32'h10408000;
      2307: inst = 32'hc4043a2;
      2308: inst = 32'h8220000;
      2309: inst = 32'h10408000;
      2310: inst = 32'hc4043a3;
      2311: inst = 32'h8220000;
      2312: inst = 32'h10408000;
      2313: inst = 32'hc4043a4;
      2314: inst = 32'h8220000;
      2315: inst = 32'h10408000;
      2316: inst = 32'hc4043a5;
      2317: inst = 32'h8220000;
      2318: inst = 32'h10408000;
      2319: inst = 32'hc4043a6;
      2320: inst = 32'h8220000;
      2321: inst = 32'h10408000;
      2322: inst = 32'hc4043b1;
      2323: inst = 32'h8220000;
      2324: inst = 32'h10408000;
      2325: inst = 32'hc4043b2;
      2326: inst = 32'h8220000;
      2327: inst = 32'h10408000;
      2328: inst = 32'hc4043b3;
      2329: inst = 32'h8220000;
      2330: inst = 32'h10408000;
      2331: inst = 32'hc4043b4;
      2332: inst = 32'h8220000;
      2333: inst = 32'h10408000;
      2334: inst = 32'hc4043b5;
      2335: inst = 32'h8220000;
      2336: inst = 32'h10408000;
      2337: inst = 32'hc4043b6;
      2338: inst = 32'h8220000;
      2339: inst = 32'h10408000;
      2340: inst = 32'hc4043b7;
      2341: inst = 32'h8220000;
      2342: inst = 32'h10408000;
      2343: inst = 32'hc4043b8;
      2344: inst = 32'h8220000;
      2345: inst = 32'h10408000;
      2346: inst = 32'hc4043b9;
      2347: inst = 32'h8220000;
      2348: inst = 32'h10408000;
      2349: inst = 32'hc4043ba;
      2350: inst = 32'h8220000;
      2351: inst = 32'h10408000;
      2352: inst = 32'hc4043bb;
      2353: inst = 32'h8220000;
      2354: inst = 32'h10408000;
      2355: inst = 32'hc4043e4;
      2356: inst = 32'h8220000;
      2357: inst = 32'h10408000;
      2358: inst = 32'hc4043e5;
      2359: inst = 32'h8220000;
      2360: inst = 32'h10408000;
      2361: inst = 32'hc4043e6;
      2362: inst = 32'h8220000;
      2363: inst = 32'h10408000;
      2364: inst = 32'hc4043e7;
      2365: inst = 32'h8220000;
      2366: inst = 32'h10408000;
      2367: inst = 32'hc4043e8;
      2368: inst = 32'h8220000;
      2369: inst = 32'h10408000;
      2370: inst = 32'hc4043e9;
      2371: inst = 32'h8220000;
      2372: inst = 32'h10408000;
      2373: inst = 32'hc4043ea;
      2374: inst = 32'h8220000;
      2375: inst = 32'h10408000;
      2376: inst = 32'hc4043eb;
      2377: inst = 32'h8220000;
      2378: inst = 32'h10408000;
      2379: inst = 32'hc4043ec;
      2380: inst = 32'h8220000;
      2381: inst = 32'h10408000;
      2382: inst = 32'hc4043ed;
      2383: inst = 32'h8220000;
      2384: inst = 32'h10408000;
      2385: inst = 32'hc4043ee;
      2386: inst = 32'h8220000;
      2387: inst = 32'h10408000;
      2388: inst = 32'hc4043ef;
      2389: inst = 32'h8220000;
      2390: inst = 32'h10408000;
      2391: inst = 32'hc4043f0;
      2392: inst = 32'h8220000;
      2393: inst = 32'h10408000;
      2394: inst = 32'hc4043f1;
      2395: inst = 32'h8220000;
      2396: inst = 32'h10408000;
      2397: inst = 32'hc4043f2;
      2398: inst = 32'h8220000;
      2399: inst = 32'h10408000;
      2400: inst = 32'hc4043f3;
      2401: inst = 32'h8220000;
      2402: inst = 32'h10408000;
      2403: inst = 32'hc4043f4;
      2404: inst = 32'h8220000;
      2405: inst = 32'h10408000;
      2406: inst = 32'hc4043f5;
      2407: inst = 32'h8220000;
      2408: inst = 32'h10408000;
      2409: inst = 32'hc4043f6;
      2410: inst = 32'h8220000;
      2411: inst = 32'h10408000;
      2412: inst = 32'hc4043f7;
      2413: inst = 32'h8220000;
      2414: inst = 32'h10408000;
      2415: inst = 32'hc4043f8;
      2416: inst = 32'h8220000;
      2417: inst = 32'h10408000;
      2418: inst = 32'hc4043f9;
      2419: inst = 32'h8220000;
      2420: inst = 32'h10408000;
      2421: inst = 32'hc4043fa;
      2422: inst = 32'h8220000;
      2423: inst = 32'h10408000;
      2424: inst = 32'hc4043fb;
      2425: inst = 32'h8220000;
      2426: inst = 32'h10408000;
      2427: inst = 32'hc4043fc;
      2428: inst = 32'h8220000;
      2429: inst = 32'h10408000;
      2430: inst = 32'hc4043fd;
      2431: inst = 32'h8220000;
      2432: inst = 32'h10408000;
      2433: inst = 32'hc4043fe;
      2434: inst = 32'h8220000;
      2435: inst = 32'h10408000;
      2436: inst = 32'hc4043ff;
      2437: inst = 32'h8220000;
      2438: inst = 32'h10408000;
      2439: inst = 32'hc404400;
      2440: inst = 32'h8220000;
      2441: inst = 32'h10408000;
      2442: inst = 32'hc404401;
      2443: inst = 32'h8220000;
      2444: inst = 32'h10408000;
      2445: inst = 32'hc404402;
      2446: inst = 32'h8220000;
      2447: inst = 32'h10408000;
      2448: inst = 32'hc404403;
      2449: inst = 32'h8220000;
      2450: inst = 32'h10408000;
      2451: inst = 32'hc404404;
      2452: inst = 32'h8220000;
      2453: inst = 32'h10408000;
      2454: inst = 32'hc404405;
      2455: inst = 32'h8220000;
      2456: inst = 32'h10408000;
      2457: inst = 32'hc404412;
      2458: inst = 32'h8220000;
      2459: inst = 32'h10408000;
      2460: inst = 32'hc404413;
      2461: inst = 32'h8220000;
      2462: inst = 32'h10408000;
      2463: inst = 32'hc404414;
      2464: inst = 32'h8220000;
      2465: inst = 32'h10408000;
      2466: inst = 32'hc404415;
      2467: inst = 32'h8220000;
      2468: inst = 32'h10408000;
      2469: inst = 32'hc404416;
      2470: inst = 32'h8220000;
      2471: inst = 32'h10408000;
      2472: inst = 32'hc404417;
      2473: inst = 32'h8220000;
      2474: inst = 32'h10408000;
      2475: inst = 32'hc404418;
      2476: inst = 32'h8220000;
      2477: inst = 32'h10408000;
      2478: inst = 32'hc404419;
      2479: inst = 32'h8220000;
      2480: inst = 32'h10408000;
      2481: inst = 32'hc40441a;
      2482: inst = 32'h8220000;
      2483: inst = 32'h10408000;
      2484: inst = 32'hc40441b;
      2485: inst = 32'h8220000;
      2486: inst = 32'h10408000;
      2487: inst = 32'hc404444;
      2488: inst = 32'h8220000;
      2489: inst = 32'h10408000;
      2490: inst = 32'hc404445;
      2491: inst = 32'h8220000;
      2492: inst = 32'h10408000;
      2493: inst = 32'hc404446;
      2494: inst = 32'h8220000;
      2495: inst = 32'h10408000;
      2496: inst = 32'hc404447;
      2497: inst = 32'h8220000;
      2498: inst = 32'h10408000;
      2499: inst = 32'hc404448;
      2500: inst = 32'h8220000;
      2501: inst = 32'h10408000;
      2502: inst = 32'hc404449;
      2503: inst = 32'h8220000;
      2504: inst = 32'h10408000;
      2505: inst = 32'hc40444a;
      2506: inst = 32'h8220000;
      2507: inst = 32'h10408000;
      2508: inst = 32'hc40444b;
      2509: inst = 32'h8220000;
      2510: inst = 32'h10408000;
      2511: inst = 32'hc40444c;
      2512: inst = 32'h8220000;
      2513: inst = 32'h10408000;
      2514: inst = 32'hc40444d;
      2515: inst = 32'h8220000;
      2516: inst = 32'h10408000;
      2517: inst = 32'hc40444e;
      2518: inst = 32'h8220000;
      2519: inst = 32'h10408000;
      2520: inst = 32'hc40444f;
      2521: inst = 32'h8220000;
      2522: inst = 32'h10408000;
      2523: inst = 32'hc404450;
      2524: inst = 32'h8220000;
      2525: inst = 32'h10408000;
      2526: inst = 32'hc404451;
      2527: inst = 32'h8220000;
      2528: inst = 32'h10408000;
      2529: inst = 32'hc404452;
      2530: inst = 32'h8220000;
      2531: inst = 32'h10408000;
      2532: inst = 32'hc404453;
      2533: inst = 32'h8220000;
      2534: inst = 32'h10408000;
      2535: inst = 32'hc404454;
      2536: inst = 32'h8220000;
      2537: inst = 32'h10408000;
      2538: inst = 32'hc404455;
      2539: inst = 32'h8220000;
      2540: inst = 32'h10408000;
      2541: inst = 32'hc404456;
      2542: inst = 32'h8220000;
      2543: inst = 32'h10408000;
      2544: inst = 32'hc404457;
      2545: inst = 32'h8220000;
      2546: inst = 32'h10408000;
      2547: inst = 32'hc404458;
      2548: inst = 32'h8220000;
      2549: inst = 32'h10408000;
      2550: inst = 32'hc404459;
      2551: inst = 32'h8220000;
      2552: inst = 32'h10408000;
      2553: inst = 32'hc40445a;
      2554: inst = 32'h8220000;
      2555: inst = 32'h10408000;
      2556: inst = 32'hc40445b;
      2557: inst = 32'h8220000;
      2558: inst = 32'h10408000;
      2559: inst = 32'hc40445c;
      2560: inst = 32'h8220000;
      2561: inst = 32'h10408000;
      2562: inst = 32'hc40445d;
      2563: inst = 32'h8220000;
      2564: inst = 32'h10408000;
      2565: inst = 32'hc40445e;
      2566: inst = 32'h8220000;
      2567: inst = 32'h10408000;
      2568: inst = 32'hc40445f;
      2569: inst = 32'h8220000;
      2570: inst = 32'h10408000;
      2571: inst = 32'hc404460;
      2572: inst = 32'h8220000;
      2573: inst = 32'h10408000;
      2574: inst = 32'hc404461;
      2575: inst = 32'h8220000;
      2576: inst = 32'h10408000;
      2577: inst = 32'hc404462;
      2578: inst = 32'h8220000;
      2579: inst = 32'h10408000;
      2580: inst = 32'hc404463;
      2581: inst = 32'h8220000;
      2582: inst = 32'h10408000;
      2583: inst = 32'hc404464;
      2584: inst = 32'h8220000;
      2585: inst = 32'h10408000;
      2586: inst = 32'hc404465;
      2587: inst = 32'h8220000;
      2588: inst = 32'h10408000;
      2589: inst = 32'hc404466;
      2590: inst = 32'h8220000;
      2591: inst = 32'h10408000;
      2592: inst = 32'hc404467;
      2593: inst = 32'h8220000;
      2594: inst = 32'h10408000;
      2595: inst = 32'hc404468;
      2596: inst = 32'h8220000;
      2597: inst = 32'h10408000;
      2598: inst = 32'hc404469;
      2599: inst = 32'h8220000;
      2600: inst = 32'h10408000;
      2601: inst = 32'hc40446e;
      2602: inst = 32'h8220000;
      2603: inst = 32'h10408000;
      2604: inst = 32'hc40446f;
      2605: inst = 32'h8220000;
      2606: inst = 32'h10408000;
      2607: inst = 32'hc404470;
      2608: inst = 32'h8220000;
      2609: inst = 32'h10408000;
      2610: inst = 32'hc404471;
      2611: inst = 32'h8220000;
      2612: inst = 32'h10408000;
      2613: inst = 32'hc404472;
      2614: inst = 32'h8220000;
      2615: inst = 32'h10408000;
      2616: inst = 32'hc404473;
      2617: inst = 32'h8220000;
      2618: inst = 32'h10408000;
      2619: inst = 32'hc404474;
      2620: inst = 32'h8220000;
      2621: inst = 32'h10408000;
      2622: inst = 32'hc404475;
      2623: inst = 32'h8220000;
      2624: inst = 32'h10408000;
      2625: inst = 32'hc404476;
      2626: inst = 32'h8220000;
      2627: inst = 32'h10408000;
      2628: inst = 32'hc404477;
      2629: inst = 32'h8220000;
      2630: inst = 32'h10408000;
      2631: inst = 32'hc404478;
      2632: inst = 32'h8220000;
      2633: inst = 32'h10408000;
      2634: inst = 32'hc404479;
      2635: inst = 32'h8220000;
      2636: inst = 32'h10408000;
      2637: inst = 32'hc40447a;
      2638: inst = 32'h8220000;
      2639: inst = 32'h10408000;
      2640: inst = 32'hc40447b;
      2641: inst = 32'h8220000;
      2642: inst = 32'h10408000;
      2643: inst = 32'hc4044a4;
      2644: inst = 32'h8220000;
      2645: inst = 32'h10408000;
      2646: inst = 32'hc4044a5;
      2647: inst = 32'h8220000;
      2648: inst = 32'h10408000;
      2649: inst = 32'hc4044a6;
      2650: inst = 32'h8220000;
      2651: inst = 32'h10408000;
      2652: inst = 32'hc4044a7;
      2653: inst = 32'h8220000;
      2654: inst = 32'h10408000;
      2655: inst = 32'hc4044a8;
      2656: inst = 32'h8220000;
      2657: inst = 32'h10408000;
      2658: inst = 32'hc4044a9;
      2659: inst = 32'h8220000;
      2660: inst = 32'h10408000;
      2661: inst = 32'hc4044aa;
      2662: inst = 32'h8220000;
      2663: inst = 32'h10408000;
      2664: inst = 32'hc4044ab;
      2665: inst = 32'h8220000;
      2666: inst = 32'h10408000;
      2667: inst = 32'hc4044ac;
      2668: inst = 32'h8220000;
      2669: inst = 32'h10408000;
      2670: inst = 32'hc4044ad;
      2671: inst = 32'h8220000;
      2672: inst = 32'h10408000;
      2673: inst = 32'hc4044ae;
      2674: inst = 32'h8220000;
      2675: inst = 32'h10408000;
      2676: inst = 32'hc4044af;
      2677: inst = 32'h8220000;
      2678: inst = 32'h10408000;
      2679: inst = 32'hc4044b0;
      2680: inst = 32'h8220000;
      2681: inst = 32'h10408000;
      2682: inst = 32'hc4044b1;
      2683: inst = 32'h8220000;
      2684: inst = 32'h10408000;
      2685: inst = 32'hc4044b6;
      2686: inst = 32'h8220000;
      2687: inst = 32'h10408000;
      2688: inst = 32'hc4044b7;
      2689: inst = 32'h8220000;
      2690: inst = 32'h10408000;
      2691: inst = 32'hc4044b8;
      2692: inst = 32'h8220000;
      2693: inst = 32'h10408000;
      2694: inst = 32'hc4044b9;
      2695: inst = 32'h8220000;
      2696: inst = 32'h10408000;
      2697: inst = 32'hc4044ba;
      2698: inst = 32'h8220000;
      2699: inst = 32'h10408000;
      2700: inst = 32'hc4044bb;
      2701: inst = 32'h8220000;
      2702: inst = 32'h10408000;
      2703: inst = 32'hc4044bc;
      2704: inst = 32'h8220000;
      2705: inst = 32'h10408000;
      2706: inst = 32'hc4044bd;
      2707: inst = 32'h8220000;
      2708: inst = 32'h10408000;
      2709: inst = 32'hc4044be;
      2710: inst = 32'h8220000;
      2711: inst = 32'h10408000;
      2712: inst = 32'hc4044bf;
      2713: inst = 32'h8220000;
      2714: inst = 32'h10408000;
      2715: inst = 32'hc4044c0;
      2716: inst = 32'h8220000;
      2717: inst = 32'h10408000;
      2718: inst = 32'hc4044c1;
      2719: inst = 32'h8220000;
      2720: inst = 32'h10408000;
      2721: inst = 32'hc4044c2;
      2722: inst = 32'h8220000;
      2723: inst = 32'h10408000;
      2724: inst = 32'hc4044c3;
      2725: inst = 32'h8220000;
      2726: inst = 32'h10408000;
      2727: inst = 32'hc4044c4;
      2728: inst = 32'h8220000;
      2729: inst = 32'h10408000;
      2730: inst = 32'hc4044c5;
      2731: inst = 32'h8220000;
      2732: inst = 32'h10408000;
      2733: inst = 32'hc4044c6;
      2734: inst = 32'h8220000;
      2735: inst = 32'h10408000;
      2736: inst = 32'hc4044c7;
      2737: inst = 32'h8220000;
      2738: inst = 32'h10408000;
      2739: inst = 32'hc4044c8;
      2740: inst = 32'h8220000;
      2741: inst = 32'h10408000;
      2742: inst = 32'hc4044c9;
      2743: inst = 32'h8220000;
      2744: inst = 32'h10408000;
      2745: inst = 32'hc4044ca;
      2746: inst = 32'h8220000;
      2747: inst = 32'h10408000;
      2748: inst = 32'hc4044cd;
      2749: inst = 32'h8220000;
      2750: inst = 32'h10408000;
      2751: inst = 32'hc4044ce;
      2752: inst = 32'h8220000;
      2753: inst = 32'h10408000;
      2754: inst = 32'hc4044cf;
      2755: inst = 32'h8220000;
      2756: inst = 32'h10408000;
      2757: inst = 32'hc4044d0;
      2758: inst = 32'h8220000;
      2759: inst = 32'h10408000;
      2760: inst = 32'hc4044d1;
      2761: inst = 32'h8220000;
      2762: inst = 32'h10408000;
      2763: inst = 32'hc4044d2;
      2764: inst = 32'h8220000;
      2765: inst = 32'h10408000;
      2766: inst = 32'hc4044d3;
      2767: inst = 32'h8220000;
      2768: inst = 32'h10408000;
      2769: inst = 32'hc4044d4;
      2770: inst = 32'h8220000;
      2771: inst = 32'h10408000;
      2772: inst = 32'hc4044d5;
      2773: inst = 32'h8220000;
      2774: inst = 32'h10408000;
      2775: inst = 32'hc4044d6;
      2776: inst = 32'h8220000;
      2777: inst = 32'h10408000;
      2778: inst = 32'hc4044d7;
      2779: inst = 32'h8220000;
      2780: inst = 32'h10408000;
      2781: inst = 32'hc4044d8;
      2782: inst = 32'h8220000;
      2783: inst = 32'h10408000;
      2784: inst = 32'hc4044d9;
      2785: inst = 32'h8220000;
      2786: inst = 32'h10408000;
      2787: inst = 32'hc4044da;
      2788: inst = 32'h8220000;
      2789: inst = 32'h10408000;
      2790: inst = 32'hc4044db;
      2791: inst = 32'h8220000;
      2792: inst = 32'h10408000;
      2793: inst = 32'hc404504;
      2794: inst = 32'h8220000;
      2795: inst = 32'h10408000;
      2796: inst = 32'hc404505;
      2797: inst = 32'h8220000;
      2798: inst = 32'h10408000;
      2799: inst = 32'hc404506;
      2800: inst = 32'h8220000;
      2801: inst = 32'h10408000;
      2802: inst = 32'hc404507;
      2803: inst = 32'h8220000;
      2804: inst = 32'h10408000;
      2805: inst = 32'hc404508;
      2806: inst = 32'h8220000;
      2807: inst = 32'h10408000;
      2808: inst = 32'hc404509;
      2809: inst = 32'h8220000;
      2810: inst = 32'h10408000;
      2811: inst = 32'hc40450a;
      2812: inst = 32'h8220000;
      2813: inst = 32'h10408000;
      2814: inst = 32'hc40450b;
      2815: inst = 32'h8220000;
      2816: inst = 32'h10408000;
      2817: inst = 32'hc40450c;
      2818: inst = 32'h8220000;
      2819: inst = 32'h10408000;
      2820: inst = 32'hc40450d;
      2821: inst = 32'h8220000;
      2822: inst = 32'h10408000;
      2823: inst = 32'hc40450e;
      2824: inst = 32'h8220000;
      2825: inst = 32'h10408000;
      2826: inst = 32'hc40450f;
      2827: inst = 32'h8220000;
      2828: inst = 32'h10408000;
      2829: inst = 32'hc404510;
      2830: inst = 32'h8220000;
      2831: inst = 32'h10408000;
      2832: inst = 32'hc404511;
      2833: inst = 32'h8220000;
      2834: inst = 32'h10408000;
      2835: inst = 32'hc404512;
      2836: inst = 32'h8220000;
      2837: inst = 32'h10408000;
      2838: inst = 32'hc404515;
      2839: inst = 32'h8220000;
      2840: inst = 32'h10408000;
      2841: inst = 32'hc404516;
      2842: inst = 32'h8220000;
      2843: inst = 32'h10408000;
      2844: inst = 32'hc404517;
      2845: inst = 32'h8220000;
      2846: inst = 32'h10408000;
      2847: inst = 32'hc404518;
      2848: inst = 32'h8220000;
      2849: inst = 32'h10408000;
      2850: inst = 32'hc404519;
      2851: inst = 32'h8220000;
      2852: inst = 32'h10408000;
      2853: inst = 32'hc40451a;
      2854: inst = 32'h8220000;
      2855: inst = 32'h10408000;
      2856: inst = 32'hc40451b;
      2857: inst = 32'h8220000;
      2858: inst = 32'h10408000;
      2859: inst = 32'hc40451c;
      2860: inst = 32'h8220000;
      2861: inst = 32'h10408000;
      2862: inst = 32'hc40451d;
      2863: inst = 32'h8220000;
      2864: inst = 32'h10408000;
      2865: inst = 32'hc40451e;
      2866: inst = 32'h8220000;
      2867: inst = 32'h10408000;
      2868: inst = 32'hc40451f;
      2869: inst = 32'h8220000;
      2870: inst = 32'h10408000;
      2871: inst = 32'hc404520;
      2872: inst = 32'h8220000;
      2873: inst = 32'h10408000;
      2874: inst = 32'hc404521;
      2875: inst = 32'h8220000;
      2876: inst = 32'h10408000;
      2877: inst = 32'hc404522;
      2878: inst = 32'h8220000;
      2879: inst = 32'h10408000;
      2880: inst = 32'hc404523;
      2881: inst = 32'h8220000;
      2882: inst = 32'h10408000;
      2883: inst = 32'hc404524;
      2884: inst = 32'h8220000;
      2885: inst = 32'h10408000;
      2886: inst = 32'hc404525;
      2887: inst = 32'h8220000;
      2888: inst = 32'h10408000;
      2889: inst = 32'hc404526;
      2890: inst = 32'h8220000;
      2891: inst = 32'h10408000;
      2892: inst = 32'hc404527;
      2893: inst = 32'h8220000;
      2894: inst = 32'h10408000;
      2895: inst = 32'hc404528;
      2896: inst = 32'h8220000;
      2897: inst = 32'h10408000;
      2898: inst = 32'hc404529;
      2899: inst = 32'h8220000;
      2900: inst = 32'h10408000;
      2901: inst = 32'hc40452a;
      2902: inst = 32'h8220000;
      2903: inst = 32'h10408000;
      2904: inst = 32'hc40452b;
      2905: inst = 32'h8220000;
      2906: inst = 32'h10408000;
      2907: inst = 32'hc40452c;
      2908: inst = 32'h8220000;
      2909: inst = 32'h10408000;
      2910: inst = 32'hc40452d;
      2911: inst = 32'h8220000;
      2912: inst = 32'h10408000;
      2913: inst = 32'hc40452e;
      2914: inst = 32'h8220000;
      2915: inst = 32'h10408000;
      2916: inst = 32'hc40452f;
      2917: inst = 32'h8220000;
      2918: inst = 32'h10408000;
      2919: inst = 32'hc404530;
      2920: inst = 32'h8220000;
      2921: inst = 32'h10408000;
      2922: inst = 32'hc404531;
      2923: inst = 32'h8220000;
      2924: inst = 32'h10408000;
      2925: inst = 32'hc404532;
      2926: inst = 32'h8220000;
      2927: inst = 32'h10408000;
      2928: inst = 32'hc404533;
      2929: inst = 32'h8220000;
      2930: inst = 32'h10408000;
      2931: inst = 32'hc404534;
      2932: inst = 32'h8220000;
      2933: inst = 32'h10408000;
      2934: inst = 32'hc404535;
      2935: inst = 32'h8220000;
      2936: inst = 32'h10408000;
      2937: inst = 32'hc404536;
      2938: inst = 32'h8220000;
      2939: inst = 32'h10408000;
      2940: inst = 32'hc404537;
      2941: inst = 32'h8220000;
      2942: inst = 32'h10408000;
      2943: inst = 32'hc404538;
      2944: inst = 32'h8220000;
      2945: inst = 32'h10408000;
      2946: inst = 32'hc404539;
      2947: inst = 32'h8220000;
      2948: inst = 32'h10408000;
      2949: inst = 32'hc40453a;
      2950: inst = 32'h8220000;
      2951: inst = 32'h10408000;
      2952: inst = 32'hc40453b;
      2953: inst = 32'h8220000;
      2954: inst = 32'h10408000;
      2955: inst = 32'hc404564;
      2956: inst = 32'h8220000;
      2957: inst = 32'h10408000;
      2958: inst = 32'hc404565;
      2959: inst = 32'h8220000;
      2960: inst = 32'h10408000;
      2961: inst = 32'hc404566;
      2962: inst = 32'h8220000;
      2963: inst = 32'h10408000;
      2964: inst = 32'hc404567;
      2965: inst = 32'h8220000;
      2966: inst = 32'h10408000;
      2967: inst = 32'hc404568;
      2968: inst = 32'h8220000;
      2969: inst = 32'h10408000;
      2970: inst = 32'hc404569;
      2971: inst = 32'h8220000;
      2972: inst = 32'h10408000;
      2973: inst = 32'hc40456a;
      2974: inst = 32'h8220000;
      2975: inst = 32'h10408000;
      2976: inst = 32'hc40456b;
      2977: inst = 32'h8220000;
      2978: inst = 32'h10408000;
      2979: inst = 32'hc40456c;
      2980: inst = 32'h8220000;
      2981: inst = 32'h10408000;
      2982: inst = 32'hc40456d;
      2983: inst = 32'h8220000;
      2984: inst = 32'h10408000;
      2985: inst = 32'hc40456e;
      2986: inst = 32'h8220000;
      2987: inst = 32'h10408000;
      2988: inst = 32'hc40456f;
      2989: inst = 32'h8220000;
      2990: inst = 32'h10408000;
      2991: inst = 32'hc404570;
      2992: inst = 32'h8220000;
      2993: inst = 32'h10408000;
      2994: inst = 32'hc404571;
      2995: inst = 32'h8220000;
      2996: inst = 32'h10408000;
      2997: inst = 32'hc404572;
      2998: inst = 32'h8220000;
      2999: inst = 32'h10408000;
      3000: inst = 32'hc404573;
      3001: inst = 32'h8220000;
      3002: inst = 32'h10408000;
      3003: inst = 32'hc404574;
      3004: inst = 32'h8220000;
      3005: inst = 32'h10408000;
      3006: inst = 32'hc404575;
      3007: inst = 32'h8220000;
      3008: inst = 32'h10408000;
      3009: inst = 32'hc404576;
      3010: inst = 32'h8220000;
      3011: inst = 32'h10408000;
      3012: inst = 32'hc404577;
      3013: inst = 32'h8220000;
      3014: inst = 32'h10408000;
      3015: inst = 32'hc404578;
      3016: inst = 32'h8220000;
      3017: inst = 32'h10408000;
      3018: inst = 32'hc404579;
      3019: inst = 32'h8220000;
      3020: inst = 32'h10408000;
      3021: inst = 32'hc40457a;
      3022: inst = 32'h8220000;
      3023: inst = 32'h10408000;
      3024: inst = 32'hc40457b;
      3025: inst = 32'h8220000;
      3026: inst = 32'h10408000;
      3027: inst = 32'hc40457c;
      3028: inst = 32'h8220000;
      3029: inst = 32'h10408000;
      3030: inst = 32'hc40457d;
      3031: inst = 32'h8220000;
      3032: inst = 32'h10408000;
      3033: inst = 32'hc40457e;
      3034: inst = 32'h8220000;
      3035: inst = 32'h10408000;
      3036: inst = 32'hc40457f;
      3037: inst = 32'h8220000;
      3038: inst = 32'h10408000;
      3039: inst = 32'hc404580;
      3040: inst = 32'h8220000;
      3041: inst = 32'h10408000;
      3042: inst = 32'hc404581;
      3043: inst = 32'h8220000;
      3044: inst = 32'h10408000;
      3045: inst = 32'hc404582;
      3046: inst = 32'h8220000;
      3047: inst = 32'h10408000;
      3048: inst = 32'hc404583;
      3049: inst = 32'h8220000;
      3050: inst = 32'h10408000;
      3051: inst = 32'hc404584;
      3052: inst = 32'h8220000;
      3053: inst = 32'h10408000;
      3054: inst = 32'hc404585;
      3055: inst = 32'h8220000;
      3056: inst = 32'h10408000;
      3057: inst = 32'hc404586;
      3058: inst = 32'h8220000;
      3059: inst = 32'h10408000;
      3060: inst = 32'hc404587;
      3061: inst = 32'h8220000;
      3062: inst = 32'h10408000;
      3063: inst = 32'hc404588;
      3064: inst = 32'h8220000;
      3065: inst = 32'h10408000;
      3066: inst = 32'hc404589;
      3067: inst = 32'h8220000;
      3068: inst = 32'h10408000;
      3069: inst = 32'hc40458a;
      3070: inst = 32'h8220000;
      3071: inst = 32'h10408000;
      3072: inst = 32'hc40458b;
      3073: inst = 32'h8220000;
      3074: inst = 32'h10408000;
      3075: inst = 32'hc40458c;
      3076: inst = 32'h8220000;
      3077: inst = 32'h10408000;
      3078: inst = 32'hc40458d;
      3079: inst = 32'h8220000;
      3080: inst = 32'h10408000;
      3081: inst = 32'hc40458e;
      3082: inst = 32'h8220000;
      3083: inst = 32'h10408000;
      3084: inst = 32'hc40458f;
      3085: inst = 32'h8220000;
      3086: inst = 32'h10408000;
      3087: inst = 32'hc404590;
      3088: inst = 32'h8220000;
      3089: inst = 32'h10408000;
      3090: inst = 32'hc404591;
      3091: inst = 32'h8220000;
      3092: inst = 32'h10408000;
      3093: inst = 32'hc404592;
      3094: inst = 32'h8220000;
      3095: inst = 32'h10408000;
      3096: inst = 32'hc404593;
      3097: inst = 32'h8220000;
      3098: inst = 32'h10408000;
      3099: inst = 32'hc404594;
      3100: inst = 32'h8220000;
      3101: inst = 32'h10408000;
      3102: inst = 32'hc404595;
      3103: inst = 32'h8220000;
      3104: inst = 32'h10408000;
      3105: inst = 32'hc404596;
      3106: inst = 32'h8220000;
      3107: inst = 32'h10408000;
      3108: inst = 32'hc404597;
      3109: inst = 32'h8220000;
      3110: inst = 32'h10408000;
      3111: inst = 32'hc404598;
      3112: inst = 32'h8220000;
      3113: inst = 32'h10408000;
      3114: inst = 32'hc404599;
      3115: inst = 32'h8220000;
      3116: inst = 32'h10408000;
      3117: inst = 32'hc40459a;
      3118: inst = 32'h8220000;
      3119: inst = 32'h10408000;
      3120: inst = 32'hc40459b;
      3121: inst = 32'h8220000;
      3122: inst = 32'h10408000;
      3123: inst = 32'hc4045c4;
      3124: inst = 32'h8220000;
      3125: inst = 32'h10408000;
      3126: inst = 32'hc4045c5;
      3127: inst = 32'h8220000;
      3128: inst = 32'h10408000;
      3129: inst = 32'hc4045c6;
      3130: inst = 32'h8220000;
      3131: inst = 32'h10408000;
      3132: inst = 32'hc4045c7;
      3133: inst = 32'h8220000;
      3134: inst = 32'h10408000;
      3135: inst = 32'hc4045c8;
      3136: inst = 32'h8220000;
      3137: inst = 32'h10408000;
      3138: inst = 32'hc4045c9;
      3139: inst = 32'h8220000;
      3140: inst = 32'h10408000;
      3141: inst = 32'hc4045ca;
      3142: inst = 32'h8220000;
      3143: inst = 32'h10408000;
      3144: inst = 32'hc4045cb;
      3145: inst = 32'h8220000;
      3146: inst = 32'h10408000;
      3147: inst = 32'hc4045cc;
      3148: inst = 32'h8220000;
      3149: inst = 32'h10408000;
      3150: inst = 32'hc4045cd;
      3151: inst = 32'h8220000;
      3152: inst = 32'h10408000;
      3153: inst = 32'hc4045ce;
      3154: inst = 32'h8220000;
      3155: inst = 32'h10408000;
      3156: inst = 32'hc4045cf;
      3157: inst = 32'h8220000;
      3158: inst = 32'h10408000;
      3159: inst = 32'hc4045d0;
      3160: inst = 32'h8220000;
      3161: inst = 32'h10408000;
      3162: inst = 32'hc4045d1;
      3163: inst = 32'h8220000;
      3164: inst = 32'h10408000;
      3165: inst = 32'hc4045d2;
      3166: inst = 32'h8220000;
      3167: inst = 32'h10408000;
      3168: inst = 32'hc4045d3;
      3169: inst = 32'h8220000;
      3170: inst = 32'h10408000;
      3171: inst = 32'hc4045d4;
      3172: inst = 32'h8220000;
      3173: inst = 32'h10408000;
      3174: inst = 32'hc4045d5;
      3175: inst = 32'h8220000;
      3176: inst = 32'h10408000;
      3177: inst = 32'hc4045d6;
      3178: inst = 32'h8220000;
      3179: inst = 32'h10408000;
      3180: inst = 32'hc4045d7;
      3181: inst = 32'h8220000;
      3182: inst = 32'h10408000;
      3183: inst = 32'hc4045d8;
      3184: inst = 32'h8220000;
      3185: inst = 32'h10408000;
      3186: inst = 32'hc4045d9;
      3187: inst = 32'h8220000;
      3188: inst = 32'h10408000;
      3189: inst = 32'hc4045da;
      3190: inst = 32'h8220000;
      3191: inst = 32'h10408000;
      3192: inst = 32'hc4045db;
      3193: inst = 32'h8220000;
      3194: inst = 32'h10408000;
      3195: inst = 32'hc4045dc;
      3196: inst = 32'h8220000;
      3197: inst = 32'h10408000;
      3198: inst = 32'hc4045dd;
      3199: inst = 32'h8220000;
      3200: inst = 32'h10408000;
      3201: inst = 32'hc4045de;
      3202: inst = 32'h8220000;
      3203: inst = 32'h10408000;
      3204: inst = 32'hc4045df;
      3205: inst = 32'h8220000;
      3206: inst = 32'h10408000;
      3207: inst = 32'hc4045e0;
      3208: inst = 32'h8220000;
      3209: inst = 32'h10408000;
      3210: inst = 32'hc4045e1;
      3211: inst = 32'h8220000;
      3212: inst = 32'h10408000;
      3213: inst = 32'hc4045e2;
      3214: inst = 32'h8220000;
      3215: inst = 32'h10408000;
      3216: inst = 32'hc4045e3;
      3217: inst = 32'h8220000;
      3218: inst = 32'h10408000;
      3219: inst = 32'hc4045e4;
      3220: inst = 32'h8220000;
      3221: inst = 32'h10408000;
      3222: inst = 32'hc4045e5;
      3223: inst = 32'h8220000;
      3224: inst = 32'h10408000;
      3225: inst = 32'hc4045e6;
      3226: inst = 32'h8220000;
      3227: inst = 32'h10408000;
      3228: inst = 32'hc4045e7;
      3229: inst = 32'h8220000;
      3230: inst = 32'h10408000;
      3231: inst = 32'hc4045e8;
      3232: inst = 32'h8220000;
      3233: inst = 32'h10408000;
      3234: inst = 32'hc4045e9;
      3235: inst = 32'h8220000;
      3236: inst = 32'h10408000;
      3237: inst = 32'hc4045ea;
      3238: inst = 32'h8220000;
      3239: inst = 32'h10408000;
      3240: inst = 32'hc4045eb;
      3241: inst = 32'h8220000;
      3242: inst = 32'h10408000;
      3243: inst = 32'hc4045ec;
      3244: inst = 32'h8220000;
      3245: inst = 32'h10408000;
      3246: inst = 32'hc4045ed;
      3247: inst = 32'h8220000;
      3248: inst = 32'h10408000;
      3249: inst = 32'hc4045ee;
      3250: inst = 32'h8220000;
      3251: inst = 32'h10408000;
      3252: inst = 32'hc4045ef;
      3253: inst = 32'h8220000;
      3254: inst = 32'h10408000;
      3255: inst = 32'hc4045f0;
      3256: inst = 32'h8220000;
      3257: inst = 32'h10408000;
      3258: inst = 32'hc4045f1;
      3259: inst = 32'h8220000;
      3260: inst = 32'h10408000;
      3261: inst = 32'hc4045f2;
      3262: inst = 32'h8220000;
      3263: inst = 32'h10408000;
      3264: inst = 32'hc4045f3;
      3265: inst = 32'h8220000;
      3266: inst = 32'h10408000;
      3267: inst = 32'hc4045f4;
      3268: inst = 32'h8220000;
      3269: inst = 32'h10408000;
      3270: inst = 32'hc4045f5;
      3271: inst = 32'h8220000;
      3272: inst = 32'h10408000;
      3273: inst = 32'hc4045f6;
      3274: inst = 32'h8220000;
      3275: inst = 32'h10408000;
      3276: inst = 32'hc4045f7;
      3277: inst = 32'h8220000;
      3278: inst = 32'h10408000;
      3279: inst = 32'hc4045f8;
      3280: inst = 32'h8220000;
      3281: inst = 32'h10408000;
      3282: inst = 32'hc4045f9;
      3283: inst = 32'h8220000;
      3284: inst = 32'h10408000;
      3285: inst = 32'hc4045fa;
      3286: inst = 32'h8220000;
      3287: inst = 32'h10408000;
      3288: inst = 32'hc4045fb;
      3289: inst = 32'h8220000;
      3290: inst = 32'h10408000;
      3291: inst = 32'hc404624;
      3292: inst = 32'h8220000;
      3293: inst = 32'h10408000;
      3294: inst = 32'hc404625;
      3295: inst = 32'h8220000;
      3296: inst = 32'h10408000;
      3297: inst = 32'hc404626;
      3298: inst = 32'h8220000;
      3299: inst = 32'h10408000;
      3300: inst = 32'hc404627;
      3301: inst = 32'h8220000;
      3302: inst = 32'h10408000;
      3303: inst = 32'hc404628;
      3304: inst = 32'h8220000;
      3305: inst = 32'h10408000;
      3306: inst = 32'hc404629;
      3307: inst = 32'h8220000;
      3308: inst = 32'h10408000;
      3309: inst = 32'hc40462a;
      3310: inst = 32'h8220000;
      3311: inst = 32'h10408000;
      3312: inst = 32'hc40462b;
      3313: inst = 32'h8220000;
      3314: inst = 32'h10408000;
      3315: inst = 32'hc40462c;
      3316: inst = 32'h8220000;
      3317: inst = 32'h10408000;
      3318: inst = 32'hc40462d;
      3319: inst = 32'h8220000;
      3320: inst = 32'h10408000;
      3321: inst = 32'hc40462e;
      3322: inst = 32'h8220000;
      3323: inst = 32'h10408000;
      3324: inst = 32'hc40462f;
      3325: inst = 32'h8220000;
      3326: inst = 32'h10408000;
      3327: inst = 32'hc404630;
      3328: inst = 32'h8220000;
      3329: inst = 32'h10408000;
      3330: inst = 32'hc404631;
      3331: inst = 32'h8220000;
      3332: inst = 32'h10408000;
      3333: inst = 32'hc404632;
      3334: inst = 32'h8220000;
      3335: inst = 32'h10408000;
      3336: inst = 32'hc404633;
      3337: inst = 32'h8220000;
      3338: inst = 32'h10408000;
      3339: inst = 32'hc404634;
      3340: inst = 32'h8220000;
      3341: inst = 32'h10408000;
      3342: inst = 32'hc404635;
      3343: inst = 32'h8220000;
      3344: inst = 32'h10408000;
      3345: inst = 32'hc404636;
      3346: inst = 32'h8220000;
      3347: inst = 32'h10408000;
      3348: inst = 32'hc404637;
      3349: inst = 32'h8220000;
      3350: inst = 32'h10408000;
      3351: inst = 32'hc404638;
      3352: inst = 32'h8220000;
      3353: inst = 32'h10408000;
      3354: inst = 32'hc404639;
      3355: inst = 32'h8220000;
      3356: inst = 32'h10408000;
      3357: inst = 32'hc40463a;
      3358: inst = 32'h8220000;
      3359: inst = 32'h10408000;
      3360: inst = 32'hc40463b;
      3361: inst = 32'h8220000;
      3362: inst = 32'h10408000;
      3363: inst = 32'hc40463c;
      3364: inst = 32'h8220000;
      3365: inst = 32'h10408000;
      3366: inst = 32'hc40463d;
      3367: inst = 32'h8220000;
      3368: inst = 32'h10408000;
      3369: inst = 32'hc40463e;
      3370: inst = 32'h8220000;
      3371: inst = 32'h10408000;
      3372: inst = 32'hc40463f;
      3373: inst = 32'h8220000;
      3374: inst = 32'h10408000;
      3375: inst = 32'hc404640;
      3376: inst = 32'h8220000;
      3377: inst = 32'h10408000;
      3378: inst = 32'hc404641;
      3379: inst = 32'h8220000;
      3380: inst = 32'h10408000;
      3381: inst = 32'hc404642;
      3382: inst = 32'h8220000;
      3383: inst = 32'h10408000;
      3384: inst = 32'hc404643;
      3385: inst = 32'h8220000;
      3386: inst = 32'h10408000;
      3387: inst = 32'hc404644;
      3388: inst = 32'h8220000;
      3389: inst = 32'h10408000;
      3390: inst = 32'hc404645;
      3391: inst = 32'h8220000;
      3392: inst = 32'h10408000;
      3393: inst = 32'hc404646;
      3394: inst = 32'h8220000;
      3395: inst = 32'h10408000;
      3396: inst = 32'hc404647;
      3397: inst = 32'h8220000;
      3398: inst = 32'h10408000;
      3399: inst = 32'hc404648;
      3400: inst = 32'h8220000;
      3401: inst = 32'h10408000;
      3402: inst = 32'hc404649;
      3403: inst = 32'h8220000;
      3404: inst = 32'h10408000;
      3405: inst = 32'hc40464a;
      3406: inst = 32'h8220000;
      3407: inst = 32'h10408000;
      3408: inst = 32'hc40464b;
      3409: inst = 32'h8220000;
      3410: inst = 32'h10408000;
      3411: inst = 32'hc40464c;
      3412: inst = 32'h8220000;
      3413: inst = 32'h10408000;
      3414: inst = 32'hc40464d;
      3415: inst = 32'h8220000;
      3416: inst = 32'h10408000;
      3417: inst = 32'hc40464e;
      3418: inst = 32'h8220000;
      3419: inst = 32'h10408000;
      3420: inst = 32'hc40464f;
      3421: inst = 32'h8220000;
      3422: inst = 32'h10408000;
      3423: inst = 32'hc404650;
      3424: inst = 32'h8220000;
      3425: inst = 32'h10408000;
      3426: inst = 32'hc404651;
      3427: inst = 32'h8220000;
      3428: inst = 32'h10408000;
      3429: inst = 32'hc404652;
      3430: inst = 32'h8220000;
      3431: inst = 32'h10408000;
      3432: inst = 32'hc404653;
      3433: inst = 32'h8220000;
      3434: inst = 32'h10408000;
      3435: inst = 32'hc404654;
      3436: inst = 32'h8220000;
      3437: inst = 32'h10408000;
      3438: inst = 32'hc404655;
      3439: inst = 32'h8220000;
      3440: inst = 32'h10408000;
      3441: inst = 32'hc404656;
      3442: inst = 32'h8220000;
      3443: inst = 32'h10408000;
      3444: inst = 32'hc404657;
      3445: inst = 32'h8220000;
      3446: inst = 32'h10408000;
      3447: inst = 32'hc404658;
      3448: inst = 32'h8220000;
      3449: inst = 32'h10408000;
      3450: inst = 32'hc404659;
      3451: inst = 32'h8220000;
      3452: inst = 32'h10408000;
      3453: inst = 32'hc40465a;
      3454: inst = 32'h8220000;
      3455: inst = 32'h10408000;
      3456: inst = 32'hc40465b;
      3457: inst = 32'h8220000;
      3458: inst = 32'h10408000;
      3459: inst = 32'hc404684;
      3460: inst = 32'h8220000;
      3461: inst = 32'h10408000;
      3462: inst = 32'hc404685;
      3463: inst = 32'h8220000;
      3464: inst = 32'h10408000;
      3465: inst = 32'hc404686;
      3466: inst = 32'h8220000;
      3467: inst = 32'h10408000;
      3468: inst = 32'hc404687;
      3469: inst = 32'h8220000;
      3470: inst = 32'h10408000;
      3471: inst = 32'hc404688;
      3472: inst = 32'h8220000;
      3473: inst = 32'h10408000;
      3474: inst = 32'hc404689;
      3475: inst = 32'h8220000;
      3476: inst = 32'h10408000;
      3477: inst = 32'hc40468a;
      3478: inst = 32'h8220000;
      3479: inst = 32'h10408000;
      3480: inst = 32'hc40468b;
      3481: inst = 32'h8220000;
      3482: inst = 32'h10408000;
      3483: inst = 32'hc40468c;
      3484: inst = 32'h8220000;
      3485: inst = 32'h10408000;
      3486: inst = 32'hc40468d;
      3487: inst = 32'h8220000;
      3488: inst = 32'h10408000;
      3489: inst = 32'hc40468e;
      3490: inst = 32'h8220000;
      3491: inst = 32'h10408000;
      3492: inst = 32'hc40468f;
      3493: inst = 32'h8220000;
      3494: inst = 32'h10408000;
      3495: inst = 32'hc404690;
      3496: inst = 32'h8220000;
      3497: inst = 32'h10408000;
      3498: inst = 32'hc404691;
      3499: inst = 32'h8220000;
      3500: inst = 32'h10408000;
      3501: inst = 32'hc404692;
      3502: inst = 32'h8220000;
      3503: inst = 32'h10408000;
      3504: inst = 32'hc404693;
      3505: inst = 32'h8220000;
      3506: inst = 32'h10408000;
      3507: inst = 32'hc404694;
      3508: inst = 32'h8220000;
      3509: inst = 32'h10408000;
      3510: inst = 32'hc404695;
      3511: inst = 32'h8220000;
      3512: inst = 32'h10408000;
      3513: inst = 32'hc404696;
      3514: inst = 32'h8220000;
      3515: inst = 32'h10408000;
      3516: inst = 32'hc404697;
      3517: inst = 32'h8220000;
      3518: inst = 32'h10408000;
      3519: inst = 32'hc404698;
      3520: inst = 32'h8220000;
      3521: inst = 32'h10408000;
      3522: inst = 32'hc404699;
      3523: inst = 32'h8220000;
      3524: inst = 32'h10408000;
      3525: inst = 32'hc40469a;
      3526: inst = 32'h8220000;
      3527: inst = 32'h10408000;
      3528: inst = 32'hc40469b;
      3529: inst = 32'h8220000;
      3530: inst = 32'h10408000;
      3531: inst = 32'hc40469c;
      3532: inst = 32'h8220000;
      3533: inst = 32'h10408000;
      3534: inst = 32'hc40469d;
      3535: inst = 32'h8220000;
      3536: inst = 32'h10408000;
      3537: inst = 32'hc40469e;
      3538: inst = 32'h8220000;
      3539: inst = 32'h10408000;
      3540: inst = 32'hc40469f;
      3541: inst = 32'h8220000;
      3542: inst = 32'h10408000;
      3543: inst = 32'hc4046a0;
      3544: inst = 32'h8220000;
      3545: inst = 32'h10408000;
      3546: inst = 32'hc4046a1;
      3547: inst = 32'h8220000;
      3548: inst = 32'h10408000;
      3549: inst = 32'hc4046a2;
      3550: inst = 32'h8220000;
      3551: inst = 32'h10408000;
      3552: inst = 32'hc4046a3;
      3553: inst = 32'h8220000;
      3554: inst = 32'h10408000;
      3555: inst = 32'hc4046a4;
      3556: inst = 32'h8220000;
      3557: inst = 32'h10408000;
      3558: inst = 32'hc4046a5;
      3559: inst = 32'h8220000;
      3560: inst = 32'h10408000;
      3561: inst = 32'hc4046a6;
      3562: inst = 32'h8220000;
      3563: inst = 32'h10408000;
      3564: inst = 32'hc4046a7;
      3565: inst = 32'h8220000;
      3566: inst = 32'h10408000;
      3567: inst = 32'hc4046a8;
      3568: inst = 32'h8220000;
      3569: inst = 32'h10408000;
      3570: inst = 32'hc4046a9;
      3571: inst = 32'h8220000;
      3572: inst = 32'h10408000;
      3573: inst = 32'hc4046aa;
      3574: inst = 32'h8220000;
      3575: inst = 32'h10408000;
      3576: inst = 32'hc4046ab;
      3577: inst = 32'h8220000;
      3578: inst = 32'h10408000;
      3579: inst = 32'hc4046ac;
      3580: inst = 32'h8220000;
      3581: inst = 32'h10408000;
      3582: inst = 32'hc4046ad;
      3583: inst = 32'h8220000;
      3584: inst = 32'h10408000;
      3585: inst = 32'hc4046ae;
      3586: inst = 32'h8220000;
      3587: inst = 32'h10408000;
      3588: inst = 32'hc4046af;
      3589: inst = 32'h8220000;
      3590: inst = 32'h10408000;
      3591: inst = 32'hc4046b0;
      3592: inst = 32'h8220000;
      3593: inst = 32'h10408000;
      3594: inst = 32'hc4046b1;
      3595: inst = 32'h8220000;
      3596: inst = 32'h10408000;
      3597: inst = 32'hc4046b2;
      3598: inst = 32'h8220000;
      3599: inst = 32'h10408000;
      3600: inst = 32'hc4046b3;
      3601: inst = 32'h8220000;
      3602: inst = 32'h10408000;
      3603: inst = 32'hc4046b4;
      3604: inst = 32'h8220000;
      3605: inst = 32'h10408000;
      3606: inst = 32'hc4046b5;
      3607: inst = 32'h8220000;
      3608: inst = 32'h10408000;
      3609: inst = 32'hc4046b6;
      3610: inst = 32'h8220000;
      3611: inst = 32'h10408000;
      3612: inst = 32'hc4046b7;
      3613: inst = 32'h8220000;
      3614: inst = 32'h10408000;
      3615: inst = 32'hc4046b8;
      3616: inst = 32'h8220000;
      3617: inst = 32'h10408000;
      3618: inst = 32'hc4046b9;
      3619: inst = 32'h8220000;
      3620: inst = 32'h10408000;
      3621: inst = 32'hc4046ba;
      3622: inst = 32'h8220000;
      3623: inst = 32'h10408000;
      3624: inst = 32'hc4046bb;
      3625: inst = 32'h8220000;
      3626: inst = 32'h10408000;
      3627: inst = 32'hc4046e4;
      3628: inst = 32'h8220000;
      3629: inst = 32'h10408000;
      3630: inst = 32'hc4046e5;
      3631: inst = 32'h8220000;
      3632: inst = 32'h10408000;
      3633: inst = 32'hc4046e6;
      3634: inst = 32'h8220000;
      3635: inst = 32'h10408000;
      3636: inst = 32'hc4046e7;
      3637: inst = 32'h8220000;
      3638: inst = 32'h10408000;
      3639: inst = 32'hc4046e8;
      3640: inst = 32'h8220000;
      3641: inst = 32'h10408000;
      3642: inst = 32'hc4046e9;
      3643: inst = 32'h8220000;
      3644: inst = 32'h10408000;
      3645: inst = 32'hc4046ea;
      3646: inst = 32'h8220000;
      3647: inst = 32'h10408000;
      3648: inst = 32'hc4046eb;
      3649: inst = 32'h8220000;
      3650: inst = 32'h10408000;
      3651: inst = 32'hc4046ec;
      3652: inst = 32'h8220000;
      3653: inst = 32'h10408000;
      3654: inst = 32'hc4046ed;
      3655: inst = 32'h8220000;
      3656: inst = 32'h10408000;
      3657: inst = 32'hc4046ee;
      3658: inst = 32'h8220000;
      3659: inst = 32'h10408000;
      3660: inst = 32'hc404700;
      3661: inst = 32'h8220000;
      3662: inst = 32'h10408000;
      3663: inst = 32'hc404701;
      3664: inst = 32'h8220000;
      3665: inst = 32'h10408000;
      3666: inst = 32'hc404702;
      3667: inst = 32'h8220000;
      3668: inst = 32'h10408000;
      3669: inst = 32'hc404703;
      3670: inst = 32'h8220000;
      3671: inst = 32'h10408000;
      3672: inst = 32'hc404704;
      3673: inst = 32'h8220000;
      3674: inst = 32'h10408000;
      3675: inst = 32'hc404705;
      3676: inst = 32'h8220000;
      3677: inst = 32'h10408000;
      3678: inst = 32'hc404706;
      3679: inst = 32'h8220000;
      3680: inst = 32'h10408000;
      3681: inst = 32'hc404707;
      3682: inst = 32'h8220000;
      3683: inst = 32'h10408000;
      3684: inst = 32'hc404708;
      3685: inst = 32'h8220000;
      3686: inst = 32'h10408000;
      3687: inst = 32'hc404709;
      3688: inst = 32'h8220000;
      3689: inst = 32'h10408000;
      3690: inst = 32'hc40470a;
      3691: inst = 32'h8220000;
      3692: inst = 32'h10408000;
      3693: inst = 32'hc40470b;
      3694: inst = 32'h8220000;
      3695: inst = 32'h10408000;
      3696: inst = 32'hc40470c;
      3697: inst = 32'h8220000;
      3698: inst = 32'h10408000;
      3699: inst = 32'hc40470d;
      3700: inst = 32'h8220000;
      3701: inst = 32'h10408000;
      3702: inst = 32'hc40470e;
      3703: inst = 32'h8220000;
      3704: inst = 32'h10408000;
      3705: inst = 32'hc40470f;
      3706: inst = 32'h8220000;
      3707: inst = 32'h10408000;
      3708: inst = 32'hc404710;
      3709: inst = 32'h8220000;
      3710: inst = 32'h10408000;
      3711: inst = 32'hc404711;
      3712: inst = 32'h8220000;
      3713: inst = 32'h10408000;
      3714: inst = 32'hc404712;
      3715: inst = 32'h8220000;
      3716: inst = 32'h10408000;
      3717: inst = 32'hc404713;
      3718: inst = 32'h8220000;
      3719: inst = 32'h10408000;
      3720: inst = 32'hc404714;
      3721: inst = 32'h8220000;
      3722: inst = 32'h10408000;
      3723: inst = 32'hc404715;
      3724: inst = 32'h8220000;
      3725: inst = 32'h10408000;
      3726: inst = 32'hc404716;
      3727: inst = 32'h8220000;
      3728: inst = 32'h10408000;
      3729: inst = 32'hc404717;
      3730: inst = 32'h8220000;
      3731: inst = 32'h10408000;
      3732: inst = 32'hc404718;
      3733: inst = 32'h8220000;
      3734: inst = 32'h10408000;
      3735: inst = 32'hc404719;
      3736: inst = 32'h8220000;
      3737: inst = 32'h10408000;
      3738: inst = 32'hc40471a;
      3739: inst = 32'h8220000;
      3740: inst = 32'h10408000;
      3741: inst = 32'hc40471b;
      3742: inst = 32'h8220000;
      3743: inst = 32'h10408000;
      3744: inst = 32'hc404744;
      3745: inst = 32'h8220000;
      3746: inst = 32'h10408000;
      3747: inst = 32'hc404745;
      3748: inst = 32'h8220000;
      3749: inst = 32'h10408000;
      3750: inst = 32'hc404746;
      3751: inst = 32'h8220000;
      3752: inst = 32'h10408000;
      3753: inst = 32'hc404747;
      3754: inst = 32'h8220000;
      3755: inst = 32'h10408000;
      3756: inst = 32'hc404748;
      3757: inst = 32'h8220000;
      3758: inst = 32'h10408000;
      3759: inst = 32'hc404749;
      3760: inst = 32'h8220000;
      3761: inst = 32'h10408000;
      3762: inst = 32'hc40474a;
      3763: inst = 32'h8220000;
      3764: inst = 32'h10408000;
      3765: inst = 32'hc40474b;
      3766: inst = 32'h8220000;
      3767: inst = 32'h10408000;
      3768: inst = 32'hc40474c;
      3769: inst = 32'h8220000;
      3770: inst = 32'h10408000;
      3771: inst = 32'hc40474d;
      3772: inst = 32'h8220000;
      3773: inst = 32'h10408000;
      3774: inst = 32'hc40474e;
      3775: inst = 32'h8220000;
      3776: inst = 32'h10408000;
      3777: inst = 32'hc404760;
      3778: inst = 32'h8220000;
      3779: inst = 32'h10408000;
      3780: inst = 32'hc404761;
      3781: inst = 32'h8220000;
      3782: inst = 32'h10408000;
      3783: inst = 32'hc404762;
      3784: inst = 32'h8220000;
      3785: inst = 32'h10408000;
      3786: inst = 32'hc404763;
      3787: inst = 32'h8220000;
      3788: inst = 32'h10408000;
      3789: inst = 32'hc404764;
      3790: inst = 32'h8220000;
      3791: inst = 32'h10408000;
      3792: inst = 32'hc404765;
      3793: inst = 32'h8220000;
      3794: inst = 32'h10408000;
      3795: inst = 32'hc404766;
      3796: inst = 32'h8220000;
      3797: inst = 32'h10408000;
      3798: inst = 32'hc404767;
      3799: inst = 32'h8220000;
      3800: inst = 32'h10408000;
      3801: inst = 32'hc404768;
      3802: inst = 32'h8220000;
      3803: inst = 32'h10408000;
      3804: inst = 32'hc404769;
      3805: inst = 32'h8220000;
      3806: inst = 32'h10408000;
      3807: inst = 32'hc40476a;
      3808: inst = 32'h8220000;
      3809: inst = 32'h10408000;
      3810: inst = 32'hc40476b;
      3811: inst = 32'h8220000;
      3812: inst = 32'h10408000;
      3813: inst = 32'hc40476c;
      3814: inst = 32'h8220000;
      3815: inst = 32'h10408000;
      3816: inst = 32'hc40476d;
      3817: inst = 32'h8220000;
      3818: inst = 32'h10408000;
      3819: inst = 32'hc40476e;
      3820: inst = 32'h8220000;
      3821: inst = 32'h10408000;
      3822: inst = 32'hc40476f;
      3823: inst = 32'h8220000;
      3824: inst = 32'h10408000;
      3825: inst = 32'hc404770;
      3826: inst = 32'h8220000;
      3827: inst = 32'h10408000;
      3828: inst = 32'hc404771;
      3829: inst = 32'h8220000;
      3830: inst = 32'h10408000;
      3831: inst = 32'hc404772;
      3832: inst = 32'h8220000;
      3833: inst = 32'h10408000;
      3834: inst = 32'hc404773;
      3835: inst = 32'h8220000;
      3836: inst = 32'h10408000;
      3837: inst = 32'hc404774;
      3838: inst = 32'h8220000;
      3839: inst = 32'h10408000;
      3840: inst = 32'hc404775;
      3841: inst = 32'h8220000;
      3842: inst = 32'h10408000;
      3843: inst = 32'hc404776;
      3844: inst = 32'h8220000;
      3845: inst = 32'h10408000;
      3846: inst = 32'hc404777;
      3847: inst = 32'h8220000;
      3848: inst = 32'h10408000;
      3849: inst = 32'hc404778;
      3850: inst = 32'h8220000;
      3851: inst = 32'h10408000;
      3852: inst = 32'hc404779;
      3853: inst = 32'h8220000;
      3854: inst = 32'h10408000;
      3855: inst = 32'hc40477a;
      3856: inst = 32'h8220000;
      3857: inst = 32'h10408000;
      3858: inst = 32'hc40477b;
      3859: inst = 32'h8220000;
      3860: inst = 32'h10408000;
      3861: inst = 32'hc4047a4;
      3862: inst = 32'h8220000;
      3863: inst = 32'h10408000;
      3864: inst = 32'hc4047a5;
      3865: inst = 32'h8220000;
      3866: inst = 32'h10408000;
      3867: inst = 32'hc4047a6;
      3868: inst = 32'h8220000;
      3869: inst = 32'h10408000;
      3870: inst = 32'hc4047a7;
      3871: inst = 32'h8220000;
      3872: inst = 32'h10408000;
      3873: inst = 32'hc4047a8;
      3874: inst = 32'h8220000;
      3875: inst = 32'h10408000;
      3876: inst = 32'hc4047a9;
      3877: inst = 32'h8220000;
      3878: inst = 32'h10408000;
      3879: inst = 32'hc4047aa;
      3880: inst = 32'h8220000;
      3881: inst = 32'h10408000;
      3882: inst = 32'hc4047ab;
      3883: inst = 32'h8220000;
      3884: inst = 32'h10408000;
      3885: inst = 32'hc4047ac;
      3886: inst = 32'h8220000;
      3887: inst = 32'h10408000;
      3888: inst = 32'hc4047ad;
      3889: inst = 32'h8220000;
      3890: inst = 32'h10408000;
      3891: inst = 32'hc4047ae;
      3892: inst = 32'h8220000;
      3893: inst = 32'h10408000;
      3894: inst = 32'hc4047c0;
      3895: inst = 32'h8220000;
      3896: inst = 32'h10408000;
      3897: inst = 32'hc4047c1;
      3898: inst = 32'h8220000;
      3899: inst = 32'h10408000;
      3900: inst = 32'hc4047c2;
      3901: inst = 32'h8220000;
      3902: inst = 32'h10408000;
      3903: inst = 32'hc4047c3;
      3904: inst = 32'h8220000;
      3905: inst = 32'h10408000;
      3906: inst = 32'hc4047c4;
      3907: inst = 32'h8220000;
      3908: inst = 32'h10408000;
      3909: inst = 32'hc4047c5;
      3910: inst = 32'h8220000;
      3911: inst = 32'h10408000;
      3912: inst = 32'hc4047c6;
      3913: inst = 32'h8220000;
      3914: inst = 32'h10408000;
      3915: inst = 32'hc4047c7;
      3916: inst = 32'h8220000;
      3917: inst = 32'h10408000;
      3918: inst = 32'hc4047c8;
      3919: inst = 32'h8220000;
      3920: inst = 32'h10408000;
      3921: inst = 32'hc4047c9;
      3922: inst = 32'h8220000;
      3923: inst = 32'h10408000;
      3924: inst = 32'hc4047ca;
      3925: inst = 32'h8220000;
      3926: inst = 32'h10408000;
      3927: inst = 32'hc4047cb;
      3928: inst = 32'h8220000;
      3929: inst = 32'h10408000;
      3930: inst = 32'hc4047cc;
      3931: inst = 32'h8220000;
      3932: inst = 32'h10408000;
      3933: inst = 32'hc4047cd;
      3934: inst = 32'h8220000;
      3935: inst = 32'h10408000;
      3936: inst = 32'hc4047ce;
      3937: inst = 32'h8220000;
      3938: inst = 32'h10408000;
      3939: inst = 32'hc4047cf;
      3940: inst = 32'h8220000;
      3941: inst = 32'h10408000;
      3942: inst = 32'hc4047d0;
      3943: inst = 32'h8220000;
      3944: inst = 32'h10408000;
      3945: inst = 32'hc4047d1;
      3946: inst = 32'h8220000;
      3947: inst = 32'h10408000;
      3948: inst = 32'hc4047d2;
      3949: inst = 32'h8220000;
      3950: inst = 32'h10408000;
      3951: inst = 32'hc4047d3;
      3952: inst = 32'h8220000;
      3953: inst = 32'h10408000;
      3954: inst = 32'hc4047d4;
      3955: inst = 32'h8220000;
      3956: inst = 32'h10408000;
      3957: inst = 32'hc4047d5;
      3958: inst = 32'h8220000;
      3959: inst = 32'h10408000;
      3960: inst = 32'hc4047d6;
      3961: inst = 32'h8220000;
      3962: inst = 32'h10408000;
      3963: inst = 32'hc4047d7;
      3964: inst = 32'h8220000;
      3965: inst = 32'h10408000;
      3966: inst = 32'hc4047d8;
      3967: inst = 32'h8220000;
      3968: inst = 32'h10408000;
      3969: inst = 32'hc4047d9;
      3970: inst = 32'h8220000;
      3971: inst = 32'h10408000;
      3972: inst = 32'hc4047da;
      3973: inst = 32'h8220000;
      3974: inst = 32'h10408000;
      3975: inst = 32'hc4047db;
      3976: inst = 32'h8220000;
      3977: inst = 32'h10408000;
      3978: inst = 32'hc404804;
      3979: inst = 32'h8220000;
      3980: inst = 32'h10408000;
      3981: inst = 32'hc404805;
      3982: inst = 32'h8220000;
      3983: inst = 32'h10408000;
      3984: inst = 32'hc404806;
      3985: inst = 32'h8220000;
      3986: inst = 32'h10408000;
      3987: inst = 32'hc404807;
      3988: inst = 32'h8220000;
      3989: inst = 32'h10408000;
      3990: inst = 32'hc404808;
      3991: inst = 32'h8220000;
      3992: inst = 32'h10408000;
      3993: inst = 32'hc404809;
      3994: inst = 32'h8220000;
      3995: inst = 32'h10408000;
      3996: inst = 32'hc40480a;
      3997: inst = 32'h8220000;
      3998: inst = 32'h10408000;
      3999: inst = 32'hc40480b;
      4000: inst = 32'h8220000;
      4001: inst = 32'h10408000;
      4002: inst = 32'hc40480c;
      4003: inst = 32'h8220000;
      4004: inst = 32'h10408000;
      4005: inst = 32'hc40480d;
      4006: inst = 32'h8220000;
      4007: inst = 32'h10408000;
      4008: inst = 32'hc40480e;
      4009: inst = 32'h8220000;
      4010: inst = 32'h10408000;
      4011: inst = 32'hc404820;
      4012: inst = 32'h8220000;
      4013: inst = 32'h10408000;
      4014: inst = 32'hc404821;
      4015: inst = 32'h8220000;
      4016: inst = 32'h10408000;
      4017: inst = 32'hc404822;
      4018: inst = 32'h8220000;
      4019: inst = 32'h10408000;
      4020: inst = 32'hc404823;
      4021: inst = 32'h8220000;
      4022: inst = 32'h10408000;
      4023: inst = 32'hc404824;
      4024: inst = 32'h8220000;
      4025: inst = 32'h10408000;
      4026: inst = 32'hc404825;
      4027: inst = 32'h8220000;
      4028: inst = 32'h10408000;
      4029: inst = 32'hc404826;
      4030: inst = 32'h8220000;
      4031: inst = 32'h10408000;
      4032: inst = 32'hc404827;
      4033: inst = 32'h8220000;
      4034: inst = 32'h10408000;
      4035: inst = 32'hc404828;
      4036: inst = 32'h8220000;
      4037: inst = 32'h10408000;
      4038: inst = 32'hc404829;
      4039: inst = 32'h8220000;
      4040: inst = 32'h10408000;
      4041: inst = 32'hc40482a;
      4042: inst = 32'h8220000;
      4043: inst = 32'h10408000;
      4044: inst = 32'hc40482b;
      4045: inst = 32'h8220000;
      4046: inst = 32'h10408000;
      4047: inst = 32'hc40482c;
      4048: inst = 32'h8220000;
      4049: inst = 32'h10408000;
      4050: inst = 32'hc40482d;
      4051: inst = 32'h8220000;
      4052: inst = 32'h10408000;
      4053: inst = 32'hc40482e;
      4054: inst = 32'h8220000;
      4055: inst = 32'h10408000;
      4056: inst = 32'hc40482f;
      4057: inst = 32'h8220000;
      4058: inst = 32'h10408000;
      4059: inst = 32'hc404830;
      4060: inst = 32'h8220000;
      4061: inst = 32'h10408000;
      4062: inst = 32'hc404831;
      4063: inst = 32'h8220000;
      4064: inst = 32'h10408000;
      4065: inst = 32'hc404832;
      4066: inst = 32'h8220000;
      4067: inst = 32'h10408000;
      4068: inst = 32'hc404833;
      4069: inst = 32'h8220000;
      4070: inst = 32'h10408000;
      4071: inst = 32'hc404834;
      4072: inst = 32'h8220000;
      4073: inst = 32'h10408000;
      4074: inst = 32'hc404835;
      4075: inst = 32'h8220000;
      4076: inst = 32'h10408000;
      4077: inst = 32'hc404836;
      4078: inst = 32'h8220000;
      4079: inst = 32'h10408000;
      4080: inst = 32'hc404837;
      4081: inst = 32'h8220000;
      4082: inst = 32'h10408000;
      4083: inst = 32'hc404838;
      4084: inst = 32'h8220000;
      4085: inst = 32'h10408000;
      4086: inst = 32'hc404839;
      4087: inst = 32'h8220000;
      4088: inst = 32'h10408000;
      4089: inst = 32'hc40483a;
      4090: inst = 32'h8220000;
      4091: inst = 32'h10408000;
      4092: inst = 32'hc40483b;
      4093: inst = 32'h8220000;
      4094: inst = 32'h10408000;
      4095: inst = 32'hc404864;
      4096: inst = 32'h8220000;
      4097: inst = 32'h10408000;
      4098: inst = 32'hc404865;
      4099: inst = 32'h8220000;
      4100: inst = 32'h10408000;
      4101: inst = 32'hc404866;
      4102: inst = 32'h8220000;
      4103: inst = 32'h10408000;
      4104: inst = 32'hc404867;
      4105: inst = 32'h8220000;
      4106: inst = 32'h10408000;
      4107: inst = 32'hc404868;
      4108: inst = 32'h8220000;
      4109: inst = 32'h10408000;
      4110: inst = 32'hc404869;
      4111: inst = 32'h8220000;
      4112: inst = 32'h10408000;
      4113: inst = 32'hc40486a;
      4114: inst = 32'h8220000;
      4115: inst = 32'h10408000;
      4116: inst = 32'hc40486b;
      4117: inst = 32'h8220000;
      4118: inst = 32'h10408000;
      4119: inst = 32'hc40486c;
      4120: inst = 32'h8220000;
      4121: inst = 32'h10408000;
      4122: inst = 32'hc40486d;
      4123: inst = 32'h8220000;
      4124: inst = 32'h10408000;
      4125: inst = 32'hc40486e;
      4126: inst = 32'h8220000;
      4127: inst = 32'h10408000;
      4128: inst = 32'hc404880;
      4129: inst = 32'h8220000;
      4130: inst = 32'h10408000;
      4131: inst = 32'hc404881;
      4132: inst = 32'h8220000;
      4133: inst = 32'h10408000;
      4134: inst = 32'hc404882;
      4135: inst = 32'h8220000;
      4136: inst = 32'h10408000;
      4137: inst = 32'hc404883;
      4138: inst = 32'h8220000;
      4139: inst = 32'h10408000;
      4140: inst = 32'hc404884;
      4141: inst = 32'h8220000;
      4142: inst = 32'h10408000;
      4143: inst = 32'hc404885;
      4144: inst = 32'h8220000;
      4145: inst = 32'h10408000;
      4146: inst = 32'hc404886;
      4147: inst = 32'h8220000;
      4148: inst = 32'h10408000;
      4149: inst = 32'hc404887;
      4150: inst = 32'h8220000;
      4151: inst = 32'h10408000;
      4152: inst = 32'hc404888;
      4153: inst = 32'h8220000;
      4154: inst = 32'h10408000;
      4155: inst = 32'hc404889;
      4156: inst = 32'h8220000;
      4157: inst = 32'h10408000;
      4158: inst = 32'hc40488a;
      4159: inst = 32'h8220000;
      4160: inst = 32'h10408000;
      4161: inst = 32'hc40488b;
      4162: inst = 32'h8220000;
      4163: inst = 32'h10408000;
      4164: inst = 32'hc40488c;
      4165: inst = 32'h8220000;
      4166: inst = 32'h10408000;
      4167: inst = 32'hc40488d;
      4168: inst = 32'h8220000;
      4169: inst = 32'h10408000;
      4170: inst = 32'hc40488e;
      4171: inst = 32'h8220000;
      4172: inst = 32'h10408000;
      4173: inst = 32'hc40488f;
      4174: inst = 32'h8220000;
      4175: inst = 32'h10408000;
      4176: inst = 32'hc404890;
      4177: inst = 32'h8220000;
      4178: inst = 32'h10408000;
      4179: inst = 32'hc404891;
      4180: inst = 32'h8220000;
      4181: inst = 32'h10408000;
      4182: inst = 32'hc404892;
      4183: inst = 32'h8220000;
      4184: inst = 32'h10408000;
      4185: inst = 32'hc404893;
      4186: inst = 32'h8220000;
      4187: inst = 32'h10408000;
      4188: inst = 32'hc404894;
      4189: inst = 32'h8220000;
      4190: inst = 32'h10408000;
      4191: inst = 32'hc404895;
      4192: inst = 32'h8220000;
      4193: inst = 32'h10408000;
      4194: inst = 32'hc404896;
      4195: inst = 32'h8220000;
      4196: inst = 32'h10408000;
      4197: inst = 32'hc404897;
      4198: inst = 32'h8220000;
      4199: inst = 32'h10408000;
      4200: inst = 32'hc404898;
      4201: inst = 32'h8220000;
      4202: inst = 32'h10408000;
      4203: inst = 32'hc404899;
      4204: inst = 32'h8220000;
      4205: inst = 32'h10408000;
      4206: inst = 32'hc40489a;
      4207: inst = 32'h8220000;
      4208: inst = 32'h10408000;
      4209: inst = 32'hc40489b;
      4210: inst = 32'h8220000;
      4211: inst = 32'h10408000;
      4212: inst = 32'hc4048c4;
      4213: inst = 32'h8220000;
      4214: inst = 32'h10408000;
      4215: inst = 32'hc4048c5;
      4216: inst = 32'h8220000;
      4217: inst = 32'h10408000;
      4218: inst = 32'hc4048c6;
      4219: inst = 32'h8220000;
      4220: inst = 32'h10408000;
      4221: inst = 32'hc4048c7;
      4222: inst = 32'h8220000;
      4223: inst = 32'h10408000;
      4224: inst = 32'hc4048c8;
      4225: inst = 32'h8220000;
      4226: inst = 32'h10408000;
      4227: inst = 32'hc4048c9;
      4228: inst = 32'h8220000;
      4229: inst = 32'h10408000;
      4230: inst = 32'hc4048ca;
      4231: inst = 32'h8220000;
      4232: inst = 32'h10408000;
      4233: inst = 32'hc4048cb;
      4234: inst = 32'h8220000;
      4235: inst = 32'h10408000;
      4236: inst = 32'hc4048cc;
      4237: inst = 32'h8220000;
      4238: inst = 32'h10408000;
      4239: inst = 32'hc4048cd;
      4240: inst = 32'h8220000;
      4241: inst = 32'h10408000;
      4242: inst = 32'hc4048ce;
      4243: inst = 32'h8220000;
      4244: inst = 32'h10408000;
      4245: inst = 32'hc4048e0;
      4246: inst = 32'h8220000;
      4247: inst = 32'h10408000;
      4248: inst = 32'hc4048e1;
      4249: inst = 32'h8220000;
      4250: inst = 32'h10408000;
      4251: inst = 32'hc4048e2;
      4252: inst = 32'h8220000;
      4253: inst = 32'h10408000;
      4254: inst = 32'hc4048e3;
      4255: inst = 32'h8220000;
      4256: inst = 32'h10408000;
      4257: inst = 32'hc4048e4;
      4258: inst = 32'h8220000;
      4259: inst = 32'h10408000;
      4260: inst = 32'hc4048e5;
      4261: inst = 32'h8220000;
      4262: inst = 32'h10408000;
      4263: inst = 32'hc4048e6;
      4264: inst = 32'h8220000;
      4265: inst = 32'h10408000;
      4266: inst = 32'hc4048e7;
      4267: inst = 32'h8220000;
      4268: inst = 32'h10408000;
      4269: inst = 32'hc4048e8;
      4270: inst = 32'h8220000;
      4271: inst = 32'h10408000;
      4272: inst = 32'hc4048e9;
      4273: inst = 32'h8220000;
      4274: inst = 32'h10408000;
      4275: inst = 32'hc4048ea;
      4276: inst = 32'h8220000;
      4277: inst = 32'h10408000;
      4278: inst = 32'hc4048eb;
      4279: inst = 32'h8220000;
      4280: inst = 32'h10408000;
      4281: inst = 32'hc4048ec;
      4282: inst = 32'h8220000;
      4283: inst = 32'h10408000;
      4284: inst = 32'hc4048ed;
      4285: inst = 32'h8220000;
      4286: inst = 32'h10408000;
      4287: inst = 32'hc4048ee;
      4288: inst = 32'h8220000;
      4289: inst = 32'h10408000;
      4290: inst = 32'hc4048ef;
      4291: inst = 32'h8220000;
      4292: inst = 32'h10408000;
      4293: inst = 32'hc4048f0;
      4294: inst = 32'h8220000;
      4295: inst = 32'h10408000;
      4296: inst = 32'hc4048f1;
      4297: inst = 32'h8220000;
      4298: inst = 32'h10408000;
      4299: inst = 32'hc4048f2;
      4300: inst = 32'h8220000;
      4301: inst = 32'h10408000;
      4302: inst = 32'hc4048f3;
      4303: inst = 32'h8220000;
      4304: inst = 32'h10408000;
      4305: inst = 32'hc4048f4;
      4306: inst = 32'h8220000;
      4307: inst = 32'h10408000;
      4308: inst = 32'hc4048f5;
      4309: inst = 32'h8220000;
      4310: inst = 32'h10408000;
      4311: inst = 32'hc4048f6;
      4312: inst = 32'h8220000;
      4313: inst = 32'h10408000;
      4314: inst = 32'hc4048f7;
      4315: inst = 32'h8220000;
      4316: inst = 32'h10408000;
      4317: inst = 32'hc4048f8;
      4318: inst = 32'h8220000;
      4319: inst = 32'h10408000;
      4320: inst = 32'hc4048f9;
      4321: inst = 32'h8220000;
      4322: inst = 32'h10408000;
      4323: inst = 32'hc4048fa;
      4324: inst = 32'h8220000;
      4325: inst = 32'h10408000;
      4326: inst = 32'hc4048fb;
      4327: inst = 32'h8220000;
      4328: inst = 32'h10408000;
      4329: inst = 32'hc404924;
      4330: inst = 32'h8220000;
      4331: inst = 32'h10408000;
      4332: inst = 32'hc404925;
      4333: inst = 32'h8220000;
      4334: inst = 32'h10408000;
      4335: inst = 32'hc404926;
      4336: inst = 32'h8220000;
      4337: inst = 32'h10408000;
      4338: inst = 32'hc404927;
      4339: inst = 32'h8220000;
      4340: inst = 32'h10408000;
      4341: inst = 32'hc404928;
      4342: inst = 32'h8220000;
      4343: inst = 32'h10408000;
      4344: inst = 32'hc404929;
      4345: inst = 32'h8220000;
      4346: inst = 32'h10408000;
      4347: inst = 32'hc40492a;
      4348: inst = 32'h8220000;
      4349: inst = 32'h10408000;
      4350: inst = 32'hc40492b;
      4351: inst = 32'h8220000;
      4352: inst = 32'h10408000;
      4353: inst = 32'hc40492c;
      4354: inst = 32'h8220000;
      4355: inst = 32'h10408000;
      4356: inst = 32'hc40492d;
      4357: inst = 32'h8220000;
      4358: inst = 32'h10408000;
      4359: inst = 32'hc40492e;
      4360: inst = 32'h8220000;
      4361: inst = 32'h10408000;
      4362: inst = 32'hc404940;
      4363: inst = 32'h8220000;
      4364: inst = 32'h10408000;
      4365: inst = 32'hc404941;
      4366: inst = 32'h8220000;
      4367: inst = 32'h10408000;
      4368: inst = 32'hc404942;
      4369: inst = 32'h8220000;
      4370: inst = 32'h10408000;
      4371: inst = 32'hc404943;
      4372: inst = 32'h8220000;
      4373: inst = 32'h10408000;
      4374: inst = 32'hc404944;
      4375: inst = 32'h8220000;
      4376: inst = 32'h10408000;
      4377: inst = 32'hc404945;
      4378: inst = 32'h8220000;
      4379: inst = 32'h10408000;
      4380: inst = 32'hc404946;
      4381: inst = 32'h8220000;
      4382: inst = 32'h10408000;
      4383: inst = 32'hc404947;
      4384: inst = 32'h8220000;
      4385: inst = 32'h10408000;
      4386: inst = 32'hc404948;
      4387: inst = 32'h8220000;
      4388: inst = 32'h10408000;
      4389: inst = 32'hc404949;
      4390: inst = 32'h8220000;
      4391: inst = 32'h10408000;
      4392: inst = 32'hc40494a;
      4393: inst = 32'h8220000;
      4394: inst = 32'h10408000;
      4395: inst = 32'hc40494b;
      4396: inst = 32'h8220000;
      4397: inst = 32'h10408000;
      4398: inst = 32'hc40494c;
      4399: inst = 32'h8220000;
      4400: inst = 32'h10408000;
      4401: inst = 32'hc40494d;
      4402: inst = 32'h8220000;
      4403: inst = 32'h10408000;
      4404: inst = 32'hc40494e;
      4405: inst = 32'h8220000;
      4406: inst = 32'h10408000;
      4407: inst = 32'hc40494f;
      4408: inst = 32'h8220000;
      4409: inst = 32'h10408000;
      4410: inst = 32'hc404950;
      4411: inst = 32'h8220000;
      4412: inst = 32'h10408000;
      4413: inst = 32'hc404951;
      4414: inst = 32'h8220000;
      4415: inst = 32'h10408000;
      4416: inst = 32'hc404952;
      4417: inst = 32'h8220000;
      4418: inst = 32'h10408000;
      4419: inst = 32'hc404953;
      4420: inst = 32'h8220000;
      4421: inst = 32'h10408000;
      4422: inst = 32'hc404954;
      4423: inst = 32'h8220000;
      4424: inst = 32'h10408000;
      4425: inst = 32'hc404955;
      4426: inst = 32'h8220000;
      4427: inst = 32'h10408000;
      4428: inst = 32'hc404956;
      4429: inst = 32'h8220000;
      4430: inst = 32'h10408000;
      4431: inst = 32'hc404957;
      4432: inst = 32'h8220000;
      4433: inst = 32'h10408000;
      4434: inst = 32'hc404958;
      4435: inst = 32'h8220000;
      4436: inst = 32'h10408000;
      4437: inst = 32'hc404959;
      4438: inst = 32'h8220000;
      4439: inst = 32'h10408000;
      4440: inst = 32'hc40495a;
      4441: inst = 32'h8220000;
      4442: inst = 32'h10408000;
      4443: inst = 32'hc40495b;
      4444: inst = 32'h8220000;
      4445: inst = 32'h10408000;
      4446: inst = 32'hc404984;
      4447: inst = 32'h8220000;
      4448: inst = 32'h10408000;
      4449: inst = 32'hc404985;
      4450: inst = 32'h8220000;
      4451: inst = 32'h10408000;
      4452: inst = 32'hc404986;
      4453: inst = 32'h8220000;
      4454: inst = 32'h10408000;
      4455: inst = 32'hc404987;
      4456: inst = 32'h8220000;
      4457: inst = 32'h10408000;
      4458: inst = 32'hc404988;
      4459: inst = 32'h8220000;
      4460: inst = 32'h10408000;
      4461: inst = 32'hc404989;
      4462: inst = 32'h8220000;
      4463: inst = 32'h10408000;
      4464: inst = 32'hc40498a;
      4465: inst = 32'h8220000;
      4466: inst = 32'h10408000;
      4467: inst = 32'hc40498b;
      4468: inst = 32'h8220000;
      4469: inst = 32'h10408000;
      4470: inst = 32'hc40498c;
      4471: inst = 32'h8220000;
      4472: inst = 32'h10408000;
      4473: inst = 32'hc40498d;
      4474: inst = 32'h8220000;
      4475: inst = 32'h10408000;
      4476: inst = 32'hc40498e;
      4477: inst = 32'h8220000;
      4478: inst = 32'h10408000;
      4479: inst = 32'hc4049a0;
      4480: inst = 32'h8220000;
      4481: inst = 32'h10408000;
      4482: inst = 32'hc4049a1;
      4483: inst = 32'h8220000;
      4484: inst = 32'h10408000;
      4485: inst = 32'hc4049a2;
      4486: inst = 32'h8220000;
      4487: inst = 32'h10408000;
      4488: inst = 32'hc4049a3;
      4489: inst = 32'h8220000;
      4490: inst = 32'h10408000;
      4491: inst = 32'hc4049a4;
      4492: inst = 32'h8220000;
      4493: inst = 32'h10408000;
      4494: inst = 32'hc4049a5;
      4495: inst = 32'h8220000;
      4496: inst = 32'h10408000;
      4497: inst = 32'hc4049a6;
      4498: inst = 32'h8220000;
      4499: inst = 32'h10408000;
      4500: inst = 32'hc4049a7;
      4501: inst = 32'h8220000;
      4502: inst = 32'h10408000;
      4503: inst = 32'hc4049a8;
      4504: inst = 32'h8220000;
      4505: inst = 32'h10408000;
      4506: inst = 32'hc4049a9;
      4507: inst = 32'h8220000;
      4508: inst = 32'h10408000;
      4509: inst = 32'hc4049aa;
      4510: inst = 32'h8220000;
      4511: inst = 32'h10408000;
      4512: inst = 32'hc4049ab;
      4513: inst = 32'h8220000;
      4514: inst = 32'h10408000;
      4515: inst = 32'hc4049ac;
      4516: inst = 32'h8220000;
      4517: inst = 32'h10408000;
      4518: inst = 32'hc4049ad;
      4519: inst = 32'h8220000;
      4520: inst = 32'h10408000;
      4521: inst = 32'hc4049ae;
      4522: inst = 32'h8220000;
      4523: inst = 32'h10408000;
      4524: inst = 32'hc4049af;
      4525: inst = 32'h8220000;
      4526: inst = 32'h10408000;
      4527: inst = 32'hc4049b0;
      4528: inst = 32'h8220000;
      4529: inst = 32'h10408000;
      4530: inst = 32'hc4049b1;
      4531: inst = 32'h8220000;
      4532: inst = 32'h10408000;
      4533: inst = 32'hc4049b2;
      4534: inst = 32'h8220000;
      4535: inst = 32'h10408000;
      4536: inst = 32'hc4049b3;
      4537: inst = 32'h8220000;
      4538: inst = 32'h10408000;
      4539: inst = 32'hc4049b4;
      4540: inst = 32'h8220000;
      4541: inst = 32'h10408000;
      4542: inst = 32'hc4049b5;
      4543: inst = 32'h8220000;
      4544: inst = 32'h10408000;
      4545: inst = 32'hc4049b6;
      4546: inst = 32'h8220000;
      4547: inst = 32'h10408000;
      4548: inst = 32'hc4049b7;
      4549: inst = 32'h8220000;
      4550: inst = 32'h10408000;
      4551: inst = 32'hc4049b8;
      4552: inst = 32'h8220000;
      4553: inst = 32'h10408000;
      4554: inst = 32'hc4049b9;
      4555: inst = 32'h8220000;
      4556: inst = 32'h10408000;
      4557: inst = 32'hc4049ba;
      4558: inst = 32'h8220000;
      4559: inst = 32'h10408000;
      4560: inst = 32'hc4049bb;
      4561: inst = 32'h8220000;
      4562: inst = 32'h10408000;
      4563: inst = 32'hc4049e4;
      4564: inst = 32'h8220000;
      4565: inst = 32'h10408000;
      4566: inst = 32'hc4049e5;
      4567: inst = 32'h8220000;
      4568: inst = 32'h10408000;
      4569: inst = 32'hc4049e6;
      4570: inst = 32'h8220000;
      4571: inst = 32'h10408000;
      4572: inst = 32'hc4049e7;
      4573: inst = 32'h8220000;
      4574: inst = 32'h10408000;
      4575: inst = 32'hc4049e8;
      4576: inst = 32'h8220000;
      4577: inst = 32'h10408000;
      4578: inst = 32'hc4049e9;
      4579: inst = 32'h8220000;
      4580: inst = 32'h10408000;
      4581: inst = 32'hc4049ea;
      4582: inst = 32'h8220000;
      4583: inst = 32'h10408000;
      4584: inst = 32'hc4049eb;
      4585: inst = 32'h8220000;
      4586: inst = 32'h10408000;
      4587: inst = 32'hc4049ec;
      4588: inst = 32'h8220000;
      4589: inst = 32'h10408000;
      4590: inst = 32'hc4049ed;
      4591: inst = 32'h8220000;
      4592: inst = 32'h10408000;
      4593: inst = 32'hc4049ee;
      4594: inst = 32'h8220000;
      4595: inst = 32'h10408000;
      4596: inst = 32'hc404a00;
      4597: inst = 32'h8220000;
      4598: inst = 32'h10408000;
      4599: inst = 32'hc404a01;
      4600: inst = 32'h8220000;
      4601: inst = 32'h10408000;
      4602: inst = 32'hc404a02;
      4603: inst = 32'h8220000;
      4604: inst = 32'h10408000;
      4605: inst = 32'hc404a03;
      4606: inst = 32'h8220000;
      4607: inst = 32'h10408000;
      4608: inst = 32'hc404a04;
      4609: inst = 32'h8220000;
      4610: inst = 32'h10408000;
      4611: inst = 32'hc404a05;
      4612: inst = 32'h8220000;
      4613: inst = 32'h10408000;
      4614: inst = 32'hc404a06;
      4615: inst = 32'h8220000;
      4616: inst = 32'h10408000;
      4617: inst = 32'hc404a07;
      4618: inst = 32'h8220000;
      4619: inst = 32'h10408000;
      4620: inst = 32'hc404a0f;
      4621: inst = 32'h8220000;
      4622: inst = 32'h10408000;
      4623: inst = 32'hc404a10;
      4624: inst = 32'h8220000;
      4625: inst = 32'h10408000;
      4626: inst = 32'hc404a11;
      4627: inst = 32'h8220000;
      4628: inst = 32'h10408000;
      4629: inst = 32'hc404a12;
      4630: inst = 32'h8220000;
      4631: inst = 32'h10408000;
      4632: inst = 32'hc404a13;
      4633: inst = 32'h8220000;
      4634: inst = 32'h10408000;
      4635: inst = 32'hc404a14;
      4636: inst = 32'h8220000;
      4637: inst = 32'h10408000;
      4638: inst = 32'hc404a15;
      4639: inst = 32'h8220000;
      4640: inst = 32'h10408000;
      4641: inst = 32'hc404a16;
      4642: inst = 32'h8220000;
      4643: inst = 32'h10408000;
      4644: inst = 32'hc404a17;
      4645: inst = 32'h8220000;
      4646: inst = 32'h10408000;
      4647: inst = 32'hc404a18;
      4648: inst = 32'h8220000;
      4649: inst = 32'h10408000;
      4650: inst = 32'hc404a19;
      4651: inst = 32'h8220000;
      4652: inst = 32'h10408000;
      4653: inst = 32'hc404a1a;
      4654: inst = 32'h8220000;
      4655: inst = 32'h10408000;
      4656: inst = 32'hc404a1b;
      4657: inst = 32'h8220000;
      4658: inst = 32'h10408000;
      4659: inst = 32'hc404a44;
      4660: inst = 32'h8220000;
      4661: inst = 32'h10408000;
      4662: inst = 32'hc404a45;
      4663: inst = 32'h8220000;
      4664: inst = 32'h10408000;
      4665: inst = 32'hc404a46;
      4666: inst = 32'h8220000;
      4667: inst = 32'h10408000;
      4668: inst = 32'hc404a47;
      4669: inst = 32'h8220000;
      4670: inst = 32'h10408000;
      4671: inst = 32'hc404a48;
      4672: inst = 32'h8220000;
      4673: inst = 32'h10408000;
      4674: inst = 32'hc404a49;
      4675: inst = 32'h8220000;
      4676: inst = 32'h10408000;
      4677: inst = 32'hc404a4a;
      4678: inst = 32'h8220000;
      4679: inst = 32'h10408000;
      4680: inst = 32'hc404a4b;
      4681: inst = 32'h8220000;
      4682: inst = 32'h10408000;
      4683: inst = 32'hc404a4c;
      4684: inst = 32'h8220000;
      4685: inst = 32'h10408000;
      4686: inst = 32'hc404a4d;
      4687: inst = 32'h8220000;
      4688: inst = 32'h10408000;
      4689: inst = 32'hc404a4e;
      4690: inst = 32'h8220000;
      4691: inst = 32'h10408000;
      4692: inst = 32'hc404a60;
      4693: inst = 32'h8220000;
      4694: inst = 32'h10408000;
      4695: inst = 32'hc404a61;
      4696: inst = 32'h8220000;
      4697: inst = 32'h10408000;
      4698: inst = 32'hc404a62;
      4699: inst = 32'h8220000;
      4700: inst = 32'h10408000;
      4701: inst = 32'hc404a63;
      4702: inst = 32'h8220000;
      4703: inst = 32'h10408000;
      4704: inst = 32'hc404a64;
      4705: inst = 32'h8220000;
      4706: inst = 32'h10408000;
      4707: inst = 32'hc404a65;
      4708: inst = 32'h8220000;
      4709: inst = 32'h10408000;
      4710: inst = 32'hc404a66;
      4711: inst = 32'h8220000;
      4712: inst = 32'h10408000;
      4713: inst = 32'hc404a70;
      4714: inst = 32'h8220000;
      4715: inst = 32'h10408000;
      4716: inst = 32'hc404a71;
      4717: inst = 32'h8220000;
      4718: inst = 32'h10408000;
      4719: inst = 32'hc404a72;
      4720: inst = 32'h8220000;
      4721: inst = 32'h10408000;
      4722: inst = 32'hc404a73;
      4723: inst = 32'h8220000;
      4724: inst = 32'h10408000;
      4725: inst = 32'hc404a74;
      4726: inst = 32'h8220000;
      4727: inst = 32'h10408000;
      4728: inst = 32'hc404a75;
      4729: inst = 32'h8220000;
      4730: inst = 32'h10408000;
      4731: inst = 32'hc404a76;
      4732: inst = 32'h8220000;
      4733: inst = 32'h10408000;
      4734: inst = 32'hc404a77;
      4735: inst = 32'h8220000;
      4736: inst = 32'h10408000;
      4737: inst = 32'hc404a78;
      4738: inst = 32'h8220000;
      4739: inst = 32'h10408000;
      4740: inst = 32'hc404a79;
      4741: inst = 32'h8220000;
      4742: inst = 32'h10408000;
      4743: inst = 32'hc404a7a;
      4744: inst = 32'h8220000;
      4745: inst = 32'h10408000;
      4746: inst = 32'hc404a7b;
      4747: inst = 32'h8220000;
      4748: inst = 32'h10408000;
      4749: inst = 32'hc404aa4;
      4750: inst = 32'h8220000;
      4751: inst = 32'h10408000;
      4752: inst = 32'hc404aa5;
      4753: inst = 32'h8220000;
      4754: inst = 32'h10408000;
      4755: inst = 32'hc404aa6;
      4756: inst = 32'h8220000;
      4757: inst = 32'h10408000;
      4758: inst = 32'hc404aa7;
      4759: inst = 32'h8220000;
      4760: inst = 32'h10408000;
      4761: inst = 32'hc404aa8;
      4762: inst = 32'h8220000;
      4763: inst = 32'h10408000;
      4764: inst = 32'hc404aa9;
      4765: inst = 32'h8220000;
      4766: inst = 32'h10408000;
      4767: inst = 32'hc404aaa;
      4768: inst = 32'h8220000;
      4769: inst = 32'h10408000;
      4770: inst = 32'hc404aab;
      4771: inst = 32'h8220000;
      4772: inst = 32'h10408000;
      4773: inst = 32'hc404aac;
      4774: inst = 32'h8220000;
      4775: inst = 32'h10408000;
      4776: inst = 32'hc404aad;
      4777: inst = 32'h8220000;
      4778: inst = 32'h10408000;
      4779: inst = 32'hc404aae;
      4780: inst = 32'h8220000;
      4781: inst = 32'h10408000;
      4782: inst = 32'hc404ac0;
      4783: inst = 32'h8220000;
      4784: inst = 32'h10408000;
      4785: inst = 32'hc404ac1;
      4786: inst = 32'h8220000;
      4787: inst = 32'h10408000;
      4788: inst = 32'hc404ac2;
      4789: inst = 32'h8220000;
      4790: inst = 32'h10408000;
      4791: inst = 32'hc404ac3;
      4792: inst = 32'h8220000;
      4793: inst = 32'h10408000;
      4794: inst = 32'hc404ac4;
      4795: inst = 32'h8220000;
      4796: inst = 32'h10408000;
      4797: inst = 32'hc404ac5;
      4798: inst = 32'h8220000;
      4799: inst = 32'h10408000;
      4800: inst = 32'hc404ac6;
      4801: inst = 32'h8220000;
      4802: inst = 32'h10408000;
      4803: inst = 32'hc404ad0;
      4804: inst = 32'h8220000;
      4805: inst = 32'h10408000;
      4806: inst = 32'hc404ad1;
      4807: inst = 32'h8220000;
      4808: inst = 32'h10408000;
      4809: inst = 32'hc404ad2;
      4810: inst = 32'h8220000;
      4811: inst = 32'h10408000;
      4812: inst = 32'hc404ad3;
      4813: inst = 32'h8220000;
      4814: inst = 32'h10408000;
      4815: inst = 32'hc404ad4;
      4816: inst = 32'h8220000;
      4817: inst = 32'h10408000;
      4818: inst = 32'hc404ad5;
      4819: inst = 32'h8220000;
      4820: inst = 32'h10408000;
      4821: inst = 32'hc404ad6;
      4822: inst = 32'h8220000;
      4823: inst = 32'h10408000;
      4824: inst = 32'hc404ad7;
      4825: inst = 32'h8220000;
      4826: inst = 32'h10408000;
      4827: inst = 32'hc404ad8;
      4828: inst = 32'h8220000;
      4829: inst = 32'h10408000;
      4830: inst = 32'hc404ad9;
      4831: inst = 32'h8220000;
      4832: inst = 32'h10408000;
      4833: inst = 32'hc404ada;
      4834: inst = 32'h8220000;
      4835: inst = 32'h10408000;
      4836: inst = 32'hc404adb;
      4837: inst = 32'h8220000;
      4838: inst = 32'h10408000;
      4839: inst = 32'hc404b04;
      4840: inst = 32'h8220000;
      4841: inst = 32'h10408000;
      4842: inst = 32'hc404b05;
      4843: inst = 32'h8220000;
      4844: inst = 32'h10408000;
      4845: inst = 32'hc404b06;
      4846: inst = 32'h8220000;
      4847: inst = 32'h10408000;
      4848: inst = 32'hc404b07;
      4849: inst = 32'h8220000;
      4850: inst = 32'h10408000;
      4851: inst = 32'hc404b08;
      4852: inst = 32'h8220000;
      4853: inst = 32'h10408000;
      4854: inst = 32'hc404b09;
      4855: inst = 32'h8220000;
      4856: inst = 32'h10408000;
      4857: inst = 32'hc404b0a;
      4858: inst = 32'h8220000;
      4859: inst = 32'h10408000;
      4860: inst = 32'hc404b0b;
      4861: inst = 32'h8220000;
      4862: inst = 32'h10408000;
      4863: inst = 32'hc404b0c;
      4864: inst = 32'h8220000;
      4865: inst = 32'h10408000;
      4866: inst = 32'hc404b0d;
      4867: inst = 32'h8220000;
      4868: inst = 32'h10408000;
      4869: inst = 32'hc404b0e;
      4870: inst = 32'h8220000;
      4871: inst = 32'h10408000;
      4872: inst = 32'hc404b20;
      4873: inst = 32'h8220000;
      4874: inst = 32'h10408000;
      4875: inst = 32'hc404b21;
      4876: inst = 32'h8220000;
      4877: inst = 32'h10408000;
      4878: inst = 32'hc404b22;
      4879: inst = 32'h8220000;
      4880: inst = 32'h10408000;
      4881: inst = 32'hc404b23;
      4882: inst = 32'h8220000;
      4883: inst = 32'h10408000;
      4884: inst = 32'hc404b24;
      4885: inst = 32'h8220000;
      4886: inst = 32'h10408000;
      4887: inst = 32'hc404b25;
      4888: inst = 32'h8220000;
      4889: inst = 32'h10408000;
      4890: inst = 32'hc404b26;
      4891: inst = 32'h8220000;
      4892: inst = 32'h10408000;
      4893: inst = 32'hc404b30;
      4894: inst = 32'h8220000;
      4895: inst = 32'h10408000;
      4896: inst = 32'hc404b31;
      4897: inst = 32'h8220000;
      4898: inst = 32'h10408000;
      4899: inst = 32'hc404b32;
      4900: inst = 32'h8220000;
      4901: inst = 32'h10408000;
      4902: inst = 32'hc404b33;
      4903: inst = 32'h8220000;
      4904: inst = 32'h10408000;
      4905: inst = 32'hc404b34;
      4906: inst = 32'h8220000;
      4907: inst = 32'h10408000;
      4908: inst = 32'hc404b35;
      4909: inst = 32'h8220000;
      4910: inst = 32'h10408000;
      4911: inst = 32'hc404b36;
      4912: inst = 32'h8220000;
      4913: inst = 32'h10408000;
      4914: inst = 32'hc404b37;
      4915: inst = 32'h8220000;
      4916: inst = 32'h10408000;
      4917: inst = 32'hc404b38;
      4918: inst = 32'h8220000;
      4919: inst = 32'h10408000;
      4920: inst = 32'hc404b39;
      4921: inst = 32'h8220000;
      4922: inst = 32'h10408000;
      4923: inst = 32'hc404b3a;
      4924: inst = 32'h8220000;
      4925: inst = 32'h10408000;
      4926: inst = 32'hc404b3b;
      4927: inst = 32'h8220000;
      4928: inst = 32'h10408000;
      4929: inst = 32'hc404b64;
      4930: inst = 32'h8220000;
      4931: inst = 32'h10408000;
      4932: inst = 32'hc404b65;
      4933: inst = 32'h8220000;
      4934: inst = 32'h10408000;
      4935: inst = 32'hc404b66;
      4936: inst = 32'h8220000;
      4937: inst = 32'h10408000;
      4938: inst = 32'hc404b67;
      4939: inst = 32'h8220000;
      4940: inst = 32'h10408000;
      4941: inst = 32'hc404b68;
      4942: inst = 32'h8220000;
      4943: inst = 32'h10408000;
      4944: inst = 32'hc404b69;
      4945: inst = 32'h8220000;
      4946: inst = 32'h10408000;
      4947: inst = 32'hc404b6a;
      4948: inst = 32'h8220000;
      4949: inst = 32'h10408000;
      4950: inst = 32'hc404b6b;
      4951: inst = 32'h8220000;
      4952: inst = 32'h10408000;
      4953: inst = 32'hc404b6c;
      4954: inst = 32'h8220000;
      4955: inst = 32'h10408000;
      4956: inst = 32'hc404b6d;
      4957: inst = 32'h8220000;
      4958: inst = 32'h10408000;
      4959: inst = 32'hc404b6e;
      4960: inst = 32'h8220000;
      4961: inst = 32'h10408000;
      4962: inst = 32'hc404b80;
      4963: inst = 32'h8220000;
      4964: inst = 32'h10408000;
      4965: inst = 32'hc404b81;
      4966: inst = 32'h8220000;
      4967: inst = 32'h10408000;
      4968: inst = 32'hc404b82;
      4969: inst = 32'h8220000;
      4970: inst = 32'h10408000;
      4971: inst = 32'hc404b83;
      4972: inst = 32'h8220000;
      4973: inst = 32'h10408000;
      4974: inst = 32'hc404b84;
      4975: inst = 32'h8220000;
      4976: inst = 32'h10408000;
      4977: inst = 32'hc404b85;
      4978: inst = 32'h8220000;
      4979: inst = 32'h10408000;
      4980: inst = 32'hc404b86;
      4981: inst = 32'h8220000;
      4982: inst = 32'h10408000;
      4983: inst = 32'hc404b90;
      4984: inst = 32'h8220000;
      4985: inst = 32'h10408000;
      4986: inst = 32'hc404b91;
      4987: inst = 32'h8220000;
      4988: inst = 32'h10408000;
      4989: inst = 32'hc404b92;
      4990: inst = 32'h8220000;
      4991: inst = 32'h10408000;
      4992: inst = 32'hc404b93;
      4993: inst = 32'h8220000;
      4994: inst = 32'h10408000;
      4995: inst = 32'hc404b94;
      4996: inst = 32'h8220000;
      4997: inst = 32'h10408000;
      4998: inst = 32'hc404b95;
      4999: inst = 32'h8220000;
      5000: inst = 32'h10408000;
      5001: inst = 32'hc404b96;
      5002: inst = 32'h8220000;
      5003: inst = 32'h10408000;
      5004: inst = 32'hc404b97;
      5005: inst = 32'h8220000;
      5006: inst = 32'h10408000;
      5007: inst = 32'hc404b98;
      5008: inst = 32'h8220000;
      5009: inst = 32'h10408000;
      5010: inst = 32'hc404b99;
      5011: inst = 32'h8220000;
      5012: inst = 32'h10408000;
      5013: inst = 32'hc404b9a;
      5014: inst = 32'h8220000;
      5015: inst = 32'h10408000;
      5016: inst = 32'hc404b9b;
      5017: inst = 32'h8220000;
      5018: inst = 32'h10408000;
      5019: inst = 32'hc404bc4;
      5020: inst = 32'h8220000;
      5021: inst = 32'h10408000;
      5022: inst = 32'hc404bc5;
      5023: inst = 32'h8220000;
      5024: inst = 32'h10408000;
      5025: inst = 32'hc404bc6;
      5026: inst = 32'h8220000;
      5027: inst = 32'h10408000;
      5028: inst = 32'hc404bc7;
      5029: inst = 32'h8220000;
      5030: inst = 32'h10408000;
      5031: inst = 32'hc404bc8;
      5032: inst = 32'h8220000;
      5033: inst = 32'h10408000;
      5034: inst = 32'hc404bc9;
      5035: inst = 32'h8220000;
      5036: inst = 32'h10408000;
      5037: inst = 32'hc404bca;
      5038: inst = 32'h8220000;
      5039: inst = 32'h10408000;
      5040: inst = 32'hc404bcb;
      5041: inst = 32'h8220000;
      5042: inst = 32'h10408000;
      5043: inst = 32'hc404bcc;
      5044: inst = 32'h8220000;
      5045: inst = 32'h10408000;
      5046: inst = 32'hc404bcd;
      5047: inst = 32'h8220000;
      5048: inst = 32'h10408000;
      5049: inst = 32'hc404bce;
      5050: inst = 32'h8220000;
      5051: inst = 32'h10408000;
      5052: inst = 32'hc404be0;
      5053: inst = 32'h8220000;
      5054: inst = 32'h10408000;
      5055: inst = 32'hc404be1;
      5056: inst = 32'h8220000;
      5057: inst = 32'h10408000;
      5058: inst = 32'hc404be2;
      5059: inst = 32'h8220000;
      5060: inst = 32'h10408000;
      5061: inst = 32'hc404be3;
      5062: inst = 32'h8220000;
      5063: inst = 32'h10408000;
      5064: inst = 32'hc404be4;
      5065: inst = 32'h8220000;
      5066: inst = 32'h10408000;
      5067: inst = 32'hc404be5;
      5068: inst = 32'h8220000;
      5069: inst = 32'h10408000;
      5070: inst = 32'hc404be6;
      5071: inst = 32'h8220000;
      5072: inst = 32'h10408000;
      5073: inst = 32'hc404bf0;
      5074: inst = 32'h8220000;
      5075: inst = 32'h10408000;
      5076: inst = 32'hc404bf1;
      5077: inst = 32'h8220000;
      5078: inst = 32'h10408000;
      5079: inst = 32'hc404bf2;
      5080: inst = 32'h8220000;
      5081: inst = 32'h10408000;
      5082: inst = 32'hc404bf3;
      5083: inst = 32'h8220000;
      5084: inst = 32'h10408000;
      5085: inst = 32'hc404bf4;
      5086: inst = 32'h8220000;
      5087: inst = 32'h10408000;
      5088: inst = 32'hc404bf5;
      5089: inst = 32'h8220000;
      5090: inst = 32'h10408000;
      5091: inst = 32'hc404bf6;
      5092: inst = 32'h8220000;
      5093: inst = 32'h10408000;
      5094: inst = 32'hc404bf7;
      5095: inst = 32'h8220000;
      5096: inst = 32'h10408000;
      5097: inst = 32'hc404bf8;
      5098: inst = 32'h8220000;
      5099: inst = 32'h10408000;
      5100: inst = 32'hc404bf9;
      5101: inst = 32'h8220000;
      5102: inst = 32'h10408000;
      5103: inst = 32'hc404c26;
      5104: inst = 32'h8220000;
      5105: inst = 32'h10408000;
      5106: inst = 32'hc404c27;
      5107: inst = 32'h8220000;
      5108: inst = 32'h10408000;
      5109: inst = 32'hc404c28;
      5110: inst = 32'h8220000;
      5111: inst = 32'h10408000;
      5112: inst = 32'hc404c29;
      5113: inst = 32'h8220000;
      5114: inst = 32'h10408000;
      5115: inst = 32'hc404c2a;
      5116: inst = 32'h8220000;
      5117: inst = 32'h10408000;
      5118: inst = 32'hc404c2b;
      5119: inst = 32'h8220000;
      5120: inst = 32'h10408000;
      5121: inst = 32'hc404c2c;
      5122: inst = 32'h8220000;
      5123: inst = 32'h10408000;
      5124: inst = 32'hc404c2d;
      5125: inst = 32'h8220000;
      5126: inst = 32'h10408000;
      5127: inst = 32'hc404c2e;
      5128: inst = 32'h8220000;
      5129: inst = 32'h10408000;
      5130: inst = 32'hc404c40;
      5131: inst = 32'h8220000;
      5132: inst = 32'h10408000;
      5133: inst = 32'hc404c41;
      5134: inst = 32'h8220000;
      5135: inst = 32'h10408000;
      5136: inst = 32'hc404c42;
      5137: inst = 32'h8220000;
      5138: inst = 32'h10408000;
      5139: inst = 32'hc404c43;
      5140: inst = 32'h8220000;
      5141: inst = 32'h10408000;
      5142: inst = 32'hc404c44;
      5143: inst = 32'h8220000;
      5144: inst = 32'h10408000;
      5145: inst = 32'hc404c45;
      5146: inst = 32'h8220000;
      5147: inst = 32'h10408000;
      5148: inst = 32'hc404c46;
      5149: inst = 32'h8220000;
      5150: inst = 32'h10408000;
      5151: inst = 32'hc404c4f;
      5152: inst = 32'h8220000;
      5153: inst = 32'h10408000;
      5154: inst = 32'hc404c50;
      5155: inst = 32'h8220000;
      5156: inst = 32'h10408000;
      5157: inst = 32'hc404c51;
      5158: inst = 32'h8220000;
      5159: inst = 32'h10408000;
      5160: inst = 32'hc404c52;
      5161: inst = 32'h8220000;
      5162: inst = 32'h10408000;
      5163: inst = 32'hc404c53;
      5164: inst = 32'h8220000;
      5165: inst = 32'h10408000;
      5166: inst = 32'hc404c54;
      5167: inst = 32'h8220000;
      5168: inst = 32'h10408000;
      5169: inst = 32'hc404c55;
      5170: inst = 32'h8220000;
      5171: inst = 32'h10408000;
      5172: inst = 32'hc404c56;
      5173: inst = 32'h8220000;
      5174: inst = 32'h10408000;
      5175: inst = 32'hc404c57;
      5176: inst = 32'h8220000;
      5177: inst = 32'h10408000;
      5178: inst = 32'hc404c58;
      5179: inst = 32'h8220000;
      5180: inst = 32'h10408000;
      5181: inst = 32'hc404c59;
      5182: inst = 32'h8220000;
      5183: inst = 32'h10408000;
      5184: inst = 32'hc404c5a;
      5185: inst = 32'h8220000;
      5186: inst = 32'h10408000;
      5187: inst = 32'hc404c5b;
      5188: inst = 32'h8220000;
      5189: inst = 32'h10408000;
      5190: inst = 32'hc404c5c;
      5191: inst = 32'h8220000;
      5192: inst = 32'h10408000;
      5193: inst = 32'hc404c5d;
      5194: inst = 32'h8220000;
      5195: inst = 32'h10408000;
      5196: inst = 32'hc404c5e;
      5197: inst = 32'h8220000;
      5198: inst = 32'h10408000;
      5199: inst = 32'hc404c5f;
      5200: inst = 32'h8220000;
      5201: inst = 32'h10408000;
      5202: inst = 32'hc404c60;
      5203: inst = 32'h8220000;
      5204: inst = 32'h10408000;
      5205: inst = 32'hc404c61;
      5206: inst = 32'h8220000;
      5207: inst = 32'h10408000;
      5208: inst = 32'hc404c62;
      5209: inst = 32'h8220000;
      5210: inst = 32'h10408000;
      5211: inst = 32'hc404c63;
      5212: inst = 32'h8220000;
      5213: inst = 32'h10408000;
      5214: inst = 32'hc404c64;
      5215: inst = 32'h8220000;
      5216: inst = 32'h10408000;
      5217: inst = 32'hc404c65;
      5218: inst = 32'h8220000;
      5219: inst = 32'h10408000;
      5220: inst = 32'hc404c66;
      5221: inst = 32'h8220000;
      5222: inst = 32'h10408000;
      5223: inst = 32'hc404c67;
      5224: inst = 32'h8220000;
      5225: inst = 32'h10408000;
      5226: inst = 32'hc404c68;
      5227: inst = 32'h8220000;
      5228: inst = 32'h10408000;
      5229: inst = 32'hc404c69;
      5230: inst = 32'h8220000;
      5231: inst = 32'h10408000;
      5232: inst = 32'hc404c6a;
      5233: inst = 32'h8220000;
      5234: inst = 32'h10408000;
      5235: inst = 32'hc404c6b;
      5236: inst = 32'h8220000;
      5237: inst = 32'h10408000;
      5238: inst = 32'hc404c6c;
      5239: inst = 32'h8220000;
      5240: inst = 32'h10408000;
      5241: inst = 32'hc404c6d;
      5242: inst = 32'h8220000;
      5243: inst = 32'h10408000;
      5244: inst = 32'hc404c6e;
      5245: inst = 32'h8220000;
      5246: inst = 32'h10408000;
      5247: inst = 32'hc404c6f;
      5248: inst = 32'h8220000;
      5249: inst = 32'h10408000;
      5250: inst = 32'hc404c70;
      5251: inst = 32'h8220000;
      5252: inst = 32'h10408000;
      5253: inst = 32'hc404c71;
      5254: inst = 32'h8220000;
      5255: inst = 32'h10408000;
      5256: inst = 32'hc404c72;
      5257: inst = 32'h8220000;
      5258: inst = 32'h10408000;
      5259: inst = 32'hc404c73;
      5260: inst = 32'h8220000;
      5261: inst = 32'h10408000;
      5262: inst = 32'hc404c74;
      5263: inst = 32'h8220000;
      5264: inst = 32'h10408000;
      5265: inst = 32'hc404c75;
      5266: inst = 32'h8220000;
      5267: inst = 32'h10408000;
      5268: inst = 32'hc404c76;
      5269: inst = 32'h8220000;
      5270: inst = 32'h10408000;
      5271: inst = 32'hc404c77;
      5272: inst = 32'h8220000;
      5273: inst = 32'h10408000;
      5274: inst = 32'hc404c78;
      5275: inst = 32'h8220000;
      5276: inst = 32'h10408000;
      5277: inst = 32'hc404c79;
      5278: inst = 32'h8220000;
      5279: inst = 32'h10408000;
      5280: inst = 32'hc404c7a;
      5281: inst = 32'h8220000;
      5282: inst = 32'h10408000;
      5283: inst = 32'hc404c7b;
      5284: inst = 32'h8220000;
      5285: inst = 32'h10408000;
      5286: inst = 32'hc404c7c;
      5287: inst = 32'h8220000;
      5288: inst = 32'h10408000;
      5289: inst = 32'hc404c7d;
      5290: inst = 32'h8220000;
      5291: inst = 32'h10408000;
      5292: inst = 32'hc404c7e;
      5293: inst = 32'h8220000;
      5294: inst = 32'h10408000;
      5295: inst = 32'hc404c7f;
      5296: inst = 32'h8220000;
      5297: inst = 32'h10408000;
      5298: inst = 32'hc404c80;
      5299: inst = 32'h8220000;
      5300: inst = 32'h10408000;
      5301: inst = 32'hc404c81;
      5302: inst = 32'h8220000;
      5303: inst = 32'h10408000;
      5304: inst = 32'hc404c82;
      5305: inst = 32'h8220000;
      5306: inst = 32'h10408000;
      5307: inst = 32'hc404c83;
      5308: inst = 32'h8220000;
      5309: inst = 32'h10408000;
      5310: inst = 32'hc404c84;
      5311: inst = 32'h8220000;
      5312: inst = 32'h10408000;
      5313: inst = 32'hc404c85;
      5314: inst = 32'h8220000;
      5315: inst = 32'h10408000;
      5316: inst = 32'hc404c86;
      5317: inst = 32'h8220000;
      5318: inst = 32'h10408000;
      5319: inst = 32'hc404c87;
      5320: inst = 32'h8220000;
      5321: inst = 32'h10408000;
      5322: inst = 32'hc404c88;
      5323: inst = 32'h8220000;
      5324: inst = 32'h10408000;
      5325: inst = 32'hc404c89;
      5326: inst = 32'h8220000;
      5327: inst = 32'h10408000;
      5328: inst = 32'hc404c8a;
      5329: inst = 32'h8220000;
      5330: inst = 32'h10408000;
      5331: inst = 32'hc404c8b;
      5332: inst = 32'h8220000;
      5333: inst = 32'h10408000;
      5334: inst = 32'hc404c8c;
      5335: inst = 32'h8220000;
      5336: inst = 32'h10408000;
      5337: inst = 32'hc404c8d;
      5338: inst = 32'h8220000;
      5339: inst = 32'h10408000;
      5340: inst = 32'hc404c8e;
      5341: inst = 32'h8220000;
      5342: inst = 32'h10408000;
      5343: inst = 32'hc404ca0;
      5344: inst = 32'h8220000;
      5345: inst = 32'h10408000;
      5346: inst = 32'hc404ca1;
      5347: inst = 32'h8220000;
      5348: inst = 32'h10408000;
      5349: inst = 32'hc404cb7;
      5350: inst = 32'h8220000;
      5351: inst = 32'h10408000;
      5352: inst = 32'hc404cb8;
      5353: inst = 32'h8220000;
      5354: inst = 32'h10408000;
      5355: inst = 32'hc404cb9;
      5356: inst = 32'h8220000;
      5357: inst = 32'h10408000;
      5358: inst = 32'hc404cba;
      5359: inst = 32'h8220000;
      5360: inst = 32'h10408000;
      5361: inst = 32'hc404cbb;
      5362: inst = 32'h8220000;
      5363: inst = 32'h10408000;
      5364: inst = 32'hc404cbc;
      5365: inst = 32'h8220000;
      5366: inst = 32'h10408000;
      5367: inst = 32'hc404cbd;
      5368: inst = 32'h8220000;
      5369: inst = 32'h10408000;
      5370: inst = 32'hc404cbe;
      5371: inst = 32'h8220000;
      5372: inst = 32'h10408000;
      5373: inst = 32'hc404cbf;
      5374: inst = 32'h8220000;
      5375: inst = 32'h10408000;
      5376: inst = 32'hc404cc0;
      5377: inst = 32'h8220000;
      5378: inst = 32'h10408000;
      5379: inst = 32'hc404cc1;
      5380: inst = 32'h8220000;
      5381: inst = 32'h10408000;
      5382: inst = 32'hc404cc2;
      5383: inst = 32'h8220000;
      5384: inst = 32'h10408000;
      5385: inst = 32'hc404cc3;
      5386: inst = 32'h8220000;
      5387: inst = 32'h10408000;
      5388: inst = 32'hc404cc4;
      5389: inst = 32'h8220000;
      5390: inst = 32'h10408000;
      5391: inst = 32'hc404cc5;
      5392: inst = 32'h8220000;
      5393: inst = 32'h10408000;
      5394: inst = 32'hc404cc6;
      5395: inst = 32'h8220000;
      5396: inst = 32'h10408000;
      5397: inst = 32'hc404cc7;
      5398: inst = 32'h8220000;
      5399: inst = 32'h10408000;
      5400: inst = 32'hc404cc8;
      5401: inst = 32'h8220000;
      5402: inst = 32'h10408000;
      5403: inst = 32'hc404cc9;
      5404: inst = 32'h8220000;
      5405: inst = 32'h10408000;
      5406: inst = 32'hc404cca;
      5407: inst = 32'h8220000;
      5408: inst = 32'h10408000;
      5409: inst = 32'hc404ccb;
      5410: inst = 32'h8220000;
      5411: inst = 32'h10408000;
      5412: inst = 32'hc404ccc;
      5413: inst = 32'h8220000;
      5414: inst = 32'h10408000;
      5415: inst = 32'hc404ccd;
      5416: inst = 32'h8220000;
      5417: inst = 32'h10408000;
      5418: inst = 32'hc404cce;
      5419: inst = 32'h8220000;
      5420: inst = 32'h10408000;
      5421: inst = 32'hc404ccf;
      5422: inst = 32'h8220000;
      5423: inst = 32'h10408000;
      5424: inst = 32'hc404cd0;
      5425: inst = 32'h8220000;
      5426: inst = 32'h10408000;
      5427: inst = 32'hc404cd1;
      5428: inst = 32'h8220000;
      5429: inst = 32'h10408000;
      5430: inst = 32'hc404cd2;
      5431: inst = 32'h8220000;
      5432: inst = 32'h10408000;
      5433: inst = 32'hc404cd3;
      5434: inst = 32'h8220000;
      5435: inst = 32'h10408000;
      5436: inst = 32'hc404cd4;
      5437: inst = 32'h8220000;
      5438: inst = 32'h10408000;
      5439: inst = 32'hc404cd5;
      5440: inst = 32'h8220000;
      5441: inst = 32'h10408000;
      5442: inst = 32'hc404cd6;
      5443: inst = 32'h8220000;
      5444: inst = 32'h10408000;
      5445: inst = 32'hc404cd7;
      5446: inst = 32'h8220000;
      5447: inst = 32'h10408000;
      5448: inst = 32'hc404cd8;
      5449: inst = 32'h8220000;
      5450: inst = 32'h10408000;
      5451: inst = 32'hc404cd9;
      5452: inst = 32'h8220000;
      5453: inst = 32'h10408000;
      5454: inst = 32'hc404cda;
      5455: inst = 32'h8220000;
      5456: inst = 32'h10408000;
      5457: inst = 32'hc404cdb;
      5458: inst = 32'h8220000;
      5459: inst = 32'h10408000;
      5460: inst = 32'hc404cdc;
      5461: inst = 32'h8220000;
      5462: inst = 32'h10408000;
      5463: inst = 32'hc404cdd;
      5464: inst = 32'h8220000;
      5465: inst = 32'h10408000;
      5466: inst = 32'hc404cde;
      5467: inst = 32'h8220000;
      5468: inst = 32'h10408000;
      5469: inst = 32'hc404cdf;
      5470: inst = 32'h8220000;
      5471: inst = 32'h10408000;
      5472: inst = 32'hc404ce0;
      5473: inst = 32'h8220000;
      5474: inst = 32'h10408000;
      5475: inst = 32'hc404ce1;
      5476: inst = 32'h8220000;
      5477: inst = 32'h10408000;
      5478: inst = 32'hc404ce2;
      5479: inst = 32'h8220000;
      5480: inst = 32'h10408000;
      5481: inst = 32'hc404ce3;
      5482: inst = 32'h8220000;
      5483: inst = 32'h10408000;
      5484: inst = 32'hc404ce4;
      5485: inst = 32'h8220000;
      5486: inst = 32'h10408000;
      5487: inst = 32'hc404ce5;
      5488: inst = 32'h8220000;
      5489: inst = 32'h10408000;
      5490: inst = 32'hc404ce6;
      5491: inst = 32'h8220000;
      5492: inst = 32'h10408000;
      5493: inst = 32'hc404ce7;
      5494: inst = 32'h8220000;
      5495: inst = 32'h10408000;
      5496: inst = 32'hc404ce8;
      5497: inst = 32'h8220000;
      5498: inst = 32'h10408000;
      5499: inst = 32'hc404ce9;
      5500: inst = 32'h8220000;
      5501: inst = 32'h10408000;
      5502: inst = 32'hc404cea;
      5503: inst = 32'h8220000;
      5504: inst = 32'h10408000;
      5505: inst = 32'hc404ceb;
      5506: inst = 32'h8220000;
      5507: inst = 32'h10408000;
      5508: inst = 32'hc404cec;
      5509: inst = 32'h8220000;
      5510: inst = 32'h10408000;
      5511: inst = 32'hc404ced;
      5512: inst = 32'h8220000;
      5513: inst = 32'h10408000;
      5514: inst = 32'hc404cee;
      5515: inst = 32'h8220000;
      5516: inst = 32'h10408000;
      5517: inst = 32'hc404d17;
      5518: inst = 32'h8220000;
      5519: inst = 32'h10408000;
      5520: inst = 32'hc404d18;
      5521: inst = 32'h8220000;
      5522: inst = 32'h10408000;
      5523: inst = 32'hc404d19;
      5524: inst = 32'h8220000;
      5525: inst = 32'h10408000;
      5526: inst = 32'hc404d1a;
      5527: inst = 32'h8220000;
      5528: inst = 32'h10408000;
      5529: inst = 32'hc404d1b;
      5530: inst = 32'h8220000;
      5531: inst = 32'h10408000;
      5532: inst = 32'hc404d1c;
      5533: inst = 32'h8220000;
      5534: inst = 32'h10408000;
      5535: inst = 32'hc404d1d;
      5536: inst = 32'h8220000;
      5537: inst = 32'h10408000;
      5538: inst = 32'hc404d1e;
      5539: inst = 32'h8220000;
      5540: inst = 32'h10408000;
      5541: inst = 32'hc404d1f;
      5542: inst = 32'h8220000;
      5543: inst = 32'h10408000;
      5544: inst = 32'hc404d20;
      5545: inst = 32'h8220000;
      5546: inst = 32'h10408000;
      5547: inst = 32'hc404d21;
      5548: inst = 32'h8220000;
      5549: inst = 32'h10408000;
      5550: inst = 32'hc404d22;
      5551: inst = 32'h8220000;
      5552: inst = 32'h10408000;
      5553: inst = 32'hc404d23;
      5554: inst = 32'h8220000;
      5555: inst = 32'h10408000;
      5556: inst = 32'hc404d24;
      5557: inst = 32'h8220000;
      5558: inst = 32'h10408000;
      5559: inst = 32'hc404d25;
      5560: inst = 32'h8220000;
      5561: inst = 32'h10408000;
      5562: inst = 32'hc404d26;
      5563: inst = 32'h8220000;
      5564: inst = 32'h10408000;
      5565: inst = 32'hc404d27;
      5566: inst = 32'h8220000;
      5567: inst = 32'h10408000;
      5568: inst = 32'hc404d28;
      5569: inst = 32'h8220000;
      5570: inst = 32'h10408000;
      5571: inst = 32'hc404d29;
      5572: inst = 32'h8220000;
      5573: inst = 32'h10408000;
      5574: inst = 32'hc404d2a;
      5575: inst = 32'h8220000;
      5576: inst = 32'h10408000;
      5577: inst = 32'hc404d2b;
      5578: inst = 32'h8220000;
      5579: inst = 32'h10408000;
      5580: inst = 32'hc404d2c;
      5581: inst = 32'h8220000;
      5582: inst = 32'h10408000;
      5583: inst = 32'hc404d2d;
      5584: inst = 32'h8220000;
      5585: inst = 32'h10408000;
      5586: inst = 32'hc404d2e;
      5587: inst = 32'h8220000;
      5588: inst = 32'h10408000;
      5589: inst = 32'hc404d2f;
      5590: inst = 32'h8220000;
      5591: inst = 32'h10408000;
      5592: inst = 32'hc404d30;
      5593: inst = 32'h8220000;
      5594: inst = 32'h10408000;
      5595: inst = 32'hc404d31;
      5596: inst = 32'h8220000;
      5597: inst = 32'h10408000;
      5598: inst = 32'hc404d32;
      5599: inst = 32'h8220000;
      5600: inst = 32'h10408000;
      5601: inst = 32'hc404d33;
      5602: inst = 32'h8220000;
      5603: inst = 32'h10408000;
      5604: inst = 32'hc404d34;
      5605: inst = 32'h8220000;
      5606: inst = 32'h10408000;
      5607: inst = 32'hc404d35;
      5608: inst = 32'h8220000;
      5609: inst = 32'h10408000;
      5610: inst = 32'hc404d36;
      5611: inst = 32'h8220000;
      5612: inst = 32'h10408000;
      5613: inst = 32'hc404d37;
      5614: inst = 32'h8220000;
      5615: inst = 32'h10408000;
      5616: inst = 32'hc404d38;
      5617: inst = 32'h8220000;
      5618: inst = 32'h10408000;
      5619: inst = 32'hc404d39;
      5620: inst = 32'h8220000;
      5621: inst = 32'h10408000;
      5622: inst = 32'hc404d3a;
      5623: inst = 32'h8220000;
      5624: inst = 32'h10408000;
      5625: inst = 32'hc404d3b;
      5626: inst = 32'h8220000;
      5627: inst = 32'h10408000;
      5628: inst = 32'hc404d3c;
      5629: inst = 32'h8220000;
      5630: inst = 32'h10408000;
      5631: inst = 32'hc404d3d;
      5632: inst = 32'h8220000;
      5633: inst = 32'h10408000;
      5634: inst = 32'hc404d3e;
      5635: inst = 32'h8220000;
      5636: inst = 32'h10408000;
      5637: inst = 32'hc404d3f;
      5638: inst = 32'h8220000;
      5639: inst = 32'h10408000;
      5640: inst = 32'hc404d40;
      5641: inst = 32'h8220000;
      5642: inst = 32'h10408000;
      5643: inst = 32'hc404d41;
      5644: inst = 32'h8220000;
      5645: inst = 32'h10408000;
      5646: inst = 32'hc404d42;
      5647: inst = 32'h8220000;
      5648: inst = 32'h10408000;
      5649: inst = 32'hc404d43;
      5650: inst = 32'h8220000;
      5651: inst = 32'h10408000;
      5652: inst = 32'hc404d44;
      5653: inst = 32'h8220000;
      5654: inst = 32'h10408000;
      5655: inst = 32'hc404d45;
      5656: inst = 32'h8220000;
      5657: inst = 32'h10408000;
      5658: inst = 32'hc404d46;
      5659: inst = 32'h8220000;
      5660: inst = 32'h10408000;
      5661: inst = 32'hc404d47;
      5662: inst = 32'h8220000;
      5663: inst = 32'h10408000;
      5664: inst = 32'hc404d48;
      5665: inst = 32'h8220000;
      5666: inst = 32'h10408000;
      5667: inst = 32'hc404d49;
      5668: inst = 32'h8220000;
      5669: inst = 32'h10408000;
      5670: inst = 32'hc404d4a;
      5671: inst = 32'h8220000;
      5672: inst = 32'h10408000;
      5673: inst = 32'hc404d4b;
      5674: inst = 32'h8220000;
      5675: inst = 32'h10408000;
      5676: inst = 32'hc404d4c;
      5677: inst = 32'h8220000;
      5678: inst = 32'h10408000;
      5679: inst = 32'hc404d4d;
      5680: inst = 32'h8220000;
      5681: inst = 32'h10408000;
      5682: inst = 32'hc404d4e;
      5683: inst = 32'h8220000;
      5684: inst = 32'h10408000;
      5685: inst = 32'hc404d77;
      5686: inst = 32'h8220000;
      5687: inst = 32'h10408000;
      5688: inst = 32'hc404d78;
      5689: inst = 32'h8220000;
      5690: inst = 32'h10408000;
      5691: inst = 32'hc404d79;
      5692: inst = 32'h8220000;
      5693: inst = 32'h10408000;
      5694: inst = 32'hc404d7a;
      5695: inst = 32'h8220000;
      5696: inst = 32'h10408000;
      5697: inst = 32'hc404d7b;
      5698: inst = 32'h8220000;
      5699: inst = 32'h10408000;
      5700: inst = 32'hc404d7c;
      5701: inst = 32'h8220000;
      5702: inst = 32'h10408000;
      5703: inst = 32'hc404d7d;
      5704: inst = 32'h8220000;
      5705: inst = 32'h10408000;
      5706: inst = 32'hc404d7e;
      5707: inst = 32'h8220000;
      5708: inst = 32'h10408000;
      5709: inst = 32'hc404d7f;
      5710: inst = 32'h8220000;
      5711: inst = 32'h10408000;
      5712: inst = 32'hc404d80;
      5713: inst = 32'h8220000;
      5714: inst = 32'h10408000;
      5715: inst = 32'hc404d81;
      5716: inst = 32'h8220000;
      5717: inst = 32'h10408000;
      5718: inst = 32'hc404d82;
      5719: inst = 32'h8220000;
      5720: inst = 32'h10408000;
      5721: inst = 32'hc404d83;
      5722: inst = 32'h8220000;
      5723: inst = 32'h10408000;
      5724: inst = 32'hc404d84;
      5725: inst = 32'h8220000;
      5726: inst = 32'h10408000;
      5727: inst = 32'hc404d85;
      5728: inst = 32'h8220000;
      5729: inst = 32'h10408000;
      5730: inst = 32'hc404d86;
      5731: inst = 32'h8220000;
      5732: inst = 32'h10408000;
      5733: inst = 32'hc404d87;
      5734: inst = 32'h8220000;
      5735: inst = 32'h10408000;
      5736: inst = 32'hc404d88;
      5737: inst = 32'h8220000;
      5738: inst = 32'h10408000;
      5739: inst = 32'hc404d89;
      5740: inst = 32'h8220000;
      5741: inst = 32'h10408000;
      5742: inst = 32'hc404d8a;
      5743: inst = 32'h8220000;
      5744: inst = 32'h10408000;
      5745: inst = 32'hc404d8b;
      5746: inst = 32'h8220000;
      5747: inst = 32'h10408000;
      5748: inst = 32'hc404d8c;
      5749: inst = 32'h8220000;
      5750: inst = 32'h10408000;
      5751: inst = 32'hc404d8d;
      5752: inst = 32'h8220000;
      5753: inst = 32'h10408000;
      5754: inst = 32'hc404d8e;
      5755: inst = 32'h8220000;
      5756: inst = 32'h10408000;
      5757: inst = 32'hc404d8f;
      5758: inst = 32'h8220000;
      5759: inst = 32'h10408000;
      5760: inst = 32'hc404d90;
      5761: inst = 32'h8220000;
      5762: inst = 32'h10408000;
      5763: inst = 32'hc404d91;
      5764: inst = 32'h8220000;
      5765: inst = 32'h10408000;
      5766: inst = 32'hc404d92;
      5767: inst = 32'h8220000;
      5768: inst = 32'h10408000;
      5769: inst = 32'hc404d93;
      5770: inst = 32'h8220000;
      5771: inst = 32'h10408000;
      5772: inst = 32'hc404d94;
      5773: inst = 32'h8220000;
      5774: inst = 32'h10408000;
      5775: inst = 32'hc404d95;
      5776: inst = 32'h8220000;
      5777: inst = 32'h10408000;
      5778: inst = 32'hc404d96;
      5779: inst = 32'h8220000;
      5780: inst = 32'h10408000;
      5781: inst = 32'hc404d97;
      5782: inst = 32'h8220000;
      5783: inst = 32'h10408000;
      5784: inst = 32'hc404d98;
      5785: inst = 32'h8220000;
      5786: inst = 32'h10408000;
      5787: inst = 32'hc404d99;
      5788: inst = 32'h8220000;
      5789: inst = 32'h10408000;
      5790: inst = 32'hc404d9a;
      5791: inst = 32'h8220000;
      5792: inst = 32'h10408000;
      5793: inst = 32'hc404d9b;
      5794: inst = 32'h8220000;
      5795: inst = 32'h10408000;
      5796: inst = 32'hc404d9c;
      5797: inst = 32'h8220000;
      5798: inst = 32'h10408000;
      5799: inst = 32'hc404d9d;
      5800: inst = 32'h8220000;
      5801: inst = 32'h10408000;
      5802: inst = 32'hc404d9e;
      5803: inst = 32'h8220000;
      5804: inst = 32'h10408000;
      5805: inst = 32'hc404d9f;
      5806: inst = 32'h8220000;
      5807: inst = 32'h10408000;
      5808: inst = 32'hc404da0;
      5809: inst = 32'h8220000;
      5810: inst = 32'h10408000;
      5811: inst = 32'hc404da1;
      5812: inst = 32'h8220000;
      5813: inst = 32'h10408000;
      5814: inst = 32'hc404da2;
      5815: inst = 32'h8220000;
      5816: inst = 32'h10408000;
      5817: inst = 32'hc404da3;
      5818: inst = 32'h8220000;
      5819: inst = 32'h10408000;
      5820: inst = 32'hc404da4;
      5821: inst = 32'h8220000;
      5822: inst = 32'h10408000;
      5823: inst = 32'hc404da5;
      5824: inst = 32'h8220000;
      5825: inst = 32'h10408000;
      5826: inst = 32'hc404da6;
      5827: inst = 32'h8220000;
      5828: inst = 32'h10408000;
      5829: inst = 32'hc404da7;
      5830: inst = 32'h8220000;
      5831: inst = 32'h10408000;
      5832: inst = 32'hc404da8;
      5833: inst = 32'h8220000;
      5834: inst = 32'h10408000;
      5835: inst = 32'hc404da9;
      5836: inst = 32'h8220000;
      5837: inst = 32'h10408000;
      5838: inst = 32'hc404daa;
      5839: inst = 32'h8220000;
      5840: inst = 32'h10408000;
      5841: inst = 32'hc404dab;
      5842: inst = 32'h8220000;
      5843: inst = 32'h10408000;
      5844: inst = 32'hc404dac;
      5845: inst = 32'h8220000;
      5846: inst = 32'h10408000;
      5847: inst = 32'hc404dad;
      5848: inst = 32'h8220000;
      5849: inst = 32'h10408000;
      5850: inst = 32'hc404dae;
      5851: inst = 32'h8220000;
      5852: inst = 32'h10408000;
      5853: inst = 32'hc404dd7;
      5854: inst = 32'h8220000;
      5855: inst = 32'h10408000;
      5856: inst = 32'hc404dd8;
      5857: inst = 32'h8220000;
      5858: inst = 32'h10408000;
      5859: inst = 32'hc404dd9;
      5860: inst = 32'h8220000;
      5861: inst = 32'h10408000;
      5862: inst = 32'hc404dda;
      5863: inst = 32'h8220000;
      5864: inst = 32'h10408000;
      5865: inst = 32'hc404ddb;
      5866: inst = 32'h8220000;
      5867: inst = 32'h10408000;
      5868: inst = 32'hc404ddc;
      5869: inst = 32'h8220000;
      5870: inst = 32'h10408000;
      5871: inst = 32'hc404ddd;
      5872: inst = 32'h8220000;
      5873: inst = 32'h10408000;
      5874: inst = 32'hc404dde;
      5875: inst = 32'h8220000;
      5876: inst = 32'h10408000;
      5877: inst = 32'hc404ddf;
      5878: inst = 32'h8220000;
      5879: inst = 32'h10408000;
      5880: inst = 32'hc404de0;
      5881: inst = 32'h8220000;
      5882: inst = 32'h10408000;
      5883: inst = 32'hc404de1;
      5884: inst = 32'h8220000;
      5885: inst = 32'h10408000;
      5886: inst = 32'hc404de2;
      5887: inst = 32'h8220000;
      5888: inst = 32'h10408000;
      5889: inst = 32'hc404de3;
      5890: inst = 32'h8220000;
      5891: inst = 32'h10408000;
      5892: inst = 32'hc404de4;
      5893: inst = 32'h8220000;
      5894: inst = 32'h10408000;
      5895: inst = 32'hc404de5;
      5896: inst = 32'h8220000;
      5897: inst = 32'h10408000;
      5898: inst = 32'hc404de6;
      5899: inst = 32'h8220000;
      5900: inst = 32'h10408000;
      5901: inst = 32'hc404de7;
      5902: inst = 32'h8220000;
      5903: inst = 32'h10408000;
      5904: inst = 32'hc404de8;
      5905: inst = 32'h8220000;
      5906: inst = 32'h10408000;
      5907: inst = 32'hc404de9;
      5908: inst = 32'h8220000;
      5909: inst = 32'h10408000;
      5910: inst = 32'hc404dea;
      5911: inst = 32'h8220000;
      5912: inst = 32'h10408000;
      5913: inst = 32'hc404deb;
      5914: inst = 32'h8220000;
      5915: inst = 32'h10408000;
      5916: inst = 32'hc404dec;
      5917: inst = 32'h8220000;
      5918: inst = 32'h10408000;
      5919: inst = 32'hc404ded;
      5920: inst = 32'h8220000;
      5921: inst = 32'h10408000;
      5922: inst = 32'hc404dee;
      5923: inst = 32'h8220000;
      5924: inst = 32'h10408000;
      5925: inst = 32'hc404def;
      5926: inst = 32'h8220000;
      5927: inst = 32'h10408000;
      5928: inst = 32'hc404df0;
      5929: inst = 32'h8220000;
      5930: inst = 32'h10408000;
      5931: inst = 32'hc404df1;
      5932: inst = 32'h8220000;
      5933: inst = 32'h10408000;
      5934: inst = 32'hc404df2;
      5935: inst = 32'h8220000;
      5936: inst = 32'h10408000;
      5937: inst = 32'hc404df3;
      5938: inst = 32'h8220000;
      5939: inst = 32'h10408000;
      5940: inst = 32'hc404df4;
      5941: inst = 32'h8220000;
      5942: inst = 32'h10408000;
      5943: inst = 32'hc404df5;
      5944: inst = 32'h8220000;
      5945: inst = 32'h10408000;
      5946: inst = 32'hc404df6;
      5947: inst = 32'h8220000;
      5948: inst = 32'h10408000;
      5949: inst = 32'hc404df7;
      5950: inst = 32'h8220000;
      5951: inst = 32'h10408000;
      5952: inst = 32'hc404df8;
      5953: inst = 32'h8220000;
      5954: inst = 32'h10408000;
      5955: inst = 32'hc404df9;
      5956: inst = 32'h8220000;
      5957: inst = 32'h10408000;
      5958: inst = 32'hc404dfa;
      5959: inst = 32'h8220000;
      5960: inst = 32'h10408000;
      5961: inst = 32'hc404dfb;
      5962: inst = 32'h8220000;
      5963: inst = 32'h10408000;
      5964: inst = 32'hc404dfc;
      5965: inst = 32'h8220000;
      5966: inst = 32'h10408000;
      5967: inst = 32'hc404dfd;
      5968: inst = 32'h8220000;
      5969: inst = 32'h10408000;
      5970: inst = 32'hc404dfe;
      5971: inst = 32'h8220000;
      5972: inst = 32'h10408000;
      5973: inst = 32'hc404dff;
      5974: inst = 32'h8220000;
      5975: inst = 32'h10408000;
      5976: inst = 32'hc404e00;
      5977: inst = 32'h8220000;
      5978: inst = 32'h10408000;
      5979: inst = 32'hc404e01;
      5980: inst = 32'h8220000;
      5981: inst = 32'h10408000;
      5982: inst = 32'hc404e02;
      5983: inst = 32'h8220000;
      5984: inst = 32'h10408000;
      5985: inst = 32'hc404e03;
      5986: inst = 32'h8220000;
      5987: inst = 32'h10408000;
      5988: inst = 32'hc404e04;
      5989: inst = 32'h8220000;
      5990: inst = 32'h10408000;
      5991: inst = 32'hc404e05;
      5992: inst = 32'h8220000;
      5993: inst = 32'h10408000;
      5994: inst = 32'hc404e06;
      5995: inst = 32'h8220000;
      5996: inst = 32'h10408000;
      5997: inst = 32'hc404e07;
      5998: inst = 32'h8220000;
      5999: inst = 32'h10408000;
      6000: inst = 32'hc404e08;
      6001: inst = 32'h8220000;
      6002: inst = 32'h10408000;
      6003: inst = 32'hc404e09;
      6004: inst = 32'h8220000;
      6005: inst = 32'h10408000;
      6006: inst = 32'hc404e0a;
      6007: inst = 32'h8220000;
      6008: inst = 32'h10408000;
      6009: inst = 32'hc404e0b;
      6010: inst = 32'h8220000;
      6011: inst = 32'h10408000;
      6012: inst = 32'hc404e0c;
      6013: inst = 32'h8220000;
      6014: inst = 32'h10408000;
      6015: inst = 32'hc404e0d;
      6016: inst = 32'h8220000;
      6017: inst = 32'h10408000;
      6018: inst = 32'hc404e0e;
      6019: inst = 32'h8220000;
      6020: inst = 32'h10408000;
      6021: inst = 32'hc404e37;
      6022: inst = 32'h8220000;
      6023: inst = 32'h10408000;
      6024: inst = 32'hc404e38;
      6025: inst = 32'h8220000;
      6026: inst = 32'h10408000;
      6027: inst = 32'hc404e39;
      6028: inst = 32'h8220000;
      6029: inst = 32'h10408000;
      6030: inst = 32'hc404e3a;
      6031: inst = 32'h8220000;
      6032: inst = 32'h10408000;
      6033: inst = 32'hc404e3b;
      6034: inst = 32'h8220000;
      6035: inst = 32'h10408000;
      6036: inst = 32'hc404e3c;
      6037: inst = 32'h8220000;
      6038: inst = 32'h10408000;
      6039: inst = 32'hc404e3d;
      6040: inst = 32'h8220000;
      6041: inst = 32'h10408000;
      6042: inst = 32'hc404e3e;
      6043: inst = 32'h8220000;
      6044: inst = 32'h10408000;
      6045: inst = 32'hc404e3f;
      6046: inst = 32'h8220000;
      6047: inst = 32'h10408000;
      6048: inst = 32'hc404e40;
      6049: inst = 32'h8220000;
      6050: inst = 32'h10408000;
      6051: inst = 32'hc404e41;
      6052: inst = 32'h8220000;
      6053: inst = 32'h10408000;
      6054: inst = 32'hc404e42;
      6055: inst = 32'h8220000;
      6056: inst = 32'h10408000;
      6057: inst = 32'hc404e43;
      6058: inst = 32'h8220000;
      6059: inst = 32'h10408000;
      6060: inst = 32'hc404e44;
      6061: inst = 32'h8220000;
      6062: inst = 32'h10408000;
      6063: inst = 32'hc404e45;
      6064: inst = 32'h8220000;
      6065: inst = 32'h10408000;
      6066: inst = 32'hc404e46;
      6067: inst = 32'h8220000;
      6068: inst = 32'h10408000;
      6069: inst = 32'hc404e47;
      6070: inst = 32'h8220000;
      6071: inst = 32'h10408000;
      6072: inst = 32'hc404e48;
      6073: inst = 32'h8220000;
      6074: inst = 32'h10408000;
      6075: inst = 32'hc404e49;
      6076: inst = 32'h8220000;
      6077: inst = 32'h10408000;
      6078: inst = 32'hc404e4a;
      6079: inst = 32'h8220000;
      6080: inst = 32'h10408000;
      6081: inst = 32'hc404e4b;
      6082: inst = 32'h8220000;
      6083: inst = 32'h10408000;
      6084: inst = 32'hc404e4c;
      6085: inst = 32'h8220000;
      6086: inst = 32'h10408000;
      6087: inst = 32'hc404e4d;
      6088: inst = 32'h8220000;
      6089: inst = 32'h10408000;
      6090: inst = 32'hc404e4e;
      6091: inst = 32'h8220000;
      6092: inst = 32'h10408000;
      6093: inst = 32'hc404e4f;
      6094: inst = 32'h8220000;
      6095: inst = 32'h10408000;
      6096: inst = 32'hc404e50;
      6097: inst = 32'h8220000;
      6098: inst = 32'h10408000;
      6099: inst = 32'hc404e51;
      6100: inst = 32'h8220000;
      6101: inst = 32'h10408000;
      6102: inst = 32'hc404e52;
      6103: inst = 32'h8220000;
      6104: inst = 32'h10408000;
      6105: inst = 32'hc404e53;
      6106: inst = 32'h8220000;
      6107: inst = 32'h10408000;
      6108: inst = 32'hc404e54;
      6109: inst = 32'h8220000;
      6110: inst = 32'h10408000;
      6111: inst = 32'hc404e55;
      6112: inst = 32'h8220000;
      6113: inst = 32'h10408000;
      6114: inst = 32'hc404e56;
      6115: inst = 32'h8220000;
      6116: inst = 32'h10408000;
      6117: inst = 32'hc404e57;
      6118: inst = 32'h8220000;
      6119: inst = 32'h10408000;
      6120: inst = 32'hc404e58;
      6121: inst = 32'h8220000;
      6122: inst = 32'h10408000;
      6123: inst = 32'hc404e59;
      6124: inst = 32'h8220000;
      6125: inst = 32'h10408000;
      6126: inst = 32'hc404e5a;
      6127: inst = 32'h8220000;
      6128: inst = 32'h10408000;
      6129: inst = 32'hc404e5b;
      6130: inst = 32'h8220000;
      6131: inst = 32'h10408000;
      6132: inst = 32'hc404e5c;
      6133: inst = 32'h8220000;
      6134: inst = 32'h10408000;
      6135: inst = 32'hc404e5d;
      6136: inst = 32'h8220000;
      6137: inst = 32'h10408000;
      6138: inst = 32'hc404e5e;
      6139: inst = 32'h8220000;
      6140: inst = 32'h10408000;
      6141: inst = 32'hc404e5f;
      6142: inst = 32'h8220000;
      6143: inst = 32'h10408000;
      6144: inst = 32'hc404e60;
      6145: inst = 32'h8220000;
      6146: inst = 32'h10408000;
      6147: inst = 32'hc404e61;
      6148: inst = 32'h8220000;
      6149: inst = 32'h10408000;
      6150: inst = 32'hc404e62;
      6151: inst = 32'h8220000;
      6152: inst = 32'h10408000;
      6153: inst = 32'hc404e63;
      6154: inst = 32'h8220000;
      6155: inst = 32'h10408000;
      6156: inst = 32'hc404e64;
      6157: inst = 32'h8220000;
      6158: inst = 32'h10408000;
      6159: inst = 32'hc404e65;
      6160: inst = 32'h8220000;
      6161: inst = 32'h10408000;
      6162: inst = 32'hc404e66;
      6163: inst = 32'h8220000;
      6164: inst = 32'h10408000;
      6165: inst = 32'hc404e67;
      6166: inst = 32'h8220000;
      6167: inst = 32'h10408000;
      6168: inst = 32'hc404e68;
      6169: inst = 32'h8220000;
      6170: inst = 32'h10408000;
      6171: inst = 32'hc404e69;
      6172: inst = 32'h8220000;
      6173: inst = 32'h10408000;
      6174: inst = 32'hc404e6a;
      6175: inst = 32'h8220000;
      6176: inst = 32'h10408000;
      6177: inst = 32'hc404e6b;
      6178: inst = 32'h8220000;
      6179: inst = 32'h10408000;
      6180: inst = 32'hc404e6c;
      6181: inst = 32'h8220000;
      6182: inst = 32'h10408000;
      6183: inst = 32'hc404e6d;
      6184: inst = 32'h8220000;
      6185: inst = 32'h10408000;
      6186: inst = 32'hc404e6e;
      6187: inst = 32'h8220000;
      6188: inst = 32'h10408000;
      6189: inst = 32'hc404e97;
      6190: inst = 32'h8220000;
      6191: inst = 32'h10408000;
      6192: inst = 32'hc404e98;
      6193: inst = 32'h8220000;
      6194: inst = 32'h10408000;
      6195: inst = 32'hc404e99;
      6196: inst = 32'h8220000;
      6197: inst = 32'h10408000;
      6198: inst = 32'hc404e9a;
      6199: inst = 32'h8220000;
      6200: inst = 32'h10408000;
      6201: inst = 32'hc404e9b;
      6202: inst = 32'h8220000;
      6203: inst = 32'h10408000;
      6204: inst = 32'hc404e9c;
      6205: inst = 32'h8220000;
      6206: inst = 32'h10408000;
      6207: inst = 32'hc404e9d;
      6208: inst = 32'h8220000;
      6209: inst = 32'h10408000;
      6210: inst = 32'hc404e9e;
      6211: inst = 32'h8220000;
      6212: inst = 32'h10408000;
      6213: inst = 32'hc404ea8;
      6214: inst = 32'h8220000;
      6215: inst = 32'h10408000;
      6216: inst = 32'hc404ea9;
      6217: inst = 32'h8220000;
      6218: inst = 32'h10408000;
      6219: inst = 32'hc404eaa;
      6220: inst = 32'h8220000;
      6221: inst = 32'h10408000;
      6222: inst = 32'hc404eab;
      6223: inst = 32'h8220000;
      6224: inst = 32'h10408000;
      6225: inst = 32'hc404eac;
      6226: inst = 32'h8220000;
      6227: inst = 32'h10408000;
      6228: inst = 32'hc404ead;
      6229: inst = 32'h8220000;
      6230: inst = 32'h10408000;
      6231: inst = 32'hc404eae;
      6232: inst = 32'h8220000;
      6233: inst = 32'h10408000;
      6234: inst = 32'hc404eaf;
      6235: inst = 32'h8220000;
      6236: inst = 32'h10408000;
      6237: inst = 32'hc404eb0;
      6238: inst = 32'h8220000;
      6239: inst = 32'h10408000;
      6240: inst = 32'hc404eb1;
      6241: inst = 32'h8220000;
      6242: inst = 32'h10408000;
      6243: inst = 32'hc404eb2;
      6244: inst = 32'h8220000;
      6245: inst = 32'h10408000;
      6246: inst = 32'hc404eb3;
      6247: inst = 32'h8220000;
      6248: inst = 32'h10408000;
      6249: inst = 32'hc404eb4;
      6250: inst = 32'h8220000;
      6251: inst = 32'h10408000;
      6252: inst = 32'hc404eb5;
      6253: inst = 32'h8220000;
      6254: inst = 32'h10408000;
      6255: inst = 32'hc404eb6;
      6256: inst = 32'h8220000;
      6257: inst = 32'h10408000;
      6258: inst = 32'hc404eb7;
      6259: inst = 32'h8220000;
      6260: inst = 32'h10408000;
      6261: inst = 32'hc404ec1;
      6262: inst = 32'h8220000;
      6263: inst = 32'h10408000;
      6264: inst = 32'hc404ec2;
      6265: inst = 32'h8220000;
      6266: inst = 32'h10408000;
      6267: inst = 32'hc404ec3;
      6268: inst = 32'h8220000;
      6269: inst = 32'h10408000;
      6270: inst = 32'hc404ec4;
      6271: inst = 32'h8220000;
      6272: inst = 32'h10408000;
      6273: inst = 32'hc404ec5;
      6274: inst = 32'h8220000;
      6275: inst = 32'h10408000;
      6276: inst = 32'hc404ec6;
      6277: inst = 32'h8220000;
      6278: inst = 32'h10408000;
      6279: inst = 32'hc404ec7;
      6280: inst = 32'h8220000;
      6281: inst = 32'h10408000;
      6282: inst = 32'hc404ec8;
      6283: inst = 32'h8220000;
      6284: inst = 32'h10408000;
      6285: inst = 32'hc404ec9;
      6286: inst = 32'h8220000;
      6287: inst = 32'h10408000;
      6288: inst = 32'hc404eca;
      6289: inst = 32'h8220000;
      6290: inst = 32'h10408000;
      6291: inst = 32'hc404ecb;
      6292: inst = 32'h8220000;
      6293: inst = 32'h10408000;
      6294: inst = 32'hc404ecc;
      6295: inst = 32'h8220000;
      6296: inst = 32'h10408000;
      6297: inst = 32'hc404ecd;
      6298: inst = 32'h8220000;
      6299: inst = 32'h10408000;
      6300: inst = 32'hc404ece;
      6301: inst = 32'h8220000;
      6302: inst = 32'h10408000;
      6303: inst = 32'hc404ef7;
      6304: inst = 32'h8220000;
      6305: inst = 32'h10408000;
      6306: inst = 32'hc404ef8;
      6307: inst = 32'h8220000;
      6308: inst = 32'h10408000;
      6309: inst = 32'hc404ef9;
      6310: inst = 32'h8220000;
      6311: inst = 32'h10408000;
      6312: inst = 32'hc404efa;
      6313: inst = 32'h8220000;
      6314: inst = 32'h10408000;
      6315: inst = 32'hc404efb;
      6316: inst = 32'h8220000;
      6317: inst = 32'h10408000;
      6318: inst = 32'hc404efc;
      6319: inst = 32'h8220000;
      6320: inst = 32'h10408000;
      6321: inst = 32'hc404efd;
      6322: inst = 32'h8220000;
      6323: inst = 32'h10408000;
      6324: inst = 32'hc404efe;
      6325: inst = 32'h8220000;
      6326: inst = 32'h10408000;
      6327: inst = 32'hc404f08;
      6328: inst = 32'h8220000;
      6329: inst = 32'h10408000;
      6330: inst = 32'hc404f09;
      6331: inst = 32'h8220000;
      6332: inst = 32'h10408000;
      6333: inst = 32'hc404f0a;
      6334: inst = 32'h8220000;
      6335: inst = 32'h10408000;
      6336: inst = 32'hc404f0b;
      6337: inst = 32'h8220000;
      6338: inst = 32'h10408000;
      6339: inst = 32'hc404f0c;
      6340: inst = 32'h8220000;
      6341: inst = 32'h10408000;
      6342: inst = 32'hc404f0d;
      6343: inst = 32'h8220000;
      6344: inst = 32'h10408000;
      6345: inst = 32'hc404f0e;
      6346: inst = 32'h8220000;
      6347: inst = 32'h10408000;
      6348: inst = 32'hc404f0f;
      6349: inst = 32'h8220000;
      6350: inst = 32'h10408000;
      6351: inst = 32'hc404f10;
      6352: inst = 32'h8220000;
      6353: inst = 32'h10408000;
      6354: inst = 32'hc404f11;
      6355: inst = 32'h8220000;
      6356: inst = 32'h10408000;
      6357: inst = 32'hc404f12;
      6358: inst = 32'h8220000;
      6359: inst = 32'h10408000;
      6360: inst = 32'hc404f13;
      6361: inst = 32'h8220000;
      6362: inst = 32'h10408000;
      6363: inst = 32'hc404f14;
      6364: inst = 32'h8220000;
      6365: inst = 32'h10408000;
      6366: inst = 32'hc404f15;
      6367: inst = 32'h8220000;
      6368: inst = 32'h10408000;
      6369: inst = 32'hc404f16;
      6370: inst = 32'h8220000;
      6371: inst = 32'h10408000;
      6372: inst = 32'hc404f17;
      6373: inst = 32'h8220000;
      6374: inst = 32'h10408000;
      6375: inst = 32'hc404f21;
      6376: inst = 32'h8220000;
      6377: inst = 32'h10408000;
      6378: inst = 32'hc404f22;
      6379: inst = 32'h8220000;
      6380: inst = 32'h10408000;
      6381: inst = 32'hc404f23;
      6382: inst = 32'h8220000;
      6383: inst = 32'h10408000;
      6384: inst = 32'hc404f24;
      6385: inst = 32'h8220000;
      6386: inst = 32'h10408000;
      6387: inst = 32'hc404f25;
      6388: inst = 32'h8220000;
      6389: inst = 32'h10408000;
      6390: inst = 32'hc404f26;
      6391: inst = 32'h8220000;
      6392: inst = 32'h10408000;
      6393: inst = 32'hc404f27;
      6394: inst = 32'h8220000;
      6395: inst = 32'h10408000;
      6396: inst = 32'hc404f28;
      6397: inst = 32'h8220000;
      6398: inst = 32'h10408000;
      6399: inst = 32'hc404f29;
      6400: inst = 32'h8220000;
      6401: inst = 32'h10408000;
      6402: inst = 32'hc404f2a;
      6403: inst = 32'h8220000;
      6404: inst = 32'h10408000;
      6405: inst = 32'hc404f2b;
      6406: inst = 32'h8220000;
      6407: inst = 32'h10408000;
      6408: inst = 32'hc404f2c;
      6409: inst = 32'h8220000;
      6410: inst = 32'h10408000;
      6411: inst = 32'hc404f2d;
      6412: inst = 32'h8220000;
      6413: inst = 32'h10408000;
      6414: inst = 32'hc404f2e;
      6415: inst = 32'h8220000;
      6416: inst = 32'h10408000;
      6417: inst = 32'hc404f57;
      6418: inst = 32'h8220000;
      6419: inst = 32'h10408000;
      6420: inst = 32'hc404f58;
      6421: inst = 32'h8220000;
      6422: inst = 32'h10408000;
      6423: inst = 32'hc404f59;
      6424: inst = 32'h8220000;
      6425: inst = 32'h10408000;
      6426: inst = 32'hc404f5a;
      6427: inst = 32'h8220000;
      6428: inst = 32'h10408000;
      6429: inst = 32'hc404f5b;
      6430: inst = 32'h8220000;
      6431: inst = 32'h10408000;
      6432: inst = 32'hc404f5c;
      6433: inst = 32'h8220000;
      6434: inst = 32'h10408000;
      6435: inst = 32'hc404f5d;
      6436: inst = 32'h8220000;
      6437: inst = 32'h10408000;
      6438: inst = 32'hc404f5e;
      6439: inst = 32'h8220000;
      6440: inst = 32'h10408000;
      6441: inst = 32'hc404f68;
      6442: inst = 32'h8220000;
      6443: inst = 32'h10408000;
      6444: inst = 32'hc404f69;
      6445: inst = 32'h8220000;
      6446: inst = 32'h10408000;
      6447: inst = 32'hc404f6a;
      6448: inst = 32'h8220000;
      6449: inst = 32'h10408000;
      6450: inst = 32'hc404f6b;
      6451: inst = 32'h8220000;
      6452: inst = 32'h10408000;
      6453: inst = 32'hc404f6c;
      6454: inst = 32'h8220000;
      6455: inst = 32'h10408000;
      6456: inst = 32'hc404f6d;
      6457: inst = 32'h8220000;
      6458: inst = 32'h10408000;
      6459: inst = 32'hc404f6e;
      6460: inst = 32'h8220000;
      6461: inst = 32'h10408000;
      6462: inst = 32'hc404f6f;
      6463: inst = 32'h8220000;
      6464: inst = 32'h10408000;
      6465: inst = 32'hc404f70;
      6466: inst = 32'h8220000;
      6467: inst = 32'h10408000;
      6468: inst = 32'hc404f71;
      6469: inst = 32'h8220000;
      6470: inst = 32'h10408000;
      6471: inst = 32'hc404f72;
      6472: inst = 32'h8220000;
      6473: inst = 32'h10408000;
      6474: inst = 32'hc404f73;
      6475: inst = 32'h8220000;
      6476: inst = 32'h10408000;
      6477: inst = 32'hc404f74;
      6478: inst = 32'h8220000;
      6479: inst = 32'h10408000;
      6480: inst = 32'hc404f75;
      6481: inst = 32'h8220000;
      6482: inst = 32'h10408000;
      6483: inst = 32'hc404f76;
      6484: inst = 32'h8220000;
      6485: inst = 32'h10408000;
      6486: inst = 32'hc404f77;
      6487: inst = 32'h8220000;
      6488: inst = 32'h10408000;
      6489: inst = 32'hc404f81;
      6490: inst = 32'h8220000;
      6491: inst = 32'h10408000;
      6492: inst = 32'hc404f82;
      6493: inst = 32'h8220000;
      6494: inst = 32'h10408000;
      6495: inst = 32'hc404f83;
      6496: inst = 32'h8220000;
      6497: inst = 32'h10408000;
      6498: inst = 32'hc404f84;
      6499: inst = 32'h8220000;
      6500: inst = 32'h10408000;
      6501: inst = 32'hc404f85;
      6502: inst = 32'h8220000;
      6503: inst = 32'h10408000;
      6504: inst = 32'hc404f86;
      6505: inst = 32'h8220000;
      6506: inst = 32'h10408000;
      6507: inst = 32'hc404f87;
      6508: inst = 32'h8220000;
      6509: inst = 32'h10408000;
      6510: inst = 32'hc404f88;
      6511: inst = 32'h8220000;
      6512: inst = 32'h10408000;
      6513: inst = 32'hc404f89;
      6514: inst = 32'h8220000;
      6515: inst = 32'h10408000;
      6516: inst = 32'hc404f8a;
      6517: inst = 32'h8220000;
      6518: inst = 32'h10408000;
      6519: inst = 32'hc404f8b;
      6520: inst = 32'h8220000;
      6521: inst = 32'h10408000;
      6522: inst = 32'hc404f8c;
      6523: inst = 32'h8220000;
      6524: inst = 32'h10408000;
      6525: inst = 32'hc404f8d;
      6526: inst = 32'h8220000;
      6527: inst = 32'h10408000;
      6528: inst = 32'hc404f8e;
      6529: inst = 32'h8220000;
      6530: inst = 32'h10408000;
      6531: inst = 32'hc404fb7;
      6532: inst = 32'h8220000;
      6533: inst = 32'h10408000;
      6534: inst = 32'hc404fb8;
      6535: inst = 32'h8220000;
      6536: inst = 32'h10408000;
      6537: inst = 32'hc404fb9;
      6538: inst = 32'h8220000;
      6539: inst = 32'h10408000;
      6540: inst = 32'hc404fba;
      6541: inst = 32'h8220000;
      6542: inst = 32'h10408000;
      6543: inst = 32'hc404fbb;
      6544: inst = 32'h8220000;
      6545: inst = 32'h10408000;
      6546: inst = 32'hc404fbc;
      6547: inst = 32'h8220000;
      6548: inst = 32'h10408000;
      6549: inst = 32'hc404fbd;
      6550: inst = 32'h8220000;
      6551: inst = 32'h10408000;
      6552: inst = 32'hc404fbe;
      6553: inst = 32'h8220000;
      6554: inst = 32'h10408000;
      6555: inst = 32'hc404fc8;
      6556: inst = 32'h8220000;
      6557: inst = 32'h10408000;
      6558: inst = 32'hc404fc9;
      6559: inst = 32'h8220000;
      6560: inst = 32'h10408000;
      6561: inst = 32'hc404fca;
      6562: inst = 32'h8220000;
      6563: inst = 32'h10408000;
      6564: inst = 32'hc404fcb;
      6565: inst = 32'h8220000;
      6566: inst = 32'h10408000;
      6567: inst = 32'hc404fcc;
      6568: inst = 32'h8220000;
      6569: inst = 32'h10408000;
      6570: inst = 32'hc404fcd;
      6571: inst = 32'h8220000;
      6572: inst = 32'h10408000;
      6573: inst = 32'hc404fce;
      6574: inst = 32'h8220000;
      6575: inst = 32'h10408000;
      6576: inst = 32'hc404fcf;
      6577: inst = 32'h8220000;
      6578: inst = 32'h10408000;
      6579: inst = 32'hc404fd0;
      6580: inst = 32'h8220000;
      6581: inst = 32'h10408000;
      6582: inst = 32'hc404fd1;
      6583: inst = 32'h8220000;
      6584: inst = 32'h10408000;
      6585: inst = 32'hc404fd2;
      6586: inst = 32'h8220000;
      6587: inst = 32'h10408000;
      6588: inst = 32'hc404fd3;
      6589: inst = 32'h8220000;
      6590: inst = 32'h10408000;
      6591: inst = 32'hc404fd4;
      6592: inst = 32'h8220000;
      6593: inst = 32'h10408000;
      6594: inst = 32'hc404fd5;
      6595: inst = 32'h8220000;
      6596: inst = 32'h10408000;
      6597: inst = 32'hc404fd6;
      6598: inst = 32'h8220000;
      6599: inst = 32'h10408000;
      6600: inst = 32'hc404fd7;
      6601: inst = 32'h8220000;
      6602: inst = 32'h10408000;
      6603: inst = 32'hc404fe1;
      6604: inst = 32'h8220000;
      6605: inst = 32'h10408000;
      6606: inst = 32'hc404fe2;
      6607: inst = 32'h8220000;
      6608: inst = 32'h10408000;
      6609: inst = 32'hc404fe3;
      6610: inst = 32'h8220000;
      6611: inst = 32'h10408000;
      6612: inst = 32'hc404fe4;
      6613: inst = 32'h8220000;
      6614: inst = 32'h10408000;
      6615: inst = 32'hc404fe5;
      6616: inst = 32'h8220000;
      6617: inst = 32'h10408000;
      6618: inst = 32'hc404fe6;
      6619: inst = 32'h8220000;
      6620: inst = 32'h10408000;
      6621: inst = 32'hc404fe7;
      6622: inst = 32'h8220000;
      6623: inst = 32'h10408000;
      6624: inst = 32'hc404fe8;
      6625: inst = 32'h8220000;
      6626: inst = 32'h10408000;
      6627: inst = 32'hc404fe9;
      6628: inst = 32'h8220000;
      6629: inst = 32'h10408000;
      6630: inst = 32'hc404fea;
      6631: inst = 32'h8220000;
      6632: inst = 32'h10408000;
      6633: inst = 32'hc404feb;
      6634: inst = 32'h8220000;
      6635: inst = 32'h10408000;
      6636: inst = 32'hc404fec;
      6637: inst = 32'h8220000;
      6638: inst = 32'h10408000;
      6639: inst = 32'hc404fed;
      6640: inst = 32'h8220000;
      6641: inst = 32'h10408000;
      6642: inst = 32'hc404fee;
      6643: inst = 32'h8220000;
      6644: inst = 32'h10408000;
      6645: inst = 32'hc405017;
      6646: inst = 32'h8220000;
      6647: inst = 32'h10408000;
      6648: inst = 32'hc405018;
      6649: inst = 32'h8220000;
      6650: inst = 32'h10408000;
      6651: inst = 32'hc405019;
      6652: inst = 32'h8220000;
      6653: inst = 32'h10408000;
      6654: inst = 32'hc40501a;
      6655: inst = 32'h8220000;
      6656: inst = 32'h10408000;
      6657: inst = 32'hc40501b;
      6658: inst = 32'h8220000;
      6659: inst = 32'h10408000;
      6660: inst = 32'hc40501c;
      6661: inst = 32'h8220000;
      6662: inst = 32'h10408000;
      6663: inst = 32'hc40501d;
      6664: inst = 32'h8220000;
      6665: inst = 32'h10408000;
      6666: inst = 32'hc40501e;
      6667: inst = 32'h8220000;
      6668: inst = 32'h10408000;
      6669: inst = 32'hc405028;
      6670: inst = 32'h8220000;
      6671: inst = 32'h10408000;
      6672: inst = 32'hc405029;
      6673: inst = 32'h8220000;
      6674: inst = 32'h10408000;
      6675: inst = 32'hc40502a;
      6676: inst = 32'h8220000;
      6677: inst = 32'h10408000;
      6678: inst = 32'hc40502b;
      6679: inst = 32'h8220000;
      6680: inst = 32'h10408000;
      6681: inst = 32'hc40502c;
      6682: inst = 32'h8220000;
      6683: inst = 32'h10408000;
      6684: inst = 32'hc40502d;
      6685: inst = 32'h8220000;
      6686: inst = 32'h10408000;
      6687: inst = 32'hc40502e;
      6688: inst = 32'h8220000;
      6689: inst = 32'h10408000;
      6690: inst = 32'hc40502f;
      6691: inst = 32'h8220000;
      6692: inst = 32'h10408000;
      6693: inst = 32'hc405030;
      6694: inst = 32'h8220000;
      6695: inst = 32'h10408000;
      6696: inst = 32'hc405031;
      6697: inst = 32'h8220000;
      6698: inst = 32'h10408000;
      6699: inst = 32'hc405032;
      6700: inst = 32'h8220000;
      6701: inst = 32'h10408000;
      6702: inst = 32'hc405033;
      6703: inst = 32'h8220000;
      6704: inst = 32'h10408000;
      6705: inst = 32'hc405034;
      6706: inst = 32'h8220000;
      6707: inst = 32'h10408000;
      6708: inst = 32'hc405035;
      6709: inst = 32'h8220000;
      6710: inst = 32'h10408000;
      6711: inst = 32'hc405036;
      6712: inst = 32'h8220000;
      6713: inst = 32'h10408000;
      6714: inst = 32'hc405037;
      6715: inst = 32'h8220000;
      6716: inst = 32'h10408000;
      6717: inst = 32'hc405041;
      6718: inst = 32'h8220000;
      6719: inst = 32'h10408000;
      6720: inst = 32'hc405042;
      6721: inst = 32'h8220000;
      6722: inst = 32'h10408000;
      6723: inst = 32'hc405043;
      6724: inst = 32'h8220000;
      6725: inst = 32'h10408000;
      6726: inst = 32'hc405044;
      6727: inst = 32'h8220000;
      6728: inst = 32'h10408000;
      6729: inst = 32'hc405045;
      6730: inst = 32'h8220000;
      6731: inst = 32'h10408000;
      6732: inst = 32'hc405046;
      6733: inst = 32'h8220000;
      6734: inst = 32'h10408000;
      6735: inst = 32'hc405047;
      6736: inst = 32'h8220000;
      6737: inst = 32'h10408000;
      6738: inst = 32'hc405048;
      6739: inst = 32'h8220000;
      6740: inst = 32'h10408000;
      6741: inst = 32'hc405049;
      6742: inst = 32'h8220000;
      6743: inst = 32'h10408000;
      6744: inst = 32'hc40504a;
      6745: inst = 32'h8220000;
      6746: inst = 32'h10408000;
      6747: inst = 32'hc40504b;
      6748: inst = 32'h8220000;
      6749: inst = 32'h10408000;
      6750: inst = 32'hc40504c;
      6751: inst = 32'h8220000;
      6752: inst = 32'h10408000;
      6753: inst = 32'hc40504d;
      6754: inst = 32'h8220000;
      6755: inst = 32'h10408000;
      6756: inst = 32'hc40504e;
      6757: inst = 32'h8220000;
      6758: inst = 32'h10408000;
      6759: inst = 32'hc405077;
      6760: inst = 32'h8220000;
      6761: inst = 32'h10408000;
      6762: inst = 32'hc405078;
      6763: inst = 32'h8220000;
      6764: inst = 32'h10408000;
      6765: inst = 32'hc405079;
      6766: inst = 32'h8220000;
      6767: inst = 32'h10408000;
      6768: inst = 32'hc40507a;
      6769: inst = 32'h8220000;
      6770: inst = 32'h10408000;
      6771: inst = 32'hc40507b;
      6772: inst = 32'h8220000;
      6773: inst = 32'h10408000;
      6774: inst = 32'hc40507c;
      6775: inst = 32'h8220000;
      6776: inst = 32'h10408000;
      6777: inst = 32'hc40507d;
      6778: inst = 32'h8220000;
      6779: inst = 32'h10408000;
      6780: inst = 32'hc40507e;
      6781: inst = 32'h8220000;
      6782: inst = 32'h10408000;
      6783: inst = 32'hc405088;
      6784: inst = 32'h8220000;
      6785: inst = 32'h10408000;
      6786: inst = 32'hc405089;
      6787: inst = 32'h8220000;
      6788: inst = 32'h10408000;
      6789: inst = 32'hc40508a;
      6790: inst = 32'h8220000;
      6791: inst = 32'h10408000;
      6792: inst = 32'hc40508b;
      6793: inst = 32'h8220000;
      6794: inst = 32'h10408000;
      6795: inst = 32'hc40508c;
      6796: inst = 32'h8220000;
      6797: inst = 32'h10408000;
      6798: inst = 32'hc40508d;
      6799: inst = 32'h8220000;
      6800: inst = 32'h10408000;
      6801: inst = 32'hc40508e;
      6802: inst = 32'h8220000;
      6803: inst = 32'h10408000;
      6804: inst = 32'hc40508f;
      6805: inst = 32'h8220000;
      6806: inst = 32'h10408000;
      6807: inst = 32'hc405090;
      6808: inst = 32'h8220000;
      6809: inst = 32'h10408000;
      6810: inst = 32'hc405091;
      6811: inst = 32'h8220000;
      6812: inst = 32'h10408000;
      6813: inst = 32'hc405092;
      6814: inst = 32'h8220000;
      6815: inst = 32'h10408000;
      6816: inst = 32'hc405093;
      6817: inst = 32'h8220000;
      6818: inst = 32'h10408000;
      6819: inst = 32'hc405094;
      6820: inst = 32'h8220000;
      6821: inst = 32'h10408000;
      6822: inst = 32'hc405095;
      6823: inst = 32'h8220000;
      6824: inst = 32'h10408000;
      6825: inst = 32'hc405096;
      6826: inst = 32'h8220000;
      6827: inst = 32'h10408000;
      6828: inst = 32'hc405097;
      6829: inst = 32'h8220000;
      6830: inst = 32'h10408000;
      6831: inst = 32'hc4050a1;
      6832: inst = 32'h8220000;
      6833: inst = 32'h10408000;
      6834: inst = 32'hc4050a2;
      6835: inst = 32'h8220000;
      6836: inst = 32'h10408000;
      6837: inst = 32'hc4050a3;
      6838: inst = 32'h8220000;
      6839: inst = 32'h10408000;
      6840: inst = 32'hc4050a4;
      6841: inst = 32'h8220000;
      6842: inst = 32'h10408000;
      6843: inst = 32'hc4050a5;
      6844: inst = 32'h8220000;
      6845: inst = 32'h10408000;
      6846: inst = 32'hc4050a6;
      6847: inst = 32'h8220000;
      6848: inst = 32'h10408000;
      6849: inst = 32'hc4050a7;
      6850: inst = 32'h8220000;
      6851: inst = 32'h10408000;
      6852: inst = 32'hc4050a8;
      6853: inst = 32'h8220000;
      6854: inst = 32'h10408000;
      6855: inst = 32'hc4050a9;
      6856: inst = 32'h8220000;
      6857: inst = 32'h10408000;
      6858: inst = 32'hc4050aa;
      6859: inst = 32'h8220000;
      6860: inst = 32'h10408000;
      6861: inst = 32'hc4050ab;
      6862: inst = 32'h8220000;
      6863: inst = 32'h10408000;
      6864: inst = 32'hc4050ac;
      6865: inst = 32'h8220000;
      6866: inst = 32'h10408000;
      6867: inst = 32'hc4050ad;
      6868: inst = 32'h8220000;
      6869: inst = 32'h10408000;
      6870: inst = 32'hc4050ae;
      6871: inst = 32'h8220000;
      6872: inst = 32'h10408000;
      6873: inst = 32'hc4050d7;
      6874: inst = 32'h8220000;
      6875: inst = 32'h10408000;
      6876: inst = 32'hc4050d8;
      6877: inst = 32'h8220000;
      6878: inst = 32'h10408000;
      6879: inst = 32'hc4050d9;
      6880: inst = 32'h8220000;
      6881: inst = 32'h10408000;
      6882: inst = 32'hc4050da;
      6883: inst = 32'h8220000;
      6884: inst = 32'h10408000;
      6885: inst = 32'hc4050db;
      6886: inst = 32'h8220000;
      6887: inst = 32'h10408000;
      6888: inst = 32'hc4050dc;
      6889: inst = 32'h8220000;
      6890: inst = 32'h10408000;
      6891: inst = 32'hc4050dd;
      6892: inst = 32'h8220000;
      6893: inst = 32'h10408000;
      6894: inst = 32'hc4050de;
      6895: inst = 32'h8220000;
      6896: inst = 32'h10408000;
      6897: inst = 32'hc4050e8;
      6898: inst = 32'h8220000;
      6899: inst = 32'h10408000;
      6900: inst = 32'hc4050e9;
      6901: inst = 32'h8220000;
      6902: inst = 32'h10408000;
      6903: inst = 32'hc4050ea;
      6904: inst = 32'h8220000;
      6905: inst = 32'h10408000;
      6906: inst = 32'hc4050eb;
      6907: inst = 32'h8220000;
      6908: inst = 32'h10408000;
      6909: inst = 32'hc4050ec;
      6910: inst = 32'h8220000;
      6911: inst = 32'h10408000;
      6912: inst = 32'hc4050ed;
      6913: inst = 32'h8220000;
      6914: inst = 32'h10408000;
      6915: inst = 32'hc4050ee;
      6916: inst = 32'h8220000;
      6917: inst = 32'h10408000;
      6918: inst = 32'hc4050ef;
      6919: inst = 32'h8220000;
      6920: inst = 32'h10408000;
      6921: inst = 32'hc4050f0;
      6922: inst = 32'h8220000;
      6923: inst = 32'h10408000;
      6924: inst = 32'hc4050f1;
      6925: inst = 32'h8220000;
      6926: inst = 32'h10408000;
      6927: inst = 32'hc4050f2;
      6928: inst = 32'h8220000;
      6929: inst = 32'h10408000;
      6930: inst = 32'hc4050f3;
      6931: inst = 32'h8220000;
      6932: inst = 32'h10408000;
      6933: inst = 32'hc4050f4;
      6934: inst = 32'h8220000;
      6935: inst = 32'h10408000;
      6936: inst = 32'hc4050f5;
      6937: inst = 32'h8220000;
      6938: inst = 32'h10408000;
      6939: inst = 32'hc4050f6;
      6940: inst = 32'h8220000;
      6941: inst = 32'h10408000;
      6942: inst = 32'hc4050f7;
      6943: inst = 32'h8220000;
      6944: inst = 32'h10408000;
      6945: inst = 32'hc405101;
      6946: inst = 32'h8220000;
      6947: inst = 32'h10408000;
      6948: inst = 32'hc405102;
      6949: inst = 32'h8220000;
      6950: inst = 32'h10408000;
      6951: inst = 32'hc405103;
      6952: inst = 32'h8220000;
      6953: inst = 32'h10408000;
      6954: inst = 32'hc405104;
      6955: inst = 32'h8220000;
      6956: inst = 32'h10408000;
      6957: inst = 32'hc405105;
      6958: inst = 32'h8220000;
      6959: inst = 32'h10408000;
      6960: inst = 32'hc405106;
      6961: inst = 32'h8220000;
      6962: inst = 32'h10408000;
      6963: inst = 32'hc405107;
      6964: inst = 32'h8220000;
      6965: inst = 32'h10408000;
      6966: inst = 32'hc405108;
      6967: inst = 32'h8220000;
      6968: inst = 32'h10408000;
      6969: inst = 32'hc405109;
      6970: inst = 32'h8220000;
      6971: inst = 32'h10408000;
      6972: inst = 32'hc40510a;
      6973: inst = 32'h8220000;
      6974: inst = 32'h10408000;
      6975: inst = 32'hc40510b;
      6976: inst = 32'h8220000;
      6977: inst = 32'h10408000;
      6978: inst = 32'hc40510c;
      6979: inst = 32'h8220000;
      6980: inst = 32'h10408000;
      6981: inst = 32'hc40510d;
      6982: inst = 32'h8220000;
      6983: inst = 32'h10408000;
      6984: inst = 32'hc40510e;
      6985: inst = 32'h8220000;
      6986: inst = 32'h10408000;
      6987: inst = 32'hc405137;
      6988: inst = 32'h8220000;
      6989: inst = 32'h10408000;
      6990: inst = 32'hc405138;
      6991: inst = 32'h8220000;
      6992: inst = 32'h10408000;
      6993: inst = 32'hc405139;
      6994: inst = 32'h8220000;
      6995: inst = 32'h10408000;
      6996: inst = 32'hc40513a;
      6997: inst = 32'h8220000;
      6998: inst = 32'h10408000;
      6999: inst = 32'hc40513b;
      7000: inst = 32'h8220000;
      7001: inst = 32'h10408000;
      7002: inst = 32'hc40513c;
      7003: inst = 32'h8220000;
      7004: inst = 32'h10408000;
      7005: inst = 32'hc40513d;
      7006: inst = 32'h8220000;
      7007: inst = 32'h10408000;
      7008: inst = 32'hc40513e;
      7009: inst = 32'h8220000;
      7010: inst = 32'h10408000;
      7011: inst = 32'hc405148;
      7012: inst = 32'h8220000;
      7013: inst = 32'h10408000;
      7014: inst = 32'hc405149;
      7015: inst = 32'h8220000;
      7016: inst = 32'h10408000;
      7017: inst = 32'hc40514a;
      7018: inst = 32'h8220000;
      7019: inst = 32'h10408000;
      7020: inst = 32'hc40514b;
      7021: inst = 32'h8220000;
      7022: inst = 32'h10408000;
      7023: inst = 32'hc40514c;
      7024: inst = 32'h8220000;
      7025: inst = 32'h10408000;
      7026: inst = 32'hc40514d;
      7027: inst = 32'h8220000;
      7028: inst = 32'h10408000;
      7029: inst = 32'hc40514e;
      7030: inst = 32'h8220000;
      7031: inst = 32'h10408000;
      7032: inst = 32'hc40514f;
      7033: inst = 32'h8220000;
      7034: inst = 32'h10408000;
      7035: inst = 32'hc405150;
      7036: inst = 32'h8220000;
      7037: inst = 32'h10408000;
      7038: inst = 32'hc405151;
      7039: inst = 32'h8220000;
      7040: inst = 32'h10408000;
      7041: inst = 32'hc405152;
      7042: inst = 32'h8220000;
      7043: inst = 32'h10408000;
      7044: inst = 32'hc405153;
      7045: inst = 32'h8220000;
      7046: inst = 32'h10408000;
      7047: inst = 32'hc405154;
      7048: inst = 32'h8220000;
      7049: inst = 32'h10408000;
      7050: inst = 32'hc405155;
      7051: inst = 32'h8220000;
      7052: inst = 32'h10408000;
      7053: inst = 32'hc405156;
      7054: inst = 32'h8220000;
      7055: inst = 32'h10408000;
      7056: inst = 32'hc405157;
      7057: inst = 32'h8220000;
      7058: inst = 32'h10408000;
      7059: inst = 32'hc405161;
      7060: inst = 32'h8220000;
      7061: inst = 32'h10408000;
      7062: inst = 32'hc405162;
      7063: inst = 32'h8220000;
      7064: inst = 32'h10408000;
      7065: inst = 32'hc405163;
      7066: inst = 32'h8220000;
      7067: inst = 32'h10408000;
      7068: inst = 32'hc405164;
      7069: inst = 32'h8220000;
      7070: inst = 32'h10408000;
      7071: inst = 32'hc405165;
      7072: inst = 32'h8220000;
      7073: inst = 32'h10408000;
      7074: inst = 32'hc405166;
      7075: inst = 32'h8220000;
      7076: inst = 32'h10408000;
      7077: inst = 32'hc405167;
      7078: inst = 32'h8220000;
      7079: inst = 32'h10408000;
      7080: inst = 32'hc405168;
      7081: inst = 32'h8220000;
      7082: inst = 32'h10408000;
      7083: inst = 32'hc405169;
      7084: inst = 32'h8220000;
      7085: inst = 32'h10408000;
      7086: inst = 32'hc40516a;
      7087: inst = 32'h8220000;
      7088: inst = 32'h10408000;
      7089: inst = 32'hc40516b;
      7090: inst = 32'h8220000;
      7091: inst = 32'h10408000;
      7092: inst = 32'hc40516c;
      7093: inst = 32'h8220000;
      7094: inst = 32'h10408000;
      7095: inst = 32'hc40516d;
      7096: inst = 32'h8220000;
      7097: inst = 32'h10408000;
      7098: inst = 32'hc40516e;
      7099: inst = 32'h8220000;
      7100: inst = 32'h10408000;
      7101: inst = 32'hc405197;
      7102: inst = 32'h8220000;
      7103: inst = 32'h10408000;
      7104: inst = 32'hc405198;
      7105: inst = 32'h8220000;
      7106: inst = 32'h10408000;
      7107: inst = 32'hc405199;
      7108: inst = 32'h8220000;
      7109: inst = 32'h10408000;
      7110: inst = 32'hc40519a;
      7111: inst = 32'h8220000;
      7112: inst = 32'h10408000;
      7113: inst = 32'hc40519b;
      7114: inst = 32'h8220000;
      7115: inst = 32'h10408000;
      7116: inst = 32'hc40519c;
      7117: inst = 32'h8220000;
      7118: inst = 32'h10408000;
      7119: inst = 32'hc40519d;
      7120: inst = 32'h8220000;
      7121: inst = 32'h10408000;
      7122: inst = 32'hc4051aa;
      7123: inst = 32'h8220000;
      7124: inst = 32'h10408000;
      7125: inst = 32'hc4051ab;
      7126: inst = 32'h8220000;
      7127: inst = 32'h10408000;
      7128: inst = 32'hc4051ac;
      7129: inst = 32'h8220000;
      7130: inst = 32'h10408000;
      7131: inst = 32'hc4051ad;
      7132: inst = 32'h8220000;
      7133: inst = 32'h10408000;
      7134: inst = 32'hc4051ae;
      7135: inst = 32'h8220000;
      7136: inst = 32'h10408000;
      7137: inst = 32'hc4051af;
      7138: inst = 32'h8220000;
      7139: inst = 32'h10408000;
      7140: inst = 32'hc4051b0;
      7141: inst = 32'h8220000;
      7142: inst = 32'h10408000;
      7143: inst = 32'hc4051b1;
      7144: inst = 32'h8220000;
      7145: inst = 32'h10408000;
      7146: inst = 32'hc4051b2;
      7147: inst = 32'h8220000;
      7148: inst = 32'h10408000;
      7149: inst = 32'hc4051b3;
      7150: inst = 32'h8220000;
      7151: inst = 32'h10408000;
      7152: inst = 32'hc4051b4;
      7153: inst = 32'h8220000;
      7154: inst = 32'h10408000;
      7155: inst = 32'hc4051b5;
      7156: inst = 32'h8220000;
      7157: inst = 32'h10408000;
      7158: inst = 32'hc4051c2;
      7159: inst = 32'h8220000;
      7160: inst = 32'h10408000;
      7161: inst = 32'hc4051c3;
      7162: inst = 32'h8220000;
      7163: inst = 32'h10408000;
      7164: inst = 32'hc4051c4;
      7165: inst = 32'h8220000;
      7166: inst = 32'h10408000;
      7167: inst = 32'hc4051c5;
      7168: inst = 32'h8220000;
      7169: inst = 32'h10408000;
      7170: inst = 32'hc4051c6;
      7171: inst = 32'h8220000;
      7172: inst = 32'h10408000;
      7173: inst = 32'hc4051c7;
      7174: inst = 32'h8220000;
      7175: inst = 32'h10408000;
      7176: inst = 32'hc4051c8;
      7177: inst = 32'h8220000;
      7178: inst = 32'h10408000;
      7179: inst = 32'hc4051c9;
      7180: inst = 32'h8220000;
      7181: inst = 32'h10408000;
      7182: inst = 32'hc4051ca;
      7183: inst = 32'h8220000;
      7184: inst = 32'h10408000;
      7185: inst = 32'hc4051cb;
      7186: inst = 32'h8220000;
      7187: inst = 32'h10408000;
      7188: inst = 32'hc4051cc;
      7189: inst = 32'h8220000;
      7190: inst = 32'h10408000;
      7191: inst = 32'hc4051cd;
      7192: inst = 32'h8220000;
      7193: inst = 32'h10408000;
      7194: inst = 32'hc4051ce;
      7195: inst = 32'h8220000;
      7196: inst = 32'h10408000;
      7197: inst = 32'hc4051f7;
      7198: inst = 32'h8220000;
      7199: inst = 32'h10408000;
      7200: inst = 32'hc4051f8;
      7201: inst = 32'h8220000;
      7202: inst = 32'h10408000;
      7203: inst = 32'hc4051f9;
      7204: inst = 32'h8220000;
      7205: inst = 32'h10408000;
      7206: inst = 32'hc4051fa;
      7207: inst = 32'h8220000;
      7208: inst = 32'h10408000;
      7209: inst = 32'hc4051fb;
      7210: inst = 32'h8220000;
      7211: inst = 32'h10408000;
      7212: inst = 32'hc4051fc;
      7213: inst = 32'h8220000;
      7214: inst = 32'h10408000;
      7215: inst = 32'hc40520a;
      7216: inst = 32'h8220000;
      7217: inst = 32'h10408000;
      7218: inst = 32'hc40520b;
      7219: inst = 32'h8220000;
      7220: inst = 32'h10408000;
      7221: inst = 32'hc40520c;
      7222: inst = 32'h8220000;
      7223: inst = 32'h10408000;
      7224: inst = 32'hc40520d;
      7225: inst = 32'h8220000;
      7226: inst = 32'h10408000;
      7227: inst = 32'hc40520e;
      7228: inst = 32'h8220000;
      7229: inst = 32'h10408000;
      7230: inst = 32'hc40520f;
      7231: inst = 32'h8220000;
      7232: inst = 32'h10408000;
      7233: inst = 32'hc405210;
      7234: inst = 32'h8220000;
      7235: inst = 32'h10408000;
      7236: inst = 32'hc405211;
      7237: inst = 32'h8220000;
      7238: inst = 32'h10408000;
      7239: inst = 32'hc405212;
      7240: inst = 32'h8220000;
      7241: inst = 32'h10408000;
      7242: inst = 32'hc405213;
      7243: inst = 32'h8220000;
      7244: inst = 32'h10408000;
      7245: inst = 32'hc405214;
      7246: inst = 32'h8220000;
      7247: inst = 32'h10408000;
      7248: inst = 32'hc405215;
      7249: inst = 32'h8220000;
      7250: inst = 32'h10408000;
      7251: inst = 32'hc405223;
      7252: inst = 32'h8220000;
      7253: inst = 32'h10408000;
      7254: inst = 32'hc405224;
      7255: inst = 32'h8220000;
      7256: inst = 32'h10408000;
      7257: inst = 32'hc405225;
      7258: inst = 32'h8220000;
      7259: inst = 32'h10408000;
      7260: inst = 32'hc405226;
      7261: inst = 32'h8220000;
      7262: inst = 32'h10408000;
      7263: inst = 32'hc405227;
      7264: inst = 32'h8220000;
      7265: inst = 32'h10408000;
      7266: inst = 32'hc405228;
      7267: inst = 32'h8220000;
      7268: inst = 32'h10408000;
      7269: inst = 32'hc405229;
      7270: inst = 32'h8220000;
      7271: inst = 32'h10408000;
      7272: inst = 32'hc40522a;
      7273: inst = 32'h8220000;
      7274: inst = 32'h10408000;
      7275: inst = 32'hc40522b;
      7276: inst = 32'h8220000;
      7277: inst = 32'h10408000;
      7278: inst = 32'hc40522c;
      7279: inst = 32'h8220000;
      7280: inst = 32'h10408000;
      7281: inst = 32'hc40522d;
      7282: inst = 32'h8220000;
      7283: inst = 32'h10408000;
      7284: inst = 32'hc40522e;
      7285: inst = 32'h8220000;
      7286: inst = 32'h10408000;
      7287: inst = 32'hc405257;
      7288: inst = 32'h8220000;
      7289: inst = 32'h10408000;
      7290: inst = 32'hc405258;
      7291: inst = 32'h8220000;
      7292: inst = 32'h10408000;
      7293: inst = 32'hc405259;
      7294: inst = 32'h8220000;
      7295: inst = 32'h10408000;
      7296: inst = 32'hc40525a;
      7297: inst = 32'h8220000;
      7298: inst = 32'h10408000;
      7299: inst = 32'hc40525b;
      7300: inst = 32'h8220000;
      7301: inst = 32'h10408000;
      7302: inst = 32'hc40526a;
      7303: inst = 32'h8220000;
      7304: inst = 32'h10408000;
      7305: inst = 32'hc40526b;
      7306: inst = 32'h8220000;
      7307: inst = 32'h10408000;
      7308: inst = 32'hc40526c;
      7309: inst = 32'h8220000;
      7310: inst = 32'h10408000;
      7311: inst = 32'hc40526d;
      7312: inst = 32'h8220000;
      7313: inst = 32'h10408000;
      7314: inst = 32'hc40526e;
      7315: inst = 32'h8220000;
      7316: inst = 32'h10408000;
      7317: inst = 32'hc40526f;
      7318: inst = 32'h8220000;
      7319: inst = 32'h10408000;
      7320: inst = 32'hc405270;
      7321: inst = 32'h8220000;
      7322: inst = 32'h10408000;
      7323: inst = 32'hc405271;
      7324: inst = 32'h8220000;
      7325: inst = 32'h10408000;
      7326: inst = 32'hc405272;
      7327: inst = 32'h8220000;
      7328: inst = 32'h10408000;
      7329: inst = 32'hc405273;
      7330: inst = 32'h8220000;
      7331: inst = 32'h10408000;
      7332: inst = 32'hc405274;
      7333: inst = 32'h8220000;
      7334: inst = 32'h10408000;
      7335: inst = 32'hc405275;
      7336: inst = 32'h8220000;
      7337: inst = 32'h10408000;
      7338: inst = 32'hc405284;
      7339: inst = 32'h8220000;
      7340: inst = 32'h10408000;
      7341: inst = 32'hc405285;
      7342: inst = 32'h8220000;
      7343: inst = 32'h10408000;
      7344: inst = 32'hc405286;
      7345: inst = 32'h8220000;
      7346: inst = 32'h10408000;
      7347: inst = 32'hc405287;
      7348: inst = 32'h8220000;
      7349: inst = 32'h10408000;
      7350: inst = 32'hc405288;
      7351: inst = 32'h8220000;
      7352: inst = 32'h10408000;
      7353: inst = 32'hc405289;
      7354: inst = 32'h8220000;
      7355: inst = 32'h10408000;
      7356: inst = 32'hc40528a;
      7357: inst = 32'h8220000;
      7358: inst = 32'h10408000;
      7359: inst = 32'hc40528b;
      7360: inst = 32'h8220000;
      7361: inst = 32'h10408000;
      7362: inst = 32'hc40528c;
      7363: inst = 32'h8220000;
      7364: inst = 32'h10408000;
      7365: inst = 32'hc40528d;
      7366: inst = 32'h8220000;
      7367: inst = 32'h10408000;
      7368: inst = 32'hc40528e;
      7369: inst = 32'h8220000;
      7370: inst = 32'h10408000;
      7371: inst = 32'hc4052b7;
      7372: inst = 32'h8220000;
      7373: inst = 32'h10408000;
      7374: inst = 32'hc4052b8;
      7375: inst = 32'h8220000;
      7376: inst = 32'h10408000;
      7377: inst = 32'hc4052b9;
      7378: inst = 32'h8220000;
      7379: inst = 32'h10408000;
      7380: inst = 32'hc4052ba;
      7381: inst = 32'h8220000;
      7382: inst = 32'h10408000;
      7383: inst = 32'hc4052bb;
      7384: inst = 32'h8220000;
      7385: inst = 32'h10408000;
      7386: inst = 32'hc4052ca;
      7387: inst = 32'h8220000;
      7388: inst = 32'h10408000;
      7389: inst = 32'hc4052cb;
      7390: inst = 32'h8220000;
      7391: inst = 32'h10408000;
      7392: inst = 32'hc4052cc;
      7393: inst = 32'h8220000;
      7394: inst = 32'h10408000;
      7395: inst = 32'hc4052cd;
      7396: inst = 32'h8220000;
      7397: inst = 32'h10408000;
      7398: inst = 32'hc4052ce;
      7399: inst = 32'h8220000;
      7400: inst = 32'h10408000;
      7401: inst = 32'hc4052cf;
      7402: inst = 32'h8220000;
      7403: inst = 32'h10408000;
      7404: inst = 32'hc4052d0;
      7405: inst = 32'h8220000;
      7406: inst = 32'h10408000;
      7407: inst = 32'hc4052d1;
      7408: inst = 32'h8220000;
      7409: inst = 32'h10408000;
      7410: inst = 32'hc4052d2;
      7411: inst = 32'h8220000;
      7412: inst = 32'h10408000;
      7413: inst = 32'hc4052d3;
      7414: inst = 32'h8220000;
      7415: inst = 32'h10408000;
      7416: inst = 32'hc4052d4;
      7417: inst = 32'h8220000;
      7418: inst = 32'h10408000;
      7419: inst = 32'hc4052d5;
      7420: inst = 32'h8220000;
      7421: inst = 32'h10408000;
      7422: inst = 32'hc4052e4;
      7423: inst = 32'h8220000;
      7424: inst = 32'h10408000;
      7425: inst = 32'hc4052e5;
      7426: inst = 32'h8220000;
      7427: inst = 32'h10408000;
      7428: inst = 32'hc4052e6;
      7429: inst = 32'h8220000;
      7430: inst = 32'h10408000;
      7431: inst = 32'hc4052e7;
      7432: inst = 32'h8220000;
      7433: inst = 32'h10408000;
      7434: inst = 32'hc4052e8;
      7435: inst = 32'h8220000;
      7436: inst = 32'h10408000;
      7437: inst = 32'hc4052e9;
      7438: inst = 32'h8220000;
      7439: inst = 32'h10408000;
      7440: inst = 32'hc4052ea;
      7441: inst = 32'h8220000;
      7442: inst = 32'h10408000;
      7443: inst = 32'hc4052eb;
      7444: inst = 32'h8220000;
      7445: inst = 32'h10408000;
      7446: inst = 32'hc4052ec;
      7447: inst = 32'h8220000;
      7448: inst = 32'h10408000;
      7449: inst = 32'hc4052ed;
      7450: inst = 32'h8220000;
      7451: inst = 32'h10408000;
      7452: inst = 32'hc4052ee;
      7453: inst = 32'h8220000;
      7454: inst = 32'hc2094b2;
      7455: inst = 32'h10408000;
      7456: inst = 32'hc403feb;
      7457: inst = 32'h8220000;
      7458: inst = 32'h10408000;
      7459: inst = 32'hc40404b;
      7460: inst = 32'h8220000;
      7461: inst = 32'h10408000;
      7462: inst = 32'hc4040ab;
      7463: inst = 32'h8220000;
      7464: inst = 32'h10408000;
      7465: inst = 32'hc40410b;
      7466: inst = 32'h8220000;
      7467: inst = 32'h10408000;
      7468: inst = 32'hc40416b;
      7469: inst = 32'h8220000;
      7470: inst = 32'h10408000;
      7471: inst = 32'hc4041cb;
      7472: inst = 32'h8220000;
      7473: inst = 32'h10408000;
      7474: inst = 32'hc40422b;
      7475: inst = 32'h8220000;
      7476: inst = 32'h10408000;
      7477: inst = 32'hc40428b;
      7478: inst = 32'h8220000;
      7479: inst = 32'hc20b596;
      7480: inst = 32'h10408000;
      7481: inst = 32'hc4041da;
      7482: inst = 32'h8220000;
      7483: inst = 32'h10408000;
      7484: inst = 32'hc4041db;
      7485: inst = 32'h8220000;
      7486: inst = 32'h10408000;
      7487: inst = 32'hc4041dc;
      7488: inst = 32'h8220000;
      7489: inst = 32'h10408000;
      7490: inst = 32'hc4041dd;
      7491: inst = 32'h8220000;
      7492: inst = 32'h10408000;
      7493: inst = 32'hc4041de;
      7494: inst = 32'h8220000;
      7495: inst = 32'h10408000;
      7496: inst = 32'hc4041df;
      7497: inst = 32'h8220000;
      7498: inst = 32'h10408000;
      7499: inst = 32'hc4041e0;
      7500: inst = 32'h8220000;
      7501: inst = 32'h10408000;
      7502: inst = 32'hc4041e1;
      7503: inst = 32'h8220000;
      7504: inst = 32'h10408000;
      7505: inst = 32'hc4041e2;
      7506: inst = 32'h8220000;
      7507: inst = 32'h10408000;
      7508: inst = 32'hc4041e3;
      7509: inst = 32'h8220000;
      7510: inst = 32'h10408000;
      7511: inst = 32'hc4041e4;
      7512: inst = 32'h8220000;
      7513: inst = 32'h10408000;
      7514: inst = 32'hc4041e5;
      7515: inst = 32'h8220000;
      7516: inst = 32'h10408000;
      7517: inst = 32'hc4041e6;
      7518: inst = 32'h8220000;
      7519: inst = 32'h10408000;
      7520: inst = 32'hc4041e7;
      7521: inst = 32'h8220000;
      7522: inst = 32'h10408000;
      7523: inst = 32'hc4041e8;
      7524: inst = 32'h8220000;
      7525: inst = 32'h10408000;
      7526: inst = 32'hc4041e9;
      7527: inst = 32'h8220000;
      7528: inst = 32'h10408000;
      7529: inst = 32'hc4041ea;
      7530: inst = 32'h8220000;
      7531: inst = 32'h10408000;
      7532: inst = 32'hc4041eb;
      7533: inst = 32'h8220000;
      7534: inst = 32'h10408000;
      7535: inst = 32'hc4041ec;
      7536: inst = 32'h8220000;
      7537: inst = 32'h10408000;
      7538: inst = 32'hc4041ed;
      7539: inst = 32'h8220000;
      7540: inst = 32'h10408000;
      7541: inst = 32'hc4041ee;
      7542: inst = 32'h8220000;
      7543: inst = 32'h10408000;
      7544: inst = 32'hc4041ef;
      7545: inst = 32'h8220000;
      7546: inst = 32'h10408000;
      7547: inst = 32'hc4041f0;
      7548: inst = 32'h8220000;
      7549: inst = 32'h10408000;
      7550: inst = 32'hc4041f1;
      7551: inst = 32'h8220000;
      7552: inst = 32'h10408000;
      7553: inst = 32'hc4041f2;
      7554: inst = 32'h8220000;
      7555: inst = 32'h10408000;
      7556: inst = 32'hc4041f3;
      7557: inst = 32'h8220000;
      7558: inst = 32'h10408000;
      7559: inst = 32'hc4041f4;
      7560: inst = 32'h8220000;
      7561: inst = 32'h10408000;
      7562: inst = 32'hc4041f5;
      7563: inst = 32'h8220000;
      7564: inst = 32'h10408000;
      7565: inst = 32'hc4041f6;
      7566: inst = 32'h8220000;
      7567: inst = 32'h10408000;
      7568: inst = 32'hc4041f7;
      7569: inst = 32'h8220000;
      7570: inst = 32'h10408000;
      7571: inst = 32'hc4041f8;
      7572: inst = 32'h8220000;
      7573: inst = 32'h10408000;
      7574: inst = 32'hc4041f9;
      7575: inst = 32'h8220000;
      7576: inst = 32'h10408000;
      7577: inst = 32'hc4041fa;
      7578: inst = 32'h8220000;
      7579: inst = 32'h10408000;
      7580: inst = 32'hc4041fb;
      7581: inst = 32'h8220000;
      7582: inst = 32'h10408000;
      7583: inst = 32'hc4041fc;
      7584: inst = 32'h8220000;
      7585: inst = 32'h10408000;
      7586: inst = 32'hc4041fd;
      7587: inst = 32'h8220000;
      7588: inst = 32'h10408000;
      7589: inst = 32'hc4041fe;
      7590: inst = 32'h8220000;
      7591: inst = 32'h10408000;
      7592: inst = 32'hc4041ff;
      7593: inst = 32'h8220000;
      7594: inst = 32'h10408000;
      7595: inst = 32'hc404200;
      7596: inst = 32'h8220000;
      7597: inst = 32'h10408000;
      7598: inst = 32'hc404201;
      7599: inst = 32'h8220000;
      7600: inst = 32'h10408000;
      7601: inst = 32'hc404202;
      7602: inst = 32'h8220000;
      7603: inst = 32'h10408000;
      7604: inst = 32'hc404203;
      7605: inst = 32'h8220000;
      7606: inst = 32'h10408000;
      7607: inst = 32'hc404204;
      7608: inst = 32'h8220000;
      7609: inst = 32'h10408000;
      7610: inst = 32'hc404205;
      7611: inst = 32'h8220000;
      7612: inst = 32'h10408000;
      7613: inst = 32'hc404bfa;
      7614: inst = 32'h8220000;
      7615: inst = 32'h10408000;
      7616: inst = 32'hc404bfb;
      7617: inst = 32'h8220000;
      7618: inst = 32'h10408000;
      7619: inst = 32'hc404bfc;
      7620: inst = 32'h8220000;
      7621: inst = 32'h10408000;
      7622: inst = 32'hc404bfd;
      7623: inst = 32'h8220000;
      7624: inst = 32'h10408000;
      7625: inst = 32'hc404bfe;
      7626: inst = 32'h8220000;
      7627: inst = 32'h10408000;
      7628: inst = 32'hc404bff;
      7629: inst = 32'h8220000;
      7630: inst = 32'h10408000;
      7631: inst = 32'hc404c00;
      7632: inst = 32'h8220000;
      7633: inst = 32'h10408000;
      7634: inst = 32'hc404c01;
      7635: inst = 32'h8220000;
      7636: inst = 32'h10408000;
      7637: inst = 32'hc404c02;
      7638: inst = 32'h8220000;
      7639: inst = 32'h10408000;
      7640: inst = 32'hc404c03;
      7641: inst = 32'h8220000;
      7642: inst = 32'h10408000;
      7643: inst = 32'hc404c04;
      7644: inst = 32'h8220000;
      7645: inst = 32'h10408000;
      7646: inst = 32'hc404c05;
      7647: inst = 32'h8220000;
      7648: inst = 32'h10408000;
      7649: inst = 32'hc404c06;
      7650: inst = 32'h8220000;
      7651: inst = 32'h10408000;
      7652: inst = 32'hc404c07;
      7653: inst = 32'h8220000;
      7654: inst = 32'h10408000;
      7655: inst = 32'hc404c08;
      7656: inst = 32'h8220000;
      7657: inst = 32'h10408000;
      7658: inst = 32'hc404c09;
      7659: inst = 32'h8220000;
      7660: inst = 32'h10408000;
      7661: inst = 32'hc404c0a;
      7662: inst = 32'h8220000;
      7663: inst = 32'h10408000;
      7664: inst = 32'hc404c0b;
      7665: inst = 32'h8220000;
      7666: inst = 32'h10408000;
      7667: inst = 32'hc404c0c;
      7668: inst = 32'h8220000;
      7669: inst = 32'h10408000;
      7670: inst = 32'hc404c0d;
      7671: inst = 32'h8220000;
      7672: inst = 32'h10408000;
      7673: inst = 32'hc404c0e;
      7674: inst = 32'h8220000;
      7675: inst = 32'h10408000;
      7676: inst = 32'hc404c0f;
      7677: inst = 32'h8220000;
      7678: inst = 32'h10408000;
      7679: inst = 32'hc404c10;
      7680: inst = 32'h8220000;
      7681: inst = 32'h10408000;
      7682: inst = 32'hc404c11;
      7683: inst = 32'h8220000;
      7684: inst = 32'h10408000;
      7685: inst = 32'hc404c12;
      7686: inst = 32'h8220000;
      7687: inst = 32'h10408000;
      7688: inst = 32'hc404c13;
      7689: inst = 32'h8220000;
      7690: inst = 32'h10408000;
      7691: inst = 32'hc404c14;
      7692: inst = 32'h8220000;
      7693: inst = 32'h10408000;
      7694: inst = 32'hc404c15;
      7695: inst = 32'h8220000;
      7696: inst = 32'h10408000;
      7697: inst = 32'hc404c16;
      7698: inst = 32'h8220000;
      7699: inst = 32'h10408000;
      7700: inst = 32'hc404c17;
      7701: inst = 32'h8220000;
      7702: inst = 32'h10408000;
      7703: inst = 32'hc404c18;
      7704: inst = 32'h8220000;
      7705: inst = 32'h10408000;
      7706: inst = 32'hc404c19;
      7707: inst = 32'h8220000;
      7708: inst = 32'h10408000;
      7709: inst = 32'hc404c1a;
      7710: inst = 32'h8220000;
      7711: inst = 32'h10408000;
      7712: inst = 32'hc404c1b;
      7713: inst = 32'h8220000;
      7714: inst = 32'h10408000;
      7715: inst = 32'hc404c1c;
      7716: inst = 32'h8220000;
      7717: inst = 32'h10408000;
      7718: inst = 32'hc404c1d;
      7719: inst = 32'h8220000;
      7720: inst = 32'h10408000;
      7721: inst = 32'hc404c1e;
      7722: inst = 32'h8220000;
      7723: inst = 32'h10408000;
      7724: inst = 32'hc404c1f;
      7725: inst = 32'h8220000;
      7726: inst = 32'h10408000;
      7727: inst = 32'hc404c20;
      7728: inst = 32'h8220000;
      7729: inst = 32'h10408000;
      7730: inst = 32'hc404c21;
      7731: inst = 32'h8220000;
      7732: inst = 32'h10408000;
      7733: inst = 32'hc404c22;
      7734: inst = 32'h8220000;
      7735: inst = 32'h10408000;
      7736: inst = 32'hc404c23;
      7737: inst = 32'h8220000;
      7738: inst = 32'h10408000;
      7739: inst = 32'hc404c24;
      7740: inst = 32'h8220000;
      7741: inst = 32'h10408000;
      7742: inst = 32'hc404c25;
      7743: inst = 32'h8220000;
      7744: inst = 32'hc20ffff;
      7745: inst = 32'h10408000;
      7746: inst = 32'hc40423c;
      7747: inst = 32'h8220000;
      7748: inst = 32'h10408000;
      7749: inst = 32'hc40423d;
      7750: inst = 32'h8220000;
      7751: inst = 32'h10408000;
      7752: inst = 32'hc40423e;
      7753: inst = 32'h8220000;
      7754: inst = 32'h10408000;
      7755: inst = 32'hc40423f;
      7756: inst = 32'h8220000;
      7757: inst = 32'h10408000;
      7758: inst = 32'hc404240;
      7759: inst = 32'h8220000;
      7760: inst = 32'h10408000;
      7761: inst = 32'hc404241;
      7762: inst = 32'h8220000;
      7763: inst = 32'h10408000;
      7764: inst = 32'hc404242;
      7765: inst = 32'h8220000;
      7766: inst = 32'h10408000;
      7767: inst = 32'hc404243;
      7768: inst = 32'h8220000;
      7769: inst = 32'h10408000;
      7770: inst = 32'hc404244;
      7771: inst = 32'h8220000;
      7772: inst = 32'h10408000;
      7773: inst = 32'hc404245;
      7774: inst = 32'h8220000;
      7775: inst = 32'h10408000;
      7776: inst = 32'hc404246;
      7777: inst = 32'h8220000;
      7778: inst = 32'h10408000;
      7779: inst = 32'hc404247;
      7780: inst = 32'h8220000;
      7781: inst = 32'h10408000;
      7782: inst = 32'hc404248;
      7783: inst = 32'h8220000;
      7784: inst = 32'h10408000;
      7785: inst = 32'hc404249;
      7786: inst = 32'h8220000;
      7787: inst = 32'h10408000;
      7788: inst = 32'hc40424a;
      7789: inst = 32'h8220000;
      7790: inst = 32'h10408000;
      7791: inst = 32'hc40424b;
      7792: inst = 32'h8220000;
      7793: inst = 32'h10408000;
      7794: inst = 32'hc40424c;
      7795: inst = 32'h8220000;
      7796: inst = 32'h10408000;
      7797: inst = 32'hc40424d;
      7798: inst = 32'h8220000;
      7799: inst = 32'h10408000;
      7800: inst = 32'hc40424e;
      7801: inst = 32'h8220000;
      7802: inst = 32'h10408000;
      7803: inst = 32'hc40424f;
      7804: inst = 32'h8220000;
      7805: inst = 32'h10408000;
      7806: inst = 32'hc404250;
      7807: inst = 32'h8220000;
      7808: inst = 32'h10408000;
      7809: inst = 32'hc404251;
      7810: inst = 32'h8220000;
      7811: inst = 32'h10408000;
      7812: inst = 32'hc404252;
      7813: inst = 32'h8220000;
      7814: inst = 32'h10408000;
      7815: inst = 32'hc404253;
      7816: inst = 32'h8220000;
      7817: inst = 32'h10408000;
      7818: inst = 32'hc404254;
      7819: inst = 32'h8220000;
      7820: inst = 32'h10408000;
      7821: inst = 32'hc404255;
      7822: inst = 32'h8220000;
      7823: inst = 32'h10408000;
      7824: inst = 32'hc404256;
      7825: inst = 32'h8220000;
      7826: inst = 32'h10408000;
      7827: inst = 32'hc404257;
      7828: inst = 32'h8220000;
      7829: inst = 32'h10408000;
      7830: inst = 32'hc404258;
      7831: inst = 32'h8220000;
      7832: inst = 32'h10408000;
      7833: inst = 32'hc404259;
      7834: inst = 32'h8220000;
      7835: inst = 32'h10408000;
      7836: inst = 32'hc40425a;
      7837: inst = 32'h8220000;
      7838: inst = 32'h10408000;
      7839: inst = 32'hc40425b;
      7840: inst = 32'h8220000;
      7841: inst = 32'h10408000;
      7842: inst = 32'hc40425c;
      7843: inst = 32'h8220000;
      7844: inst = 32'h10408000;
      7845: inst = 32'hc40425d;
      7846: inst = 32'h8220000;
      7847: inst = 32'h10408000;
      7848: inst = 32'hc40425e;
      7849: inst = 32'h8220000;
      7850: inst = 32'h10408000;
      7851: inst = 32'hc40425f;
      7852: inst = 32'h8220000;
      7853: inst = 32'h10408000;
      7854: inst = 32'hc404260;
      7855: inst = 32'h8220000;
      7856: inst = 32'h10408000;
      7857: inst = 32'hc404261;
      7858: inst = 32'h8220000;
      7859: inst = 32'h10408000;
      7860: inst = 32'hc404262;
      7861: inst = 32'h8220000;
      7862: inst = 32'h10408000;
      7863: inst = 32'hc404263;
      7864: inst = 32'h8220000;
      7865: inst = 32'h10408000;
      7866: inst = 32'hc40429c;
      7867: inst = 32'h8220000;
      7868: inst = 32'h10408000;
      7869: inst = 32'hc40429d;
      7870: inst = 32'h8220000;
      7871: inst = 32'h10408000;
      7872: inst = 32'hc40429e;
      7873: inst = 32'h8220000;
      7874: inst = 32'h10408000;
      7875: inst = 32'hc40429f;
      7876: inst = 32'h8220000;
      7877: inst = 32'h10408000;
      7878: inst = 32'hc4042a0;
      7879: inst = 32'h8220000;
      7880: inst = 32'h10408000;
      7881: inst = 32'hc4042a1;
      7882: inst = 32'h8220000;
      7883: inst = 32'h10408000;
      7884: inst = 32'hc4042a2;
      7885: inst = 32'h8220000;
      7886: inst = 32'h10408000;
      7887: inst = 32'hc4042a3;
      7888: inst = 32'h8220000;
      7889: inst = 32'h10408000;
      7890: inst = 32'hc4042a4;
      7891: inst = 32'h8220000;
      7892: inst = 32'h10408000;
      7893: inst = 32'hc4042a5;
      7894: inst = 32'h8220000;
      7895: inst = 32'h10408000;
      7896: inst = 32'hc4042a6;
      7897: inst = 32'h8220000;
      7898: inst = 32'h10408000;
      7899: inst = 32'hc4042a7;
      7900: inst = 32'h8220000;
      7901: inst = 32'h10408000;
      7902: inst = 32'hc4042a8;
      7903: inst = 32'h8220000;
      7904: inst = 32'h10408000;
      7905: inst = 32'hc4042a9;
      7906: inst = 32'h8220000;
      7907: inst = 32'h10408000;
      7908: inst = 32'hc4042aa;
      7909: inst = 32'h8220000;
      7910: inst = 32'h10408000;
      7911: inst = 32'hc4042ab;
      7912: inst = 32'h8220000;
      7913: inst = 32'h10408000;
      7914: inst = 32'hc4042ac;
      7915: inst = 32'h8220000;
      7916: inst = 32'h10408000;
      7917: inst = 32'hc4042ad;
      7918: inst = 32'h8220000;
      7919: inst = 32'h10408000;
      7920: inst = 32'hc4042ae;
      7921: inst = 32'h8220000;
      7922: inst = 32'h10408000;
      7923: inst = 32'hc4042af;
      7924: inst = 32'h8220000;
      7925: inst = 32'h10408000;
      7926: inst = 32'hc4042b0;
      7927: inst = 32'h8220000;
      7928: inst = 32'h10408000;
      7929: inst = 32'hc4042b1;
      7930: inst = 32'h8220000;
      7931: inst = 32'h10408000;
      7932: inst = 32'hc4042b2;
      7933: inst = 32'h8220000;
      7934: inst = 32'h10408000;
      7935: inst = 32'hc4042b3;
      7936: inst = 32'h8220000;
      7937: inst = 32'h10408000;
      7938: inst = 32'hc4042b4;
      7939: inst = 32'h8220000;
      7940: inst = 32'h10408000;
      7941: inst = 32'hc4042b5;
      7942: inst = 32'h8220000;
      7943: inst = 32'h10408000;
      7944: inst = 32'hc4042b6;
      7945: inst = 32'h8220000;
      7946: inst = 32'h10408000;
      7947: inst = 32'hc4042b7;
      7948: inst = 32'h8220000;
      7949: inst = 32'h10408000;
      7950: inst = 32'hc4042b8;
      7951: inst = 32'h8220000;
      7952: inst = 32'h10408000;
      7953: inst = 32'hc4042b9;
      7954: inst = 32'h8220000;
      7955: inst = 32'h10408000;
      7956: inst = 32'hc4042ba;
      7957: inst = 32'h8220000;
      7958: inst = 32'h10408000;
      7959: inst = 32'hc4042bb;
      7960: inst = 32'h8220000;
      7961: inst = 32'h10408000;
      7962: inst = 32'hc4042bc;
      7963: inst = 32'h8220000;
      7964: inst = 32'h10408000;
      7965: inst = 32'hc4042bd;
      7966: inst = 32'h8220000;
      7967: inst = 32'h10408000;
      7968: inst = 32'hc4042be;
      7969: inst = 32'h8220000;
      7970: inst = 32'h10408000;
      7971: inst = 32'hc4042bf;
      7972: inst = 32'h8220000;
      7973: inst = 32'h10408000;
      7974: inst = 32'hc4042c0;
      7975: inst = 32'h8220000;
      7976: inst = 32'h10408000;
      7977: inst = 32'hc4042c1;
      7978: inst = 32'h8220000;
      7979: inst = 32'h10408000;
      7980: inst = 32'hc4042c2;
      7981: inst = 32'h8220000;
      7982: inst = 32'h10408000;
      7983: inst = 32'hc4042c3;
      7984: inst = 32'h8220000;
      7985: inst = 32'h10408000;
      7986: inst = 32'hc4042fc;
      7987: inst = 32'h8220000;
      7988: inst = 32'h10408000;
      7989: inst = 32'hc4042fd;
      7990: inst = 32'h8220000;
      7991: inst = 32'h10408000;
      7992: inst = 32'hc4042fe;
      7993: inst = 32'h8220000;
      7994: inst = 32'h10408000;
      7995: inst = 32'hc4042ff;
      7996: inst = 32'h8220000;
      7997: inst = 32'h10408000;
      7998: inst = 32'hc404300;
      7999: inst = 32'h8220000;
      8000: inst = 32'h10408000;
      8001: inst = 32'hc404301;
      8002: inst = 32'h8220000;
      8003: inst = 32'h10408000;
      8004: inst = 32'hc404302;
      8005: inst = 32'h8220000;
      8006: inst = 32'h10408000;
      8007: inst = 32'hc404303;
      8008: inst = 32'h8220000;
      8009: inst = 32'h10408000;
      8010: inst = 32'hc404304;
      8011: inst = 32'h8220000;
      8012: inst = 32'h10408000;
      8013: inst = 32'hc404305;
      8014: inst = 32'h8220000;
      8015: inst = 32'h10408000;
      8016: inst = 32'hc404306;
      8017: inst = 32'h8220000;
      8018: inst = 32'h10408000;
      8019: inst = 32'hc404307;
      8020: inst = 32'h8220000;
      8021: inst = 32'h10408000;
      8022: inst = 32'hc404308;
      8023: inst = 32'h8220000;
      8024: inst = 32'h10408000;
      8025: inst = 32'hc404309;
      8026: inst = 32'h8220000;
      8027: inst = 32'h10408000;
      8028: inst = 32'hc40430a;
      8029: inst = 32'h8220000;
      8030: inst = 32'h10408000;
      8031: inst = 32'hc40430b;
      8032: inst = 32'h8220000;
      8033: inst = 32'h10408000;
      8034: inst = 32'hc40430c;
      8035: inst = 32'h8220000;
      8036: inst = 32'h10408000;
      8037: inst = 32'hc40430d;
      8038: inst = 32'h8220000;
      8039: inst = 32'h10408000;
      8040: inst = 32'hc40430e;
      8041: inst = 32'h8220000;
      8042: inst = 32'h10408000;
      8043: inst = 32'hc40430f;
      8044: inst = 32'h8220000;
      8045: inst = 32'h10408000;
      8046: inst = 32'hc404310;
      8047: inst = 32'h8220000;
      8048: inst = 32'h10408000;
      8049: inst = 32'hc404311;
      8050: inst = 32'h8220000;
      8051: inst = 32'h10408000;
      8052: inst = 32'hc404312;
      8053: inst = 32'h8220000;
      8054: inst = 32'h10408000;
      8055: inst = 32'hc404313;
      8056: inst = 32'h8220000;
      8057: inst = 32'h10408000;
      8058: inst = 32'hc404314;
      8059: inst = 32'h8220000;
      8060: inst = 32'h10408000;
      8061: inst = 32'hc404315;
      8062: inst = 32'h8220000;
      8063: inst = 32'h10408000;
      8064: inst = 32'hc404316;
      8065: inst = 32'h8220000;
      8066: inst = 32'h10408000;
      8067: inst = 32'hc404317;
      8068: inst = 32'h8220000;
      8069: inst = 32'h10408000;
      8070: inst = 32'hc404318;
      8071: inst = 32'h8220000;
      8072: inst = 32'h10408000;
      8073: inst = 32'hc404319;
      8074: inst = 32'h8220000;
      8075: inst = 32'h10408000;
      8076: inst = 32'hc40431a;
      8077: inst = 32'h8220000;
      8078: inst = 32'h10408000;
      8079: inst = 32'hc40431b;
      8080: inst = 32'h8220000;
      8081: inst = 32'h10408000;
      8082: inst = 32'hc40431c;
      8083: inst = 32'h8220000;
      8084: inst = 32'h10408000;
      8085: inst = 32'hc40431d;
      8086: inst = 32'h8220000;
      8087: inst = 32'h10408000;
      8088: inst = 32'hc40431e;
      8089: inst = 32'h8220000;
      8090: inst = 32'h10408000;
      8091: inst = 32'hc40431f;
      8092: inst = 32'h8220000;
      8093: inst = 32'h10408000;
      8094: inst = 32'hc404320;
      8095: inst = 32'h8220000;
      8096: inst = 32'h10408000;
      8097: inst = 32'hc404321;
      8098: inst = 32'h8220000;
      8099: inst = 32'h10408000;
      8100: inst = 32'hc404322;
      8101: inst = 32'h8220000;
      8102: inst = 32'h10408000;
      8103: inst = 32'hc404323;
      8104: inst = 32'h8220000;
      8105: inst = 32'h10408000;
      8106: inst = 32'hc40435c;
      8107: inst = 32'h8220000;
      8108: inst = 32'h10408000;
      8109: inst = 32'hc40435d;
      8110: inst = 32'h8220000;
      8111: inst = 32'h10408000;
      8112: inst = 32'hc40435e;
      8113: inst = 32'h8220000;
      8114: inst = 32'h10408000;
      8115: inst = 32'hc40435f;
      8116: inst = 32'h8220000;
      8117: inst = 32'h10408000;
      8118: inst = 32'hc404360;
      8119: inst = 32'h8220000;
      8120: inst = 32'h10408000;
      8121: inst = 32'hc404361;
      8122: inst = 32'h8220000;
      8123: inst = 32'h10408000;
      8124: inst = 32'hc404362;
      8125: inst = 32'h8220000;
      8126: inst = 32'h10408000;
      8127: inst = 32'hc404363;
      8128: inst = 32'h8220000;
      8129: inst = 32'h10408000;
      8130: inst = 32'hc404364;
      8131: inst = 32'h8220000;
      8132: inst = 32'h10408000;
      8133: inst = 32'hc404365;
      8134: inst = 32'h8220000;
      8135: inst = 32'h10408000;
      8136: inst = 32'hc404366;
      8137: inst = 32'h8220000;
      8138: inst = 32'h10408000;
      8139: inst = 32'hc404367;
      8140: inst = 32'h8220000;
      8141: inst = 32'h10408000;
      8142: inst = 32'hc404368;
      8143: inst = 32'h8220000;
      8144: inst = 32'h10408000;
      8145: inst = 32'hc404369;
      8146: inst = 32'h8220000;
      8147: inst = 32'h10408000;
      8148: inst = 32'hc40436a;
      8149: inst = 32'h8220000;
      8150: inst = 32'h10408000;
      8151: inst = 32'hc40436b;
      8152: inst = 32'h8220000;
      8153: inst = 32'h10408000;
      8154: inst = 32'hc40436c;
      8155: inst = 32'h8220000;
      8156: inst = 32'h10408000;
      8157: inst = 32'hc40436d;
      8158: inst = 32'h8220000;
      8159: inst = 32'h10408000;
      8160: inst = 32'hc40436e;
      8161: inst = 32'h8220000;
      8162: inst = 32'h10408000;
      8163: inst = 32'hc40436f;
      8164: inst = 32'h8220000;
      8165: inst = 32'h10408000;
      8166: inst = 32'hc404370;
      8167: inst = 32'h8220000;
      8168: inst = 32'h10408000;
      8169: inst = 32'hc404371;
      8170: inst = 32'h8220000;
      8171: inst = 32'h10408000;
      8172: inst = 32'hc404372;
      8173: inst = 32'h8220000;
      8174: inst = 32'h10408000;
      8175: inst = 32'hc404373;
      8176: inst = 32'h8220000;
      8177: inst = 32'h10408000;
      8178: inst = 32'hc404374;
      8179: inst = 32'h8220000;
      8180: inst = 32'h10408000;
      8181: inst = 32'hc404375;
      8182: inst = 32'h8220000;
      8183: inst = 32'h10408000;
      8184: inst = 32'hc404376;
      8185: inst = 32'h8220000;
      8186: inst = 32'h10408000;
      8187: inst = 32'hc404377;
      8188: inst = 32'h8220000;
      8189: inst = 32'h10408000;
      8190: inst = 32'hc404378;
      8191: inst = 32'h8220000;
      8192: inst = 32'h10408000;
      8193: inst = 32'hc404379;
      8194: inst = 32'h8220000;
      8195: inst = 32'h10408000;
      8196: inst = 32'hc40437a;
      8197: inst = 32'h8220000;
      8198: inst = 32'h10408000;
      8199: inst = 32'hc40437b;
      8200: inst = 32'h8220000;
      8201: inst = 32'h10408000;
      8202: inst = 32'hc40437c;
      8203: inst = 32'h8220000;
      8204: inst = 32'h10408000;
      8205: inst = 32'hc40437d;
      8206: inst = 32'h8220000;
      8207: inst = 32'h10408000;
      8208: inst = 32'hc40437e;
      8209: inst = 32'h8220000;
      8210: inst = 32'h10408000;
      8211: inst = 32'hc40437f;
      8212: inst = 32'h8220000;
      8213: inst = 32'h10408000;
      8214: inst = 32'hc404380;
      8215: inst = 32'h8220000;
      8216: inst = 32'h10408000;
      8217: inst = 32'hc404381;
      8218: inst = 32'h8220000;
      8219: inst = 32'h10408000;
      8220: inst = 32'hc404382;
      8221: inst = 32'h8220000;
      8222: inst = 32'h10408000;
      8223: inst = 32'hc404383;
      8224: inst = 32'h8220000;
      8225: inst = 32'h10408000;
      8226: inst = 32'hc4043bc;
      8227: inst = 32'h8220000;
      8228: inst = 32'h10408000;
      8229: inst = 32'hc4043bd;
      8230: inst = 32'h8220000;
      8231: inst = 32'h10408000;
      8232: inst = 32'hc4043be;
      8233: inst = 32'h8220000;
      8234: inst = 32'h10408000;
      8235: inst = 32'hc4043bf;
      8236: inst = 32'h8220000;
      8237: inst = 32'h10408000;
      8238: inst = 32'hc4043c0;
      8239: inst = 32'h8220000;
      8240: inst = 32'h10408000;
      8241: inst = 32'hc4043c1;
      8242: inst = 32'h8220000;
      8243: inst = 32'h10408000;
      8244: inst = 32'hc4043c2;
      8245: inst = 32'h8220000;
      8246: inst = 32'h10408000;
      8247: inst = 32'hc4043c3;
      8248: inst = 32'h8220000;
      8249: inst = 32'h10408000;
      8250: inst = 32'hc4043c4;
      8251: inst = 32'h8220000;
      8252: inst = 32'h10408000;
      8253: inst = 32'hc4043c5;
      8254: inst = 32'h8220000;
      8255: inst = 32'h10408000;
      8256: inst = 32'hc4043c6;
      8257: inst = 32'h8220000;
      8258: inst = 32'h10408000;
      8259: inst = 32'hc4043c7;
      8260: inst = 32'h8220000;
      8261: inst = 32'h10408000;
      8262: inst = 32'hc4043c8;
      8263: inst = 32'h8220000;
      8264: inst = 32'h10408000;
      8265: inst = 32'hc4043c9;
      8266: inst = 32'h8220000;
      8267: inst = 32'h10408000;
      8268: inst = 32'hc4043ca;
      8269: inst = 32'h8220000;
      8270: inst = 32'h10408000;
      8271: inst = 32'hc4043cb;
      8272: inst = 32'h8220000;
      8273: inst = 32'h10408000;
      8274: inst = 32'hc4043cc;
      8275: inst = 32'h8220000;
      8276: inst = 32'h10408000;
      8277: inst = 32'hc4043cd;
      8278: inst = 32'h8220000;
      8279: inst = 32'h10408000;
      8280: inst = 32'hc4043ce;
      8281: inst = 32'h8220000;
      8282: inst = 32'h10408000;
      8283: inst = 32'hc4043cf;
      8284: inst = 32'h8220000;
      8285: inst = 32'h10408000;
      8286: inst = 32'hc4043d0;
      8287: inst = 32'h8220000;
      8288: inst = 32'h10408000;
      8289: inst = 32'hc4043d1;
      8290: inst = 32'h8220000;
      8291: inst = 32'h10408000;
      8292: inst = 32'hc4043d2;
      8293: inst = 32'h8220000;
      8294: inst = 32'h10408000;
      8295: inst = 32'hc4043d3;
      8296: inst = 32'h8220000;
      8297: inst = 32'h10408000;
      8298: inst = 32'hc4043d4;
      8299: inst = 32'h8220000;
      8300: inst = 32'h10408000;
      8301: inst = 32'hc4043d5;
      8302: inst = 32'h8220000;
      8303: inst = 32'h10408000;
      8304: inst = 32'hc4043d6;
      8305: inst = 32'h8220000;
      8306: inst = 32'h10408000;
      8307: inst = 32'hc4043d7;
      8308: inst = 32'h8220000;
      8309: inst = 32'h10408000;
      8310: inst = 32'hc4043d8;
      8311: inst = 32'h8220000;
      8312: inst = 32'h10408000;
      8313: inst = 32'hc4043d9;
      8314: inst = 32'h8220000;
      8315: inst = 32'h10408000;
      8316: inst = 32'hc4043da;
      8317: inst = 32'h8220000;
      8318: inst = 32'h10408000;
      8319: inst = 32'hc4043db;
      8320: inst = 32'h8220000;
      8321: inst = 32'h10408000;
      8322: inst = 32'hc4043dc;
      8323: inst = 32'h8220000;
      8324: inst = 32'h10408000;
      8325: inst = 32'hc4043dd;
      8326: inst = 32'h8220000;
      8327: inst = 32'h10408000;
      8328: inst = 32'hc4043de;
      8329: inst = 32'h8220000;
      8330: inst = 32'h10408000;
      8331: inst = 32'hc4043df;
      8332: inst = 32'h8220000;
      8333: inst = 32'h10408000;
      8334: inst = 32'hc4043e0;
      8335: inst = 32'h8220000;
      8336: inst = 32'h10408000;
      8337: inst = 32'hc4043e1;
      8338: inst = 32'h8220000;
      8339: inst = 32'h10408000;
      8340: inst = 32'hc4043e2;
      8341: inst = 32'h8220000;
      8342: inst = 32'h10408000;
      8343: inst = 32'hc4043e3;
      8344: inst = 32'h8220000;
      8345: inst = 32'h10408000;
      8346: inst = 32'hc40441c;
      8347: inst = 32'h8220000;
      8348: inst = 32'h10408000;
      8349: inst = 32'hc40441d;
      8350: inst = 32'h8220000;
      8351: inst = 32'h10408000;
      8352: inst = 32'hc40441e;
      8353: inst = 32'h8220000;
      8354: inst = 32'h10408000;
      8355: inst = 32'hc40441f;
      8356: inst = 32'h8220000;
      8357: inst = 32'h10408000;
      8358: inst = 32'hc404420;
      8359: inst = 32'h8220000;
      8360: inst = 32'h10408000;
      8361: inst = 32'hc404421;
      8362: inst = 32'h8220000;
      8363: inst = 32'h10408000;
      8364: inst = 32'hc404422;
      8365: inst = 32'h8220000;
      8366: inst = 32'h10408000;
      8367: inst = 32'hc404423;
      8368: inst = 32'h8220000;
      8369: inst = 32'h10408000;
      8370: inst = 32'hc404424;
      8371: inst = 32'h8220000;
      8372: inst = 32'h10408000;
      8373: inst = 32'hc404425;
      8374: inst = 32'h8220000;
      8375: inst = 32'h10408000;
      8376: inst = 32'hc404426;
      8377: inst = 32'h8220000;
      8378: inst = 32'h10408000;
      8379: inst = 32'hc404427;
      8380: inst = 32'h8220000;
      8381: inst = 32'h10408000;
      8382: inst = 32'hc404428;
      8383: inst = 32'h8220000;
      8384: inst = 32'h10408000;
      8385: inst = 32'hc404429;
      8386: inst = 32'h8220000;
      8387: inst = 32'h10408000;
      8388: inst = 32'hc40442a;
      8389: inst = 32'h8220000;
      8390: inst = 32'h10408000;
      8391: inst = 32'hc40442b;
      8392: inst = 32'h8220000;
      8393: inst = 32'h10408000;
      8394: inst = 32'hc40442c;
      8395: inst = 32'h8220000;
      8396: inst = 32'h10408000;
      8397: inst = 32'hc40442d;
      8398: inst = 32'h8220000;
      8399: inst = 32'h10408000;
      8400: inst = 32'hc40442e;
      8401: inst = 32'h8220000;
      8402: inst = 32'h10408000;
      8403: inst = 32'hc40442f;
      8404: inst = 32'h8220000;
      8405: inst = 32'h10408000;
      8406: inst = 32'hc404430;
      8407: inst = 32'h8220000;
      8408: inst = 32'h10408000;
      8409: inst = 32'hc404431;
      8410: inst = 32'h8220000;
      8411: inst = 32'h10408000;
      8412: inst = 32'hc404432;
      8413: inst = 32'h8220000;
      8414: inst = 32'h10408000;
      8415: inst = 32'hc404433;
      8416: inst = 32'h8220000;
      8417: inst = 32'h10408000;
      8418: inst = 32'hc404434;
      8419: inst = 32'h8220000;
      8420: inst = 32'h10408000;
      8421: inst = 32'hc404435;
      8422: inst = 32'h8220000;
      8423: inst = 32'h10408000;
      8424: inst = 32'hc404436;
      8425: inst = 32'h8220000;
      8426: inst = 32'h10408000;
      8427: inst = 32'hc404437;
      8428: inst = 32'h8220000;
      8429: inst = 32'h10408000;
      8430: inst = 32'hc404438;
      8431: inst = 32'h8220000;
      8432: inst = 32'h10408000;
      8433: inst = 32'hc404439;
      8434: inst = 32'h8220000;
      8435: inst = 32'h10408000;
      8436: inst = 32'hc40443a;
      8437: inst = 32'h8220000;
      8438: inst = 32'h10408000;
      8439: inst = 32'hc40443b;
      8440: inst = 32'h8220000;
      8441: inst = 32'h10408000;
      8442: inst = 32'hc40443c;
      8443: inst = 32'h8220000;
      8444: inst = 32'h10408000;
      8445: inst = 32'hc40443d;
      8446: inst = 32'h8220000;
      8447: inst = 32'h10408000;
      8448: inst = 32'hc40443e;
      8449: inst = 32'h8220000;
      8450: inst = 32'h10408000;
      8451: inst = 32'hc40443f;
      8452: inst = 32'h8220000;
      8453: inst = 32'h10408000;
      8454: inst = 32'hc404440;
      8455: inst = 32'h8220000;
      8456: inst = 32'h10408000;
      8457: inst = 32'hc404441;
      8458: inst = 32'h8220000;
      8459: inst = 32'h10408000;
      8460: inst = 32'hc404442;
      8461: inst = 32'h8220000;
      8462: inst = 32'h10408000;
      8463: inst = 32'hc404443;
      8464: inst = 32'h8220000;
      8465: inst = 32'h10408000;
      8466: inst = 32'hc40447c;
      8467: inst = 32'h8220000;
      8468: inst = 32'h10408000;
      8469: inst = 32'hc40447d;
      8470: inst = 32'h8220000;
      8471: inst = 32'h10408000;
      8472: inst = 32'hc40447e;
      8473: inst = 32'h8220000;
      8474: inst = 32'h10408000;
      8475: inst = 32'hc40447f;
      8476: inst = 32'h8220000;
      8477: inst = 32'h10408000;
      8478: inst = 32'hc404480;
      8479: inst = 32'h8220000;
      8480: inst = 32'h10408000;
      8481: inst = 32'hc404481;
      8482: inst = 32'h8220000;
      8483: inst = 32'h10408000;
      8484: inst = 32'hc404482;
      8485: inst = 32'h8220000;
      8486: inst = 32'h10408000;
      8487: inst = 32'hc404483;
      8488: inst = 32'h8220000;
      8489: inst = 32'h10408000;
      8490: inst = 32'hc404484;
      8491: inst = 32'h8220000;
      8492: inst = 32'h10408000;
      8493: inst = 32'hc404485;
      8494: inst = 32'h8220000;
      8495: inst = 32'h10408000;
      8496: inst = 32'hc404486;
      8497: inst = 32'h8220000;
      8498: inst = 32'h10408000;
      8499: inst = 32'hc404487;
      8500: inst = 32'h8220000;
      8501: inst = 32'h10408000;
      8502: inst = 32'hc404488;
      8503: inst = 32'h8220000;
      8504: inst = 32'h10408000;
      8505: inst = 32'hc404489;
      8506: inst = 32'h8220000;
      8507: inst = 32'h10408000;
      8508: inst = 32'hc40448a;
      8509: inst = 32'h8220000;
      8510: inst = 32'h10408000;
      8511: inst = 32'hc40448b;
      8512: inst = 32'h8220000;
      8513: inst = 32'h10408000;
      8514: inst = 32'hc40448c;
      8515: inst = 32'h8220000;
      8516: inst = 32'h10408000;
      8517: inst = 32'hc40448d;
      8518: inst = 32'h8220000;
      8519: inst = 32'h10408000;
      8520: inst = 32'hc40448e;
      8521: inst = 32'h8220000;
      8522: inst = 32'h10408000;
      8523: inst = 32'hc40448f;
      8524: inst = 32'h8220000;
      8525: inst = 32'h10408000;
      8526: inst = 32'hc404490;
      8527: inst = 32'h8220000;
      8528: inst = 32'h10408000;
      8529: inst = 32'hc404491;
      8530: inst = 32'h8220000;
      8531: inst = 32'h10408000;
      8532: inst = 32'hc404492;
      8533: inst = 32'h8220000;
      8534: inst = 32'h10408000;
      8535: inst = 32'hc404493;
      8536: inst = 32'h8220000;
      8537: inst = 32'h10408000;
      8538: inst = 32'hc404494;
      8539: inst = 32'h8220000;
      8540: inst = 32'h10408000;
      8541: inst = 32'hc404495;
      8542: inst = 32'h8220000;
      8543: inst = 32'h10408000;
      8544: inst = 32'hc404496;
      8545: inst = 32'h8220000;
      8546: inst = 32'h10408000;
      8547: inst = 32'hc404497;
      8548: inst = 32'h8220000;
      8549: inst = 32'h10408000;
      8550: inst = 32'hc404498;
      8551: inst = 32'h8220000;
      8552: inst = 32'h10408000;
      8553: inst = 32'hc404499;
      8554: inst = 32'h8220000;
      8555: inst = 32'h10408000;
      8556: inst = 32'hc40449a;
      8557: inst = 32'h8220000;
      8558: inst = 32'h10408000;
      8559: inst = 32'hc40449b;
      8560: inst = 32'h8220000;
      8561: inst = 32'h10408000;
      8562: inst = 32'hc40449c;
      8563: inst = 32'h8220000;
      8564: inst = 32'h10408000;
      8565: inst = 32'hc40449d;
      8566: inst = 32'h8220000;
      8567: inst = 32'h10408000;
      8568: inst = 32'hc40449e;
      8569: inst = 32'h8220000;
      8570: inst = 32'h10408000;
      8571: inst = 32'hc40449f;
      8572: inst = 32'h8220000;
      8573: inst = 32'h10408000;
      8574: inst = 32'hc4044a0;
      8575: inst = 32'h8220000;
      8576: inst = 32'h10408000;
      8577: inst = 32'hc4044a1;
      8578: inst = 32'h8220000;
      8579: inst = 32'h10408000;
      8580: inst = 32'hc4044a2;
      8581: inst = 32'h8220000;
      8582: inst = 32'h10408000;
      8583: inst = 32'hc4044a3;
      8584: inst = 32'h8220000;
      8585: inst = 32'h10408000;
      8586: inst = 32'hc4044dc;
      8587: inst = 32'h8220000;
      8588: inst = 32'h10408000;
      8589: inst = 32'hc4044dd;
      8590: inst = 32'h8220000;
      8591: inst = 32'h10408000;
      8592: inst = 32'hc4044de;
      8593: inst = 32'h8220000;
      8594: inst = 32'h10408000;
      8595: inst = 32'hc4044df;
      8596: inst = 32'h8220000;
      8597: inst = 32'h10408000;
      8598: inst = 32'hc4044e0;
      8599: inst = 32'h8220000;
      8600: inst = 32'h10408000;
      8601: inst = 32'hc4044e1;
      8602: inst = 32'h8220000;
      8603: inst = 32'h10408000;
      8604: inst = 32'hc4044e2;
      8605: inst = 32'h8220000;
      8606: inst = 32'h10408000;
      8607: inst = 32'hc4044e3;
      8608: inst = 32'h8220000;
      8609: inst = 32'h10408000;
      8610: inst = 32'hc4044e4;
      8611: inst = 32'h8220000;
      8612: inst = 32'h10408000;
      8613: inst = 32'hc4044e5;
      8614: inst = 32'h8220000;
      8615: inst = 32'h10408000;
      8616: inst = 32'hc4044e6;
      8617: inst = 32'h8220000;
      8618: inst = 32'h10408000;
      8619: inst = 32'hc4044e7;
      8620: inst = 32'h8220000;
      8621: inst = 32'h10408000;
      8622: inst = 32'hc4044e8;
      8623: inst = 32'h8220000;
      8624: inst = 32'h10408000;
      8625: inst = 32'hc4044e9;
      8626: inst = 32'h8220000;
      8627: inst = 32'h10408000;
      8628: inst = 32'hc4044ea;
      8629: inst = 32'h8220000;
      8630: inst = 32'h10408000;
      8631: inst = 32'hc4044eb;
      8632: inst = 32'h8220000;
      8633: inst = 32'h10408000;
      8634: inst = 32'hc4044ec;
      8635: inst = 32'h8220000;
      8636: inst = 32'h10408000;
      8637: inst = 32'hc4044ed;
      8638: inst = 32'h8220000;
      8639: inst = 32'h10408000;
      8640: inst = 32'hc4044ee;
      8641: inst = 32'h8220000;
      8642: inst = 32'h10408000;
      8643: inst = 32'hc4044ef;
      8644: inst = 32'h8220000;
      8645: inst = 32'h10408000;
      8646: inst = 32'hc4044f0;
      8647: inst = 32'h8220000;
      8648: inst = 32'h10408000;
      8649: inst = 32'hc4044f1;
      8650: inst = 32'h8220000;
      8651: inst = 32'h10408000;
      8652: inst = 32'hc4044f2;
      8653: inst = 32'h8220000;
      8654: inst = 32'h10408000;
      8655: inst = 32'hc4044f3;
      8656: inst = 32'h8220000;
      8657: inst = 32'h10408000;
      8658: inst = 32'hc4044f4;
      8659: inst = 32'h8220000;
      8660: inst = 32'h10408000;
      8661: inst = 32'hc4044f5;
      8662: inst = 32'h8220000;
      8663: inst = 32'h10408000;
      8664: inst = 32'hc4044f6;
      8665: inst = 32'h8220000;
      8666: inst = 32'h10408000;
      8667: inst = 32'hc4044f7;
      8668: inst = 32'h8220000;
      8669: inst = 32'h10408000;
      8670: inst = 32'hc4044f8;
      8671: inst = 32'h8220000;
      8672: inst = 32'h10408000;
      8673: inst = 32'hc4044f9;
      8674: inst = 32'h8220000;
      8675: inst = 32'h10408000;
      8676: inst = 32'hc4044fa;
      8677: inst = 32'h8220000;
      8678: inst = 32'h10408000;
      8679: inst = 32'hc4044fb;
      8680: inst = 32'h8220000;
      8681: inst = 32'h10408000;
      8682: inst = 32'hc4044fc;
      8683: inst = 32'h8220000;
      8684: inst = 32'h10408000;
      8685: inst = 32'hc4044fd;
      8686: inst = 32'h8220000;
      8687: inst = 32'h10408000;
      8688: inst = 32'hc4044fe;
      8689: inst = 32'h8220000;
      8690: inst = 32'h10408000;
      8691: inst = 32'hc4044ff;
      8692: inst = 32'h8220000;
      8693: inst = 32'h10408000;
      8694: inst = 32'hc404500;
      8695: inst = 32'h8220000;
      8696: inst = 32'h10408000;
      8697: inst = 32'hc404501;
      8698: inst = 32'h8220000;
      8699: inst = 32'h10408000;
      8700: inst = 32'hc404502;
      8701: inst = 32'h8220000;
      8702: inst = 32'h10408000;
      8703: inst = 32'hc404503;
      8704: inst = 32'h8220000;
      8705: inst = 32'h10408000;
      8706: inst = 32'hc40453c;
      8707: inst = 32'h8220000;
      8708: inst = 32'h10408000;
      8709: inst = 32'hc40453d;
      8710: inst = 32'h8220000;
      8711: inst = 32'h10408000;
      8712: inst = 32'hc40453e;
      8713: inst = 32'h8220000;
      8714: inst = 32'h10408000;
      8715: inst = 32'hc40453f;
      8716: inst = 32'h8220000;
      8717: inst = 32'h10408000;
      8718: inst = 32'hc404540;
      8719: inst = 32'h8220000;
      8720: inst = 32'h10408000;
      8721: inst = 32'hc404541;
      8722: inst = 32'h8220000;
      8723: inst = 32'h10408000;
      8724: inst = 32'hc404542;
      8725: inst = 32'h8220000;
      8726: inst = 32'h10408000;
      8727: inst = 32'hc404543;
      8728: inst = 32'h8220000;
      8729: inst = 32'h10408000;
      8730: inst = 32'hc404544;
      8731: inst = 32'h8220000;
      8732: inst = 32'h10408000;
      8733: inst = 32'hc404545;
      8734: inst = 32'h8220000;
      8735: inst = 32'h10408000;
      8736: inst = 32'hc404546;
      8737: inst = 32'h8220000;
      8738: inst = 32'h10408000;
      8739: inst = 32'hc404547;
      8740: inst = 32'h8220000;
      8741: inst = 32'h10408000;
      8742: inst = 32'hc404548;
      8743: inst = 32'h8220000;
      8744: inst = 32'h10408000;
      8745: inst = 32'hc404549;
      8746: inst = 32'h8220000;
      8747: inst = 32'h10408000;
      8748: inst = 32'hc40454a;
      8749: inst = 32'h8220000;
      8750: inst = 32'h10408000;
      8751: inst = 32'hc40454b;
      8752: inst = 32'h8220000;
      8753: inst = 32'h10408000;
      8754: inst = 32'hc40454c;
      8755: inst = 32'h8220000;
      8756: inst = 32'h10408000;
      8757: inst = 32'hc40454d;
      8758: inst = 32'h8220000;
      8759: inst = 32'h10408000;
      8760: inst = 32'hc40454e;
      8761: inst = 32'h8220000;
      8762: inst = 32'h10408000;
      8763: inst = 32'hc40454f;
      8764: inst = 32'h8220000;
      8765: inst = 32'h10408000;
      8766: inst = 32'hc404550;
      8767: inst = 32'h8220000;
      8768: inst = 32'h10408000;
      8769: inst = 32'hc404551;
      8770: inst = 32'h8220000;
      8771: inst = 32'h10408000;
      8772: inst = 32'hc404552;
      8773: inst = 32'h8220000;
      8774: inst = 32'h10408000;
      8775: inst = 32'hc404553;
      8776: inst = 32'h8220000;
      8777: inst = 32'h10408000;
      8778: inst = 32'hc404554;
      8779: inst = 32'h8220000;
      8780: inst = 32'h10408000;
      8781: inst = 32'hc404555;
      8782: inst = 32'h8220000;
      8783: inst = 32'h10408000;
      8784: inst = 32'hc404556;
      8785: inst = 32'h8220000;
      8786: inst = 32'h10408000;
      8787: inst = 32'hc404557;
      8788: inst = 32'h8220000;
      8789: inst = 32'h10408000;
      8790: inst = 32'hc404558;
      8791: inst = 32'h8220000;
      8792: inst = 32'h10408000;
      8793: inst = 32'hc404559;
      8794: inst = 32'h8220000;
      8795: inst = 32'h10408000;
      8796: inst = 32'hc40455a;
      8797: inst = 32'h8220000;
      8798: inst = 32'h10408000;
      8799: inst = 32'hc40455b;
      8800: inst = 32'h8220000;
      8801: inst = 32'h10408000;
      8802: inst = 32'hc40455c;
      8803: inst = 32'h8220000;
      8804: inst = 32'h10408000;
      8805: inst = 32'hc40455d;
      8806: inst = 32'h8220000;
      8807: inst = 32'h10408000;
      8808: inst = 32'hc40455e;
      8809: inst = 32'h8220000;
      8810: inst = 32'h10408000;
      8811: inst = 32'hc40455f;
      8812: inst = 32'h8220000;
      8813: inst = 32'h10408000;
      8814: inst = 32'hc404560;
      8815: inst = 32'h8220000;
      8816: inst = 32'h10408000;
      8817: inst = 32'hc404561;
      8818: inst = 32'h8220000;
      8819: inst = 32'h10408000;
      8820: inst = 32'hc404562;
      8821: inst = 32'h8220000;
      8822: inst = 32'h10408000;
      8823: inst = 32'hc404563;
      8824: inst = 32'h8220000;
      8825: inst = 32'h10408000;
      8826: inst = 32'hc40459c;
      8827: inst = 32'h8220000;
      8828: inst = 32'h10408000;
      8829: inst = 32'hc40459d;
      8830: inst = 32'h8220000;
      8831: inst = 32'h10408000;
      8832: inst = 32'hc40459e;
      8833: inst = 32'h8220000;
      8834: inst = 32'h10408000;
      8835: inst = 32'hc40459f;
      8836: inst = 32'h8220000;
      8837: inst = 32'h10408000;
      8838: inst = 32'hc4045a0;
      8839: inst = 32'h8220000;
      8840: inst = 32'h10408000;
      8841: inst = 32'hc4045a1;
      8842: inst = 32'h8220000;
      8843: inst = 32'h10408000;
      8844: inst = 32'hc4045a2;
      8845: inst = 32'h8220000;
      8846: inst = 32'h10408000;
      8847: inst = 32'hc4045a3;
      8848: inst = 32'h8220000;
      8849: inst = 32'h10408000;
      8850: inst = 32'hc4045a4;
      8851: inst = 32'h8220000;
      8852: inst = 32'h10408000;
      8853: inst = 32'hc4045a5;
      8854: inst = 32'h8220000;
      8855: inst = 32'h10408000;
      8856: inst = 32'hc4045a6;
      8857: inst = 32'h8220000;
      8858: inst = 32'h10408000;
      8859: inst = 32'hc4045a7;
      8860: inst = 32'h8220000;
      8861: inst = 32'h10408000;
      8862: inst = 32'hc4045a8;
      8863: inst = 32'h8220000;
      8864: inst = 32'h10408000;
      8865: inst = 32'hc4045a9;
      8866: inst = 32'h8220000;
      8867: inst = 32'h10408000;
      8868: inst = 32'hc4045aa;
      8869: inst = 32'h8220000;
      8870: inst = 32'h10408000;
      8871: inst = 32'hc4045ab;
      8872: inst = 32'h8220000;
      8873: inst = 32'h10408000;
      8874: inst = 32'hc4045ac;
      8875: inst = 32'h8220000;
      8876: inst = 32'h10408000;
      8877: inst = 32'hc4045ad;
      8878: inst = 32'h8220000;
      8879: inst = 32'h10408000;
      8880: inst = 32'hc4045ae;
      8881: inst = 32'h8220000;
      8882: inst = 32'h10408000;
      8883: inst = 32'hc4045af;
      8884: inst = 32'h8220000;
      8885: inst = 32'h10408000;
      8886: inst = 32'hc4045b0;
      8887: inst = 32'h8220000;
      8888: inst = 32'h10408000;
      8889: inst = 32'hc4045b1;
      8890: inst = 32'h8220000;
      8891: inst = 32'h10408000;
      8892: inst = 32'hc4045b2;
      8893: inst = 32'h8220000;
      8894: inst = 32'h10408000;
      8895: inst = 32'hc4045b3;
      8896: inst = 32'h8220000;
      8897: inst = 32'h10408000;
      8898: inst = 32'hc4045b4;
      8899: inst = 32'h8220000;
      8900: inst = 32'h10408000;
      8901: inst = 32'hc4045b5;
      8902: inst = 32'h8220000;
      8903: inst = 32'h10408000;
      8904: inst = 32'hc4045b6;
      8905: inst = 32'h8220000;
      8906: inst = 32'h10408000;
      8907: inst = 32'hc4045b7;
      8908: inst = 32'h8220000;
      8909: inst = 32'h10408000;
      8910: inst = 32'hc4045b8;
      8911: inst = 32'h8220000;
      8912: inst = 32'h10408000;
      8913: inst = 32'hc4045b9;
      8914: inst = 32'h8220000;
      8915: inst = 32'h10408000;
      8916: inst = 32'hc4045ba;
      8917: inst = 32'h8220000;
      8918: inst = 32'h10408000;
      8919: inst = 32'hc4045bb;
      8920: inst = 32'h8220000;
      8921: inst = 32'h10408000;
      8922: inst = 32'hc4045bc;
      8923: inst = 32'h8220000;
      8924: inst = 32'h10408000;
      8925: inst = 32'hc4045bd;
      8926: inst = 32'h8220000;
      8927: inst = 32'h10408000;
      8928: inst = 32'hc4045be;
      8929: inst = 32'h8220000;
      8930: inst = 32'h10408000;
      8931: inst = 32'hc4045bf;
      8932: inst = 32'h8220000;
      8933: inst = 32'h10408000;
      8934: inst = 32'hc4045c0;
      8935: inst = 32'h8220000;
      8936: inst = 32'h10408000;
      8937: inst = 32'hc4045c1;
      8938: inst = 32'h8220000;
      8939: inst = 32'h10408000;
      8940: inst = 32'hc4045c2;
      8941: inst = 32'h8220000;
      8942: inst = 32'h10408000;
      8943: inst = 32'hc4045c3;
      8944: inst = 32'h8220000;
      8945: inst = 32'h10408000;
      8946: inst = 32'hc4045fc;
      8947: inst = 32'h8220000;
      8948: inst = 32'h10408000;
      8949: inst = 32'hc4045fd;
      8950: inst = 32'h8220000;
      8951: inst = 32'h10408000;
      8952: inst = 32'hc4045fe;
      8953: inst = 32'h8220000;
      8954: inst = 32'h10408000;
      8955: inst = 32'hc4045ff;
      8956: inst = 32'h8220000;
      8957: inst = 32'h10408000;
      8958: inst = 32'hc404600;
      8959: inst = 32'h8220000;
      8960: inst = 32'h10408000;
      8961: inst = 32'hc404601;
      8962: inst = 32'h8220000;
      8963: inst = 32'h10408000;
      8964: inst = 32'hc404602;
      8965: inst = 32'h8220000;
      8966: inst = 32'h10408000;
      8967: inst = 32'hc404603;
      8968: inst = 32'h8220000;
      8969: inst = 32'h10408000;
      8970: inst = 32'hc404604;
      8971: inst = 32'h8220000;
      8972: inst = 32'h10408000;
      8973: inst = 32'hc404605;
      8974: inst = 32'h8220000;
      8975: inst = 32'h10408000;
      8976: inst = 32'hc404606;
      8977: inst = 32'h8220000;
      8978: inst = 32'h10408000;
      8979: inst = 32'hc404607;
      8980: inst = 32'h8220000;
      8981: inst = 32'h10408000;
      8982: inst = 32'hc404608;
      8983: inst = 32'h8220000;
      8984: inst = 32'h10408000;
      8985: inst = 32'hc404609;
      8986: inst = 32'h8220000;
      8987: inst = 32'h10408000;
      8988: inst = 32'hc40460a;
      8989: inst = 32'h8220000;
      8990: inst = 32'h10408000;
      8991: inst = 32'hc40460b;
      8992: inst = 32'h8220000;
      8993: inst = 32'h10408000;
      8994: inst = 32'hc40460c;
      8995: inst = 32'h8220000;
      8996: inst = 32'h10408000;
      8997: inst = 32'hc40460d;
      8998: inst = 32'h8220000;
      8999: inst = 32'h10408000;
      9000: inst = 32'hc40460e;
      9001: inst = 32'h8220000;
      9002: inst = 32'h10408000;
      9003: inst = 32'hc40460f;
      9004: inst = 32'h8220000;
      9005: inst = 32'h10408000;
      9006: inst = 32'hc404610;
      9007: inst = 32'h8220000;
      9008: inst = 32'h10408000;
      9009: inst = 32'hc404611;
      9010: inst = 32'h8220000;
      9011: inst = 32'h10408000;
      9012: inst = 32'hc404612;
      9013: inst = 32'h8220000;
      9014: inst = 32'h10408000;
      9015: inst = 32'hc404613;
      9016: inst = 32'h8220000;
      9017: inst = 32'h10408000;
      9018: inst = 32'hc404614;
      9019: inst = 32'h8220000;
      9020: inst = 32'h10408000;
      9021: inst = 32'hc404615;
      9022: inst = 32'h8220000;
      9023: inst = 32'h10408000;
      9024: inst = 32'hc404616;
      9025: inst = 32'h8220000;
      9026: inst = 32'h10408000;
      9027: inst = 32'hc404617;
      9028: inst = 32'h8220000;
      9029: inst = 32'h10408000;
      9030: inst = 32'hc404618;
      9031: inst = 32'h8220000;
      9032: inst = 32'h10408000;
      9033: inst = 32'hc404619;
      9034: inst = 32'h8220000;
      9035: inst = 32'h10408000;
      9036: inst = 32'hc40461a;
      9037: inst = 32'h8220000;
      9038: inst = 32'h10408000;
      9039: inst = 32'hc40461b;
      9040: inst = 32'h8220000;
      9041: inst = 32'h10408000;
      9042: inst = 32'hc40461c;
      9043: inst = 32'h8220000;
      9044: inst = 32'h10408000;
      9045: inst = 32'hc40461d;
      9046: inst = 32'h8220000;
      9047: inst = 32'h10408000;
      9048: inst = 32'hc40461e;
      9049: inst = 32'h8220000;
      9050: inst = 32'h10408000;
      9051: inst = 32'hc40461f;
      9052: inst = 32'h8220000;
      9053: inst = 32'h10408000;
      9054: inst = 32'hc404620;
      9055: inst = 32'h8220000;
      9056: inst = 32'h10408000;
      9057: inst = 32'hc404621;
      9058: inst = 32'h8220000;
      9059: inst = 32'h10408000;
      9060: inst = 32'hc404622;
      9061: inst = 32'h8220000;
      9062: inst = 32'h10408000;
      9063: inst = 32'hc404623;
      9064: inst = 32'h8220000;
      9065: inst = 32'h10408000;
      9066: inst = 32'hc40465c;
      9067: inst = 32'h8220000;
      9068: inst = 32'h10408000;
      9069: inst = 32'hc40465d;
      9070: inst = 32'h8220000;
      9071: inst = 32'h10408000;
      9072: inst = 32'hc40465e;
      9073: inst = 32'h8220000;
      9074: inst = 32'h10408000;
      9075: inst = 32'hc40465f;
      9076: inst = 32'h8220000;
      9077: inst = 32'h10408000;
      9078: inst = 32'hc404660;
      9079: inst = 32'h8220000;
      9080: inst = 32'h10408000;
      9081: inst = 32'hc404661;
      9082: inst = 32'h8220000;
      9083: inst = 32'h10408000;
      9084: inst = 32'hc404662;
      9085: inst = 32'h8220000;
      9086: inst = 32'h10408000;
      9087: inst = 32'hc404663;
      9088: inst = 32'h8220000;
      9089: inst = 32'h10408000;
      9090: inst = 32'hc404664;
      9091: inst = 32'h8220000;
      9092: inst = 32'h10408000;
      9093: inst = 32'hc404665;
      9094: inst = 32'h8220000;
      9095: inst = 32'h10408000;
      9096: inst = 32'hc404666;
      9097: inst = 32'h8220000;
      9098: inst = 32'h10408000;
      9099: inst = 32'hc404667;
      9100: inst = 32'h8220000;
      9101: inst = 32'h10408000;
      9102: inst = 32'hc404668;
      9103: inst = 32'h8220000;
      9104: inst = 32'h10408000;
      9105: inst = 32'hc404669;
      9106: inst = 32'h8220000;
      9107: inst = 32'h10408000;
      9108: inst = 32'hc40466a;
      9109: inst = 32'h8220000;
      9110: inst = 32'h10408000;
      9111: inst = 32'hc40466b;
      9112: inst = 32'h8220000;
      9113: inst = 32'h10408000;
      9114: inst = 32'hc40466c;
      9115: inst = 32'h8220000;
      9116: inst = 32'h10408000;
      9117: inst = 32'hc40466d;
      9118: inst = 32'h8220000;
      9119: inst = 32'h10408000;
      9120: inst = 32'hc40466e;
      9121: inst = 32'h8220000;
      9122: inst = 32'h10408000;
      9123: inst = 32'hc40466f;
      9124: inst = 32'h8220000;
      9125: inst = 32'h10408000;
      9126: inst = 32'hc404670;
      9127: inst = 32'h8220000;
      9128: inst = 32'h10408000;
      9129: inst = 32'hc404671;
      9130: inst = 32'h8220000;
      9131: inst = 32'h10408000;
      9132: inst = 32'hc404672;
      9133: inst = 32'h8220000;
      9134: inst = 32'h10408000;
      9135: inst = 32'hc404673;
      9136: inst = 32'h8220000;
      9137: inst = 32'h10408000;
      9138: inst = 32'hc404674;
      9139: inst = 32'h8220000;
      9140: inst = 32'h10408000;
      9141: inst = 32'hc404675;
      9142: inst = 32'h8220000;
      9143: inst = 32'h10408000;
      9144: inst = 32'hc404676;
      9145: inst = 32'h8220000;
      9146: inst = 32'h10408000;
      9147: inst = 32'hc404677;
      9148: inst = 32'h8220000;
      9149: inst = 32'h10408000;
      9150: inst = 32'hc404678;
      9151: inst = 32'h8220000;
      9152: inst = 32'h10408000;
      9153: inst = 32'hc404679;
      9154: inst = 32'h8220000;
      9155: inst = 32'h10408000;
      9156: inst = 32'hc40467a;
      9157: inst = 32'h8220000;
      9158: inst = 32'h10408000;
      9159: inst = 32'hc40467b;
      9160: inst = 32'h8220000;
      9161: inst = 32'h10408000;
      9162: inst = 32'hc40467c;
      9163: inst = 32'h8220000;
      9164: inst = 32'h10408000;
      9165: inst = 32'hc40467d;
      9166: inst = 32'h8220000;
      9167: inst = 32'h10408000;
      9168: inst = 32'hc40467e;
      9169: inst = 32'h8220000;
      9170: inst = 32'h10408000;
      9171: inst = 32'hc40467f;
      9172: inst = 32'h8220000;
      9173: inst = 32'h10408000;
      9174: inst = 32'hc404680;
      9175: inst = 32'h8220000;
      9176: inst = 32'h10408000;
      9177: inst = 32'hc404681;
      9178: inst = 32'h8220000;
      9179: inst = 32'h10408000;
      9180: inst = 32'hc404682;
      9181: inst = 32'h8220000;
      9182: inst = 32'h10408000;
      9183: inst = 32'hc404683;
      9184: inst = 32'h8220000;
      9185: inst = 32'h10408000;
      9186: inst = 32'hc4046bc;
      9187: inst = 32'h8220000;
      9188: inst = 32'h10408000;
      9189: inst = 32'hc4046bd;
      9190: inst = 32'h8220000;
      9191: inst = 32'h10408000;
      9192: inst = 32'hc4046be;
      9193: inst = 32'h8220000;
      9194: inst = 32'h10408000;
      9195: inst = 32'hc4046bf;
      9196: inst = 32'h8220000;
      9197: inst = 32'h10408000;
      9198: inst = 32'hc4046c0;
      9199: inst = 32'h8220000;
      9200: inst = 32'h10408000;
      9201: inst = 32'hc4046c1;
      9202: inst = 32'h8220000;
      9203: inst = 32'h10408000;
      9204: inst = 32'hc4046c2;
      9205: inst = 32'h8220000;
      9206: inst = 32'h10408000;
      9207: inst = 32'hc4046c3;
      9208: inst = 32'h8220000;
      9209: inst = 32'h10408000;
      9210: inst = 32'hc4046c4;
      9211: inst = 32'h8220000;
      9212: inst = 32'h10408000;
      9213: inst = 32'hc4046c5;
      9214: inst = 32'h8220000;
      9215: inst = 32'h10408000;
      9216: inst = 32'hc4046c6;
      9217: inst = 32'h8220000;
      9218: inst = 32'h10408000;
      9219: inst = 32'hc4046c7;
      9220: inst = 32'h8220000;
      9221: inst = 32'h10408000;
      9222: inst = 32'hc4046c8;
      9223: inst = 32'h8220000;
      9224: inst = 32'h10408000;
      9225: inst = 32'hc4046c9;
      9226: inst = 32'h8220000;
      9227: inst = 32'h10408000;
      9228: inst = 32'hc4046ca;
      9229: inst = 32'h8220000;
      9230: inst = 32'h10408000;
      9231: inst = 32'hc4046cb;
      9232: inst = 32'h8220000;
      9233: inst = 32'h10408000;
      9234: inst = 32'hc4046cc;
      9235: inst = 32'h8220000;
      9236: inst = 32'h10408000;
      9237: inst = 32'hc4046cd;
      9238: inst = 32'h8220000;
      9239: inst = 32'h10408000;
      9240: inst = 32'hc4046ce;
      9241: inst = 32'h8220000;
      9242: inst = 32'h10408000;
      9243: inst = 32'hc4046cf;
      9244: inst = 32'h8220000;
      9245: inst = 32'h10408000;
      9246: inst = 32'hc4046d0;
      9247: inst = 32'h8220000;
      9248: inst = 32'h10408000;
      9249: inst = 32'hc4046d1;
      9250: inst = 32'h8220000;
      9251: inst = 32'h10408000;
      9252: inst = 32'hc4046d2;
      9253: inst = 32'h8220000;
      9254: inst = 32'h10408000;
      9255: inst = 32'hc4046d3;
      9256: inst = 32'h8220000;
      9257: inst = 32'h10408000;
      9258: inst = 32'hc4046d4;
      9259: inst = 32'h8220000;
      9260: inst = 32'h10408000;
      9261: inst = 32'hc4046d5;
      9262: inst = 32'h8220000;
      9263: inst = 32'h10408000;
      9264: inst = 32'hc4046d6;
      9265: inst = 32'h8220000;
      9266: inst = 32'h10408000;
      9267: inst = 32'hc4046d7;
      9268: inst = 32'h8220000;
      9269: inst = 32'h10408000;
      9270: inst = 32'hc4046d8;
      9271: inst = 32'h8220000;
      9272: inst = 32'h10408000;
      9273: inst = 32'hc4046d9;
      9274: inst = 32'h8220000;
      9275: inst = 32'h10408000;
      9276: inst = 32'hc4046da;
      9277: inst = 32'h8220000;
      9278: inst = 32'h10408000;
      9279: inst = 32'hc4046db;
      9280: inst = 32'h8220000;
      9281: inst = 32'h10408000;
      9282: inst = 32'hc4046dc;
      9283: inst = 32'h8220000;
      9284: inst = 32'h10408000;
      9285: inst = 32'hc4046dd;
      9286: inst = 32'h8220000;
      9287: inst = 32'h10408000;
      9288: inst = 32'hc4046de;
      9289: inst = 32'h8220000;
      9290: inst = 32'h10408000;
      9291: inst = 32'hc4046df;
      9292: inst = 32'h8220000;
      9293: inst = 32'h10408000;
      9294: inst = 32'hc4046e0;
      9295: inst = 32'h8220000;
      9296: inst = 32'h10408000;
      9297: inst = 32'hc4046e1;
      9298: inst = 32'h8220000;
      9299: inst = 32'h10408000;
      9300: inst = 32'hc4046e2;
      9301: inst = 32'h8220000;
      9302: inst = 32'h10408000;
      9303: inst = 32'hc4046e3;
      9304: inst = 32'h8220000;
      9305: inst = 32'h10408000;
      9306: inst = 32'hc40471c;
      9307: inst = 32'h8220000;
      9308: inst = 32'h10408000;
      9309: inst = 32'hc40471d;
      9310: inst = 32'h8220000;
      9311: inst = 32'h10408000;
      9312: inst = 32'hc40471e;
      9313: inst = 32'h8220000;
      9314: inst = 32'h10408000;
      9315: inst = 32'hc40471f;
      9316: inst = 32'h8220000;
      9317: inst = 32'h10408000;
      9318: inst = 32'hc404720;
      9319: inst = 32'h8220000;
      9320: inst = 32'h10408000;
      9321: inst = 32'hc404721;
      9322: inst = 32'h8220000;
      9323: inst = 32'h10408000;
      9324: inst = 32'hc404722;
      9325: inst = 32'h8220000;
      9326: inst = 32'h10408000;
      9327: inst = 32'hc404723;
      9328: inst = 32'h8220000;
      9329: inst = 32'h10408000;
      9330: inst = 32'hc404724;
      9331: inst = 32'h8220000;
      9332: inst = 32'h10408000;
      9333: inst = 32'hc404725;
      9334: inst = 32'h8220000;
      9335: inst = 32'h10408000;
      9336: inst = 32'hc404726;
      9337: inst = 32'h8220000;
      9338: inst = 32'h10408000;
      9339: inst = 32'hc404727;
      9340: inst = 32'h8220000;
      9341: inst = 32'h10408000;
      9342: inst = 32'hc404728;
      9343: inst = 32'h8220000;
      9344: inst = 32'h10408000;
      9345: inst = 32'hc404729;
      9346: inst = 32'h8220000;
      9347: inst = 32'h10408000;
      9348: inst = 32'hc40472a;
      9349: inst = 32'h8220000;
      9350: inst = 32'h10408000;
      9351: inst = 32'hc40472b;
      9352: inst = 32'h8220000;
      9353: inst = 32'h10408000;
      9354: inst = 32'hc40472c;
      9355: inst = 32'h8220000;
      9356: inst = 32'h10408000;
      9357: inst = 32'hc40472d;
      9358: inst = 32'h8220000;
      9359: inst = 32'h10408000;
      9360: inst = 32'hc40472e;
      9361: inst = 32'h8220000;
      9362: inst = 32'h10408000;
      9363: inst = 32'hc40472f;
      9364: inst = 32'h8220000;
      9365: inst = 32'h10408000;
      9366: inst = 32'hc404730;
      9367: inst = 32'h8220000;
      9368: inst = 32'h10408000;
      9369: inst = 32'hc404731;
      9370: inst = 32'h8220000;
      9371: inst = 32'h10408000;
      9372: inst = 32'hc404732;
      9373: inst = 32'h8220000;
      9374: inst = 32'h10408000;
      9375: inst = 32'hc404733;
      9376: inst = 32'h8220000;
      9377: inst = 32'h10408000;
      9378: inst = 32'hc404734;
      9379: inst = 32'h8220000;
      9380: inst = 32'h10408000;
      9381: inst = 32'hc404735;
      9382: inst = 32'h8220000;
      9383: inst = 32'h10408000;
      9384: inst = 32'hc404736;
      9385: inst = 32'h8220000;
      9386: inst = 32'h10408000;
      9387: inst = 32'hc404737;
      9388: inst = 32'h8220000;
      9389: inst = 32'h10408000;
      9390: inst = 32'hc404738;
      9391: inst = 32'h8220000;
      9392: inst = 32'h10408000;
      9393: inst = 32'hc404739;
      9394: inst = 32'h8220000;
      9395: inst = 32'h10408000;
      9396: inst = 32'hc40473a;
      9397: inst = 32'h8220000;
      9398: inst = 32'h10408000;
      9399: inst = 32'hc40473b;
      9400: inst = 32'h8220000;
      9401: inst = 32'h10408000;
      9402: inst = 32'hc40473c;
      9403: inst = 32'h8220000;
      9404: inst = 32'h10408000;
      9405: inst = 32'hc40473d;
      9406: inst = 32'h8220000;
      9407: inst = 32'h10408000;
      9408: inst = 32'hc40473e;
      9409: inst = 32'h8220000;
      9410: inst = 32'h10408000;
      9411: inst = 32'hc40473f;
      9412: inst = 32'h8220000;
      9413: inst = 32'h10408000;
      9414: inst = 32'hc404740;
      9415: inst = 32'h8220000;
      9416: inst = 32'h10408000;
      9417: inst = 32'hc404741;
      9418: inst = 32'h8220000;
      9419: inst = 32'h10408000;
      9420: inst = 32'hc404742;
      9421: inst = 32'h8220000;
      9422: inst = 32'h10408000;
      9423: inst = 32'hc404743;
      9424: inst = 32'h8220000;
      9425: inst = 32'h10408000;
      9426: inst = 32'hc40477c;
      9427: inst = 32'h8220000;
      9428: inst = 32'h10408000;
      9429: inst = 32'hc40477d;
      9430: inst = 32'h8220000;
      9431: inst = 32'h10408000;
      9432: inst = 32'hc40477e;
      9433: inst = 32'h8220000;
      9434: inst = 32'h10408000;
      9435: inst = 32'hc40477f;
      9436: inst = 32'h8220000;
      9437: inst = 32'h10408000;
      9438: inst = 32'hc404780;
      9439: inst = 32'h8220000;
      9440: inst = 32'h10408000;
      9441: inst = 32'hc404781;
      9442: inst = 32'h8220000;
      9443: inst = 32'h10408000;
      9444: inst = 32'hc404782;
      9445: inst = 32'h8220000;
      9446: inst = 32'h10408000;
      9447: inst = 32'hc404783;
      9448: inst = 32'h8220000;
      9449: inst = 32'h10408000;
      9450: inst = 32'hc404784;
      9451: inst = 32'h8220000;
      9452: inst = 32'h10408000;
      9453: inst = 32'hc404785;
      9454: inst = 32'h8220000;
      9455: inst = 32'h10408000;
      9456: inst = 32'hc404786;
      9457: inst = 32'h8220000;
      9458: inst = 32'h10408000;
      9459: inst = 32'hc404787;
      9460: inst = 32'h8220000;
      9461: inst = 32'h10408000;
      9462: inst = 32'hc404788;
      9463: inst = 32'h8220000;
      9464: inst = 32'h10408000;
      9465: inst = 32'hc404789;
      9466: inst = 32'h8220000;
      9467: inst = 32'h10408000;
      9468: inst = 32'hc40478a;
      9469: inst = 32'h8220000;
      9470: inst = 32'h10408000;
      9471: inst = 32'hc40478b;
      9472: inst = 32'h8220000;
      9473: inst = 32'h10408000;
      9474: inst = 32'hc40478c;
      9475: inst = 32'h8220000;
      9476: inst = 32'h10408000;
      9477: inst = 32'hc40478d;
      9478: inst = 32'h8220000;
      9479: inst = 32'h10408000;
      9480: inst = 32'hc40478e;
      9481: inst = 32'h8220000;
      9482: inst = 32'h10408000;
      9483: inst = 32'hc40478f;
      9484: inst = 32'h8220000;
      9485: inst = 32'h10408000;
      9486: inst = 32'hc404790;
      9487: inst = 32'h8220000;
      9488: inst = 32'h10408000;
      9489: inst = 32'hc404791;
      9490: inst = 32'h8220000;
      9491: inst = 32'h10408000;
      9492: inst = 32'hc404792;
      9493: inst = 32'h8220000;
      9494: inst = 32'h10408000;
      9495: inst = 32'hc404793;
      9496: inst = 32'h8220000;
      9497: inst = 32'h10408000;
      9498: inst = 32'hc404794;
      9499: inst = 32'h8220000;
      9500: inst = 32'h10408000;
      9501: inst = 32'hc404795;
      9502: inst = 32'h8220000;
      9503: inst = 32'h10408000;
      9504: inst = 32'hc404796;
      9505: inst = 32'h8220000;
      9506: inst = 32'h10408000;
      9507: inst = 32'hc404797;
      9508: inst = 32'h8220000;
      9509: inst = 32'h10408000;
      9510: inst = 32'hc404798;
      9511: inst = 32'h8220000;
      9512: inst = 32'h10408000;
      9513: inst = 32'hc404799;
      9514: inst = 32'h8220000;
      9515: inst = 32'h10408000;
      9516: inst = 32'hc40479a;
      9517: inst = 32'h8220000;
      9518: inst = 32'h10408000;
      9519: inst = 32'hc40479b;
      9520: inst = 32'h8220000;
      9521: inst = 32'h10408000;
      9522: inst = 32'hc40479c;
      9523: inst = 32'h8220000;
      9524: inst = 32'h10408000;
      9525: inst = 32'hc40479d;
      9526: inst = 32'h8220000;
      9527: inst = 32'h10408000;
      9528: inst = 32'hc40479e;
      9529: inst = 32'h8220000;
      9530: inst = 32'h10408000;
      9531: inst = 32'hc40479f;
      9532: inst = 32'h8220000;
      9533: inst = 32'h10408000;
      9534: inst = 32'hc4047a0;
      9535: inst = 32'h8220000;
      9536: inst = 32'h10408000;
      9537: inst = 32'hc4047a1;
      9538: inst = 32'h8220000;
      9539: inst = 32'h10408000;
      9540: inst = 32'hc4047a2;
      9541: inst = 32'h8220000;
      9542: inst = 32'h10408000;
      9543: inst = 32'hc4047a3;
      9544: inst = 32'h8220000;
      9545: inst = 32'h10408000;
      9546: inst = 32'hc4047dc;
      9547: inst = 32'h8220000;
      9548: inst = 32'h10408000;
      9549: inst = 32'hc4047dd;
      9550: inst = 32'h8220000;
      9551: inst = 32'h10408000;
      9552: inst = 32'hc4047de;
      9553: inst = 32'h8220000;
      9554: inst = 32'h10408000;
      9555: inst = 32'hc4047df;
      9556: inst = 32'h8220000;
      9557: inst = 32'h10408000;
      9558: inst = 32'hc4047e0;
      9559: inst = 32'h8220000;
      9560: inst = 32'h10408000;
      9561: inst = 32'hc4047e1;
      9562: inst = 32'h8220000;
      9563: inst = 32'h10408000;
      9564: inst = 32'hc4047e2;
      9565: inst = 32'h8220000;
      9566: inst = 32'h10408000;
      9567: inst = 32'hc4047e3;
      9568: inst = 32'h8220000;
      9569: inst = 32'h10408000;
      9570: inst = 32'hc4047e4;
      9571: inst = 32'h8220000;
      9572: inst = 32'h10408000;
      9573: inst = 32'hc4047e5;
      9574: inst = 32'h8220000;
      9575: inst = 32'h10408000;
      9576: inst = 32'hc4047e6;
      9577: inst = 32'h8220000;
      9578: inst = 32'h10408000;
      9579: inst = 32'hc4047e7;
      9580: inst = 32'h8220000;
      9581: inst = 32'h10408000;
      9582: inst = 32'hc4047e8;
      9583: inst = 32'h8220000;
      9584: inst = 32'h10408000;
      9585: inst = 32'hc4047e9;
      9586: inst = 32'h8220000;
      9587: inst = 32'h10408000;
      9588: inst = 32'hc4047ea;
      9589: inst = 32'h8220000;
      9590: inst = 32'h10408000;
      9591: inst = 32'hc4047eb;
      9592: inst = 32'h8220000;
      9593: inst = 32'h10408000;
      9594: inst = 32'hc4047ec;
      9595: inst = 32'h8220000;
      9596: inst = 32'h10408000;
      9597: inst = 32'hc4047ed;
      9598: inst = 32'h8220000;
      9599: inst = 32'h10408000;
      9600: inst = 32'hc4047ee;
      9601: inst = 32'h8220000;
      9602: inst = 32'h10408000;
      9603: inst = 32'hc4047ef;
      9604: inst = 32'h8220000;
      9605: inst = 32'h10408000;
      9606: inst = 32'hc4047f0;
      9607: inst = 32'h8220000;
      9608: inst = 32'h10408000;
      9609: inst = 32'hc4047f1;
      9610: inst = 32'h8220000;
      9611: inst = 32'h10408000;
      9612: inst = 32'hc4047f2;
      9613: inst = 32'h8220000;
      9614: inst = 32'h10408000;
      9615: inst = 32'hc4047f3;
      9616: inst = 32'h8220000;
      9617: inst = 32'h10408000;
      9618: inst = 32'hc4047f4;
      9619: inst = 32'h8220000;
      9620: inst = 32'h10408000;
      9621: inst = 32'hc4047f5;
      9622: inst = 32'h8220000;
      9623: inst = 32'h10408000;
      9624: inst = 32'hc4047f6;
      9625: inst = 32'h8220000;
      9626: inst = 32'h10408000;
      9627: inst = 32'hc4047f7;
      9628: inst = 32'h8220000;
      9629: inst = 32'h10408000;
      9630: inst = 32'hc4047f8;
      9631: inst = 32'h8220000;
      9632: inst = 32'h10408000;
      9633: inst = 32'hc4047f9;
      9634: inst = 32'h8220000;
      9635: inst = 32'h10408000;
      9636: inst = 32'hc4047fa;
      9637: inst = 32'h8220000;
      9638: inst = 32'h10408000;
      9639: inst = 32'hc4047fb;
      9640: inst = 32'h8220000;
      9641: inst = 32'h10408000;
      9642: inst = 32'hc4047fc;
      9643: inst = 32'h8220000;
      9644: inst = 32'h10408000;
      9645: inst = 32'hc4047fd;
      9646: inst = 32'h8220000;
      9647: inst = 32'h10408000;
      9648: inst = 32'hc4047fe;
      9649: inst = 32'h8220000;
      9650: inst = 32'h10408000;
      9651: inst = 32'hc4047ff;
      9652: inst = 32'h8220000;
      9653: inst = 32'h10408000;
      9654: inst = 32'hc404800;
      9655: inst = 32'h8220000;
      9656: inst = 32'h10408000;
      9657: inst = 32'hc404801;
      9658: inst = 32'h8220000;
      9659: inst = 32'h10408000;
      9660: inst = 32'hc404802;
      9661: inst = 32'h8220000;
      9662: inst = 32'h10408000;
      9663: inst = 32'hc404803;
      9664: inst = 32'h8220000;
      9665: inst = 32'h10408000;
      9666: inst = 32'hc40483c;
      9667: inst = 32'h8220000;
      9668: inst = 32'h10408000;
      9669: inst = 32'hc40483d;
      9670: inst = 32'h8220000;
      9671: inst = 32'h10408000;
      9672: inst = 32'hc40483e;
      9673: inst = 32'h8220000;
      9674: inst = 32'h10408000;
      9675: inst = 32'hc40483f;
      9676: inst = 32'h8220000;
      9677: inst = 32'h10408000;
      9678: inst = 32'hc404840;
      9679: inst = 32'h8220000;
      9680: inst = 32'h10408000;
      9681: inst = 32'hc404841;
      9682: inst = 32'h8220000;
      9683: inst = 32'h10408000;
      9684: inst = 32'hc404842;
      9685: inst = 32'h8220000;
      9686: inst = 32'h10408000;
      9687: inst = 32'hc404843;
      9688: inst = 32'h8220000;
      9689: inst = 32'h10408000;
      9690: inst = 32'hc404844;
      9691: inst = 32'h8220000;
      9692: inst = 32'h10408000;
      9693: inst = 32'hc404845;
      9694: inst = 32'h8220000;
      9695: inst = 32'h10408000;
      9696: inst = 32'hc404846;
      9697: inst = 32'h8220000;
      9698: inst = 32'h10408000;
      9699: inst = 32'hc404847;
      9700: inst = 32'h8220000;
      9701: inst = 32'h10408000;
      9702: inst = 32'hc404848;
      9703: inst = 32'h8220000;
      9704: inst = 32'h10408000;
      9705: inst = 32'hc404849;
      9706: inst = 32'h8220000;
      9707: inst = 32'h10408000;
      9708: inst = 32'hc40484a;
      9709: inst = 32'h8220000;
      9710: inst = 32'h10408000;
      9711: inst = 32'hc40484b;
      9712: inst = 32'h8220000;
      9713: inst = 32'h10408000;
      9714: inst = 32'hc40484c;
      9715: inst = 32'h8220000;
      9716: inst = 32'h10408000;
      9717: inst = 32'hc40484d;
      9718: inst = 32'h8220000;
      9719: inst = 32'h10408000;
      9720: inst = 32'hc40484e;
      9721: inst = 32'h8220000;
      9722: inst = 32'h10408000;
      9723: inst = 32'hc40484f;
      9724: inst = 32'h8220000;
      9725: inst = 32'h10408000;
      9726: inst = 32'hc404850;
      9727: inst = 32'h8220000;
      9728: inst = 32'h10408000;
      9729: inst = 32'hc404851;
      9730: inst = 32'h8220000;
      9731: inst = 32'h10408000;
      9732: inst = 32'hc404852;
      9733: inst = 32'h8220000;
      9734: inst = 32'h10408000;
      9735: inst = 32'hc404853;
      9736: inst = 32'h8220000;
      9737: inst = 32'h10408000;
      9738: inst = 32'hc404854;
      9739: inst = 32'h8220000;
      9740: inst = 32'h10408000;
      9741: inst = 32'hc404855;
      9742: inst = 32'h8220000;
      9743: inst = 32'h10408000;
      9744: inst = 32'hc404856;
      9745: inst = 32'h8220000;
      9746: inst = 32'h10408000;
      9747: inst = 32'hc404857;
      9748: inst = 32'h8220000;
      9749: inst = 32'h10408000;
      9750: inst = 32'hc404858;
      9751: inst = 32'h8220000;
      9752: inst = 32'h10408000;
      9753: inst = 32'hc404859;
      9754: inst = 32'h8220000;
      9755: inst = 32'h10408000;
      9756: inst = 32'hc40485a;
      9757: inst = 32'h8220000;
      9758: inst = 32'h10408000;
      9759: inst = 32'hc40485b;
      9760: inst = 32'h8220000;
      9761: inst = 32'h10408000;
      9762: inst = 32'hc40485c;
      9763: inst = 32'h8220000;
      9764: inst = 32'h10408000;
      9765: inst = 32'hc40485d;
      9766: inst = 32'h8220000;
      9767: inst = 32'h10408000;
      9768: inst = 32'hc40485e;
      9769: inst = 32'h8220000;
      9770: inst = 32'h10408000;
      9771: inst = 32'hc40485f;
      9772: inst = 32'h8220000;
      9773: inst = 32'h10408000;
      9774: inst = 32'hc404860;
      9775: inst = 32'h8220000;
      9776: inst = 32'h10408000;
      9777: inst = 32'hc404861;
      9778: inst = 32'h8220000;
      9779: inst = 32'h10408000;
      9780: inst = 32'hc404862;
      9781: inst = 32'h8220000;
      9782: inst = 32'h10408000;
      9783: inst = 32'hc404863;
      9784: inst = 32'h8220000;
      9785: inst = 32'h10408000;
      9786: inst = 32'hc40489c;
      9787: inst = 32'h8220000;
      9788: inst = 32'h10408000;
      9789: inst = 32'hc40489d;
      9790: inst = 32'h8220000;
      9791: inst = 32'h10408000;
      9792: inst = 32'hc40489e;
      9793: inst = 32'h8220000;
      9794: inst = 32'h10408000;
      9795: inst = 32'hc40489f;
      9796: inst = 32'h8220000;
      9797: inst = 32'h10408000;
      9798: inst = 32'hc4048a0;
      9799: inst = 32'h8220000;
      9800: inst = 32'h10408000;
      9801: inst = 32'hc4048a1;
      9802: inst = 32'h8220000;
      9803: inst = 32'h10408000;
      9804: inst = 32'hc4048a2;
      9805: inst = 32'h8220000;
      9806: inst = 32'h10408000;
      9807: inst = 32'hc4048a3;
      9808: inst = 32'h8220000;
      9809: inst = 32'h10408000;
      9810: inst = 32'hc4048a4;
      9811: inst = 32'h8220000;
      9812: inst = 32'h10408000;
      9813: inst = 32'hc4048a5;
      9814: inst = 32'h8220000;
      9815: inst = 32'h10408000;
      9816: inst = 32'hc4048a6;
      9817: inst = 32'h8220000;
      9818: inst = 32'h10408000;
      9819: inst = 32'hc4048a7;
      9820: inst = 32'h8220000;
      9821: inst = 32'h10408000;
      9822: inst = 32'hc4048a8;
      9823: inst = 32'h8220000;
      9824: inst = 32'h10408000;
      9825: inst = 32'hc4048a9;
      9826: inst = 32'h8220000;
      9827: inst = 32'h10408000;
      9828: inst = 32'hc4048aa;
      9829: inst = 32'h8220000;
      9830: inst = 32'h10408000;
      9831: inst = 32'hc4048ab;
      9832: inst = 32'h8220000;
      9833: inst = 32'h10408000;
      9834: inst = 32'hc4048ac;
      9835: inst = 32'h8220000;
      9836: inst = 32'h10408000;
      9837: inst = 32'hc4048ad;
      9838: inst = 32'h8220000;
      9839: inst = 32'h10408000;
      9840: inst = 32'hc4048ae;
      9841: inst = 32'h8220000;
      9842: inst = 32'h10408000;
      9843: inst = 32'hc4048af;
      9844: inst = 32'h8220000;
      9845: inst = 32'h10408000;
      9846: inst = 32'hc4048b0;
      9847: inst = 32'h8220000;
      9848: inst = 32'h10408000;
      9849: inst = 32'hc4048b1;
      9850: inst = 32'h8220000;
      9851: inst = 32'h10408000;
      9852: inst = 32'hc4048b2;
      9853: inst = 32'h8220000;
      9854: inst = 32'h10408000;
      9855: inst = 32'hc4048b3;
      9856: inst = 32'h8220000;
      9857: inst = 32'h10408000;
      9858: inst = 32'hc4048b4;
      9859: inst = 32'h8220000;
      9860: inst = 32'h10408000;
      9861: inst = 32'hc4048b5;
      9862: inst = 32'h8220000;
      9863: inst = 32'h10408000;
      9864: inst = 32'hc4048b6;
      9865: inst = 32'h8220000;
      9866: inst = 32'h10408000;
      9867: inst = 32'hc4048b7;
      9868: inst = 32'h8220000;
      9869: inst = 32'h10408000;
      9870: inst = 32'hc4048b8;
      9871: inst = 32'h8220000;
      9872: inst = 32'h10408000;
      9873: inst = 32'hc4048b9;
      9874: inst = 32'h8220000;
      9875: inst = 32'h10408000;
      9876: inst = 32'hc4048ba;
      9877: inst = 32'h8220000;
      9878: inst = 32'h10408000;
      9879: inst = 32'hc4048bb;
      9880: inst = 32'h8220000;
      9881: inst = 32'h10408000;
      9882: inst = 32'hc4048bc;
      9883: inst = 32'h8220000;
      9884: inst = 32'h10408000;
      9885: inst = 32'hc4048bd;
      9886: inst = 32'h8220000;
      9887: inst = 32'h10408000;
      9888: inst = 32'hc4048be;
      9889: inst = 32'h8220000;
      9890: inst = 32'h10408000;
      9891: inst = 32'hc4048bf;
      9892: inst = 32'h8220000;
      9893: inst = 32'h10408000;
      9894: inst = 32'hc4048c0;
      9895: inst = 32'h8220000;
      9896: inst = 32'h10408000;
      9897: inst = 32'hc4048c1;
      9898: inst = 32'h8220000;
      9899: inst = 32'h10408000;
      9900: inst = 32'hc4048c2;
      9901: inst = 32'h8220000;
      9902: inst = 32'h10408000;
      9903: inst = 32'hc4048c3;
      9904: inst = 32'h8220000;
      9905: inst = 32'h10408000;
      9906: inst = 32'hc4048fc;
      9907: inst = 32'h8220000;
      9908: inst = 32'h10408000;
      9909: inst = 32'hc4048fd;
      9910: inst = 32'h8220000;
      9911: inst = 32'h10408000;
      9912: inst = 32'hc4048fe;
      9913: inst = 32'h8220000;
      9914: inst = 32'h10408000;
      9915: inst = 32'hc4048ff;
      9916: inst = 32'h8220000;
      9917: inst = 32'h10408000;
      9918: inst = 32'hc404900;
      9919: inst = 32'h8220000;
      9920: inst = 32'h10408000;
      9921: inst = 32'hc404901;
      9922: inst = 32'h8220000;
      9923: inst = 32'h10408000;
      9924: inst = 32'hc404902;
      9925: inst = 32'h8220000;
      9926: inst = 32'h10408000;
      9927: inst = 32'hc404903;
      9928: inst = 32'h8220000;
      9929: inst = 32'h10408000;
      9930: inst = 32'hc404904;
      9931: inst = 32'h8220000;
      9932: inst = 32'h10408000;
      9933: inst = 32'hc404905;
      9934: inst = 32'h8220000;
      9935: inst = 32'h10408000;
      9936: inst = 32'hc404906;
      9937: inst = 32'h8220000;
      9938: inst = 32'h10408000;
      9939: inst = 32'hc404907;
      9940: inst = 32'h8220000;
      9941: inst = 32'h10408000;
      9942: inst = 32'hc404908;
      9943: inst = 32'h8220000;
      9944: inst = 32'h10408000;
      9945: inst = 32'hc404909;
      9946: inst = 32'h8220000;
      9947: inst = 32'h10408000;
      9948: inst = 32'hc40490a;
      9949: inst = 32'h8220000;
      9950: inst = 32'h10408000;
      9951: inst = 32'hc40490b;
      9952: inst = 32'h8220000;
      9953: inst = 32'h10408000;
      9954: inst = 32'hc40490c;
      9955: inst = 32'h8220000;
      9956: inst = 32'h10408000;
      9957: inst = 32'hc40490d;
      9958: inst = 32'h8220000;
      9959: inst = 32'h10408000;
      9960: inst = 32'hc40490e;
      9961: inst = 32'h8220000;
      9962: inst = 32'h10408000;
      9963: inst = 32'hc40490f;
      9964: inst = 32'h8220000;
      9965: inst = 32'h10408000;
      9966: inst = 32'hc404910;
      9967: inst = 32'h8220000;
      9968: inst = 32'h10408000;
      9969: inst = 32'hc404911;
      9970: inst = 32'h8220000;
      9971: inst = 32'h10408000;
      9972: inst = 32'hc404912;
      9973: inst = 32'h8220000;
      9974: inst = 32'h10408000;
      9975: inst = 32'hc404913;
      9976: inst = 32'h8220000;
      9977: inst = 32'h10408000;
      9978: inst = 32'hc404914;
      9979: inst = 32'h8220000;
      9980: inst = 32'h10408000;
      9981: inst = 32'hc404915;
      9982: inst = 32'h8220000;
      9983: inst = 32'h10408000;
      9984: inst = 32'hc404916;
      9985: inst = 32'h8220000;
      9986: inst = 32'h10408000;
      9987: inst = 32'hc404917;
      9988: inst = 32'h8220000;
      9989: inst = 32'h10408000;
      9990: inst = 32'hc404918;
      9991: inst = 32'h8220000;
      9992: inst = 32'h10408000;
      9993: inst = 32'hc404919;
      9994: inst = 32'h8220000;
      9995: inst = 32'h10408000;
      9996: inst = 32'hc40491a;
      9997: inst = 32'h8220000;
      9998: inst = 32'h10408000;
      9999: inst = 32'hc40491b;
      10000: inst = 32'h8220000;
      10001: inst = 32'h10408000;
      10002: inst = 32'hc40491c;
      10003: inst = 32'h8220000;
      10004: inst = 32'h10408000;
      10005: inst = 32'hc40491d;
      10006: inst = 32'h8220000;
      10007: inst = 32'h10408000;
      10008: inst = 32'hc40491e;
      10009: inst = 32'h8220000;
      10010: inst = 32'h10408000;
      10011: inst = 32'hc40491f;
      10012: inst = 32'h8220000;
      10013: inst = 32'h10408000;
      10014: inst = 32'hc404920;
      10015: inst = 32'h8220000;
      10016: inst = 32'h10408000;
      10017: inst = 32'hc404921;
      10018: inst = 32'h8220000;
      10019: inst = 32'h10408000;
      10020: inst = 32'hc404922;
      10021: inst = 32'h8220000;
      10022: inst = 32'h10408000;
      10023: inst = 32'hc404923;
      10024: inst = 32'h8220000;
      10025: inst = 32'h10408000;
      10026: inst = 32'hc40495c;
      10027: inst = 32'h8220000;
      10028: inst = 32'h10408000;
      10029: inst = 32'hc40495d;
      10030: inst = 32'h8220000;
      10031: inst = 32'h10408000;
      10032: inst = 32'hc40495e;
      10033: inst = 32'h8220000;
      10034: inst = 32'h10408000;
      10035: inst = 32'hc40495f;
      10036: inst = 32'h8220000;
      10037: inst = 32'h10408000;
      10038: inst = 32'hc404960;
      10039: inst = 32'h8220000;
      10040: inst = 32'h10408000;
      10041: inst = 32'hc404961;
      10042: inst = 32'h8220000;
      10043: inst = 32'h10408000;
      10044: inst = 32'hc404962;
      10045: inst = 32'h8220000;
      10046: inst = 32'h10408000;
      10047: inst = 32'hc404963;
      10048: inst = 32'h8220000;
      10049: inst = 32'h10408000;
      10050: inst = 32'hc404964;
      10051: inst = 32'h8220000;
      10052: inst = 32'h10408000;
      10053: inst = 32'hc404965;
      10054: inst = 32'h8220000;
      10055: inst = 32'h10408000;
      10056: inst = 32'hc404966;
      10057: inst = 32'h8220000;
      10058: inst = 32'h10408000;
      10059: inst = 32'hc404967;
      10060: inst = 32'h8220000;
      10061: inst = 32'h10408000;
      10062: inst = 32'hc404968;
      10063: inst = 32'h8220000;
      10064: inst = 32'h10408000;
      10065: inst = 32'hc404969;
      10066: inst = 32'h8220000;
      10067: inst = 32'h10408000;
      10068: inst = 32'hc40496a;
      10069: inst = 32'h8220000;
      10070: inst = 32'h10408000;
      10071: inst = 32'hc40496b;
      10072: inst = 32'h8220000;
      10073: inst = 32'h10408000;
      10074: inst = 32'hc40496c;
      10075: inst = 32'h8220000;
      10076: inst = 32'h10408000;
      10077: inst = 32'hc40496d;
      10078: inst = 32'h8220000;
      10079: inst = 32'h10408000;
      10080: inst = 32'hc40496e;
      10081: inst = 32'h8220000;
      10082: inst = 32'h10408000;
      10083: inst = 32'hc40496f;
      10084: inst = 32'h8220000;
      10085: inst = 32'h10408000;
      10086: inst = 32'hc404970;
      10087: inst = 32'h8220000;
      10088: inst = 32'h10408000;
      10089: inst = 32'hc404971;
      10090: inst = 32'h8220000;
      10091: inst = 32'h10408000;
      10092: inst = 32'hc404972;
      10093: inst = 32'h8220000;
      10094: inst = 32'h10408000;
      10095: inst = 32'hc404973;
      10096: inst = 32'h8220000;
      10097: inst = 32'h10408000;
      10098: inst = 32'hc404974;
      10099: inst = 32'h8220000;
      10100: inst = 32'h10408000;
      10101: inst = 32'hc404975;
      10102: inst = 32'h8220000;
      10103: inst = 32'h10408000;
      10104: inst = 32'hc404976;
      10105: inst = 32'h8220000;
      10106: inst = 32'h10408000;
      10107: inst = 32'hc404977;
      10108: inst = 32'h8220000;
      10109: inst = 32'h10408000;
      10110: inst = 32'hc404978;
      10111: inst = 32'h8220000;
      10112: inst = 32'h10408000;
      10113: inst = 32'hc404979;
      10114: inst = 32'h8220000;
      10115: inst = 32'h10408000;
      10116: inst = 32'hc40497a;
      10117: inst = 32'h8220000;
      10118: inst = 32'h10408000;
      10119: inst = 32'hc40497b;
      10120: inst = 32'h8220000;
      10121: inst = 32'h10408000;
      10122: inst = 32'hc40497c;
      10123: inst = 32'h8220000;
      10124: inst = 32'h10408000;
      10125: inst = 32'hc40497d;
      10126: inst = 32'h8220000;
      10127: inst = 32'h10408000;
      10128: inst = 32'hc40497e;
      10129: inst = 32'h8220000;
      10130: inst = 32'h10408000;
      10131: inst = 32'hc40497f;
      10132: inst = 32'h8220000;
      10133: inst = 32'h10408000;
      10134: inst = 32'hc404980;
      10135: inst = 32'h8220000;
      10136: inst = 32'h10408000;
      10137: inst = 32'hc404981;
      10138: inst = 32'h8220000;
      10139: inst = 32'h10408000;
      10140: inst = 32'hc404982;
      10141: inst = 32'h8220000;
      10142: inst = 32'h10408000;
      10143: inst = 32'hc404983;
      10144: inst = 32'h8220000;
      10145: inst = 32'h10408000;
      10146: inst = 32'hc404992;
      10147: inst = 32'h8220000;
      10148: inst = 32'h10408000;
      10149: inst = 32'hc4049bc;
      10150: inst = 32'h8220000;
      10151: inst = 32'h10408000;
      10152: inst = 32'hc4049bd;
      10153: inst = 32'h8220000;
      10154: inst = 32'h10408000;
      10155: inst = 32'hc4049be;
      10156: inst = 32'h8220000;
      10157: inst = 32'h10408000;
      10158: inst = 32'hc4049bf;
      10159: inst = 32'h8220000;
      10160: inst = 32'h10408000;
      10161: inst = 32'hc4049c0;
      10162: inst = 32'h8220000;
      10163: inst = 32'h10408000;
      10164: inst = 32'hc4049c1;
      10165: inst = 32'h8220000;
      10166: inst = 32'h10408000;
      10167: inst = 32'hc4049c2;
      10168: inst = 32'h8220000;
      10169: inst = 32'h10408000;
      10170: inst = 32'hc4049c3;
      10171: inst = 32'h8220000;
      10172: inst = 32'h10408000;
      10173: inst = 32'hc4049c4;
      10174: inst = 32'h8220000;
      10175: inst = 32'h10408000;
      10176: inst = 32'hc4049c5;
      10177: inst = 32'h8220000;
      10178: inst = 32'h10408000;
      10179: inst = 32'hc4049c6;
      10180: inst = 32'h8220000;
      10181: inst = 32'h10408000;
      10182: inst = 32'hc4049c7;
      10183: inst = 32'h8220000;
      10184: inst = 32'h10408000;
      10185: inst = 32'hc4049c8;
      10186: inst = 32'h8220000;
      10187: inst = 32'h10408000;
      10188: inst = 32'hc4049c9;
      10189: inst = 32'h8220000;
      10190: inst = 32'h10408000;
      10191: inst = 32'hc4049ca;
      10192: inst = 32'h8220000;
      10193: inst = 32'h10408000;
      10194: inst = 32'hc4049cb;
      10195: inst = 32'h8220000;
      10196: inst = 32'h10408000;
      10197: inst = 32'hc4049cc;
      10198: inst = 32'h8220000;
      10199: inst = 32'h10408000;
      10200: inst = 32'hc4049cd;
      10201: inst = 32'h8220000;
      10202: inst = 32'h10408000;
      10203: inst = 32'hc4049ce;
      10204: inst = 32'h8220000;
      10205: inst = 32'h10408000;
      10206: inst = 32'hc4049cf;
      10207: inst = 32'h8220000;
      10208: inst = 32'h10408000;
      10209: inst = 32'hc4049d0;
      10210: inst = 32'h8220000;
      10211: inst = 32'h10408000;
      10212: inst = 32'hc4049d1;
      10213: inst = 32'h8220000;
      10214: inst = 32'h10408000;
      10215: inst = 32'hc4049d2;
      10216: inst = 32'h8220000;
      10217: inst = 32'h10408000;
      10218: inst = 32'hc4049d3;
      10219: inst = 32'h8220000;
      10220: inst = 32'h10408000;
      10221: inst = 32'hc4049d4;
      10222: inst = 32'h8220000;
      10223: inst = 32'h10408000;
      10224: inst = 32'hc4049d5;
      10225: inst = 32'h8220000;
      10226: inst = 32'h10408000;
      10227: inst = 32'hc4049d6;
      10228: inst = 32'h8220000;
      10229: inst = 32'h10408000;
      10230: inst = 32'hc4049d7;
      10231: inst = 32'h8220000;
      10232: inst = 32'h10408000;
      10233: inst = 32'hc4049d8;
      10234: inst = 32'h8220000;
      10235: inst = 32'h10408000;
      10236: inst = 32'hc4049d9;
      10237: inst = 32'h8220000;
      10238: inst = 32'h10408000;
      10239: inst = 32'hc4049da;
      10240: inst = 32'h8220000;
      10241: inst = 32'h10408000;
      10242: inst = 32'hc4049db;
      10243: inst = 32'h8220000;
      10244: inst = 32'h10408000;
      10245: inst = 32'hc4049dc;
      10246: inst = 32'h8220000;
      10247: inst = 32'h10408000;
      10248: inst = 32'hc4049dd;
      10249: inst = 32'h8220000;
      10250: inst = 32'h10408000;
      10251: inst = 32'hc4049de;
      10252: inst = 32'h8220000;
      10253: inst = 32'h10408000;
      10254: inst = 32'hc4049df;
      10255: inst = 32'h8220000;
      10256: inst = 32'h10408000;
      10257: inst = 32'hc4049e0;
      10258: inst = 32'h8220000;
      10259: inst = 32'h10408000;
      10260: inst = 32'hc4049e1;
      10261: inst = 32'h8220000;
      10262: inst = 32'h10408000;
      10263: inst = 32'hc4049e2;
      10264: inst = 32'h8220000;
      10265: inst = 32'h10408000;
      10266: inst = 32'hc4049e3;
      10267: inst = 32'h8220000;
      10268: inst = 32'h10408000;
      10269: inst = 32'hc4049f2;
      10270: inst = 32'h8220000;
      10271: inst = 32'h10408000;
      10272: inst = 32'hc404a1c;
      10273: inst = 32'h8220000;
      10274: inst = 32'h10408000;
      10275: inst = 32'hc404a1d;
      10276: inst = 32'h8220000;
      10277: inst = 32'h10408000;
      10278: inst = 32'hc404a1e;
      10279: inst = 32'h8220000;
      10280: inst = 32'h10408000;
      10281: inst = 32'hc404a1f;
      10282: inst = 32'h8220000;
      10283: inst = 32'h10408000;
      10284: inst = 32'hc404a20;
      10285: inst = 32'h8220000;
      10286: inst = 32'h10408000;
      10287: inst = 32'hc404a21;
      10288: inst = 32'h8220000;
      10289: inst = 32'h10408000;
      10290: inst = 32'hc404a22;
      10291: inst = 32'h8220000;
      10292: inst = 32'h10408000;
      10293: inst = 32'hc404a23;
      10294: inst = 32'h8220000;
      10295: inst = 32'h10408000;
      10296: inst = 32'hc404a24;
      10297: inst = 32'h8220000;
      10298: inst = 32'h10408000;
      10299: inst = 32'hc404a25;
      10300: inst = 32'h8220000;
      10301: inst = 32'h10408000;
      10302: inst = 32'hc404a26;
      10303: inst = 32'h8220000;
      10304: inst = 32'h10408000;
      10305: inst = 32'hc404a27;
      10306: inst = 32'h8220000;
      10307: inst = 32'h10408000;
      10308: inst = 32'hc404a28;
      10309: inst = 32'h8220000;
      10310: inst = 32'h10408000;
      10311: inst = 32'hc404a29;
      10312: inst = 32'h8220000;
      10313: inst = 32'h10408000;
      10314: inst = 32'hc404a2a;
      10315: inst = 32'h8220000;
      10316: inst = 32'h10408000;
      10317: inst = 32'hc404a2b;
      10318: inst = 32'h8220000;
      10319: inst = 32'h10408000;
      10320: inst = 32'hc404a2c;
      10321: inst = 32'h8220000;
      10322: inst = 32'h10408000;
      10323: inst = 32'hc404a2d;
      10324: inst = 32'h8220000;
      10325: inst = 32'h10408000;
      10326: inst = 32'hc404a2e;
      10327: inst = 32'h8220000;
      10328: inst = 32'h10408000;
      10329: inst = 32'hc404a2f;
      10330: inst = 32'h8220000;
      10331: inst = 32'h10408000;
      10332: inst = 32'hc404a30;
      10333: inst = 32'h8220000;
      10334: inst = 32'h10408000;
      10335: inst = 32'hc404a31;
      10336: inst = 32'h8220000;
      10337: inst = 32'h10408000;
      10338: inst = 32'hc404a32;
      10339: inst = 32'h8220000;
      10340: inst = 32'h10408000;
      10341: inst = 32'hc404a33;
      10342: inst = 32'h8220000;
      10343: inst = 32'h10408000;
      10344: inst = 32'hc404a34;
      10345: inst = 32'h8220000;
      10346: inst = 32'h10408000;
      10347: inst = 32'hc404a35;
      10348: inst = 32'h8220000;
      10349: inst = 32'h10408000;
      10350: inst = 32'hc404a36;
      10351: inst = 32'h8220000;
      10352: inst = 32'h10408000;
      10353: inst = 32'hc404a37;
      10354: inst = 32'h8220000;
      10355: inst = 32'h10408000;
      10356: inst = 32'hc404a38;
      10357: inst = 32'h8220000;
      10358: inst = 32'h10408000;
      10359: inst = 32'hc404a39;
      10360: inst = 32'h8220000;
      10361: inst = 32'h10408000;
      10362: inst = 32'hc404a3a;
      10363: inst = 32'h8220000;
      10364: inst = 32'h10408000;
      10365: inst = 32'hc404a3b;
      10366: inst = 32'h8220000;
      10367: inst = 32'h10408000;
      10368: inst = 32'hc404a3c;
      10369: inst = 32'h8220000;
      10370: inst = 32'h10408000;
      10371: inst = 32'hc404a3d;
      10372: inst = 32'h8220000;
      10373: inst = 32'h10408000;
      10374: inst = 32'hc404a3e;
      10375: inst = 32'h8220000;
      10376: inst = 32'h10408000;
      10377: inst = 32'hc404a3f;
      10378: inst = 32'h8220000;
      10379: inst = 32'h10408000;
      10380: inst = 32'hc404a40;
      10381: inst = 32'h8220000;
      10382: inst = 32'h10408000;
      10383: inst = 32'hc404a41;
      10384: inst = 32'h8220000;
      10385: inst = 32'h10408000;
      10386: inst = 32'hc404a42;
      10387: inst = 32'h8220000;
      10388: inst = 32'h10408000;
      10389: inst = 32'hc404a43;
      10390: inst = 32'h8220000;
      10391: inst = 32'h10408000;
      10392: inst = 32'hc404a52;
      10393: inst = 32'h8220000;
      10394: inst = 32'h10408000;
      10395: inst = 32'hc404a7c;
      10396: inst = 32'h8220000;
      10397: inst = 32'h10408000;
      10398: inst = 32'hc404a7d;
      10399: inst = 32'h8220000;
      10400: inst = 32'h10408000;
      10401: inst = 32'hc404a7e;
      10402: inst = 32'h8220000;
      10403: inst = 32'h10408000;
      10404: inst = 32'hc404a7f;
      10405: inst = 32'h8220000;
      10406: inst = 32'h10408000;
      10407: inst = 32'hc404a80;
      10408: inst = 32'h8220000;
      10409: inst = 32'h10408000;
      10410: inst = 32'hc404a81;
      10411: inst = 32'h8220000;
      10412: inst = 32'h10408000;
      10413: inst = 32'hc404a82;
      10414: inst = 32'h8220000;
      10415: inst = 32'h10408000;
      10416: inst = 32'hc404a83;
      10417: inst = 32'h8220000;
      10418: inst = 32'h10408000;
      10419: inst = 32'hc404a84;
      10420: inst = 32'h8220000;
      10421: inst = 32'h10408000;
      10422: inst = 32'hc404a85;
      10423: inst = 32'h8220000;
      10424: inst = 32'h10408000;
      10425: inst = 32'hc404a86;
      10426: inst = 32'h8220000;
      10427: inst = 32'h10408000;
      10428: inst = 32'hc404a87;
      10429: inst = 32'h8220000;
      10430: inst = 32'h10408000;
      10431: inst = 32'hc404a88;
      10432: inst = 32'h8220000;
      10433: inst = 32'h10408000;
      10434: inst = 32'hc404a89;
      10435: inst = 32'h8220000;
      10436: inst = 32'h10408000;
      10437: inst = 32'hc404a8a;
      10438: inst = 32'h8220000;
      10439: inst = 32'h10408000;
      10440: inst = 32'hc404a8b;
      10441: inst = 32'h8220000;
      10442: inst = 32'h10408000;
      10443: inst = 32'hc404a8c;
      10444: inst = 32'h8220000;
      10445: inst = 32'h10408000;
      10446: inst = 32'hc404a8d;
      10447: inst = 32'h8220000;
      10448: inst = 32'h10408000;
      10449: inst = 32'hc404a8e;
      10450: inst = 32'h8220000;
      10451: inst = 32'h10408000;
      10452: inst = 32'hc404a8f;
      10453: inst = 32'h8220000;
      10454: inst = 32'h10408000;
      10455: inst = 32'hc404a90;
      10456: inst = 32'h8220000;
      10457: inst = 32'h10408000;
      10458: inst = 32'hc404a91;
      10459: inst = 32'h8220000;
      10460: inst = 32'h10408000;
      10461: inst = 32'hc404a92;
      10462: inst = 32'h8220000;
      10463: inst = 32'h10408000;
      10464: inst = 32'hc404a93;
      10465: inst = 32'h8220000;
      10466: inst = 32'h10408000;
      10467: inst = 32'hc404a94;
      10468: inst = 32'h8220000;
      10469: inst = 32'h10408000;
      10470: inst = 32'hc404a95;
      10471: inst = 32'h8220000;
      10472: inst = 32'h10408000;
      10473: inst = 32'hc404a96;
      10474: inst = 32'h8220000;
      10475: inst = 32'h10408000;
      10476: inst = 32'hc404a97;
      10477: inst = 32'h8220000;
      10478: inst = 32'h10408000;
      10479: inst = 32'hc404a98;
      10480: inst = 32'h8220000;
      10481: inst = 32'h10408000;
      10482: inst = 32'hc404a99;
      10483: inst = 32'h8220000;
      10484: inst = 32'h10408000;
      10485: inst = 32'hc404a9a;
      10486: inst = 32'h8220000;
      10487: inst = 32'h10408000;
      10488: inst = 32'hc404a9b;
      10489: inst = 32'h8220000;
      10490: inst = 32'h10408000;
      10491: inst = 32'hc404a9c;
      10492: inst = 32'h8220000;
      10493: inst = 32'h10408000;
      10494: inst = 32'hc404a9d;
      10495: inst = 32'h8220000;
      10496: inst = 32'h10408000;
      10497: inst = 32'hc404a9e;
      10498: inst = 32'h8220000;
      10499: inst = 32'h10408000;
      10500: inst = 32'hc404a9f;
      10501: inst = 32'h8220000;
      10502: inst = 32'h10408000;
      10503: inst = 32'hc404aa0;
      10504: inst = 32'h8220000;
      10505: inst = 32'h10408000;
      10506: inst = 32'hc404aa1;
      10507: inst = 32'h8220000;
      10508: inst = 32'h10408000;
      10509: inst = 32'hc404aa2;
      10510: inst = 32'h8220000;
      10511: inst = 32'h10408000;
      10512: inst = 32'hc404aa3;
      10513: inst = 32'h8220000;
      10514: inst = 32'h10408000;
      10515: inst = 32'hc404ab4;
      10516: inst = 32'h8220000;
      10517: inst = 32'h10408000;
      10518: inst = 32'hc404adc;
      10519: inst = 32'h8220000;
      10520: inst = 32'h10408000;
      10521: inst = 32'hc404add;
      10522: inst = 32'h8220000;
      10523: inst = 32'h10408000;
      10524: inst = 32'hc404ade;
      10525: inst = 32'h8220000;
      10526: inst = 32'h10408000;
      10527: inst = 32'hc404adf;
      10528: inst = 32'h8220000;
      10529: inst = 32'h10408000;
      10530: inst = 32'hc404ae0;
      10531: inst = 32'h8220000;
      10532: inst = 32'h10408000;
      10533: inst = 32'hc404ae1;
      10534: inst = 32'h8220000;
      10535: inst = 32'h10408000;
      10536: inst = 32'hc404ae2;
      10537: inst = 32'h8220000;
      10538: inst = 32'h10408000;
      10539: inst = 32'hc404ae3;
      10540: inst = 32'h8220000;
      10541: inst = 32'h10408000;
      10542: inst = 32'hc404ae4;
      10543: inst = 32'h8220000;
      10544: inst = 32'h10408000;
      10545: inst = 32'hc404ae5;
      10546: inst = 32'h8220000;
      10547: inst = 32'h10408000;
      10548: inst = 32'hc404ae6;
      10549: inst = 32'h8220000;
      10550: inst = 32'h10408000;
      10551: inst = 32'hc404ae7;
      10552: inst = 32'h8220000;
      10553: inst = 32'h10408000;
      10554: inst = 32'hc404ae8;
      10555: inst = 32'h8220000;
      10556: inst = 32'h10408000;
      10557: inst = 32'hc404ae9;
      10558: inst = 32'h8220000;
      10559: inst = 32'h10408000;
      10560: inst = 32'hc404aea;
      10561: inst = 32'h8220000;
      10562: inst = 32'h10408000;
      10563: inst = 32'hc404aeb;
      10564: inst = 32'h8220000;
      10565: inst = 32'h10408000;
      10566: inst = 32'hc404aec;
      10567: inst = 32'h8220000;
      10568: inst = 32'h10408000;
      10569: inst = 32'hc404aed;
      10570: inst = 32'h8220000;
      10571: inst = 32'h10408000;
      10572: inst = 32'hc404aee;
      10573: inst = 32'h8220000;
      10574: inst = 32'h10408000;
      10575: inst = 32'hc404aef;
      10576: inst = 32'h8220000;
      10577: inst = 32'h10408000;
      10578: inst = 32'hc404af0;
      10579: inst = 32'h8220000;
      10580: inst = 32'h10408000;
      10581: inst = 32'hc404af1;
      10582: inst = 32'h8220000;
      10583: inst = 32'h10408000;
      10584: inst = 32'hc404af2;
      10585: inst = 32'h8220000;
      10586: inst = 32'h10408000;
      10587: inst = 32'hc404af3;
      10588: inst = 32'h8220000;
      10589: inst = 32'h10408000;
      10590: inst = 32'hc404af4;
      10591: inst = 32'h8220000;
      10592: inst = 32'h10408000;
      10593: inst = 32'hc404af5;
      10594: inst = 32'h8220000;
      10595: inst = 32'h10408000;
      10596: inst = 32'hc404af6;
      10597: inst = 32'h8220000;
      10598: inst = 32'h10408000;
      10599: inst = 32'hc404af7;
      10600: inst = 32'h8220000;
      10601: inst = 32'h10408000;
      10602: inst = 32'hc404af8;
      10603: inst = 32'h8220000;
      10604: inst = 32'h10408000;
      10605: inst = 32'hc404af9;
      10606: inst = 32'h8220000;
      10607: inst = 32'h10408000;
      10608: inst = 32'hc404afa;
      10609: inst = 32'h8220000;
      10610: inst = 32'h10408000;
      10611: inst = 32'hc404afb;
      10612: inst = 32'h8220000;
      10613: inst = 32'h10408000;
      10614: inst = 32'hc404afc;
      10615: inst = 32'h8220000;
      10616: inst = 32'h10408000;
      10617: inst = 32'hc404afd;
      10618: inst = 32'h8220000;
      10619: inst = 32'h10408000;
      10620: inst = 32'hc404afe;
      10621: inst = 32'h8220000;
      10622: inst = 32'h10408000;
      10623: inst = 32'hc404aff;
      10624: inst = 32'h8220000;
      10625: inst = 32'h10408000;
      10626: inst = 32'hc404b00;
      10627: inst = 32'h8220000;
      10628: inst = 32'h10408000;
      10629: inst = 32'hc404b01;
      10630: inst = 32'h8220000;
      10631: inst = 32'h10408000;
      10632: inst = 32'hc404b02;
      10633: inst = 32'h8220000;
      10634: inst = 32'h10408000;
      10635: inst = 32'hc404b03;
      10636: inst = 32'h8220000;
      10637: inst = 32'h10408000;
      10638: inst = 32'hc404b14;
      10639: inst = 32'h8220000;
      10640: inst = 32'h10408000;
      10641: inst = 32'hc404b3c;
      10642: inst = 32'h8220000;
      10643: inst = 32'h10408000;
      10644: inst = 32'hc404b3d;
      10645: inst = 32'h8220000;
      10646: inst = 32'h10408000;
      10647: inst = 32'hc404b3e;
      10648: inst = 32'h8220000;
      10649: inst = 32'h10408000;
      10650: inst = 32'hc404b3f;
      10651: inst = 32'h8220000;
      10652: inst = 32'h10408000;
      10653: inst = 32'hc404b40;
      10654: inst = 32'h8220000;
      10655: inst = 32'h10408000;
      10656: inst = 32'hc404b41;
      10657: inst = 32'h8220000;
      10658: inst = 32'h10408000;
      10659: inst = 32'hc404b42;
      10660: inst = 32'h8220000;
      10661: inst = 32'h10408000;
      10662: inst = 32'hc404b43;
      10663: inst = 32'h8220000;
      10664: inst = 32'h10408000;
      10665: inst = 32'hc404b44;
      10666: inst = 32'h8220000;
      10667: inst = 32'h10408000;
      10668: inst = 32'hc404b45;
      10669: inst = 32'h8220000;
      10670: inst = 32'h10408000;
      10671: inst = 32'hc404b46;
      10672: inst = 32'h8220000;
      10673: inst = 32'h10408000;
      10674: inst = 32'hc404b47;
      10675: inst = 32'h8220000;
      10676: inst = 32'h10408000;
      10677: inst = 32'hc404b48;
      10678: inst = 32'h8220000;
      10679: inst = 32'h10408000;
      10680: inst = 32'hc404b49;
      10681: inst = 32'h8220000;
      10682: inst = 32'h10408000;
      10683: inst = 32'hc404b4a;
      10684: inst = 32'h8220000;
      10685: inst = 32'h10408000;
      10686: inst = 32'hc404b4b;
      10687: inst = 32'h8220000;
      10688: inst = 32'h10408000;
      10689: inst = 32'hc404b4c;
      10690: inst = 32'h8220000;
      10691: inst = 32'h10408000;
      10692: inst = 32'hc404b4d;
      10693: inst = 32'h8220000;
      10694: inst = 32'h10408000;
      10695: inst = 32'hc404b4e;
      10696: inst = 32'h8220000;
      10697: inst = 32'h10408000;
      10698: inst = 32'hc404b4f;
      10699: inst = 32'h8220000;
      10700: inst = 32'h10408000;
      10701: inst = 32'hc404b50;
      10702: inst = 32'h8220000;
      10703: inst = 32'h10408000;
      10704: inst = 32'hc404b51;
      10705: inst = 32'h8220000;
      10706: inst = 32'h10408000;
      10707: inst = 32'hc404b52;
      10708: inst = 32'h8220000;
      10709: inst = 32'h10408000;
      10710: inst = 32'hc404b53;
      10711: inst = 32'h8220000;
      10712: inst = 32'h10408000;
      10713: inst = 32'hc404b54;
      10714: inst = 32'h8220000;
      10715: inst = 32'h10408000;
      10716: inst = 32'hc404b55;
      10717: inst = 32'h8220000;
      10718: inst = 32'h10408000;
      10719: inst = 32'hc404b56;
      10720: inst = 32'h8220000;
      10721: inst = 32'h10408000;
      10722: inst = 32'hc404b57;
      10723: inst = 32'h8220000;
      10724: inst = 32'h10408000;
      10725: inst = 32'hc404b58;
      10726: inst = 32'h8220000;
      10727: inst = 32'h10408000;
      10728: inst = 32'hc404b59;
      10729: inst = 32'h8220000;
      10730: inst = 32'h10408000;
      10731: inst = 32'hc404b5a;
      10732: inst = 32'h8220000;
      10733: inst = 32'h10408000;
      10734: inst = 32'hc404b5b;
      10735: inst = 32'h8220000;
      10736: inst = 32'h10408000;
      10737: inst = 32'hc404b5c;
      10738: inst = 32'h8220000;
      10739: inst = 32'h10408000;
      10740: inst = 32'hc404b5d;
      10741: inst = 32'h8220000;
      10742: inst = 32'h10408000;
      10743: inst = 32'hc404b5e;
      10744: inst = 32'h8220000;
      10745: inst = 32'h10408000;
      10746: inst = 32'hc404b5f;
      10747: inst = 32'h8220000;
      10748: inst = 32'h10408000;
      10749: inst = 32'hc404b60;
      10750: inst = 32'h8220000;
      10751: inst = 32'h10408000;
      10752: inst = 32'hc404b61;
      10753: inst = 32'h8220000;
      10754: inst = 32'h10408000;
      10755: inst = 32'hc404b62;
      10756: inst = 32'h8220000;
      10757: inst = 32'h10408000;
      10758: inst = 32'hc404b63;
      10759: inst = 32'h8220000;
      10760: inst = 32'h10408000;
      10761: inst = 32'hc404b9c;
      10762: inst = 32'h8220000;
      10763: inst = 32'h10408000;
      10764: inst = 32'hc404b9d;
      10765: inst = 32'h8220000;
      10766: inst = 32'h10408000;
      10767: inst = 32'hc404b9e;
      10768: inst = 32'h8220000;
      10769: inst = 32'h10408000;
      10770: inst = 32'hc404b9f;
      10771: inst = 32'h8220000;
      10772: inst = 32'h10408000;
      10773: inst = 32'hc404ba0;
      10774: inst = 32'h8220000;
      10775: inst = 32'h10408000;
      10776: inst = 32'hc404ba1;
      10777: inst = 32'h8220000;
      10778: inst = 32'h10408000;
      10779: inst = 32'hc404ba2;
      10780: inst = 32'h8220000;
      10781: inst = 32'h10408000;
      10782: inst = 32'hc404ba3;
      10783: inst = 32'h8220000;
      10784: inst = 32'h10408000;
      10785: inst = 32'hc404ba4;
      10786: inst = 32'h8220000;
      10787: inst = 32'h10408000;
      10788: inst = 32'hc404ba5;
      10789: inst = 32'h8220000;
      10790: inst = 32'h10408000;
      10791: inst = 32'hc404ba6;
      10792: inst = 32'h8220000;
      10793: inst = 32'h10408000;
      10794: inst = 32'hc404ba7;
      10795: inst = 32'h8220000;
      10796: inst = 32'h10408000;
      10797: inst = 32'hc404ba8;
      10798: inst = 32'h8220000;
      10799: inst = 32'h10408000;
      10800: inst = 32'hc404ba9;
      10801: inst = 32'h8220000;
      10802: inst = 32'h10408000;
      10803: inst = 32'hc404baa;
      10804: inst = 32'h8220000;
      10805: inst = 32'h10408000;
      10806: inst = 32'hc404bab;
      10807: inst = 32'h8220000;
      10808: inst = 32'h10408000;
      10809: inst = 32'hc404bac;
      10810: inst = 32'h8220000;
      10811: inst = 32'h10408000;
      10812: inst = 32'hc404bad;
      10813: inst = 32'h8220000;
      10814: inst = 32'h10408000;
      10815: inst = 32'hc404bae;
      10816: inst = 32'h8220000;
      10817: inst = 32'h10408000;
      10818: inst = 32'hc404baf;
      10819: inst = 32'h8220000;
      10820: inst = 32'h10408000;
      10821: inst = 32'hc404bb0;
      10822: inst = 32'h8220000;
      10823: inst = 32'h10408000;
      10824: inst = 32'hc404bb1;
      10825: inst = 32'h8220000;
      10826: inst = 32'h10408000;
      10827: inst = 32'hc404bb2;
      10828: inst = 32'h8220000;
      10829: inst = 32'h10408000;
      10830: inst = 32'hc404bb3;
      10831: inst = 32'h8220000;
      10832: inst = 32'h10408000;
      10833: inst = 32'hc404bb4;
      10834: inst = 32'h8220000;
      10835: inst = 32'h10408000;
      10836: inst = 32'hc404bb5;
      10837: inst = 32'h8220000;
      10838: inst = 32'h10408000;
      10839: inst = 32'hc404bb6;
      10840: inst = 32'h8220000;
      10841: inst = 32'h10408000;
      10842: inst = 32'hc404bb7;
      10843: inst = 32'h8220000;
      10844: inst = 32'h10408000;
      10845: inst = 32'hc404bb8;
      10846: inst = 32'h8220000;
      10847: inst = 32'h10408000;
      10848: inst = 32'hc404bb9;
      10849: inst = 32'h8220000;
      10850: inst = 32'h10408000;
      10851: inst = 32'hc404bba;
      10852: inst = 32'h8220000;
      10853: inst = 32'h10408000;
      10854: inst = 32'hc404bbb;
      10855: inst = 32'h8220000;
      10856: inst = 32'h10408000;
      10857: inst = 32'hc404bbc;
      10858: inst = 32'h8220000;
      10859: inst = 32'h10408000;
      10860: inst = 32'hc404bbd;
      10861: inst = 32'h8220000;
      10862: inst = 32'h10408000;
      10863: inst = 32'hc404bbe;
      10864: inst = 32'h8220000;
      10865: inst = 32'h10408000;
      10866: inst = 32'hc404bbf;
      10867: inst = 32'h8220000;
      10868: inst = 32'h10408000;
      10869: inst = 32'hc404bc0;
      10870: inst = 32'h8220000;
      10871: inst = 32'h10408000;
      10872: inst = 32'hc404bc1;
      10873: inst = 32'h8220000;
      10874: inst = 32'h10408000;
      10875: inst = 32'hc404bc2;
      10876: inst = 32'h8220000;
      10877: inst = 32'h10408000;
      10878: inst = 32'hc404bc3;
      10879: inst = 32'h8220000;
      10880: inst = 32'hc20ee75;
      10881: inst = 32'h10408000;
      10882: inst = 32'hc4042ea;
      10883: inst = 32'h8220000;
      10884: inst = 32'h10408000;
      10885: inst = 32'hc4043a7;
      10886: inst = 32'h8220000;
      10887: inst = 32'hc20d42c;
      10888: inst = 32'h10408000;
      10889: inst = 32'hc4042eb;
      10890: inst = 32'h8220000;
      10891: inst = 32'h10408000;
      10892: inst = 32'hc4042ec;
      10893: inst = 32'h8220000;
      10894: inst = 32'h10408000;
      10895: inst = 32'hc4043a8;
      10896: inst = 32'h8220000;
      10897: inst = 32'hc20ee55;
      10898: inst = 32'h10408000;
      10899: inst = 32'hc4042ed;
      10900: inst = 32'h8220000;
      10901: inst = 32'h10408000;
      10902: inst = 32'hc4043b0;
      10903: inst = 32'h8220000;
      10904: inst = 32'hc20e571;
      10905: inst = 32'h10408000;
      10906: inst = 32'hc404349;
      10907: inst = 32'h8220000;
      10908: inst = 32'h10408000;
      10909: inst = 32'hc40434e;
      10910: inst = 32'h8220000;
      10911: inst = 32'h10408000;
      10912: inst = 32'hc404406;
      10913: inst = 32'h8220000;
      10914: inst = 32'h10408000;
      10915: inst = 32'hc404411;
      10916: inst = 32'h8220000;
      10917: inst = 32'hc20cb28;
      10918: inst = 32'h10408000;
      10919: inst = 32'hc40434a;
      10920: inst = 32'h8220000;
      10921: inst = 32'h10408000;
      10922: inst = 32'hc40434d;
      10923: inst = 32'h8220000;
      10924: inst = 32'h10408000;
      10925: inst = 32'hc404407;
      10926: inst = 32'h8220000;
      10927: inst = 32'h10408000;
      10928: inst = 32'hc404410;
      10929: inst = 32'h8220000;
      10930: inst = 32'hc20cac7;
      10931: inst = 32'h10408000;
      10932: inst = 32'hc40434b;
      10933: inst = 32'h8220000;
      10934: inst = 32'h10408000;
      10935: inst = 32'hc40434c;
      10936: inst = 32'h8220000;
      10937: inst = 32'h10408000;
      10938: inst = 32'hc4043a9;
      10939: inst = 32'h8220000;
      10940: inst = 32'h10408000;
      10941: inst = 32'hc4043aa;
      10942: inst = 32'h8220000;
      10943: inst = 32'h10408000;
      10944: inst = 32'hc4043ab;
      10945: inst = 32'h8220000;
      10946: inst = 32'h10408000;
      10947: inst = 32'hc4043ac;
      10948: inst = 32'h8220000;
      10949: inst = 32'h10408000;
      10950: inst = 32'hc4043ad;
      10951: inst = 32'h8220000;
      10952: inst = 32'h10408000;
      10953: inst = 32'hc4043ae;
      10954: inst = 32'h8220000;
      10955: inst = 32'h10408000;
      10956: inst = 32'hc404408;
      10957: inst = 32'h8220000;
      10958: inst = 32'h10408000;
      10959: inst = 32'hc404409;
      10960: inst = 32'h8220000;
      10961: inst = 32'h10408000;
      10962: inst = 32'hc40440a;
      10963: inst = 32'h8220000;
      10964: inst = 32'h10408000;
      10965: inst = 32'hc40440b;
      10966: inst = 32'h8220000;
      10967: inst = 32'h10408000;
      10968: inst = 32'hc40440c;
      10969: inst = 32'h8220000;
      10970: inst = 32'h10408000;
      10971: inst = 32'hc40440d;
      10972: inst = 32'h8220000;
      10973: inst = 32'h10408000;
      10974: inst = 32'hc40440e;
      10975: inst = 32'h8220000;
      10976: inst = 32'h10408000;
      10977: inst = 32'hc40440f;
      10978: inst = 32'h8220000;
      10979: inst = 32'hc20d40c;
      10980: inst = 32'h10408000;
      10981: inst = 32'hc4043af;
      10982: inst = 32'h8220000;
      10983: inst = 32'hc20ee8e;
      10984: inst = 32'h10408000;
      10985: inst = 32'hc40446a;
      10986: inst = 32'h8220000;
      10987: inst = 32'h10408000;
      10988: inst = 32'hc4044b5;
      10989: inst = 32'h8220000;
      10990: inst = 32'hc20ee48;
      10991: inst = 32'h10408000;
      10992: inst = 32'hc40446b;
      10993: inst = 32'h8220000;
      10994: inst = 32'h10408000;
      10995: inst = 32'hc40446c;
      10996: inst = 32'h8220000;
      10997: inst = 32'h10408000;
      10998: inst = 32'hc4044b3;
      10999: inst = 32'h8220000;
      11000: inst = 32'h10408000;
      11001: inst = 32'hc4044b4;
      11002: inst = 32'h8220000;
      11003: inst = 32'hc20ee90;
      11004: inst = 32'h10408000;
      11005: inst = 32'hc40446d;
      11006: inst = 32'h8220000;
      11007: inst = 32'h10408000;
      11008: inst = 32'hc4044b2;
      11009: inst = 32'h8220000;
      11010: inst = 32'hc20eeb5;
      11011: inst = 32'h10408000;
      11012: inst = 32'hc4044cb;
      11013: inst = 32'h8220000;
      11014: inst = 32'h10408000;
      11015: inst = 32'hc4044cc;
      11016: inst = 32'h8220000;
      11017: inst = 32'h10408000;
      11018: inst = 32'hc404513;
      11019: inst = 32'h8220000;
      11020: inst = 32'h10408000;
      11021: inst = 32'hc404514;
      11022: inst = 32'h8220000;
      11023: inst = 32'hc20c2e2;
      11024: inst = 32'h10408000;
      11025: inst = 32'hc4046ef;
      11026: inst = 32'h8220000;
      11027: inst = 32'h10408000;
      11028: inst = 32'hc4046f0;
      11029: inst = 32'h8220000;
      11030: inst = 32'h10408000;
      11031: inst = 32'hc4046f1;
      11032: inst = 32'h8220000;
      11033: inst = 32'h10408000;
      11034: inst = 32'hc4046f2;
      11035: inst = 32'h8220000;
      11036: inst = 32'h10408000;
      11037: inst = 32'hc4046f3;
      11038: inst = 32'h8220000;
      11039: inst = 32'h10408000;
      11040: inst = 32'hc4046f4;
      11041: inst = 32'h8220000;
      11042: inst = 32'h10408000;
      11043: inst = 32'hc4046f5;
      11044: inst = 32'h8220000;
      11045: inst = 32'h10408000;
      11046: inst = 32'hc4046f6;
      11047: inst = 32'h8220000;
      11048: inst = 32'h10408000;
      11049: inst = 32'hc4046f7;
      11050: inst = 32'h8220000;
      11051: inst = 32'h10408000;
      11052: inst = 32'hc4046f8;
      11053: inst = 32'h8220000;
      11054: inst = 32'h10408000;
      11055: inst = 32'hc4046f9;
      11056: inst = 32'h8220000;
      11057: inst = 32'h10408000;
      11058: inst = 32'hc4046fa;
      11059: inst = 32'h8220000;
      11060: inst = 32'h10408000;
      11061: inst = 32'hc4046fb;
      11062: inst = 32'h8220000;
      11063: inst = 32'h10408000;
      11064: inst = 32'hc4046fc;
      11065: inst = 32'h8220000;
      11066: inst = 32'h10408000;
      11067: inst = 32'hc4046fd;
      11068: inst = 32'h8220000;
      11069: inst = 32'h10408000;
      11070: inst = 32'hc4046fe;
      11071: inst = 32'h8220000;
      11072: inst = 32'h10408000;
      11073: inst = 32'hc4046ff;
      11074: inst = 32'h8220000;
      11075: inst = 32'h10408000;
      11076: inst = 32'hc40474f;
      11077: inst = 32'h8220000;
      11078: inst = 32'h10408000;
      11079: inst = 32'hc40475f;
      11080: inst = 32'h8220000;
      11081: inst = 32'h10408000;
      11082: inst = 32'hc4047af;
      11083: inst = 32'h8220000;
      11084: inst = 32'h10408000;
      11085: inst = 32'hc4047bf;
      11086: inst = 32'h8220000;
      11087: inst = 32'h10408000;
      11088: inst = 32'hc40480f;
      11089: inst = 32'h8220000;
      11090: inst = 32'h10408000;
      11091: inst = 32'hc40481f;
      11092: inst = 32'h8220000;
      11093: inst = 32'h10408000;
      11094: inst = 32'hc40486f;
      11095: inst = 32'h8220000;
      11096: inst = 32'h10408000;
      11097: inst = 32'hc40487f;
      11098: inst = 32'h8220000;
      11099: inst = 32'h10408000;
      11100: inst = 32'hc4048cf;
      11101: inst = 32'h8220000;
      11102: inst = 32'h10408000;
      11103: inst = 32'hc4048df;
      11104: inst = 32'h8220000;
      11105: inst = 32'h10408000;
      11106: inst = 32'hc40492f;
      11107: inst = 32'h8220000;
      11108: inst = 32'h10408000;
      11109: inst = 32'hc40493f;
      11110: inst = 32'h8220000;
      11111: inst = 32'h10408000;
      11112: inst = 32'hc40498f;
      11113: inst = 32'h8220000;
      11114: inst = 32'h10408000;
      11115: inst = 32'hc40499f;
      11116: inst = 32'h8220000;
      11117: inst = 32'h10408000;
      11118: inst = 32'hc4049ef;
      11119: inst = 32'h8220000;
      11120: inst = 32'h10408000;
      11121: inst = 32'hc4049ff;
      11122: inst = 32'h8220000;
      11123: inst = 32'h10408000;
      11124: inst = 32'hc404a4f;
      11125: inst = 32'h8220000;
      11126: inst = 32'h10408000;
      11127: inst = 32'hc404a5f;
      11128: inst = 32'h8220000;
      11129: inst = 32'h10408000;
      11130: inst = 32'hc404aaf;
      11131: inst = 32'h8220000;
      11132: inst = 32'h10408000;
      11133: inst = 32'hc404abf;
      11134: inst = 32'h8220000;
      11135: inst = 32'h10408000;
      11136: inst = 32'hc404b0f;
      11137: inst = 32'h8220000;
      11138: inst = 32'h10408000;
      11139: inst = 32'hc404b1f;
      11140: inst = 32'h8220000;
      11141: inst = 32'h10408000;
      11142: inst = 32'hc404b6f;
      11143: inst = 32'h8220000;
      11144: inst = 32'h10408000;
      11145: inst = 32'hc404b7f;
      11146: inst = 32'h8220000;
      11147: inst = 32'h10408000;
      11148: inst = 32'hc404bcf;
      11149: inst = 32'h8220000;
      11150: inst = 32'h10408000;
      11151: inst = 32'hc404bdf;
      11152: inst = 32'h8220000;
      11153: inst = 32'h10408000;
      11154: inst = 32'hc404c2f;
      11155: inst = 32'h8220000;
      11156: inst = 32'h10408000;
      11157: inst = 32'hc404c3f;
      11158: inst = 32'h8220000;
      11159: inst = 32'h10408000;
      11160: inst = 32'hc404c8f;
      11161: inst = 32'h8220000;
      11162: inst = 32'h10408000;
      11163: inst = 32'hc404c9f;
      11164: inst = 32'h8220000;
      11165: inst = 32'h10408000;
      11166: inst = 32'hc404cef;
      11167: inst = 32'h8220000;
      11168: inst = 32'h10408000;
      11169: inst = 32'hc404cff;
      11170: inst = 32'h8220000;
      11171: inst = 32'h10408000;
      11172: inst = 32'hc404d4f;
      11173: inst = 32'h8220000;
      11174: inst = 32'h10408000;
      11175: inst = 32'hc404d5f;
      11176: inst = 32'h8220000;
      11177: inst = 32'h10408000;
      11178: inst = 32'hc404daf;
      11179: inst = 32'h8220000;
      11180: inst = 32'h10408000;
      11181: inst = 32'hc404dbf;
      11182: inst = 32'h8220000;
      11183: inst = 32'h10408000;
      11184: inst = 32'hc404e0f;
      11185: inst = 32'h8220000;
      11186: inst = 32'h10408000;
      11187: inst = 32'hc404e1f;
      11188: inst = 32'h8220000;
      11189: inst = 32'h10408000;
      11190: inst = 32'hc404e6f;
      11191: inst = 32'h8220000;
      11192: inst = 32'h10408000;
      11193: inst = 32'hc404e7f;
      11194: inst = 32'h8220000;
      11195: inst = 32'h10408000;
      11196: inst = 32'hc404ecf;
      11197: inst = 32'h8220000;
      11198: inst = 32'h10408000;
      11199: inst = 32'hc404edf;
      11200: inst = 32'h8220000;
      11201: inst = 32'h10408000;
      11202: inst = 32'hc404f2f;
      11203: inst = 32'h8220000;
      11204: inst = 32'h10408000;
      11205: inst = 32'hc404f3f;
      11206: inst = 32'h8220000;
      11207: inst = 32'h10408000;
      11208: inst = 32'hc404f8f;
      11209: inst = 32'h8220000;
      11210: inst = 32'h10408000;
      11211: inst = 32'hc404f9f;
      11212: inst = 32'h8220000;
      11213: inst = 32'h10408000;
      11214: inst = 32'hc404fef;
      11215: inst = 32'h8220000;
      11216: inst = 32'h10408000;
      11217: inst = 32'hc404fff;
      11218: inst = 32'h8220000;
      11219: inst = 32'h10408000;
      11220: inst = 32'hc40504f;
      11221: inst = 32'h8220000;
      11222: inst = 32'h10408000;
      11223: inst = 32'hc40505f;
      11224: inst = 32'h8220000;
      11225: inst = 32'h10408000;
      11226: inst = 32'hc4050af;
      11227: inst = 32'h8220000;
      11228: inst = 32'h10408000;
      11229: inst = 32'hc4050bf;
      11230: inst = 32'h8220000;
      11231: inst = 32'h10408000;
      11232: inst = 32'hc40510f;
      11233: inst = 32'h8220000;
      11234: inst = 32'h10408000;
      11235: inst = 32'hc40511f;
      11236: inst = 32'h8220000;
      11237: inst = 32'h10408000;
      11238: inst = 32'hc40516f;
      11239: inst = 32'h8220000;
      11240: inst = 32'h10408000;
      11241: inst = 32'hc40517f;
      11242: inst = 32'h8220000;
      11243: inst = 32'h10408000;
      11244: inst = 32'hc4051cf;
      11245: inst = 32'h8220000;
      11246: inst = 32'h10408000;
      11247: inst = 32'hc4051df;
      11248: inst = 32'h8220000;
      11249: inst = 32'h10408000;
      11250: inst = 32'hc40522f;
      11251: inst = 32'h8220000;
      11252: inst = 32'h10408000;
      11253: inst = 32'hc40523f;
      11254: inst = 32'h8220000;
      11255: inst = 32'h10408000;
      11256: inst = 32'hc40528f;
      11257: inst = 32'h8220000;
      11258: inst = 32'h10408000;
      11259: inst = 32'hc40529f;
      11260: inst = 32'h8220000;
      11261: inst = 32'h10408000;
      11262: inst = 32'hc4052ef;
      11263: inst = 32'h8220000;
      11264: inst = 32'h10408000;
      11265: inst = 32'hc4052f0;
      11266: inst = 32'h8220000;
      11267: inst = 32'h10408000;
      11268: inst = 32'hc4052f1;
      11269: inst = 32'h8220000;
      11270: inst = 32'h10408000;
      11271: inst = 32'hc4052f2;
      11272: inst = 32'h8220000;
      11273: inst = 32'h10408000;
      11274: inst = 32'hc4052f3;
      11275: inst = 32'h8220000;
      11276: inst = 32'h10408000;
      11277: inst = 32'hc4052f4;
      11278: inst = 32'h8220000;
      11279: inst = 32'h10408000;
      11280: inst = 32'hc4052f5;
      11281: inst = 32'h8220000;
      11282: inst = 32'h10408000;
      11283: inst = 32'hc4052f6;
      11284: inst = 32'h8220000;
      11285: inst = 32'h10408000;
      11286: inst = 32'hc4052f7;
      11287: inst = 32'h8220000;
      11288: inst = 32'h10408000;
      11289: inst = 32'hc4052f8;
      11290: inst = 32'h8220000;
      11291: inst = 32'h10408000;
      11292: inst = 32'hc4052f9;
      11293: inst = 32'h8220000;
      11294: inst = 32'h10408000;
      11295: inst = 32'hc4052fa;
      11296: inst = 32'h8220000;
      11297: inst = 32'h10408000;
      11298: inst = 32'hc4052fb;
      11299: inst = 32'h8220000;
      11300: inst = 32'h10408000;
      11301: inst = 32'hc4052fc;
      11302: inst = 32'h8220000;
      11303: inst = 32'h10408000;
      11304: inst = 32'hc4052fd;
      11305: inst = 32'h8220000;
      11306: inst = 32'h10408000;
      11307: inst = 32'hc4052fe;
      11308: inst = 32'h8220000;
      11309: inst = 32'h10408000;
      11310: inst = 32'hc4052ff;
      11311: inst = 32'h8220000;
      11312: inst = 32'hc20dbc5;
      11313: inst = 32'h10408000;
      11314: inst = 32'hc404750;
      11315: inst = 32'h8220000;
      11316: inst = 32'h10408000;
      11317: inst = 32'hc404751;
      11318: inst = 32'h8220000;
      11319: inst = 32'h10408000;
      11320: inst = 32'hc404752;
      11321: inst = 32'h8220000;
      11322: inst = 32'h10408000;
      11323: inst = 32'hc404753;
      11324: inst = 32'h8220000;
      11325: inst = 32'h10408000;
      11326: inst = 32'hc404754;
      11327: inst = 32'h8220000;
      11328: inst = 32'h10408000;
      11329: inst = 32'hc404755;
      11330: inst = 32'h8220000;
      11331: inst = 32'h10408000;
      11332: inst = 32'hc404756;
      11333: inst = 32'h8220000;
      11334: inst = 32'h10408000;
      11335: inst = 32'hc404757;
      11336: inst = 32'h8220000;
      11337: inst = 32'h10408000;
      11338: inst = 32'hc404758;
      11339: inst = 32'h8220000;
      11340: inst = 32'h10408000;
      11341: inst = 32'hc404759;
      11342: inst = 32'h8220000;
      11343: inst = 32'h10408000;
      11344: inst = 32'hc40475a;
      11345: inst = 32'h8220000;
      11346: inst = 32'h10408000;
      11347: inst = 32'hc40475b;
      11348: inst = 32'h8220000;
      11349: inst = 32'h10408000;
      11350: inst = 32'hc40475c;
      11351: inst = 32'h8220000;
      11352: inst = 32'h10408000;
      11353: inst = 32'hc40475d;
      11354: inst = 32'h8220000;
      11355: inst = 32'h10408000;
      11356: inst = 32'hc40475e;
      11357: inst = 32'h8220000;
      11358: inst = 32'h10408000;
      11359: inst = 32'hc4047b0;
      11360: inst = 32'h8220000;
      11361: inst = 32'h10408000;
      11362: inst = 32'hc4047b1;
      11363: inst = 32'h8220000;
      11364: inst = 32'h10408000;
      11365: inst = 32'hc4047b2;
      11366: inst = 32'h8220000;
      11367: inst = 32'h10408000;
      11368: inst = 32'hc4047b3;
      11369: inst = 32'h8220000;
      11370: inst = 32'h10408000;
      11371: inst = 32'hc4047b4;
      11372: inst = 32'h8220000;
      11373: inst = 32'h10408000;
      11374: inst = 32'hc4047b5;
      11375: inst = 32'h8220000;
      11376: inst = 32'h10408000;
      11377: inst = 32'hc4047b6;
      11378: inst = 32'h8220000;
      11379: inst = 32'h10408000;
      11380: inst = 32'hc4047b7;
      11381: inst = 32'h8220000;
      11382: inst = 32'h10408000;
      11383: inst = 32'hc4047b8;
      11384: inst = 32'h8220000;
      11385: inst = 32'h10408000;
      11386: inst = 32'hc4047b9;
      11387: inst = 32'h8220000;
      11388: inst = 32'h10408000;
      11389: inst = 32'hc4047ba;
      11390: inst = 32'h8220000;
      11391: inst = 32'h10408000;
      11392: inst = 32'hc4047bb;
      11393: inst = 32'h8220000;
      11394: inst = 32'h10408000;
      11395: inst = 32'hc4047bc;
      11396: inst = 32'h8220000;
      11397: inst = 32'h10408000;
      11398: inst = 32'hc4047bd;
      11399: inst = 32'h8220000;
      11400: inst = 32'h10408000;
      11401: inst = 32'hc4047be;
      11402: inst = 32'h8220000;
      11403: inst = 32'h10408000;
      11404: inst = 32'hc404810;
      11405: inst = 32'h8220000;
      11406: inst = 32'h10408000;
      11407: inst = 32'hc404811;
      11408: inst = 32'h8220000;
      11409: inst = 32'h10408000;
      11410: inst = 32'hc404812;
      11411: inst = 32'h8220000;
      11412: inst = 32'h10408000;
      11413: inst = 32'hc404813;
      11414: inst = 32'h8220000;
      11415: inst = 32'h10408000;
      11416: inst = 32'hc404814;
      11417: inst = 32'h8220000;
      11418: inst = 32'h10408000;
      11419: inst = 32'hc404815;
      11420: inst = 32'h8220000;
      11421: inst = 32'h10408000;
      11422: inst = 32'hc404816;
      11423: inst = 32'h8220000;
      11424: inst = 32'h10408000;
      11425: inst = 32'hc404817;
      11426: inst = 32'h8220000;
      11427: inst = 32'h10408000;
      11428: inst = 32'hc404818;
      11429: inst = 32'h8220000;
      11430: inst = 32'h10408000;
      11431: inst = 32'hc404819;
      11432: inst = 32'h8220000;
      11433: inst = 32'h10408000;
      11434: inst = 32'hc40481a;
      11435: inst = 32'h8220000;
      11436: inst = 32'h10408000;
      11437: inst = 32'hc40481b;
      11438: inst = 32'h8220000;
      11439: inst = 32'h10408000;
      11440: inst = 32'hc40481c;
      11441: inst = 32'h8220000;
      11442: inst = 32'h10408000;
      11443: inst = 32'hc40481d;
      11444: inst = 32'h8220000;
      11445: inst = 32'h10408000;
      11446: inst = 32'hc40481e;
      11447: inst = 32'h8220000;
      11448: inst = 32'h10408000;
      11449: inst = 32'hc404870;
      11450: inst = 32'h8220000;
      11451: inst = 32'h10408000;
      11452: inst = 32'hc404871;
      11453: inst = 32'h8220000;
      11454: inst = 32'h10408000;
      11455: inst = 32'hc404872;
      11456: inst = 32'h8220000;
      11457: inst = 32'h10408000;
      11458: inst = 32'hc404873;
      11459: inst = 32'h8220000;
      11460: inst = 32'h10408000;
      11461: inst = 32'hc404874;
      11462: inst = 32'h8220000;
      11463: inst = 32'h10408000;
      11464: inst = 32'hc404875;
      11465: inst = 32'h8220000;
      11466: inst = 32'h10408000;
      11467: inst = 32'hc404876;
      11468: inst = 32'h8220000;
      11469: inst = 32'h10408000;
      11470: inst = 32'hc404877;
      11471: inst = 32'h8220000;
      11472: inst = 32'h10408000;
      11473: inst = 32'hc404878;
      11474: inst = 32'h8220000;
      11475: inst = 32'h10408000;
      11476: inst = 32'hc404879;
      11477: inst = 32'h8220000;
      11478: inst = 32'h10408000;
      11479: inst = 32'hc40487a;
      11480: inst = 32'h8220000;
      11481: inst = 32'h10408000;
      11482: inst = 32'hc40487b;
      11483: inst = 32'h8220000;
      11484: inst = 32'h10408000;
      11485: inst = 32'hc40487c;
      11486: inst = 32'h8220000;
      11487: inst = 32'h10408000;
      11488: inst = 32'hc40487d;
      11489: inst = 32'h8220000;
      11490: inst = 32'h10408000;
      11491: inst = 32'hc40487e;
      11492: inst = 32'h8220000;
      11493: inst = 32'h10408000;
      11494: inst = 32'hc4048d0;
      11495: inst = 32'h8220000;
      11496: inst = 32'h10408000;
      11497: inst = 32'hc4048d1;
      11498: inst = 32'h8220000;
      11499: inst = 32'h10408000;
      11500: inst = 32'hc4048d2;
      11501: inst = 32'h8220000;
      11502: inst = 32'h10408000;
      11503: inst = 32'hc4048d3;
      11504: inst = 32'h8220000;
      11505: inst = 32'h10408000;
      11506: inst = 32'hc4048d4;
      11507: inst = 32'h8220000;
      11508: inst = 32'h10408000;
      11509: inst = 32'hc4048d5;
      11510: inst = 32'h8220000;
      11511: inst = 32'h10408000;
      11512: inst = 32'hc4048d6;
      11513: inst = 32'h8220000;
      11514: inst = 32'h10408000;
      11515: inst = 32'hc4048d7;
      11516: inst = 32'h8220000;
      11517: inst = 32'h10408000;
      11518: inst = 32'hc4048d8;
      11519: inst = 32'h8220000;
      11520: inst = 32'h10408000;
      11521: inst = 32'hc4048d9;
      11522: inst = 32'h8220000;
      11523: inst = 32'h10408000;
      11524: inst = 32'hc4048da;
      11525: inst = 32'h8220000;
      11526: inst = 32'h10408000;
      11527: inst = 32'hc4048db;
      11528: inst = 32'h8220000;
      11529: inst = 32'h10408000;
      11530: inst = 32'hc4048dc;
      11531: inst = 32'h8220000;
      11532: inst = 32'h10408000;
      11533: inst = 32'hc4048dd;
      11534: inst = 32'h8220000;
      11535: inst = 32'h10408000;
      11536: inst = 32'hc4048de;
      11537: inst = 32'h8220000;
      11538: inst = 32'h10408000;
      11539: inst = 32'hc404930;
      11540: inst = 32'h8220000;
      11541: inst = 32'h10408000;
      11542: inst = 32'hc404931;
      11543: inst = 32'h8220000;
      11544: inst = 32'h10408000;
      11545: inst = 32'hc404936;
      11546: inst = 32'h8220000;
      11547: inst = 32'h10408000;
      11548: inst = 32'hc404937;
      11549: inst = 32'h8220000;
      11550: inst = 32'h10408000;
      11551: inst = 32'hc404938;
      11552: inst = 32'h8220000;
      11553: inst = 32'h10408000;
      11554: inst = 32'hc404939;
      11555: inst = 32'h8220000;
      11556: inst = 32'h10408000;
      11557: inst = 32'hc40493a;
      11558: inst = 32'h8220000;
      11559: inst = 32'h10408000;
      11560: inst = 32'hc40493b;
      11561: inst = 32'h8220000;
      11562: inst = 32'h10408000;
      11563: inst = 32'hc40493c;
      11564: inst = 32'h8220000;
      11565: inst = 32'h10408000;
      11566: inst = 32'hc40493d;
      11567: inst = 32'h8220000;
      11568: inst = 32'h10408000;
      11569: inst = 32'hc40493e;
      11570: inst = 32'h8220000;
      11571: inst = 32'h10408000;
      11572: inst = 32'hc404990;
      11573: inst = 32'h8220000;
      11574: inst = 32'h10408000;
      11575: inst = 32'hc404991;
      11576: inst = 32'h8220000;
      11577: inst = 32'h10408000;
      11578: inst = 32'hc404996;
      11579: inst = 32'h8220000;
      11580: inst = 32'h10408000;
      11581: inst = 32'hc404997;
      11582: inst = 32'h8220000;
      11583: inst = 32'h10408000;
      11584: inst = 32'hc404998;
      11585: inst = 32'h8220000;
      11586: inst = 32'h10408000;
      11587: inst = 32'hc404999;
      11588: inst = 32'h8220000;
      11589: inst = 32'h10408000;
      11590: inst = 32'hc40499a;
      11591: inst = 32'h8220000;
      11592: inst = 32'h10408000;
      11593: inst = 32'hc40499b;
      11594: inst = 32'h8220000;
      11595: inst = 32'h10408000;
      11596: inst = 32'hc40499c;
      11597: inst = 32'h8220000;
      11598: inst = 32'h10408000;
      11599: inst = 32'hc40499d;
      11600: inst = 32'h8220000;
      11601: inst = 32'h10408000;
      11602: inst = 32'hc40499e;
      11603: inst = 32'h8220000;
      11604: inst = 32'h10408000;
      11605: inst = 32'hc4049f0;
      11606: inst = 32'h8220000;
      11607: inst = 32'h10408000;
      11608: inst = 32'hc4049f1;
      11609: inst = 32'h8220000;
      11610: inst = 32'h10408000;
      11611: inst = 32'hc4049f6;
      11612: inst = 32'h8220000;
      11613: inst = 32'h10408000;
      11614: inst = 32'hc4049f7;
      11615: inst = 32'h8220000;
      11616: inst = 32'h10408000;
      11617: inst = 32'hc4049f8;
      11618: inst = 32'h8220000;
      11619: inst = 32'h10408000;
      11620: inst = 32'hc4049f9;
      11621: inst = 32'h8220000;
      11622: inst = 32'h10408000;
      11623: inst = 32'hc4049fa;
      11624: inst = 32'h8220000;
      11625: inst = 32'h10408000;
      11626: inst = 32'hc4049fb;
      11627: inst = 32'h8220000;
      11628: inst = 32'h10408000;
      11629: inst = 32'hc4049fc;
      11630: inst = 32'h8220000;
      11631: inst = 32'h10408000;
      11632: inst = 32'hc4049fd;
      11633: inst = 32'h8220000;
      11634: inst = 32'h10408000;
      11635: inst = 32'hc4049fe;
      11636: inst = 32'h8220000;
      11637: inst = 32'h10408000;
      11638: inst = 32'hc404a50;
      11639: inst = 32'h8220000;
      11640: inst = 32'h10408000;
      11641: inst = 32'hc404a51;
      11642: inst = 32'h8220000;
      11643: inst = 32'h10408000;
      11644: inst = 32'hc404a56;
      11645: inst = 32'h8220000;
      11646: inst = 32'h10408000;
      11647: inst = 32'hc404a57;
      11648: inst = 32'h8220000;
      11649: inst = 32'h10408000;
      11650: inst = 32'hc404a58;
      11651: inst = 32'h8220000;
      11652: inst = 32'h10408000;
      11653: inst = 32'hc404a59;
      11654: inst = 32'h8220000;
      11655: inst = 32'h10408000;
      11656: inst = 32'hc404a5a;
      11657: inst = 32'h8220000;
      11658: inst = 32'h10408000;
      11659: inst = 32'hc404a5b;
      11660: inst = 32'h8220000;
      11661: inst = 32'h10408000;
      11662: inst = 32'hc404a5c;
      11663: inst = 32'h8220000;
      11664: inst = 32'h10408000;
      11665: inst = 32'hc404a5d;
      11666: inst = 32'h8220000;
      11667: inst = 32'h10408000;
      11668: inst = 32'hc404a5e;
      11669: inst = 32'h8220000;
      11670: inst = 32'h10408000;
      11671: inst = 32'hc404ab0;
      11672: inst = 32'h8220000;
      11673: inst = 32'h10408000;
      11674: inst = 32'hc404ab1;
      11675: inst = 32'h8220000;
      11676: inst = 32'h10408000;
      11677: inst = 32'hc404ab6;
      11678: inst = 32'h8220000;
      11679: inst = 32'h10408000;
      11680: inst = 32'hc404ab7;
      11681: inst = 32'h8220000;
      11682: inst = 32'h10408000;
      11683: inst = 32'hc404ab8;
      11684: inst = 32'h8220000;
      11685: inst = 32'h10408000;
      11686: inst = 32'hc404ab9;
      11687: inst = 32'h8220000;
      11688: inst = 32'h10408000;
      11689: inst = 32'hc404aba;
      11690: inst = 32'h8220000;
      11691: inst = 32'h10408000;
      11692: inst = 32'hc404abb;
      11693: inst = 32'h8220000;
      11694: inst = 32'h10408000;
      11695: inst = 32'hc404abc;
      11696: inst = 32'h8220000;
      11697: inst = 32'h10408000;
      11698: inst = 32'hc404abd;
      11699: inst = 32'h8220000;
      11700: inst = 32'h10408000;
      11701: inst = 32'hc404abe;
      11702: inst = 32'h8220000;
      11703: inst = 32'h10408000;
      11704: inst = 32'hc404b10;
      11705: inst = 32'h8220000;
      11706: inst = 32'h10408000;
      11707: inst = 32'hc404b11;
      11708: inst = 32'h8220000;
      11709: inst = 32'h10408000;
      11710: inst = 32'hc404b16;
      11711: inst = 32'h8220000;
      11712: inst = 32'h10408000;
      11713: inst = 32'hc404b17;
      11714: inst = 32'h8220000;
      11715: inst = 32'h10408000;
      11716: inst = 32'hc404b18;
      11717: inst = 32'h8220000;
      11718: inst = 32'h10408000;
      11719: inst = 32'hc404b19;
      11720: inst = 32'h8220000;
      11721: inst = 32'h10408000;
      11722: inst = 32'hc404b1a;
      11723: inst = 32'h8220000;
      11724: inst = 32'h10408000;
      11725: inst = 32'hc404b1b;
      11726: inst = 32'h8220000;
      11727: inst = 32'h10408000;
      11728: inst = 32'hc404b1c;
      11729: inst = 32'h8220000;
      11730: inst = 32'h10408000;
      11731: inst = 32'hc404b1d;
      11732: inst = 32'h8220000;
      11733: inst = 32'h10408000;
      11734: inst = 32'hc404b1e;
      11735: inst = 32'h8220000;
      11736: inst = 32'h10408000;
      11737: inst = 32'hc404b70;
      11738: inst = 32'h8220000;
      11739: inst = 32'h10408000;
      11740: inst = 32'hc404b71;
      11741: inst = 32'h8220000;
      11742: inst = 32'h10408000;
      11743: inst = 32'hc404b76;
      11744: inst = 32'h8220000;
      11745: inst = 32'h10408000;
      11746: inst = 32'hc404b77;
      11747: inst = 32'h8220000;
      11748: inst = 32'h10408000;
      11749: inst = 32'hc404b78;
      11750: inst = 32'h8220000;
      11751: inst = 32'h10408000;
      11752: inst = 32'hc404b79;
      11753: inst = 32'h8220000;
      11754: inst = 32'h10408000;
      11755: inst = 32'hc404b7a;
      11756: inst = 32'h8220000;
      11757: inst = 32'h10408000;
      11758: inst = 32'hc404b7b;
      11759: inst = 32'h8220000;
      11760: inst = 32'h10408000;
      11761: inst = 32'hc404b7c;
      11762: inst = 32'h8220000;
      11763: inst = 32'h10408000;
      11764: inst = 32'hc404b7d;
      11765: inst = 32'h8220000;
      11766: inst = 32'h10408000;
      11767: inst = 32'hc404b7e;
      11768: inst = 32'h8220000;
      11769: inst = 32'h10408000;
      11770: inst = 32'hc404bd0;
      11771: inst = 32'h8220000;
      11772: inst = 32'h10408000;
      11773: inst = 32'hc404bd1;
      11774: inst = 32'h8220000;
      11775: inst = 32'h10408000;
      11776: inst = 32'hc404bd2;
      11777: inst = 32'h8220000;
      11778: inst = 32'h10408000;
      11779: inst = 32'hc404bd3;
      11780: inst = 32'h8220000;
      11781: inst = 32'h10408000;
      11782: inst = 32'hc404bd4;
      11783: inst = 32'h8220000;
      11784: inst = 32'h10408000;
      11785: inst = 32'hc404bd5;
      11786: inst = 32'h8220000;
      11787: inst = 32'h10408000;
      11788: inst = 32'hc404bd6;
      11789: inst = 32'h8220000;
      11790: inst = 32'h10408000;
      11791: inst = 32'hc404bd7;
      11792: inst = 32'h8220000;
      11793: inst = 32'h10408000;
      11794: inst = 32'hc404bd8;
      11795: inst = 32'h8220000;
      11796: inst = 32'h10408000;
      11797: inst = 32'hc404bd9;
      11798: inst = 32'h8220000;
      11799: inst = 32'h10408000;
      11800: inst = 32'hc404bda;
      11801: inst = 32'h8220000;
      11802: inst = 32'h10408000;
      11803: inst = 32'hc404bdb;
      11804: inst = 32'h8220000;
      11805: inst = 32'h10408000;
      11806: inst = 32'hc404bdc;
      11807: inst = 32'h8220000;
      11808: inst = 32'h10408000;
      11809: inst = 32'hc404bdd;
      11810: inst = 32'h8220000;
      11811: inst = 32'h10408000;
      11812: inst = 32'hc404bde;
      11813: inst = 32'h8220000;
      11814: inst = 32'h10408000;
      11815: inst = 32'hc404c30;
      11816: inst = 32'h8220000;
      11817: inst = 32'h10408000;
      11818: inst = 32'hc404c31;
      11819: inst = 32'h8220000;
      11820: inst = 32'h10408000;
      11821: inst = 32'hc404c32;
      11822: inst = 32'h8220000;
      11823: inst = 32'h10408000;
      11824: inst = 32'hc404c33;
      11825: inst = 32'h8220000;
      11826: inst = 32'h10408000;
      11827: inst = 32'hc404c34;
      11828: inst = 32'h8220000;
      11829: inst = 32'h10408000;
      11830: inst = 32'hc404c35;
      11831: inst = 32'h8220000;
      11832: inst = 32'h10408000;
      11833: inst = 32'hc404c36;
      11834: inst = 32'h8220000;
      11835: inst = 32'h10408000;
      11836: inst = 32'hc404c37;
      11837: inst = 32'h8220000;
      11838: inst = 32'h10408000;
      11839: inst = 32'hc404c38;
      11840: inst = 32'h8220000;
      11841: inst = 32'h10408000;
      11842: inst = 32'hc404c39;
      11843: inst = 32'h8220000;
      11844: inst = 32'h10408000;
      11845: inst = 32'hc404c3a;
      11846: inst = 32'h8220000;
      11847: inst = 32'h10408000;
      11848: inst = 32'hc404c3b;
      11849: inst = 32'h8220000;
      11850: inst = 32'h10408000;
      11851: inst = 32'hc404c3c;
      11852: inst = 32'h8220000;
      11853: inst = 32'h10408000;
      11854: inst = 32'hc404c3d;
      11855: inst = 32'h8220000;
      11856: inst = 32'h10408000;
      11857: inst = 32'hc404c3e;
      11858: inst = 32'h8220000;
      11859: inst = 32'h10408000;
      11860: inst = 32'hc404c90;
      11861: inst = 32'h8220000;
      11862: inst = 32'h10408000;
      11863: inst = 32'hc404c91;
      11864: inst = 32'h8220000;
      11865: inst = 32'h10408000;
      11866: inst = 32'hc404c92;
      11867: inst = 32'h8220000;
      11868: inst = 32'h10408000;
      11869: inst = 32'hc404c93;
      11870: inst = 32'h8220000;
      11871: inst = 32'h10408000;
      11872: inst = 32'hc404c94;
      11873: inst = 32'h8220000;
      11874: inst = 32'h10408000;
      11875: inst = 32'hc404c95;
      11876: inst = 32'h8220000;
      11877: inst = 32'h10408000;
      11878: inst = 32'hc404c96;
      11879: inst = 32'h8220000;
      11880: inst = 32'h10408000;
      11881: inst = 32'hc404c97;
      11882: inst = 32'h8220000;
      11883: inst = 32'h10408000;
      11884: inst = 32'hc404c98;
      11885: inst = 32'h8220000;
      11886: inst = 32'h10408000;
      11887: inst = 32'hc404c99;
      11888: inst = 32'h8220000;
      11889: inst = 32'h10408000;
      11890: inst = 32'hc404c9a;
      11891: inst = 32'h8220000;
      11892: inst = 32'h10408000;
      11893: inst = 32'hc404c9b;
      11894: inst = 32'h8220000;
      11895: inst = 32'h10408000;
      11896: inst = 32'hc404c9c;
      11897: inst = 32'h8220000;
      11898: inst = 32'h10408000;
      11899: inst = 32'hc404c9d;
      11900: inst = 32'h8220000;
      11901: inst = 32'h10408000;
      11902: inst = 32'hc404c9e;
      11903: inst = 32'h8220000;
      11904: inst = 32'h10408000;
      11905: inst = 32'hc404cf0;
      11906: inst = 32'h8220000;
      11907: inst = 32'h10408000;
      11908: inst = 32'hc404cf1;
      11909: inst = 32'h8220000;
      11910: inst = 32'h10408000;
      11911: inst = 32'hc404cf2;
      11912: inst = 32'h8220000;
      11913: inst = 32'h10408000;
      11914: inst = 32'hc404cf3;
      11915: inst = 32'h8220000;
      11916: inst = 32'h10408000;
      11917: inst = 32'hc404cf4;
      11918: inst = 32'h8220000;
      11919: inst = 32'h10408000;
      11920: inst = 32'hc404cf5;
      11921: inst = 32'h8220000;
      11922: inst = 32'h10408000;
      11923: inst = 32'hc404cf6;
      11924: inst = 32'h8220000;
      11925: inst = 32'h10408000;
      11926: inst = 32'hc404cf7;
      11927: inst = 32'h8220000;
      11928: inst = 32'h10408000;
      11929: inst = 32'hc404cf8;
      11930: inst = 32'h8220000;
      11931: inst = 32'h10408000;
      11932: inst = 32'hc404cf9;
      11933: inst = 32'h8220000;
      11934: inst = 32'h10408000;
      11935: inst = 32'hc404cfa;
      11936: inst = 32'h8220000;
      11937: inst = 32'h10408000;
      11938: inst = 32'hc404cfe;
      11939: inst = 32'h8220000;
      11940: inst = 32'h10408000;
      11941: inst = 32'hc404d50;
      11942: inst = 32'h8220000;
      11943: inst = 32'h10408000;
      11944: inst = 32'hc404d51;
      11945: inst = 32'h8220000;
      11946: inst = 32'h10408000;
      11947: inst = 32'hc404d52;
      11948: inst = 32'h8220000;
      11949: inst = 32'h10408000;
      11950: inst = 32'hc404d53;
      11951: inst = 32'h8220000;
      11952: inst = 32'h10408000;
      11953: inst = 32'hc404d54;
      11954: inst = 32'h8220000;
      11955: inst = 32'h10408000;
      11956: inst = 32'hc404d55;
      11957: inst = 32'h8220000;
      11958: inst = 32'h10408000;
      11959: inst = 32'hc404d56;
      11960: inst = 32'h8220000;
      11961: inst = 32'h10408000;
      11962: inst = 32'hc404d57;
      11963: inst = 32'h8220000;
      11964: inst = 32'h10408000;
      11965: inst = 32'hc404d58;
      11966: inst = 32'h8220000;
      11967: inst = 32'h10408000;
      11968: inst = 32'hc404d59;
      11969: inst = 32'h8220000;
      11970: inst = 32'h10408000;
      11971: inst = 32'hc404d5a;
      11972: inst = 32'h8220000;
      11973: inst = 32'h10408000;
      11974: inst = 32'hc404d5c;
      11975: inst = 32'h8220000;
      11976: inst = 32'h10408000;
      11977: inst = 32'hc404d5d;
      11978: inst = 32'h8220000;
      11979: inst = 32'h10408000;
      11980: inst = 32'hc404d5e;
      11981: inst = 32'h8220000;
      11982: inst = 32'h10408000;
      11983: inst = 32'hc404db0;
      11984: inst = 32'h8220000;
      11985: inst = 32'h10408000;
      11986: inst = 32'hc404db1;
      11987: inst = 32'h8220000;
      11988: inst = 32'h10408000;
      11989: inst = 32'hc404db2;
      11990: inst = 32'h8220000;
      11991: inst = 32'h10408000;
      11992: inst = 32'hc404db3;
      11993: inst = 32'h8220000;
      11994: inst = 32'h10408000;
      11995: inst = 32'hc404db4;
      11996: inst = 32'h8220000;
      11997: inst = 32'h10408000;
      11998: inst = 32'hc404db5;
      11999: inst = 32'h8220000;
      12000: inst = 32'h10408000;
      12001: inst = 32'hc404db6;
      12002: inst = 32'h8220000;
      12003: inst = 32'h10408000;
      12004: inst = 32'hc404db7;
      12005: inst = 32'h8220000;
      12006: inst = 32'h10408000;
      12007: inst = 32'hc404db8;
      12008: inst = 32'h8220000;
      12009: inst = 32'h10408000;
      12010: inst = 32'hc404db9;
      12011: inst = 32'h8220000;
      12012: inst = 32'h10408000;
      12013: inst = 32'hc404dba;
      12014: inst = 32'h8220000;
      12015: inst = 32'h10408000;
      12016: inst = 32'hc404dbb;
      12017: inst = 32'h8220000;
      12018: inst = 32'h10408000;
      12019: inst = 32'hc404dbc;
      12020: inst = 32'h8220000;
      12021: inst = 32'h10408000;
      12022: inst = 32'hc404dbd;
      12023: inst = 32'h8220000;
      12024: inst = 32'h10408000;
      12025: inst = 32'hc404dbe;
      12026: inst = 32'h8220000;
      12027: inst = 32'h10408000;
      12028: inst = 32'hc404e10;
      12029: inst = 32'h8220000;
      12030: inst = 32'h10408000;
      12031: inst = 32'hc404e11;
      12032: inst = 32'h8220000;
      12033: inst = 32'h10408000;
      12034: inst = 32'hc404e12;
      12035: inst = 32'h8220000;
      12036: inst = 32'h10408000;
      12037: inst = 32'hc404e13;
      12038: inst = 32'h8220000;
      12039: inst = 32'h10408000;
      12040: inst = 32'hc404e14;
      12041: inst = 32'h8220000;
      12042: inst = 32'h10408000;
      12043: inst = 32'hc404e15;
      12044: inst = 32'h8220000;
      12045: inst = 32'h10408000;
      12046: inst = 32'hc404e16;
      12047: inst = 32'h8220000;
      12048: inst = 32'h10408000;
      12049: inst = 32'hc404e17;
      12050: inst = 32'h8220000;
      12051: inst = 32'h10408000;
      12052: inst = 32'hc404e18;
      12053: inst = 32'h8220000;
      12054: inst = 32'h10408000;
      12055: inst = 32'hc404e19;
      12056: inst = 32'h8220000;
      12057: inst = 32'h10408000;
      12058: inst = 32'hc404e1a;
      12059: inst = 32'h8220000;
      12060: inst = 32'h10408000;
      12061: inst = 32'hc404e1b;
      12062: inst = 32'h8220000;
      12063: inst = 32'h10408000;
      12064: inst = 32'hc404e1c;
      12065: inst = 32'h8220000;
      12066: inst = 32'h10408000;
      12067: inst = 32'hc404e1d;
      12068: inst = 32'h8220000;
      12069: inst = 32'h10408000;
      12070: inst = 32'hc404e1e;
      12071: inst = 32'h8220000;
      12072: inst = 32'h10408000;
      12073: inst = 32'hc404e70;
      12074: inst = 32'h8220000;
      12075: inst = 32'h10408000;
      12076: inst = 32'hc404e71;
      12077: inst = 32'h8220000;
      12078: inst = 32'h10408000;
      12079: inst = 32'hc404e72;
      12080: inst = 32'h8220000;
      12081: inst = 32'h10408000;
      12082: inst = 32'hc404e73;
      12083: inst = 32'h8220000;
      12084: inst = 32'h10408000;
      12085: inst = 32'hc404e74;
      12086: inst = 32'h8220000;
      12087: inst = 32'h10408000;
      12088: inst = 32'hc404e75;
      12089: inst = 32'h8220000;
      12090: inst = 32'h10408000;
      12091: inst = 32'hc404e76;
      12092: inst = 32'h8220000;
      12093: inst = 32'h10408000;
      12094: inst = 32'hc404e77;
      12095: inst = 32'h8220000;
      12096: inst = 32'h10408000;
      12097: inst = 32'hc404e78;
      12098: inst = 32'h8220000;
      12099: inst = 32'h10408000;
      12100: inst = 32'hc404e79;
      12101: inst = 32'h8220000;
      12102: inst = 32'h10408000;
      12103: inst = 32'hc404e7a;
      12104: inst = 32'h8220000;
      12105: inst = 32'h10408000;
      12106: inst = 32'hc404e7b;
      12107: inst = 32'h8220000;
      12108: inst = 32'h10408000;
      12109: inst = 32'hc404e7c;
      12110: inst = 32'h8220000;
      12111: inst = 32'h10408000;
      12112: inst = 32'hc404e7d;
      12113: inst = 32'h8220000;
      12114: inst = 32'h10408000;
      12115: inst = 32'hc404e7e;
      12116: inst = 32'h8220000;
      12117: inst = 32'h10408000;
      12118: inst = 32'hc404ed0;
      12119: inst = 32'h8220000;
      12120: inst = 32'h10408000;
      12121: inst = 32'hc404ed1;
      12122: inst = 32'h8220000;
      12123: inst = 32'h10408000;
      12124: inst = 32'hc404ed2;
      12125: inst = 32'h8220000;
      12126: inst = 32'h10408000;
      12127: inst = 32'hc404ed3;
      12128: inst = 32'h8220000;
      12129: inst = 32'h10408000;
      12130: inst = 32'hc404ed4;
      12131: inst = 32'h8220000;
      12132: inst = 32'h10408000;
      12133: inst = 32'hc404ed5;
      12134: inst = 32'h8220000;
      12135: inst = 32'h10408000;
      12136: inst = 32'hc404ed6;
      12137: inst = 32'h8220000;
      12138: inst = 32'h10408000;
      12139: inst = 32'hc404ed7;
      12140: inst = 32'h8220000;
      12141: inst = 32'h10408000;
      12142: inst = 32'hc404ed8;
      12143: inst = 32'h8220000;
      12144: inst = 32'h10408000;
      12145: inst = 32'hc404ed9;
      12146: inst = 32'h8220000;
      12147: inst = 32'h10408000;
      12148: inst = 32'hc404eda;
      12149: inst = 32'h8220000;
      12150: inst = 32'h10408000;
      12151: inst = 32'hc404edb;
      12152: inst = 32'h8220000;
      12153: inst = 32'h10408000;
      12154: inst = 32'hc404edc;
      12155: inst = 32'h8220000;
      12156: inst = 32'h10408000;
      12157: inst = 32'hc404edd;
      12158: inst = 32'h8220000;
      12159: inst = 32'h10408000;
      12160: inst = 32'hc404ede;
      12161: inst = 32'h8220000;
      12162: inst = 32'h10408000;
      12163: inst = 32'hc404f30;
      12164: inst = 32'h8220000;
      12165: inst = 32'h10408000;
      12166: inst = 32'hc404f31;
      12167: inst = 32'h8220000;
      12168: inst = 32'h10408000;
      12169: inst = 32'hc404f32;
      12170: inst = 32'h8220000;
      12171: inst = 32'h10408000;
      12172: inst = 32'hc404f33;
      12173: inst = 32'h8220000;
      12174: inst = 32'h10408000;
      12175: inst = 32'hc404f34;
      12176: inst = 32'h8220000;
      12177: inst = 32'h10408000;
      12178: inst = 32'hc404f35;
      12179: inst = 32'h8220000;
      12180: inst = 32'h10408000;
      12181: inst = 32'hc404f36;
      12182: inst = 32'h8220000;
      12183: inst = 32'h10408000;
      12184: inst = 32'hc404f37;
      12185: inst = 32'h8220000;
      12186: inst = 32'h10408000;
      12187: inst = 32'hc404f38;
      12188: inst = 32'h8220000;
      12189: inst = 32'h10408000;
      12190: inst = 32'hc404f39;
      12191: inst = 32'h8220000;
      12192: inst = 32'h10408000;
      12193: inst = 32'hc404f3a;
      12194: inst = 32'h8220000;
      12195: inst = 32'h10408000;
      12196: inst = 32'hc404f3b;
      12197: inst = 32'h8220000;
      12198: inst = 32'h10408000;
      12199: inst = 32'hc404f3c;
      12200: inst = 32'h8220000;
      12201: inst = 32'h10408000;
      12202: inst = 32'hc404f3d;
      12203: inst = 32'h8220000;
      12204: inst = 32'h10408000;
      12205: inst = 32'hc404f3e;
      12206: inst = 32'h8220000;
      12207: inst = 32'h10408000;
      12208: inst = 32'hc404f90;
      12209: inst = 32'h8220000;
      12210: inst = 32'h10408000;
      12211: inst = 32'hc404f91;
      12212: inst = 32'h8220000;
      12213: inst = 32'h10408000;
      12214: inst = 32'hc404f92;
      12215: inst = 32'h8220000;
      12216: inst = 32'h10408000;
      12217: inst = 32'hc404f93;
      12218: inst = 32'h8220000;
      12219: inst = 32'h10408000;
      12220: inst = 32'hc404f94;
      12221: inst = 32'h8220000;
      12222: inst = 32'h10408000;
      12223: inst = 32'hc404f95;
      12224: inst = 32'h8220000;
      12225: inst = 32'h10408000;
      12226: inst = 32'hc404f96;
      12227: inst = 32'h8220000;
      12228: inst = 32'h10408000;
      12229: inst = 32'hc404f97;
      12230: inst = 32'h8220000;
      12231: inst = 32'h10408000;
      12232: inst = 32'hc404f98;
      12233: inst = 32'h8220000;
      12234: inst = 32'h10408000;
      12235: inst = 32'hc404f99;
      12236: inst = 32'h8220000;
      12237: inst = 32'h10408000;
      12238: inst = 32'hc404f9a;
      12239: inst = 32'h8220000;
      12240: inst = 32'h10408000;
      12241: inst = 32'hc404f9b;
      12242: inst = 32'h8220000;
      12243: inst = 32'h10408000;
      12244: inst = 32'hc404f9c;
      12245: inst = 32'h8220000;
      12246: inst = 32'h10408000;
      12247: inst = 32'hc404f9d;
      12248: inst = 32'h8220000;
      12249: inst = 32'h10408000;
      12250: inst = 32'hc404f9e;
      12251: inst = 32'h8220000;
      12252: inst = 32'h10408000;
      12253: inst = 32'hc404ff0;
      12254: inst = 32'h8220000;
      12255: inst = 32'h10408000;
      12256: inst = 32'hc404ff1;
      12257: inst = 32'h8220000;
      12258: inst = 32'h10408000;
      12259: inst = 32'hc404ff2;
      12260: inst = 32'h8220000;
      12261: inst = 32'h10408000;
      12262: inst = 32'hc404ff3;
      12263: inst = 32'h8220000;
      12264: inst = 32'h10408000;
      12265: inst = 32'hc404ff4;
      12266: inst = 32'h8220000;
      12267: inst = 32'h10408000;
      12268: inst = 32'hc404ff5;
      12269: inst = 32'h8220000;
      12270: inst = 32'h10408000;
      12271: inst = 32'hc404ff6;
      12272: inst = 32'h8220000;
      12273: inst = 32'h10408000;
      12274: inst = 32'hc404ff7;
      12275: inst = 32'h8220000;
      12276: inst = 32'h10408000;
      12277: inst = 32'hc404ff8;
      12278: inst = 32'h8220000;
      12279: inst = 32'h10408000;
      12280: inst = 32'hc404ff9;
      12281: inst = 32'h8220000;
      12282: inst = 32'h10408000;
      12283: inst = 32'hc404ffa;
      12284: inst = 32'h8220000;
      12285: inst = 32'h10408000;
      12286: inst = 32'hc404ffb;
      12287: inst = 32'h8220000;
      12288: inst = 32'h10408000;
      12289: inst = 32'hc404ffc;
      12290: inst = 32'h8220000;
      12291: inst = 32'h10408000;
      12292: inst = 32'hc404ffd;
      12293: inst = 32'h8220000;
      12294: inst = 32'h10408000;
      12295: inst = 32'hc404ffe;
      12296: inst = 32'h8220000;
      12297: inst = 32'h10408000;
      12298: inst = 32'hc405050;
      12299: inst = 32'h8220000;
      12300: inst = 32'h10408000;
      12301: inst = 32'hc405051;
      12302: inst = 32'h8220000;
      12303: inst = 32'h10408000;
      12304: inst = 32'hc405052;
      12305: inst = 32'h8220000;
      12306: inst = 32'h10408000;
      12307: inst = 32'hc405053;
      12308: inst = 32'h8220000;
      12309: inst = 32'h10408000;
      12310: inst = 32'hc405054;
      12311: inst = 32'h8220000;
      12312: inst = 32'h10408000;
      12313: inst = 32'hc405055;
      12314: inst = 32'h8220000;
      12315: inst = 32'h10408000;
      12316: inst = 32'hc405056;
      12317: inst = 32'h8220000;
      12318: inst = 32'h10408000;
      12319: inst = 32'hc405057;
      12320: inst = 32'h8220000;
      12321: inst = 32'h10408000;
      12322: inst = 32'hc405058;
      12323: inst = 32'h8220000;
      12324: inst = 32'h10408000;
      12325: inst = 32'hc405059;
      12326: inst = 32'h8220000;
      12327: inst = 32'h10408000;
      12328: inst = 32'hc40505a;
      12329: inst = 32'h8220000;
      12330: inst = 32'h10408000;
      12331: inst = 32'hc40505b;
      12332: inst = 32'h8220000;
      12333: inst = 32'h10408000;
      12334: inst = 32'hc40505c;
      12335: inst = 32'h8220000;
      12336: inst = 32'h10408000;
      12337: inst = 32'hc40505d;
      12338: inst = 32'h8220000;
      12339: inst = 32'h10408000;
      12340: inst = 32'hc40505e;
      12341: inst = 32'h8220000;
      12342: inst = 32'h10408000;
      12343: inst = 32'hc4050b0;
      12344: inst = 32'h8220000;
      12345: inst = 32'h10408000;
      12346: inst = 32'hc4050b1;
      12347: inst = 32'h8220000;
      12348: inst = 32'h10408000;
      12349: inst = 32'hc4050b2;
      12350: inst = 32'h8220000;
      12351: inst = 32'h10408000;
      12352: inst = 32'hc4050b3;
      12353: inst = 32'h8220000;
      12354: inst = 32'h10408000;
      12355: inst = 32'hc4050b4;
      12356: inst = 32'h8220000;
      12357: inst = 32'h10408000;
      12358: inst = 32'hc4050b5;
      12359: inst = 32'h8220000;
      12360: inst = 32'h10408000;
      12361: inst = 32'hc4050b6;
      12362: inst = 32'h8220000;
      12363: inst = 32'h10408000;
      12364: inst = 32'hc4050b7;
      12365: inst = 32'h8220000;
      12366: inst = 32'h10408000;
      12367: inst = 32'hc4050b8;
      12368: inst = 32'h8220000;
      12369: inst = 32'h10408000;
      12370: inst = 32'hc4050b9;
      12371: inst = 32'h8220000;
      12372: inst = 32'h10408000;
      12373: inst = 32'hc4050ba;
      12374: inst = 32'h8220000;
      12375: inst = 32'h10408000;
      12376: inst = 32'hc4050bb;
      12377: inst = 32'h8220000;
      12378: inst = 32'h10408000;
      12379: inst = 32'hc4050bc;
      12380: inst = 32'h8220000;
      12381: inst = 32'h10408000;
      12382: inst = 32'hc4050bd;
      12383: inst = 32'h8220000;
      12384: inst = 32'h10408000;
      12385: inst = 32'hc4050be;
      12386: inst = 32'h8220000;
      12387: inst = 32'h10408000;
      12388: inst = 32'hc405110;
      12389: inst = 32'h8220000;
      12390: inst = 32'h10408000;
      12391: inst = 32'hc405111;
      12392: inst = 32'h8220000;
      12393: inst = 32'h10408000;
      12394: inst = 32'hc405112;
      12395: inst = 32'h8220000;
      12396: inst = 32'h10408000;
      12397: inst = 32'hc405113;
      12398: inst = 32'h8220000;
      12399: inst = 32'h10408000;
      12400: inst = 32'hc405114;
      12401: inst = 32'h8220000;
      12402: inst = 32'h10408000;
      12403: inst = 32'hc405115;
      12404: inst = 32'h8220000;
      12405: inst = 32'h10408000;
      12406: inst = 32'hc405116;
      12407: inst = 32'h8220000;
      12408: inst = 32'h10408000;
      12409: inst = 32'hc405117;
      12410: inst = 32'h8220000;
      12411: inst = 32'h10408000;
      12412: inst = 32'hc405118;
      12413: inst = 32'h8220000;
      12414: inst = 32'h10408000;
      12415: inst = 32'hc405119;
      12416: inst = 32'h8220000;
      12417: inst = 32'h10408000;
      12418: inst = 32'hc40511a;
      12419: inst = 32'h8220000;
      12420: inst = 32'h10408000;
      12421: inst = 32'hc40511b;
      12422: inst = 32'h8220000;
      12423: inst = 32'h10408000;
      12424: inst = 32'hc40511c;
      12425: inst = 32'h8220000;
      12426: inst = 32'h10408000;
      12427: inst = 32'hc40511d;
      12428: inst = 32'h8220000;
      12429: inst = 32'h10408000;
      12430: inst = 32'hc40511e;
      12431: inst = 32'h8220000;
      12432: inst = 32'h10408000;
      12433: inst = 32'hc405170;
      12434: inst = 32'h8220000;
      12435: inst = 32'h10408000;
      12436: inst = 32'hc405171;
      12437: inst = 32'h8220000;
      12438: inst = 32'h10408000;
      12439: inst = 32'hc405172;
      12440: inst = 32'h8220000;
      12441: inst = 32'h10408000;
      12442: inst = 32'hc405173;
      12443: inst = 32'h8220000;
      12444: inst = 32'h10408000;
      12445: inst = 32'hc405174;
      12446: inst = 32'h8220000;
      12447: inst = 32'h10408000;
      12448: inst = 32'hc405175;
      12449: inst = 32'h8220000;
      12450: inst = 32'h10408000;
      12451: inst = 32'hc405176;
      12452: inst = 32'h8220000;
      12453: inst = 32'h10408000;
      12454: inst = 32'hc405177;
      12455: inst = 32'h8220000;
      12456: inst = 32'h10408000;
      12457: inst = 32'hc405178;
      12458: inst = 32'h8220000;
      12459: inst = 32'h10408000;
      12460: inst = 32'hc405179;
      12461: inst = 32'h8220000;
      12462: inst = 32'h10408000;
      12463: inst = 32'hc40517a;
      12464: inst = 32'h8220000;
      12465: inst = 32'h10408000;
      12466: inst = 32'hc40517b;
      12467: inst = 32'h8220000;
      12468: inst = 32'h10408000;
      12469: inst = 32'hc40517c;
      12470: inst = 32'h8220000;
      12471: inst = 32'h10408000;
      12472: inst = 32'hc40517d;
      12473: inst = 32'h8220000;
      12474: inst = 32'h10408000;
      12475: inst = 32'hc40517e;
      12476: inst = 32'h8220000;
      12477: inst = 32'h10408000;
      12478: inst = 32'hc4051d0;
      12479: inst = 32'h8220000;
      12480: inst = 32'h10408000;
      12481: inst = 32'hc4051d1;
      12482: inst = 32'h8220000;
      12483: inst = 32'h10408000;
      12484: inst = 32'hc4051d2;
      12485: inst = 32'h8220000;
      12486: inst = 32'h10408000;
      12487: inst = 32'hc4051d3;
      12488: inst = 32'h8220000;
      12489: inst = 32'h10408000;
      12490: inst = 32'hc4051d4;
      12491: inst = 32'h8220000;
      12492: inst = 32'h10408000;
      12493: inst = 32'hc4051d5;
      12494: inst = 32'h8220000;
      12495: inst = 32'h10408000;
      12496: inst = 32'hc4051d6;
      12497: inst = 32'h8220000;
      12498: inst = 32'h10408000;
      12499: inst = 32'hc4051d7;
      12500: inst = 32'h8220000;
      12501: inst = 32'h10408000;
      12502: inst = 32'hc4051d8;
      12503: inst = 32'h8220000;
      12504: inst = 32'h10408000;
      12505: inst = 32'hc4051d9;
      12506: inst = 32'h8220000;
      12507: inst = 32'h10408000;
      12508: inst = 32'hc4051da;
      12509: inst = 32'h8220000;
      12510: inst = 32'h10408000;
      12511: inst = 32'hc4051db;
      12512: inst = 32'h8220000;
      12513: inst = 32'h10408000;
      12514: inst = 32'hc4051dc;
      12515: inst = 32'h8220000;
      12516: inst = 32'h10408000;
      12517: inst = 32'hc4051dd;
      12518: inst = 32'h8220000;
      12519: inst = 32'h10408000;
      12520: inst = 32'hc4051de;
      12521: inst = 32'h8220000;
      12522: inst = 32'h10408000;
      12523: inst = 32'hc405230;
      12524: inst = 32'h8220000;
      12525: inst = 32'h10408000;
      12526: inst = 32'hc405231;
      12527: inst = 32'h8220000;
      12528: inst = 32'h10408000;
      12529: inst = 32'hc405232;
      12530: inst = 32'h8220000;
      12531: inst = 32'h10408000;
      12532: inst = 32'hc405233;
      12533: inst = 32'h8220000;
      12534: inst = 32'h10408000;
      12535: inst = 32'hc405234;
      12536: inst = 32'h8220000;
      12537: inst = 32'h10408000;
      12538: inst = 32'hc405235;
      12539: inst = 32'h8220000;
      12540: inst = 32'h10408000;
      12541: inst = 32'hc405236;
      12542: inst = 32'h8220000;
      12543: inst = 32'h10408000;
      12544: inst = 32'hc405237;
      12545: inst = 32'h8220000;
      12546: inst = 32'h10408000;
      12547: inst = 32'hc405238;
      12548: inst = 32'h8220000;
      12549: inst = 32'h10408000;
      12550: inst = 32'hc405239;
      12551: inst = 32'h8220000;
      12552: inst = 32'h10408000;
      12553: inst = 32'hc40523a;
      12554: inst = 32'h8220000;
      12555: inst = 32'h10408000;
      12556: inst = 32'hc40523b;
      12557: inst = 32'h8220000;
      12558: inst = 32'h10408000;
      12559: inst = 32'hc40523c;
      12560: inst = 32'h8220000;
      12561: inst = 32'h10408000;
      12562: inst = 32'hc40523d;
      12563: inst = 32'h8220000;
      12564: inst = 32'h10408000;
      12565: inst = 32'hc40523e;
      12566: inst = 32'h8220000;
      12567: inst = 32'h10408000;
      12568: inst = 32'hc405290;
      12569: inst = 32'h8220000;
      12570: inst = 32'h10408000;
      12571: inst = 32'hc405291;
      12572: inst = 32'h8220000;
      12573: inst = 32'h10408000;
      12574: inst = 32'hc405292;
      12575: inst = 32'h8220000;
      12576: inst = 32'h10408000;
      12577: inst = 32'hc405293;
      12578: inst = 32'h8220000;
      12579: inst = 32'h10408000;
      12580: inst = 32'hc405294;
      12581: inst = 32'h8220000;
      12582: inst = 32'h10408000;
      12583: inst = 32'hc405295;
      12584: inst = 32'h8220000;
      12585: inst = 32'h10408000;
      12586: inst = 32'hc405296;
      12587: inst = 32'h8220000;
      12588: inst = 32'h10408000;
      12589: inst = 32'hc405297;
      12590: inst = 32'h8220000;
      12591: inst = 32'h10408000;
      12592: inst = 32'hc405298;
      12593: inst = 32'h8220000;
      12594: inst = 32'h10408000;
      12595: inst = 32'hc405299;
      12596: inst = 32'h8220000;
      12597: inst = 32'h10408000;
      12598: inst = 32'hc40529a;
      12599: inst = 32'h8220000;
      12600: inst = 32'h10408000;
      12601: inst = 32'hc40529b;
      12602: inst = 32'h8220000;
      12603: inst = 32'h10408000;
      12604: inst = 32'hc40529c;
      12605: inst = 32'h8220000;
      12606: inst = 32'h10408000;
      12607: inst = 32'hc40529d;
      12608: inst = 32'h8220000;
      12609: inst = 32'h10408000;
      12610: inst = 32'hc40529e;
      12611: inst = 32'h8220000;
      12612: inst = 32'hc20ef7c;
      12613: inst = 32'h10408000;
      12614: inst = 32'hc404932;
      12615: inst = 32'h8220000;
      12616: inst = 32'h10408000;
      12617: inst = 32'hc404933;
      12618: inst = 32'h8220000;
      12619: inst = 32'h10408000;
      12620: inst = 32'hc404934;
      12621: inst = 32'h8220000;
      12622: inst = 32'h10408000;
      12623: inst = 32'hc404935;
      12624: inst = 32'h8220000;
      12625: inst = 32'h10408000;
      12626: inst = 32'hc404993;
      12627: inst = 32'h8220000;
      12628: inst = 32'h10408000;
      12629: inst = 32'hc404994;
      12630: inst = 32'h8220000;
      12631: inst = 32'h10408000;
      12632: inst = 32'hc404995;
      12633: inst = 32'h8220000;
      12634: inst = 32'h10408000;
      12635: inst = 32'hc4049f3;
      12636: inst = 32'h8220000;
      12637: inst = 32'h10408000;
      12638: inst = 32'hc4049f4;
      12639: inst = 32'h8220000;
      12640: inst = 32'h10408000;
      12641: inst = 32'hc4049f5;
      12642: inst = 32'h8220000;
      12643: inst = 32'h10408000;
      12644: inst = 32'hc404a53;
      12645: inst = 32'h8220000;
      12646: inst = 32'h10408000;
      12647: inst = 32'hc404a54;
      12648: inst = 32'h8220000;
      12649: inst = 32'h10408000;
      12650: inst = 32'hc404a55;
      12651: inst = 32'h8220000;
      12652: inst = 32'h10408000;
      12653: inst = 32'hc404ab2;
      12654: inst = 32'h8220000;
      12655: inst = 32'h10408000;
      12656: inst = 32'hc404ab3;
      12657: inst = 32'h8220000;
      12658: inst = 32'h10408000;
      12659: inst = 32'hc404ab5;
      12660: inst = 32'h8220000;
      12661: inst = 32'h10408000;
      12662: inst = 32'hc404b12;
      12663: inst = 32'h8220000;
      12664: inst = 32'h10408000;
      12665: inst = 32'hc404b13;
      12666: inst = 32'h8220000;
      12667: inst = 32'h10408000;
      12668: inst = 32'hc404b15;
      12669: inst = 32'h8220000;
      12670: inst = 32'h10408000;
      12671: inst = 32'hc404b72;
      12672: inst = 32'h8220000;
      12673: inst = 32'h10408000;
      12674: inst = 32'hc404b73;
      12675: inst = 32'h8220000;
      12676: inst = 32'h10408000;
      12677: inst = 32'hc404b74;
      12678: inst = 32'h8220000;
      12679: inst = 32'h10408000;
      12680: inst = 32'hc404b75;
      12681: inst = 32'h8220000;
      12682: inst = 32'hc20eed7;
      12683: inst = 32'h10408000;
      12684: inst = 32'hc404a08;
      12685: inst = 32'h8220000;
      12686: inst = 32'h10408000;
      12687: inst = 32'hc404a0e;
      12688: inst = 32'h8220000;
      12689: inst = 32'hc20e6fa;
      12690: inst = 32'h10408000;
      12691: inst = 32'hc404a09;
      12692: inst = 32'h8220000;
      12693: inst = 32'h10408000;
      12694: inst = 32'hc404a0d;
      12695: inst = 32'h8220000;
      12696: inst = 32'h10408000;
      12697: inst = 32'hc404be7;
      12698: inst = 32'h8220000;
      12699: inst = 32'hc20e6fb;
      12700: inst = 32'h10408000;
      12701: inst = 32'hc404a0a;
      12702: inst = 32'h8220000;
      12703: inst = 32'h10408000;
      12704: inst = 32'hc404a0c;
      12705: inst = 32'h8220000;
      12706: inst = 32'h10408000;
      12707: inst = 32'hc404ac7;
      12708: inst = 32'h8220000;
      12709: inst = 32'h10408000;
      12710: inst = 32'hc404acf;
      12711: inst = 32'h8220000;
      12712: inst = 32'h10408000;
      12713: inst = 32'hc404b87;
      12714: inst = 32'h8220000;
      12715: inst = 32'h10408000;
      12716: inst = 32'hc404b8f;
      12717: inst = 32'h8220000;
      12718: inst = 32'h10408000;
      12719: inst = 32'hc404c4d;
      12720: inst = 32'h8220000;
      12721: inst = 32'hc20defb;
      12722: inst = 32'h10408000;
      12723: inst = 32'hc404a0b;
      12724: inst = 32'h8220000;
      12725: inst = 32'h10408000;
      12726: inst = 32'hc404a68;
      12727: inst = 32'h8220000;
      12728: inst = 32'h10408000;
      12729: inst = 32'hc404a69;
      12730: inst = 32'h8220000;
      12731: inst = 32'h10408000;
      12732: inst = 32'hc404a6a;
      12733: inst = 32'h8220000;
      12734: inst = 32'h10408000;
      12735: inst = 32'hc404a6b;
      12736: inst = 32'h8220000;
      12737: inst = 32'h10408000;
      12738: inst = 32'hc404a6c;
      12739: inst = 32'h8220000;
      12740: inst = 32'h10408000;
      12741: inst = 32'hc404a6d;
      12742: inst = 32'h8220000;
      12743: inst = 32'h10408000;
      12744: inst = 32'hc404a6e;
      12745: inst = 32'h8220000;
      12746: inst = 32'h10408000;
      12747: inst = 32'hc404ac8;
      12748: inst = 32'h8220000;
      12749: inst = 32'h10408000;
      12750: inst = 32'hc404ac9;
      12751: inst = 32'h8220000;
      12752: inst = 32'h10408000;
      12753: inst = 32'hc404aca;
      12754: inst = 32'h8220000;
      12755: inst = 32'h10408000;
      12756: inst = 32'hc404acb;
      12757: inst = 32'h8220000;
      12758: inst = 32'h10408000;
      12759: inst = 32'hc404acc;
      12760: inst = 32'h8220000;
      12761: inst = 32'h10408000;
      12762: inst = 32'hc404acd;
      12763: inst = 32'h8220000;
      12764: inst = 32'h10408000;
      12765: inst = 32'hc404ace;
      12766: inst = 32'h8220000;
      12767: inst = 32'h10408000;
      12768: inst = 32'hc404b27;
      12769: inst = 32'h8220000;
      12770: inst = 32'h10408000;
      12771: inst = 32'hc404b2a;
      12772: inst = 32'h8220000;
      12773: inst = 32'h10408000;
      12774: inst = 32'hc404b2d;
      12775: inst = 32'h8220000;
      12776: inst = 32'h10408000;
      12777: inst = 32'hc404b2e;
      12778: inst = 32'h8220000;
      12779: inst = 32'h10408000;
      12780: inst = 32'hc404b2f;
      12781: inst = 32'h8220000;
      12782: inst = 32'h10408000;
      12783: inst = 32'hc404b8a;
      12784: inst = 32'h8220000;
      12785: inst = 32'h10408000;
      12786: inst = 32'hc404b8d;
      12787: inst = 32'h8220000;
      12788: inst = 32'h10408000;
      12789: inst = 32'hc404b8e;
      12790: inst = 32'h8220000;
      12791: inst = 32'h10408000;
      12792: inst = 32'hc404be8;
      12793: inst = 32'h8220000;
      12794: inst = 32'h10408000;
      12795: inst = 32'hc404be9;
      12796: inst = 32'h8220000;
      12797: inst = 32'h10408000;
      12798: inst = 32'hc404bea;
      12799: inst = 32'h8220000;
      12800: inst = 32'h10408000;
      12801: inst = 32'hc404beb;
      12802: inst = 32'h8220000;
      12803: inst = 32'h10408000;
      12804: inst = 32'hc404bec;
      12805: inst = 32'h8220000;
      12806: inst = 32'h10408000;
      12807: inst = 32'hc404bed;
      12808: inst = 32'h8220000;
      12809: inst = 32'h10408000;
      12810: inst = 32'hc404bee;
      12811: inst = 32'h8220000;
      12812: inst = 32'h10408000;
      12813: inst = 32'hc404c49;
      12814: inst = 32'h8220000;
      12815: inst = 32'h10408000;
      12816: inst = 32'hc404c4b;
      12817: inst = 32'h8220000;
      12818: inst = 32'h10408000;
      12819: inst = 32'hc404ca9;
      12820: inst = 32'h8220000;
      12821: inst = 32'h10408000;
      12822: inst = 32'hc404cab;
      12823: inst = 32'h8220000;
      12824: inst = 32'hc20eed8;
      12825: inst = 32'h10408000;
      12826: inst = 32'hc404a67;
      12827: inst = 32'h8220000;
      12828: inst = 32'h10408000;
      12829: inst = 32'hc404a6f;
      12830: inst = 32'h8220000;
      12831: inst = 32'hc204a69;
      12832: inst = 32'h10408000;
      12833: inst = 32'hc404b28;
      12834: inst = 32'h8220000;
      12835: inst = 32'h10408000;
      12836: inst = 32'hc404b29;
      12837: inst = 32'h8220000;
      12838: inst = 32'h10408000;
      12839: inst = 32'hc404b2b;
      12840: inst = 32'h8220000;
      12841: inst = 32'h10408000;
      12842: inst = 32'hc404b2c;
      12843: inst = 32'h8220000;
      12844: inst = 32'h10408000;
      12845: inst = 32'hc404b88;
      12846: inst = 32'h8220000;
      12847: inst = 32'h10408000;
      12848: inst = 32'hc404b89;
      12849: inst = 32'h8220000;
      12850: inst = 32'h10408000;
      12851: inst = 32'hc404b8b;
      12852: inst = 32'h8220000;
      12853: inst = 32'h10408000;
      12854: inst = 32'hc404b8c;
      12855: inst = 32'h8220000;
      12856: inst = 32'h10408000;
      12857: inst = 32'hc404c48;
      12858: inst = 32'h8220000;
      12859: inst = 32'h10408000;
      12860: inst = 32'hc404c4a;
      12861: inst = 32'h8220000;
      12862: inst = 32'h10408000;
      12863: inst = 32'hc404c4c;
      12864: inst = 32'h8220000;
      12865: inst = 32'h10408000;
      12866: inst = 32'hc404ca8;
      12867: inst = 32'h8220000;
      12868: inst = 32'h10408000;
      12869: inst = 32'hc404caa;
      12870: inst = 32'h8220000;
      12871: inst = 32'h10408000;
      12872: inst = 32'hc404cac;
      12873: inst = 32'h8220000;
      12874: inst = 32'h10408000;
      12875: inst = 32'hc405085;
      12876: inst = 32'h8220000;
      12877: inst = 32'h10408000;
      12878: inst = 32'hc40509a;
      12879: inst = 32'h8220000;
      12880: inst = 32'h10408000;
      12881: inst = 32'hc4050e4;
      12882: inst = 32'h8220000;
      12883: inst = 32'h10408000;
      12884: inst = 32'hc4050e5;
      12885: inst = 32'h8220000;
      12886: inst = 32'h10408000;
      12887: inst = 32'hc4050fa;
      12888: inst = 32'h8220000;
      12889: inst = 32'h10408000;
      12890: inst = 32'hc4050fb;
      12891: inst = 32'h8220000;
      12892: inst = 32'h10408000;
      12893: inst = 32'hc405143;
      12894: inst = 32'h8220000;
      12895: inst = 32'h10408000;
      12896: inst = 32'hc405144;
      12897: inst = 32'h8220000;
      12898: inst = 32'h10408000;
      12899: inst = 32'hc405145;
      12900: inst = 32'h8220000;
      12901: inst = 32'h10408000;
      12902: inst = 32'hc40515a;
      12903: inst = 32'h8220000;
      12904: inst = 32'h10408000;
      12905: inst = 32'hc40515b;
      12906: inst = 32'h8220000;
      12907: inst = 32'h10408000;
      12908: inst = 32'hc40515c;
      12909: inst = 32'h8220000;
      12910: inst = 32'h10408000;
      12911: inst = 32'hc4051a2;
      12912: inst = 32'h8220000;
      12913: inst = 32'h10408000;
      12914: inst = 32'hc4051a3;
      12915: inst = 32'h8220000;
      12916: inst = 32'h10408000;
      12917: inst = 32'hc4051a4;
      12918: inst = 32'h8220000;
      12919: inst = 32'h10408000;
      12920: inst = 32'hc4051a5;
      12921: inst = 32'h8220000;
      12922: inst = 32'h10408000;
      12923: inst = 32'hc4051ba;
      12924: inst = 32'h8220000;
      12925: inst = 32'h10408000;
      12926: inst = 32'hc4051bb;
      12927: inst = 32'h8220000;
      12928: inst = 32'h10408000;
      12929: inst = 32'hc4051bc;
      12930: inst = 32'h8220000;
      12931: inst = 32'h10408000;
      12932: inst = 32'hc4051bd;
      12933: inst = 32'h8220000;
      12934: inst = 32'h10408000;
      12935: inst = 32'hc405202;
      12936: inst = 32'h8220000;
      12937: inst = 32'h10408000;
      12938: inst = 32'hc405203;
      12939: inst = 32'h8220000;
      12940: inst = 32'h10408000;
      12941: inst = 32'hc405204;
      12942: inst = 32'h8220000;
      12943: inst = 32'h10408000;
      12944: inst = 32'hc405205;
      12945: inst = 32'h8220000;
      12946: inst = 32'h10408000;
      12947: inst = 32'hc40521a;
      12948: inst = 32'h8220000;
      12949: inst = 32'h10408000;
      12950: inst = 32'hc40521b;
      12951: inst = 32'h8220000;
      12952: inst = 32'h10408000;
      12953: inst = 32'hc40521c;
      12954: inst = 32'h8220000;
      12955: inst = 32'h10408000;
      12956: inst = 32'hc40521d;
      12957: inst = 32'h8220000;
      12958: inst = 32'h10408000;
      12959: inst = 32'hc405262;
      12960: inst = 32'h8220000;
      12961: inst = 32'h10408000;
      12962: inst = 32'hc405263;
      12963: inst = 32'h8220000;
      12964: inst = 32'h10408000;
      12965: inst = 32'hc405264;
      12966: inst = 32'h8220000;
      12967: inst = 32'h10408000;
      12968: inst = 32'hc405265;
      12969: inst = 32'h8220000;
      12970: inst = 32'h10408000;
      12971: inst = 32'hc40527a;
      12972: inst = 32'h8220000;
      12973: inst = 32'h10408000;
      12974: inst = 32'hc40527b;
      12975: inst = 32'h8220000;
      12976: inst = 32'h10408000;
      12977: inst = 32'hc40527c;
      12978: inst = 32'h8220000;
      12979: inst = 32'h10408000;
      12980: inst = 32'hc40527d;
      12981: inst = 32'h8220000;
      12982: inst = 32'h10408000;
      12983: inst = 32'hc4052c2;
      12984: inst = 32'h8220000;
      12985: inst = 32'h10408000;
      12986: inst = 32'hc4052c3;
      12987: inst = 32'h8220000;
      12988: inst = 32'h10408000;
      12989: inst = 32'hc4052c4;
      12990: inst = 32'h8220000;
      12991: inst = 32'h10408000;
      12992: inst = 32'hc4052db;
      12993: inst = 32'h8220000;
      12994: inst = 32'h10408000;
      12995: inst = 32'hc4052dc;
      12996: inst = 32'h8220000;
      12997: inst = 32'h10408000;
      12998: inst = 32'hc4052dd;
      12999: inst = 32'h8220000;
      13000: inst = 32'h10408000;
      13001: inst = 32'hc405322;
      13002: inst = 32'h8220000;
      13003: inst = 32'h10408000;
      13004: inst = 32'hc405323;
      13005: inst = 32'h8220000;
      13006: inst = 32'h10408000;
      13007: inst = 32'hc405324;
      13008: inst = 32'h8220000;
      13009: inst = 32'h10408000;
      13010: inst = 32'hc40533b;
      13011: inst = 32'h8220000;
      13012: inst = 32'h10408000;
      13013: inst = 32'hc40533c;
      13014: inst = 32'h8220000;
      13015: inst = 32'h10408000;
      13016: inst = 32'hc40533d;
      13017: inst = 32'h8220000;
      13018: inst = 32'h10408000;
      13019: inst = 32'hc40537f;
      13020: inst = 32'h8220000;
      13021: inst = 32'h10408000;
      13022: inst = 32'hc405382;
      13023: inst = 32'h8220000;
      13024: inst = 32'h10408000;
      13025: inst = 32'hc405383;
      13026: inst = 32'h8220000;
      13027: inst = 32'h10408000;
      13028: inst = 32'hc405384;
      13029: inst = 32'h8220000;
      13030: inst = 32'h10408000;
      13031: inst = 32'hc40539b;
      13032: inst = 32'h8220000;
      13033: inst = 32'h10408000;
      13034: inst = 32'hc40539c;
      13035: inst = 32'h8220000;
      13036: inst = 32'h10408000;
      13037: inst = 32'hc40539d;
      13038: inst = 32'h8220000;
      13039: inst = 32'h10408000;
      13040: inst = 32'hc4053a0;
      13041: inst = 32'h8220000;
      13042: inst = 32'h10408000;
      13043: inst = 32'hc4053de;
      13044: inst = 32'h8220000;
      13045: inst = 32'h10408000;
      13046: inst = 32'hc4053df;
      13047: inst = 32'h8220000;
      13048: inst = 32'h10408000;
      13049: inst = 32'hc4053e2;
      13050: inst = 32'h8220000;
      13051: inst = 32'h10408000;
      13052: inst = 32'hc4053e3;
      13053: inst = 32'h8220000;
      13054: inst = 32'h10408000;
      13055: inst = 32'hc4053fc;
      13056: inst = 32'h8220000;
      13057: inst = 32'h10408000;
      13058: inst = 32'hc4053fd;
      13059: inst = 32'h8220000;
      13060: inst = 32'h10408000;
      13061: inst = 32'hc405400;
      13062: inst = 32'h8220000;
      13063: inst = 32'h10408000;
      13064: inst = 32'hc405401;
      13065: inst = 32'h8220000;
      13066: inst = 32'h10408000;
      13067: inst = 32'hc40543d;
      13068: inst = 32'h8220000;
      13069: inst = 32'h10408000;
      13070: inst = 32'hc40543e;
      13071: inst = 32'h8220000;
      13072: inst = 32'h10408000;
      13073: inst = 32'hc40543f;
      13074: inst = 32'h8220000;
      13075: inst = 32'h10408000;
      13076: inst = 32'hc405442;
      13077: inst = 32'h8220000;
      13078: inst = 32'h10408000;
      13079: inst = 32'hc405443;
      13080: inst = 32'h8220000;
      13081: inst = 32'h10408000;
      13082: inst = 32'hc40545c;
      13083: inst = 32'h8220000;
      13084: inst = 32'h10408000;
      13085: inst = 32'hc40545d;
      13086: inst = 32'h8220000;
      13087: inst = 32'h10408000;
      13088: inst = 32'hc405460;
      13089: inst = 32'h8220000;
      13090: inst = 32'h10408000;
      13091: inst = 32'hc405461;
      13092: inst = 32'h8220000;
      13093: inst = 32'h10408000;
      13094: inst = 32'hc405462;
      13095: inst = 32'h8220000;
      13096: inst = 32'h10408000;
      13097: inst = 32'hc40549d;
      13098: inst = 32'h8220000;
      13099: inst = 32'h10408000;
      13100: inst = 32'hc40549e;
      13101: inst = 32'h8220000;
      13102: inst = 32'h10408000;
      13103: inst = 32'hc4054a0;
      13104: inst = 32'h8220000;
      13105: inst = 32'h10408000;
      13106: inst = 32'hc4054a1;
      13107: inst = 32'h8220000;
      13108: inst = 32'h10408000;
      13109: inst = 32'hc4054a2;
      13110: inst = 32'h8220000;
      13111: inst = 32'h10408000;
      13112: inst = 32'hc4054a3;
      13113: inst = 32'h8220000;
      13114: inst = 32'h10408000;
      13115: inst = 32'hc4054bc;
      13116: inst = 32'h8220000;
      13117: inst = 32'h10408000;
      13118: inst = 32'hc4054bd;
      13119: inst = 32'h8220000;
      13120: inst = 32'h10408000;
      13121: inst = 32'hc4054be;
      13122: inst = 32'h8220000;
      13123: inst = 32'h10408000;
      13124: inst = 32'hc4054bf;
      13125: inst = 32'h8220000;
      13126: inst = 32'h10408000;
      13127: inst = 32'hc4054c1;
      13128: inst = 32'h8220000;
      13129: inst = 32'h10408000;
      13130: inst = 32'hc4054c2;
      13131: inst = 32'h8220000;
      13132: inst = 32'h10408000;
      13133: inst = 32'hc4054fc;
      13134: inst = 32'h8220000;
      13135: inst = 32'h10408000;
      13136: inst = 32'hc4054fd;
      13137: inst = 32'h8220000;
      13138: inst = 32'h10408000;
      13139: inst = 32'hc4054fe;
      13140: inst = 32'h8220000;
      13141: inst = 32'h10408000;
      13142: inst = 32'hc405502;
      13143: inst = 32'h8220000;
      13144: inst = 32'h10408000;
      13145: inst = 32'hc40551d;
      13146: inst = 32'h8220000;
      13147: inst = 32'h10408000;
      13148: inst = 32'hc405521;
      13149: inst = 32'h8220000;
      13150: inst = 32'h10408000;
      13151: inst = 32'hc405522;
      13152: inst = 32'h8220000;
      13153: inst = 32'h10408000;
      13154: inst = 32'hc405523;
      13155: inst = 32'h8220000;
      13156: inst = 32'h10408000;
      13157: inst = 32'hc40555b;
      13158: inst = 32'h8220000;
      13159: inst = 32'h10408000;
      13160: inst = 32'hc40555c;
      13161: inst = 32'h8220000;
      13162: inst = 32'h10408000;
      13163: inst = 32'hc40555d;
      13164: inst = 32'h8220000;
      13165: inst = 32'h10408000;
      13166: inst = 32'hc405562;
      13167: inst = 32'h8220000;
      13168: inst = 32'h10408000;
      13169: inst = 32'hc40557d;
      13170: inst = 32'h8220000;
      13171: inst = 32'h10408000;
      13172: inst = 32'hc405582;
      13173: inst = 32'h8220000;
      13174: inst = 32'h10408000;
      13175: inst = 32'hc405583;
      13176: inst = 32'h8220000;
      13177: inst = 32'h10408000;
      13178: inst = 32'hc405584;
      13179: inst = 32'h8220000;
      13180: inst = 32'h10408000;
      13181: inst = 32'hc4055ba;
      13182: inst = 32'h8220000;
      13183: inst = 32'h10408000;
      13184: inst = 32'hc4055bb;
      13185: inst = 32'h8220000;
      13186: inst = 32'h10408000;
      13187: inst = 32'hc4055bc;
      13188: inst = 32'h8220000;
      13189: inst = 32'h10408000;
      13190: inst = 32'hc4055bd;
      13191: inst = 32'h8220000;
      13192: inst = 32'h10408000;
      13193: inst = 32'hc4055c2;
      13194: inst = 32'h8220000;
      13195: inst = 32'h10408000;
      13196: inst = 32'hc4055dd;
      13197: inst = 32'h8220000;
      13198: inst = 32'h10408000;
      13199: inst = 32'hc4055e2;
      13200: inst = 32'h8220000;
      13201: inst = 32'h10408000;
      13202: inst = 32'hc4055e3;
      13203: inst = 32'h8220000;
      13204: inst = 32'h10408000;
      13205: inst = 32'hc4055e4;
      13206: inst = 32'h8220000;
      13207: inst = 32'h10408000;
      13208: inst = 32'hc4055e5;
      13209: inst = 32'h8220000;
      13210: inst = 32'h10408000;
      13211: inst = 32'hc40561a;
      13212: inst = 32'h8220000;
      13213: inst = 32'h10408000;
      13214: inst = 32'hc40561b;
      13215: inst = 32'h8220000;
      13216: inst = 32'h10408000;
      13217: inst = 32'hc40561c;
      13218: inst = 32'h8220000;
      13219: inst = 32'h10408000;
      13220: inst = 32'hc40561d;
      13221: inst = 32'h8220000;
      13222: inst = 32'h10408000;
      13223: inst = 32'hc405642;
      13224: inst = 32'h8220000;
      13225: inst = 32'h10408000;
      13226: inst = 32'hc405643;
      13227: inst = 32'h8220000;
      13228: inst = 32'h10408000;
      13229: inst = 32'hc405644;
      13230: inst = 32'h8220000;
      13231: inst = 32'h10408000;
      13232: inst = 32'hc405645;
      13233: inst = 32'h8220000;
      13234: inst = 32'h10408000;
      13235: inst = 32'hc405679;
      13236: inst = 32'h8220000;
      13237: inst = 32'h10408000;
      13238: inst = 32'hc40567a;
      13239: inst = 32'h8220000;
      13240: inst = 32'h10408000;
      13241: inst = 32'hc40567b;
      13242: inst = 32'h8220000;
      13243: inst = 32'h10408000;
      13244: inst = 32'hc40567c;
      13245: inst = 32'h8220000;
      13246: inst = 32'h10408000;
      13247: inst = 32'hc4056a3;
      13248: inst = 32'h8220000;
      13249: inst = 32'h10408000;
      13250: inst = 32'hc4056a4;
      13251: inst = 32'h8220000;
      13252: inst = 32'h10408000;
      13253: inst = 32'hc4056a5;
      13254: inst = 32'h8220000;
      13255: inst = 32'h10408000;
      13256: inst = 32'hc4056a6;
      13257: inst = 32'h8220000;
      13258: inst = 32'hc20e6d9;
      13259: inst = 32'h10408000;
      13260: inst = 32'hc404bef;
      13261: inst = 32'h8220000;
      13262: inst = 32'h10408000;
      13263: inst = 32'hc404c4e;
      13264: inst = 32'h8220000;
      13265: inst = 32'hc20eeb7;
      13266: inst = 32'h10408000;
      13267: inst = 32'hc404c47;
      13268: inst = 32'h8220000;
      13269: inst = 32'hc20d615;
      13270: inst = 32'h10408000;
      13271: inst = 32'hc404ca2;
      13272: inst = 32'h8220000;
      13273: inst = 32'h10408000;
      13274: inst = 32'hc404d00;
      13275: inst = 32'h8220000;
      13276: inst = 32'hc209c91;
      13277: inst = 32'h10408000;
      13278: inst = 32'hc404ca3;
      13279: inst = 32'h8220000;
      13280: inst = 32'h10408000;
      13281: inst = 32'hc404d01;
      13282: inst = 32'h8220000;
      13283: inst = 32'hc207bf0;
      13284: inst = 32'h10408000;
      13285: inst = 32'hc404ca4;
      13286: inst = 32'h8220000;
      13287: inst = 32'h10408000;
      13288: inst = 32'hc404ca5;
      13289: inst = 32'h8220000;
      13290: inst = 32'h10408000;
      13291: inst = 32'hc404ca6;
      13292: inst = 32'h8220000;
      13293: inst = 32'h10408000;
      13294: inst = 32'hc404ca7;
      13295: inst = 32'h8220000;
      13296: inst = 32'h10408000;
      13297: inst = 32'hc404d02;
      13298: inst = 32'h8220000;
      13299: inst = 32'h10408000;
      13300: inst = 32'hc404d03;
      13301: inst = 32'h8220000;
      13302: inst = 32'h10408000;
      13303: inst = 32'hc404d04;
      13304: inst = 32'h8220000;
      13305: inst = 32'h10408000;
      13306: inst = 32'hc404d05;
      13307: inst = 32'h8220000;
      13308: inst = 32'h10408000;
      13309: inst = 32'hc404d06;
      13310: inst = 32'h8220000;
      13311: inst = 32'h10408000;
      13312: inst = 32'hc404d07;
      13313: inst = 32'h8220000;
      13314: inst = 32'h10408000;
      13315: inst = 32'hc404d08;
      13316: inst = 32'h8220000;
      13317: inst = 32'h10408000;
      13318: inst = 32'hc404d09;
      13319: inst = 32'h8220000;
      13320: inst = 32'h10408000;
      13321: inst = 32'hc404d0a;
      13322: inst = 32'h8220000;
      13323: inst = 32'h10408000;
      13324: inst = 32'hc404d0b;
      13325: inst = 32'h8220000;
      13326: inst = 32'h10408000;
      13327: inst = 32'hc404d0c;
      13328: inst = 32'h8220000;
      13329: inst = 32'h10408000;
      13330: inst = 32'hc404d0d;
      13331: inst = 32'h8220000;
      13332: inst = 32'h10408000;
      13333: inst = 32'hc404d0e;
      13334: inst = 32'h8220000;
      13335: inst = 32'h10408000;
      13336: inst = 32'hc404d0f;
      13337: inst = 32'h8220000;
      13338: inst = 32'h10408000;
      13339: inst = 32'hc404d10;
      13340: inst = 32'h8220000;
      13341: inst = 32'h10408000;
      13342: inst = 32'hc404d11;
      13343: inst = 32'h8220000;
      13344: inst = 32'h10408000;
      13345: inst = 32'hc404d12;
      13346: inst = 32'h8220000;
      13347: inst = 32'h10408000;
      13348: inst = 32'hc404d13;
      13349: inst = 32'h8220000;
      13350: inst = 32'h10408000;
      13351: inst = 32'hc404d14;
      13352: inst = 32'h8220000;
      13353: inst = 32'h10408000;
      13354: inst = 32'hc4055c3;
      13355: inst = 32'h8220000;
      13356: inst = 32'h10408000;
      13357: inst = 32'hc4055dc;
      13358: inst = 32'h8220000;
      13359: inst = 32'hc20ad55;
      13360: inst = 32'h10408000;
      13361: inst = 32'hc404cad;
      13362: inst = 32'h8220000;
      13363: inst = 32'hc208410;
      13364: inst = 32'h10408000;
      13365: inst = 32'hc404cae;
      13366: inst = 32'h8220000;
      13367: inst = 32'h10408000;
      13368: inst = 32'hc404caf;
      13369: inst = 32'h8220000;
      13370: inst = 32'h10408000;
      13371: inst = 32'hc404cb0;
      13372: inst = 32'h8220000;
      13373: inst = 32'h10408000;
      13374: inst = 32'hc404cb1;
      13375: inst = 32'h8220000;
      13376: inst = 32'h10408000;
      13377: inst = 32'hc404cb2;
      13378: inst = 32'h8220000;
      13379: inst = 32'h10408000;
      13380: inst = 32'hc404cb3;
      13381: inst = 32'h8220000;
      13382: inst = 32'h10408000;
      13383: inst = 32'hc404cb4;
      13384: inst = 32'h8220000;
      13385: inst = 32'h10408000;
      13386: inst = 32'hc404cb5;
      13387: inst = 32'h8220000;
      13388: inst = 32'h10408000;
      13389: inst = 32'hc40537d;
      13390: inst = 32'h8220000;
      13391: inst = 32'h10408000;
      13392: inst = 32'hc405385;
      13393: inst = 32'h8220000;
      13394: inst = 32'h10408000;
      13395: inst = 32'hc40539a;
      13396: inst = 32'h8220000;
      13397: inst = 32'h10408000;
      13398: inst = 32'hc4053a2;
      13399: inst = 32'h8220000;
      13400: inst = 32'h10408000;
      13401: inst = 32'hc4054a4;
      13402: inst = 32'h8220000;
      13403: inst = 32'h10408000;
      13404: inst = 32'hc4054bb;
      13405: inst = 32'h8220000;
      13406: inst = 32'h10408000;
      13407: inst = 32'hc405741;
      13408: inst = 32'h8220000;
      13409: inst = 32'h10408000;
      13410: inst = 32'hc40575e;
      13411: inst = 32'h8220000;
      13412: inst = 32'hc209470;
      13413: inst = 32'h10408000;
      13414: inst = 32'hc404cb6;
      13415: inst = 32'h8220000;
      13416: inst = 32'h10408000;
      13417: inst = 32'hc404d15;
      13418: inst = 32'h8220000;
      13419: inst = 32'hc20a534;
      13420: inst = 32'h10408000;
      13421: inst = 32'hc404cfb;
      13422: inst = 32'h8220000;
      13423: inst = 32'hc208c51;
      13424: inst = 32'h10408000;
      13425: inst = 32'hc404cfc;
      13426: inst = 32'h8220000;
      13427: inst = 32'h10408000;
      13428: inst = 32'hc404cfd;
      13429: inst = 32'h8220000;
      13430: inst = 32'h10408000;
      13431: inst = 32'hc4053da;
      13432: inst = 32'h8220000;
      13433: inst = 32'h10408000;
      13434: inst = 32'hc4053dc;
      13435: inst = 32'h8220000;
      13436: inst = 32'h10408000;
      13437: inst = 32'hc405403;
      13438: inst = 32'h8220000;
      13439: inst = 32'h10408000;
      13440: inst = 32'hc405405;
      13441: inst = 32'h8220000;
      13442: inst = 32'h10408000;
      13443: inst = 32'hc4054fa;
      13444: inst = 32'h8220000;
      13445: inst = 32'h10408000;
      13446: inst = 32'hc405525;
      13447: inst = 32'h8220000;
      13448: inst = 32'h10408000;
      13449: inst = 32'hc405557;
      13450: inst = 32'h8220000;
      13451: inst = 32'h10408000;
      13452: inst = 32'hc40555f;
      13453: inst = 32'h8220000;
      13454: inst = 32'h10408000;
      13455: inst = 32'hc405580;
      13456: inst = 32'h8220000;
      13457: inst = 32'h10408000;
      13458: inst = 32'hc405588;
      13459: inst = 32'h8220000;
      13460: inst = 32'h10408000;
      13461: inst = 32'hc405618;
      13462: inst = 32'h8220000;
      13463: inst = 32'h10408000;
      13464: inst = 32'hc405627;
      13465: inst = 32'h8220000;
      13466: inst = 32'h10408000;
      13467: inst = 32'hc405638;
      13468: inst = 32'h8220000;
      13469: inst = 32'h10408000;
      13470: inst = 32'hc405647;
      13471: inst = 32'h8220000;
      13472: inst = 32'h10408000;
      13473: inst = 32'hc40570b;
      13474: inst = 32'h8220000;
      13475: inst = 32'hc206b6d;
      13476: inst = 32'h10408000;
      13477: inst = 32'hc404d16;
      13478: inst = 32'h8220000;
      13479: inst = 32'h10408000;
      13480: inst = 32'hc404d75;
      13481: inst = 32'h8220000;
      13482: inst = 32'h10408000;
      13483: inst = 32'hc404d76;
      13484: inst = 32'h8220000;
      13485: inst = 32'h10408000;
      13486: inst = 32'hc404dd5;
      13487: inst = 32'h8220000;
      13488: inst = 32'h10408000;
      13489: inst = 32'hc404dd6;
      13490: inst = 32'h8220000;
      13491: inst = 32'h10408000;
      13492: inst = 32'hc404e35;
      13493: inst = 32'h8220000;
      13494: inst = 32'h10408000;
      13495: inst = 32'hc404e36;
      13496: inst = 32'h8220000;
      13497: inst = 32'h10408000;
      13498: inst = 32'hc404e95;
      13499: inst = 32'h8220000;
      13500: inst = 32'h10408000;
      13501: inst = 32'hc404e96;
      13502: inst = 32'h8220000;
      13503: inst = 32'h10408000;
      13504: inst = 32'hc404ef5;
      13505: inst = 32'h8220000;
      13506: inst = 32'h10408000;
      13507: inst = 32'hc404ef6;
      13508: inst = 32'h8220000;
      13509: inst = 32'h10408000;
      13510: inst = 32'hc404f55;
      13511: inst = 32'h8220000;
      13512: inst = 32'h10408000;
      13513: inst = 32'hc404f56;
      13514: inst = 32'h8220000;
      13515: inst = 32'h10408000;
      13516: inst = 32'hc404fb5;
      13517: inst = 32'h8220000;
      13518: inst = 32'h10408000;
      13519: inst = 32'hc404fb6;
      13520: inst = 32'h8220000;
      13521: inst = 32'h10408000;
      13522: inst = 32'hc405015;
      13523: inst = 32'h8220000;
      13524: inst = 32'h10408000;
      13525: inst = 32'hc405016;
      13526: inst = 32'h8220000;
      13527: inst = 32'h10408000;
      13528: inst = 32'hc405075;
      13529: inst = 32'h8220000;
      13530: inst = 32'h10408000;
      13531: inst = 32'hc405076;
      13532: inst = 32'h8220000;
      13533: inst = 32'h10408000;
      13534: inst = 32'hc4050d5;
      13535: inst = 32'h8220000;
      13536: inst = 32'h10408000;
      13537: inst = 32'hc4050d6;
      13538: inst = 32'h8220000;
      13539: inst = 32'h10408000;
      13540: inst = 32'hc405135;
      13541: inst = 32'h8220000;
      13542: inst = 32'h10408000;
      13543: inst = 32'hc405136;
      13544: inst = 32'h8220000;
      13545: inst = 32'h10408000;
      13546: inst = 32'hc405195;
      13547: inst = 32'h8220000;
      13548: inst = 32'h10408000;
      13549: inst = 32'hc405196;
      13550: inst = 32'h8220000;
      13551: inst = 32'h10408000;
      13552: inst = 32'hc4051f5;
      13553: inst = 32'h8220000;
      13554: inst = 32'h10408000;
      13555: inst = 32'hc4051f6;
      13556: inst = 32'h8220000;
      13557: inst = 32'h10408000;
      13558: inst = 32'hc405255;
      13559: inst = 32'h8220000;
      13560: inst = 32'h10408000;
      13561: inst = 32'hc405256;
      13562: inst = 32'h8220000;
      13563: inst = 32'h10408000;
      13564: inst = 32'hc4052b5;
      13565: inst = 32'h8220000;
      13566: inst = 32'h10408000;
      13567: inst = 32'hc4052b6;
      13568: inst = 32'h8220000;
      13569: inst = 32'h10408000;
      13570: inst = 32'hc405325;
      13571: inst = 32'h8220000;
      13572: inst = 32'h10408000;
      13573: inst = 32'hc40533a;
      13574: inst = 32'h8220000;
      13575: inst = 32'hc20c638;
      13576: inst = 32'h10408000;
      13577: inst = 32'hc404d5b;
      13578: inst = 32'h8220000;
      13579: inst = 32'hc208c71;
      13580: inst = 32'h10408000;
      13581: inst = 32'hc404d60;
      13582: inst = 32'h8220000;
      13583: inst = 32'h10408000;
      13584: inst = 32'hc404d61;
      13585: inst = 32'h8220000;
      13586: inst = 32'h10408000;
      13587: inst = 32'hc404d62;
      13588: inst = 32'h8220000;
      13589: inst = 32'h10408000;
      13590: inst = 32'hc404d63;
      13591: inst = 32'h8220000;
      13592: inst = 32'h10408000;
      13593: inst = 32'hc404d64;
      13594: inst = 32'h8220000;
      13595: inst = 32'h10408000;
      13596: inst = 32'hc404d65;
      13597: inst = 32'h8220000;
      13598: inst = 32'h10408000;
      13599: inst = 32'hc404d66;
      13600: inst = 32'h8220000;
      13601: inst = 32'h10408000;
      13602: inst = 32'hc404d67;
      13603: inst = 32'h8220000;
      13604: inst = 32'h10408000;
      13605: inst = 32'hc404d68;
      13606: inst = 32'h8220000;
      13607: inst = 32'h10408000;
      13608: inst = 32'hc404d69;
      13609: inst = 32'h8220000;
      13610: inst = 32'h10408000;
      13611: inst = 32'hc404d6a;
      13612: inst = 32'h8220000;
      13613: inst = 32'h10408000;
      13614: inst = 32'hc404d6b;
      13615: inst = 32'h8220000;
      13616: inst = 32'h10408000;
      13617: inst = 32'hc404d6c;
      13618: inst = 32'h8220000;
      13619: inst = 32'h10408000;
      13620: inst = 32'hc404d6d;
      13621: inst = 32'h8220000;
      13622: inst = 32'h10408000;
      13623: inst = 32'hc404d6e;
      13624: inst = 32'h8220000;
      13625: inst = 32'h10408000;
      13626: inst = 32'hc404d6f;
      13627: inst = 32'h8220000;
      13628: inst = 32'h10408000;
      13629: inst = 32'hc404d70;
      13630: inst = 32'h8220000;
      13631: inst = 32'h10408000;
      13632: inst = 32'hc404d71;
      13633: inst = 32'h8220000;
      13634: inst = 32'h10408000;
      13635: inst = 32'hc404d72;
      13636: inst = 32'h8220000;
      13637: inst = 32'h10408000;
      13638: inst = 32'hc404d73;
      13639: inst = 32'h8220000;
      13640: inst = 32'h10408000;
      13641: inst = 32'hc404d74;
      13642: inst = 32'h8220000;
      13643: inst = 32'h10408000;
      13644: inst = 32'hc404dc0;
      13645: inst = 32'h8220000;
      13646: inst = 32'h10408000;
      13647: inst = 32'hc404dca;
      13648: inst = 32'h8220000;
      13649: inst = 32'h10408000;
      13650: inst = 32'hc404dd4;
      13651: inst = 32'h8220000;
      13652: inst = 32'h10408000;
      13653: inst = 32'hc404e20;
      13654: inst = 32'h8220000;
      13655: inst = 32'h10408000;
      13656: inst = 32'hc404e2a;
      13657: inst = 32'h8220000;
      13658: inst = 32'h10408000;
      13659: inst = 32'hc404e34;
      13660: inst = 32'h8220000;
      13661: inst = 32'h10408000;
      13662: inst = 32'hc404e80;
      13663: inst = 32'h8220000;
      13664: inst = 32'h10408000;
      13665: inst = 32'hc404e8a;
      13666: inst = 32'h8220000;
      13667: inst = 32'h10408000;
      13668: inst = 32'hc404e94;
      13669: inst = 32'h8220000;
      13670: inst = 32'h10408000;
      13671: inst = 32'hc404ee0;
      13672: inst = 32'h8220000;
      13673: inst = 32'h10408000;
      13674: inst = 32'hc404eea;
      13675: inst = 32'h8220000;
      13676: inst = 32'h10408000;
      13677: inst = 32'hc404ef4;
      13678: inst = 32'h8220000;
      13679: inst = 32'h10408000;
      13680: inst = 32'hc404f40;
      13681: inst = 32'h8220000;
      13682: inst = 32'h10408000;
      13683: inst = 32'hc404f4a;
      13684: inst = 32'h8220000;
      13685: inst = 32'h10408000;
      13686: inst = 32'hc404f54;
      13687: inst = 32'h8220000;
      13688: inst = 32'h10408000;
      13689: inst = 32'hc404fa0;
      13690: inst = 32'h8220000;
      13691: inst = 32'h10408000;
      13692: inst = 32'hc404faa;
      13693: inst = 32'h8220000;
      13694: inst = 32'h10408000;
      13695: inst = 32'hc404fb4;
      13696: inst = 32'h8220000;
      13697: inst = 32'h10408000;
      13698: inst = 32'hc405000;
      13699: inst = 32'h8220000;
      13700: inst = 32'h10408000;
      13701: inst = 32'hc40500a;
      13702: inst = 32'h8220000;
      13703: inst = 32'h10408000;
      13704: inst = 32'hc405014;
      13705: inst = 32'h8220000;
      13706: inst = 32'h10408000;
      13707: inst = 32'hc405060;
      13708: inst = 32'h8220000;
      13709: inst = 32'h10408000;
      13710: inst = 32'hc40506a;
      13711: inst = 32'h8220000;
      13712: inst = 32'h10408000;
      13713: inst = 32'hc405074;
      13714: inst = 32'h8220000;
      13715: inst = 32'h10408000;
      13716: inst = 32'hc4050c0;
      13717: inst = 32'h8220000;
      13718: inst = 32'h10408000;
      13719: inst = 32'hc4050ca;
      13720: inst = 32'h8220000;
      13721: inst = 32'h10408000;
      13722: inst = 32'hc4050d4;
      13723: inst = 32'h8220000;
      13724: inst = 32'h10408000;
      13725: inst = 32'hc405120;
      13726: inst = 32'h8220000;
      13727: inst = 32'h10408000;
      13728: inst = 32'hc40512a;
      13729: inst = 32'h8220000;
      13730: inst = 32'h10408000;
      13731: inst = 32'hc405134;
      13732: inst = 32'h8220000;
      13733: inst = 32'h10408000;
      13734: inst = 32'hc405180;
      13735: inst = 32'h8220000;
      13736: inst = 32'h10408000;
      13737: inst = 32'hc40518a;
      13738: inst = 32'h8220000;
      13739: inst = 32'h10408000;
      13740: inst = 32'hc405194;
      13741: inst = 32'h8220000;
      13742: inst = 32'h10408000;
      13743: inst = 32'hc4051a8;
      13744: inst = 32'h8220000;
      13745: inst = 32'h10408000;
      13746: inst = 32'hc4051a9;
      13747: inst = 32'h8220000;
      13748: inst = 32'h10408000;
      13749: inst = 32'hc4051b7;
      13750: inst = 32'h8220000;
      13751: inst = 32'h10408000;
      13752: inst = 32'hc4051e0;
      13753: inst = 32'h8220000;
      13754: inst = 32'h10408000;
      13755: inst = 32'hc4051ea;
      13756: inst = 32'h8220000;
      13757: inst = 32'h10408000;
      13758: inst = 32'hc4051f4;
      13759: inst = 32'h8220000;
      13760: inst = 32'h10408000;
      13761: inst = 32'hc405208;
      13762: inst = 32'h8220000;
      13763: inst = 32'h10408000;
      13764: inst = 32'hc405217;
      13765: inst = 32'h8220000;
      13766: inst = 32'h10408000;
      13767: inst = 32'hc405240;
      13768: inst = 32'h8220000;
      13769: inst = 32'h10408000;
      13770: inst = 32'hc40524a;
      13771: inst = 32'h8220000;
      13772: inst = 32'h10408000;
      13773: inst = 32'hc405254;
      13774: inst = 32'h8220000;
      13775: inst = 32'h10408000;
      13776: inst = 32'hc40525e;
      13777: inst = 32'h8220000;
      13778: inst = 32'h10408000;
      13779: inst = 32'hc405268;
      13780: inst = 32'h8220000;
      13781: inst = 32'h10408000;
      13782: inst = 32'hc405277;
      13783: inst = 32'h8220000;
      13784: inst = 32'h10408000;
      13785: inst = 32'hc405281;
      13786: inst = 32'h8220000;
      13787: inst = 32'h10408000;
      13788: inst = 32'hc4052a0;
      13789: inst = 32'h8220000;
      13790: inst = 32'h10408000;
      13791: inst = 32'hc4052a1;
      13792: inst = 32'h8220000;
      13793: inst = 32'h10408000;
      13794: inst = 32'hc4052a2;
      13795: inst = 32'h8220000;
      13796: inst = 32'h10408000;
      13797: inst = 32'hc4052a3;
      13798: inst = 32'h8220000;
      13799: inst = 32'h10408000;
      13800: inst = 32'hc4052a4;
      13801: inst = 32'h8220000;
      13802: inst = 32'h10408000;
      13803: inst = 32'hc4052a5;
      13804: inst = 32'h8220000;
      13805: inst = 32'h10408000;
      13806: inst = 32'hc4052a6;
      13807: inst = 32'h8220000;
      13808: inst = 32'h10408000;
      13809: inst = 32'hc4052a7;
      13810: inst = 32'h8220000;
      13811: inst = 32'h10408000;
      13812: inst = 32'hc4052a8;
      13813: inst = 32'h8220000;
      13814: inst = 32'h10408000;
      13815: inst = 32'hc4052a9;
      13816: inst = 32'h8220000;
      13817: inst = 32'h10408000;
      13818: inst = 32'hc4052aa;
      13819: inst = 32'h8220000;
      13820: inst = 32'h10408000;
      13821: inst = 32'hc4052ab;
      13822: inst = 32'h8220000;
      13823: inst = 32'h10408000;
      13824: inst = 32'hc4052ac;
      13825: inst = 32'h8220000;
      13826: inst = 32'h10408000;
      13827: inst = 32'hc4052ad;
      13828: inst = 32'h8220000;
      13829: inst = 32'h10408000;
      13830: inst = 32'hc4052ae;
      13831: inst = 32'h8220000;
      13832: inst = 32'h10408000;
      13833: inst = 32'hc4052af;
      13834: inst = 32'h8220000;
      13835: inst = 32'h10408000;
      13836: inst = 32'hc4052b0;
      13837: inst = 32'h8220000;
      13838: inst = 32'h10408000;
      13839: inst = 32'hc4052b1;
      13840: inst = 32'h8220000;
      13841: inst = 32'h10408000;
      13842: inst = 32'hc4052b2;
      13843: inst = 32'h8220000;
      13844: inst = 32'h10408000;
      13845: inst = 32'hc4052b3;
      13846: inst = 32'h8220000;
      13847: inst = 32'h10408000;
      13848: inst = 32'hc4052b4;
      13849: inst = 32'h8220000;
      13850: inst = 32'h10408000;
      13851: inst = 32'hc4052bd;
      13852: inst = 32'h8220000;
      13853: inst = 32'h10408000;
      13854: inst = 32'hc4052be;
      13855: inst = 32'h8220000;
      13856: inst = 32'h10408000;
      13857: inst = 32'hc4052c8;
      13858: inst = 32'h8220000;
      13859: inst = 32'h10408000;
      13860: inst = 32'hc4052d7;
      13861: inst = 32'h8220000;
      13862: inst = 32'h10408000;
      13863: inst = 32'hc4052e1;
      13864: inst = 32'h8220000;
      13865: inst = 32'h10408000;
      13866: inst = 32'hc4052e2;
      13867: inst = 32'h8220000;
      13868: inst = 32'h10408000;
      13869: inst = 32'hc40531c;
      13870: inst = 32'h8220000;
      13871: inst = 32'h10408000;
      13872: inst = 32'hc40531d;
      13873: inst = 32'h8220000;
      13874: inst = 32'h10408000;
      13875: inst = 32'hc40531e;
      13876: inst = 32'h8220000;
      13877: inst = 32'h10408000;
      13878: inst = 32'hc40531f;
      13879: inst = 32'h8220000;
      13880: inst = 32'h10408000;
      13881: inst = 32'hc405320;
      13882: inst = 32'h8220000;
      13883: inst = 32'h10408000;
      13884: inst = 32'hc405326;
      13885: inst = 32'h8220000;
      13886: inst = 32'h10408000;
      13887: inst = 32'hc405327;
      13888: inst = 32'h8220000;
      13889: inst = 32'h10408000;
      13890: inst = 32'hc405328;
      13891: inst = 32'h8220000;
      13892: inst = 32'h10408000;
      13893: inst = 32'hc405337;
      13894: inst = 32'h8220000;
      13895: inst = 32'h10408000;
      13896: inst = 32'hc405338;
      13897: inst = 32'h8220000;
      13898: inst = 32'h10408000;
      13899: inst = 32'hc405339;
      13900: inst = 32'h8220000;
      13901: inst = 32'h10408000;
      13902: inst = 32'hc40533f;
      13903: inst = 32'h8220000;
      13904: inst = 32'h10408000;
      13905: inst = 32'hc405340;
      13906: inst = 32'h8220000;
      13907: inst = 32'h10408000;
      13908: inst = 32'hc405341;
      13909: inst = 32'h8220000;
      13910: inst = 32'h10408000;
      13911: inst = 32'hc405342;
      13912: inst = 32'h8220000;
      13913: inst = 32'h10408000;
      13914: inst = 32'hc405343;
      13915: inst = 32'h8220000;
      13916: inst = 32'h10408000;
      13917: inst = 32'hc40537b;
      13918: inst = 32'h8220000;
      13919: inst = 32'h10408000;
      13920: inst = 32'hc40537c;
      13921: inst = 32'h8220000;
      13922: inst = 32'h10408000;
      13923: inst = 32'hc405386;
      13924: inst = 32'h8220000;
      13925: inst = 32'h10408000;
      13926: inst = 32'hc405387;
      13927: inst = 32'h8220000;
      13928: inst = 32'h10408000;
      13929: inst = 32'hc405388;
      13930: inst = 32'h8220000;
      13931: inst = 32'h10408000;
      13932: inst = 32'hc405397;
      13933: inst = 32'h8220000;
      13934: inst = 32'h10408000;
      13935: inst = 32'hc405398;
      13936: inst = 32'h8220000;
      13937: inst = 32'h10408000;
      13938: inst = 32'hc405399;
      13939: inst = 32'h8220000;
      13940: inst = 32'h10408000;
      13941: inst = 32'hc4053a3;
      13942: inst = 32'h8220000;
      13943: inst = 32'h10408000;
      13944: inst = 32'hc4053a4;
      13945: inst = 32'h8220000;
      13946: inst = 32'h10408000;
      13947: inst = 32'hc4053db;
      13948: inst = 32'h8220000;
      13949: inst = 32'h10408000;
      13950: inst = 32'hc4053e5;
      13951: inst = 32'h8220000;
      13952: inst = 32'h10408000;
      13953: inst = 32'hc4053e6;
      13954: inst = 32'h8220000;
      13955: inst = 32'h10408000;
      13956: inst = 32'hc4053e7;
      13957: inst = 32'h8220000;
      13958: inst = 32'h10408000;
      13959: inst = 32'hc4053f8;
      13960: inst = 32'h8220000;
      13961: inst = 32'h10408000;
      13962: inst = 32'hc4053f9;
      13963: inst = 32'h8220000;
      13964: inst = 32'h10408000;
      13965: inst = 32'hc4053fa;
      13966: inst = 32'h8220000;
      13967: inst = 32'h10408000;
      13968: inst = 32'hc405404;
      13969: inst = 32'h8220000;
      13970: inst = 32'h10408000;
      13971: inst = 32'hc40543a;
      13972: inst = 32'h8220000;
      13973: inst = 32'h10408000;
      13974: inst = 32'hc40543b;
      13975: inst = 32'h8220000;
      13976: inst = 32'h10408000;
      13977: inst = 32'hc405445;
      13978: inst = 32'h8220000;
      13979: inst = 32'h10408000;
      13980: inst = 32'hc405446;
      13981: inst = 32'h8220000;
      13982: inst = 32'h10408000;
      13983: inst = 32'hc405447;
      13984: inst = 32'h8220000;
      13985: inst = 32'h10408000;
      13986: inst = 32'hc405458;
      13987: inst = 32'h8220000;
      13988: inst = 32'h10408000;
      13989: inst = 32'hc405459;
      13990: inst = 32'h8220000;
      13991: inst = 32'h10408000;
      13992: inst = 32'hc40545a;
      13993: inst = 32'h8220000;
      13994: inst = 32'h10408000;
      13995: inst = 32'hc405464;
      13996: inst = 32'h8220000;
      13997: inst = 32'h10408000;
      13998: inst = 32'hc405465;
      13999: inst = 32'h8220000;
      14000: inst = 32'h10408000;
      14001: inst = 32'hc405499;
      14002: inst = 32'h8220000;
      14003: inst = 32'h10408000;
      14004: inst = 32'hc40549a;
      14005: inst = 32'h8220000;
      14006: inst = 32'h10408000;
      14007: inst = 32'hc4054a5;
      14008: inst = 32'h8220000;
      14009: inst = 32'h10408000;
      14010: inst = 32'hc4054a6;
      14011: inst = 32'h8220000;
      14012: inst = 32'h10408000;
      14013: inst = 32'hc4054a7;
      14014: inst = 32'h8220000;
      14015: inst = 32'h10408000;
      14016: inst = 32'hc4054b8;
      14017: inst = 32'h8220000;
      14018: inst = 32'h10408000;
      14019: inst = 32'hc4054b9;
      14020: inst = 32'h8220000;
      14021: inst = 32'h10408000;
      14022: inst = 32'hc4054ba;
      14023: inst = 32'h8220000;
      14024: inst = 32'h10408000;
      14025: inst = 32'hc4054c5;
      14026: inst = 32'h8220000;
      14027: inst = 32'h10408000;
      14028: inst = 32'hc4054c6;
      14029: inst = 32'h8220000;
      14030: inst = 32'h10408000;
      14031: inst = 32'hc4054f8;
      14032: inst = 32'h8220000;
      14033: inst = 32'h10408000;
      14034: inst = 32'hc4054f9;
      14035: inst = 32'h8220000;
      14036: inst = 32'h10408000;
      14037: inst = 32'hc405500;
      14038: inst = 32'h8220000;
      14039: inst = 32'h10408000;
      14040: inst = 32'hc405504;
      14041: inst = 32'h8220000;
      14042: inst = 32'h10408000;
      14043: inst = 32'hc405505;
      14044: inst = 32'h8220000;
      14045: inst = 32'h10408000;
      14046: inst = 32'hc405506;
      14047: inst = 32'h8220000;
      14048: inst = 32'h10408000;
      14049: inst = 32'hc405507;
      14050: inst = 32'h8220000;
      14051: inst = 32'h10408000;
      14052: inst = 32'hc405518;
      14053: inst = 32'h8220000;
      14054: inst = 32'h10408000;
      14055: inst = 32'hc405519;
      14056: inst = 32'h8220000;
      14057: inst = 32'h10408000;
      14058: inst = 32'hc40551a;
      14059: inst = 32'h8220000;
      14060: inst = 32'h10408000;
      14061: inst = 32'hc40551b;
      14062: inst = 32'h8220000;
      14063: inst = 32'h10408000;
      14064: inst = 32'hc40551f;
      14065: inst = 32'h8220000;
      14066: inst = 32'h10408000;
      14067: inst = 32'hc405526;
      14068: inst = 32'h8220000;
      14069: inst = 32'h10408000;
      14070: inst = 32'hc405527;
      14071: inst = 32'h8220000;
      14072: inst = 32'h10408000;
      14073: inst = 32'hc405558;
      14074: inst = 32'h8220000;
      14075: inst = 32'h10408000;
      14076: inst = 32'hc405559;
      14077: inst = 32'h8220000;
      14078: inst = 32'h10408000;
      14079: inst = 32'hc405560;
      14080: inst = 32'h8220000;
      14081: inst = 32'h10408000;
      14082: inst = 32'hc405564;
      14083: inst = 32'h8220000;
      14084: inst = 32'h10408000;
      14085: inst = 32'hc405565;
      14086: inst = 32'h8220000;
      14087: inst = 32'h10408000;
      14088: inst = 32'hc405566;
      14089: inst = 32'h8220000;
      14090: inst = 32'h10408000;
      14091: inst = 32'hc405567;
      14092: inst = 32'h8220000;
      14093: inst = 32'h10408000;
      14094: inst = 32'hc405578;
      14095: inst = 32'h8220000;
      14096: inst = 32'h10408000;
      14097: inst = 32'hc405579;
      14098: inst = 32'h8220000;
      14099: inst = 32'h10408000;
      14100: inst = 32'hc40557a;
      14101: inst = 32'h8220000;
      14102: inst = 32'h10408000;
      14103: inst = 32'hc40557b;
      14104: inst = 32'h8220000;
      14105: inst = 32'h10408000;
      14106: inst = 32'hc40557f;
      14107: inst = 32'h8220000;
      14108: inst = 32'h10408000;
      14109: inst = 32'hc405586;
      14110: inst = 32'h8220000;
      14111: inst = 32'h10408000;
      14112: inst = 32'hc405587;
      14113: inst = 32'h8220000;
      14114: inst = 32'h10408000;
      14115: inst = 32'hc4055b7;
      14116: inst = 32'h8220000;
      14117: inst = 32'h10408000;
      14118: inst = 32'hc4055b8;
      14119: inst = 32'h8220000;
      14120: inst = 32'h10408000;
      14121: inst = 32'hc4055bf;
      14122: inst = 32'h8220000;
      14123: inst = 32'h10408000;
      14124: inst = 32'hc4055c0;
      14125: inst = 32'h8220000;
      14126: inst = 32'h10408000;
      14127: inst = 32'hc4055c4;
      14128: inst = 32'h8220000;
      14129: inst = 32'h10408000;
      14130: inst = 32'hc4055c5;
      14131: inst = 32'h8220000;
      14132: inst = 32'h10408000;
      14133: inst = 32'hc4055c6;
      14134: inst = 32'h8220000;
      14135: inst = 32'h10408000;
      14136: inst = 32'hc4055c7;
      14137: inst = 32'h8220000;
      14138: inst = 32'h10408000;
      14139: inst = 32'hc4055d8;
      14140: inst = 32'h8220000;
      14141: inst = 32'h10408000;
      14142: inst = 32'hc4055d9;
      14143: inst = 32'h8220000;
      14144: inst = 32'h10408000;
      14145: inst = 32'hc4055da;
      14146: inst = 32'h8220000;
      14147: inst = 32'h10408000;
      14148: inst = 32'hc4055db;
      14149: inst = 32'h8220000;
      14150: inst = 32'h10408000;
      14151: inst = 32'hc4055df;
      14152: inst = 32'h8220000;
      14153: inst = 32'h10408000;
      14154: inst = 32'hc4055e0;
      14155: inst = 32'h8220000;
      14156: inst = 32'h10408000;
      14157: inst = 32'hc4055e7;
      14158: inst = 32'h8220000;
      14159: inst = 32'h10408000;
      14160: inst = 32'hc4055e8;
      14161: inst = 32'h8220000;
      14162: inst = 32'h10408000;
      14163: inst = 32'hc405616;
      14164: inst = 32'h8220000;
      14165: inst = 32'h10408000;
      14166: inst = 32'hc405617;
      14167: inst = 32'h8220000;
      14168: inst = 32'h10408000;
      14169: inst = 32'hc40561f;
      14170: inst = 32'h8220000;
      14171: inst = 32'h10408000;
      14172: inst = 32'hc405620;
      14173: inst = 32'h8220000;
      14174: inst = 32'h10408000;
      14175: inst = 32'hc405623;
      14176: inst = 32'h8220000;
      14177: inst = 32'h10408000;
      14178: inst = 32'hc405624;
      14179: inst = 32'h8220000;
      14180: inst = 32'h10408000;
      14181: inst = 32'hc405625;
      14182: inst = 32'h8220000;
      14183: inst = 32'h10408000;
      14184: inst = 32'hc405626;
      14185: inst = 32'h8220000;
      14186: inst = 32'h10408000;
      14187: inst = 32'hc405639;
      14188: inst = 32'h8220000;
      14189: inst = 32'h10408000;
      14190: inst = 32'hc40563a;
      14191: inst = 32'h8220000;
      14192: inst = 32'h10408000;
      14193: inst = 32'hc40563b;
      14194: inst = 32'h8220000;
      14195: inst = 32'h10408000;
      14196: inst = 32'hc40563c;
      14197: inst = 32'h8220000;
      14198: inst = 32'h10408000;
      14199: inst = 32'hc40563f;
      14200: inst = 32'h8220000;
      14201: inst = 32'h10408000;
      14202: inst = 32'hc405640;
      14203: inst = 32'h8220000;
      14204: inst = 32'h10408000;
      14205: inst = 32'hc405648;
      14206: inst = 32'h8220000;
      14207: inst = 32'h10408000;
      14208: inst = 32'hc405649;
      14209: inst = 32'h8220000;
      14210: inst = 32'h10408000;
      14211: inst = 32'hc405675;
      14212: inst = 32'h8220000;
      14213: inst = 32'h10408000;
      14214: inst = 32'hc405676;
      14215: inst = 32'h8220000;
      14216: inst = 32'h10408000;
      14217: inst = 32'hc405677;
      14218: inst = 32'h8220000;
      14219: inst = 32'h10408000;
      14220: inst = 32'hc40567e;
      14221: inst = 32'h8220000;
      14222: inst = 32'h10408000;
      14223: inst = 32'hc40567f;
      14224: inst = 32'h8220000;
      14225: inst = 32'h10408000;
      14226: inst = 32'hc405680;
      14227: inst = 32'h8220000;
      14228: inst = 32'h10408000;
      14229: inst = 32'hc405683;
      14230: inst = 32'h8220000;
      14231: inst = 32'h10408000;
      14232: inst = 32'hc405684;
      14233: inst = 32'h8220000;
      14234: inst = 32'h10408000;
      14235: inst = 32'hc405685;
      14236: inst = 32'h8220000;
      14237: inst = 32'h10408000;
      14238: inst = 32'hc405686;
      14239: inst = 32'h8220000;
      14240: inst = 32'h10408000;
      14241: inst = 32'hc405699;
      14242: inst = 32'h8220000;
      14243: inst = 32'h10408000;
      14244: inst = 32'hc40569a;
      14245: inst = 32'h8220000;
      14246: inst = 32'h10408000;
      14247: inst = 32'hc40569b;
      14248: inst = 32'h8220000;
      14249: inst = 32'h10408000;
      14250: inst = 32'hc40569c;
      14251: inst = 32'h8220000;
      14252: inst = 32'h10408000;
      14253: inst = 32'hc40569f;
      14254: inst = 32'h8220000;
      14255: inst = 32'h10408000;
      14256: inst = 32'hc4056a0;
      14257: inst = 32'h8220000;
      14258: inst = 32'h10408000;
      14259: inst = 32'hc4056a1;
      14260: inst = 32'h8220000;
      14261: inst = 32'h10408000;
      14262: inst = 32'hc4056a8;
      14263: inst = 32'h8220000;
      14264: inst = 32'h10408000;
      14265: inst = 32'hc4056a9;
      14266: inst = 32'h8220000;
      14267: inst = 32'h10408000;
      14268: inst = 32'hc4056aa;
      14269: inst = 32'h8220000;
      14270: inst = 32'h10408000;
      14271: inst = 32'hc4056d4;
      14272: inst = 32'h8220000;
      14273: inst = 32'h10408000;
      14274: inst = 32'hc4056d5;
      14275: inst = 32'h8220000;
      14276: inst = 32'h10408000;
      14277: inst = 32'hc4056d6;
      14278: inst = 32'h8220000;
      14279: inst = 32'h10408000;
      14280: inst = 32'hc4056d7;
      14281: inst = 32'h8220000;
      14282: inst = 32'h10408000;
      14283: inst = 32'hc4056d8;
      14284: inst = 32'h8220000;
      14285: inst = 32'h10408000;
      14286: inst = 32'hc4056d9;
      14287: inst = 32'h8220000;
      14288: inst = 32'h10408000;
      14289: inst = 32'hc4056da;
      14290: inst = 32'h8220000;
      14291: inst = 32'h10408000;
      14292: inst = 32'hc4056db;
      14293: inst = 32'h8220000;
      14294: inst = 32'h10408000;
      14295: inst = 32'hc4056dc;
      14296: inst = 32'h8220000;
      14297: inst = 32'h10408000;
      14298: inst = 32'hc4056dd;
      14299: inst = 32'h8220000;
      14300: inst = 32'h10408000;
      14301: inst = 32'hc4056de;
      14302: inst = 32'h8220000;
      14303: inst = 32'h10408000;
      14304: inst = 32'hc4056df;
      14305: inst = 32'h8220000;
      14306: inst = 32'h10408000;
      14307: inst = 32'hc4056e0;
      14308: inst = 32'h8220000;
      14309: inst = 32'h10408000;
      14310: inst = 32'hc4056e3;
      14311: inst = 32'h8220000;
      14312: inst = 32'h10408000;
      14313: inst = 32'hc4056e4;
      14314: inst = 32'h8220000;
      14315: inst = 32'h10408000;
      14316: inst = 32'hc4056e5;
      14317: inst = 32'h8220000;
      14318: inst = 32'h10408000;
      14319: inst = 32'hc4056e6;
      14320: inst = 32'h8220000;
      14321: inst = 32'h10408000;
      14322: inst = 32'hc4056f9;
      14323: inst = 32'h8220000;
      14324: inst = 32'h10408000;
      14325: inst = 32'hc4056fa;
      14326: inst = 32'h8220000;
      14327: inst = 32'h10408000;
      14328: inst = 32'hc4056fb;
      14329: inst = 32'h8220000;
      14330: inst = 32'h10408000;
      14331: inst = 32'hc4056fc;
      14332: inst = 32'h8220000;
      14333: inst = 32'h10408000;
      14334: inst = 32'hc4056ff;
      14335: inst = 32'h8220000;
      14336: inst = 32'h10408000;
      14337: inst = 32'hc405700;
      14338: inst = 32'h8220000;
      14339: inst = 32'h10408000;
      14340: inst = 32'hc405701;
      14341: inst = 32'h8220000;
      14342: inst = 32'h10408000;
      14343: inst = 32'hc405702;
      14344: inst = 32'h8220000;
      14345: inst = 32'h10408000;
      14346: inst = 32'hc405703;
      14347: inst = 32'h8220000;
      14348: inst = 32'h10408000;
      14349: inst = 32'hc405704;
      14350: inst = 32'h8220000;
      14351: inst = 32'h10408000;
      14352: inst = 32'hc405705;
      14353: inst = 32'h8220000;
      14354: inst = 32'h10408000;
      14355: inst = 32'hc405706;
      14356: inst = 32'h8220000;
      14357: inst = 32'h10408000;
      14358: inst = 32'hc405707;
      14359: inst = 32'h8220000;
      14360: inst = 32'h10408000;
      14361: inst = 32'hc405708;
      14362: inst = 32'h8220000;
      14363: inst = 32'h10408000;
      14364: inst = 32'hc405709;
      14365: inst = 32'h8220000;
      14366: inst = 32'h10408000;
      14367: inst = 32'hc40570a;
      14368: inst = 32'h8220000;
      14369: inst = 32'h10408000;
      14370: inst = 32'hc405734;
      14371: inst = 32'h8220000;
      14372: inst = 32'h10408000;
      14373: inst = 32'hc405735;
      14374: inst = 32'h8220000;
      14375: inst = 32'h10408000;
      14376: inst = 32'hc405736;
      14377: inst = 32'h8220000;
      14378: inst = 32'h10408000;
      14379: inst = 32'hc405737;
      14380: inst = 32'h8220000;
      14381: inst = 32'h10408000;
      14382: inst = 32'hc405738;
      14383: inst = 32'h8220000;
      14384: inst = 32'h10408000;
      14385: inst = 32'hc405739;
      14386: inst = 32'h8220000;
      14387: inst = 32'h10408000;
      14388: inst = 32'hc40573a;
      14389: inst = 32'h8220000;
      14390: inst = 32'h10408000;
      14391: inst = 32'hc40573b;
      14392: inst = 32'h8220000;
      14393: inst = 32'h10408000;
      14394: inst = 32'hc40573c;
      14395: inst = 32'h8220000;
      14396: inst = 32'h10408000;
      14397: inst = 32'hc40573d;
      14398: inst = 32'h8220000;
      14399: inst = 32'h10408000;
      14400: inst = 32'hc40573e;
      14401: inst = 32'h8220000;
      14402: inst = 32'h10408000;
      14403: inst = 32'hc40573f;
      14404: inst = 32'h8220000;
      14405: inst = 32'h10408000;
      14406: inst = 32'hc405740;
      14407: inst = 32'h8220000;
      14408: inst = 32'h10408000;
      14409: inst = 32'hc405742;
      14410: inst = 32'h8220000;
      14411: inst = 32'h10408000;
      14412: inst = 32'hc405743;
      14413: inst = 32'h8220000;
      14414: inst = 32'h10408000;
      14415: inst = 32'hc405744;
      14416: inst = 32'h8220000;
      14417: inst = 32'h10408000;
      14418: inst = 32'hc405745;
      14419: inst = 32'h8220000;
      14420: inst = 32'h10408000;
      14421: inst = 32'hc405746;
      14422: inst = 32'h8220000;
      14423: inst = 32'h10408000;
      14424: inst = 32'hc405759;
      14425: inst = 32'h8220000;
      14426: inst = 32'h10408000;
      14427: inst = 32'hc40575a;
      14428: inst = 32'h8220000;
      14429: inst = 32'h10408000;
      14430: inst = 32'hc40575b;
      14431: inst = 32'h8220000;
      14432: inst = 32'h10408000;
      14433: inst = 32'hc40575c;
      14434: inst = 32'h8220000;
      14435: inst = 32'h10408000;
      14436: inst = 32'hc40575d;
      14437: inst = 32'h8220000;
      14438: inst = 32'h10408000;
      14439: inst = 32'hc40575f;
      14440: inst = 32'h8220000;
      14441: inst = 32'h10408000;
      14442: inst = 32'hc405760;
      14443: inst = 32'h8220000;
      14444: inst = 32'h10408000;
      14445: inst = 32'hc405761;
      14446: inst = 32'h8220000;
      14447: inst = 32'h10408000;
      14448: inst = 32'hc405762;
      14449: inst = 32'h8220000;
      14450: inst = 32'h10408000;
      14451: inst = 32'hc405763;
      14452: inst = 32'h8220000;
      14453: inst = 32'h10408000;
      14454: inst = 32'hc405764;
      14455: inst = 32'h8220000;
      14456: inst = 32'h10408000;
      14457: inst = 32'hc405765;
      14458: inst = 32'h8220000;
      14459: inst = 32'h10408000;
      14460: inst = 32'hc405766;
      14461: inst = 32'h8220000;
      14462: inst = 32'h10408000;
      14463: inst = 32'hc405767;
      14464: inst = 32'h8220000;
      14465: inst = 32'h10408000;
      14466: inst = 32'hc405768;
      14467: inst = 32'h8220000;
      14468: inst = 32'h10408000;
      14469: inst = 32'hc405769;
      14470: inst = 32'h8220000;
      14471: inst = 32'h10408000;
      14472: inst = 32'hc40576a;
      14473: inst = 32'h8220000;
      14474: inst = 32'h10408000;
      14475: inst = 32'hc40576b;
      14476: inst = 32'h8220000;
      14477: inst = 32'h10408000;
      14478: inst = 32'hc405793;
      14479: inst = 32'h8220000;
      14480: inst = 32'h10408000;
      14481: inst = 32'hc405794;
      14482: inst = 32'h8220000;
      14483: inst = 32'h10408000;
      14484: inst = 32'hc405795;
      14485: inst = 32'h8220000;
      14486: inst = 32'h10408000;
      14487: inst = 32'hc405796;
      14488: inst = 32'h8220000;
      14489: inst = 32'h10408000;
      14490: inst = 32'hc405797;
      14491: inst = 32'h8220000;
      14492: inst = 32'h10408000;
      14493: inst = 32'hc405798;
      14494: inst = 32'h8220000;
      14495: inst = 32'h10408000;
      14496: inst = 32'hc405799;
      14497: inst = 32'h8220000;
      14498: inst = 32'h10408000;
      14499: inst = 32'hc40579a;
      14500: inst = 32'h8220000;
      14501: inst = 32'h10408000;
      14502: inst = 32'hc40579b;
      14503: inst = 32'h8220000;
      14504: inst = 32'h10408000;
      14505: inst = 32'hc40579c;
      14506: inst = 32'h8220000;
      14507: inst = 32'h10408000;
      14508: inst = 32'hc40579d;
      14509: inst = 32'h8220000;
      14510: inst = 32'h10408000;
      14511: inst = 32'hc40579e;
      14512: inst = 32'h8220000;
      14513: inst = 32'h10408000;
      14514: inst = 32'hc40579f;
      14515: inst = 32'h8220000;
      14516: inst = 32'h10408000;
      14517: inst = 32'hc4057a0;
      14518: inst = 32'h8220000;
      14519: inst = 32'h10408000;
      14520: inst = 32'hc4057a1;
      14521: inst = 32'h8220000;
      14522: inst = 32'h10408000;
      14523: inst = 32'hc4057a2;
      14524: inst = 32'h8220000;
      14525: inst = 32'h10408000;
      14526: inst = 32'hc4057a3;
      14527: inst = 32'h8220000;
      14528: inst = 32'h10408000;
      14529: inst = 32'hc4057a4;
      14530: inst = 32'h8220000;
      14531: inst = 32'h10408000;
      14532: inst = 32'hc4057a5;
      14533: inst = 32'h8220000;
      14534: inst = 32'h10408000;
      14535: inst = 32'hc4057a6;
      14536: inst = 32'h8220000;
      14537: inst = 32'h10408000;
      14538: inst = 32'hc4057b9;
      14539: inst = 32'h8220000;
      14540: inst = 32'h10408000;
      14541: inst = 32'hc4057ba;
      14542: inst = 32'h8220000;
      14543: inst = 32'h10408000;
      14544: inst = 32'hc4057bb;
      14545: inst = 32'h8220000;
      14546: inst = 32'h10408000;
      14547: inst = 32'hc4057bc;
      14548: inst = 32'h8220000;
      14549: inst = 32'h10408000;
      14550: inst = 32'hc4057bd;
      14551: inst = 32'h8220000;
      14552: inst = 32'h10408000;
      14553: inst = 32'hc4057be;
      14554: inst = 32'h8220000;
      14555: inst = 32'h10408000;
      14556: inst = 32'hc4057bf;
      14557: inst = 32'h8220000;
      14558: inst = 32'h10408000;
      14559: inst = 32'hc4057c0;
      14560: inst = 32'h8220000;
      14561: inst = 32'h10408000;
      14562: inst = 32'hc4057c1;
      14563: inst = 32'h8220000;
      14564: inst = 32'h10408000;
      14565: inst = 32'hc4057c2;
      14566: inst = 32'h8220000;
      14567: inst = 32'h10408000;
      14568: inst = 32'hc4057c3;
      14569: inst = 32'h8220000;
      14570: inst = 32'h10408000;
      14571: inst = 32'hc4057c4;
      14572: inst = 32'h8220000;
      14573: inst = 32'h10408000;
      14574: inst = 32'hc4057c5;
      14575: inst = 32'h8220000;
      14576: inst = 32'h10408000;
      14577: inst = 32'hc4057c6;
      14578: inst = 32'h8220000;
      14579: inst = 32'h10408000;
      14580: inst = 32'hc4057c7;
      14581: inst = 32'h8220000;
      14582: inst = 32'h10408000;
      14583: inst = 32'hc4057c8;
      14584: inst = 32'h8220000;
      14585: inst = 32'h10408000;
      14586: inst = 32'hc4057c9;
      14587: inst = 32'h8220000;
      14588: inst = 32'h10408000;
      14589: inst = 32'hc4057ca;
      14590: inst = 32'h8220000;
      14591: inst = 32'h10408000;
      14592: inst = 32'hc4057cb;
      14593: inst = 32'h8220000;
      14594: inst = 32'h10408000;
      14595: inst = 32'hc4057cc;
      14596: inst = 32'h8220000;
      14597: inst = 32'hc20bdd7;
      14598: inst = 32'h10408000;
      14599: inst = 32'hc404dc1;
      14600: inst = 32'h8220000;
      14601: inst = 32'h10408000;
      14602: inst = 32'hc404dc2;
      14603: inst = 32'h8220000;
      14604: inst = 32'h10408000;
      14605: inst = 32'hc404dc3;
      14606: inst = 32'h8220000;
      14607: inst = 32'h10408000;
      14608: inst = 32'hc404dc4;
      14609: inst = 32'h8220000;
      14610: inst = 32'h10408000;
      14611: inst = 32'hc404dc5;
      14612: inst = 32'h8220000;
      14613: inst = 32'h10408000;
      14614: inst = 32'hc404dc6;
      14615: inst = 32'h8220000;
      14616: inst = 32'h10408000;
      14617: inst = 32'hc404dc7;
      14618: inst = 32'h8220000;
      14619: inst = 32'h10408000;
      14620: inst = 32'hc404dc8;
      14621: inst = 32'h8220000;
      14622: inst = 32'h10408000;
      14623: inst = 32'hc404dc9;
      14624: inst = 32'h8220000;
      14625: inst = 32'h10408000;
      14626: inst = 32'hc404dcb;
      14627: inst = 32'h8220000;
      14628: inst = 32'h10408000;
      14629: inst = 32'hc404dcc;
      14630: inst = 32'h8220000;
      14631: inst = 32'h10408000;
      14632: inst = 32'hc404dcd;
      14633: inst = 32'h8220000;
      14634: inst = 32'h10408000;
      14635: inst = 32'hc404dce;
      14636: inst = 32'h8220000;
      14637: inst = 32'h10408000;
      14638: inst = 32'hc404dcf;
      14639: inst = 32'h8220000;
      14640: inst = 32'h10408000;
      14641: inst = 32'hc404dd0;
      14642: inst = 32'h8220000;
      14643: inst = 32'h10408000;
      14644: inst = 32'hc404dd1;
      14645: inst = 32'h8220000;
      14646: inst = 32'h10408000;
      14647: inst = 32'hc404dd2;
      14648: inst = 32'h8220000;
      14649: inst = 32'h10408000;
      14650: inst = 32'hc404dd3;
      14651: inst = 32'h8220000;
      14652: inst = 32'h10408000;
      14653: inst = 32'hc404e21;
      14654: inst = 32'h8220000;
      14655: inst = 32'h10408000;
      14656: inst = 32'hc404e22;
      14657: inst = 32'h8220000;
      14658: inst = 32'h10408000;
      14659: inst = 32'hc404e23;
      14660: inst = 32'h8220000;
      14661: inst = 32'h10408000;
      14662: inst = 32'hc404e24;
      14663: inst = 32'h8220000;
      14664: inst = 32'h10408000;
      14665: inst = 32'hc404e25;
      14666: inst = 32'h8220000;
      14667: inst = 32'h10408000;
      14668: inst = 32'hc404e26;
      14669: inst = 32'h8220000;
      14670: inst = 32'h10408000;
      14671: inst = 32'hc404e27;
      14672: inst = 32'h8220000;
      14673: inst = 32'h10408000;
      14674: inst = 32'hc404e28;
      14675: inst = 32'h8220000;
      14676: inst = 32'h10408000;
      14677: inst = 32'hc404e29;
      14678: inst = 32'h8220000;
      14679: inst = 32'h10408000;
      14680: inst = 32'hc404e2b;
      14681: inst = 32'h8220000;
      14682: inst = 32'h10408000;
      14683: inst = 32'hc404e2c;
      14684: inst = 32'h8220000;
      14685: inst = 32'h10408000;
      14686: inst = 32'hc404e2d;
      14687: inst = 32'h8220000;
      14688: inst = 32'h10408000;
      14689: inst = 32'hc404e2e;
      14690: inst = 32'h8220000;
      14691: inst = 32'h10408000;
      14692: inst = 32'hc404e2f;
      14693: inst = 32'h8220000;
      14694: inst = 32'h10408000;
      14695: inst = 32'hc404e30;
      14696: inst = 32'h8220000;
      14697: inst = 32'h10408000;
      14698: inst = 32'hc404e31;
      14699: inst = 32'h8220000;
      14700: inst = 32'h10408000;
      14701: inst = 32'hc404e32;
      14702: inst = 32'h8220000;
      14703: inst = 32'h10408000;
      14704: inst = 32'hc404e33;
      14705: inst = 32'h8220000;
      14706: inst = 32'h10408000;
      14707: inst = 32'hc404e81;
      14708: inst = 32'h8220000;
      14709: inst = 32'h10408000;
      14710: inst = 32'hc404e82;
      14711: inst = 32'h8220000;
      14712: inst = 32'h10408000;
      14713: inst = 32'hc404e83;
      14714: inst = 32'h8220000;
      14715: inst = 32'h10408000;
      14716: inst = 32'hc404e84;
      14717: inst = 32'h8220000;
      14718: inst = 32'h10408000;
      14719: inst = 32'hc404e85;
      14720: inst = 32'h8220000;
      14721: inst = 32'h10408000;
      14722: inst = 32'hc404e86;
      14723: inst = 32'h8220000;
      14724: inst = 32'h10408000;
      14725: inst = 32'hc404e87;
      14726: inst = 32'h8220000;
      14727: inst = 32'h10408000;
      14728: inst = 32'hc404e88;
      14729: inst = 32'h8220000;
      14730: inst = 32'h10408000;
      14731: inst = 32'hc404e89;
      14732: inst = 32'h8220000;
      14733: inst = 32'h10408000;
      14734: inst = 32'hc404e8b;
      14735: inst = 32'h8220000;
      14736: inst = 32'h10408000;
      14737: inst = 32'hc404e8c;
      14738: inst = 32'h8220000;
      14739: inst = 32'h10408000;
      14740: inst = 32'hc404e8d;
      14741: inst = 32'h8220000;
      14742: inst = 32'h10408000;
      14743: inst = 32'hc404e8e;
      14744: inst = 32'h8220000;
      14745: inst = 32'h10408000;
      14746: inst = 32'hc404e8f;
      14747: inst = 32'h8220000;
      14748: inst = 32'h10408000;
      14749: inst = 32'hc404e90;
      14750: inst = 32'h8220000;
      14751: inst = 32'h10408000;
      14752: inst = 32'hc404e91;
      14753: inst = 32'h8220000;
      14754: inst = 32'h10408000;
      14755: inst = 32'hc404e92;
      14756: inst = 32'h8220000;
      14757: inst = 32'h10408000;
      14758: inst = 32'hc404e93;
      14759: inst = 32'h8220000;
      14760: inst = 32'h10408000;
      14761: inst = 32'hc404ee1;
      14762: inst = 32'h8220000;
      14763: inst = 32'h10408000;
      14764: inst = 32'hc404ee2;
      14765: inst = 32'h8220000;
      14766: inst = 32'h10408000;
      14767: inst = 32'hc404ee3;
      14768: inst = 32'h8220000;
      14769: inst = 32'h10408000;
      14770: inst = 32'hc404ee4;
      14771: inst = 32'h8220000;
      14772: inst = 32'h10408000;
      14773: inst = 32'hc404ee5;
      14774: inst = 32'h8220000;
      14775: inst = 32'h10408000;
      14776: inst = 32'hc404ee6;
      14777: inst = 32'h8220000;
      14778: inst = 32'h10408000;
      14779: inst = 32'hc404ee7;
      14780: inst = 32'h8220000;
      14781: inst = 32'h10408000;
      14782: inst = 32'hc404ee8;
      14783: inst = 32'h8220000;
      14784: inst = 32'h10408000;
      14785: inst = 32'hc404ee9;
      14786: inst = 32'h8220000;
      14787: inst = 32'h10408000;
      14788: inst = 32'hc404eeb;
      14789: inst = 32'h8220000;
      14790: inst = 32'h10408000;
      14791: inst = 32'hc404eec;
      14792: inst = 32'h8220000;
      14793: inst = 32'h10408000;
      14794: inst = 32'hc404eed;
      14795: inst = 32'h8220000;
      14796: inst = 32'h10408000;
      14797: inst = 32'hc404eee;
      14798: inst = 32'h8220000;
      14799: inst = 32'h10408000;
      14800: inst = 32'hc404eef;
      14801: inst = 32'h8220000;
      14802: inst = 32'h10408000;
      14803: inst = 32'hc404ef0;
      14804: inst = 32'h8220000;
      14805: inst = 32'h10408000;
      14806: inst = 32'hc404ef1;
      14807: inst = 32'h8220000;
      14808: inst = 32'h10408000;
      14809: inst = 32'hc404ef2;
      14810: inst = 32'h8220000;
      14811: inst = 32'h10408000;
      14812: inst = 32'hc404ef3;
      14813: inst = 32'h8220000;
      14814: inst = 32'h10408000;
      14815: inst = 32'hc404f41;
      14816: inst = 32'h8220000;
      14817: inst = 32'h10408000;
      14818: inst = 32'hc404f42;
      14819: inst = 32'h8220000;
      14820: inst = 32'h10408000;
      14821: inst = 32'hc404f43;
      14822: inst = 32'h8220000;
      14823: inst = 32'h10408000;
      14824: inst = 32'hc404f44;
      14825: inst = 32'h8220000;
      14826: inst = 32'h10408000;
      14827: inst = 32'hc404f45;
      14828: inst = 32'h8220000;
      14829: inst = 32'h10408000;
      14830: inst = 32'hc404f46;
      14831: inst = 32'h8220000;
      14832: inst = 32'h10408000;
      14833: inst = 32'hc404f47;
      14834: inst = 32'h8220000;
      14835: inst = 32'h10408000;
      14836: inst = 32'hc404f48;
      14837: inst = 32'h8220000;
      14838: inst = 32'h10408000;
      14839: inst = 32'hc404f49;
      14840: inst = 32'h8220000;
      14841: inst = 32'h10408000;
      14842: inst = 32'hc404f4b;
      14843: inst = 32'h8220000;
      14844: inst = 32'h10408000;
      14845: inst = 32'hc404f4c;
      14846: inst = 32'h8220000;
      14847: inst = 32'h10408000;
      14848: inst = 32'hc404f4d;
      14849: inst = 32'h8220000;
      14850: inst = 32'h10408000;
      14851: inst = 32'hc404f4e;
      14852: inst = 32'h8220000;
      14853: inst = 32'h10408000;
      14854: inst = 32'hc404f4f;
      14855: inst = 32'h8220000;
      14856: inst = 32'h10408000;
      14857: inst = 32'hc404f50;
      14858: inst = 32'h8220000;
      14859: inst = 32'h10408000;
      14860: inst = 32'hc404f51;
      14861: inst = 32'h8220000;
      14862: inst = 32'h10408000;
      14863: inst = 32'hc404f52;
      14864: inst = 32'h8220000;
      14865: inst = 32'h10408000;
      14866: inst = 32'hc404f53;
      14867: inst = 32'h8220000;
      14868: inst = 32'h10408000;
      14869: inst = 32'hc404fa1;
      14870: inst = 32'h8220000;
      14871: inst = 32'h10408000;
      14872: inst = 32'hc404fa2;
      14873: inst = 32'h8220000;
      14874: inst = 32'h10408000;
      14875: inst = 32'hc404fa3;
      14876: inst = 32'h8220000;
      14877: inst = 32'h10408000;
      14878: inst = 32'hc404fa4;
      14879: inst = 32'h8220000;
      14880: inst = 32'h10408000;
      14881: inst = 32'hc404fa5;
      14882: inst = 32'h8220000;
      14883: inst = 32'h10408000;
      14884: inst = 32'hc404fa6;
      14885: inst = 32'h8220000;
      14886: inst = 32'h10408000;
      14887: inst = 32'hc404fa7;
      14888: inst = 32'h8220000;
      14889: inst = 32'h10408000;
      14890: inst = 32'hc404fa9;
      14891: inst = 32'h8220000;
      14892: inst = 32'h10408000;
      14893: inst = 32'hc404fab;
      14894: inst = 32'h8220000;
      14895: inst = 32'h10408000;
      14896: inst = 32'hc404fad;
      14897: inst = 32'h8220000;
      14898: inst = 32'h10408000;
      14899: inst = 32'hc404fae;
      14900: inst = 32'h8220000;
      14901: inst = 32'h10408000;
      14902: inst = 32'hc404faf;
      14903: inst = 32'h8220000;
      14904: inst = 32'h10408000;
      14905: inst = 32'hc404fb0;
      14906: inst = 32'h8220000;
      14907: inst = 32'h10408000;
      14908: inst = 32'hc404fb1;
      14909: inst = 32'h8220000;
      14910: inst = 32'h10408000;
      14911: inst = 32'hc404fb2;
      14912: inst = 32'h8220000;
      14913: inst = 32'h10408000;
      14914: inst = 32'hc404fb3;
      14915: inst = 32'h8220000;
      14916: inst = 32'h10408000;
      14917: inst = 32'hc405001;
      14918: inst = 32'h8220000;
      14919: inst = 32'h10408000;
      14920: inst = 32'hc405002;
      14921: inst = 32'h8220000;
      14922: inst = 32'h10408000;
      14923: inst = 32'hc405003;
      14924: inst = 32'h8220000;
      14925: inst = 32'h10408000;
      14926: inst = 32'hc405004;
      14927: inst = 32'h8220000;
      14928: inst = 32'h10408000;
      14929: inst = 32'hc405005;
      14930: inst = 32'h8220000;
      14931: inst = 32'h10408000;
      14932: inst = 32'hc405006;
      14933: inst = 32'h8220000;
      14934: inst = 32'h10408000;
      14935: inst = 32'hc405007;
      14936: inst = 32'h8220000;
      14937: inst = 32'h10408000;
      14938: inst = 32'hc405009;
      14939: inst = 32'h8220000;
      14940: inst = 32'h10408000;
      14941: inst = 32'hc40500b;
      14942: inst = 32'h8220000;
      14943: inst = 32'h10408000;
      14944: inst = 32'hc40500d;
      14945: inst = 32'h8220000;
      14946: inst = 32'h10408000;
      14947: inst = 32'hc40500e;
      14948: inst = 32'h8220000;
      14949: inst = 32'h10408000;
      14950: inst = 32'hc40500f;
      14951: inst = 32'h8220000;
      14952: inst = 32'h10408000;
      14953: inst = 32'hc405010;
      14954: inst = 32'h8220000;
      14955: inst = 32'h10408000;
      14956: inst = 32'hc405011;
      14957: inst = 32'h8220000;
      14958: inst = 32'h10408000;
      14959: inst = 32'hc405012;
      14960: inst = 32'h8220000;
      14961: inst = 32'h10408000;
      14962: inst = 32'hc405013;
      14963: inst = 32'h8220000;
      14964: inst = 32'h10408000;
      14965: inst = 32'hc405061;
      14966: inst = 32'h8220000;
      14967: inst = 32'h10408000;
      14968: inst = 32'hc405062;
      14969: inst = 32'h8220000;
      14970: inst = 32'h10408000;
      14971: inst = 32'hc405063;
      14972: inst = 32'h8220000;
      14973: inst = 32'h10408000;
      14974: inst = 32'hc405064;
      14975: inst = 32'h8220000;
      14976: inst = 32'h10408000;
      14977: inst = 32'hc405065;
      14978: inst = 32'h8220000;
      14979: inst = 32'h10408000;
      14980: inst = 32'hc405066;
      14981: inst = 32'h8220000;
      14982: inst = 32'h10408000;
      14983: inst = 32'hc405067;
      14984: inst = 32'h8220000;
      14985: inst = 32'h10408000;
      14986: inst = 32'hc405068;
      14987: inst = 32'h8220000;
      14988: inst = 32'h10408000;
      14989: inst = 32'hc405069;
      14990: inst = 32'h8220000;
      14991: inst = 32'h10408000;
      14992: inst = 32'hc40506b;
      14993: inst = 32'h8220000;
      14994: inst = 32'h10408000;
      14995: inst = 32'hc40506c;
      14996: inst = 32'h8220000;
      14997: inst = 32'h10408000;
      14998: inst = 32'hc40506d;
      14999: inst = 32'h8220000;
      15000: inst = 32'h10408000;
      15001: inst = 32'hc40506e;
      15002: inst = 32'h8220000;
      15003: inst = 32'h10408000;
      15004: inst = 32'hc40506f;
      15005: inst = 32'h8220000;
      15006: inst = 32'h10408000;
      15007: inst = 32'hc405070;
      15008: inst = 32'h8220000;
      15009: inst = 32'h10408000;
      15010: inst = 32'hc405071;
      15011: inst = 32'h8220000;
      15012: inst = 32'h10408000;
      15013: inst = 32'hc405072;
      15014: inst = 32'h8220000;
      15015: inst = 32'h10408000;
      15016: inst = 32'hc405073;
      15017: inst = 32'h8220000;
      15018: inst = 32'h10408000;
      15019: inst = 32'hc4050c1;
      15020: inst = 32'h8220000;
      15021: inst = 32'h10408000;
      15022: inst = 32'hc4050c2;
      15023: inst = 32'h8220000;
      15024: inst = 32'h10408000;
      15025: inst = 32'hc4050c3;
      15026: inst = 32'h8220000;
      15027: inst = 32'h10408000;
      15028: inst = 32'hc4050c4;
      15029: inst = 32'h8220000;
      15030: inst = 32'h10408000;
      15031: inst = 32'hc4050c5;
      15032: inst = 32'h8220000;
      15033: inst = 32'h10408000;
      15034: inst = 32'hc4050c6;
      15035: inst = 32'h8220000;
      15036: inst = 32'h10408000;
      15037: inst = 32'hc4050c7;
      15038: inst = 32'h8220000;
      15039: inst = 32'h10408000;
      15040: inst = 32'hc4050c8;
      15041: inst = 32'h8220000;
      15042: inst = 32'h10408000;
      15043: inst = 32'hc4050c9;
      15044: inst = 32'h8220000;
      15045: inst = 32'h10408000;
      15046: inst = 32'hc4050cb;
      15047: inst = 32'h8220000;
      15048: inst = 32'h10408000;
      15049: inst = 32'hc4050cc;
      15050: inst = 32'h8220000;
      15051: inst = 32'h10408000;
      15052: inst = 32'hc4050cd;
      15053: inst = 32'h8220000;
      15054: inst = 32'h10408000;
      15055: inst = 32'hc4050ce;
      15056: inst = 32'h8220000;
      15057: inst = 32'h10408000;
      15058: inst = 32'hc4050cf;
      15059: inst = 32'h8220000;
      15060: inst = 32'h10408000;
      15061: inst = 32'hc4050d0;
      15062: inst = 32'h8220000;
      15063: inst = 32'h10408000;
      15064: inst = 32'hc4050d1;
      15065: inst = 32'h8220000;
      15066: inst = 32'h10408000;
      15067: inst = 32'hc4050d2;
      15068: inst = 32'h8220000;
      15069: inst = 32'h10408000;
      15070: inst = 32'hc4050d3;
      15071: inst = 32'h8220000;
      15072: inst = 32'h10408000;
      15073: inst = 32'hc405121;
      15074: inst = 32'h8220000;
      15075: inst = 32'h10408000;
      15076: inst = 32'hc405122;
      15077: inst = 32'h8220000;
      15078: inst = 32'h10408000;
      15079: inst = 32'hc405123;
      15080: inst = 32'h8220000;
      15081: inst = 32'h10408000;
      15082: inst = 32'hc405124;
      15083: inst = 32'h8220000;
      15084: inst = 32'h10408000;
      15085: inst = 32'hc405125;
      15086: inst = 32'h8220000;
      15087: inst = 32'h10408000;
      15088: inst = 32'hc405126;
      15089: inst = 32'h8220000;
      15090: inst = 32'h10408000;
      15091: inst = 32'hc405127;
      15092: inst = 32'h8220000;
      15093: inst = 32'h10408000;
      15094: inst = 32'hc405128;
      15095: inst = 32'h8220000;
      15096: inst = 32'h10408000;
      15097: inst = 32'hc405129;
      15098: inst = 32'h8220000;
      15099: inst = 32'h10408000;
      15100: inst = 32'hc40512b;
      15101: inst = 32'h8220000;
      15102: inst = 32'h10408000;
      15103: inst = 32'hc40512c;
      15104: inst = 32'h8220000;
      15105: inst = 32'h10408000;
      15106: inst = 32'hc40512d;
      15107: inst = 32'h8220000;
      15108: inst = 32'h10408000;
      15109: inst = 32'hc40512e;
      15110: inst = 32'h8220000;
      15111: inst = 32'h10408000;
      15112: inst = 32'hc40512f;
      15113: inst = 32'h8220000;
      15114: inst = 32'h10408000;
      15115: inst = 32'hc405130;
      15116: inst = 32'h8220000;
      15117: inst = 32'h10408000;
      15118: inst = 32'hc405131;
      15119: inst = 32'h8220000;
      15120: inst = 32'h10408000;
      15121: inst = 32'hc405132;
      15122: inst = 32'h8220000;
      15123: inst = 32'h10408000;
      15124: inst = 32'hc405133;
      15125: inst = 32'h8220000;
      15126: inst = 32'h10408000;
      15127: inst = 32'hc405181;
      15128: inst = 32'h8220000;
      15129: inst = 32'h10408000;
      15130: inst = 32'hc405182;
      15131: inst = 32'h8220000;
      15132: inst = 32'h10408000;
      15133: inst = 32'hc405183;
      15134: inst = 32'h8220000;
      15135: inst = 32'h10408000;
      15136: inst = 32'hc405184;
      15137: inst = 32'h8220000;
      15138: inst = 32'h10408000;
      15139: inst = 32'hc405185;
      15140: inst = 32'h8220000;
      15141: inst = 32'h10408000;
      15142: inst = 32'hc405186;
      15143: inst = 32'h8220000;
      15144: inst = 32'h10408000;
      15145: inst = 32'hc405187;
      15146: inst = 32'h8220000;
      15147: inst = 32'h10408000;
      15148: inst = 32'hc405188;
      15149: inst = 32'h8220000;
      15150: inst = 32'h10408000;
      15151: inst = 32'hc405189;
      15152: inst = 32'h8220000;
      15153: inst = 32'h10408000;
      15154: inst = 32'hc40518b;
      15155: inst = 32'h8220000;
      15156: inst = 32'h10408000;
      15157: inst = 32'hc40518c;
      15158: inst = 32'h8220000;
      15159: inst = 32'h10408000;
      15160: inst = 32'hc40518d;
      15161: inst = 32'h8220000;
      15162: inst = 32'h10408000;
      15163: inst = 32'hc40518e;
      15164: inst = 32'h8220000;
      15165: inst = 32'h10408000;
      15166: inst = 32'hc40518f;
      15167: inst = 32'h8220000;
      15168: inst = 32'h10408000;
      15169: inst = 32'hc405190;
      15170: inst = 32'h8220000;
      15171: inst = 32'h10408000;
      15172: inst = 32'hc405191;
      15173: inst = 32'h8220000;
      15174: inst = 32'h10408000;
      15175: inst = 32'hc405192;
      15176: inst = 32'h8220000;
      15177: inst = 32'h10408000;
      15178: inst = 32'hc405193;
      15179: inst = 32'h8220000;
      15180: inst = 32'h10408000;
      15181: inst = 32'hc4051e1;
      15182: inst = 32'h8220000;
      15183: inst = 32'h10408000;
      15184: inst = 32'hc4051e2;
      15185: inst = 32'h8220000;
      15186: inst = 32'h10408000;
      15187: inst = 32'hc4051e3;
      15188: inst = 32'h8220000;
      15189: inst = 32'h10408000;
      15190: inst = 32'hc4051e4;
      15191: inst = 32'h8220000;
      15192: inst = 32'h10408000;
      15193: inst = 32'hc4051e5;
      15194: inst = 32'h8220000;
      15195: inst = 32'h10408000;
      15196: inst = 32'hc4051e6;
      15197: inst = 32'h8220000;
      15198: inst = 32'h10408000;
      15199: inst = 32'hc4051e7;
      15200: inst = 32'h8220000;
      15201: inst = 32'h10408000;
      15202: inst = 32'hc4051e8;
      15203: inst = 32'h8220000;
      15204: inst = 32'h10408000;
      15205: inst = 32'hc4051e9;
      15206: inst = 32'h8220000;
      15207: inst = 32'h10408000;
      15208: inst = 32'hc4051eb;
      15209: inst = 32'h8220000;
      15210: inst = 32'h10408000;
      15211: inst = 32'hc4051ec;
      15212: inst = 32'h8220000;
      15213: inst = 32'h10408000;
      15214: inst = 32'hc4051ed;
      15215: inst = 32'h8220000;
      15216: inst = 32'h10408000;
      15217: inst = 32'hc4051ee;
      15218: inst = 32'h8220000;
      15219: inst = 32'h10408000;
      15220: inst = 32'hc4051ef;
      15221: inst = 32'h8220000;
      15222: inst = 32'h10408000;
      15223: inst = 32'hc4051f0;
      15224: inst = 32'h8220000;
      15225: inst = 32'h10408000;
      15226: inst = 32'hc4051f1;
      15227: inst = 32'h8220000;
      15228: inst = 32'h10408000;
      15229: inst = 32'hc4051f2;
      15230: inst = 32'h8220000;
      15231: inst = 32'h10408000;
      15232: inst = 32'hc4051f3;
      15233: inst = 32'h8220000;
      15234: inst = 32'h10408000;
      15235: inst = 32'hc405241;
      15236: inst = 32'h8220000;
      15237: inst = 32'h10408000;
      15238: inst = 32'hc405242;
      15239: inst = 32'h8220000;
      15240: inst = 32'h10408000;
      15241: inst = 32'hc405243;
      15242: inst = 32'h8220000;
      15243: inst = 32'h10408000;
      15244: inst = 32'hc405244;
      15245: inst = 32'h8220000;
      15246: inst = 32'h10408000;
      15247: inst = 32'hc405245;
      15248: inst = 32'h8220000;
      15249: inst = 32'h10408000;
      15250: inst = 32'hc405246;
      15251: inst = 32'h8220000;
      15252: inst = 32'h10408000;
      15253: inst = 32'hc405247;
      15254: inst = 32'h8220000;
      15255: inst = 32'h10408000;
      15256: inst = 32'hc405248;
      15257: inst = 32'h8220000;
      15258: inst = 32'h10408000;
      15259: inst = 32'hc405249;
      15260: inst = 32'h8220000;
      15261: inst = 32'h10408000;
      15262: inst = 32'hc40524b;
      15263: inst = 32'h8220000;
      15264: inst = 32'h10408000;
      15265: inst = 32'hc40524c;
      15266: inst = 32'h8220000;
      15267: inst = 32'h10408000;
      15268: inst = 32'hc40524d;
      15269: inst = 32'h8220000;
      15270: inst = 32'h10408000;
      15271: inst = 32'hc40524e;
      15272: inst = 32'h8220000;
      15273: inst = 32'h10408000;
      15274: inst = 32'hc40524f;
      15275: inst = 32'h8220000;
      15276: inst = 32'h10408000;
      15277: inst = 32'hc405250;
      15278: inst = 32'h8220000;
      15279: inst = 32'h10408000;
      15280: inst = 32'hc405251;
      15281: inst = 32'h8220000;
      15282: inst = 32'h10408000;
      15283: inst = 32'hc405252;
      15284: inst = 32'h8220000;
      15285: inst = 32'h10408000;
      15286: inst = 32'hc405253;
      15287: inst = 32'h8220000;
      15288: inst = 32'hc20bd73;
      15289: inst = 32'h10408000;
      15290: inst = 32'hc404e9f;
      15291: inst = 32'h8220000;
      15292: inst = 32'h10408000;
      15293: inst = 32'hc404ec0;
      15294: inst = 32'h8220000;
      15295: inst = 32'hc205aed;
      15296: inst = 32'h10408000;
      15297: inst = 32'hc404ea0;
      15298: inst = 32'h8220000;
      15299: inst = 32'h10408000;
      15300: inst = 32'hc404ea1;
      15301: inst = 32'h8220000;
      15302: inst = 32'h10408000;
      15303: inst = 32'hc404ea2;
      15304: inst = 32'h8220000;
      15305: inst = 32'h10408000;
      15306: inst = 32'hc404ea3;
      15307: inst = 32'h8220000;
      15308: inst = 32'h10408000;
      15309: inst = 32'hc404ea4;
      15310: inst = 32'h8220000;
      15311: inst = 32'h10408000;
      15312: inst = 32'hc404ebb;
      15313: inst = 32'h8220000;
      15314: inst = 32'h10408000;
      15315: inst = 32'hc404ebc;
      15316: inst = 32'h8220000;
      15317: inst = 32'h10408000;
      15318: inst = 32'hc404ebd;
      15319: inst = 32'h8220000;
      15320: inst = 32'h10408000;
      15321: inst = 32'hc404ebe;
      15322: inst = 32'h8220000;
      15323: inst = 32'h10408000;
      15324: inst = 32'hc404ebf;
      15325: inst = 32'h8220000;
      15326: inst = 32'h10408000;
      15327: inst = 32'hc404f00;
      15328: inst = 32'h8220000;
      15329: inst = 32'h10408000;
      15330: inst = 32'hc404f01;
      15331: inst = 32'h8220000;
      15332: inst = 32'h10408000;
      15333: inst = 32'hc404f02;
      15334: inst = 32'h8220000;
      15335: inst = 32'h10408000;
      15336: inst = 32'hc404f03;
      15337: inst = 32'h8220000;
      15338: inst = 32'h10408000;
      15339: inst = 32'hc404f04;
      15340: inst = 32'h8220000;
      15341: inst = 32'h10408000;
      15342: inst = 32'hc404f05;
      15343: inst = 32'h8220000;
      15344: inst = 32'h10408000;
      15345: inst = 32'hc404f1a;
      15346: inst = 32'h8220000;
      15347: inst = 32'h10408000;
      15348: inst = 32'hc404f1b;
      15349: inst = 32'h8220000;
      15350: inst = 32'h10408000;
      15351: inst = 32'hc404f1c;
      15352: inst = 32'h8220000;
      15353: inst = 32'h10408000;
      15354: inst = 32'hc404f1d;
      15355: inst = 32'h8220000;
      15356: inst = 32'h10408000;
      15357: inst = 32'hc404f1e;
      15358: inst = 32'h8220000;
      15359: inst = 32'h10408000;
      15360: inst = 32'hc404f1f;
      15361: inst = 32'h8220000;
      15362: inst = 32'h10408000;
      15363: inst = 32'hc404f60;
      15364: inst = 32'h8220000;
      15365: inst = 32'h10408000;
      15366: inst = 32'hc404f61;
      15367: inst = 32'h8220000;
      15368: inst = 32'h10408000;
      15369: inst = 32'hc404f62;
      15370: inst = 32'h8220000;
      15371: inst = 32'h10408000;
      15372: inst = 32'hc404f63;
      15373: inst = 32'h8220000;
      15374: inst = 32'h10408000;
      15375: inst = 32'hc404f64;
      15376: inst = 32'h8220000;
      15377: inst = 32'h10408000;
      15378: inst = 32'hc404f65;
      15379: inst = 32'h8220000;
      15380: inst = 32'h10408000;
      15381: inst = 32'hc404f66;
      15382: inst = 32'h8220000;
      15383: inst = 32'h10408000;
      15384: inst = 32'hc404f67;
      15385: inst = 32'h8220000;
      15386: inst = 32'h10408000;
      15387: inst = 32'hc404f78;
      15388: inst = 32'h8220000;
      15389: inst = 32'h10408000;
      15390: inst = 32'hc404f79;
      15391: inst = 32'h8220000;
      15392: inst = 32'h10408000;
      15393: inst = 32'hc404f7a;
      15394: inst = 32'h8220000;
      15395: inst = 32'h10408000;
      15396: inst = 32'hc404f7b;
      15397: inst = 32'h8220000;
      15398: inst = 32'h10408000;
      15399: inst = 32'hc404f7c;
      15400: inst = 32'h8220000;
      15401: inst = 32'h10408000;
      15402: inst = 32'hc404f7d;
      15403: inst = 32'h8220000;
      15404: inst = 32'h10408000;
      15405: inst = 32'hc404f7e;
      15406: inst = 32'h8220000;
      15407: inst = 32'h10408000;
      15408: inst = 32'hc404f7f;
      15409: inst = 32'h8220000;
      15410: inst = 32'h10408000;
      15411: inst = 32'hc404fc0;
      15412: inst = 32'h8220000;
      15413: inst = 32'h10408000;
      15414: inst = 32'hc404fc1;
      15415: inst = 32'h8220000;
      15416: inst = 32'h10408000;
      15417: inst = 32'hc404fc2;
      15418: inst = 32'h8220000;
      15419: inst = 32'h10408000;
      15420: inst = 32'hc404fc3;
      15421: inst = 32'h8220000;
      15422: inst = 32'h10408000;
      15423: inst = 32'hc404fc4;
      15424: inst = 32'h8220000;
      15425: inst = 32'h10408000;
      15426: inst = 32'hc404fc6;
      15427: inst = 32'h8220000;
      15428: inst = 32'h10408000;
      15429: inst = 32'hc404fc7;
      15430: inst = 32'h8220000;
      15431: inst = 32'h10408000;
      15432: inst = 32'hc404fd8;
      15433: inst = 32'h8220000;
      15434: inst = 32'h10408000;
      15435: inst = 32'hc404fd9;
      15436: inst = 32'h8220000;
      15437: inst = 32'h10408000;
      15438: inst = 32'hc404fdb;
      15439: inst = 32'h8220000;
      15440: inst = 32'h10408000;
      15441: inst = 32'hc404fdc;
      15442: inst = 32'h8220000;
      15443: inst = 32'h10408000;
      15444: inst = 32'hc404fdd;
      15445: inst = 32'h8220000;
      15446: inst = 32'h10408000;
      15447: inst = 32'hc404fde;
      15448: inst = 32'h8220000;
      15449: inst = 32'h10408000;
      15450: inst = 32'hc404fdf;
      15451: inst = 32'h8220000;
      15452: inst = 32'h10408000;
      15453: inst = 32'hc405020;
      15454: inst = 32'h8220000;
      15455: inst = 32'h10408000;
      15456: inst = 32'hc405021;
      15457: inst = 32'h8220000;
      15458: inst = 32'h10408000;
      15459: inst = 32'hc405022;
      15460: inst = 32'h8220000;
      15461: inst = 32'h10408000;
      15462: inst = 32'hc405023;
      15463: inst = 32'h8220000;
      15464: inst = 32'h10408000;
      15465: inst = 32'hc405026;
      15466: inst = 32'h8220000;
      15467: inst = 32'h10408000;
      15468: inst = 32'hc405027;
      15469: inst = 32'h8220000;
      15470: inst = 32'h10408000;
      15471: inst = 32'hc405038;
      15472: inst = 32'h8220000;
      15473: inst = 32'h10408000;
      15474: inst = 32'hc405039;
      15475: inst = 32'h8220000;
      15476: inst = 32'h10408000;
      15477: inst = 32'hc40503c;
      15478: inst = 32'h8220000;
      15479: inst = 32'h10408000;
      15480: inst = 32'hc40503d;
      15481: inst = 32'h8220000;
      15482: inst = 32'h10408000;
      15483: inst = 32'hc40503e;
      15484: inst = 32'h8220000;
      15485: inst = 32'h10408000;
      15486: inst = 32'hc40503f;
      15487: inst = 32'h8220000;
      15488: inst = 32'h10408000;
      15489: inst = 32'hc40507f;
      15490: inst = 32'h8220000;
      15491: inst = 32'h10408000;
      15492: inst = 32'hc405080;
      15493: inst = 32'h8220000;
      15494: inst = 32'h10408000;
      15495: inst = 32'hc405081;
      15496: inst = 32'h8220000;
      15497: inst = 32'h10408000;
      15498: inst = 32'hc405082;
      15499: inst = 32'h8220000;
      15500: inst = 32'h10408000;
      15501: inst = 32'hc405086;
      15502: inst = 32'h8220000;
      15503: inst = 32'h10408000;
      15504: inst = 32'hc405087;
      15505: inst = 32'h8220000;
      15506: inst = 32'h10408000;
      15507: inst = 32'hc405098;
      15508: inst = 32'h8220000;
      15509: inst = 32'h10408000;
      15510: inst = 32'hc405099;
      15511: inst = 32'h8220000;
      15512: inst = 32'h10408000;
      15513: inst = 32'hc40509d;
      15514: inst = 32'h8220000;
      15515: inst = 32'h10408000;
      15516: inst = 32'hc40509e;
      15517: inst = 32'h8220000;
      15518: inst = 32'h10408000;
      15519: inst = 32'hc40509f;
      15520: inst = 32'h8220000;
      15521: inst = 32'h10408000;
      15522: inst = 32'hc4050a0;
      15523: inst = 32'h8220000;
      15524: inst = 32'h10408000;
      15525: inst = 32'hc4050df;
      15526: inst = 32'h8220000;
      15527: inst = 32'h10408000;
      15528: inst = 32'hc4050e0;
      15529: inst = 32'h8220000;
      15530: inst = 32'h10408000;
      15531: inst = 32'hc4050e1;
      15532: inst = 32'h8220000;
      15533: inst = 32'h10408000;
      15534: inst = 32'hc4050e2;
      15535: inst = 32'h8220000;
      15536: inst = 32'h10408000;
      15537: inst = 32'hc4050e6;
      15538: inst = 32'h8220000;
      15539: inst = 32'h10408000;
      15540: inst = 32'hc4050e7;
      15541: inst = 32'h8220000;
      15542: inst = 32'h10408000;
      15543: inst = 32'hc4050f8;
      15544: inst = 32'h8220000;
      15545: inst = 32'h10408000;
      15546: inst = 32'hc4050f9;
      15547: inst = 32'h8220000;
      15548: inst = 32'h10408000;
      15549: inst = 32'hc4050fd;
      15550: inst = 32'h8220000;
      15551: inst = 32'h10408000;
      15552: inst = 32'hc4050fe;
      15553: inst = 32'h8220000;
      15554: inst = 32'h10408000;
      15555: inst = 32'hc4050ff;
      15556: inst = 32'h8220000;
      15557: inst = 32'h10408000;
      15558: inst = 32'hc405100;
      15559: inst = 32'h8220000;
      15560: inst = 32'h10408000;
      15561: inst = 32'hc40513f;
      15562: inst = 32'h8220000;
      15563: inst = 32'h10408000;
      15564: inst = 32'hc405140;
      15565: inst = 32'h8220000;
      15566: inst = 32'h10408000;
      15567: inst = 32'hc405141;
      15568: inst = 32'h8220000;
      15569: inst = 32'h10408000;
      15570: inst = 32'hc405146;
      15571: inst = 32'h8220000;
      15572: inst = 32'h10408000;
      15573: inst = 32'hc405147;
      15574: inst = 32'h8220000;
      15575: inst = 32'h10408000;
      15576: inst = 32'hc405158;
      15577: inst = 32'h8220000;
      15578: inst = 32'h10408000;
      15579: inst = 32'hc405159;
      15580: inst = 32'h8220000;
      15581: inst = 32'h10408000;
      15582: inst = 32'hc40515e;
      15583: inst = 32'h8220000;
      15584: inst = 32'h10408000;
      15585: inst = 32'hc40515f;
      15586: inst = 32'h8220000;
      15587: inst = 32'h10408000;
      15588: inst = 32'hc405160;
      15589: inst = 32'h8220000;
      15590: inst = 32'h10408000;
      15591: inst = 32'hc40519f;
      15592: inst = 32'h8220000;
      15593: inst = 32'h10408000;
      15594: inst = 32'hc4051a0;
      15595: inst = 32'h8220000;
      15596: inst = 32'h10408000;
      15597: inst = 32'hc4051a6;
      15598: inst = 32'h8220000;
      15599: inst = 32'h10408000;
      15600: inst = 32'hc4051a7;
      15601: inst = 32'h8220000;
      15602: inst = 32'h10408000;
      15603: inst = 32'hc4051b8;
      15604: inst = 32'h8220000;
      15605: inst = 32'h10408000;
      15606: inst = 32'hc4051b9;
      15607: inst = 32'h8220000;
      15608: inst = 32'h10408000;
      15609: inst = 32'hc4051bf;
      15610: inst = 32'h8220000;
      15611: inst = 32'h10408000;
      15612: inst = 32'hc4051c0;
      15613: inst = 32'h8220000;
      15614: inst = 32'h10408000;
      15615: inst = 32'hc4051ff;
      15616: inst = 32'h8220000;
      15617: inst = 32'h10408000;
      15618: inst = 32'hc405200;
      15619: inst = 32'h8220000;
      15620: inst = 32'h10408000;
      15621: inst = 32'hc405206;
      15622: inst = 32'h8220000;
      15623: inst = 32'h10408000;
      15624: inst = 32'hc405207;
      15625: inst = 32'h8220000;
      15626: inst = 32'h10408000;
      15627: inst = 32'hc405218;
      15628: inst = 32'h8220000;
      15629: inst = 32'h10408000;
      15630: inst = 32'hc405219;
      15631: inst = 32'h8220000;
      15632: inst = 32'h10408000;
      15633: inst = 32'hc40521f;
      15634: inst = 32'h8220000;
      15635: inst = 32'h10408000;
      15636: inst = 32'hc405220;
      15637: inst = 32'h8220000;
      15638: inst = 32'h10408000;
      15639: inst = 32'hc40525f;
      15640: inst = 32'h8220000;
      15641: inst = 32'h10408000;
      15642: inst = 32'hc405260;
      15643: inst = 32'h8220000;
      15644: inst = 32'h10408000;
      15645: inst = 32'hc405266;
      15646: inst = 32'h8220000;
      15647: inst = 32'h10408000;
      15648: inst = 32'hc405267;
      15649: inst = 32'h8220000;
      15650: inst = 32'h10408000;
      15651: inst = 32'hc405278;
      15652: inst = 32'h8220000;
      15653: inst = 32'h10408000;
      15654: inst = 32'hc405279;
      15655: inst = 32'h8220000;
      15656: inst = 32'h10408000;
      15657: inst = 32'hc40527f;
      15658: inst = 32'h8220000;
      15659: inst = 32'h10408000;
      15660: inst = 32'hc405280;
      15661: inst = 32'h8220000;
      15662: inst = 32'h10408000;
      15663: inst = 32'hc4052bf;
      15664: inst = 32'h8220000;
      15665: inst = 32'h10408000;
      15666: inst = 32'hc4052c0;
      15667: inst = 32'h8220000;
      15668: inst = 32'h10408000;
      15669: inst = 32'hc4052c6;
      15670: inst = 32'h8220000;
      15671: inst = 32'h10408000;
      15672: inst = 32'hc4052c7;
      15673: inst = 32'h8220000;
      15674: inst = 32'h10408000;
      15675: inst = 32'hc4052d8;
      15676: inst = 32'h8220000;
      15677: inst = 32'h10408000;
      15678: inst = 32'hc4052d9;
      15679: inst = 32'h8220000;
      15680: inst = 32'h10408000;
      15681: inst = 32'hc4052df;
      15682: inst = 32'h8220000;
      15683: inst = 32'h10408000;
      15684: inst = 32'hc4052e0;
      15685: inst = 32'h8220000;
      15686: inst = 32'hc207bae;
      15687: inst = 32'h10408000;
      15688: inst = 32'hc404ea5;
      15689: inst = 32'h8220000;
      15690: inst = 32'h10408000;
      15691: inst = 32'hc404eba;
      15692: inst = 32'h8220000;
      15693: inst = 32'hc20c5b4;
      15694: inst = 32'h10408000;
      15695: inst = 32'hc404ea6;
      15696: inst = 32'h8220000;
      15697: inst = 32'h10408000;
      15698: inst = 32'hc404eb9;
      15699: inst = 32'h8220000;
      15700: inst = 32'hc20d5f4;
      15701: inst = 32'h10408000;
      15702: inst = 32'hc404ea7;
      15703: inst = 32'h8220000;
      15704: inst = 32'h10408000;
      15705: inst = 32'hc404eb8;
      15706: inst = 32'h8220000;
      15707: inst = 32'hc20a4b1;
      15708: inst = 32'h10408000;
      15709: inst = 32'hc404eff;
      15710: inst = 32'h8220000;
      15711: inst = 32'h10408000;
      15712: inst = 32'hc404f20;
      15713: inst = 32'h8220000;
      15714: inst = 32'h10408000;
      15715: inst = 32'hc404fbf;
      15716: inst = 32'h8220000;
      15717: inst = 32'h10408000;
      15718: inst = 32'hc404fe0;
      15719: inst = 32'h8220000;
      15720: inst = 32'hc2062ed;
      15721: inst = 32'h10408000;
      15722: inst = 32'hc404f06;
      15723: inst = 32'h8220000;
      15724: inst = 32'h10408000;
      15725: inst = 32'hc404f19;
      15726: inst = 32'h8220000;
      15727: inst = 32'hc209450;
      15728: inst = 32'h10408000;
      15729: inst = 32'hc404f07;
      15730: inst = 32'h8220000;
      15731: inst = 32'h10408000;
      15732: inst = 32'hc404f18;
      15733: inst = 32'h8220000;
      15734: inst = 32'h10408000;
      15735: inst = 32'hc405209;
      15736: inst = 32'h8220000;
      15737: inst = 32'h10408000;
      15738: inst = 32'hc405216;
      15739: inst = 32'h8220000;
      15740: inst = 32'hc20a4d1;
      15741: inst = 32'h10408000;
      15742: inst = 32'hc404f5f;
      15743: inst = 32'h8220000;
      15744: inst = 32'h10408000;
      15745: inst = 32'hc404f80;
      15746: inst = 32'h8220000;
      15747: inst = 32'hc204a49;
      15748: inst = 32'h10408000;
      15749: inst = 32'hc404fa8;
      15750: inst = 32'h8220000;
      15751: inst = 32'h10408000;
      15752: inst = 32'hc404fac;
      15753: inst = 32'h8220000;
      15754: inst = 32'h10408000;
      15755: inst = 32'hc405008;
      15756: inst = 32'h8220000;
      15757: inst = 32'h10408000;
      15758: inst = 32'hc40500c;
      15759: inst = 32'h8220000;
      15760: inst = 32'hc205acb;
      15761: inst = 32'h10408000;
      15762: inst = 32'hc404fc5;
      15763: inst = 32'h8220000;
      15764: inst = 32'h10408000;
      15765: inst = 32'hc404fda;
      15766: inst = 32'h8220000;
      15767: inst = 32'h10408000;
      15768: inst = 32'hc405336;
      15769: inst = 32'h8220000;
      15770: inst = 32'h10408000;
      15771: inst = 32'hc405380;
      15772: inst = 32'h8220000;
      15773: inst = 32'h10408000;
      15774: inst = 32'hc40539f;
      15775: inst = 32'h8220000;
      15776: inst = 32'h10408000;
      15777: inst = 32'hc4053dd;
      15778: inst = 32'h8220000;
      15779: inst = 32'h10408000;
      15780: inst = 32'hc405402;
      15781: inst = 32'h8220000;
      15782: inst = 32'hc20630d;
      15783: inst = 32'h10408000;
      15784: inst = 32'hc40501f;
      15785: inst = 32'h8220000;
      15786: inst = 32'h10408000;
      15787: inst = 32'hc405040;
      15788: inst = 32'h8220000;
      15789: inst = 32'hc205aec;
      15790: inst = 32'h10408000;
      15791: inst = 32'hc405024;
      15792: inst = 32'h8220000;
      15793: inst = 32'h10408000;
      15794: inst = 32'hc40503b;
      15795: inst = 32'h8220000;
      15796: inst = 32'h10408000;
      15797: inst = 32'hc405083;
      15798: inst = 32'h8220000;
      15799: inst = 32'h10408000;
      15800: inst = 32'hc40509c;
      15801: inst = 32'h8220000;
      15802: inst = 32'h10408000;
      15803: inst = 32'hc4051a1;
      15804: inst = 32'h8220000;
      15805: inst = 32'h10408000;
      15806: inst = 32'hc4051be;
      15807: inst = 32'h8220000;
      15808: inst = 32'h10408000;
      15809: inst = 32'hc405329;
      15810: inst = 32'h8220000;
      15811: inst = 32'h10408000;
      15812: inst = 32'hc405568;
      15813: inst = 32'h8220000;
      15814: inst = 32'h10408000;
      15815: inst = 32'hc405577;
      15816: inst = 32'h8220000;
      15817: inst = 32'h10408000;
      15818: inst = 32'hc4057a7;
      15819: inst = 32'h8220000;
      15820: inst = 32'h10408000;
      15821: inst = 32'hc4057b8;
      15822: inst = 32'h8220000;
      15823: inst = 32'hc205269;
      15824: inst = 32'h10408000;
      15825: inst = 32'hc405025;
      15826: inst = 32'h8220000;
      15827: inst = 32'h10408000;
      15828: inst = 32'hc40503a;
      15829: inst = 32'h8220000;
      15830: inst = 32'h10408000;
      15831: inst = 32'hc40537e;
      15832: inst = 32'h8220000;
      15833: inst = 32'h10408000;
      15834: inst = 32'hc4053a1;
      15835: inst = 32'h8220000;
      15836: inst = 32'h10408000;
      15837: inst = 32'hc40549c;
      15838: inst = 32'h8220000;
      15839: inst = 32'h10408000;
      15840: inst = 32'hc4054c3;
      15841: inst = 32'h8220000;
      15842: inst = 32'hc20528a;
      15843: inst = 32'h10408000;
      15844: inst = 32'hc405084;
      15845: inst = 32'h8220000;
      15846: inst = 32'h10408000;
      15847: inst = 32'hc40509b;
      15848: inst = 32'h8220000;
      15849: inst = 32'h10408000;
      15850: inst = 32'hc4050e3;
      15851: inst = 32'h8220000;
      15852: inst = 32'h10408000;
      15853: inst = 32'hc4050fc;
      15854: inst = 32'h8220000;
      15855: inst = 32'h10408000;
      15856: inst = 32'hc4052c5;
      15857: inst = 32'h8220000;
      15858: inst = 32'h10408000;
      15859: inst = 32'hc4052da;
      15860: inst = 32'h8220000;
      15861: inst = 32'h10408000;
      15862: inst = 32'hc4053e9;
      15863: inst = 32'h8220000;
      15864: inst = 32'h10408000;
      15865: inst = 32'hc4053f6;
      15866: inst = 32'h8220000;
      15867: inst = 32'h10408000;
      15868: inst = 32'hc405449;
      15869: inst = 32'h8220000;
      15870: inst = 32'h10408000;
      15871: inst = 32'hc405456;
      15872: inst = 32'h8220000;
      15873: inst = 32'h10408000;
      15874: inst = 32'hc4054a9;
      15875: inst = 32'h8220000;
      15876: inst = 32'h10408000;
      15877: inst = 32'hc4054b6;
      15878: inst = 32'h8220000;
      15879: inst = 32'h10408000;
      15880: inst = 32'hc405509;
      15881: inst = 32'h8220000;
      15882: inst = 32'h10408000;
      15883: inst = 32'hc405516;
      15884: inst = 32'h8220000;
      15885: inst = 32'h10408000;
      15886: inst = 32'hc40555e;
      15887: inst = 32'h8220000;
      15888: inst = 32'h10408000;
      15889: inst = 32'hc405569;
      15890: inst = 32'h8220000;
      15891: inst = 32'h10408000;
      15892: inst = 32'hc405576;
      15893: inst = 32'h8220000;
      15894: inst = 32'h10408000;
      15895: inst = 32'hc405581;
      15896: inst = 32'h8220000;
      15897: inst = 32'h10408000;
      15898: inst = 32'hc4055c9;
      15899: inst = 32'h8220000;
      15900: inst = 32'h10408000;
      15901: inst = 32'hc4055d6;
      15902: inst = 32'h8220000;
      15903: inst = 32'h10408000;
      15904: inst = 32'hc405628;
      15905: inst = 32'h8220000;
      15906: inst = 32'h10408000;
      15907: inst = 32'hc405629;
      15908: inst = 32'h8220000;
      15909: inst = 32'h10408000;
      15910: inst = 32'hc405636;
      15911: inst = 32'h8220000;
      15912: inst = 32'h10408000;
      15913: inst = 32'hc405637;
      15914: inst = 32'h8220000;
      15915: inst = 32'h10408000;
      15916: inst = 32'hc40567d;
      15917: inst = 32'h8220000;
      15918: inst = 32'h10408000;
      15919: inst = 32'hc405688;
      15920: inst = 32'h8220000;
      15921: inst = 32'h10408000;
      15922: inst = 32'hc405689;
      15923: inst = 32'h8220000;
      15924: inst = 32'h10408000;
      15925: inst = 32'hc405696;
      15926: inst = 32'h8220000;
      15927: inst = 32'h10408000;
      15928: inst = 32'hc405697;
      15929: inst = 32'h8220000;
      15930: inst = 32'h10408000;
      15931: inst = 32'hc4056a2;
      15932: inst = 32'h8220000;
      15933: inst = 32'h10408000;
      15934: inst = 32'hc4056e8;
      15935: inst = 32'h8220000;
      15936: inst = 32'h10408000;
      15937: inst = 32'hc4056e9;
      15938: inst = 32'h8220000;
      15939: inst = 32'h10408000;
      15940: inst = 32'hc4056f6;
      15941: inst = 32'h8220000;
      15942: inst = 32'h10408000;
      15943: inst = 32'hc4056f7;
      15944: inst = 32'h8220000;
      15945: inst = 32'h10408000;
      15946: inst = 32'hc405748;
      15947: inst = 32'h8220000;
      15948: inst = 32'h10408000;
      15949: inst = 32'hc405749;
      15950: inst = 32'h8220000;
      15951: inst = 32'h10408000;
      15952: inst = 32'hc405756;
      15953: inst = 32'h8220000;
      15954: inst = 32'h10408000;
      15955: inst = 32'hc405757;
      15956: inst = 32'h8220000;
      15957: inst = 32'h10408000;
      15958: inst = 32'hc4057a8;
      15959: inst = 32'h8220000;
      15960: inst = 32'h10408000;
      15961: inst = 32'hc4057a9;
      15962: inst = 32'h8220000;
      15963: inst = 32'h10408000;
      15964: inst = 32'hc4057b6;
      15965: inst = 32'h8220000;
      15966: inst = 32'h10408000;
      15967: inst = 32'hc4057b7;
      15968: inst = 32'h8220000;
      15969: inst = 32'hc205aab;
      15970: inst = 32'h10408000;
      15971: inst = 32'hc405142;
      15972: inst = 32'h8220000;
      15973: inst = 32'h10408000;
      15974: inst = 32'hc40515d;
      15975: inst = 32'h8220000;
      15976: inst = 32'hc20cdd4;
      15977: inst = 32'h10408000;
      15978: inst = 32'hc40519e;
      15979: inst = 32'h8220000;
      15980: inst = 32'h10408000;
      15981: inst = 32'hc4051c1;
      15982: inst = 32'h8220000;
      15983: inst = 32'hc209471;
      15984: inst = 32'h10408000;
      15985: inst = 32'hc4051b6;
      15986: inst = 32'h8220000;
      15987: inst = 32'hc20de55;
      15988: inst = 32'h10408000;
      15989: inst = 32'hc4051fd;
      15990: inst = 32'h8220000;
      15991: inst = 32'h10408000;
      15992: inst = 32'hc405222;
      15993: inst = 32'h8220000;
      15994: inst = 32'hc209492;
      15995: inst = 32'h10408000;
      15996: inst = 32'hc4051fe;
      15997: inst = 32'h8220000;
      15998: inst = 32'h10408000;
      15999: inst = 32'hc405221;
      16000: inst = 32'h8220000;
      16001: inst = 32'hc205acc;
      16002: inst = 32'h10408000;
      16003: inst = 32'hc405201;
      16004: inst = 32'h8220000;
      16005: inst = 32'h10408000;
      16006: inst = 32'hc40521e;
      16007: inst = 32'h8220000;
      16008: inst = 32'h10408000;
      16009: inst = 32'hc405261;
      16010: inst = 32'h8220000;
      16011: inst = 32'h10408000;
      16012: inst = 32'hc40527e;
      16013: inst = 32'h8220000;
      16014: inst = 32'h10408000;
      16015: inst = 32'hc4052c1;
      16016: inst = 32'h8220000;
      16017: inst = 32'h10408000;
      16018: inst = 32'hc4052de;
      16019: inst = 32'h8220000;
      16020: inst = 32'hc20e696;
      16021: inst = 32'h10408000;
      16022: inst = 32'hc40525c;
      16023: inst = 32'h8220000;
      16024: inst = 32'h10408000;
      16025: inst = 32'hc405283;
      16026: inst = 32'h8220000;
      16027: inst = 32'hc209cb2;
      16028: inst = 32'h10408000;
      16029: inst = 32'hc40525d;
      16030: inst = 32'h8220000;
      16031: inst = 32'h10408000;
      16032: inst = 32'hc405282;
      16033: inst = 32'h8220000;
      16034: inst = 32'hc208c2f;
      16035: inst = 32'h10408000;
      16036: inst = 32'hc405269;
      16037: inst = 32'h8220000;
      16038: inst = 32'h10408000;
      16039: inst = 32'hc405276;
      16040: inst = 32'h8220000;
      16041: inst = 32'hc20ad33;
      16042: inst = 32'h10408000;
      16043: inst = 32'hc4052bc;
      16044: inst = 32'h8220000;
      16045: inst = 32'h10408000;
      16046: inst = 32'hc4052e3;
      16047: inst = 32'h8220000;
      16048: inst = 32'hc2083ee;
      16049: inst = 32'h10408000;
      16050: inst = 32'hc4052c9;
      16051: inst = 32'h8220000;
      16052: inst = 32'h10408000;
      16053: inst = 32'hc4052d6;
      16054: inst = 32'h8220000;
      16055: inst = 32'hc206b50;
      16056: inst = 32'h10408000;
      16057: inst = 32'hc405300;
      16058: inst = 32'h8220000;
      16059: inst = 32'h10408000;
      16060: inst = 32'hc405301;
      16061: inst = 32'h8220000;
      16062: inst = 32'h10408000;
      16063: inst = 32'hc405302;
      16064: inst = 32'h8220000;
      16065: inst = 32'h10408000;
      16066: inst = 32'hc405303;
      16067: inst = 32'h8220000;
      16068: inst = 32'h10408000;
      16069: inst = 32'hc405304;
      16070: inst = 32'h8220000;
      16071: inst = 32'h10408000;
      16072: inst = 32'hc405305;
      16073: inst = 32'h8220000;
      16074: inst = 32'h10408000;
      16075: inst = 32'hc405306;
      16076: inst = 32'h8220000;
      16077: inst = 32'h10408000;
      16078: inst = 32'hc405307;
      16079: inst = 32'h8220000;
      16080: inst = 32'h10408000;
      16081: inst = 32'hc405308;
      16082: inst = 32'h8220000;
      16083: inst = 32'h10408000;
      16084: inst = 32'hc405309;
      16085: inst = 32'h8220000;
      16086: inst = 32'h10408000;
      16087: inst = 32'hc40530a;
      16088: inst = 32'h8220000;
      16089: inst = 32'h10408000;
      16090: inst = 32'hc40530b;
      16091: inst = 32'h8220000;
      16092: inst = 32'h10408000;
      16093: inst = 32'hc40530c;
      16094: inst = 32'h8220000;
      16095: inst = 32'h10408000;
      16096: inst = 32'hc40530d;
      16097: inst = 32'h8220000;
      16098: inst = 32'h10408000;
      16099: inst = 32'hc40530e;
      16100: inst = 32'h8220000;
      16101: inst = 32'h10408000;
      16102: inst = 32'hc40530f;
      16103: inst = 32'h8220000;
      16104: inst = 32'h10408000;
      16105: inst = 32'hc405310;
      16106: inst = 32'h8220000;
      16107: inst = 32'h10408000;
      16108: inst = 32'hc405311;
      16109: inst = 32'h8220000;
      16110: inst = 32'h10408000;
      16111: inst = 32'hc405312;
      16112: inst = 32'h8220000;
      16113: inst = 32'h10408000;
      16114: inst = 32'hc405313;
      16115: inst = 32'h8220000;
      16116: inst = 32'h10408000;
      16117: inst = 32'hc405314;
      16118: inst = 32'h8220000;
      16119: inst = 32'h10408000;
      16120: inst = 32'hc405315;
      16121: inst = 32'h8220000;
      16122: inst = 32'h10408000;
      16123: inst = 32'hc405316;
      16124: inst = 32'h8220000;
      16125: inst = 32'h10408000;
      16126: inst = 32'hc405317;
      16127: inst = 32'h8220000;
      16128: inst = 32'h10408000;
      16129: inst = 32'hc405318;
      16130: inst = 32'h8220000;
      16131: inst = 32'h10408000;
      16132: inst = 32'hc405319;
      16133: inst = 32'h8220000;
      16134: inst = 32'h10408000;
      16135: inst = 32'hc40531a;
      16136: inst = 32'h8220000;
      16137: inst = 32'h10408000;
      16138: inst = 32'hc40532a;
      16139: inst = 32'h8220000;
      16140: inst = 32'h10408000;
      16141: inst = 32'hc40532b;
      16142: inst = 32'h8220000;
      16143: inst = 32'h10408000;
      16144: inst = 32'hc40532c;
      16145: inst = 32'h8220000;
      16146: inst = 32'h10408000;
      16147: inst = 32'hc40532d;
      16148: inst = 32'h8220000;
      16149: inst = 32'h10408000;
      16150: inst = 32'hc40532e;
      16151: inst = 32'h8220000;
      16152: inst = 32'h10408000;
      16153: inst = 32'hc40532f;
      16154: inst = 32'h8220000;
      16155: inst = 32'h10408000;
      16156: inst = 32'hc405330;
      16157: inst = 32'h8220000;
      16158: inst = 32'h10408000;
      16159: inst = 32'hc405331;
      16160: inst = 32'h8220000;
      16161: inst = 32'h10408000;
      16162: inst = 32'hc405332;
      16163: inst = 32'h8220000;
      16164: inst = 32'h10408000;
      16165: inst = 32'hc405333;
      16166: inst = 32'h8220000;
      16167: inst = 32'h10408000;
      16168: inst = 32'hc405334;
      16169: inst = 32'h8220000;
      16170: inst = 32'h10408000;
      16171: inst = 32'hc405335;
      16172: inst = 32'h8220000;
      16173: inst = 32'h10408000;
      16174: inst = 32'hc405345;
      16175: inst = 32'h8220000;
      16176: inst = 32'h10408000;
      16177: inst = 32'hc405346;
      16178: inst = 32'h8220000;
      16179: inst = 32'h10408000;
      16180: inst = 32'hc405347;
      16181: inst = 32'h8220000;
      16182: inst = 32'h10408000;
      16183: inst = 32'hc405348;
      16184: inst = 32'h8220000;
      16185: inst = 32'h10408000;
      16186: inst = 32'hc405349;
      16187: inst = 32'h8220000;
      16188: inst = 32'h10408000;
      16189: inst = 32'hc40534a;
      16190: inst = 32'h8220000;
      16191: inst = 32'h10408000;
      16192: inst = 32'hc40534b;
      16193: inst = 32'h8220000;
      16194: inst = 32'h10408000;
      16195: inst = 32'hc40534c;
      16196: inst = 32'h8220000;
      16197: inst = 32'h10408000;
      16198: inst = 32'hc40534d;
      16199: inst = 32'h8220000;
      16200: inst = 32'h10408000;
      16201: inst = 32'hc40534e;
      16202: inst = 32'h8220000;
      16203: inst = 32'h10408000;
      16204: inst = 32'hc40534f;
      16205: inst = 32'h8220000;
      16206: inst = 32'h10408000;
      16207: inst = 32'hc405350;
      16208: inst = 32'h8220000;
      16209: inst = 32'h10408000;
      16210: inst = 32'hc405351;
      16211: inst = 32'h8220000;
      16212: inst = 32'h10408000;
      16213: inst = 32'hc405352;
      16214: inst = 32'h8220000;
      16215: inst = 32'h10408000;
      16216: inst = 32'hc405353;
      16217: inst = 32'h8220000;
      16218: inst = 32'h10408000;
      16219: inst = 32'hc405354;
      16220: inst = 32'h8220000;
      16221: inst = 32'h10408000;
      16222: inst = 32'hc405355;
      16223: inst = 32'h8220000;
      16224: inst = 32'h10408000;
      16225: inst = 32'hc405356;
      16226: inst = 32'h8220000;
      16227: inst = 32'h10408000;
      16228: inst = 32'hc405357;
      16229: inst = 32'h8220000;
      16230: inst = 32'h10408000;
      16231: inst = 32'hc405358;
      16232: inst = 32'h8220000;
      16233: inst = 32'h10408000;
      16234: inst = 32'hc405359;
      16235: inst = 32'h8220000;
      16236: inst = 32'h10408000;
      16237: inst = 32'hc40535a;
      16238: inst = 32'h8220000;
      16239: inst = 32'h10408000;
      16240: inst = 32'hc40535b;
      16241: inst = 32'h8220000;
      16242: inst = 32'h10408000;
      16243: inst = 32'hc40535c;
      16244: inst = 32'h8220000;
      16245: inst = 32'h10408000;
      16246: inst = 32'hc40535d;
      16247: inst = 32'h8220000;
      16248: inst = 32'h10408000;
      16249: inst = 32'hc40535e;
      16250: inst = 32'h8220000;
      16251: inst = 32'h10408000;
      16252: inst = 32'hc40535f;
      16253: inst = 32'h8220000;
      16254: inst = 32'h10408000;
      16255: inst = 32'hc405360;
      16256: inst = 32'h8220000;
      16257: inst = 32'h10408000;
      16258: inst = 32'hc405361;
      16259: inst = 32'h8220000;
      16260: inst = 32'h10408000;
      16261: inst = 32'hc405362;
      16262: inst = 32'h8220000;
      16263: inst = 32'h10408000;
      16264: inst = 32'hc405363;
      16265: inst = 32'h8220000;
      16266: inst = 32'h10408000;
      16267: inst = 32'hc405364;
      16268: inst = 32'h8220000;
      16269: inst = 32'h10408000;
      16270: inst = 32'hc405365;
      16271: inst = 32'h8220000;
      16272: inst = 32'h10408000;
      16273: inst = 32'hc405366;
      16274: inst = 32'h8220000;
      16275: inst = 32'h10408000;
      16276: inst = 32'hc405367;
      16277: inst = 32'h8220000;
      16278: inst = 32'h10408000;
      16279: inst = 32'hc405368;
      16280: inst = 32'h8220000;
      16281: inst = 32'h10408000;
      16282: inst = 32'hc405369;
      16283: inst = 32'h8220000;
      16284: inst = 32'h10408000;
      16285: inst = 32'hc40536a;
      16286: inst = 32'h8220000;
      16287: inst = 32'h10408000;
      16288: inst = 32'hc40536b;
      16289: inst = 32'h8220000;
      16290: inst = 32'h10408000;
      16291: inst = 32'hc40536c;
      16292: inst = 32'h8220000;
      16293: inst = 32'h10408000;
      16294: inst = 32'hc40536d;
      16295: inst = 32'h8220000;
      16296: inst = 32'h10408000;
      16297: inst = 32'hc40536e;
      16298: inst = 32'h8220000;
      16299: inst = 32'h10408000;
      16300: inst = 32'hc40536f;
      16301: inst = 32'h8220000;
      16302: inst = 32'h10408000;
      16303: inst = 32'hc405370;
      16304: inst = 32'h8220000;
      16305: inst = 32'h10408000;
      16306: inst = 32'hc405371;
      16307: inst = 32'h8220000;
      16308: inst = 32'h10408000;
      16309: inst = 32'hc405372;
      16310: inst = 32'h8220000;
      16311: inst = 32'h10408000;
      16312: inst = 32'hc405373;
      16313: inst = 32'h8220000;
      16314: inst = 32'h10408000;
      16315: inst = 32'hc405374;
      16316: inst = 32'h8220000;
      16317: inst = 32'h10408000;
      16318: inst = 32'hc405375;
      16319: inst = 32'h8220000;
      16320: inst = 32'h10408000;
      16321: inst = 32'hc405376;
      16322: inst = 32'h8220000;
      16323: inst = 32'h10408000;
      16324: inst = 32'hc405377;
      16325: inst = 32'h8220000;
      16326: inst = 32'h10408000;
      16327: inst = 32'hc405378;
      16328: inst = 32'h8220000;
      16329: inst = 32'h10408000;
      16330: inst = 32'hc405379;
      16331: inst = 32'h8220000;
      16332: inst = 32'h10408000;
      16333: inst = 32'hc40538a;
      16334: inst = 32'h8220000;
      16335: inst = 32'h10408000;
      16336: inst = 32'hc40538b;
      16337: inst = 32'h8220000;
      16338: inst = 32'h10408000;
      16339: inst = 32'hc40538c;
      16340: inst = 32'h8220000;
      16341: inst = 32'h10408000;
      16342: inst = 32'hc40538d;
      16343: inst = 32'h8220000;
      16344: inst = 32'h10408000;
      16345: inst = 32'hc40538e;
      16346: inst = 32'h8220000;
      16347: inst = 32'h10408000;
      16348: inst = 32'hc40538f;
      16349: inst = 32'h8220000;
      16350: inst = 32'h10408000;
      16351: inst = 32'hc405390;
      16352: inst = 32'h8220000;
      16353: inst = 32'h10408000;
      16354: inst = 32'hc405391;
      16355: inst = 32'h8220000;
      16356: inst = 32'h10408000;
      16357: inst = 32'hc405392;
      16358: inst = 32'h8220000;
      16359: inst = 32'h10408000;
      16360: inst = 32'hc405393;
      16361: inst = 32'h8220000;
      16362: inst = 32'h10408000;
      16363: inst = 32'hc405394;
      16364: inst = 32'h8220000;
      16365: inst = 32'h10408000;
      16366: inst = 32'hc405395;
      16367: inst = 32'h8220000;
      16368: inst = 32'h10408000;
      16369: inst = 32'hc4053a6;
      16370: inst = 32'h8220000;
      16371: inst = 32'h10408000;
      16372: inst = 32'hc4053a7;
      16373: inst = 32'h8220000;
      16374: inst = 32'h10408000;
      16375: inst = 32'hc4053a8;
      16376: inst = 32'h8220000;
      16377: inst = 32'h10408000;
      16378: inst = 32'hc4053a9;
      16379: inst = 32'h8220000;
      16380: inst = 32'h10408000;
      16381: inst = 32'hc4053aa;
      16382: inst = 32'h8220000;
      16383: inst = 32'h10408000;
      16384: inst = 32'hc4053ab;
      16385: inst = 32'h8220000;
      16386: inst = 32'h10408000;
      16387: inst = 32'hc4053ac;
      16388: inst = 32'h8220000;
      16389: inst = 32'h10408000;
      16390: inst = 32'hc4053ad;
      16391: inst = 32'h8220000;
      16392: inst = 32'h10408000;
      16393: inst = 32'hc4053ae;
      16394: inst = 32'h8220000;
      16395: inst = 32'h10408000;
      16396: inst = 32'hc4053af;
      16397: inst = 32'h8220000;
      16398: inst = 32'h10408000;
      16399: inst = 32'hc4053b0;
      16400: inst = 32'h8220000;
      16401: inst = 32'h10408000;
      16402: inst = 32'hc4053b1;
      16403: inst = 32'h8220000;
      16404: inst = 32'h10408000;
      16405: inst = 32'hc4053b2;
      16406: inst = 32'h8220000;
      16407: inst = 32'h10408000;
      16408: inst = 32'hc4053b3;
      16409: inst = 32'h8220000;
      16410: inst = 32'h10408000;
      16411: inst = 32'hc4053b4;
      16412: inst = 32'h8220000;
      16413: inst = 32'h10408000;
      16414: inst = 32'hc4053b5;
      16415: inst = 32'h8220000;
      16416: inst = 32'h10408000;
      16417: inst = 32'hc4053b6;
      16418: inst = 32'h8220000;
      16419: inst = 32'h10408000;
      16420: inst = 32'hc4053b7;
      16421: inst = 32'h8220000;
      16422: inst = 32'h10408000;
      16423: inst = 32'hc4053b8;
      16424: inst = 32'h8220000;
      16425: inst = 32'h10408000;
      16426: inst = 32'hc4053b9;
      16427: inst = 32'h8220000;
      16428: inst = 32'h10408000;
      16429: inst = 32'hc4053ba;
      16430: inst = 32'h8220000;
      16431: inst = 32'h10408000;
      16432: inst = 32'hc4053bb;
      16433: inst = 32'h8220000;
      16434: inst = 32'h10408000;
      16435: inst = 32'hc4053bc;
      16436: inst = 32'h8220000;
      16437: inst = 32'h10408000;
      16438: inst = 32'hc4053bd;
      16439: inst = 32'h8220000;
      16440: inst = 32'h10408000;
      16441: inst = 32'hc4053be;
      16442: inst = 32'h8220000;
      16443: inst = 32'h10408000;
      16444: inst = 32'hc4053bf;
      16445: inst = 32'h8220000;
      16446: inst = 32'h10408000;
      16447: inst = 32'hc4053c0;
      16448: inst = 32'h8220000;
      16449: inst = 32'h10408000;
      16450: inst = 32'hc4053c1;
      16451: inst = 32'h8220000;
      16452: inst = 32'h10408000;
      16453: inst = 32'hc4053c2;
      16454: inst = 32'h8220000;
      16455: inst = 32'h10408000;
      16456: inst = 32'hc4053c3;
      16457: inst = 32'h8220000;
      16458: inst = 32'h10408000;
      16459: inst = 32'hc4053c4;
      16460: inst = 32'h8220000;
      16461: inst = 32'h10408000;
      16462: inst = 32'hc4053c5;
      16463: inst = 32'h8220000;
      16464: inst = 32'h10408000;
      16465: inst = 32'hc4053c6;
      16466: inst = 32'h8220000;
      16467: inst = 32'h10408000;
      16468: inst = 32'hc4053c7;
      16469: inst = 32'h8220000;
      16470: inst = 32'h10408000;
      16471: inst = 32'hc4053c8;
      16472: inst = 32'h8220000;
      16473: inst = 32'h10408000;
      16474: inst = 32'hc4053c9;
      16475: inst = 32'h8220000;
      16476: inst = 32'h10408000;
      16477: inst = 32'hc4053ca;
      16478: inst = 32'h8220000;
      16479: inst = 32'h10408000;
      16480: inst = 32'hc4053cb;
      16481: inst = 32'h8220000;
      16482: inst = 32'h10408000;
      16483: inst = 32'hc4053cc;
      16484: inst = 32'h8220000;
      16485: inst = 32'h10408000;
      16486: inst = 32'hc4053cd;
      16487: inst = 32'h8220000;
      16488: inst = 32'h10408000;
      16489: inst = 32'hc4053ce;
      16490: inst = 32'h8220000;
      16491: inst = 32'h10408000;
      16492: inst = 32'hc4053cf;
      16493: inst = 32'h8220000;
      16494: inst = 32'h10408000;
      16495: inst = 32'hc4053d0;
      16496: inst = 32'h8220000;
      16497: inst = 32'h10408000;
      16498: inst = 32'hc4053d1;
      16499: inst = 32'h8220000;
      16500: inst = 32'h10408000;
      16501: inst = 32'hc4053d2;
      16502: inst = 32'h8220000;
      16503: inst = 32'h10408000;
      16504: inst = 32'hc4053d3;
      16505: inst = 32'h8220000;
      16506: inst = 32'h10408000;
      16507: inst = 32'hc4053d4;
      16508: inst = 32'h8220000;
      16509: inst = 32'h10408000;
      16510: inst = 32'hc4053d5;
      16511: inst = 32'h8220000;
      16512: inst = 32'h10408000;
      16513: inst = 32'hc4053d6;
      16514: inst = 32'h8220000;
      16515: inst = 32'h10408000;
      16516: inst = 32'hc4053d7;
      16517: inst = 32'h8220000;
      16518: inst = 32'h10408000;
      16519: inst = 32'hc4053d8;
      16520: inst = 32'h8220000;
      16521: inst = 32'h10408000;
      16522: inst = 32'hc4053ea;
      16523: inst = 32'h8220000;
      16524: inst = 32'h10408000;
      16525: inst = 32'hc4053eb;
      16526: inst = 32'h8220000;
      16527: inst = 32'h10408000;
      16528: inst = 32'hc4053ec;
      16529: inst = 32'h8220000;
      16530: inst = 32'h10408000;
      16531: inst = 32'hc4053ed;
      16532: inst = 32'h8220000;
      16533: inst = 32'h10408000;
      16534: inst = 32'hc4053ee;
      16535: inst = 32'h8220000;
      16536: inst = 32'h10408000;
      16537: inst = 32'hc4053ef;
      16538: inst = 32'h8220000;
      16539: inst = 32'h10408000;
      16540: inst = 32'hc4053f0;
      16541: inst = 32'h8220000;
      16542: inst = 32'h10408000;
      16543: inst = 32'hc4053f1;
      16544: inst = 32'h8220000;
      16545: inst = 32'h10408000;
      16546: inst = 32'hc4053f2;
      16547: inst = 32'h8220000;
      16548: inst = 32'h10408000;
      16549: inst = 32'hc4053f3;
      16550: inst = 32'h8220000;
      16551: inst = 32'h10408000;
      16552: inst = 32'hc4053f4;
      16553: inst = 32'h8220000;
      16554: inst = 32'h10408000;
      16555: inst = 32'hc4053f5;
      16556: inst = 32'h8220000;
      16557: inst = 32'h10408000;
      16558: inst = 32'hc405407;
      16559: inst = 32'h8220000;
      16560: inst = 32'h10408000;
      16561: inst = 32'hc405408;
      16562: inst = 32'h8220000;
      16563: inst = 32'h10408000;
      16564: inst = 32'hc405409;
      16565: inst = 32'h8220000;
      16566: inst = 32'h10408000;
      16567: inst = 32'hc40540a;
      16568: inst = 32'h8220000;
      16569: inst = 32'h10408000;
      16570: inst = 32'hc40540b;
      16571: inst = 32'h8220000;
      16572: inst = 32'h10408000;
      16573: inst = 32'hc40540c;
      16574: inst = 32'h8220000;
      16575: inst = 32'h10408000;
      16576: inst = 32'hc40540d;
      16577: inst = 32'h8220000;
      16578: inst = 32'h10408000;
      16579: inst = 32'hc40540e;
      16580: inst = 32'h8220000;
      16581: inst = 32'h10408000;
      16582: inst = 32'hc40540f;
      16583: inst = 32'h8220000;
      16584: inst = 32'h10408000;
      16585: inst = 32'hc405410;
      16586: inst = 32'h8220000;
      16587: inst = 32'h10408000;
      16588: inst = 32'hc405411;
      16589: inst = 32'h8220000;
      16590: inst = 32'h10408000;
      16591: inst = 32'hc405412;
      16592: inst = 32'h8220000;
      16593: inst = 32'h10408000;
      16594: inst = 32'hc405413;
      16595: inst = 32'h8220000;
      16596: inst = 32'h10408000;
      16597: inst = 32'hc405414;
      16598: inst = 32'h8220000;
      16599: inst = 32'h10408000;
      16600: inst = 32'hc405415;
      16601: inst = 32'h8220000;
      16602: inst = 32'h10408000;
      16603: inst = 32'hc405416;
      16604: inst = 32'h8220000;
      16605: inst = 32'h10408000;
      16606: inst = 32'hc405417;
      16607: inst = 32'h8220000;
      16608: inst = 32'h10408000;
      16609: inst = 32'hc405418;
      16610: inst = 32'h8220000;
      16611: inst = 32'h10408000;
      16612: inst = 32'hc405419;
      16613: inst = 32'h8220000;
      16614: inst = 32'h10408000;
      16615: inst = 32'hc40541a;
      16616: inst = 32'h8220000;
      16617: inst = 32'h10408000;
      16618: inst = 32'hc40541b;
      16619: inst = 32'h8220000;
      16620: inst = 32'h10408000;
      16621: inst = 32'hc40541c;
      16622: inst = 32'h8220000;
      16623: inst = 32'h10408000;
      16624: inst = 32'hc40541d;
      16625: inst = 32'h8220000;
      16626: inst = 32'h10408000;
      16627: inst = 32'hc40541e;
      16628: inst = 32'h8220000;
      16629: inst = 32'h10408000;
      16630: inst = 32'hc40541f;
      16631: inst = 32'h8220000;
      16632: inst = 32'h10408000;
      16633: inst = 32'hc405420;
      16634: inst = 32'h8220000;
      16635: inst = 32'h10408000;
      16636: inst = 32'hc405421;
      16637: inst = 32'h8220000;
      16638: inst = 32'h10408000;
      16639: inst = 32'hc405422;
      16640: inst = 32'h8220000;
      16641: inst = 32'h10408000;
      16642: inst = 32'hc405423;
      16643: inst = 32'h8220000;
      16644: inst = 32'h10408000;
      16645: inst = 32'hc405424;
      16646: inst = 32'h8220000;
      16647: inst = 32'h10408000;
      16648: inst = 32'hc405425;
      16649: inst = 32'h8220000;
      16650: inst = 32'h10408000;
      16651: inst = 32'hc405426;
      16652: inst = 32'h8220000;
      16653: inst = 32'h10408000;
      16654: inst = 32'hc405427;
      16655: inst = 32'h8220000;
      16656: inst = 32'h10408000;
      16657: inst = 32'hc405428;
      16658: inst = 32'h8220000;
      16659: inst = 32'h10408000;
      16660: inst = 32'hc405429;
      16661: inst = 32'h8220000;
      16662: inst = 32'h10408000;
      16663: inst = 32'hc40542a;
      16664: inst = 32'h8220000;
      16665: inst = 32'h10408000;
      16666: inst = 32'hc40542b;
      16667: inst = 32'h8220000;
      16668: inst = 32'h10408000;
      16669: inst = 32'hc40542c;
      16670: inst = 32'h8220000;
      16671: inst = 32'h10408000;
      16672: inst = 32'hc40542d;
      16673: inst = 32'h8220000;
      16674: inst = 32'h10408000;
      16675: inst = 32'hc40542e;
      16676: inst = 32'h8220000;
      16677: inst = 32'h10408000;
      16678: inst = 32'hc40542f;
      16679: inst = 32'h8220000;
      16680: inst = 32'h10408000;
      16681: inst = 32'hc405430;
      16682: inst = 32'h8220000;
      16683: inst = 32'h10408000;
      16684: inst = 32'hc405431;
      16685: inst = 32'h8220000;
      16686: inst = 32'h10408000;
      16687: inst = 32'hc405432;
      16688: inst = 32'h8220000;
      16689: inst = 32'h10408000;
      16690: inst = 32'hc405433;
      16691: inst = 32'h8220000;
      16692: inst = 32'h10408000;
      16693: inst = 32'hc405434;
      16694: inst = 32'h8220000;
      16695: inst = 32'h10408000;
      16696: inst = 32'hc405435;
      16697: inst = 32'h8220000;
      16698: inst = 32'h10408000;
      16699: inst = 32'hc405436;
      16700: inst = 32'h8220000;
      16701: inst = 32'h10408000;
      16702: inst = 32'hc405437;
      16703: inst = 32'h8220000;
      16704: inst = 32'h10408000;
      16705: inst = 32'hc405438;
      16706: inst = 32'h8220000;
      16707: inst = 32'h10408000;
      16708: inst = 32'hc40544a;
      16709: inst = 32'h8220000;
      16710: inst = 32'h10408000;
      16711: inst = 32'hc40544b;
      16712: inst = 32'h8220000;
      16713: inst = 32'h10408000;
      16714: inst = 32'hc40544c;
      16715: inst = 32'h8220000;
      16716: inst = 32'h10408000;
      16717: inst = 32'hc40544d;
      16718: inst = 32'h8220000;
      16719: inst = 32'h10408000;
      16720: inst = 32'hc40544e;
      16721: inst = 32'h8220000;
      16722: inst = 32'h10408000;
      16723: inst = 32'hc40544f;
      16724: inst = 32'h8220000;
      16725: inst = 32'h10408000;
      16726: inst = 32'hc405450;
      16727: inst = 32'h8220000;
      16728: inst = 32'h10408000;
      16729: inst = 32'hc405451;
      16730: inst = 32'h8220000;
      16731: inst = 32'h10408000;
      16732: inst = 32'hc405452;
      16733: inst = 32'h8220000;
      16734: inst = 32'h10408000;
      16735: inst = 32'hc405453;
      16736: inst = 32'h8220000;
      16737: inst = 32'h10408000;
      16738: inst = 32'hc405454;
      16739: inst = 32'h8220000;
      16740: inst = 32'h10408000;
      16741: inst = 32'hc405455;
      16742: inst = 32'h8220000;
      16743: inst = 32'h10408000;
      16744: inst = 32'hc405467;
      16745: inst = 32'h8220000;
      16746: inst = 32'h10408000;
      16747: inst = 32'hc405468;
      16748: inst = 32'h8220000;
      16749: inst = 32'h10408000;
      16750: inst = 32'hc405469;
      16751: inst = 32'h8220000;
      16752: inst = 32'h10408000;
      16753: inst = 32'hc40546a;
      16754: inst = 32'h8220000;
      16755: inst = 32'h10408000;
      16756: inst = 32'hc40546b;
      16757: inst = 32'h8220000;
      16758: inst = 32'h10408000;
      16759: inst = 32'hc40546c;
      16760: inst = 32'h8220000;
      16761: inst = 32'h10408000;
      16762: inst = 32'hc40546d;
      16763: inst = 32'h8220000;
      16764: inst = 32'h10408000;
      16765: inst = 32'hc40546e;
      16766: inst = 32'h8220000;
      16767: inst = 32'h10408000;
      16768: inst = 32'hc40546f;
      16769: inst = 32'h8220000;
      16770: inst = 32'h10408000;
      16771: inst = 32'hc405470;
      16772: inst = 32'h8220000;
      16773: inst = 32'h10408000;
      16774: inst = 32'hc405471;
      16775: inst = 32'h8220000;
      16776: inst = 32'h10408000;
      16777: inst = 32'hc405472;
      16778: inst = 32'h8220000;
      16779: inst = 32'h10408000;
      16780: inst = 32'hc405473;
      16781: inst = 32'h8220000;
      16782: inst = 32'h10408000;
      16783: inst = 32'hc405474;
      16784: inst = 32'h8220000;
      16785: inst = 32'h10408000;
      16786: inst = 32'hc405475;
      16787: inst = 32'h8220000;
      16788: inst = 32'h10408000;
      16789: inst = 32'hc405476;
      16790: inst = 32'h8220000;
      16791: inst = 32'h10408000;
      16792: inst = 32'hc405477;
      16793: inst = 32'h8220000;
      16794: inst = 32'h10408000;
      16795: inst = 32'hc405478;
      16796: inst = 32'h8220000;
      16797: inst = 32'h10408000;
      16798: inst = 32'hc405479;
      16799: inst = 32'h8220000;
      16800: inst = 32'h10408000;
      16801: inst = 32'hc40547a;
      16802: inst = 32'h8220000;
      16803: inst = 32'h10408000;
      16804: inst = 32'hc40547b;
      16805: inst = 32'h8220000;
      16806: inst = 32'h10408000;
      16807: inst = 32'hc40547c;
      16808: inst = 32'h8220000;
      16809: inst = 32'h10408000;
      16810: inst = 32'hc40547d;
      16811: inst = 32'h8220000;
      16812: inst = 32'h10408000;
      16813: inst = 32'hc40547e;
      16814: inst = 32'h8220000;
      16815: inst = 32'h10408000;
      16816: inst = 32'hc40547f;
      16817: inst = 32'h8220000;
      16818: inst = 32'h10408000;
      16819: inst = 32'hc405480;
      16820: inst = 32'h8220000;
      16821: inst = 32'h10408000;
      16822: inst = 32'hc405481;
      16823: inst = 32'h8220000;
      16824: inst = 32'h10408000;
      16825: inst = 32'hc405482;
      16826: inst = 32'h8220000;
      16827: inst = 32'h10408000;
      16828: inst = 32'hc405483;
      16829: inst = 32'h8220000;
      16830: inst = 32'h10408000;
      16831: inst = 32'hc405484;
      16832: inst = 32'h8220000;
      16833: inst = 32'h10408000;
      16834: inst = 32'hc405485;
      16835: inst = 32'h8220000;
      16836: inst = 32'h10408000;
      16837: inst = 32'hc405486;
      16838: inst = 32'h8220000;
      16839: inst = 32'h10408000;
      16840: inst = 32'hc405487;
      16841: inst = 32'h8220000;
      16842: inst = 32'h10408000;
      16843: inst = 32'hc405488;
      16844: inst = 32'h8220000;
      16845: inst = 32'h10408000;
      16846: inst = 32'hc405489;
      16847: inst = 32'h8220000;
      16848: inst = 32'h10408000;
      16849: inst = 32'hc40548a;
      16850: inst = 32'h8220000;
      16851: inst = 32'h10408000;
      16852: inst = 32'hc40548b;
      16853: inst = 32'h8220000;
      16854: inst = 32'h10408000;
      16855: inst = 32'hc40548c;
      16856: inst = 32'h8220000;
      16857: inst = 32'h10408000;
      16858: inst = 32'hc40548d;
      16859: inst = 32'h8220000;
      16860: inst = 32'h10408000;
      16861: inst = 32'hc40548e;
      16862: inst = 32'h8220000;
      16863: inst = 32'h10408000;
      16864: inst = 32'hc40548f;
      16865: inst = 32'h8220000;
      16866: inst = 32'h10408000;
      16867: inst = 32'hc405490;
      16868: inst = 32'h8220000;
      16869: inst = 32'h10408000;
      16870: inst = 32'hc405491;
      16871: inst = 32'h8220000;
      16872: inst = 32'h10408000;
      16873: inst = 32'hc405492;
      16874: inst = 32'h8220000;
      16875: inst = 32'h10408000;
      16876: inst = 32'hc405493;
      16877: inst = 32'h8220000;
      16878: inst = 32'h10408000;
      16879: inst = 32'hc405494;
      16880: inst = 32'h8220000;
      16881: inst = 32'h10408000;
      16882: inst = 32'hc405495;
      16883: inst = 32'h8220000;
      16884: inst = 32'h10408000;
      16885: inst = 32'hc405496;
      16886: inst = 32'h8220000;
      16887: inst = 32'h10408000;
      16888: inst = 32'hc405497;
      16889: inst = 32'h8220000;
      16890: inst = 32'h10408000;
      16891: inst = 32'hc4054aa;
      16892: inst = 32'h8220000;
      16893: inst = 32'h10408000;
      16894: inst = 32'hc4054ab;
      16895: inst = 32'h8220000;
      16896: inst = 32'h10408000;
      16897: inst = 32'hc4054ac;
      16898: inst = 32'h8220000;
      16899: inst = 32'h10408000;
      16900: inst = 32'hc4054ad;
      16901: inst = 32'h8220000;
      16902: inst = 32'h10408000;
      16903: inst = 32'hc4054ae;
      16904: inst = 32'h8220000;
      16905: inst = 32'h10408000;
      16906: inst = 32'hc4054af;
      16907: inst = 32'h8220000;
      16908: inst = 32'h10408000;
      16909: inst = 32'hc4054b0;
      16910: inst = 32'h8220000;
      16911: inst = 32'h10408000;
      16912: inst = 32'hc4054b1;
      16913: inst = 32'h8220000;
      16914: inst = 32'h10408000;
      16915: inst = 32'hc4054b2;
      16916: inst = 32'h8220000;
      16917: inst = 32'h10408000;
      16918: inst = 32'hc4054b3;
      16919: inst = 32'h8220000;
      16920: inst = 32'h10408000;
      16921: inst = 32'hc4054b4;
      16922: inst = 32'h8220000;
      16923: inst = 32'h10408000;
      16924: inst = 32'hc4054b5;
      16925: inst = 32'h8220000;
      16926: inst = 32'h10408000;
      16927: inst = 32'hc4054c8;
      16928: inst = 32'h8220000;
      16929: inst = 32'h10408000;
      16930: inst = 32'hc4054c9;
      16931: inst = 32'h8220000;
      16932: inst = 32'h10408000;
      16933: inst = 32'hc4054ca;
      16934: inst = 32'h8220000;
      16935: inst = 32'h10408000;
      16936: inst = 32'hc4054cb;
      16937: inst = 32'h8220000;
      16938: inst = 32'h10408000;
      16939: inst = 32'hc4054cc;
      16940: inst = 32'h8220000;
      16941: inst = 32'h10408000;
      16942: inst = 32'hc4054cd;
      16943: inst = 32'h8220000;
      16944: inst = 32'h10408000;
      16945: inst = 32'hc4054ce;
      16946: inst = 32'h8220000;
      16947: inst = 32'h10408000;
      16948: inst = 32'hc4054cf;
      16949: inst = 32'h8220000;
      16950: inst = 32'h10408000;
      16951: inst = 32'hc4054d0;
      16952: inst = 32'h8220000;
      16953: inst = 32'h10408000;
      16954: inst = 32'hc4054d1;
      16955: inst = 32'h8220000;
      16956: inst = 32'h10408000;
      16957: inst = 32'hc4054d2;
      16958: inst = 32'h8220000;
      16959: inst = 32'h10408000;
      16960: inst = 32'hc4054d3;
      16961: inst = 32'h8220000;
      16962: inst = 32'h10408000;
      16963: inst = 32'hc4054d4;
      16964: inst = 32'h8220000;
      16965: inst = 32'h10408000;
      16966: inst = 32'hc4054d5;
      16967: inst = 32'h8220000;
      16968: inst = 32'h10408000;
      16969: inst = 32'hc4054d6;
      16970: inst = 32'h8220000;
      16971: inst = 32'h10408000;
      16972: inst = 32'hc4054d7;
      16973: inst = 32'h8220000;
      16974: inst = 32'h10408000;
      16975: inst = 32'hc4054d8;
      16976: inst = 32'h8220000;
      16977: inst = 32'h10408000;
      16978: inst = 32'hc4054d9;
      16979: inst = 32'h8220000;
      16980: inst = 32'h10408000;
      16981: inst = 32'hc4054da;
      16982: inst = 32'h8220000;
      16983: inst = 32'h10408000;
      16984: inst = 32'hc4054db;
      16985: inst = 32'h8220000;
      16986: inst = 32'h10408000;
      16987: inst = 32'hc4054dc;
      16988: inst = 32'h8220000;
      16989: inst = 32'h10408000;
      16990: inst = 32'hc4054dd;
      16991: inst = 32'h8220000;
      16992: inst = 32'h10408000;
      16993: inst = 32'hc4054de;
      16994: inst = 32'h8220000;
      16995: inst = 32'h10408000;
      16996: inst = 32'hc4054df;
      16997: inst = 32'h8220000;
      16998: inst = 32'h10408000;
      16999: inst = 32'hc4054e0;
      17000: inst = 32'h8220000;
      17001: inst = 32'h10408000;
      17002: inst = 32'hc4054e1;
      17003: inst = 32'h8220000;
      17004: inst = 32'h10408000;
      17005: inst = 32'hc4054e2;
      17006: inst = 32'h8220000;
      17007: inst = 32'h10408000;
      17008: inst = 32'hc4054e3;
      17009: inst = 32'h8220000;
      17010: inst = 32'h10408000;
      17011: inst = 32'hc4054e4;
      17012: inst = 32'h8220000;
      17013: inst = 32'h10408000;
      17014: inst = 32'hc4054e5;
      17015: inst = 32'h8220000;
      17016: inst = 32'h10408000;
      17017: inst = 32'hc4054e6;
      17018: inst = 32'h8220000;
      17019: inst = 32'h10408000;
      17020: inst = 32'hc4054e7;
      17021: inst = 32'h8220000;
      17022: inst = 32'h10408000;
      17023: inst = 32'hc4054e8;
      17024: inst = 32'h8220000;
      17025: inst = 32'h10408000;
      17026: inst = 32'hc4054e9;
      17027: inst = 32'h8220000;
      17028: inst = 32'h10408000;
      17029: inst = 32'hc4054ea;
      17030: inst = 32'h8220000;
      17031: inst = 32'h10408000;
      17032: inst = 32'hc4054eb;
      17033: inst = 32'h8220000;
      17034: inst = 32'h10408000;
      17035: inst = 32'hc4054ec;
      17036: inst = 32'h8220000;
      17037: inst = 32'h10408000;
      17038: inst = 32'hc4054ed;
      17039: inst = 32'h8220000;
      17040: inst = 32'h10408000;
      17041: inst = 32'hc4054ee;
      17042: inst = 32'h8220000;
      17043: inst = 32'h10408000;
      17044: inst = 32'hc4054ef;
      17045: inst = 32'h8220000;
      17046: inst = 32'h10408000;
      17047: inst = 32'hc4054f0;
      17048: inst = 32'h8220000;
      17049: inst = 32'h10408000;
      17050: inst = 32'hc4054f1;
      17051: inst = 32'h8220000;
      17052: inst = 32'h10408000;
      17053: inst = 32'hc4054f2;
      17054: inst = 32'h8220000;
      17055: inst = 32'h10408000;
      17056: inst = 32'hc4054f3;
      17057: inst = 32'h8220000;
      17058: inst = 32'h10408000;
      17059: inst = 32'hc4054f4;
      17060: inst = 32'h8220000;
      17061: inst = 32'h10408000;
      17062: inst = 32'hc4054f5;
      17063: inst = 32'h8220000;
      17064: inst = 32'h10408000;
      17065: inst = 32'hc4054f6;
      17066: inst = 32'h8220000;
      17067: inst = 32'h10408000;
      17068: inst = 32'hc40550a;
      17069: inst = 32'h8220000;
      17070: inst = 32'h10408000;
      17071: inst = 32'hc40550b;
      17072: inst = 32'h8220000;
      17073: inst = 32'h10408000;
      17074: inst = 32'hc40550c;
      17075: inst = 32'h8220000;
      17076: inst = 32'h10408000;
      17077: inst = 32'hc40550d;
      17078: inst = 32'h8220000;
      17079: inst = 32'h10408000;
      17080: inst = 32'hc40550e;
      17081: inst = 32'h8220000;
      17082: inst = 32'h10408000;
      17083: inst = 32'hc40550f;
      17084: inst = 32'h8220000;
      17085: inst = 32'h10408000;
      17086: inst = 32'hc405510;
      17087: inst = 32'h8220000;
      17088: inst = 32'h10408000;
      17089: inst = 32'hc405511;
      17090: inst = 32'h8220000;
      17091: inst = 32'h10408000;
      17092: inst = 32'hc405512;
      17093: inst = 32'h8220000;
      17094: inst = 32'h10408000;
      17095: inst = 32'hc405513;
      17096: inst = 32'h8220000;
      17097: inst = 32'h10408000;
      17098: inst = 32'hc405514;
      17099: inst = 32'h8220000;
      17100: inst = 32'h10408000;
      17101: inst = 32'hc405515;
      17102: inst = 32'h8220000;
      17103: inst = 32'h10408000;
      17104: inst = 32'hc405529;
      17105: inst = 32'h8220000;
      17106: inst = 32'h10408000;
      17107: inst = 32'hc40552a;
      17108: inst = 32'h8220000;
      17109: inst = 32'h10408000;
      17110: inst = 32'hc40552b;
      17111: inst = 32'h8220000;
      17112: inst = 32'h10408000;
      17113: inst = 32'hc40552c;
      17114: inst = 32'h8220000;
      17115: inst = 32'h10408000;
      17116: inst = 32'hc40552d;
      17117: inst = 32'h8220000;
      17118: inst = 32'h10408000;
      17119: inst = 32'hc40552e;
      17120: inst = 32'h8220000;
      17121: inst = 32'h10408000;
      17122: inst = 32'hc40552f;
      17123: inst = 32'h8220000;
      17124: inst = 32'h10408000;
      17125: inst = 32'hc405530;
      17126: inst = 32'h8220000;
      17127: inst = 32'h10408000;
      17128: inst = 32'hc405531;
      17129: inst = 32'h8220000;
      17130: inst = 32'h10408000;
      17131: inst = 32'hc405532;
      17132: inst = 32'h8220000;
      17133: inst = 32'h10408000;
      17134: inst = 32'hc405533;
      17135: inst = 32'h8220000;
      17136: inst = 32'h10408000;
      17137: inst = 32'hc405534;
      17138: inst = 32'h8220000;
      17139: inst = 32'h10408000;
      17140: inst = 32'hc405535;
      17141: inst = 32'h8220000;
      17142: inst = 32'h10408000;
      17143: inst = 32'hc405536;
      17144: inst = 32'h8220000;
      17145: inst = 32'h10408000;
      17146: inst = 32'hc405537;
      17147: inst = 32'h8220000;
      17148: inst = 32'h10408000;
      17149: inst = 32'hc405538;
      17150: inst = 32'h8220000;
      17151: inst = 32'h10408000;
      17152: inst = 32'hc405539;
      17153: inst = 32'h8220000;
      17154: inst = 32'h10408000;
      17155: inst = 32'hc40553a;
      17156: inst = 32'h8220000;
      17157: inst = 32'h10408000;
      17158: inst = 32'hc40553b;
      17159: inst = 32'h8220000;
      17160: inst = 32'h10408000;
      17161: inst = 32'hc40553c;
      17162: inst = 32'h8220000;
      17163: inst = 32'h10408000;
      17164: inst = 32'hc40553d;
      17165: inst = 32'h8220000;
      17166: inst = 32'h10408000;
      17167: inst = 32'hc40553e;
      17168: inst = 32'h8220000;
      17169: inst = 32'h10408000;
      17170: inst = 32'hc40553f;
      17171: inst = 32'h8220000;
      17172: inst = 32'h10408000;
      17173: inst = 32'hc405540;
      17174: inst = 32'h8220000;
      17175: inst = 32'h10408000;
      17176: inst = 32'hc405541;
      17177: inst = 32'h8220000;
      17178: inst = 32'h10408000;
      17179: inst = 32'hc405542;
      17180: inst = 32'h8220000;
      17181: inst = 32'h10408000;
      17182: inst = 32'hc405543;
      17183: inst = 32'h8220000;
      17184: inst = 32'h10408000;
      17185: inst = 32'hc405544;
      17186: inst = 32'h8220000;
      17187: inst = 32'h10408000;
      17188: inst = 32'hc405545;
      17189: inst = 32'h8220000;
      17190: inst = 32'h10408000;
      17191: inst = 32'hc405546;
      17192: inst = 32'h8220000;
      17193: inst = 32'h10408000;
      17194: inst = 32'hc405547;
      17195: inst = 32'h8220000;
      17196: inst = 32'h10408000;
      17197: inst = 32'hc405548;
      17198: inst = 32'h8220000;
      17199: inst = 32'h10408000;
      17200: inst = 32'hc405549;
      17201: inst = 32'h8220000;
      17202: inst = 32'h10408000;
      17203: inst = 32'hc40554a;
      17204: inst = 32'h8220000;
      17205: inst = 32'h10408000;
      17206: inst = 32'hc40554b;
      17207: inst = 32'h8220000;
      17208: inst = 32'h10408000;
      17209: inst = 32'hc40554c;
      17210: inst = 32'h8220000;
      17211: inst = 32'h10408000;
      17212: inst = 32'hc40554d;
      17213: inst = 32'h8220000;
      17214: inst = 32'h10408000;
      17215: inst = 32'hc40554e;
      17216: inst = 32'h8220000;
      17217: inst = 32'h10408000;
      17218: inst = 32'hc40554f;
      17219: inst = 32'h8220000;
      17220: inst = 32'h10408000;
      17221: inst = 32'hc405550;
      17222: inst = 32'h8220000;
      17223: inst = 32'h10408000;
      17224: inst = 32'hc405551;
      17225: inst = 32'h8220000;
      17226: inst = 32'h10408000;
      17227: inst = 32'hc405552;
      17228: inst = 32'h8220000;
      17229: inst = 32'h10408000;
      17230: inst = 32'hc405553;
      17231: inst = 32'h8220000;
      17232: inst = 32'h10408000;
      17233: inst = 32'hc405554;
      17234: inst = 32'h8220000;
      17235: inst = 32'h10408000;
      17236: inst = 32'hc405555;
      17237: inst = 32'h8220000;
      17238: inst = 32'h10408000;
      17239: inst = 32'hc40556a;
      17240: inst = 32'h8220000;
      17241: inst = 32'h10408000;
      17242: inst = 32'hc40556b;
      17243: inst = 32'h8220000;
      17244: inst = 32'h10408000;
      17245: inst = 32'hc40556c;
      17246: inst = 32'h8220000;
      17247: inst = 32'h10408000;
      17248: inst = 32'hc40556d;
      17249: inst = 32'h8220000;
      17250: inst = 32'h10408000;
      17251: inst = 32'hc40556e;
      17252: inst = 32'h8220000;
      17253: inst = 32'h10408000;
      17254: inst = 32'hc40556f;
      17255: inst = 32'h8220000;
      17256: inst = 32'h10408000;
      17257: inst = 32'hc405570;
      17258: inst = 32'h8220000;
      17259: inst = 32'h10408000;
      17260: inst = 32'hc405571;
      17261: inst = 32'h8220000;
      17262: inst = 32'h10408000;
      17263: inst = 32'hc405572;
      17264: inst = 32'h8220000;
      17265: inst = 32'h10408000;
      17266: inst = 32'hc405573;
      17267: inst = 32'h8220000;
      17268: inst = 32'h10408000;
      17269: inst = 32'hc405574;
      17270: inst = 32'h8220000;
      17271: inst = 32'h10408000;
      17272: inst = 32'hc405575;
      17273: inst = 32'h8220000;
      17274: inst = 32'h10408000;
      17275: inst = 32'hc40558a;
      17276: inst = 32'h8220000;
      17277: inst = 32'h10408000;
      17278: inst = 32'hc40558b;
      17279: inst = 32'h8220000;
      17280: inst = 32'h10408000;
      17281: inst = 32'hc40558c;
      17282: inst = 32'h8220000;
      17283: inst = 32'h10408000;
      17284: inst = 32'hc40558d;
      17285: inst = 32'h8220000;
      17286: inst = 32'h10408000;
      17287: inst = 32'hc40558e;
      17288: inst = 32'h8220000;
      17289: inst = 32'h10408000;
      17290: inst = 32'hc40558f;
      17291: inst = 32'h8220000;
      17292: inst = 32'h10408000;
      17293: inst = 32'hc405590;
      17294: inst = 32'h8220000;
      17295: inst = 32'h10408000;
      17296: inst = 32'hc405591;
      17297: inst = 32'h8220000;
      17298: inst = 32'h10408000;
      17299: inst = 32'hc405592;
      17300: inst = 32'h8220000;
      17301: inst = 32'h10408000;
      17302: inst = 32'hc405593;
      17303: inst = 32'h8220000;
      17304: inst = 32'h10408000;
      17305: inst = 32'hc405594;
      17306: inst = 32'h8220000;
      17307: inst = 32'h10408000;
      17308: inst = 32'hc405595;
      17309: inst = 32'h8220000;
      17310: inst = 32'h10408000;
      17311: inst = 32'hc405596;
      17312: inst = 32'h8220000;
      17313: inst = 32'h10408000;
      17314: inst = 32'hc405597;
      17315: inst = 32'h8220000;
      17316: inst = 32'h10408000;
      17317: inst = 32'hc405598;
      17318: inst = 32'h8220000;
      17319: inst = 32'h10408000;
      17320: inst = 32'hc405599;
      17321: inst = 32'h8220000;
      17322: inst = 32'h10408000;
      17323: inst = 32'hc40559a;
      17324: inst = 32'h8220000;
      17325: inst = 32'h10408000;
      17326: inst = 32'hc40559b;
      17327: inst = 32'h8220000;
      17328: inst = 32'h10408000;
      17329: inst = 32'hc40559c;
      17330: inst = 32'h8220000;
      17331: inst = 32'h10408000;
      17332: inst = 32'hc40559d;
      17333: inst = 32'h8220000;
      17334: inst = 32'h10408000;
      17335: inst = 32'hc40559e;
      17336: inst = 32'h8220000;
      17337: inst = 32'h10408000;
      17338: inst = 32'hc40559f;
      17339: inst = 32'h8220000;
      17340: inst = 32'h10408000;
      17341: inst = 32'hc4055a0;
      17342: inst = 32'h8220000;
      17343: inst = 32'h10408000;
      17344: inst = 32'hc4055a1;
      17345: inst = 32'h8220000;
      17346: inst = 32'h10408000;
      17347: inst = 32'hc4055a2;
      17348: inst = 32'h8220000;
      17349: inst = 32'h10408000;
      17350: inst = 32'hc4055a3;
      17351: inst = 32'h8220000;
      17352: inst = 32'h10408000;
      17353: inst = 32'hc4055a4;
      17354: inst = 32'h8220000;
      17355: inst = 32'h10408000;
      17356: inst = 32'hc4055a5;
      17357: inst = 32'h8220000;
      17358: inst = 32'h10408000;
      17359: inst = 32'hc4055a6;
      17360: inst = 32'h8220000;
      17361: inst = 32'h10408000;
      17362: inst = 32'hc4055a7;
      17363: inst = 32'h8220000;
      17364: inst = 32'h10408000;
      17365: inst = 32'hc4055a8;
      17366: inst = 32'h8220000;
      17367: inst = 32'h10408000;
      17368: inst = 32'hc4055a9;
      17369: inst = 32'h8220000;
      17370: inst = 32'h10408000;
      17371: inst = 32'hc4055aa;
      17372: inst = 32'h8220000;
      17373: inst = 32'h10408000;
      17374: inst = 32'hc4055ab;
      17375: inst = 32'h8220000;
      17376: inst = 32'h10408000;
      17377: inst = 32'hc4055ac;
      17378: inst = 32'h8220000;
      17379: inst = 32'h10408000;
      17380: inst = 32'hc4055ad;
      17381: inst = 32'h8220000;
      17382: inst = 32'h10408000;
      17383: inst = 32'hc4055ae;
      17384: inst = 32'h8220000;
      17385: inst = 32'h10408000;
      17386: inst = 32'hc4055af;
      17387: inst = 32'h8220000;
      17388: inst = 32'h10408000;
      17389: inst = 32'hc4055b0;
      17390: inst = 32'h8220000;
      17391: inst = 32'h10408000;
      17392: inst = 32'hc4055b1;
      17393: inst = 32'h8220000;
      17394: inst = 32'h10408000;
      17395: inst = 32'hc4055b2;
      17396: inst = 32'h8220000;
      17397: inst = 32'h10408000;
      17398: inst = 32'hc4055b3;
      17399: inst = 32'h8220000;
      17400: inst = 32'h10408000;
      17401: inst = 32'hc4055b4;
      17402: inst = 32'h8220000;
      17403: inst = 32'h10408000;
      17404: inst = 32'hc4055ca;
      17405: inst = 32'h8220000;
      17406: inst = 32'h10408000;
      17407: inst = 32'hc4055cb;
      17408: inst = 32'h8220000;
      17409: inst = 32'h10408000;
      17410: inst = 32'hc4055cc;
      17411: inst = 32'h8220000;
      17412: inst = 32'h10408000;
      17413: inst = 32'hc4055cd;
      17414: inst = 32'h8220000;
      17415: inst = 32'h10408000;
      17416: inst = 32'hc4055ce;
      17417: inst = 32'h8220000;
      17418: inst = 32'h10408000;
      17419: inst = 32'hc4055cf;
      17420: inst = 32'h8220000;
      17421: inst = 32'h10408000;
      17422: inst = 32'hc4055d0;
      17423: inst = 32'h8220000;
      17424: inst = 32'h10408000;
      17425: inst = 32'hc4055d1;
      17426: inst = 32'h8220000;
      17427: inst = 32'h10408000;
      17428: inst = 32'hc4055d2;
      17429: inst = 32'h8220000;
      17430: inst = 32'h10408000;
      17431: inst = 32'hc4055d3;
      17432: inst = 32'h8220000;
      17433: inst = 32'h10408000;
      17434: inst = 32'hc4055d4;
      17435: inst = 32'h8220000;
      17436: inst = 32'h10408000;
      17437: inst = 32'hc4055d5;
      17438: inst = 32'h8220000;
      17439: inst = 32'h10408000;
      17440: inst = 32'hc4055eb;
      17441: inst = 32'h8220000;
      17442: inst = 32'h10408000;
      17443: inst = 32'hc4055ec;
      17444: inst = 32'h8220000;
      17445: inst = 32'h10408000;
      17446: inst = 32'hc4055ed;
      17447: inst = 32'h8220000;
      17448: inst = 32'h10408000;
      17449: inst = 32'hc4055ee;
      17450: inst = 32'h8220000;
      17451: inst = 32'h10408000;
      17452: inst = 32'hc4055ef;
      17453: inst = 32'h8220000;
      17454: inst = 32'h10408000;
      17455: inst = 32'hc4055f0;
      17456: inst = 32'h8220000;
      17457: inst = 32'h10408000;
      17458: inst = 32'hc4055f1;
      17459: inst = 32'h8220000;
      17460: inst = 32'h10408000;
      17461: inst = 32'hc4055f2;
      17462: inst = 32'h8220000;
      17463: inst = 32'h10408000;
      17464: inst = 32'hc4055f3;
      17465: inst = 32'h8220000;
      17466: inst = 32'h10408000;
      17467: inst = 32'hc4055f4;
      17468: inst = 32'h8220000;
      17469: inst = 32'h10408000;
      17470: inst = 32'hc4055f5;
      17471: inst = 32'h8220000;
      17472: inst = 32'h10408000;
      17473: inst = 32'hc4055f6;
      17474: inst = 32'h8220000;
      17475: inst = 32'h10408000;
      17476: inst = 32'hc4055f7;
      17477: inst = 32'h8220000;
      17478: inst = 32'h10408000;
      17479: inst = 32'hc4055f8;
      17480: inst = 32'h8220000;
      17481: inst = 32'h10408000;
      17482: inst = 32'hc4055f9;
      17483: inst = 32'h8220000;
      17484: inst = 32'h10408000;
      17485: inst = 32'hc4055fa;
      17486: inst = 32'h8220000;
      17487: inst = 32'h10408000;
      17488: inst = 32'hc4055fb;
      17489: inst = 32'h8220000;
      17490: inst = 32'h10408000;
      17491: inst = 32'hc4055fc;
      17492: inst = 32'h8220000;
      17493: inst = 32'h10408000;
      17494: inst = 32'hc4055fd;
      17495: inst = 32'h8220000;
      17496: inst = 32'h10408000;
      17497: inst = 32'hc4055fe;
      17498: inst = 32'h8220000;
      17499: inst = 32'h10408000;
      17500: inst = 32'hc4055ff;
      17501: inst = 32'h8220000;
      17502: inst = 32'h10408000;
      17503: inst = 32'hc405600;
      17504: inst = 32'h8220000;
      17505: inst = 32'h10408000;
      17506: inst = 32'hc405601;
      17507: inst = 32'h8220000;
      17508: inst = 32'h10408000;
      17509: inst = 32'hc405602;
      17510: inst = 32'h8220000;
      17511: inst = 32'h10408000;
      17512: inst = 32'hc405603;
      17513: inst = 32'h8220000;
      17514: inst = 32'h10408000;
      17515: inst = 32'hc405604;
      17516: inst = 32'h8220000;
      17517: inst = 32'h10408000;
      17518: inst = 32'hc405605;
      17519: inst = 32'h8220000;
      17520: inst = 32'h10408000;
      17521: inst = 32'hc405606;
      17522: inst = 32'h8220000;
      17523: inst = 32'h10408000;
      17524: inst = 32'hc405607;
      17525: inst = 32'h8220000;
      17526: inst = 32'h10408000;
      17527: inst = 32'hc405608;
      17528: inst = 32'h8220000;
      17529: inst = 32'h10408000;
      17530: inst = 32'hc405609;
      17531: inst = 32'h8220000;
      17532: inst = 32'h10408000;
      17533: inst = 32'hc40560a;
      17534: inst = 32'h8220000;
      17535: inst = 32'h10408000;
      17536: inst = 32'hc40560b;
      17537: inst = 32'h8220000;
      17538: inst = 32'h10408000;
      17539: inst = 32'hc40560c;
      17540: inst = 32'h8220000;
      17541: inst = 32'h10408000;
      17542: inst = 32'hc40560d;
      17543: inst = 32'h8220000;
      17544: inst = 32'h10408000;
      17545: inst = 32'hc40560e;
      17546: inst = 32'h8220000;
      17547: inst = 32'h10408000;
      17548: inst = 32'hc40560f;
      17549: inst = 32'h8220000;
      17550: inst = 32'h10408000;
      17551: inst = 32'hc405610;
      17552: inst = 32'h8220000;
      17553: inst = 32'h10408000;
      17554: inst = 32'hc405611;
      17555: inst = 32'h8220000;
      17556: inst = 32'h10408000;
      17557: inst = 32'hc405612;
      17558: inst = 32'h8220000;
      17559: inst = 32'h10408000;
      17560: inst = 32'hc405613;
      17561: inst = 32'h8220000;
      17562: inst = 32'h10408000;
      17563: inst = 32'hc405614;
      17564: inst = 32'h8220000;
      17565: inst = 32'h10408000;
      17566: inst = 32'hc40562a;
      17567: inst = 32'h8220000;
      17568: inst = 32'h10408000;
      17569: inst = 32'hc40562b;
      17570: inst = 32'h8220000;
      17571: inst = 32'h10408000;
      17572: inst = 32'hc40562c;
      17573: inst = 32'h8220000;
      17574: inst = 32'h10408000;
      17575: inst = 32'hc40562d;
      17576: inst = 32'h8220000;
      17577: inst = 32'h10408000;
      17578: inst = 32'hc40562e;
      17579: inst = 32'h8220000;
      17580: inst = 32'h10408000;
      17581: inst = 32'hc40562f;
      17582: inst = 32'h8220000;
      17583: inst = 32'h10408000;
      17584: inst = 32'hc405630;
      17585: inst = 32'h8220000;
      17586: inst = 32'h10408000;
      17587: inst = 32'hc405631;
      17588: inst = 32'h8220000;
      17589: inst = 32'h10408000;
      17590: inst = 32'hc405632;
      17591: inst = 32'h8220000;
      17592: inst = 32'h10408000;
      17593: inst = 32'hc405633;
      17594: inst = 32'h8220000;
      17595: inst = 32'h10408000;
      17596: inst = 32'hc405634;
      17597: inst = 32'h8220000;
      17598: inst = 32'h10408000;
      17599: inst = 32'hc405635;
      17600: inst = 32'h8220000;
      17601: inst = 32'h10408000;
      17602: inst = 32'hc40564b;
      17603: inst = 32'h8220000;
      17604: inst = 32'h10408000;
      17605: inst = 32'hc40564c;
      17606: inst = 32'h8220000;
      17607: inst = 32'h10408000;
      17608: inst = 32'hc40564d;
      17609: inst = 32'h8220000;
      17610: inst = 32'h10408000;
      17611: inst = 32'hc40564e;
      17612: inst = 32'h8220000;
      17613: inst = 32'h10408000;
      17614: inst = 32'hc40564f;
      17615: inst = 32'h8220000;
      17616: inst = 32'h10408000;
      17617: inst = 32'hc405650;
      17618: inst = 32'h8220000;
      17619: inst = 32'h10408000;
      17620: inst = 32'hc405651;
      17621: inst = 32'h8220000;
      17622: inst = 32'h10408000;
      17623: inst = 32'hc405652;
      17624: inst = 32'h8220000;
      17625: inst = 32'h10408000;
      17626: inst = 32'hc405653;
      17627: inst = 32'h8220000;
      17628: inst = 32'h10408000;
      17629: inst = 32'hc405654;
      17630: inst = 32'h8220000;
      17631: inst = 32'h10408000;
      17632: inst = 32'hc405655;
      17633: inst = 32'h8220000;
      17634: inst = 32'h10408000;
      17635: inst = 32'hc405656;
      17636: inst = 32'h8220000;
      17637: inst = 32'h10408000;
      17638: inst = 32'hc405657;
      17639: inst = 32'h8220000;
      17640: inst = 32'h10408000;
      17641: inst = 32'hc405658;
      17642: inst = 32'h8220000;
      17643: inst = 32'h10408000;
      17644: inst = 32'hc405659;
      17645: inst = 32'h8220000;
      17646: inst = 32'h10408000;
      17647: inst = 32'hc40565a;
      17648: inst = 32'h8220000;
      17649: inst = 32'h10408000;
      17650: inst = 32'hc40565b;
      17651: inst = 32'h8220000;
      17652: inst = 32'h10408000;
      17653: inst = 32'hc40565c;
      17654: inst = 32'h8220000;
      17655: inst = 32'h10408000;
      17656: inst = 32'hc40565d;
      17657: inst = 32'h8220000;
      17658: inst = 32'h10408000;
      17659: inst = 32'hc40565e;
      17660: inst = 32'h8220000;
      17661: inst = 32'h10408000;
      17662: inst = 32'hc40565f;
      17663: inst = 32'h8220000;
      17664: inst = 32'h10408000;
      17665: inst = 32'hc405660;
      17666: inst = 32'h8220000;
      17667: inst = 32'h10408000;
      17668: inst = 32'hc405661;
      17669: inst = 32'h8220000;
      17670: inst = 32'h10408000;
      17671: inst = 32'hc405662;
      17672: inst = 32'h8220000;
      17673: inst = 32'h10408000;
      17674: inst = 32'hc405663;
      17675: inst = 32'h8220000;
      17676: inst = 32'h10408000;
      17677: inst = 32'hc405664;
      17678: inst = 32'h8220000;
      17679: inst = 32'h10408000;
      17680: inst = 32'hc405665;
      17681: inst = 32'h8220000;
      17682: inst = 32'h10408000;
      17683: inst = 32'hc405666;
      17684: inst = 32'h8220000;
      17685: inst = 32'h10408000;
      17686: inst = 32'hc405667;
      17687: inst = 32'h8220000;
      17688: inst = 32'h10408000;
      17689: inst = 32'hc405668;
      17690: inst = 32'h8220000;
      17691: inst = 32'h10408000;
      17692: inst = 32'hc405669;
      17693: inst = 32'h8220000;
      17694: inst = 32'h10408000;
      17695: inst = 32'hc40566a;
      17696: inst = 32'h8220000;
      17697: inst = 32'h10408000;
      17698: inst = 32'hc40566b;
      17699: inst = 32'h8220000;
      17700: inst = 32'h10408000;
      17701: inst = 32'hc40566c;
      17702: inst = 32'h8220000;
      17703: inst = 32'h10408000;
      17704: inst = 32'hc40566d;
      17705: inst = 32'h8220000;
      17706: inst = 32'h10408000;
      17707: inst = 32'hc40566e;
      17708: inst = 32'h8220000;
      17709: inst = 32'h10408000;
      17710: inst = 32'hc40566f;
      17711: inst = 32'h8220000;
      17712: inst = 32'h10408000;
      17713: inst = 32'hc405670;
      17714: inst = 32'h8220000;
      17715: inst = 32'h10408000;
      17716: inst = 32'hc405671;
      17717: inst = 32'h8220000;
      17718: inst = 32'h10408000;
      17719: inst = 32'hc405672;
      17720: inst = 32'h8220000;
      17721: inst = 32'h10408000;
      17722: inst = 32'hc405673;
      17723: inst = 32'h8220000;
      17724: inst = 32'h10408000;
      17725: inst = 32'hc40568a;
      17726: inst = 32'h8220000;
      17727: inst = 32'h10408000;
      17728: inst = 32'hc40568b;
      17729: inst = 32'h8220000;
      17730: inst = 32'h10408000;
      17731: inst = 32'hc40568c;
      17732: inst = 32'h8220000;
      17733: inst = 32'h10408000;
      17734: inst = 32'hc40568d;
      17735: inst = 32'h8220000;
      17736: inst = 32'h10408000;
      17737: inst = 32'hc40568e;
      17738: inst = 32'h8220000;
      17739: inst = 32'h10408000;
      17740: inst = 32'hc40568f;
      17741: inst = 32'h8220000;
      17742: inst = 32'h10408000;
      17743: inst = 32'hc405690;
      17744: inst = 32'h8220000;
      17745: inst = 32'h10408000;
      17746: inst = 32'hc405691;
      17747: inst = 32'h8220000;
      17748: inst = 32'h10408000;
      17749: inst = 32'hc405692;
      17750: inst = 32'h8220000;
      17751: inst = 32'h10408000;
      17752: inst = 32'hc405693;
      17753: inst = 32'h8220000;
      17754: inst = 32'h10408000;
      17755: inst = 32'hc405694;
      17756: inst = 32'h8220000;
      17757: inst = 32'h10408000;
      17758: inst = 32'hc405695;
      17759: inst = 32'h8220000;
      17760: inst = 32'h10408000;
      17761: inst = 32'hc4056ac;
      17762: inst = 32'h8220000;
      17763: inst = 32'h10408000;
      17764: inst = 32'hc4056ad;
      17765: inst = 32'h8220000;
      17766: inst = 32'h10408000;
      17767: inst = 32'hc4056ae;
      17768: inst = 32'h8220000;
      17769: inst = 32'h10408000;
      17770: inst = 32'hc4056af;
      17771: inst = 32'h8220000;
      17772: inst = 32'h10408000;
      17773: inst = 32'hc4056b0;
      17774: inst = 32'h8220000;
      17775: inst = 32'h10408000;
      17776: inst = 32'hc4056b1;
      17777: inst = 32'h8220000;
      17778: inst = 32'h10408000;
      17779: inst = 32'hc4056b2;
      17780: inst = 32'h8220000;
      17781: inst = 32'h10408000;
      17782: inst = 32'hc4056b3;
      17783: inst = 32'h8220000;
      17784: inst = 32'h10408000;
      17785: inst = 32'hc4056b4;
      17786: inst = 32'h8220000;
      17787: inst = 32'h10408000;
      17788: inst = 32'hc4056b5;
      17789: inst = 32'h8220000;
      17790: inst = 32'h10408000;
      17791: inst = 32'hc4056b6;
      17792: inst = 32'h8220000;
      17793: inst = 32'h10408000;
      17794: inst = 32'hc4056b7;
      17795: inst = 32'h8220000;
      17796: inst = 32'h10408000;
      17797: inst = 32'hc4056b8;
      17798: inst = 32'h8220000;
      17799: inst = 32'h10408000;
      17800: inst = 32'hc4056b9;
      17801: inst = 32'h8220000;
      17802: inst = 32'h10408000;
      17803: inst = 32'hc4056ba;
      17804: inst = 32'h8220000;
      17805: inst = 32'h10408000;
      17806: inst = 32'hc4056bb;
      17807: inst = 32'h8220000;
      17808: inst = 32'h10408000;
      17809: inst = 32'hc4056bc;
      17810: inst = 32'h8220000;
      17811: inst = 32'h10408000;
      17812: inst = 32'hc4056bd;
      17813: inst = 32'h8220000;
      17814: inst = 32'h10408000;
      17815: inst = 32'hc4056be;
      17816: inst = 32'h8220000;
      17817: inst = 32'h10408000;
      17818: inst = 32'hc4056bf;
      17819: inst = 32'h8220000;
      17820: inst = 32'h10408000;
      17821: inst = 32'hc4056c0;
      17822: inst = 32'h8220000;
      17823: inst = 32'h10408000;
      17824: inst = 32'hc4056c1;
      17825: inst = 32'h8220000;
      17826: inst = 32'h10408000;
      17827: inst = 32'hc4056c2;
      17828: inst = 32'h8220000;
      17829: inst = 32'h10408000;
      17830: inst = 32'hc4056c3;
      17831: inst = 32'h8220000;
      17832: inst = 32'h10408000;
      17833: inst = 32'hc4056c4;
      17834: inst = 32'h8220000;
      17835: inst = 32'h10408000;
      17836: inst = 32'hc4056c5;
      17837: inst = 32'h8220000;
      17838: inst = 32'h10408000;
      17839: inst = 32'hc4056c6;
      17840: inst = 32'h8220000;
      17841: inst = 32'h10408000;
      17842: inst = 32'hc4056c7;
      17843: inst = 32'h8220000;
      17844: inst = 32'h10408000;
      17845: inst = 32'hc4056c8;
      17846: inst = 32'h8220000;
      17847: inst = 32'h10408000;
      17848: inst = 32'hc4056c9;
      17849: inst = 32'h8220000;
      17850: inst = 32'h10408000;
      17851: inst = 32'hc4056ca;
      17852: inst = 32'h8220000;
      17853: inst = 32'h10408000;
      17854: inst = 32'hc4056cb;
      17855: inst = 32'h8220000;
      17856: inst = 32'h10408000;
      17857: inst = 32'hc4056cc;
      17858: inst = 32'h8220000;
      17859: inst = 32'h10408000;
      17860: inst = 32'hc4056cd;
      17861: inst = 32'h8220000;
      17862: inst = 32'h10408000;
      17863: inst = 32'hc4056ce;
      17864: inst = 32'h8220000;
      17865: inst = 32'h10408000;
      17866: inst = 32'hc4056cf;
      17867: inst = 32'h8220000;
      17868: inst = 32'h10408000;
      17869: inst = 32'hc4056d0;
      17870: inst = 32'h8220000;
      17871: inst = 32'h10408000;
      17872: inst = 32'hc4056d1;
      17873: inst = 32'h8220000;
      17874: inst = 32'h10408000;
      17875: inst = 32'hc4056d2;
      17876: inst = 32'h8220000;
      17877: inst = 32'h10408000;
      17878: inst = 32'hc4056ea;
      17879: inst = 32'h8220000;
      17880: inst = 32'h10408000;
      17881: inst = 32'hc4056eb;
      17882: inst = 32'h8220000;
      17883: inst = 32'h10408000;
      17884: inst = 32'hc4056ec;
      17885: inst = 32'h8220000;
      17886: inst = 32'h10408000;
      17887: inst = 32'hc4056ed;
      17888: inst = 32'h8220000;
      17889: inst = 32'h10408000;
      17890: inst = 32'hc4056ee;
      17891: inst = 32'h8220000;
      17892: inst = 32'h10408000;
      17893: inst = 32'hc4056ef;
      17894: inst = 32'h8220000;
      17895: inst = 32'h10408000;
      17896: inst = 32'hc4056f0;
      17897: inst = 32'h8220000;
      17898: inst = 32'h10408000;
      17899: inst = 32'hc4056f1;
      17900: inst = 32'h8220000;
      17901: inst = 32'h10408000;
      17902: inst = 32'hc4056f2;
      17903: inst = 32'h8220000;
      17904: inst = 32'h10408000;
      17905: inst = 32'hc4056f3;
      17906: inst = 32'h8220000;
      17907: inst = 32'h10408000;
      17908: inst = 32'hc4056f4;
      17909: inst = 32'h8220000;
      17910: inst = 32'h10408000;
      17911: inst = 32'hc4056f5;
      17912: inst = 32'h8220000;
      17913: inst = 32'h10408000;
      17914: inst = 32'hc40570d;
      17915: inst = 32'h8220000;
      17916: inst = 32'h10408000;
      17917: inst = 32'hc40570e;
      17918: inst = 32'h8220000;
      17919: inst = 32'h10408000;
      17920: inst = 32'hc40570f;
      17921: inst = 32'h8220000;
      17922: inst = 32'h10408000;
      17923: inst = 32'hc405710;
      17924: inst = 32'h8220000;
      17925: inst = 32'h10408000;
      17926: inst = 32'hc405711;
      17927: inst = 32'h8220000;
      17928: inst = 32'h10408000;
      17929: inst = 32'hc405712;
      17930: inst = 32'h8220000;
      17931: inst = 32'h10408000;
      17932: inst = 32'hc405713;
      17933: inst = 32'h8220000;
      17934: inst = 32'h10408000;
      17935: inst = 32'hc405714;
      17936: inst = 32'h8220000;
      17937: inst = 32'h10408000;
      17938: inst = 32'hc405715;
      17939: inst = 32'h8220000;
      17940: inst = 32'h10408000;
      17941: inst = 32'hc405716;
      17942: inst = 32'h8220000;
      17943: inst = 32'h10408000;
      17944: inst = 32'hc405717;
      17945: inst = 32'h8220000;
      17946: inst = 32'h10408000;
      17947: inst = 32'hc405718;
      17948: inst = 32'h8220000;
      17949: inst = 32'h10408000;
      17950: inst = 32'hc405719;
      17951: inst = 32'h8220000;
      17952: inst = 32'h10408000;
      17953: inst = 32'hc40571a;
      17954: inst = 32'h8220000;
      17955: inst = 32'h10408000;
      17956: inst = 32'hc40571b;
      17957: inst = 32'h8220000;
      17958: inst = 32'h10408000;
      17959: inst = 32'hc40571c;
      17960: inst = 32'h8220000;
      17961: inst = 32'h10408000;
      17962: inst = 32'hc40571d;
      17963: inst = 32'h8220000;
      17964: inst = 32'h10408000;
      17965: inst = 32'hc40571e;
      17966: inst = 32'h8220000;
      17967: inst = 32'h10408000;
      17968: inst = 32'hc40571f;
      17969: inst = 32'h8220000;
      17970: inst = 32'h10408000;
      17971: inst = 32'hc405720;
      17972: inst = 32'h8220000;
      17973: inst = 32'h10408000;
      17974: inst = 32'hc405721;
      17975: inst = 32'h8220000;
      17976: inst = 32'h10408000;
      17977: inst = 32'hc405722;
      17978: inst = 32'h8220000;
      17979: inst = 32'h10408000;
      17980: inst = 32'hc405723;
      17981: inst = 32'h8220000;
      17982: inst = 32'h10408000;
      17983: inst = 32'hc405724;
      17984: inst = 32'h8220000;
      17985: inst = 32'h10408000;
      17986: inst = 32'hc405725;
      17987: inst = 32'h8220000;
      17988: inst = 32'h10408000;
      17989: inst = 32'hc405726;
      17990: inst = 32'h8220000;
      17991: inst = 32'h10408000;
      17992: inst = 32'hc405727;
      17993: inst = 32'h8220000;
      17994: inst = 32'h10408000;
      17995: inst = 32'hc405728;
      17996: inst = 32'h8220000;
      17997: inst = 32'h10408000;
      17998: inst = 32'hc405729;
      17999: inst = 32'h8220000;
      18000: inst = 32'h10408000;
      18001: inst = 32'hc40572a;
      18002: inst = 32'h8220000;
      18003: inst = 32'h10408000;
      18004: inst = 32'hc40572b;
      18005: inst = 32'h8220000;
      18006: inst = 32'h10408000;
      18007: inst = 32'hc40572c;
      18008: inst = 32'h8220000;
      18009: inst = 32'h10408000;
      18010: inst = 32'hc40572d;
      18011: inst = 32'h8220000;
      18012: inst = 32'h10408000;
      18013: inst = 32'hc40572e;
      18014: inst = 32'h8220000;
      18015: inst = 32'h10408000;
      18016: inst = 32'hc40572f;
      18017: inst = 32'h8220000;
      18018: inst = 32'h10408000;
      18019: inst = 32'hc405730;
      18020: inst = 32'h8220000;
      18021: inst = 32'h10408000;
      18022: inst = 32'hc405731;
      18023: inst = 32'h8220000;
      18024: inst = 32'h10408000;
      18025: inst = 32'hc40574a;
      18026: inst = 32'h8220000;
      18027: inst = 32'h10408000;
      18028: inst = 32'hc40574b;
      18029: inst = 32'h8220000;
      18030: inst = 32'h10408000;
      18031: inst = 32'hc40574c;
      18032: inst = 32'h8220000;
      18033: inst = 32'h10408000;
      18034: inst = 32'hc40574d;
      18035: inst = 32'h8220000;
      18036: inst = 32'h10408000;
      18037: inst = 32'hc40574e;
      18038: inst = 32'h8220000;
      18039: inst = 32'h10408000;
      18040: inst = 32'hc40574f;
      18041: inst = 32'h8220000;
      18042: inst = 32'h10408000;
      18043: inst = 32'hc405750;
      18044: inst = 32'h8220000;
      18045: inst = 32'h10408000;
      18046: inst = 32'hc405751;
      18047: inst = 32'h8220000;
      18048: inst = 32'h10408000;
      18049: inst = 32'hc405752;
      18050: inst = 32'h8220000;
      18051: inst = 32'h10408000;
      18052: inst = 32'hc405753;
      18053: inst = 32'h8220000;
      18054: inst = 32'h10408000;
      18055: inst = 32'hc405754;
      18056: inst = 32'h8220000;
      18057: inst = 32'h10408000;
      18058: inst = 32'hc405755;
      18059: inst = 32'h8220000;
      18060: inst = 32'h10408000;
      18061: inst = 32'hc40576e;
      18062: inst = 32'h8220000;
      18063: inst = 32'h10408000;
      18064: inst = 32'hc40576f;
      18065: inst = 32'h8220000;
      18066: inst = 32'h10408000;
      18067: inst = 32'hc405770;
      18068: inst = 32'h8220000;
      18069: inst = 32'h10408000;
      18070: inst = 32'hc405771;
      18071: inst = 32'h8220000;
      18072: inst = 32'h10408000;
      18073: inst = 32'hc405772;
      18074: inst = 32'h8220000;
      18075: inst = 32'h10408000;
      18076: inst = 32'hc405773;
      18077: inst = 32'h8220000;
      18078: inst = 32'h10408000;
      18079: inst = 32'hc405774;
      18080: inst = 32'h8220000;
      18081: inst = 32'h10408000;
      18082: inst = 32'hc405775;
      18083: inst = 32'h8220000;
      18084: inst = 32'h10408000;
      18085: inst = 32'hc405776;
      18086: inst = 32'h8220000;
      18087: inst = 32'h10408000;
      18088: inst = 32'hc405777;
      18089: inst = 32'h8220000;
      18090: inst = 32'h10408000;
      18091: inst = 32'hc405778;
      18092: inst = 32'h8220000;
      18093: inst = 32'h10408000;
      18094: inst = 32'hc405779;
      18095: inst = 32'h8220000;
      18096: inst = 32'h10408000;
      18097: inst = 32'hc40577a;
      18098: inst = 32'h8220000;
      18099: inst = 32'h10408000;
      18100: inst = 32'hc40577b;
      18101: inst = 32'h8220000;
      18102: inst = 32'h10408000;
      18103: inst = 32'hc40577c;
      18104: inst = 32'h8220000;
      18105: inst = 32'h10408000;
      18106: inst = 32'hc40577d;
      18107: inst = 32'h8220000;
      18108: inst = 32'h10408000;
      18109: inst = 32'hc40577e;
      18110: inst = 32'h8220000;
      18111: inst = 32'h10408000;
      18112: inst = 32'hc40577f;
      18113: inst = 32'h8220000;
      18114: inst = 32'h10408000;
      18115: inst = 32'hc405780;
      18116: inst = 32'h8220000;
      18117: inst = 32'h10408000;
      18118: inst = 32'hc405781;
      18119: inst = 32'h8220000;
      18120: inst = 32'h10408000;
      18121: inst = 32'hc405782;
      18122: inst = 32'h8220000;
      18123: inst = 32'h10408000;
      18124: inst = 32'hc405783;
      18125: inst = 32'h8220000;
      18126: inst = 32'h10408000;
      18127: inst = 32'hc405784;
      18128: inst = 32'h8220000;
      18129: inst = 32'h10408000;
      18130: inst = 32'hc405785;
      18131: inst = 32'h8220000;
      18132: inst = 32'h10408000;
      18133: inst = 32'hc405786;
      18134: inst = 32'h8220000;
      18135: inst = 32'h10408000;
      18136: inst = 32'hc405787;
      18137: inst = 32'h8220000;
      18138: inst = 32'h10408000;
      18139: inst = 32'hc405788;
      18140: inst = 32'h8220000;
      18141: inst = 32'h10408000;
      18142: inst = 32'hc405789;
      18143: inst = 32'h8220000;
      18144: inst = 32'h10408000;
      18145: inst = 32'hc40578a;
      18146: inst = 32'h8220000;
      18147: inst = 32'h10408000;
      18148: inst = 32'hc40578b;
      18149: inst = 32'h8220000;
      18150: inst = 32'h10408000;
      18151: inst = 32'hc40578c;
      18152: inst = 32'h8220000;
      18153: inst = 32'h10408000;
      18154: inst = 32'hc40578d;
      18155: inst = 32'h8220000;
      18156: inst = 32'h10408000;
      18157: inst = 32'hc40578e;
      18158: inst = 32'h8220000;
      18159: inst = 32'h10408000;
      18160: inst = 32'hc40578f;
      18161: inst = 32'h8220000;
      18162: inst = 32'h10408000;
      18163: inst = 32'hc405790;
      18164: inst = 32'h8220000;
      18165: inst = 32'h10408000;
      18166: inst = 32'hc405791;
      18167: inst = 32'h8220000;
      18168: inst = 32'h10408000;
      18169: inst = 32'hc4057aa;
      18170: inst = 32'h8220000;
      18171: inst = 32'h10408000;
      18172: inst = 32'hc4057ab;
      18173: inst = 32'h8220000;
      18174: inst = 32'h10408000;
      18175: inst = 32'hc4057ac;
      18176: inst = 32'h8220000;
      18177: inst = 32'h10408000;
      18178: inst = 32'hc4057ad;
      18179: inst = 32'h8220000;
      18180: inst = 32'h10408000;
      18181: inst = 32'hc4057ae;
      18182: inst = 32'h8220000;
      18183: inst = 32'h10408000;
      18184: inst = 32'hc4057af;
      18185: inst = 32'h8220000;
      18186: inst = 32'h10408000;
      18187: inst = 32'hc4057b0;
      18188: inst = 32'h8220000;
      18189: inst = 32'h10408000;
      18190: inst = 32'hc4057b1;
      18191: inst = 32'h8220000;
      18192: inst = 32'h10408000;
      18193: inst = 32'hc4057b2;
      18194: inst = 32'h8220000;
      18195: inst = 32'h10408000;
      18196: inst = 32'hc4057b3;
      18197: inst = 32'h8220000;
      18198: inst = 32'h10408000;
      18199: inst = 32'hc4057b4;
      18200: inst = 32'h8220000;
      18201: inst = 32'h10408000;
      18202: inst = 32'hc4057b5;
      18203: inst = 32'h8220000;
      18204: inst = 32'h10408000;
      18205: inst = 32'hc4057ce;
      18206: inst = 32'h8220000;
      18207: inst = 32'h10408000;
      18208: inst = 32'hc4057cf;
      18209: inst = 32'h8220000;
      18210: inst = 32'h10408000;
      18211: inst = 32'hc4057d0;
      18212: inst = 32'h8220000;
      18213: inst = 32'h10408000;
      18214: inst = 32'hc4057d1;
      18215: inst = 32'h8220000;
      18216: inst = 32'h10408000;
      18217: inst = 32'hc4057d2;
      18218: inst = 32'h8220000;
      18219: inst = 32'h10408000;
      18220: inst = 32'hc4057d3;
      18221: inst = 32'h8220000;
      18222: inst = 32'h10408000;
      18223: inst = 32'hc4057d4;
      18224: inst = 32'h8220000;
      18225: inst = 32'h10408000;
      18226: inst = 32'hc4057d5;
      18227: inst = 32'h8220000;
      18228: inst = 32'h10408000;
      18229: inst = 32'hc4057d6;
      18230: inst = 32'h8220000;
      18231: inst = 32'h10408000;
      18232: inst = 32'hc4057d7;
      18233: inst = 32'h8220000;
      18234: inst = 32'h10408000;
      18235: inst = 32'hc4057d8;
      18236: inst = 32'h8220000;
      18237: inst = 32'h10408000;
      18238: inst = 32'hc4057d9;
      18239: inst = 32'h8220000;
      18240: inst = 32'h10408000;
      18241: inst = 32'hc4057da;
      18242: inst = 32'h8220000;
      18243: inst = 32'h10408000;
      18244: inst = 32'hc4057db;
      18245: inst = 32'h8220000;
      18246: inst = 32'h10408000;
      18247: inst = 32'hc4057dc;
      18248: inst = 32'h8220000;
      18249: inst = 32'h10408000;
      18250: inst = 32'hc4057dd;
      18251: inst = 32'h8220000;
      18252: inst = 32'h10408000;
      18253: inst = 32'hc4057de;
      18254: inst = 32'h8220000;
      18255: inst = 32'h10408000;
      18256: inst = 32'hc4057df;
      18257: inst = 32'h8220000;
      18258: inst = 32'hc207bd0;
      18259: inst = 32'h10408000;
      18260: inst = 32'hc40531b;
      18261: inst = 32'h8220000;
      18262: inst = 32'h10408000;
      18263: inst = 32'hc405344;
      18264: inst = 32'h8220000;
      18265: inst = 32'hc207bcf;
      18266: inst = 32'h10408000;
      18267: inst = 32'hc405321;
      18268: inst = 32'h8220000;
      18269: inst = 32'h10408000;
      18270: inst = 32'hc40533e;
      18271: inst = 32'h8220000;
      18272: inst = 32'h10408000;
      18273: inst = 32'hc405381;
      18274: inst = 32'h8220000;
      18275: inst = 32'h10408000;
      18276: inst = 32'hc40539e;
      18277: inst = 32'h8220000;
      18278: inst = 32'h10408000;
      18279: inst = 32'hc4053e1;
      18280: inst = 32'h8220000;
      18281: inst = 32'h10408000;
      18282: inst = 32'hc4053fe;
      18283: inst = 32'h8220000;
      18284: inst = 32'h10408000;
      18285: inst = 32'hc405441;
      18286: inst = 32'h8220000;
      18287: inst = 32'h10408000;
      18288: inst = 32'hc405448;
      18289: inst = 32'h8220000;
      18290: inst = 32'h10408000;
      18291: inst = 32'hc405457;
      18292: inst = 32'h8220000;
      18293: inst = 32'h10408000;
      18294: inst = 32'hc40545e;
      18295: inst = 32'h8220000;
      18296: inst = 32'h10408000;
      18297: inst = 32'hc405501;
      18298: inst = 32'h8220000;
      18299: inst = 32'h10408000;
      18300: inst = 32'hc40551e;
      18301: inst = 32'h8220000;
      18302: inst = 32'h10408000;
      18303: inst = 32'hc405561;
      18304: inst = 32'h8220000;
      18305: inst = 32'h10408000;
      18306: inst = 32'hc40557e;
      18307: inst = 32'h8220000;
      18308: inst = 32'h10408000;
      18309: inst = 32'hc4055b9;
      18310: inst = 32'h8220000;
      18311: inst = 32'h10408000;
      18312: inst = 32'hc4055c1;
      18313: inst = 32'h8220000;
      18314: inst = 32'h10408000;
      18315: inst = 32'hc4055de;
      18316: inst = 32'h8220000;
      18317: inst = 32'h10408000;
      18318: inst = 32'hc4055e6;
      18319: inst = 32'h8220000;
      18320: inst = 32'h10408000;
      18321: inst = 32'hc40561e;
      18322: inst = 32'h8220000;
      18323: inst = 32'h10408000;
      18324: inst = 32'hc405621;
      18325: inst = 32'h8220000;
      18326: inst = 32'h10408000;
      18327: inst = 32'hc40563e;
      18328: inst = 32'h8220000;
      18329: inst = 32'h10408000;
      18330: inst = 32'hc405641;
      18331: inst = 32'h8220000;
      18332: inst = 32'h10408000;
      18333: inst = 32'hc405681;
      18334: inst = 32'h8220000;
      18335: inst = 32'h10408000;
      18336: inst = 32'hc405698;
      18337: inst = 32'h8220000;
      18338: inst = 32'h10408000;
      18339: inst = 32'hc40569e;
      18340: inst = 32'h8220000;
      18341: inst = 32'h10408000;
      18342: inst = 32'hc4056e1;
      18343: inst = 32'h8220000;
      18344: inst = 32'h10408000;
      18345: inst = 32'hc4056fe;
      18346: inst = 32'h8220000;
      18347: inst = 32'hc207390;
      18348: inst = 32'h10408000;
      18349: inst = 32'hc40537a;
      18350: inst = 32'h8220000;
      18351: inst = 32'h10408000;
      18352: inst = 32'hc4053a5;
      18353: inst = 32'h8220000;
      18354: inst = 32'hc2052aa;
      18355: inst = 32'h10408000;
      18356: inst = 32'hc405389;
      18357: inst = 32'h8220000;
      18358: inst = 32'h10408000;
      18359: inst = 32'hc405396;
      18360: inst = 32'h8220000;
      18361: inst = 32'h10408000;
      18362: inst = 32'hc4054fb;
      18363: inst = 32'h8220000;
      18364: inst = 32'h10408000;
      18365: inst = 32'hc405503;
      18366: inst = 32'h8220000;
      18367: inst = 32'h10408000;
      18368: inst = 32'hc40551c;
      18369: inst = 32'h8220000;
      18370: inst = 32'h10408000;
      18371: inst = 32'hc405524;
      18372: inst = 32'h8220000;
      18373: inst = 32'h10408000;
      18374: inst = 32'hc4055c8;
      18375: inst = 32'h8220000;
      18376: inst = 32'h10408000;
      18377: inst = 32'hc4055d7;
      18378: inst = 32'h8220000;
      18379: inst = 32'h10408000;
      18380: inst = 32'hc405619;
      18381: inst = 32'h8220000;
      18382: inst = 32'h10408000;
      18383: inst = 32'hc405622;
      18384: inst = 32'h8220000;
      18385: inst = 32'h10408000;
      18386: inst = 32'hc40563d;
      18387: inst = 32'h8220000;
      18388: inst = 32'h10408000;
      18389: inst = 32'hc405646;
      18390: inst = 32'h8220000;
      18391: inst = 32'hc206b70;
      18392: inst = 32'h10408000;
      18393: inst = 32'hc4053d9;
      18394: inst = 32'h8220000;
      18395: inst = 32'h10408000;
      18396: inst = 32'hc405406;
      18397: inst = 32'h8220000;
      18398: inst = 32'h10408000;
      18399: inst = 32'hc405556;
      18400: inst = 32'h8220000;
      18401: inst = 32'h10408000;
      18402: inst = 32'hc405589;
      18403: inst = 32'h8220000;
      18404: inst = 32'h10408000;
      18405: inst = 32'hc4055b5;
      18406: inst = 32'h8220000;
      18407: inst = 32'h10408000;
      18408: inst = 32'hc4055ea;
      18409: inst = 32'h8220000;
      18410: inst = 32'h10408000;
      18411: inst = 32'hc405732;
      18412: inst = 32'h8220000;
      18413: inst = 32'h10408000;
      18414: inst = 32'hc40576d;
      18415: inst = 32'h8220000;
      18416: inst = 32'hc20736e;
      18417: inst = 32'h10408000;
      18418: inst = 32'hc4053e0;
      18419: inst = 32'h8220000;
      18420: inst = 32'h10408000;
      18421: inst = 32'hc4053ff;
      18422: inst = 32'h8220000;
      18423: inst = 32'hc205aaa;
      18424: inst = 32'h10408000;
      18425: inst = 32'hc4053e4;
      18426: inst = 32'h8220000;
      18427: inst = 32'h10408000;
      18428: inst = 32'hc4053fb;
      18429: inst = 32'h8220000;
      18430: inst = 32'hc208431;
      18431: inst = 32'h10408000;
      18432: inst = 32'hc4053e8;
      18433: inst = 32'h8220000;
      18434: inst = 32'h10408000;
      18435: inst = 32'hc4053f7;
      18436: inst = 32'h8220000;
      18437: inst = 32'h10408000;
      18438: inst = 32'hc405439;
      18439: inst = 32'h8220000;
      18440: inst = 32'h10408000;
      18441: inst = 32'hc405466;
      18442: inst = 32'h8220000;
      18443: inst = 32'h10408000;
      18444: inst = 32'hc4055b6;
      18445: inst = 32'h8220000;
      18446: inst = 32'h10408000;
      18447: inst = 32'hc4055e9;
      18448: inst = 32'h8220000;
      18449: inst = 32'h10408000;
      18450: inst = 32'hc405733;
      18451: inst = 32'h8220000;
      18452: inst = 32'h10408000;
      18453: inst = 32'hc40576c;
      18454: inst = 32'h8220000;
      18455: inst = 32'hc206b4d;
      18456: inst = 32'h10408000;
      18457: inst = 32'hc40543c;
      18458: inst = 32'h8220000;
      18459: inst = 32'h10408000;
      18460: inst = 32'hc405444;
      18461: inst = 32'h8220000;
      18462: inst = 32'h10408000;
      18463: inst = 32'hc40545b;
      18464: inst = 32'h8220000;
      18465: inst = 32'h10408000;
      18466: inst = 32'hc405463;
      18467: inst = 32'h8220000;
      18468: inst = 32'h10408000;
      18469: inst = 32'hc405563;
      18470: inst = 32'h8220000;
      18471: inst = 32'h10408000;
      18472: inst = 32'hc40557c;
      18473: inst = 32'h8220000;
      18474: inst = 32'h10408000;
      18475: inst = 32'hc405682;
      18476: inst = 32'h8220000;
      18477: inst = 32'h10408000;
      18478: inst = 32'hc40569d;
      18479: inst = 32'h8220000;
      18480: inst = 32'hc208430;
      18481: inst = 32'h10408000;
      18482: inst = 32'hc405440;
      18483: inst = 32'h8220000;
      18484: inst = 32'h10408000;
      18485: inst = 32'hc40545f;
      18486: inst = 32'h8220000;
      18487: inst = 32'hc207bf1;
      18488: inst = 32'h10408000;
      18489: inst = 32'hc405498;
      18490: inst = 32'h8220000;
      18491: inst = 32'h10408000;
      18492: inst = 32'hc4054c7;
      18493: inst = 32'h8220000;
      18494: inst = 32'h10408000;
      18495: inst = 32'hc405615;
      18496: inst = 32'h8220000;
      18497: inst = 32'h10408000;
      18498: inst = 32'hc40564a;
      18499: inst = 32'h8220000;
      18500: inst = 32'hc207bef;
      18501: inst = 32'h10408000;
      18502: inst = 32'hc40549b;
      18503: inst = 32'h8220000;
      18504: inst = 32'h10408000;
      18505: inst = 32'hc4054c4;
      18506: inst = 32'h8220000;
      18507: inst = 32'h10408000;
      18508: inst = 32'hc405687;
      18509: inst = 32'h8220000;
      18510: inst = 32'h10408000;
      18511: inst = 32'hc4056e2;
      18512: inst = 32'h8220000;
      18513: inst = 32'h10408000;
      18514: inst = 32'hc4056fd;
      18515: inst = 32'h8220000;
      18516: inst = 32'hc205aeb;
      18517: inst = 32'h10408000;
      18518: inst = 32'hc40549f;
      18519: inst = 32'h8220000;
      18520: inst = 32'h10408000;
      18521: inst = 32'hc4054c0;
      18522: inst = 32'h8220000;
      18523: inst = 32'hc206b6e;
      18524: inst = 32'h10408000;
      18525: inst = 32'hc4054a8;
      18526: inst = 32'h8220000;
      18527: inst = 32'h10408000;
      18528: inst = 32'hc4054b7;
      18529: inst = 32'h8220000;
      18530: inst = 32'h10408000;
      18531: inst = 32'hc4056e7;
      18532: inst = 32'h8220000;
      18533: inst = 32'h10408000;
      18534: inst = 32'hc4056f8;
      18535: inst = 32'h8220000;
      18536: inst = 32'hc2073b0;
      18537: inst = 32'h10408000;
      18538: inst = 32'hc4054f7;
      18539: inst = 32'h8220000;
      18540: inst = 32'h10408000;
      18541: inst = 32'hc405528;
      18542: inst = 32'h8220000;
      18543: inst = 32'h10408000;
      18544: inst = 32'hc405674;
      18545: inst = 32'h8220000;
      18546: inst = 32'h10408000;
      18547: inst = 32'hc4056ab;
      18548: inst = 32'h8220000;
      18549: inst = 32'hc2073ae;
      18550: inst = 32'h10408000;
      18551: inst = 32'hc4054ff;
      18552: inst = 32'h8220000;
      18553: inst = 32'h10408000;
      18554: inst = 32'hc405520;
      18555: inst = 32'h8220000;
      18556: inst = 32'hc20632d;
      18557: inst = 32'h10408000;
      18558: inst = 32'hc405508;
      18559: inst = 32'h8220000;
      18560: inst = 32'h10408000;
      18561: inst = 32'hc405517;
      18562: inst = 32'h8220000;
      18563: inst = 32'h10408000;
      18564: inst = 32'hc405747;
      18565: inst = 32'h8220000;
      18566: inst = 32'h10408000;
      18567: inst = 32'hc405758;
      18568: inst = 32'h8220000;
      18569: inst = 32'hc206b2d;
      18570: inst = 32'h10408000;
      18571: inst = 32'hc40555a;
      18572: inst = 32'h8220000;
      18573: inst = 32'h10408000;
      18574: inst = 32'hc405585;
      18575: inst = 32'h8220000;
      18576: inst = 32'hc20630c;
      18577: inst = 32'h10408000;
      18578: inst = 32'hc4055be;
      18579: inst = 32'h8220000;
      18580: inst = 32'h10408000;
      18581: inst = 32'hc4055e1;
      18582: inst = 32'h8220000;
      18583: inst = 32'h10408000;
      18584: inst = 32'hc405678;
      18585: inst = 32'h8220000;
      18586: inst = 32'hc20632c;
      18587: inst = 32'h10408000;
      18588: inst = 32'hc4056a7;
      18589: inst = 32'h8220000;
      18590: inst = 32'hc206b90;
      18591: inst = 32'h10408000;
      18592: inst = 32'hc4056d3;
      18593: inst = 32'h8220000;
      18594: inst = 32'h10408000;
      18595: inst = 32'hc40570c;
      18596: inst = 32'h8220000;
      18597: inst = 32'hc207c11;
      18598: inst = 32'h10408000;
      18599: inst = 32'hc405792;
      18600: inst = 32'h8220000;
      18601: inst = 32'h10408000;
      18602: inst = 32'hc4057cd;
      18603: inst = 32'h8220000;
      18604: inst = 32'h58000000;
      18605: inst = 32'hc20ea25;
      18606: inst = 32'h10408000;
      18607: inst = 32'hc40464d;
      18608: inst = 32'h8220000;
      18609: inst = 32'h10408000;
      18610: inst = 32'hc40464e;
      18611: inst = 32'h8220000;
      18612: inst = 32'h10408000;
      18613: inst = 32'hc40464f;
      18614: inst = 32'h8220000;
      18615: inst = 32'h10408000;
      18616: inst = 32'hc404650;
      18617: inst = 32'h8220000;
      18618: inst = 32'h10408000;
      18619: inst = 32'hc404651;
      18620: inst = 32'h8220000;
      18621: inst = 32'h10408000;
      18622: inst = 32'hc404652;
      18623: inst = 32'h8220000;
      18624: inst = 32'h10408000;
      18625: inst = 32'hc404653;
      18626: inst = 32'h8220000;
      18627: inst = 32'h10408000;
      18628: inst = 32'hc404654;
      18629: inst = 32'h8220000;
      18630: inst = 32'h10408000;
      18631: inst = 32'hc404655;
      18632: inst = 32'h8220000;
      18633: inst = 32'h10408000;
      18634: inst = 32'hc404659;
      18635: inst = 32'h8220000;
      18636: inst = 32'h10408000;
      18637: inst = 32'hc40465a;
      18638: inst = 32'h8220000;
      18639: inst = 32'h10408000;
      18640: inst = 32'hc40465b;
      18641: inst = 32'h8220000;
      18642: inst = 32'h10408000;
      18643: inst = 32'hc40465c;
      18644: inst = 32'h8220000;
      18645: inst = 32'h10408000;
      18646: inst = 32'hc40465d;
      18647: inst = 32'h8220000;
      18648: inst = 32'h10408000;
      18649: inst = 32'hc40465e;
      18650: inst = 32'h8220000;
      18651: inst = 32'h10408000;
      18652: inst = 32'hc40465f;
      18653: inst = 32'h8220000;
      18654: inst = 32'h10408000;
      18655: inst = 32'hc404660;
      18656: inst = 32'h8220000;
      18657: inst = 32'h10408000;
      18658: inst = 32'hc404661;
      18659: inst = 32'h8220000;
      18660: inst = 32'h10408000;
      18661: inst = 32'hc404663;
      18662: inst = 32'h8220000;
      18663: inst = 32'h10408000;
      18664: inst = 32'hc404664;
      18665: inst = 32'h8220000;
      18666: inst = 32'h10408000;
      18667: inst = 32'hc404665;
      18668: inst = 32'h8220000;
      18669: inst = 32'h10408000;
      18670: inst = 32'hc404666;
      18671: inst = 32'h8220000;
      18672: inst = 32'h10408000;
      18673: inst = 32'hc404667;
      18674: inst = 32'h8220000;
      18675: inst = 32'h10408000;
      18676: inst = 32'hc404668;
      18677: inst = 32'h8220000;
      18678: inst = 32'h10408000;
      18679: inst = 32'hc404669;
      18680: inst = 32'h8220000;
      18681: inst = 32'h10408000;
      18682: inst = 32'hc40466a;
      18683: inst = 32'h8220000;
      18684: inst = 32'h10408000;
      18685: inst = 32'hc40466b;
      18686: inst = 32'h8220000;
      18687: inst = 32'h10408000;
      18688: inst = 32'hc404671;
      18689: inst = 32'h8220000;
      18690: inst = 32'h10408000;
      18691: inst = 32'hc404672;
      18692: inst = 32'h8220000;
      18693: inst = 32'h10408000;
      18694: inst = 32'hc404673;
      18695: inst = 32'h8220000;
      18696: inst = 32'h10408000;
      18697: inst = 32'hc404674;
      18698: inst = 32'h8220000;
      18699: inst = 32'h10408000;
      18700: inst = 32'hc404675;
      18701: inst = 32'h8220000;
      18702: inst = 32'h10408000;
      18703: inst = 32'hc404676;
      18704: inst = 32'h8220000;
      18705: inst = 32'h10408000;
      18706: inst = 32'hc404677;
      18707: inst = 32'h8220000;
      18708: inst = 32'h10408000;
      18709: inst = 32'hc404678;
      18710: inst = 32'h8220000;
      18711: inst = 32'h10408000;
      18712: inst = 32'hc404679;
      18713: inst = 32'h8220000;
      18714: inst = 32'h10408000;
      18715: inst = 32'hc40467c;
      18716: inst = 32'h8220000;
      18717: inst = 32'h10408000;
      18718: inst = 32'hc40467d;
      18719: inst = 32'h8220000;
      18720: inst = 32'h10408000;
      18721: inst = 32'hc40467e;
      18722: inst = 32'h8220000;
      18723: inst = 32'h10408000;
      18724: inst = 32'hc40467f;
      18725: inst = 32'h8220000;
      18726: inst = 32'h10408000;
      18727: inst = 32'hc404680;
      18728: inst = 32'h8220000;
      18729: inst = 32'h10408000;
      18730: inst = 32'hc404681;
      18731: inst = 32'h8220000;
      18732: inst = 32'h10408000;
      18733: inst = 32'hc404682;
      18734: inst = 32'h8220000;
      18735: inst = 32'h10408000;
      18736: inst = 32'hc404683;
      18737: inst = 32'h8220000;
      18738: inst = 32'h10408000;
      18739: inst = 32'hc404684;
      18740: inst = 32'h8220000;
      18741: inst = 32'h10408000;
      18742: inst = 32'hc404685;
      18743: inst = 32'h8220000;
      18744: inst = 32'h10408000;
      18745: inst = 32'hc40468b;
      18746: inst = 32'h8220000;
      18747: inst = 32'h10408000;
      18748: inst = 32'hc40468c;
      18749: inst = 32'h8220000;
      18750: inst = 32'h10408000;
      18751: inst = 32'hc40468d;
      18752: inst = 32'h8220000;
      18753: inst = 32'h10408000;
      18754: inst = 32'hc40468e;
      18755: inst = 32'h8220000;
      18756: inst = 32'h10408000;
      18757: inst = 32'hc40468f;
      18758: inst = 32'h8220000;
      18759: inst = 32'h10408000;
      18760: inst = 32'hc404690;
      18761: inst = 32'h8220000;
      18762: inst = 32'h10408000;
      18763: inst = 32'hc404691;
      18764: inst = 32'h8220000;
      18765: inst = 32'h10408000;
      18766: inst = 32'hc404692;
      18767: inst = 32'h8220000;
      18768: inst = 32'h10408000;
      18769: inst = 32'hc404693;
      18770: inst = 32'h8220000;
      18771: inst = 32'h10408000;
      18772: inst = 32'hc4046ac;
      18773: inst = 32'h8220000;
      18774: inst = 32'h10408000;
      18775: inst = 32'hc4046ad;
      18776: inst = 32'h8220000;
      18777: inst = 32'h10408000;
      18778: inst = 32'hc4046ae;
      18779: inst = 32'h8220000;
      18780: inst = 32'h10408000;
      18781: inst = 32'hc4046af;
      18782: inst = 32'h8220000;
      18783: inst = 32'h10408000;
      18784: inst = 32'hc4046b0;
      18785: inst = 32'h8220000;
      18786: inst = 32'h10408000;
      18787: inst = 32'hc4046b1;
      18788: inst = 32'h8220000;
      18789: inst = 32'h10408000;
      18790: inst = 32'hc4046b2;
      18791: inst = 32'h8220000;
      18792: inst = 32'h10408000;
      18793: inst = 32'hc4046b3;
      18794: inst = 32'h8220000;
      18795: inst = 32'h10408000;
      18796: inst = 32'hc4046b4;
      18797: inst = 32'h8220000;
      18798: inst = 32'h10408000;
      18799: inst = 32'hc4046b5;
      18800: inst = 32'h8220000;
      18801: inst = 32'h10408000;
      18802: inst = 32'hc4046b8;
      18803: inst = 32'h8220000;
      18804: inst = 32'h10408000;
      18805: inst = 32'hc4046b9;
      18806: inst = 32'h8220000;
      18807: inst = 32'h10408000;
      18808: inst = 32'hc4046ba;
      18809: inst = 32'h8220000;
      18810: inst = 32'h10408000;
      18811: inst = 32'hc4046bb;
      18812: inst = 32'h8220000;
      18813: inst = 32'h10408000;
      18814: inst = 32'hc4046bc;
      18815: inst = 32'h8220000;
      18816: inst = 32'h10408000;
      18817: inst = 32'hc4046bd;
      18818: inst = 32'h8220000;
      18819: inst = 32'h10408000;
      18820: inst = 32'hc4046be;
      18821: inst = 32'h8220000;
      18822: inst = 32'h10408000;
      18823: inst = 32'hc4046bf;
      18824: inst = 32'h8220000;
      18825: inst = 32'h10408000;
      18826: inst = 32'hc4046c0;
      18827: inst = 32'h8220000;
      18828: inst = 32'h10408000;
      18829: inst = 32'hc4046c1;
      18830: inst = 32'h8220000;
      18831: inst = 32'h10408000;
      18832: inst = 32'hc4046c3;
      18833: inst = 32'h8220000;
      18834: inst = 32'h10408000;
      18835: inst = 32'hc4046c4;
      18836: inst = 32'h8220000;
      18837: inst = 32'h10408000;
      18838: inst = 32'hc4046c5;
      18839: inst = 32'h8220000;
      18840: inst = 32'h10408000;
      18841: inst = 32'hc4046c6;
      18842: inst = 32'h8220000;
      18843: inst = 32'h10408000;
      18844: inst = 32'hc4046c7;
      18845: inst = 32'h8220000;
      18846: inst = 32'h10408000;
      18847: inst = 32'hc4046c8;
      18848: inst = 32'h8220000;
      18849: inst = 32'h10408000;
      18850: inst = 32'hc4046c9;
      18851: inst = 32'h8220000;
      18852: inst = 32'h10408000;
      18853: inst = 32'hc4046ca;
      18854: inst = 32'h8220000;
      18855: inst = 32'h10408000;
      18856: inst = 32'hc4046cb;
      18857: inst = 32'h8220000;
      18858: inst = 32'h10408000;
      18859: inst = 32'hc4046d0;
      18860: inst = 32'h8220000;
      18861: inst = 32'h10408000;
      18862: inst = 32'hc4046d1;
      18863: inst = 32'h8220000;
      18864: inst = 32'h10408000;
      18865: inst = 32'hc4046d2;
      18866: inst = 32'h8220000;
      18867: inst = 32'h10408000;
      18868: inst = 32'hc4046d3;
      18869: inst = 32'h8220000;
      18870: inst = 32'h10408000;
      18871: inst = 32'hc4046d4;
      18872: inst = 32'h8220000;
      18873: inst = 32'h10408000;
      18874: inst = 32'hc4046d5;
      18875: inst = 32'h8220000;
      18876: inst = 32'h10408000;
      18877: inst = 32'hc4046d6;
      18878: inst = 32'h8220000;
      18879: inst = 32'h10408000;
      18880: inst = 32'hc4046d7;
      18881: inst = 32'h8220000;
      18882: inst = 32'h10408000;
      18883: inst = 32'hc4046d8;
      18884: inst = 32'h8220000;
      18885: inst = 32'h10408000;
      18886: inst = 32'hc4046da;
      18887: inst = 32'h8220000;
      18888: inst = 32'h10408000;
      18889: inst = 32'hc4046dc;
      18890: inst = 32'h8220000;
      18891: inst = 32'h10408000;
      18892: inst = 32'hc4046dd;
      18893: inst = 32'h8220000;
      18894: inst = 32'h10408000;
      18895: inst = 32'hc4046de;
      18896: inst = 32'h8220000;
      18897: inst = 32'h10408000;
      18898: inst = 32'hc4046df;
      18899: inst = 32'h8220000;
      18900: inst = 32'h10408000;
      18901: inst = 32'hc4046e0;
      18902: inst = 32'h8220000;
      18903: inst = 32'h10408000;
      18904: inst = 32'hc4046e1;
      18905: inst = 32'h8220000;
      18906: inst = 32'h10408000;
      18907: inst = 32'hc4046e2;
      18908: inst = 32'h8220000;
      18909: inst = 32'h10408000;
      18910: inst = 32'hc4046e3;
      18911: inst = 32'h8220000;
      18912: inst = 32'h10408000;
      18913: inst = 32'hc4046e4;
      18914: inst = 32'h8220000;
      18915: inst = 32'h10408000;
      18916: inst = 32'hc4046e5;
      18917: inst = 32'h8220000;
      18918: inst = 32'h10408000;
      18919: inst = 32'hc4046ea;
      18920: inst = 32'h8220000;
      18921: inst = 32'h10408000;
      18922: inst = 32'hc4046eb;
      18923: inst = 32'h8220000;
      18924: inst = 32'h10408000;
      18925: inst = 32'hc4046ec;
      18926: inst = 32'h8220000;
      18927: inst = 32'h10408000;
      18928: inst = 32'hc4046ed;
      18929: inst = 32'h8220000;
      18930: inst = 32'h10408000;
      18931: inst = 32'hc4046ee;
      18932: inst = 32'h8220000;
      18933: inst = 32'h10408000;
      18934: inst = 32'hc4046ef;
      18935: inst = 32'h8220000;
      18936: inst = 32'h10408000;
      18937: inst = 32'hc4046f0;
      18938: inst = 32'h8220000;
      18939: inst = 32'h10408000;
      18940: inst = 32'hc4046f1;
      18941: inst = 32'h8220000;
      18942: inst = 32'h10408000;
      18943: inst = 32'hc4046f2;
      18944: inst = 32'h8220000;
      18945: inst = 32'h10408000;
      18946: inst = 32'hc4046f3;
      18947: inst = 32'h8220000;
      18948: inst = 32'h10408000;
      18949: inst = 32'hc40470b;
      18950: inst = 32'h8220000;
      18951: inst = 32'h10408000;
      18952: inst = 32'hc40470c;
      18953: inst = 32'h8220000;
      18954: inst = 32'h10408000;
      18955: inst = 32'hc40470d;
      18956: inst = 32'h8220000;
      18957: inst = 32'h10408000;
      18958: inst = 32'hc404717;
      18959: inst = 32'h8220000;
      18960: inst = 32'h10408000;
      18961: inst = 32'hc404718;
      18962: inst = 32'h8220000;
      18963: inst = 32'h10408000;
      18964: inst = 32'hc404719;
      18965: inst = 32'h8220000;
      18966: inst = 32'h10408000;
      18967: inst = 32'hc404728;
      18968: inst = 32'h8220000;
      18969: inst = 32'h10408000;
      18970: inst = 32'hc404729;
      18971: inst = 32'h8220000;
      18972: inst = 32'h10408000;
      18973: inst = 32'hc40472a;
      18974: inst = 32'h8220000;
      18975: inst = 32'h10408000;
      18976: inst = 32'hc40472b;
      18977: inst = 32'h8220000;
      18978: inst = 32'h10408000;
      18979: inst = 32'hc404730;
      18980: inst = 32'h8220000;
      18981: inst = 32'h10408000;
      18982: inst = 32'hc404731;
      18983: inst = 32'h8220000;
      18984: inst = 32'h10408000;
      18985: inst = 32'hc404735;
      18986: inst = 32'h8220000;
      18987: inst = 32'h10408000;
      18988: inst = 32'hc404736;
      18989: inst = 32'h8220000;
      18990: inst = 32'h10408000;
      18991: inst = 32'hc404737;
      18992: inst = 32'h8220000;
      18993: inst = 32'h10408000;
      18994: inst = 32'hc404739;
      18995: inst = 32'h8220000;
      18996: inst = 32'h10408000;
      18997: inst = 32'hc40473a;
      18998: inst = 32'h8220000;
      18999: inst = 32'h10408000;
      19000: inst = 32'hc404742;
      19001: inst = 32'h8220000;
      19002: inst = 32'h10408000;
      19003: inst = 32'hc404743;
      19004: inst = 32'h8220000;
      19005: inst = 32'h10408000;
      19006: inst = 32'hc404744;
      19007: inst = 32'h8220000;
      19008: inst = 32'h10408000;
      19009: inst = 32'hc404745;
      19010: inst = 32'h8220000;
      19011: inst = 32'h10408000;
      19012: inst = 32'hc404749;
      19013: inst = 32'h8220000;
      19014: inst = 32'h10408000;
      19015: inst = 32'hc40474a;
      19016: inst = 32'h8220000;
      19017: inst = 32'h10408000;
      19018: inst = 32'hc40474b;
      19019: inst = 32'h8220000;
      19020: inst = 32'h10408000;
      19021: inst = 32'hc40476b;
      19022: inst = 32'h8220000;
      19023: inst = 32'h10408000;
      19024: inst = 32'hc40476c;
      19025: inst = 32'h8220000;
      19026: inst = 32'h10408000;
      19027: inst = 32'hc404777;
      19028: inst = 32'h8220000;
      19029: inst = 32'h10408000;
      19030: inst = 32'hc404778;
      19031: inst = 32'h8220000;
      19032: inst = 32'h10408000;
      19033: inst = 32'hc404788;
      19034: inst = 32'h8220000;
      19035: inst = 32'h10408000;
      19036: inst = 32'hc404789;
      19037: inst = 32'h8220000;
      19038: inst = 32'h10408000;
      19039: inst = 32'hc40478a;
      19040: inst = 32'h8220000;
      19041: inst = 32'h10408000;
      19042: inst = 32'hc404790;
      19043: inst = 32'h8220000;
      19044: inst = 32'h10408000;
      19045: inst = 32'hc404791;
      19046: inst = 32'h8220000;
      19047: inst = 32'h10408000;
      19048: inst = 32'hc404795;
      19049: inst = 32'h8220000;
      19050: inst = 32'h10408000;
      19051: inst = 32'hc404799;
      19052: inst = 32'h8220000;
      19053: inst = 32'h10408000;
      19054: inst = 32'hc40479a;
      19055: inst = 32'h8220000;
      19056: inst = 32'h10408000;
      19057: inst = 32'hc4047a2;
      19058: inst = 32'h8220000;
      19059: inst = 32'h10408000;
      19060: inst = 32'hc4047a3;
      19061: inst = 32'h8220000;
      19062: inst = 32'h10408000;
      19063: inst = 32'hc4047a4;
      19064: inst = 32'h8220000;
      19065: inst = 32'h10408000;
      19066: inst = 32'hc4047a9;
      19067: inst = 32'h8220000;
      19068: inst = 32'h10408000;
      19069: inst = 32'hc4047aa;
      19070: inst = 32'h8220000;
      19071: inst = 32'h10408000;
      19072: inst = 32'hc4047cb;
      19073: inst = 32'h8220000;
      19074: inst = 32'h10408000;
      19075: inst = 32'hc4047cc;
      19076: inst = 32'h8220000;
      19077: inst = 32'h10408000;
      19078: inst = 32'hc4047ce;
      19079: inst = 32'h8220000;
      19080: inst = 32'h10408000;
      19081: inst = 32'hc4047cf;
      19082: inst = 32'h8220000;
      19083: inst = 32'h10408000;
      19084: inst = 32'hc4047d0;
      19085: inst = 32'h8220000;
      19086: inst = 32'h10408000;
      19087: inst = 32'hc4047d1;
      19088: inst = 32'h8220000;
      19089: inst = 32'h10408000;
      19090: inst = 32'hc4047d2;
      19091: inst = 32'h8220000;
      19092: inst = 32'h10408000;
      19093: inst = 32'hc4047d7;
      19094: inst = 32'h8220000;
      19095: inst = 32'h10408000;
      19096: inst = 32'hc4047d8;
      19097: inst = 32'h8220000;
      19098: inst = 32'h10408000;
      19099: inst = 32'hc4047da;
      19100: inst = 32'h8220000;
      19101: inst = 32'h10408000;
      19102: inst = 32'hc4047db;
      19103: inst = 32'h8220000;
      19104: inst = 32'h10408000;
      19105: inst = 32'hc4047dc;
      19106: inst = 32'h8220000;
      19107: inst = 32'h10408000;
      19108: inst = 32'hc4047dd;
      19109: inst = 32'h8220000;
      19110: inst = 32'h10408000;
      19111: inst = 32'hc4047de;
      19112: inst = 32'h8220000;
      19113: inst = 32'h10408000;
      19114: inst = 32'hc4047e7;
      19115: inst = 32'h8220000;
      19116: inst = 32'h10408000;
      19117: inst = 32'hc4047e8;
      19118: inst = 32'h8220000;
      19119: inst = 32'h10408000;
      19120: inst = 32'hc4047e9;
      19121: inst = 32'h8220000;
      19122: inst = 32'h10408000;
      19123: inst = 32'hc4047f0;
      19124: inst = 32'h8220000;
      19125: inst = 32'h10408000;
      19126: inst = 32'hc4047f1;
      19127: inst = 32'h8220000;
      19128: inst = 32'h10408000;
      19129: inst = 32'hc4047f9;
      19130: inst = 32'h8220000;
      19131: inst = 32'h10408000;
      19132: inst = 32'hc4047fa;
      19133: inst = 32'h8220000;
      19134: inst = 32'h10408000;
      19135: inst = 32'hc404800;
      19136: inst = 32'h8220000;
      19137: inst = 32'h10408000;
      19138: inst = 32'hc404801;
      19139: inst = 32'h8220000;
      19140: inst = 32'h10408000;
      19141: inst = 32'hc404802;
      19142: inst = 32'h8220000;
      19143: inst = 32'h10408000;
      19144: inst = 32'hc404803;
      19145: inst = 32'h8220000;
      19146: inst = 32'h10408000;
      19147: inst = 32'hc404809;
      19148: inst = 32'h8220000;
      19149: inst = 32'h10408000;
      19150: inst = 32'hc40480a;
      19151: inst = 32'h8220000;
      19152: inst = 32'h10408000;
      19153: inst = 32'hc40480c;
      19154: inst = 32'h8220000;
      19155: inst = 32'h10408000;
      19156: inst = 32'hc40480d;
      19157: inst = 32'h8220000;
      19158: inst = 32'h10408000;
      19159: inst = 32'hc40480e;
      19160: inst = 32'h8220000;
      19161: inst = 32'h10408000;
      19162: inst = 32'hc40480f;
      19163: inst = 32'h8220000;
      19164: inst = 32'h10408000;
      19165: inst = 32'hc404810;
      19166: inst = 32'h8220000;
      19167: inst = 32'h10408000;
      19168: inst = 32'hc404811;
      19169: inst = 32'h8220000;
      19170: inst = 32'h10408000;
      19171: inst = 32'hc40482b;
      19172: inst = 32'h8220000;
      19173: inst = 32'h10408000;
      19174: inst = 32'hc40482c;
      19175: inst = 32'h8220000;
      19176: inst = 32'h10408000;
      19177: inst = 32'hc40482e;
      19178: inst = 32'h8220000;
      19179: inst = 32'h10408000;
      19180: inst = 32'hc40482f;
      19181: inst = 32'h8220000;
      19182: inst = 32'h10408000;
      19183: inst = 32'hc404830;
      19184: inst = 32'h8220000;
      19185: inst = 32'h10408000;
      19186: inst = 32'hc404831;
      19187: inst = 32'h8220000;
      19188: inst = 32'h10408000;
      19189: inst = 32'hc404832;
      19190: inst = 32'h8220000;
      19191: inst = 32'h10408000;
      19192: inst = 32'hc404837;
      19193: inst = 32'h8220000;
      19194: inst = 32'h10408000;
      19195: inst = 32'hc404838;
      19196: inst = 32'h8220000;
      19197: inst = 32'h10408000;
      19198: inst = 32'hc40483a;
      19199: inst = 32'h8220000;
      19200: inst = 32'h10408000;
      19201: inst = 32'hc40483b;
      19202: inst = 32'h8220000;
      19203: inst = 32'h10408000;
      19204: inst = 32'hc40483c;
      19205: inst = 32'h8220000;
      19206: inst = 32'h10408000;
      19207: inst = 32'hc40483d;
      19208: inst = 32'h8220000;
      19209: inst = 32'h10408000;
      19210: inst = 32'hc40483e;
      19211: inst = 32'h8220000;
      19212: inst = 32'h10408000;
      19213: inst = 32'hc404846;
      19214: inst = 32'h8220000;
      19215: inst = 32'h10408000;
      19216: inst = 32'hc404847;
      19217: inst = 32'h8220000;
      19218: inst = 32'h10408000;
      19219: inst = 32'hc404848;
      19220: inst = 32'h8220000;
      19221: inst = 32'h10408000;
      19222: inst = 32'hc404850;
      19223: inst = 32'h8220000;
      19224: inst = 32'h10408000;
      19225: inst = 32'hc404851;
      19226: inst = 32'h8220000;
      19227: inst = 32'h10408000;
      19228: inst = 32'hc404859;
      19229: inst = 32'h8220000;
      19230: inst = 32'h10408000;
      19231: inst = 32'hc40485a;
      19232: inst = 32'h8220000;
      19233: inst = 32'h10408000;
      19234: inst = 32'hc40485f;
      19235: inst = 32'h8220000;
      19236: inst = 32'h10408000;
      19237: inst = 32'hc404860;
      19238: inst = 32'h8220000;
      19239: inst = 32'h10408000;
      19240: inst = 32'hc404861;
      19241: inst = 32'h8220000;
      19242: inst = 32'h10408000;
      19243: inst = 32'hc404862;
      19244: inst = 32'h8220000;
      19245: inst = 32'h10408000;
      19246: inst = 32'hc404869;
      19247: inst = 32'h8220000;
      19248: inst = 32'h10408000;
      19249: inst = 32'hc40486a;
      19250: inst = 32'h8220000;
      19251: inst = 32'h10408000;
      19252: inst = 32'hc40486c;
      19253: inst = 32'h8220000;
      19254: inst = 32'h10408000;
      19255: inst = 32'hc40486d;
      19256: inst = 32'h8220000;
      19257: inst = 32'h10408000;
      19258: inst = 32'hc40486e;
      19259: inst = 32'h8220000;
      19260: inst = 32'h10408000;
      19261: inst = 32'hc40486f;
      19262: inst = 32'h8220000;
      19263: inst = 32'h10408000;
      19264: inst = 32'hc404870;
      19265: inst = 32'h8220000;
      19266: inst = 32'h10408000;
      19267: inst = 32'hc404871;
      19268: inst = 32'h8220000;
      19269: inst = 32'h10408000;
      19270: inst = 32'hc404872;
      19271: inst = 32'h8220000;
      19272: inst = 32'h10408000;
      19273: inst = 32'hc40488b;
      19274: inst = 32'h8220000;
      19275: inst = 32'h10408000;
      19276: inst = 32'hc40488c;
      19277: inst = 32'h8220000;
      19278: inst = 32'h10408000;
      19279: inst = 32'hc404897;
      19280: inst = 32'h8220000;
      19281: inst = 32'h10408000;
      19282: inst = 32'hc404898;
      19283: inst = 32'h8220000;
      19284: inst = 32'h10408000;
      19285: inst = 32'hc4048a6;
      19286: inst = 32'h8220000;
      19287: inst = 32'h10408000;
      19288: inst = 32'hc4048b0;
      19289: inst = 32'h8220000;
      19290: inst = 32'h10408000;
      19291: inst = 32'hc4048b1;
      19292: inst = 32'h8220000;
      19293: inst = 32'h10408000;
      19294: inst = 32'hc4048b4;
      19295: inst = 32'h8220000;
      19296: inst = 32'h10408000;
      19297: inst = 32'hc4048b5;
      19298: inst = 32'h8220000;
      19299: inst = 32'h10408000;
      19300: inst = 32'hc4048b9;
      19301: inst = 32'h8220000;
      19302: inst = 32'h10408000;
      19303: inst = 32'hc4048ba;
      19304: inst = 32'h8220000;
      19305: inst = 32'h10408000;
      19306: inst = 32'hc4048bf;
      19307: inst = 32'h8220000;
      19308: inst = 32'h10408000;
      19309: inst = 32'hc4048c9;
      19310: inst = 32'h8220000;
      19311: inst = 32'h10408000;
      19312: inst = 32'hc4048ca;
      19313: inst = 32'h8220000;
      19314: inst = 32'h10408000;
      19315: inst = 32'hc4048d1;
      19316: inst = 32'h8220000;
      19317: inst = 32'h10408000;
      19318: inst = 32'hc4048d2;
      19319: inst = 32'h8220000;
      19320: inst = 32'h10408000;
      19321: inst = 32'hc4048d3;
      19322: inst = 32'h8220000;
      19323: inst = 32'h10408000;
      19324: inst = 32'hc4048eb;
      19325: inst = 32'h8220000;
      19326: inst = 32'h10408000;
      19327: inst = 32'hc4048ec;
      19328: inst = 32'h8220000;
      19329: inst = 32'h10408000;
      19330: inst = 32'hc4048ed;
      19331: inst = 32'h8220000;
      19332: inst = 32'h10408000;
      19333: inst = 32'hc4048ee;
      19334: inst = 32'h8220000;
      19335: inst = 32'h10408000;
      19336: inst = 32'hc4048ef;
      19337: inst = 32'h8220000;
      19338: inst = 32'h10408000;
      19339: inst = 32'hc4048f0;
      19340: inst = 32'h8220000;
      19341: inst = 32'h10408000;
      19342: inst = 32'hc4048f1;
      19343: inst = 32'h8220000;
      19344: inst = 32'h10408000;
      19345: inst = 32'hc4048f2;
      19346: inst = 32'h8220000;
      19347: inst = 32'h10408000;
      19348: inst = 32'hc4048f3;
      19349: inst = 32'h8220000;
      19350: inst = 32'h10408000;
      19351: inst = 32'hc4048f4;
      19352: inst = 32'h8220000;
      19353: inst = 32'h10408000;
      19354: inst = 32'hc4048f5;
      19355: inst = 32'h8220000;
      19356: inst = 32'h10408000;
      19357: inst = 32'hc4048f7;
      19358: inst = 32'h8220000;
      19359: inst = 32'h10408000;
      19360: inst = 32'hc4048f8;
      19361: inst = 32'h8220000;
      19362: inst = 32'h10408000;
      19363: inst = 32'hc4048f9;
      19364: inst = 32'h8220000;
      19365: inst = 32'h10408000;
      19366: inst = 32'hc4048fa;
      19367: inst = 32'h8220000;
      19368: inst = 32'h10408000;
      19369: inst = 32'hc4048fb;
      19370: inst = 32'h8220000;
      19371: inst = 32'h10408000;
      19372: inst = 32'hc4048fc;
      19373: inst = 32'h8220000;
      19374: inst = 32'h10408000;
      19375: inst = 32'hc4048fd;
      19376: inst = 32'h8220000;
      19377: inst = 32'h10408000;
      19378: inst = 32'hc4048fe;
      19379: inst = 32'h8220000;
      19380: inst = 32'h10408000;
      19381: inst = 32'hc4048ff;
      19382: inst = 32'h8220000;
      19383: inst = 32'h10408000;
      19384: inst = 32'hc404900;
      19385: inst = 32'h8220000;
      19386: inst = 32'h10408000;
      19387: inst = 32'hc404901;
      19388: inst = 32'h8220000;
      19389: inst = 32'h10408000;
      19390: inst = 32'hc404904;
      19391: inst = 32'h8220000;
      19392: inst = 32'h10408000;
      19393: inst = 32'hc404905;
      19394: inst = 32'h8220000;
      19395: inst = 32'h10408000;
      19396: inst = 32'hc404906;
      19397: inst = 32'h8220000;
      19398: inst = 32'h10408000;
      19399: inst = 32'hc404907;
      19400: inst = 32'h8220000;
      19401: inst = 32'h10408000;
      19402: inst = 32'hc404908;
      19403: inst = 32'h8220000;
      19404: inst = 32'h10408000;
      19405: inst = 32'hc404909;
      19406: inst = 32'h8220000;
      19407: inst = 32'h10408000;
      19408: inst = 32'hc40490a;
      19409: inst = 32'h8220000;
      19410: inst = 32'h10408000;
      19411: inst = 32'hc40490b;
      19412: inst = 32'h8220000;
      19413: inst = 32'h10408000;
      19414: inst = 32'hc40490c;
      19415: inst = 32'h8220000;
      19416: inst = 32'h10408000;
      19417: inst = 32'hc40490d;
      19418: inst = 32'h8220000;
      19419: inst = 32'h10408000;
      19420: inst = 32'hc404910;
      19421: inst = 32'h8220000;
      19422: inst = 32'h10408000;
      19423: inst = 32'hc404911;
      19424: inst = 32'h8220000;
      19425: inst = 32'h10408000;
      19426: inst = 32'hc404912;
      19427: inst = 32'h8220000;
      19428: inst = 32'h10408000;
      19429: inst = 32'hc404913;
      19430: inst = 32'h8220000;
      19431: inst = 32'h10408000;
      19432: inst = 32'hc404914;
      19433: inst = 32'h8220000;
      19434: inst = 32'h10408000;
      19435: inst = 32'hc404915;
      19436: inst = 32'h8220000;
      19437: inst = 32'h10408000;
      19438: inst = 32'hc404916;
      19439: inst = 32'h8220000;
      19440: inst = 32'h10408000;
      19441: inst = 32'hc404917;
      19442: inst = 32'h8220000;
      19443: inst = 32'h10408000;
      19444: inst = 32'hc404918;
      19445: inst = 32'h8220000;
      19446: inst = 32'h10408000;
      19447: inst = 32'hc404919;
      19448: inst = 32'h8220000;
      19449: inst = 32'h10408000;
      19450: inst = 32'hc40491a;
      19451: inst = 32'h8220000;
      19452: inst = 32'h10408000;
      19453: inst = 32'hc40491e;
      19454: inst = 32'h8220000;
      19455: inst = 32'h10408000;
      19456: inst = 32'hc40491f;
      19457: inst = 32'h8220000;
      19458: inst = 32'h10408000;
      19459: inst = 32'hc404920;
      19460: inst = 32'h8220000;
      19461: inst = 32'h10408000;
      19462: inst = 32'hc404921;
      19463: inst = 32'h8220000;
      19464: inst = 32'h10408000;
      19465: inst = 32'hc404922;
      19466: inst = 32'h8220000;
      19467: inst = 32'h10408000;
      19468: inst = 32'hc404923;
      19469: inst = 32'h8220000;
      19470: inst = 32'h10408000;
      19471: inst = 32'hc404924;
      19472: inst = 32'h8220000;
      19473: inst = 32'h10408000;
      19474: inst = 32'hc404925;
      19475: inst = 32'h8220000;
      19476: inst = 32'h10408000;
      19477: inst = 32'hc404926;
      19478: inst = 32'h8220000;
      19479: inst = 32'h10408000;
      19480: inst = 32'hc404927;
      19481: inst = 32'h8220000;
      19482: inst = 32'h10408000;
      19483: inst = 32'hc404929;
      19484: inst = 32'h8220000;
      19485: inst = 32'h10408000;
      19486: inst = 32'hc40492a;
      19487: inst = 32'h8220000;
      19488: inst = 32'h10408000;
      19489: inst = 32'hc40492b;
      19490: inst = 32'h8220000;
      19491: inst = 32'h10408000;
      19492: inst = 32'hc40492c;
      19493: inst = 32'h8220000;
      19494: inst = 32'h10408000;
      19495: inst = 32'hc40492d;
      19496: inst = 32'h8220000;
      19497: inst = 32'h10408000;
      19498: inst = 32'hc40492e;
      19499: inst = 32'h8220000;
      19500: inst = 32'h10408000;
      19501: inst = 32'hc40492f;
      19502: inst = 32'h8220000;
      19503: inst = 32'h10408000;
      19504: inst = 32'hc404930;
      19505: inst = 32'h8220000;
      19506: inst = 32'h10408000;
      19507: inst = 32'hc404931;
      19508: inst = 32'h8220000;
      19509: inst = 32'h10408000;
      19510: inst = 32'hc404932;
      19511: inst = 32'h8220000;
      19512: inst = 32'h10408000;
      19513: inst = 32'hc404933;
      19514: inst = 32'h8220000;
      19515: inst = 32'h10408000;
      19516: inst = 32'hc40494b;
      19517: inst = 32'h8220000;
      19518: inst = 32'h10408000;
      19519: inst = 32'hc40494c;
      19520: inst = 32'h8220000;
      19521: inst = 32'h10408000;
      19522: inst = 32'hc40494d;
      19523: inst = 32'h8220000;
      19524: inst = 32'h10408000;
      19525: inst = 32'hc40494e;
      19526: inst = 32'h8220000;
      19527: inst = 32'h10408000;
      19528: inst = 32'hc40494f;
      19529: inst = 32'h8220000;
      19530: inst = 32'h10408000;
      19531: inst = 32'hc404950;
      19532: inst = 32'h8220000;
      19533: inst = 32'h10408000;
      19534: inst = 32'hc404951;
      19535: inst = 32'h8220000;
      19536: inst = 32'h10408000;
      19537: inst = 32'hc404952;
      19538: inst = 32'h8220000;
      19539: inst = 32'h10408000;
      19540: inst = 32'hc404953;
      19541: inst = 32'h8220000;
      19542: inst = 32'h10408000;
      19543: inst = 32'hc404954;
      19544: inst = 32'h8220000;
      19545: inst = 32'h10408000;
      19546: inst = 32'hc404957;
      19547: inst = 32'h8220000;
      19548: inst = 32'h10408000;
      19549: inst = 32'hc404958;
      19550: inst = 32'h8220000;
      19551: inst = 32'h10408000;
      19552: inst = 32'hc404959;
      19553: inst = 32'h8220000;
      19554: inst = 32'h10408000;
      19555: inst = 32'hc40495a;
      19556: inst = 32'h8220000;
      19557: inst = 32'h10408000;
      19558: inst = 32'hc40495b;
      19559: inst = 32'h8220000;
      19560: inst = 32'h10408000;
      19561: inst = 32'hc40495c;
      19562: inst = 32'h8220000;
      19563: inst = 32'h10408000;
      19564: inst = 32'hc40495d;
      19565: inst = 32'h8220000;
      19566: inst = 32'h10408000;
      19567: inst = 32'hc40495e;
      19568: inst = 32'h8220000;
      19569: inst = 32'h10408000;
      19570: inst = 32'hc40495f;
      19571: inst = 32'h8220000;
      19572: inst = 32'h10408000;
      19573: inst = 32'hc404960;
      19574: inst = 32'h8220000;
      19575: inst = 32'h10408000;
      19576: inst = 32'hc404961;
      19577: inst = 32'h8220000;
      19578: inst = 32'h10408000;
      19579: inst = 32'hc404963;
      19580: inst = 32'h8220000;
      19581: inst = 32'h10408000;
      19582: inst = 32'hc404964;
      19583: inst = 32'h8220000;
      19584: inst = 32'h10408000;
      19585: inst = 32'hc404965;
      19586: inst = 32'h8220000;
      19587: inst = 32'h10408000;
      19588: inst = 32'hc404966;
      19589: inst = 32'h8220000;
      19590: inst = 32'h10408000;
      19591: inst = 32'hc404967;
      19592: inst = 32'h8220000;
      19593: inst = 32'h10408000;
      19594: inst = 32'hc404968;
      19595: inst = 32'h8220000;
      19596: inst = 32'h10408000;
      19597: inst = 32'hc404969;
      19598: inst = 32'h8220000;
      19599: inst = 32'h10408000;
      19600: inst = 32'hc40496a;
      19601: inst = 32'h8220000;
      19602: inst = 32'h10408000;
      19603: inst = 32'hc40496b;
      19604: inst = 32'h8220000;
      19605: inst = 32'h10408000;
      19606: inst = 32'hc40496c;
      19607: inst = 32'h8220000;
      19608: inst = 32'h10408000;
      19609: inst = 32'hc40496d;
      19610: inst = 32'h8220000;
      19611: inst = 32'h10408000;
      19612: inst = 32'hc404970;
      19613: inst = 32'h8220000;
      19614: inst = 32'h10408000;
      19615: inst = 32'hc404971;
      19616: inst = 32'h8220000;
      19617: inst = 32'h10408000;
      19618: inst = 32'hc404972;
      19619: inst = 32'h8220000;
      19620: inst = 32'h10408000;
      19621: inst = 32'hc404973;
      19622: inst = 32'h8220000;
      19623: inst = 32'h10408000;
      19624: inst = 32'hc404974;
      19625: inst = 32'h8220000;
      19626: inst = 32'h10408000;
      19627: inst = 32'hc404975;
      19628: inst = 32'h8220000;
      19629: inst = 32'h10408000;
      19630: inst = 32'hc404976;
      19631: inst = 32'h8220000;
      19632: inst = 32'h10408000;
      19633: inst = 32'hc404977;
      19634: inst = 32'h8220000;
      19635: inst = 32'h10408000;
      19636: inst = 32'hc404978;
      19637: inst = 32'h8220000;
      19638: inst = 32'h10408000;
      19639: inst = 32'hc404979;
      19640: inst = 32'h8220000;
      19641: inst = 32'h10408000;
      19642: inst = 32'hc40497d;
      19643: inst = 32'h8220000;
      19644: inst = 32'h10408000;
      19645: inst = 32'hc40497e;
      19646: inst = 32'h8220000;
      19647: inst = 32'h10408000;
      19648: inst = 32'hc40497f;
      19649: inst = 32'h8220000;
      19650: inst = 32'h10408000;
      19651: inst = 32'hc404980;
      19652: inst = 32'h8220000;
      19653: inst = 32'h10408000;
      19654: inst = 32'hc404981;
      19655: inst = 32'h8220000;
      19656: inst = 32'h10408000;
      19657: inst = 32'hc404982;
      19658: inst = 32'h8220000;
      19659: inst = 32'h10408000;
      19660: inst = 32'hc404983;
      19661: inst = 32'h8220000;
      19662: inst = 32'h10408000;
      19663: inst = 32'hc404984;
      19664: inst = 32'h8220000;
      19665: inst = 32'h10408000;
      19666: inst = 32'hc404985;
      19667: inst = 32'h8220000;
      19668: inst = 32'h10408000;
      19669: inst = 32'hc404986;
      19670: inst = 32'h8220000;
      19671: inst = 32'h10408000;
      19672: inst = 32'hc404987;
      19673: inst = 32'h8220000;
      19674: inst = 32'h10408000;
      19675: inst = 32'hc404989;
      19676: inst = 32'h8220000;
      19677: inst = 32'h10408000;
      19678: inst = 32'hc40498a;
      19679: inst = 32'h8220000;
      19680: inst = 32'h10408000;
      19681: inst = 32'hc40498b;
      19682: inst = 32'h8220000;
      19683: inst = 32'h10408000;
      19684: inst = 32'hc40498c;
      19685: inst = 32'h8220000;
      19686: inst = 32'h10408000;
      19687: inst = 32'hc40498d;
      19688: inst = 32'h8220000;
      19689: inst = 32'h10408000;
      19690: inst = 32'hc40498e;
      19691: inst = 32'h8220000;
      19692: inst = 32'h10408000;
      19693: inst = 32'hc40498f;
      19694: inst = 32'h8220000;
      19695: inst = 32'h10408000;
      19696: inst = 32'hc404990;
      19697: inst = 32'h8220000;
      19698: inst = 32'h10408000;
      19699: inst = 32'hc404991;
      19700: inst = 32'h8220000;
      19701: inst = 32'h10408000;
      19702: inst = 32'hc404992;
      19703: inst = 32'h8220000;
      19704: inst = 32'h10408000;
      19705: inst = 32'hc404993;
      19706: inst = 32'h8220000;
      19707: inst = 32'h10408000;
      19708: inst = 32'hc404dcd;
      19709: inst = 32'h8220000;
      19710: inst = 32'h10408000;
      19711: inst = 32'hc404dce;
      19712: inst = 32'h8220000;
      19713: inst = 32'h10408000;
      19714: inst = 32'hc404dcf;
      19715: inst = 32'h8220000;
      19716: inst = 32'h10408000;
      19717: inst = 32'hc404dd0;
      19718: inst = 32'h8220000;
      19719: inst = 32'h10408000;
      19720: inst = 32'hc404dd1;
      19721: inst = 32'h8220000;
      19722: inst = 32'h10408000;
      19723: inst = 32'hc404dd2;
      19724: inst = 32'h8220000;
      19725: inst = 32'h10408000;
      19726: inst = 32'hc404dd3;
      19727: inst = 32'h8220000;
      19728: inst = 32'h10408000;
      19729: inst = 32'hc404dd4;
      19730: inst = 32'h8220000;
      19731: inst = 32'h10408000;
      19732: inst = 32'hc404dd5;
      19733: inst = 32'h8220000;
      19734: inst = 32'h10408000;
      19735: inst = 32'hc404dd7;
      19736: inst = 32'h8220000;
      19737: inst = 32'h10408000;
      19738: inst = 32'hc404dd8;
      19739: inst = 32'h8220000;
      19740: inst = 32'h10408000;
      19741: inst = 32'hc404dd9;
      19742: inst = 32'h8220000;
      19743: inst = 32'h10408000;
      19744: inst = 32'hc404dda;
      19745: inst = 32'h8220000;
      19746: inst = 32'h10408000;
      19747: inst = 32'hc404ddb;
      19748: inst = 32'h8220000;
      19749: inst = 32'h10408000;
      19750: inst = 32'hc404ddc;
      19751: inst = 32'h8220000;
      19752: inst = 32'h10408000;
      19753: inst = 32'hc404ddd;
      19754: inst = 32'h8220000;
      19755: inst = 32'h10408000;
      19756: inst = 32'hc404dde;
      19757: inst = 32'h8220000;
      19758: inst = 32'h10408000;
      19759: inst = 32'hc404ddf;
      19760: inst = 32'h8220000;
      19761: inst = 32'h10408000;
      19762: inst = 32'hc404de0;
      19763: inst = 32'h8220000;
      19764: inst = 32'h10408000;
      19765: inst = 32'hc404de1;
      19766: inst = 32'h8220000;
      19767: inst = 32'h10408000;
      19768: inst = 32'hc404de2;
      19769: inst = 32'h8220000;
      19770: inst = 32'h10408000;
      19771: inst = 32'hc404de4;
      19772: inst = 32'h8220000;
      19773: inst = 32'h10408000;
      19774: inst = 32'hc404de5;
      19775: inst = 32'h8220000;
      19776: inst = 32'h10408000;
      19777: inst = 32'hc404de6;
      19778: inst = 32'h8220000;
      19779: inst = 32'h10408000;
      19780: inst = 32'hc404de7;
      19781: inst = 32'h8220000;
      19782: inst = 32'h10408000;
      19783: inst = 32'hc404de8;
      19784: inst = 32'h8220000;
      19785: inst = 32'h10408000;
      19786: inst = 32'hc404de9;
      19787: inst = 32'h8220000;
      19788: inst = 32'h10408000;
      19789: inst = 32'hc404dea;
      19790: inst = 32'h8220000;
      19791: inst = 32'h10408000;
      19792: inst = 32'hc404deb;
      19793: inst = 32'h8220000;
      19794: inst = 32'h10408000;
      19795: inst = 32'hc404dec;
      19796: inst = 32'h8220000;
      19797: inst = 32'h10408000;
      19798: inst = 32'hc404ded;
      19799: inst = 32'h8220000;
      19800: inst = 32'h10408000;
      19801: inst = 32'hc404df0;
      19802: inst = 32'h8220000;
      19803: inst = 32'h10408000;
      19804: inst = 32'hc404df1;
      19805: inst = 32'h8220000;
      19806: inst = 32'h10408000;
      19807: inst = 32'hc404df2;
      19808: inst = 32'h8220000;
      19809: inst = 32'h10408000;
      19810: inst = 32'hc404dfc;
      19811: inst = 32'h8220000;
      19812: inst = 32'h10408000;
      19813: inst = 32'hc404dfd;
      19814: inst = 32'h8220000;
      19815: inst = 32'h10408000;
      19816: inst = 32'hc404dfe;
      19817: inst = 32'h8220000;
      19818: inst = 32'h10408000;
      19819: inst = 32'hc404dff;
      19820: inst = 32'h8220000;
      19821: inst = 32'h10408000;
      19822: inst = 32'hc404e00;
      19823: inst = 32'h8220000;
      19824: inst = 32'h10408000;
      19825: inst = 32'hc404e01;
      19826: inst = 32'h8220000;
      19827: inst = 32'h10408000;
      19828: inst = 32'hc404e02;
      19829: inst = 32'h8220000;
      19830: inst = 32'h10408000;
      19831: inst = 32'hc404e03;
      19832: inst = 32'h8220000;
      19833: inst = 32'h10408000;
      19834: inst = 32'hc404e04;
      19835: inst = 32'h8220000;
      19836: inst = 32'h10408000;
      19837: inst = 32'hc404e05;
      19838: inst = 32'h8220000;
      19839: inst = 32'h10408000;
      19840: inst = 32'hc404e06;
      19841: inst = 32'h8220000;
      19842: inst = 32'h10408000;
      19843: inst = 32'hc404e07;
      19844: inst = 32'h8220000;
      19845: inst = 32'h10408000;
      19846: inst = 32'hc404e0b;
      19847: inst = 32'h8220000;
      19848: inst = 32'h10408000;
      19849: inst = 32'hc404e0c;
      19850: inst = 32'h8220000;
      19851: inst = 32'h10408000;
      19852: inst = 32'hc404e0d;
      19853: inst = 32'h8220000;
      19854: inst = 32'h10408000;
      19855: inst = 32'hc404e0e;
      19856: inst = 32'h8220000;
      19857: inst = 32'h10408000;
      19858: inst = 32'hc404e0f;
      19859: inst = 32'h8220000;
      19860: inst = 32'h10408000;
      19861: inst = 32'hc404e10;
      19862: inst = 32'h8220000;
      19863: inst = 32'h10408000;
      19864: inst = 32'hc404e11;
      19865: inst = 32'h8220000;
      19866: inst = 32'h10408000;
      19867: inst = 32'hc404e12;
      19868: inst = 32'h8220000;
      19869: inst = 32'h10408000;
      19870: inst = 32'hc404e13;
      19871: inst = 32'h8220000;
      19872: inst = 32'h10408000;
      19873: inst = 32'hc404e2c;
      19874: inst = 32'h8220000;
      19875: inst = 32'h10408000;
      19876: inst = 32'hc404e2d;
      19877: inst = 32'h8220000;
      19878: inst = 32'h10408000;
      19879: inst = 32'hc404e2e;
      19880: inst = 32'h8220000;
      19881: inst = 32'h10408000;
      19882: inst = 32'hc404e2f;
      19883: inst = 32'h8220000;
      19884: inst = 32'h10408000;
      19885: inst = 32'hc404e30;
      19886: inst = 32'h8220000;
      19887: inst = 32'h10408000;
      19888: inst = 32'hc404e31;
      19889: inst = 32'h8220000;
      19890: inst = 32'h10408000;
      19891: inst = 32'hc404e32;
      19892: inst = 32'h8220000;
      19893: inst = 32'h10408000;
      19894: inst = 32'hc404e33;
      19895: inst = 32'h8220000;
      19896: inst = 32'h10408000;
      19897: inst = 32'hc404e34;
      19898: inst = 32'h8220000;
      19899: inst = 32'h10408000;
      19900: inst = 32'hc404e35;
      19901: inst = 32'h8220000;
      19902: inst = 32'h10408000;
      19903: inst = 32'hc404e38;
      19904: inst = 32'h8220000;
      19905: inst = 32'h10408000;
      19906: inst = 32'hc404e39;
      19907: inst = 32'h8220000;
      19908: inst = 32'h10408000;
      19909: inst = 32'hc404e3a;
      19910: inst = 32'h8220000;
      19911: inst = 32'h10408000;
      19912: inst = 32'hc404e3b;
      19913: inst = 32'h8220000;
      19914: inst = 32'h10408000;
      19915: inst = 32'hc404e3c;
      19916: inst = 32'h8220000;
      19917: inst = 32'h10408000;
      19918: inst = 32'hc404e3d;
      19919: inst = 32'h8220000;
      19920: inst = 32'h10408000;
      19921: inst = 32'hc404e3e;
      19922: inst = 32'h8220000;
      19923: inst = 32'h10408000;
      19924: inst = 32'hc404e3f;
      19925: inst = 32'h8220000;
      19926: inst = 32'h10408000;
      19927: inst = 32'hc404e40;
      19928: inst = 32'h8220000;
      19929: inst = 32'h10408000;
      19930: inst = 32'hc404e41;
      19931: inst = 32'h8220000;
      19932: inst = 32'h10408000;
      19933: inst = 32'hc404e42;
      19934: inst = 32'h8220000;
      19935: inst = 32'h10408000;
      19936: inst = 32'hc404e44;
      19937: inst = 32'h8220000;
      19938: inst = 32'h10408000;
      19939: inst = 32'hc404e45;
      19940: inst = 32'h8220000;
      19941: inst = 32'h10408000;
      19942: inst = 32'hc404e46;
      19943: inst = 32'h8220000;
      19944: inst = 32'h10408000;
      19945: inst = 32'hc404e47;
      19946: inst = 32'h8220000;
      19947: inst = 32'h10408000;
      19948: inst = 32'hc404e48;
      19949: inst = 32'h8220000;
      19950: inst = 32'h10408000;
      19951: inst = 32'hc404e49;
      19952: inst = 32'h8220000;
      19953: inst = 32'h10408000;
      19954: inst = 32'hc404e4a;
      19955: inst = 32'h8220000;
      19956: inst = 32'h10408000;
      19957: inst = 32'hc404e4b;
      19958: inst = 32'h8220000;
      19959: inst = 32'h10408000;
      19960: inst = 32'hc404e4c;
      19961: inst = 32'h8220000;
      19962: inst = 32'h10408000;
      19963: inst = 32'hc404e4d;
      19964: inst = 32'h8220000;
      19965: inst = 32'h10408000;
      19966: inst = 32'hc404e50;
      19967: inst = 32'h8220000;
      19968: inst = 32'h10408000;
      19969: inst = 32'hc404e51;
      19970: inst = 32'h8220000;
      19971: inst = 32'h10408000;
      19972: inst = 32'hc404e52;
      19973: inst = 32'h8220000;
      19974: inst = 32'h10408000;
      19975: inst = 32'hc404e53;
      19976: inst = 32'h8220000;
      19977: inst = 32'h10408000;
      19978: inst = 32'hc404e5c;
      19979: inst = 32'h8220000;
      19980: inst = 32'h10408000;
      19981: inst = 32'hc404e5d;
      19982: inst = 32'h8220000;
      19983: inst = 32'h10408000;
      19984: inst = 32'hc404e5e;
      19985: inst = 32'h8220000;
      19986: inst = 32'h10408000;
      19987: inst = 32'hc404e5f;
      19988: inst = 32'h8220000;
      19989: inst = 32'h10408000;
      19990: inst = 32'hc404e60;
      19991: inst = 32'h8220000;
      19992: inst = 32'h10408000;
      19993: inst = 32'hc404e61;
      19994: inst = 32'h8220000;
      19995: inst = 32'h10408000;
      19996: inst = 32'hc404e62;
      19997: inst = 32'h8220000;
      19998: inst = 32'h10408000;
      19999: inst = 32'hc404e63;
      20000: inst = 32'h8220000;
      20001: inst = 32'h10408000;
      20002: inst = 32'hc404e64;
      20003: inst = 32'h8220000;
      20004: inst = 32'h10408000;
      20005: inst = 32'hc404e65;
      20006: inst = 32'h8220000;
      20007: inst = 32'h10408000;
      20008: inst = 32'hc404e66;
      20009: inst = 32'h8220000;
      20010: inst = 32'h10408000;
      20011: inst = 32'hc404e6a;
      20012: inst = 32'h8220000;
      20013: inst = 32'h10408000;
      20014: inst = 32'hc404e6b;
      20015: inst = 32'h8220000;
      20016: inst = 32'h10408000;
      20017: inst = 32'hc404e6c;
      20018: inst = 32'h8220000;
      20019: inst = 32'h10408000;
      20020: inst = 32'hc404e6d;
      20021: inst = 32'h8220000;
      20022: inst = 32'h10408000;
      20023: inst = 32'hc404e6e;
      20024: inst = 32'h8220000;
      20025: inst = 32'h10408000;
      20026: inst = 32'hc404e6f;
      20027: inst = 32'h8220000;
      20028: inst = 32'h10408000;
      20029: inst = 32'hc404e70;
      20030: inst = 32'h8220000;
      20031: inst = 32'h10408000;
      20032: inst = 32'hc404e71;
      20033: inst = 32'h8220000;
      20034: inst = 32'h10408000;
      20035: inst = 32'hc404e72;
      20036: inst = 32'h8220000;
      20037: inst = 32'h10408000;
      20038: inst = 32'hc404e73;
      20039: inst = 32'h8220000;
      20040: inst = 32'h10408000;
      20041: inst = 32'hc404e8b;
      20042: inst = 32'h8220000;
      20043: inst = 32'h10408000;
      20044: inst = 32'hc404e8c;
      20045: inst = 32'h8220000;
      20046: inst = 32'h10408000;
      20047: inst = 32'hc404e8d;
      20048: inst = 32'h8220000;
      20049: inst = 32'h10408000;
      20050: inst = 32'hc404e99;
      20051: inst = 32'h8220000;
      20052: inst = 32'h10408000;
      20053: inst = 32'hc404e9a;
      20054: inst = 32'h8220000;
      20055: inst = 32'h10408000;
      20056: inst = 32'hc404e9b;
      20057: inst = 32'h8220000;
      20058: inst = 32'h10408000;
      20059: inst = 32'hc404e9c;
      20060: inst = 32'h8220000;
      20061: inst = 32'h10408000;
      20062: inst = 32'hc404ea4;
      20063: inst = 32'h8220000;
      20064: inst = 32'h10408000;
      20065: inst = 32'hc404ea5;
      20066: inst = 32'h8220000;
      20067: inst = 32'h10408000;
      20068: inst = 32'hc404eac;
      20069: inst = 32'h8220000;
      20070: inst = 32'h10408000;
      20071: inst = 32'hc404ead;
      20072: inst = 32'h8220000;
      20073: inst = 32'h10408000;
      20074: inst = 32'hc404eb0;
      20075: inst = 32'h8220000;
      20076: inst = 32'h10408000;
      20077: inst = 32'hc404eb1;
      20078: inst = 32'h8220000;
      20079: inst = 32'h10408000;
      20080: inst = 32'hc404eb2;
      20081: inst = 32'h8220000;
      20082: inst = 32'h10408000;
      20083: inst = 32'hc404eb3;
      20084: inst = 32'h8220000;
      20085: inst = 32'h10408000;
      20086: inst = 32'hc404eb4;
      20087: inst = 32'h8220000;
      20088: inst = 32'h10408000;
      20089: inst = 32'hc404ebc;
      20090: inst = 32'h8220000;
      20091: inst = 32'h10408000;
      20092: inst = 32'hc404ebd;
      20093: inst = 32'h8220000;
      20094: inst = 32'h10408000;
      20095: inst = 32'hc404ec2;
      20096: inst = 32'h8220000;
      20097: inst = 32'h10408000;
      20098: inst = 32'hc404ec3;
      20099: inst = 32'h8220000;
      20100: inst = 32'h10408000;
      20101: inst = 32'hc404ec4;
      20102: inst = 32'h8220000;
      20103: inst = 32'h10408000;
      20104: inst = 32'hc404ec5;
      20105: inst = 32'h8220000;
      20106: inst = 32'h10408000;
      20107: inst = 32'hc404ec9;
      20108: inst = 32'h8220000;
      20109: inst = 32'h10408000;
      20110: inst = 32'hc404eca;
      20111: inst = 32'h8220000;
      20112: inst = 32'h10408000;
      20113: inst = 32'hc404eeb;
      20114: inst = 32'h8220000;
      20115: inst = 32'h10408000;
      20116: inst = 32'hc404eec;
      20117: inst = 32'h8220000;
      20118: inst = 32'h10408000;
      20119: inst = 32'hc404efa;
      20120: inst = 32'h8220000;
      20121: inst = 32'h10408000;
      20122: inst = 32'hc404efb;
      20123: inst = 32'h8220000;
      20124: inst = 32'h10408000;
      20125: inst = 32'hc404efc;
      20126: inst = 32'h8220000;
      20127: inst = 32'h10408000;
      20128: inst = 32'hc404f04;
      20129: inst = 32'h8220000;
      20130: inst = 32'h10408000;
      20131: inst = 32'hc404f05;
      20132: inst = 32'h8220000;
      20133: inst = 32'h10408000;
      20134: inst = 32'hc404f0c;
      20135: inst = 32'h8220000;
      20136: inst = 32'h10408000;
      20137: inst = 32'hc404f0d;
      20138: inst = 32'h8220000;
      20139: inst = 32'h10408000;
      20140: inst = 32'hc404f10;
      20141: inst = 32'h8220000;
      20142: inst = 32'h10408000;
      20143: inst = 32'hc404f12;
      20144: inst = 32'h8220000;
      20145: inst = 32'h10408000;
      20146: inst = 32'hc404f13;
      20147: inst = 32'h8220000;
      20148: inst = 32'h10408000;
      20149: inst = 32'hc404f14;
      20150: inst = 32'h8220000;
      20151: inst = 32'h10408000;
      20152: inst = 32'hc404f15;
      20153: inst = 32'h8220000;
      20154: inst = 32'h10408000;
      20155: inst = 32'hc404f1c;
      20156: inst = 32'h8220000;
      20157: inst = 32'h10408000;
      20158: inst = 32'hc404f1d;
      20159: inst = 32'h8220000;
      20160: inst = 32'h10408000;
      20161: inst = 32'hc404f22;
      20162: inst = 32'h8220000;
      20163: inst = 32'h10408000;
      20164: inst = 32'hc404f23;
      20165: inst = 32'h8220000;
      20166: inst = 32'h10408000;
      20167: inst = 32'hc404f24;
      20168: inst = 32'h8220000;
      20169: inst = 32'h10408000;
      20170: inst = 32'hc404f29;
      20171: inst = 32'h8220000;
      20172: inst = 32'h10408000;
      20173: inst = 32'hc404f2a;
      20174: inst = 32'h8220000;
      20175: inst = 32'h10408000;
      20176: inst = 32'hc404f4b;
      20177: inst = 32'h8220000;
      20178: inst = 32'h10408000;
      20179: inst = 32'hc404f4c;
      20180: inst = 32'h8220000;
      20181: inst = 32'h10408000;
      20182: inst = 32'hc404f4e;
      20183: inst = 32'h8220000;
      20184: inst = 32'h10408000;
      20185: inst = 32'hc404f4f;
      20186: inst = 32'h8220000;
      20187: inst = 32'h10408000;
      20188: inst = 32'hc404f50;
      20189: inst = 32'h8220000;
      20190: inst = 32'h10408000;
      20191: inst = 32'hc404f51;
      20192: inst = 32'h8220000;
      20193: inst = 32'h10408000;
      20194: inst = 32'hc404f52;
      20195: inst = 32'h8220000;
      20196: inst = 32'h10408000;
      20197: inst = 32'hc404f5b;
      20198: inst = 32'h8220000;
      20199: inst = 32'h10408000;
      20200: inst = 32'hc404f5c;
      20201: inst = 32'h8220000;
      20202: inst = 32'h10408000;
      20203: inst = 32'hc404f5d;
      20204: inst = 32'h8220000;
      20205: inst = 32'h10408000;
      20206: inst = 32'hc404f64;
      20207: inst = 32'h8220000;
      20208: inst = 32'h10408000;
      20209: inst = 32'hc404f65;
      20210: inst = 32'h8220000;
      20211: inst = 32'h10408000;
      20212: inst = 32'hc404f6c;
      20213: inst = 32'h8220000;
      20214: inst = 32'h10408000;
      20215: inst = 32'hc404f70;
      20216: inst = 32'h8220000;
      20217: inst = 32'h10408000;
      20218: inst = 32'hc404f71;
      20219: inst = 32'h8220000;
      20220: inst = 32'h10408000;
      20221: inst = 32'hc404f72;
      20222: inst = 32'h8220000;
      20223: inst = 32'h10408000;
      20224: inst = 32'hc404f73;
      20225: inst = 32'h8220000;
      20226: inst = 32'h10408000;
      20227: inst = 32'hc404f74;
      20228: inst = 32'h8220000;
      20229: inst = 32'h10408000;
      20230: inst = 32'hc404f75;
      20231: inst = 32'h8220000;
      20232: inst = 32'h10408000;
      20233: inst = 32'hc404f76;
      20234: inst = 32'h8220000;
      20235: inst = 32'h10408000;
      20236: inst = 32'hc404f7c;
      20237: inst = 32'h8220000;
      20238: inst = 32'h10408000;
      20239: inst = 32'hc404f7d;
      20240: inst = 32'h8220000;
      20241: inst = 32'h10408000;
      20242: inst = 32'hc404f7f;
      20243: inst = 32'h8220000;
      20244: inst = 32'h10408000;
      20245: inst = 32'hc404f80;
      20246: inst = 32'h8220000;
      20247: inst = 32'h10408000;
      20248: inst = 32'hc404f81;
      20249: inst = 32'h8220000;
      20250: inst = 32'h10408000;
      20251: inst = 32'hc404f82;
      20252: inst = 32'h8220000;
      20253: inst = 32'h10408000;
      20254: inst = 32'hc404f83;
      20255: inst = 32'h8220000;
      20256: inst = 32'h10408000;
      20257: inst = 32'hc404f89;
      20258: inst = 32'h8220000;
      20259: inst = 32'h10408000;
      20260: inst = 32'hc404f8a;
      20261: inst = 32'h8220000;
      20262: inst = 32'h10408000;
      20263: inst = 32'hc404f8c;
      20264: inst = 32'h8220000;
      20265: inst = 32'h10408000;
      20266: inst = 32'hc404f8d;
      20267: inst = 32'h8220000;
      20268: inst = 32'h10408000;
      20269: inst = 32'hc404f8e;
      20270: inst = 32'h8220000;
      20271: inst = 32'h10408000;
      20272: inst = 32'hc404f8f;
      20273: inst = 32'h8220000;
      20274: inst = 32'h10408000;
      20275: inst = 32'hc404f90;
      20276: inst = 32'h8220000;
      20277: inst = 32'h10408000;
      20278: inst = 32'hc404fab;
      20279: inst = 32'h8220000;
      20280: inst = 32'h10408000;
      20281: inst = 32'hc404fac;
      20282: inst = 32'h8220000;
      20283: inst = 32'h10408000;
      20284: inst = 32'hc404fae;
      20285: inst = 32'h8220000;
      20286: inst = 32'h10408000;
      20287: inst = 32'hc404faf;
      20288: inst = 32'h8220000;
      20289: inst = 32'h10408000;
      20290: inst = 32'hc404fb0;
      20291: inst = 32'h8220000;
      20292: inst = 32'h10408000;
      20293: inst = 32'hc404fb1;
      20294: inst = 32'h8220000;
      20295: inst = 32'h10408000;
      20296: inst = 32'hc404fb2;
      20297: inst = 32'h8220000;
      20298: inst = 32'h10408000;
      20299: inst = 32'hc404fbc;
      20300: inst = 32'h8220000;
      20301: inst = 32'h10408000;
      20302: inst = 32'hc404fbd;
      20303: inst = 32'h8220000;
      20304: inst = 32'h10408000;
      20305: inst = 32'hc404fbe;
      20306: inst = 32'h8220000;
      20307: inst = 32'h10408000;
      20308: inst = 32'hc404fc4;
      20309: inst = 32'h8220000;
      20310: inst = 32'h10408000;
      20311: inst = 32'hc404fc5;
      20312: inst = 32'h8220000;
      20313: inst = 32'h10408000;
      20314: inst = 32'hc404fd0;
      20315: inst = 32'h8220000;
      20316: inst = 32'h10408000;
      20317: inst = 32'hc404fd1;
      20318: inst = 32'h8220000;
      20319: inst = 32'h10408000;
      20320: inst = 32'hc404fd2;
      20321: inst = 32'h8220000;
      20322: inst = 32'h10408000;
      20323: inst = 32'hc404fd4;
      20324: inst = 32'h8220000;
      20325: inst = 32'h10408000;
      20326: inst = 32'hc404fd5;
      20327: inst = 32'h8220000;
      20328: inst = 32'h10408000;
      20329: inst = 32'hc404fd6;
      20330: inst = 32'h8220000;
      20331: inst = 32'h10408000;
      20332: inst = 32'hc404fd7;
      20333: inst = 32'h8220000;
      20334: inst = 32'h10408000;
      20335: inst = 32'hc404fdc;
      20336: inst = 32'h8220000;
      20337: inst = 32'h10408000;
      20338: inst = 32'hc404fdd;
      20339: inst = 32'h8220000;
      20340: inst = 32'h10408000;
      20341: inst = 32'hc404fdf;
      20342: inst = 32'h8220000;
      20343: inst = 32'h10408000;
      20344: inst = 32'hc404fe0;
      20345: inst = 32'h8220000;
      20346: inst = 32'h10408000;
      20347: inst = 32'hc404fe1;
      20348: inst = 32'h8220000;
      20349: inst = 32'h10408000;
      20350: inst = 32'hc404fe2;
      20351: inst = 32'h8220000;
      20352: inst = 32'h10408000;
      20353: inst = 32'hc404fe9;
      20354: inst = 32'h8220000;
      20355: inst = 32'h10408000;
      20356: inst = 32'hc404fea;
      20357: inst = 32'h8220000;
      20358: inst = 32'h10408000;
      20359: inst = 32'hc404fec;
      20360: inst = 32'h8220000;
      20361: inst = 32'h10408000;
      20362: inst = 32'hc404fed;
      20363: inst = 32'h8220000;
      20364: inst = 32'h10408000;
      20365: inst = 32'hc404fee;
      20366: inst = 32'h8220000;
      20367: inst = 32'h10408000;
      20368: inst = 32'hc404fef;
      20369: inst = 32'h8220000;
      20370: inst = 32'h10408000;
      20371: inst = 32'hc404ff0;
      20372: inst = 32'h8220000;
      20373: inst = 32'h10408000;
      20374: inst = 32'hc40500b;
      20375: inst = 32'h8220000;
      20376: inst = 32'h10408000;
      20377: inst = 32'hc40500c;
      20378: inst = 32'h8220000;
      20379: inst = 32'h10408000;
      20380: inst = 32'hc40501d;
      20381: inst = 32'h8220000;
      20382: inst = 32'h10408000;
      20383: inst = 32'hc40501e;
      20384: inst = 32'h8220000;
      20385: inst = 32'h10408000;
      20386: inst = 32'hc40501f;
      20387: inst = 32'h8220000;
      20388: inst = 32'h10408000;
      20389: inst = 32'hc405024;
      20390: inst = 32'h8220000;
      20391: inst = 32'h10408000;
      20392: inst = 32'hc405025;
      20393: inst = 32'h8220000;
      20394: inst = 32'h10408000;
      20395: inst = 32'hc405030;
      20396: inst = 32'h8220000;
      20397: inst = 32'h10408000;
      20398: inst = 32'hc405031;
      20399: inst = 32'h8220000;
      20400: inst = 32'h10408000;
      20401: inst = 32'hc405032;
      20402: inst = 32'h8220000;
      20403: inst = 32'h10408000;
      20404: inst = 32'hc405033;
      20405: inst = 32'h8220000;
      20406: inst = 32'h10408000;
      20407: inst = 32'hc405034;
      20408: inst = 32'h8220000;
      20409: inst = 32'h10408000;
      20410: inst = 32'hc405035;
      20411: inst = 32'h8220000;
      20412: inst = 32'h10408000;
      20413: inst = 32'hc405036;
      20414: inst = 32'h8220000;
      20415: inst = 32'h10408000;
      20416: inst = 32'hc405037;
      20417: inst = 32'h8220000;
      20418: inst = 32'h10408000;
      20419: inst = 32'hc405038;
      20420: inst = 32'h8220000;
      20421: inst = 32'h10408000;
      20422: inst = 32'hc40503c;
      20423: inst = 32'h8220000;
      20424: inst = 32'h10408000;
      20425: inst = 32'hc40503d;
      20426: inst = 32'h8220000;
      20427: inst = 32'h10408000;
      20428: inst = 32'hc405049;
      20429: inst = 32'h8220000;
      20430: inst = 32'h10408000;
      20431: inst = 32'hc40504a;
      20432: inst = 32'h8220000;
      20433: inst = 32'h10408000;
      20434: inst = 32'hc40506b;
      20435: inst = 32'h8220000;
      20436: inst = 32'h10408000;
      20437: inst = 32'hc40506c;
      20438: inst = 32'h8220000;
      20439: inst = 32'h10408000;
      20440: inst = 32'hc40506d;
      20441: inst = 32'h8220000;
      20442: inst = 32'h10408000;
      20443: inst = 32'hc40506e;
      20444: inst = 32'h8220000;
      20445: inst = 32'h10408000;
      20446: inst = 32'hc40506f;
      20447: inst = 32'h8220000;
      20448: inst = 32'h10408000;
      20449: inst = 32'hc405070;
      20450: inst = 32'h8220000;
      20451: inst = 32'h10408000;
      20452: inst = 32'hc405071;
      20453: inst = 32'h8220000;
      20454: inst = 32'h10408000;
      20455: inst = 32'hc405072;
      20456: inst = 32'h8220000;
      20457: inst = 32'h10408000;
      20458: inst = 32'hc405073;
      20459: inst = 32'h8220000;
      20460: inst = 32'h10408000;
      20461: inst = 32'hc405074;
      20462: inst = 32'h8220000;
      20463: inst = 32'h10408000;
      20464: inst = 32'hc405075;
      20465: inst = 32'h8220000;
      20466: inst = 32'h10408000;
      20467: inst = 32'hc405077;
      20468: inst = 32'h8220000;
      20469: inst = 32'h10408000;
      20470: inst = 32'hc405078;
      20471: inst = 32'h8220000;
      20472: inst = 32'h10408000;
      20473: inst = 32'hc405079;
      20474: inst = 32'h8220000;
      20475: inst = 32'h10408000;
      20476: inst = 32'hc40507a;
      20477: inst = 32'h8220000;
      20478: inst = 32'h10408000;
      20479: inst = 32'hc40507b;
      20480: inst = 32'h8220000;
      20481: inst = 32'h10408000;
      20482: inst = 32'hc40507c;
      20483: inst = 32'h8220000;
      20484: inst = 32'h10408000;
      20485: inst = 32'hc40507d;
      20486: inst = 32'h8220000;
      20487: inst = 32'h10408000;
      20488: inst = 32'hc40507e;
      20489: inst = 32'h8220000;
      20490: inst = 32'h10408000;
      20491: inst = 32'hc40507f;
      20492: inst = 32'h8220000;
      20493: inst = 32'h10408000;
      20494: inst = 32'hc405080;
      20495: inst = 32'h8220000;
      20496: inst = 32'h10408000;
      20497: inst = 32'hc405084;
      20498: inst = 32'h8220000;
      20499: inst = 32'h10408000;
      20500: inst = 32'hc405085;
      20501: inst = 32'h8220000;
      20502: inst = 32'h10408000;
      20503: inst = 32'hc405086;
      20504: inst = 32'h8220000;
      20505: inst = 32'h10408000;
      20506: inst = 32'hc405087;
      20507: inst = 32'h8220000;
      20508: inst = 32'h10408000;
      20509: inst = 32'hc405088;
      20510: inst = 32'h8220000;
      20511: inst = 32'h10408000;
      20512: inst = 32'hc405089;
      20513: inst = 32'h8220000;
      20514: inst = 32'h10408000;
      20515: inst = 32'hc40508a;
      20516: inst = 32'h8220000;
      20517: inst = 32'h10408000;
      20518: inst = 32'hc40508b;
      20519: inst = 32'h8220000;
      20520: inst = 32'h10408000;
      20521: inst = 32'hc40508c;
      20522: inst = 32'h8220000;
      20523: inst = 32'h10408000;
      20524: inst = 32'hc40508d;
      20525: inst = 32'h8220000;
      20526: inst = 32'h10408000;
      20527: inst = 32'hc405090;
      20528: inst = 32'h8220000;
      20529: inst = 32'h10408000;
      20530: inst = 32'hc405091;
      20531: inst = 32'h8220000;
      20532: inst = 32'h10408000;
      20533: inst = 32'hc405096;
      20534: inst = 32'h8220000;
      20535: inst = 32'h10408000;
      20536: inst = 32'hc405097;
      20537: inst = 32'h8220000;
      20538: inst = 32'h10408000;
      20539: inst = 32'hc405098;
      20540: inst = 32'h8220000;
      20541: inst = 32'h10408000;
      20542: inst = 32'hc405099;
      20543: inst = 32'h8220000;
      20544: inst = 32'h10408000;
      20545: inst = 32'hc40509c;
      20546: inst = 32'h8220000;
      20547: inst = 32'h10408000;
      20548: inst = 32'hc40509d;
      20549: inst = 32'h8220000;
      20550: inst = 32'h10408000;
      20551: inst = 32'hc4050a9;
      20552: inst = 32'h8220000;
      20553: inst = 32'h10408000;
      20554: inst = 32'hc4050aa;
      20555: inst = 32'h8220000;
      20556: inst = 32'h10408000;
      20557: inst = 32'hc4050ab;
      20558: inst = 32'h8220000;
      20559: inst = 32'h10408000;
      20560: inst = 32'hc4050ac;
      20561: inst = 32'h8220000;
      20562: inst = 32'h10408000;
      20563: inst = 32'hc4050ad;
      20564: inst = 32'h8220000;
      20565: inst = 32'h10408000;
      20566: inst = 32'hc4050ae;
      20567: inst = 32'h8220000;
      20568: inst = 32'h10408000;
      20569: inst = 32'hc4050af;
      20570: inst = 32'h8220000;
      20571: inst = 32'h10408000;
      20572: inst = 32'hc4050b0;
      20573: inst = 32'h8220000;
      20574: inst = 32'h10408000;
      20575: inst = 32'hc4050b1;
      20576: inst = 32'h8220000;
      20577: inst = 32'h10408000;
      20578: inst = 32'hc4050b2;
      20579: inst = 32'h8220000;
      20580: inst = 32'h10408000;
      20581: inst = 32'hc4050b3;
      20582: inst = 32'h8220000;
      20583: inst = 32'h10408000;
      20584: inst = 32'hc4050cb;
      20585: inst = 32'h8220000;
      20586: inst = 32'h10408000;
      20587: inst = 32'hc4050cc;
      20588: inst = 32'h8220000;
      20589: inst = 32'h10408000;
      20590: inst = 32'hc4050cd;
      20591: inst = 32'h8220000;
      20592: inst = 32'h10408000;
      20593: inst = 32'hc4050ce;
      20594: inst = 32'h8220000;
      20595: inst = 32'h10408000;
      20596: inst = 32'hc4050cf;
      20597: inst = 32'h8220000;
      20598: inst = 32'h10408000;
      20599: inst = 32'hc4050d0;
      20600: inst = 32'h8220000;
      20601: inst = 32'h10408000;
      20602: inst = 32'hc4050d1;
      20603: inst = 32'h8220000;
      20604: inst = 32'h10408000;
      20605: inst = 32'hc4050d2;
      20606: inst = 32'h8220000;
      20607: inst = 32'h10408000;
      20608: inst = 32'hc4050d3;
      20609: inst = 32'h8220000;
      20610: inst = 32'h10408000;
      20611: inst = 32'hc4050d4;
      20612: inst = 32'h8220000;
      20613: inst = 32'h10408000;
      20614: inst = 32'hc4050d7;
      20615: inst = 32'h8220000;
      20616: inst = 32'h10408000;
      20617: inst = 32'hc4050d8;
      20618: inst = 32'h8220000;
      20619: inst = 32'h10408000;
      20620: inst = 32'hc4050d9;
      20621: inst = 32'h8220000;
      20622: inst = 32'h10408000;
      20623: inst = 32'hc4050da;
      20624: inst = 32'h8220000;
      20625: inst = 32'h10408000;
      20626: inst = 32'hc4050db;
      20627: inst = 32'h8220000;
      20628: inst = 32'h10408000;
      20629: inst = 32'hc4050dc;
      20630: inst = 32'h8220000;
      20631: inst = 32'h10408000;
      20632: inst = 32'hc4050dd;
      20633: inst = 32'h8220000;
      20634: inst = 32'h10408000;
      20635: inst = 32'hc4050de;
      20636: inst = 32'h8220000;
      20637: inst = 32'h10408000;
      20638: inst = 32'hc4050df;
      20639: inst = 32'h8220000;
      20640: inst = 32'h10408000;
      20641: inst = 32'hc4050e0;
      20642: inst = 32'h8220000;
      20643: inst = 32'h10408000;
      20644: inst = 32'hc4050e1;
      20645: inst = 32'h8220000;
      20646: inst = 32'h10408000;
      20647: inst = 32'hc4050e5;
      20648: inst = 32'h8220000;
      20649: inst = 32'h10408000;
      20650: inst = 32'hc4050e6;
      20651: inst = 32'h8220000;
      20652: inst = 32'h10408000;
      20653: inst = 32'hc4050e7;
      20654: inst = 32'h8220000;
      20655: inst = 32'h10408000;
      20656: inst = 32'hc4050e8;
      20657: inst = 32'h8220000;
      20658: inst = 32'h10408000;
      20659: inst = 32'hc4050e9;
      20660: inst = 32'h8220000;
      20661: inst = 32'h10408000;
      20662: inst = 32'hc4050ea;
      20663: inst = 32'h8220000;
      20664: inst = 32'h10408000;
      20665: inst = 32'hc4050eb;
      20666: inst = 32'h8220000;
      20667: inst = 32'h10408000;
      20668: inst = 32'hc4050ec;
      20669: inst = 32'h8220000;
      20670: inst = 32'h10408000;
      20671: inst = 32'hc4050ed;
      20672: inst = 32'h8220000;
      20673: inst = 32'h10408000;
      20674: inst = 32'hc4050f0;
      20675: inst = 32'h8220000;
      20676: inst = 32'h10408000;
      20677: inst = 32'hc4050f1;
      20678: inst = 32'h8220000;
      20679: inst = 32'h10408000;
      20680: inst = 32'hc4050f6;
      20681: inst = 32'h8220000;
      20682: inst = 32'h10408000;
      20683: inst = 32'hc4050f7;
      20684: inst = 32'h8220000;
      20685: inst = 32'h10408000;
      20686: inst = 32'hc4050f8;
      20687: inst = 32'h8220000;
      20688: inst = 32'h10408000;
      20689: inst = 32'hc4050f9;
      20690: inst = 32'h8220000;
      20691: inst = 32'h10408000;
      20692: inst = 32'hc4050fa;
      20693: inst = 32'h8220000;
      20694: inst = 32'h10408000;
      20695: inst = 32'hc4050fc;
      20696: inst = 32'h8220000;
      20697: inst = 32'h10408000;
      20698: inst = 32'hc4050fd;
      20699: inst = 32'h8220000;
      20700: inst = 32'h10408000;
      20701: inst = 32'hc405109;
      20702: inst = 32'h8220000;
      20703: inst = 32'h10408000;
      20704: inst = 32'hc40510a;
      20705: inst = 32'h8220000;
      20706: inst = 32'h10408000;
      20707: inst = 32'hc40510b;
      20708: inst = 32'h8220000;
      20709: inst = 32'h10408000;
      20710: inst = 32'hc40510c;
      20711: inst = 32'h8220000;
      20712: inst = 32'h10408000;
      20713: inst = 32'hc40510d;
      20714: inst = 32'h8220000;
      20715: inst = 32'h10408000;
      20716: inst = 32'hc40510e;
      20717: inst = 32'h8220000;
      20718: inst = 32'h10408000;
      20719: inst = 32'hc40510f;
      20720: inst = 32'h8220000;
      20721: inst = 32'h10408000;
      20722: inst = 32'hc405110;
      20723: inst = 32'h8220000;
      20724: inst = 32'h10408000;
      20725: inst = 32'hc405111;
      20726: inst = 32'h8220000;
      20727: inst = 32'h10408000;
      20728: inst = 32'hc405112;
      20729: inst = 32'h8220000;
      20730: inst = 32'h10408000;
      20731: inst = 32'hc405113;
      20732: inst = 32'h8220000;
      20733: inst = 32'h58000000;
      20734: inst = 32'hc20529c;
      20735: inst = 32'h10408000;
      20736: inst = 32'hc404224;
      20737: inst = 32'h8220000;
      20738: inst = 32'h10408000;
      20739: inst = 32'hc404225;
      20740: inst = 32'h8220000;
      20741: inst = 32'h10408000;
      20742: inst = 32'hc404226;
      20743: inst = 32'h8220000;
      20744: inst = 32'h10408000;
      20745: inst = 32'hc404227;
      20746: inst = 32'h8220000;
      20747: inst = 32'h10408000;
      20748: inst = 32'hc404228;
      20749: inst = 32'h8220000;
      20750: inst = 32'h10408000;
      20751: inst = 32'hc404229;
      20752: inst = 32'h8220000;
      20753: inst = 32'h10408000;
      20754: inst = 32'hc40422a;
      20755: inst = 32'h8220000;
      20756: inst = 32'h10408000;
      20757: inst = 32'hc40422b;
      20758: inst = 32'h8220000;
      20759: inst = 32'h10408000;
      20760: inst = 32'hc40422c;
      20761: inst = 32'h8220000;
      20762: inst = 32'h10408000;
      20763: inst = 32'hc40422d;
      20764: inst = 32'h8220000;
      20765: inst = 32'h10408000;
      20766: inst = 32'hc40422e;
      20767: inst = 32'h8220000;
      20768: inst = 32'h10408000;
      20769: inst = 32'hc40422f;
      20770: inst = 32'h8220000;
      20771: inst = 32'h10408000;
      20772: inst = 32'hc404230;
      20773: inst = 32'h8220000;
      20774: inst = 32'h10408000;
      20775: inst = 32'hc404231;
      20776: inst = 32'h8220000;
      20777: inst = 32'h10408000;
      20778: inst = 32'hc404232;
      20779: inst = 32'h8220000;
      20780: inst = 32'h10408000;
      20781: inst = 32'hc404233;
      20782: inst = 32'h8220000;
      20783: inst = 32'h10408000;
      20784: inst = 32'hc404234;
      20785: inst = 32'h8220000;
      20786: inst = 32'h10408000;
      20787: inst = 32'hc404235;
      20788: inst = 32'h8220000;
      20789: inst = 32'h10408000;
      20790: inst = 32'hc404236;
      20791: inst = 32'h8220000;
      20792: inst = 32'h10408000;
      20793: inst = 32'hc404237;
      20794: inst = 32'h8220000;
      20795: inst = 32'h10408000;
      20796: inst = 32'hc404238;
      20797: inst = 32'h8220000;
      20798: inst = 32'h10408000;
      20799: inst = 32'hc404239;
      20800: inst = 32'h8220000;
      20801: inst = 32'h10408000;
      20802: inst = 32'hc40423a;
      20803: inst = 32'h8220000;
      20804: inst = 32'h10408000;
      20805: inst = 32'hc40423b;
      20806: inst = 32'h8220000;
      20807: inst = 32'h10408000;
      20808: inst = 32'hc40423c;
      20809: inst = 32'h8220000;
      20810: inst = 32'h10408000;
      20811: inst = 32'hc40423d;
      20812: inst = 32'h8220000;
      20813: inst = 32'h10408000;
      20814: inst = 32'hc40423e;
      20815: inst = 32'h8220000;
      20816: inst = 32'h10408000;
      20817: inst = 32'hc40423f;
      20818: inst = 32'h8220000;
      20819: inst = 32'h10408000;
      20820: inst = 32'hc404240;
      20821: inst = 32'h8220000;
      20822: inst = 32'h10408000;
      20823: inst = 32'hc404241;
      20824: inst = 32'h8220000;
      20825: inst = 32'h10408000;
      20826: inst = 32'hc404242;
      20827: inst = 32'h8220000;
      20828: inst = 32'h10408000;
      20829: inst = 32'hc404243;
      20830: inst = 32'h8220000;
      20831: inst = 32'h10408000;
      20832: inst = 32'hc404244;
      20833: inst = 32'h8220000;
      20834: inst = 32'h10408000;
      20835: inst = 32'hc404245;
      20836: inst = 32'h8220000;
      20837: inst = 32'h10408000;
      20838: inst = 32'hc404246;
      20839: inst = 32'h8220000;
      20840: inst = 32'h10408000;
      20841: inst = 32'hc404247;
      20842: inst = 32'h8220000;
      20843: inst = 32'h10408000;
      20844: inst = 32'hc404248;
      20845: inst = 32'h8220000;
      20846: inst = 32'h10408000;
      20847: inst = 32'hc404249;
      20848: inst = 32'h8220000;
      20849: inst = 32'h10408000;
      20850: inst = 32'hc40424a;
      20851: inst = 32'h8220000;
      20852: inst = 32'h10408000;
      20853: inst = 32'hc40424b;
      20854: inst = 32'h8220000;
      20855: inst = 32'h10408000;
      20856: inst = 32'hc40424c;
      20857: inst = 32'h8220000;
      20858: inst = 32'h10408000;
      20859: inst = 32'hc40424d;
      20860: inst = 32'h8220000;
      20861: inst = 32'h10408000;
      20862: inst = 32'hc40424e;
      20863: inst = 32'h8220000;
      20864: inst = 32'h10408000;
      20865: inst = 32'hc40424f;
      20866: inst = 32'h8220000;
      20867: inst = 32'h10408000;
      20868: inst = 32'hc404250;
      20869: inst = 32'h8220000;
      20870: inst = 32'h10408000;
      20871: inst = 32'hc404251;
      20872: inst = 32'h8220000;
      20873: inst = 32'h10408000;
      20874: inst = 32'hc404252;
      20875: inst = 32'h8220000;
      20876: inst = 32'h10408000;
      20877: inst = 32'hc404253;
      20878: inst = 32'h8220000;
      20879: inst = 32'h10408000;
      20880: inst = 32'hc404254;
      20881: inst = 32'h8220000;
      20882: inst = 32'h10408000;
      20883: inst = 32'hc404255;
      20884: inst = 32'h8220000;
      20885: inst = 32'h10408000;
      20886: inst = 32'hc404256;
      20887: inst = 32'h8220000;
      20888: inst = 32'h10408000;
      20889: inst = 32'hc404257;
      20890: inst = 32'h8220000;
      20891: inst = 32'h10408000;
      20892: inst = 32'hc404258;
      20893: inst = 32'h8220000;
      20894: inst = 32'h10408000;
      20895: inst = 32'hc404259;
      20896: inst = 32'h8220000;
      20897: inst = 32'h10408000;
      20898: inst = 32'hc40425a;
      20899: inst = 32'h8220000;
      20900: inst = 32'h10408000;
      20901: inst = 32'hc40425b;
      20902: inst = 32'h8220000;
      20903: inst = 32'h10408000;
      20904: inst = 32'hc40425c;
      20905: inst = 32'h8220000;
      20906: inst = 32'h10408000;
      20907: inst = 32'hc40425d;
      20908: inst = 32'h8220000;
      20909: inst = 32'h10408000;
      20910: inst = 32'hc40425e;
      20911: inst = 32'h8220000;
      20912: inst = 32'h10408000;
      20913: inst = 32'hc40425f;
      20914: inst = 32'h8220000;
      20915: inst = 32'h10408000;
      20916: inst = 32'hc404260;
      20917: inst = 32'h8220000;
      20918: inst = 32'h10408000;
      20919: inst = 32'hc404261;
      20920: inst = 32'h8220000;
      20921: inst = 32'h10408000;
      20922: inst = 32'hc404262;
      20923: inst = 32'h8220000;
      20924: inst = 32'h10408000;
      20925: inst = 32'hc404263;
      20926: inst = 32'h8220000;
      20927: inst = 32'h10408000;
      20928: inst = 32'hc404264;
      20929: inst = 32'h8220000;
      20930: inst = 32'h10408000;
      20931: inst = 32'hc404265;
      20932: inst = 32'h8220000;
      20933: inst = 32'h10408000;
      20934: inst = 32'hc404266;
      20935: inst = 32'h8220000;
      20936: inst = 32'h10408000;
      20937: inst = 32'hc404267;
      20938: inst = 32'h8220000;
      20939: inst = 32'h10408000;
      20940: inst = 32'hc404268;
      20941: inst = 32'h8220000;
      20942: inst = 32'h10408000;
      20943: inst = 32'hc404269;
      20944: inst = 32'h8220000;
      20945: inst = 32'h10408000;
      20946: inst = 32'hc40426a;
      20947: inst = 32'h8220000;
      20948: inst = 32'h10408000;
      20949: inst = 32'hc40426b;
      20950: inst = 32'h8220000;
      20951: inst = 32'h10408000;
      20952: inst = 32'hc40426c;
      20953: inst = 32'h8220000;
      20954: inst = 32'h10408000;
      20955: inst = 32'hc40426d;
      20956: inst = 32'h8220000;
      20957: inst = 32'h10408000;
      20958: inst = 32'hc40426e;
      20959: inst = 32'h8220000;
      20960: inst = 32'h10408000;
      20961: inst = 32'hc40426f;
      20962: inst = 32'h8220000;
      20963: inst = 32'h10408000;
      20964: inst = 32'hc404270;
      20965: inst = 32'h8220000;
      20966: inst = 32'h10408000;
      20967: inst = 32'hc404271;
      20968: inst = 32'h8220000;
      20969: inst = 32'h10408000;
      20970: inst = 32'hc404272;
      20971: inst = 32'h8220000;
      20972: inst = 32'h10408000;
      20973: inst = 32'hc404273;
      20974: inst = 32'h8220000;
      20975: inst = 32'h10408000;
      20976: inst = 32'hc404274;
      20977: inst = 32'h8220000;
      20978: inst = 32'h10408000;
      20979: inst = 32'hc404275;
      20980: inst = 32'h8220000;
      20981: inst = 32'h10408000;
      20982: inst = 32'hc404276;
      20983: inst = 32'h8220000;
      20984: inst = 32'h10408000;
      20985: inst = 32'hc404277;
      20986: inst = 32'h8220000;
      20987: inst = 32'h10408000;
      20988: inst = 32'hc404278;
      20989: inst = 32'h8220000;
      20990: inst = 32'h10408000;
      20991: inst = 32'hc404279;
      20992: inst = 32'h8220000;
      20993: inst = 32'h10408000;
      20994: inst = 32'hc40427a;
      20995: inst = 32'h8220000;
      20996: inst = 32'h10408000;
      20997: inst = 32'hc40427b;
      20998: inst = 32'h8220000;
      20999: inst = 32'h10408000;
      21000: inst = 32'hc404284;
      21001: inst = 32'h8220000;
      21002: inst = 32'h10408000;
      21003: inst = 32'hc404285;
      21004: inst = 32'h8220000;
      21005: inst = 32'h10408000;
      21006: inst = 32'hc404286;
      21007: inst = 32'h8220000;
      21008: inst = 32'h10408000;
      21009: inst = 32'hc404287;
      21010: inst = 32'h8220000;
      21011: inst = 32'h10408000;
      21012: inst = 32'hc404288;
      21013: inst = 32'h8220000;
      21014: inst = 32'h10408000;
      21015: inst = 32'hc404289;
      21016: inst = 32'h8220000;
      21017: inst = 32'h10408000;
      21018: inst = 32'hc40428a;
      21019: inst = 32'h8220000;
      21020: inst = 32'h10408000;
      21021: inst = 32'hc40428b;
      21022: inst = 32'h8220000;
      21023: inst = 32'h10408000;
      21024: inst = 32'hc40428c;
      21025: inst = 32'h8220000;
      21026: inst = 32'h10408000;
      21027: inst = 32'hc40428d;
      21028: inst = 32'h8220000;
      21029: inst = 32'h10408000;
      21030: inst = 32'hc40428e;
      21031: inst = 32'h8220000;
      21032: inst = 32'h10408000;
      21033: inst = 32'hc40428f;
      21034: inst = 32'h8220000;
      21035: inst = 32'h10408000;
      21036: inst = 32'hc404290;
      21037: inst = 32'h8220000;
      21038: inst = 32'h10408000;
      21039: inst = 32'hc404291;
      21040: inst = 32'h8220000;
      21041: inst = 32'h10408000;
      21042: inst = 32'hc404292;
      21043: inst = 32'h8220000;
      21044: inst = 32'h10408000;
      21045: inst = 32'hc404293;
      21046: inst = 32'h8220000;
      21047: inst = 32'h10408000;
      21048: inst = 32'hc404294;
      21049: inst = 32'h8220000;
      21050: inst = 32'h10408000;
      21051: inst = 32'hc404295;
      21052: inst = 32'h8220000;
      21053: inst = 32'h10408000;
      21054: inst = 32'hc404296;
      21055: inst = 32'h8220000;
      21056: inst = 32'h10408000;
      21057: inst = 32'hc404297;
      21058: inst = 32'h8220000;
      21059: inst = 32'h10408000;
      21060: inst = 32'hc404298;
      21061: inst = 32'h8220000;
      21062: inst = 32'h10408000;
      21063: inst = 32'hc404299;
      21064: inst = 32'h8220000;
      21065: inst = 32'h10408000;
      21066: inst = 32'hc40429a;
      21067: inst = 32'h8220000;
      21068: inst = 32'h10408000;
      21069: inst = 32'hc40429b;
      21070: inst = 32'h8220000;
      21071: inst = 32'h10408000;
      21072: inst = 32'hc40429c;
      21073: inst = 32'h8220000;
      21074: inst = 32'h10408000;
      21075: inst = 32'hc40429d;
      21076: inst = 32'h8220000;
      21077: inst = 32'h10408000;
      21078: inst = 32'hc40429e;
      21079: inst = 32'h8220000;
      21080: inst = 32'h10408000;
      21081: inst = 32'hc40429f;
      21082: inst = 32'h8220000;
      21083: inst = 32'h10408000;
      21084: inst = 32'hc4042a0;
      21085: inst = 32'h8220000;
      21086: inst = 32'h10408000;
      21087: inst = 32'hc4042a1;
      21088: inst = 32'h8220000;
      21089: inst = 32'h10408000;
      21090: inst = 32'hc4042a2;
      21091: inst = 32'h8220000;
      21092: inst = 32'h10408000;
      21093: inst = 32'hc4042a3;
      21094: inst = 32'h8220000;
      21095: inst = 32'h10408000;
      21096: inst = 32'hc4042a4;
      21097: inst = 32'h8220000;
      21098: inst = 32'h10408000;
      21099: inst = 32'hc4042a5;
      21100: inst = 32'h8220000;
      21101: inst = 32'h10408000;
      21102: inst = 32'hc4042a6;
      21103: inst = 32'h8220000;
      21104: inst = 32'h10408000;
      21105: inst = 32'hc4042a7;
      21106: inst = 32'h8220000;
      21107: inst = 32'h10408000;
      21108: inst = 32'hc4042a8;
      21109: inst = 32'h8220000;
      21110: inst = 32'h10408000;
      21111: inst = 32'hc4042a9;
      21112: inst = 32'h8220000;
      21113: inst = 32'h10408000;
      21114: inst = 32'hc4042aa;
      21115: inst = 32'h8220000;
      21116: inst = 32'h10408000;
      21117: inst = 32'hc4042ab;
      21118: inst = 32'h8220000;
      21119: inst = 32'h10408000;
      21120: inst = 32'hc4042ac;
      21121: inst = 32'h8220000;
      21122: inst = 32'h10408000;
      21123: inst = 32'hc4042ad;
      21124: inst = 32'h8220000;
      21125: inst = 32'h10408000;
      21126: inst = 32'hc4042ae;
      21127: inst = 32'h8220000;
      21128: inst = 32'h10408000;
      21129: inst = 32'hc4042af;
      21130: inst = 32'h8220000;
      21131: inst = 32'h10408000;
      21132: inst = 32'hc4042b0;
      21133: inst = 32'h8220000;
      21134: inst = 32'h10408000;
      21135: inst = 32'hc4042b1;
      21136: inst = 32'h8220000;
      21137: inst = 32'h10408000;
      21138: inst = 32'hc4042b2;
      21139: inst = 32'h8220000;
      21140: inst = 32'h10408000;
      21141: inst = 32'hc4042b3;
      21142: inst = 32'h8220000;
      21143: inst = 32'h10408000;
      21144: inst = 32'hc4042b4;
      21145: inst = 32'h8220000;
      21146: inst = 32'h10408000;
      21147: inst = 32'hc4042b5;
      21148: inst = 32'h8220000;
      21149: inst = 32'h10408000;
      21150: inst = 32'hc4042b6;
      21151: inst = 32'h8220000;
      21152: inst = 32'h10408000;
      21153: inst = 32'hc4042b7;
      21154: inst = 32'h8220000;
      21155: inst = 32'h10408000;
      21156: inst = 32'hc4042b8;
      21157: inst = 32'h8220000;
      21158: inst = 32'h10408000;
      21159: inst = 32'hc4042b9;
      21160: inst = 32'h8220000;
      21161: inst = 32'h10408000;
      21162: inst = 32'hc4042ba;
      21163: inst = 32'h8220000;
      21164: inst = 32'h10408000;
      21165: inst = 32'hc4042bb;
      21166: inst = 32'h8220000;
      21167: inst = 32'h10408000;
      21168: inst = 32'hc4042bc;
      21169: inst = 32'h8220000;
      21170: inst = 32'h10408000;
      21171: inst = 32'hc4042bd;
      21172: inst = 32'h8220000;
      21173: inst = 32'h10408000;
      21174: inst = 32'hc4042be;
      21175: inst = 32'h8220000;
      21176: inst = 32'h10408000;
      21177: inst = 32'hc4042bf;
      21178: inst = 32'h8220000;
      21179: inst = 32'h10408000;
      21180: inst = 32'hc4042c0;
      21181: inst = 32'h8220000;
      21182: inst = 32'h10408000;
      21183: inst = 32'hc4042c1;
      21184: inst = 32'h8220000;
      21185: inst = 32'h10408000;
      21186: inst = 32'hc4042c2;
      21187: inst = 32'h8220000;
      21188: inst = 32'h10408000;
      21189: inst = 32'hc4042c3;
      21190: inst = 32'h8220000;
      21191: inst = 32'h10408000;
      21192: inst = 32'hc4042c4;
      21193: inst = 32'h8220000;
      21194: inst = 32'h10408000;
      21195: inst = 32'hc4042c5;
      21196: inst = 32'h8220000;
      21197: inst = 32'h10408000;
      21198: inst = 32'hc4042c6;
      21199: inst = 32'h8220000;
      21200: inst = 32'h10408000;
      21201: inst = 32'hc4042c7;
      21202: inst = 32'h8220000;
      21203: inst = 32'h10408000;
      21204: inst = 32'hc4042c8;
      21205: inst = 32'h8220000;
      21206: inst = 32'h10408000;
      21207: inst = 32'hc4042c9;
      21208: inst = 32'h8220000;
      21209: inst = 32'h10408000;
      21210: inst = 32'hc4042ca;
      21211: inst = 32'h8220000;
      21212: inst = 32'h10408000;
      21213: inst = 32'hc4042cb;
      21214: inst = 32'h8220000;
      21215: inst = 32'h10408000;
      21216: inst = 32'hc4042cc;
      21217: inst = 32'h8220000;
      21218: inst = 32'h10408000;
      21219: inst = 32'hc4042cd;
      21220: inst = 32'h8220000;
      21221: inst = 32'h10408000;
      21222: inst = 32'hc4042ce;
      21223: inst = 32'h8220000;
      21224: inst = 32'h10408000;
      21225: inst = 32'hc4042cf;
      21226: inst = 32'h8220000;
      21227: inst = 32'h10408000;
      21228: inst = 32'hc4042d0;
      21229: inst = 32'h8220000;
      21230: inst = 32'h10408000;
      21231: inst = 32'hc4042d1;
      21232: inst = 32'h8220000;
      21233: inst = 32'h10408000;
      21234: inst = 32'hc4042d2;
      21235: inst = 32'h8220000;
      21236: inst = 32'h10408000;
      21237: inst = 32'hc4042d3;
      21238: inst = 32'h8220000;
      21239: inst = 32'h10408000;
      21240: inst = 32'hc4042d4;
      21241: inst = 32'h8220000;
      21242: inst = 32'h10408000;
      21243: inst = 32'hc4042d5;
      21244: inst = 32'h8220000;
      21245: inst = 32'h10408000;
      21246: inst = 32'hc4042d6;
      21247: inst = 32'h8220000;
      21248: inst = 32'h10408000;
      21249: inst = 32'hc4042d7;
      21250: inst = 32'h8220000;
      21251: inst = 32'h10408000;
      21252: inst = 32'hc4042d8;
      21253: inst = 32'h8220000;
      21254: inst = 32'h10408000;
      21255: inst = 32'hc4042d9;
      21256: inst = 32'h8220000;
      21257: inst = 32'h10408000;
      21258: inst = 32'hc4042da;
      21259: inst = 32'h8220000;
      21260: inst = 32'h10408000;
      21261: inst = 32'hc4042db;
      21262: inst = 32'h8220000;
      21263: inst = 32'h10408000;
      21264: inst = 32'hc4042e4;
      21265: inst = 32'h8220000;
      21266: inst = 32'h10408000;
      21267: inst = 32'hc4042e5;
      21268: inst = 32'h8220000;
      21269: inst = 32'h10408000;
      21270: inst = 32'hc4042e6;
      21271: inst = 32'h8220000;
      21272: inst = 32'h10408000;
      21273: inst = 32'hc404339;
      21274: inst = 32'h8220000;
      21275: inst = 32'h10408000;
      21276: inst = 32'hc40433a;
      21277: inst = 32'h8220000;
      21278: inst = 32'h10408000;
      21279: inst = 32'hc40433b;
      21280: inst = 32'h8220000;
      21281: inst = 32'h10408000;
      21282: inst = 32'hc404344;
      21283: inst = 32'h8220000;
      21284: inst = 32'h10408000;
      21285: inst = 32'hc404345;
      21286: inst = 32'h8220000;
      21287: inst = 32'h10408000;
      21288: inst = 32'hc40439a;
      21289: inst = 32'h8220000;
      21290: inst = 32'h10408000;
      21291: inst = 32'hc40439b;
      21292: inst = 32'h8220000;
      21293: inst = 32'h10408000;
      21294: inst = 32'hc4043a4;
      21295: inst = 32'h8220000;
      21296: inst = 32'h10408000;
      21297: inst = 32'hc4043a5;
      21298: inst = 32'h8220000;
      21299: inst = 32'h10408000;
      21300: inst = 32'hc4043fa;
      21301: inst = 32'h8220000;
      21302: inst = 32'h10408000;
      21303: inst = 32'hc4043fb;
      21304: inst = 32'h8220000;
      21305: inst = 32'h10408000;
      21306: inst = 32'hc404404;
      21307: inst = 32'h8220000;
      21308: inst = 32'h10408000;
      21309: inst = 32'hc404405;
      21310: inst = 32'h8220000;
      21311: inst = 32'h10408000;
      21312: inst = 32'hc40445a;
      21313: inst = 32'h8220000;
      21314: inst = 32'h10408000;
      21315: inst = 32'hc40445b;
      21316: inst = 32'h8220000;
      21317: inst = 32'h10408000;
      21318: inst = 32'hc404464;
      21319: inst = 32'h8220000;
      21320: inst = 32'h10408000;
      21321: inst = 32'hc404465;
      21322: inst = 32'h8220000;
      21323: inst = 32'h10408000;
      21324: inst = 32'hc4044ba;
      21325: inst = 32'h8220000;
      21326: inst = 32'h10408000;
      21327: inst = 32'hc4044bb;
      21328: inst = 32'h8220000;
      21329: inst = 32'h10408000;
      21330: inst = 32'hc4044c4;
      21331: inst = 32'h8220000;
      21332: inst = 32'h10408000;
      21333: inst = 32'hc4044c5;
      21334: inst = 32'h8220000;
      21335: inst = 32'h10408000;
      21336: inst = 32'hc40451a;
      21337: inst = 32'h8220000;
      21338: inst = 32'h10408000;
      21339: inst = 32'hc40451b;
      21340: inst = 32'h8220000;
      21341: inst = 32'h10408000;
      21342: inst = 32'hc404524;
      21343: inst = 32'h8220000;
      21344: inst = 32'h10408000;
      21345: inst = 32'hc404525;
      21346: inst = 32'h8220000;
      21347: inst = 32'h10408000;
      21348: inst = 32'hc40457a;
      21349: inst = 32'h8220000;
      21350: inst = 32'h10408000;
      21351: inst = 32'hc40457b;
      21352: inst = 32'h8220000;
      21353: inst = 32'h10408000;
      21354: inst = 32'hc404584;
      21355: inst = 32'h8220000;
      21356: inst = 32'h10408000;
      21357: inst = 32'hc404585;
      21358: inst = 32'h8220000;
      21359: inst = 32'h10408000;
      21360: inst = 32'hc4045da;
      21361: inst = 32'h8220000;
      21362: inst = 32'h10408000;
      21363: inst = 32'hc4045db;
      21364: inst = 32'h8220000;
      21365: inst = 32'h10408000;
      21366: inst = 32'hc4045e4;
      21367: inst = 32'h8220000;
      21368: inst = 32'h10408000;
      21369: inst = 32'hc4045e5;
      21370: inst = 32'h8220000;
      21371: inst = 32'h10408000;
      21372: inst = 32'hc40463a;
      21373: inst = 32'h8220000;
      21374: inst = 32'h10408000;
      21375: inst = 32'hc40463b;
      21376: inst = 32'h8220000;
      21377: inst = 32'h10408000;
      21378: inst = 32'hc404644;
      21379: inst = 32'h8220000;
      21380: inst = 32'h10408000;
      21381: inst = 32'hc404645;
      21382: inst = 32'h8220000;
      21383: inst = 32'h10408000;
      21384: inst = 32'hc40469a;
      21385: inst = 32'h8220000;
      21386: inst = 32'h10408000;
      21387: inst = 32'hc40469b;
      21388: inst = 32'h8220000;
      21389: inst = 32'h10408000;
      21390: inst = 32'hc4046a4;
      21391: inst = 32'h8220000;
      21392: inst = 32'h10408000;
      21393: inst = 32'hc4046a5;
      21394: inst = 32'h8220000;
      21395: inst = 32'h10408000;
      21396: inst = 32'hc4046fa;
      21397: inst = 32'h8220000;
      21398: inst = 32'h10408000;
      21399: inst = 32'hc4046fb;
      21400: inst = 32'h8220000;
      21401: inst = 32'h10408000;
      21402: inst = 32'hc404704;
      21403: inst = 32'h8220000;
      21404: inst = 32'h10408000;
      21405: inst = 32'hc404705;
      21406: inst = 32'h8220000;
      21407: inst = 32'h10408000;
      21408: inst = 32'hc40475a;
      21409: inst = 32'h8220000;
      21410: inst = 32'h10408000;
      21411: inst = 32'hc40475b;
      21412: inst = 32'h8220000;
      21413: inst = 32'h10408000;
      21414: inst = 32'hc404764;
      21415: inst = 32'h8220000;
      21416: inst = 32'h10408000;
      21417: inst = 32'hc404765;
      21418: inst = 32'h8220000;
      21419: inst = 32'h10408000;
      21420: inst = 32'hc4047ba;
      21421: inst = 32'h8220000;
      21422: inst = 32'h10408000;
      21423: inst = 32'hc4047bb;
      21424: inst = 32'h8220000;
      21425: inst = 32'h10408000;
      21426: inst = 32'hc4047c4;
      21427: inst = 32'h8220000;
      21428: inst = 32'h10408000;
      21429: inst = 32'hc4047c5;
      21430: inst = 32'h8220000;
      21431: inst = 32'h10408000;
      21432: inst = 32'hc40481a;
      21433: inst = 32'h8220000;
      21434: inst = 32'h10408000;
      21435: inst = 32'hc40481b;
      21436: inst = 32'h8220000;
      21437: inst = 32'h10408000;
      21438: inst = 32'hc404824;
      21439: inst = 32'h8220000;
      21440: inst = 32'h10408000;
      21441: inst = 32'hc404825;
      21442: inst = 32'h8220000;
      21443: inst = 32'h10408000;
      21444: inst = 32'hc40487a;
      21445: inst = 32'h8220000;
      21446: inst = 32'h10408000;
      21447: inst = 32'hc40487b;
      21448: inst = 32'h8220000;
      21449: inst = 32'h10408000;
      21450: inst = 32'hc404884;
      21451: inst = 32'h8220000;
      21452: inst = 32'h10408000;
      21453: inst = 32'hc404885;
      21454: inst = 32'h8220000;
      21455: inst = 32'h10408000;
      21456: inst = 32'hc4048da;
      21457: inst = 32'h8220000;
      21458: inst = 32'h10408000;
      21459: inst = 32'hc4048db;
      21460: inst = 32'h8220000;
      21461: inst = 32'h10408000;
      21462: inst = 32'hc4048e4;
      21463: inst = 32'h8220000;
      21464: inst = 32'h10408000;
      21465: inst = 32'hc4048e5;
      21466: inst = 32'h8220000;
      21467: inst = 32'h10408000;
      21468: inst = 32'hc40493a;
      21469: inst = 32'h8220000;
      21470: inst = 32'h10408000;
      21471: inst = 32'hc40493b;
      21472: inst = 32'h8220000;
      21473: inst = 32'h10408000;
      21474: inst = 32'hc404944;
      21475: inst = 32'h8220000;
      21476: inst = 32'h10408000;
      21477: inst = 32'hc404945;
      21478: inst = 32'h8220000;
      21479: inst = 32'h10408000;
      21480: inst = 32'hc40499a;
      21481: inst = 32'h8220000;
      21482: inst = 32'h10408000;
      21483: inst = 32'hc40499b;
      21484: inst = 32'h8220000;
      21485: inst = 32'h10408000;
      21486: inst = 32'hc4049a4;
      21487: inst = 32'h8220000;
      21488: inst = 32'h10408000;
      21489: inst = 32'hc4049a5;
      21490: inst = 32'h8220000;
      21491: inst = 32'h10408000;
      21492: inst = 32'hc4049fa;
      21493: inst = 32'h8220000;
      21494: inst = 32'h10408000;
      21495: inst = 32'hc4049fb;
      21496: inst = 32'h8220000;
      21497: inst = 32'h10408000;
      21498: inst = 32'hc404a04;
      21499: inst = 32'h8220000;
      21500: inst = 32'h10408000;
      21501: inst = 32'hc404a05;
      21502: inst = 32'h8220000;
      21503: inst = 32'h10408000;
      21504: inst = 32'hc404a5a;
      21505: inst = 32'h8220000;
      21506: inst = 32'h10408000;
      21507: inst = 32'hc404a5b;
      21508: inst = 32'h8220000;
      21509: inst = 32'h10408000;
      21510: inst = 32'hc404a64;
      21511: inst = 32'h8220000;
      21512: inst = 32'h10408000;
      21513: inst = 32'hc404a65;
      21514: inst = 32'h8220000;
      21515: inst = 32'h10408000;
      21516: inst = 32'hc404aba;
      21517: inst = 32'h8220000;
      21518: inst = 32'h10408000;
      21519: inst = 32'hc404abb;
      21520: inst = 32'h8220000;
      21521: inst = 32'h10408000;
      21522: inst = 32'hc404ac4;
      21523: inst = 32'h8220000;
      21524: inst = 32'h10408000;
      21525: inst = 32'hc404ac5;
      21526: inst = 32'h8220000;
      21527: inst = 32'h10408000;
      21528: inst = 32'hc404b1a;
      21529: inst = 32'h8220000;
      21530: inst = 32'h10408000;
      21531: inst = 32'hc404b1b;
      21532: inst = 32'h8220000;
      21533: inst = 32'h10408000;
      21534: inst = 32'hc404b24;
      21535: inst = 32'h8220000;
      21536: inst = 32'h10408000;
      21537: inst = 32'hc404b25;
      21538: inst = 32'h8220000;
      21539: inst = 32'h10408000;
      21540: inst = 32'hc404b7a;
      21541: inst = 32'h8220000;
      21542: inst = 32'h10408000;
      21543: inst = 32'hc404b7b;
      21544: inst = 32'h8220000;
      21545: inst = 32'h10408000;
      21546: inst = 32'hc404b84;
      21547: inst = 32'h8220000;
      21548: inst = 32'h10408000;
      21549: inst = 32'hc404b85;
      21550: inst = 32'h8220000;
      21551: inst = 32'h10408000;
      21552: inst = 32'hc404bda;
      21553: inst = 32'h8220000;
      21554: inst = 32'h10408000;
      21555: inst = 32'hc404bdb;
      21556: inst = 32'h8220000;
      21557: inst = 32'h10408000;
      21558: inst = 32'hc404be4;
      21559: inst = 32'h8220000;
      21560: inst = 32'h10408000;
      21561: inst = 32'hc404be5;
      21562: inst = 32'h8220000;
      21563: inst = 32'h10408000;
      21564: inst = 32'hc404c3a;
      21565: inst = 32'h8220000;
      21566: inst = 32'h10408000;
      21567: inst = 32'hc404c3b;
      21568: inst = 32'h8220000;
      21569: inst = 32'h10408000;
      21570: inst = 32'hc404c44;
      21571: inst = 32'h8220000;
      21572: inst = 32'h10408000;
      21573: inst = 32'hc404c45;
      21574: inst = 32'h8220000;
      21575: inst = 32'h10408000;
      21576: inst = 32'hc404c9a;
      21577: inst = 32'h8220000;
      21578: inst = 32'h10408000;
      21579: inst = 32'hc404c9b;
      21580: inst = 32'h8220000;
      21581: inst = 32'h10408000;
      21582: inst = 32'hc404ca4;
      21583: inst = 32'h8220000;
      21584: inst = 32'h10408000;
      21585: inst = 32'hc404ca5;
      21586: inst = 32'h8220000;
      21587: inst = 32'h10408000;
      21588: inst = 32'hc404cfa;
      21589: inst = 32'h8220000;
      21590: inst = 32'h10408000;
      21591: inst = 32'hc404cfb;
      21592: inst = 32'h8220000;
      21593: inst = 32'h10408000;
      21594: inst = 32'hc404d04;
      21595: inst = 32'h8220000;
      21596: inst = 32'h10408000;
      21597: inst = 32'hc404d05;
      21598: inst = 32'h8220000;
      21599: inst = 32'h10408000;
      21600: inst = 32'hc404d5a;
      21601: inst = 32'h8220000;
      21602: inst = 32'h10408000;
      21603: inst = 32'hc404d5b;
      21604: inst = 32'h8220000;
      21605: inst = 32'h10408000;
      21606: inst = 32'hc404d64;
      21607: inst = 32'h8220000;
      21608: inst = 32'h10408000;
      21609: inst = 32'hc404d65;
      21610: inst = 32'h8220000;
      21611: inst = 32'h10408000;
      21612: inst = 32'hc404dba;
      21613: inst = 32'h8220000;
      21614: inst = 32'h10408000;
      21615: inst = 32'hc404dbb;
      21616: inst = 32'h8220000;
      21617: inst = 32'h10408000;
      21618: inst = 32'hc404dc4;
      21619: inst = 32'h8220000;
      21620: inst = 32'h10408000;
      21621: inst = 32'hc404dc5;
      21622: inst = 32'h8220000;
      21623: inst = 32'h10408000;
      21624: inst = 32'hc404e1a;
      21625: inst = 32'h8220000;
      21626: inst = 32'h10408000;
      21627: inst = 32'hc404e1b;
      21628: inst = 32'h8220000;
      21629: inst = 32'h10408000;
      21630: inst = 32'hc404e24;
      21631: inst = 32'h8220000;
      21632: inst = 32'h10408000;
      21633: inst = 32'hc404e25;
      21634: inst = 32'h8220000;
      21635: inst = 32'h10408000;
      21636: inst = 32'hc404e7a;
      21637: inst = 32'h8220000;
      21638: inst = 32'h10408000;
      21639: inst = 32'hc404e7b;
      21640: inst = 32'h8220000;
      21641: inst = 32'h10408000;
      21642: inst = 32'hc404e84;
      21643: inst = 32'h8220000;
      21644: inst = 32'h10408000;
      21645: inst = 32'hc404e85;
      21646: inst = 32'h8220000;
      21647: inst = 32'h10408000;
      21648: inst = 32'hc404eda;
      21649: inst = 32'h8220000;
      21650: inst = 32'h10408000;
      21651: inst = 32'hc404edb;
      21652: inst = 32'h8220000;
      21653: inst = 32'h10408000;
      21654: inst = 32'hc404ee4;
      21655: inst = 32'h8220000;
      21656: inst = 32'h10408000;
      21657: inst = 32'hc404ee5;
      21658: inst = 32'h8220000;
      21659: inst = 32'h10408000;
      21660: inst = 32'hc404f3a;
      21661: inst = 32'h8220000;
      21662: inst = 32'h10408000;
      21663: inst = 32'hc404f3b;
      21664: inst = 32'h8220000;
      21665: inst = 32'h10408000;
      21666: inst = 32'hc404f44;
      21667: inst = 32'h8220000;
      21668: inst = 32'h10408000;
      21669: inst = 32'hc404f45;
      21670: inst = 32'h8220000;
      21671: inst = 32'h10408000;
      21672: inst = 32'hc404f9a;
      21673: inst = 32'h8220000;
      21674: inst = 32'h10408000;
      21675: inst = 32'hc404f9b;
      21676: inst = 32'h8220000;
      21677: inst = 32'h10408000;
      21678: inst = 32'hc404fa4;
      21679: inst = 32'h8220000;
      21680: inst = 32'h10408000;
      21681: inst = 32'hc404fa5;
      21682: inst = 32'h8220000;
      21683: inst = 32'h10408000;
      21684: inst = 32'hc404ffa;
      21685: inst = 32'h8220000;
      21686: inst = 32'h10408000;
      21687: inst = 32'hc404ffb;
      21688: inst = 32'h8220000;
      21689: inst = 32'h10408000;
      21690: inst = 32'hc405004;
      21691: inst = 32'h8220000;
      21692: inst = 32'h10408000;
      21693: inst = 32'hc405005;
      21694: inst = 32'h8220000;
      21695: inst = 32'h10408000;
      21696: inst = 32'hc40505a;
      21697: inst = 32'h8220000;
      21698: inst = 32'h10408000;
      21699: inst = 32'hc40505b;
      21700: inst = 32'h8220000;
      21701: inst = 32'h10408000;
      21702: inst = 32'hc405064;
      21703: inst = 32'h8220000;
      21704: inst = 32'h10408000;
      21705: inst = 32'hc405065;
      21706: inst = 32'h8220000;
      21707: inst = 32'h10408000;
      21708: inst = 32'hc4050ba;
      21709: inst = 32'h8220000;
      21710: inst = 32'h10408000;
      21711: inst = 32'hc4050bb;
      21712: inst = 32'h8220000;
      21713: inst = 32'h10408000;
      21714: inst = 32'hc4050c4;
      21715: inst = 32'h8220000;
      21716: inst = 32'h10408000;
      21717: inst = 32'hc4050c5;
      21718: inst = 32'h8220000;
      21719: inst = 32'h10408000;
      21720: inst = 32'hc40511a;
      21721: inst = 32'h8220000;
      21722: inst = 32'h10408000;
      21723: inst = 32'hc40511b;
      21724: inst = 32'h8220000;
      21725: inst = 32'h10408000;
      21726: inst = 32'hc405124;
      21727: inst = 32'h8220000;
      21728: inst = 32'h10408000;
      21729: inst = 32'hc405125;
      21730: inst = 32'h8220000;
      21731: inst = 32'h10408000;
      21732: inst = 32'hc40517a;
      21733: inst = 32'h8220000;
      21734: inst = 32'h10408000;
      21735: inst = 32'hc40517b;
      21736: inst = 32'h8220000;
      21737: inst = 32'h10408000;
      21738: inst = 32'hc405184;
      21739: inst = 32'h8220000;
      21740: inst = 32'h10408000;
      21741: inst = 32'hc405185;
      21742: inst = 32'h8220000;
      21743: inst = 32'h10408000;
      21744: inst = 32'hc4051da;
      21745: inst = 32'h8220000;
      21746: inst = 32'h10408000;
      21747: inst = 32'hc4051db;
      21748: inst = 32'h8220000;
      21749: inst = 32'h10408000;
      21750: inst = 32'hc4051e4;
      21751: inst = 32'h8220000;
      21752: inst = 32'h10408000;
      21753: inst = 32'hc4051e5;
      21754: inst = 32'h8220000;
      21755: inst = 32'h10408000;
      21756: inst = 32'hc40523a;
      21757: inst = 32'h8220000;
      21758: inst = 32'h10408000;
      21759: inst = 32'hc40523b;
      21760: inst = 32'h8220000;
      21761: inst = 32'h10408000;
      21762: inst = 32'hc405244;
      21763: inst = 32'h8220000;
      21764: inst = 32'h10408000;
      21765: inst = 32'hc405245;
      21766: inst = 32'h8220000;
      21767: inst = 32'h10408000;
      21768: inst = 32'hc40529a;
      21769: inst = 32'h8220000;
      21770: inst = 32'h10408000;
      21771: inst = 32'hc40529b;
      21772: inst = 32'h8220000;
      21773: inst = 32'h10408000;
      21774: inst = 32'hc4052a4;
      21775: inst = 32'h8220000;
      21776: inst = 32'h10408000;
      21777: inst = 32'hc4052a5;
      21778: inst = 32'h8220000;
      21779: inst = 32'h10408000;
      21780: inst = 32'hc4052fa;
      21781: inst = 32'h8220000;
      21782: inst = 32'h10408000;
      21783: inst = 32'hc4052fb;
      21784: inst = 32'h8220000;
      21785: inst = 32'h10408000;
      21786: inst = 32'hc405304;
      21787: inst = 32'h8220000;
      21788: inst = 32'h10408000;
      21789: inst = 32'hc405305;
      21790: inst = 32'h8220000;
      21791: inst = 32'h10408000;
      21792: inst = 32'hc40535a;
      21793: inst = 32'h8220000;
      21794: inst = 32'h10408000;
      21795: inst = 32'hc40535b;
      21796: inst = 32'h8220000;
      21797: inst = 32'h10408000;
      21798: inst = 32'hc405364;
      21799: inst = 32'h8220000;
      21800: inst = 32'h10408000;
      21801: inst = 32'hc405365;
      21802: inst = 32'h8220000;
      21803: inst = 32'h10408000;
      21804: inst = 32'hc4053ba;
      21805: inst = 32'h8220000;
      21806: inst = 32'h10408000;
      21807: inst = 32'hc4053bb;
      21808: inst = 32'h8220000;
      21809: inst = 32'h10408000;
      21810: inst = 32'hc4053c4;
      21811: inst = 32'h8220000;
      21812: inst = 32'h10408000;
      21813: inst = 32'hc4053c5;
      21814: inst = 32'h8220000;
      21815: inst = 32'h10408000;
      21816: inst = 32'hc40541a;
      21817: inst = 32'h8220000;
      21818: inst = 32'h10408000;
      21819: inst = 32'hc40541b;
      21820: inst = 32'h8220000;
      21821: inst = 32'h10408000;
      21822: inst = 32'hc405424;
      21823: inst = 32'h8220000;
      21824: inst = 32'h10408000;
      21825: inst = 32'hc405425;
      21826: inst = 32'h8220000;
      21827: inst = 32'h10408000;
      21828: inst = 32'hc405426;
      21829: inst = 32'h8220000;
      21830: inst = 32'h10408000;
      21831: inst = 32'hc405479;
      21832: inst = 32'h8220000;
      21833: inst = 32'h10408000;
      21834: inst = 32'hc40547a;
      21835: inst = 32'h8220000;
      21836: inst = 32'h10408000;
      21837: inst = 32'hc40547b;
      21838: inst = 32'h8220000;
      21839: inst = 32'h10408000;
      21840: inst = 32'hc405484;
      21841: inst = 32'h8220000;
      21842: inst = 32'h10408000;
      21843: inst = 32'hc405485;
      21844: inst = 32'h8220000;
      21845: inst = 32'h10408000;
      21846: inst = 32'hc405486;
      21847: inst = 32'h8220000;
      21848: inst = 32'h10408000;
      21849: inst = 32'hc405487;
      21850: inst = 32'h8220000;
      21851: inst = 32'h10408000;
      21852: inst = 32'hc405488;
      21853: inst = 32'h8220000;
      21854: inst = 32'h10408000;
      21855: inst = 32'hc405489;
      21856: inst = 32'h8220000;
      21857: inst = 32'h10408000;
      21858: inst = 32'hc40548a;
      21859: inst = 32'h8220000;
      21860: inst = 32'h10408000;
      21861: inst = 32'hc40548b;
      21862: inst = 32'h8220000;
      21863: inst = 32'h10408000;
      21864: inst = 32'hc40548c;
      21865: inst = 32'h8220000;
      21866: inst = 32'h10408000;
      21867: inst = 32'hc40548d;
      21868: inst = 32'h8220000;
      21869: inst = 32'h10408000;
      21870: inst = 32'hc40548e;
      21871: inst = 32'h8220000;
      21872: inst = 32'h10408000;
      21873: inst = 32'hc40548f;
      21874: inst = 32'h8220000;
      21875: inst = 32'h10408000;
      21876: inst = 32'hc405490;
      21877: inst = 32'h8220000;
      21878: inst = 32'h10408000;
      21879: inst = 32'hc405491;
      21880: inst = 32'h8220000;
      21881: inst = 32'h10408000;
      21882: inst = 32'hc405492;
      21883: inst = 32'h8220000;
      21884: inst = 32'h10408000;
      21885: inst = 32'hc405493;
      21886: inst = 32'h8220000;
      21887: inst = 32'h10408000;
      21888: inst = 32'hc405494;
      21889: inst = 32'h8220000;
      21890: inst = 32'h10408000;
      21891: inst = 32'hc405495;
      21892: inst = 32'h8220000;
      21893: inst = 32'h10408000;
      21894: inst = 32'hc405496;
      21895: inst = 32'h8220000;
      21896: inst = 32'h10408000;
      21897: inst = 32'hc405497;
      21898: inst = 32'h8220000;
      21899: inst = 32'h10408000;
      21900: inst = 32'hc405498;
      21901: inst = 32'h8220000;
      21902: inst = 32'h10408000;
      21903: inst = 32'hc405499;
      21904: inst = 32'h8220000;
      21905: inst = 32'h10408000;
      21906: inst = 32'hc40549a;
      21907: inst = 32'h8220000;
      21908: inst = 32'h10408000;
      21909: inst = 32'hc40549b;
      21910: inst = 32'h8220000;
      21911: inst = 32'h10408000;
      21912: inst = 32'hc40549c;
      21913: inst = 32'h8220000;
      21914: inst = 32'h10408000;
      21915: inst = 32'hc40549d;
      21916: inst = 32'h8220000;
      21917: inst = 32'h10408000;
      21918: inst = 32'hc40549e;
      21919: inst = 32'h8220000;
      21920: inst = 32'h10408000;
      21921: inst = 32'hc40549f;
      21922: inst = 32'h8220000;
      21923: inst = 32'h10408000;
      21924: inst = 32'hc4054a0;
      21925: inst = 32'h8220000;
      21926: inst = 32'h10408000;
      21927: inst = 32'hc4054a1;
      21928: inst = 32'h8220000;
      21929: inst = 32'h10408000;
      21930: inst = 32'hc4054a2;
      21931: inst = 32'h8220000;
      21932: inst = 32'h10408000;
      21933: inst = 32'hc4054a3;
      21934: inst = 32'h8220000;
      21935: inst = 32'h10408000;
      21936: inst = 32'hc4054a4;
      21937: inst = 32'h8220000;
      21938: inst = 32'h10408000;
      21939: inst = 32'hc4054a5;
      21940: inst = 32'h8220000;
      21941: inst = 32'h10408000;
      21942: inst = 32'hc4054a6;
      21943: inst = 32'h8220000;
      21944: inst = 32'h10408000;
      21945: inst = 32'hc4054a7;
      21946: inst = 32'h8220000;
      21947: inst = 32'h10408000;
      21948: inst = 32'hc4054a8;
      21949: inst = 32'h8220000;
      21950: inst = 32'h10408000;
      21951: inst = 32'hc4054a9;
      21952: inst = 32'h8220000;
      21953: inst = 32'h10408000;
      21954: inst = 32'hc4054aa;
      21955: inst = 32'h8220000;
      21956: inst = 32'h10408000;
      21957: inst = 32'hc4054ab;
      21958: inst = 32'h8220000;
      21959: inst = 32'h10408000;
      21960: inst = 32'hc4054ac;
      21961: inst = 32'h8220000;
      21962: inst = 32'h10408000;
      21963: inst = 32'hc4054ad;
      21964: inst = 32'h8220000;
      21965: inst = 32'h10408000;
      21966: inst = 32'hc4054ae;
      21967: inst = 32'h8220000;
      21968: inst = 32'h10408000;
      21969: inst = 32'hc4054af;
      21970: inst = 32'h8220000;
      21971: inst = 32'h10408000;
      21972: inst = 32'hc4054b0;
      21973: inst = 32'h8220000;
      21974: inst = 32'h10408000;
      21975: inst = 32'hc4054b1;
      21976: inst = 32'h8220000;
      21977: inst = 32'h10408000;
      21978: inst = 32'hc4054b2;
      21979: inst = 32'h8220000;
      21980: inst = 32'h10408000;
      21981: inst = 32'hc4054b3;
      21982: inst = 32'h8220000;
      21983: inst = 32'h10408000;
      21984: inst = 32'hc4054b4;
      21985: inst = 32'h8220000;
      21986: inst = 32'h10408000;
      21987: inst = 32'hc4054b5;
      21988: inst = 32'h8220000;
      21989: inst = 32'h10408000;
      21990: inst = 32'hc4054b6;
      21991: inst = 32'h8220000;
      21992: inst = 32'h10408000;
      21993: inst = 32'hc4054b7;
      21994: inst = 32'h8220000;
      21995: inst = 32'h10408000;
      21996: inst = 32'hc4054b8;
      21997: inst = 32'h8220000;
      21998: inst = 32'h10408000;
      21999: inst = 32'hc4054b9;
      22000: inst = 32'h8220000;
      22001: inst = 32'h10408000;
      22002: inst = 32'hc4054ba;
      22003: inst = 32'h8220000;
      22004: inst = 32'h10408000;
      22005: inst = 32'hc4054bb;
      22006: inst = 32'h8220000;
      22007: inst = 32'h10408000;
      22008: inst = 32'hc4054bc;
      22009: inst = 32'h8220000;
      22010: inst = 32'h10408000;
      22011: inst = 32'hc4054bd;
      22012: inst = 32'h8220000;
      22013: inst = 32'h10408000;
      22014: inst = 32'hc4054be;
      22015: inst = 32'h8220000;
      22016: inst = 32'h10408000;
      22017: inst = 32'hc4054bf;
      22018: inst = 32'h8220000;
      22019: inst = 32'h10408000;
      22020: inst = 32'hc4054c0;
      22021: inst = 32'h8220000;
      22022: inst = 32'h10408000;
      22023: inst = 32'hc4054c1;
      22024: inst = 32'h8220000;
      22025: inst = 32'h10408000;
      22026: inst = 32'hc4054c2;
      22027: inst = 32'h8220000;
      22028: inst = 32'h10408000;
      22029: inst = 32'hc4054c3;
      22030: inst = 32'h8220000;
      22031: inst = 32'h10408000;
      22032: inst = 32'hc4054c4;
      22033: inst = 32'h8220000;
      22034: inst = 32'h10408000;
      22035: inst = 32'hc4054c5;
      22036: inst = 32'h8220000;
      22037: inst = 32'h10408000;
      22038: inst = 32'hc4054c6;
      22039: inst = 32'h8220000;
      22040: inst = 32'h10408000;
      22041: inst = 32'hc4054c7;
      22042: inst = 32'h8220000;
      22043: inst = 32'h10408000;
      22044: inst = 32'hc4054c8;
      22045: inst = 32'h8220000;
      22046: inst = 32'h10408000;
      22047: inst = 32'hc4054c9;
      22048: inst = 32'h8220000;
      22049: inst = 32'h10408000;
      22050: inst = 32'hc4054ca;
      22051: inst = 32'h8220000;
      22052: inst = 32'h10408000;
      22053: inst = 32'hc4054cb;
      22054: inst = 32'h8220000;
      22055: inst = 32'h10408000;
      22056: inst = 32'hc4054cc;
      22057: inst = 32'h8220000;
      22058: inst = 32'h10408000;
      22059: inst = 32'hc4054cd;
      22060: inst = 32'h8220000;
      22061: inst = 32'h10408000;
      22062: inst = 32'hc4054ce;
      22063: inst = 32'h8220000;
      22064: inst = 32'h10408000;
      22065: inst = 32'hc4054cf;
      22066: inst = 32'h8220000;
      22067: inst = 32'h10408000;
      22068: inst = 32'hc4054d0;
      22069: inst = 32'h8220000;
      22070: inst = 32'h10408000;
      22071: inst = 32'hc4054d1;
      22072: inst = 32'h8220000;
      22073: inst = 32'h10408000;
      22074: inst = 32'hc4054d2;
      22075: inst = 32'h8220000;
      22076: inst = 32'h10408000;
      22077: inst = 32'hc4054d3;
      22078: inst = 32'h8220000;
      22079: inst = 32'h10408000;
      22080: inst = 32'hc4054d4;
      22081: inst = 32'h8220000;
      22082: inst = 32'h10408000;
      22083: inst = 32'hc4054d5;
      22084: inst = 32'h8220000;
      22085: inst = 32'h10408000;
      22086: inst = 32'hc4054d6;
      22087: inst = 32'h8220000;
      22088: inst = 32'h10408000;
      22089: inst = 32'hc4054d7;
      22090: inst = 32'h8220000;
      22091: inst = 32'h10408000;
      22092: inst = 32'hc4054d8;
      22093: inst = 32'h8220000;
      22094: inst = 32'h10408000;
      22095: inst = 32'hc4054d9;
      22096: inst = 32'h8220000;
      22097: inst = 32'h10408000;
      22098: inst = 32'hc4054da;
      22099: inst = 32'h8220000;
      22100: inst = 32'h10408000;
      22101: inst = 32'hc4054db;
      22102: inst = 32'h8220000;
      22103: inst = 32'h10408000;
      22104: inst = 32'hc4054e4;
      22105: inst = 32'h8220000;
      22106: inst = 32'h10408000;
      22107: inst = 32'hc4054e5;
      22108: inst = 32'h8220000;
      22109: inst = 32'h10408000;
      22110: inst = 32'hc4054e6;
      22111: inst = 32'h8220000;
      22112: inst = 32'h10408000;
      22113: inst = 32'hc4054e7;
      22114: inst = 32'h8220000;
      22115: inst = 32'h10408000;
      22116: inst = 32'hc4054e8;
      22117: inst = 32'h8220000;
      22118: inst = 32'h10408000;
      22119: inst = 32'hc4054e9;
      22120: inst = 32'h8220000;
      22121: inst = 32'h10408000;
      22122: inst = 32'hc4054ea;
      22123: inst = 32'h8220000;
      22124: inst = 32'h10408000;
      22125: inst = 32'hc4054eb;
      22126: inst = 32'h8220000;
      22127: inst = 32'h10408000;
      22128: inst = 32'hc4054ec;
      22129: inst = 32'h8220000;
      22130: inst = 32'h10408000;
      22131: inst = 32'hc4054ed;
      22132: inst = 32'h8220000;
      22133: inst = 32'h10408000;
      22134: inst = 32'hc4054ee;
      22135: inst = 32'h8220000;
      22136: inst = 32'h10408000;
      22137: inst = 32'hc4054ef;
      22138: inst = 32'h8220000;
      22139: inst = 32'h10408000;
      22140: inst = 32'hc4054f0;
      22141: inst = 32'h8220000;
      22142: inst = 32'h10408000;
      22143: inst = 32'hc4054f1;
      22144: inst = 32'h8220000;
      22145: inst = 32'h10408000;
      22146: inst = 32'hc4054f2;
      22147: inst = 32'h8220000;
      22148: inst = 32'h10408000;
      22149: inst = 32'hc4054f3;
      22150: inst = 32'h8220000;
      22151: inst = 32'h10408000;
      22152: inst = 32'hc4054f4;
      22153: inst = 32'h8220000;
      22154: inst = 32'h10408000;
      22155: inst = 32'hc4054f5;
      22156: inst = 32'h8220000;
      22157: inst = 32'h10408000;
      22158: inst = 32'hc4054f6;
      22159: inst = 32'h8220000;
      22160: inst = 32'h10408000;
      22161: inst = 32'hc4054f7;
      22162: inst = 32'h8220000;
      22163: inst = 32'h10408000;
      22164: inst = 32'hc4054f8;
      22165: inst = 32'h8220000;
      22166: inst = 32'h10408000;
      22167: inst = 32'hc4054f9;
      22168: inst = 32'h8220000;
      22169: inst = 32'h10408000;
      22170: inst = 32'hc4054fa;
      22171: inst = 32'h8220000;
      22172: inst = 32'h10408000;
      22173: inst = 32'hc4054fb;
      22174: inst = 32'h8220000;
      22175: inst = 32'h10408000;
      22176: inst = 32'hc4054fc;
      22177: inst = 32'h8220000;
      22178: inst = 32'h10408000;
      22179: inst = 32'hc4054fd;
      22180: inst = 32'h8220000;
      22181: inst = 32'h10408000;
      22182: inst = 32'hc4054fe;
      22183: inst = 32'h8220000;
      22184: inst = 32'h10408000;
      22185: inst = 32'hc4054ff;
      22186: inst = 32'h8220000;
      22187: inst = 32'h10408000;
      22188: inst = 32'hc405500;
      22189: inst = 32'h8220000;
      22190: inst = 32'h10408000;
      22191: inst = 32'hc405501;
      22192: inst = 32'h8220000;
      22193: inst = 32'h10408000;
      22194: inst = 32'hc405502;
      22195: inst = 32'h8220000;
      22196: inst = 32'h10408000;
      22197: inst = 32'hc405503;
      22198: inst = 32'h8220000;
      22199: inst = 32'h10408000;
      22200: inst = 32'hc405504;
      22201: inst = 32'h8220000;
      22202: inst = 32'h10408000;
      22203: inst = 32'hc405505;
      22204: inst = 32'h8220000;
      22205: inst = 32'h10408000;
      22206: inst = 32'hc405506;
      22207: inst = 32'h8220000;
      22208: inst = 32'h10408000;
      22209: inst = 32'hc405507;
      22210: inst = 32'h8220000;
      22211: inst = 32'h10408000;
      22212: inst = 32'hc405508;
      22213: inst = 32'h8220000;
      22214: inst = 32'h10408000;
      22215: inst = 32'hc405509;
      22216: inst = 32'h8220000;
      22217: inst = 32'h10408000;
      22218: inst = 32'hc40550a;
      22219: inst = 32'h8220000;
      22220: inst = 32'h10408000;
      22221: inst = 32'hc40550b;
      22222: inst = 32'h8220000;
      22223: inst = 32'h10408000;
      22224: inst = 32'hc40550c;
      22225: inst = 32'h8220000;
      22226: inst = 32'h10408000;
      22227: inst = 32'hc40550d;
      22228: inst = 32'h8220000;
      22229: inst = 32'h10408000;
      22230: inst = 32'hc40550e;
      22231: inst = 32'h8220000;
      22232: inst = 32'h10408000;
      22233: inst = 32'hc40550f;
      22234: inst = 32'h8220000;
      22235: inst = 32'h10408000;
      22236: inst = 32'hc405510;
      22237: inst = 32'h8220000;
      22238: inst = 32'h10408000;
      22239: inst = 32'hc405511;
      22240: inst = 32'h8220000;
      22241: inst = 32'h10408000;
      22242: inst = 32'hc405512;
      22243: inst = 32'h8220000;
      22244: inst = 32'h10408000;
      22245: inst = 32'hc405513;
      22246: inst = 32'h8220000;
      22247: inst = 32'h10408000;
      22248: inst = 32'hc405514;
      22249: inst = 32'h8220000;
      22250: inst = 32'h10408000;
      22251: inst = 32'hc405515;
      22252: inst = 32'h8220000;
      22253: inst = 32'h10408000;
      22254: inst = 32'hc405516;
      22255: inst = 32'h8220000;
      22256: inst = 32'h10408000;
      22257: inst = 32'hc405517;
      22258: inst = 32'h8220000;
      22259: inst = 32'h10408000;
      22260: inst = 32'hc405518;
      22261: inst = 32'h8220000;
      22262: inst = 32'h10408000;
      22263: inst = 32'hc405519;
      22264: inst = 32'h8220000;
      22265: inst = 32'h10408000;
      22266: inst = 32'hc40551a;
      22267: inst = 32'h8220000;
      22268: inst = 32'h10408000;
      22269: inst = 32'hc40551b;
      22270: inst = 32'h8220000;
      22271: inst = 32'h10408000;
      22272: inst = 32'hc40551c;
      22273: inst = 32'h8220000;
      22274: inst = 32'h10408000;
      22275: inst = 32'hc40551d;
      22276: inst = 32'h8220000;
      22277: inst = 32'h10408000;
      22278: inst = 32'hc40551e;
      22279: inst = 32'h8220000;
      22280: inst = 32'h10408000;
      22281: inst = 32'hc40551f;
      22282: inst = 32'h8220000;
      22283: inst = 32'h10408000;
      22284: inst = 32'hc405520;
      22285: inst = 32'h8220000;
      22286: inst = 32'h10408000;
      22287: inst = 32'hc405521;
      22288: inst = 32'h8220000;
      22289: inst = 32'h10408000;
      22290: inst = 32'hc405522;
      22291: inst = 32'h8220000;
      22292: inst = 32'h10408000;
      22293: inst = 32'hc405523;
      22294: inst = 32'h8220000;
      22295: inst = 32'h10408000;
      22296: inst = 32'hc405524;
      22297: inst = 32'h8220000;
      22298: inst = 32'h10408000;
      22299: inst = 32'hc405525;
      22300: inst = 32'h8220000;
      22301: inst = 32'h10408000;
      22302: inst = 32'hc405526;
      22303: inst = 32'h8220000;
      22304: inst = 32'h10408000;
      22305: inst = 32'hc405527;
      22306: inst = 32'h8220000;
      22307: inst = 32'h10408000;
      22308: inst = 32'hc405528;
      22309: inst = 32'h8220000;
      22310: inst = 32'h10408000;
      22311: inst = 32'hc405529;
      22312: inst = 32'h8220000;
      22313: inst = 32'h10408000;
      22314: inst = 32'hc40552a;
      22315: inst = 32'h8220000;
      22316: inst = 32'h10408000;
      22317: inst = 32'hc40552b;
      22318: inst = 32'h8220000;
      22319: inst = 32'h10408000;
      22320: inst = 32'hc40552c;
      22321: inst = 32'h8220000;
      22322: inst = 32'h10408000;
      22323: inst = 32'hc40552d;
      22324: inst = 32'h8220000;
      22325: inst = 32'h10408000;
      22326: inst = 32'hc40552e;
      22327: inst = 32'h8220000;
      22328: inst = 32'h10408000;
      22329: inst = 32'hc40552f;
      22330: inst = 32'h8220000;
      22331: inst = 32'h10408000;
      22332: inst = 32'hc405530;
      22333: inst = 32'h8220000;
      22334: inst = 32'h10408000;
      22335: inst = 32'hc405531;
      22336: inst = 32'h8220000;
      22337: inst = 32'h10408000;
      22338: inst = 32'hc405532;
      22339: inst = 32'h8220000;
      22340: inst = 32'h10408000;
      22341: inst = 32'hc405533;
      22342: inst = 32'h8220000;
      22343: inst = 32'h10408000;
      22344: inst = 32'hc405534;
      22345: inst = 32'h8220000;
      22346: inst = 32'h10408000;
      22347: inst = 32'hc405535;
      22348: inst = 32'h8220000;
      22349: inst = 32'h10408000;
      22350: inst = 32'hc405536;
      22351: inst = 32'h8220000;
      22352: inst = 32'h10408000;
      22353: inst = 32'hc405537;
      22354: inst = 32'h8220000;
      22355: inst = 32'h10408000;
      22356: inst = 32'hc405538;
      22357: inst = 32'h8220000;
      22358: inst = 32'h10408000;
      22359: inst = 32'hc405539;
      22360: inst = 32'h8220000;
      22361: inst = 32'h10408000;
      22362: inst = 32'hc40553a;
      22363: inst = 32'h8220000;
      22364: inst = 32'h10408000;
      22365: inst = 32'hc40553b;
      22366: inst = 32'h8220000;
      22367: inst = 32'hc204a7a;
      22368: inst = 32'h10408000;
      22369: inst = 32'hc4042e7;
      22370: inst = 32'h8220000;
      22371: inst = 32'h10408000;
      22372: inst = 32'hc404338;
      22373: inst = 32'h8220000;
      22374: inst = 32'h10408000;
      22375: inst = 32'hc404346;
      22376: inst = 32'h8220000;
      22377: inst = 32'h10408000;
      22378: inst = 32'hc404399;
      22379: inst = 32'h8220000;
      22380: inst = 32'h10408000;
      22381: inst = 32'hc4053c6;
      22382: inst = 32'h8220000;
      22383: inst = 32'h10408000;
      22384: inst = 32'hc405419;
      22385: inst = 32'h8220000;
      22386: inst = 32'h10408000;
      22387: inst = 32'hc405427;
      22388: inst = 32'h8220000;
      22389: inst = 32'h10408000;
      22390: inst = 32'hc405478;
      22391: inst = 32'h8220000;
      22392: inst = 32'hc2031b0;
      22393: inst = 32'h10408000;
      22394: inst = 32'hc4042e8;
      22395: inst = 32'h8220000;
      22396: inst = 32'h10408000;
      22397: inst = 32'hc404337;
      22398: inst = 32'h8220000;
      22399: inst = 32'h10408000;
      22400: inst = 32'hc4043a6;
      22401: inst = 32'h8220000;
      22402: inst = 32'h10408000;
      22403: inst = 32'hc4043f9;
      22404: inst = 32'h8220000;
      22405: inst = 32'h10408000;
      22406: inst = 32'hc405366;
      22407: inst = 32'h8220000;
      22408: inst = 32'h10408000;
      22409: inst = 32'hc4053b9;
      22410: inst = 32'h8220000;
      22411: inst = 32'h10408000;
      22412: inst = 32'hc405428;
      22413: inst = 32'h8220000;
      22414: inst = 32'h10408000;
      22415: inst = 32'hc405477;
      22416: inst = 32'h8220000;
      22417: inst = 32'hc20296d;
      22418: inst = 32'h10408000;
      22419: inst = 32'hc4042e9;
      22420: inst = 32'h8220000;
      22421: inst = 32'h10408000;
      22422: inst = 32'hc4042ea;
      22423: inst = 32'h8220000;
      22424: inst = 32'h10408000;
      22425: inst = 32'hc4042eb;
      22426: inst = 32'h8220000;
      22427: inst = 32'h10408000;
      22428: inst = 32'hc4042ec;
      22429: inst = 32'h8220000;
      22430: inst = 32'h10408000;
      22431: inst = 32'hc4042ed;
      22432: inst = 32'h8220000;
      22433: inst = 32'h10408000;
      22434: inst = 32'hc4042ee;
      22435: inst = 32'h8220000;
      22436: inst = 32'h10408000;
      22437: inst = 32'hc4042ef;
      22438: inst = 32'h8220000;
      22439: inst = 32'h10408000;
      22440: inst = 32'hc4042f0;
      22441: inst = 32'h8220000;
      22442: inst = 32'h10408000;
      22443: inst = 32'hc4042f1;
      22444: inst = 32'h8220000;
      22445: inst = 32'h10408000;
      22446: inst = 32'hc4042f2;
      22447: inst = 32'h8220000;
      22448: inst = 32'h10408000;
      22449: inst = 32'hc4042f3;
      22450: inst = 32'h8220000;
      22451: inst = 32'h10408000;
      22452: inst = 32'hc4042f4;
      22453: inst = 32'h8220000;
      22454: inst = 32'h10408000;
      22455: inst = 32'hc4042f5;
      22456: inst = 32'h8220000;
      22457: inst = 32'h10408000;
      22458: inst = 32'hc4042f6;
      22459: inst = 32'h8220000;
      22460: inst = 32'h10408000;
      22461: inst = 32'hc4042f7;
      22462: inst = 32'h8220000;
      22463: inst = 32'h10408000;
      22464: inst = 32'hc4042f8;
      22465: inst = 32'h8220000;
      22466: inst = 32'h10408000;
      22467: inst = 32'hc4042f9;
      22468: inst = 32'h8220000;
      22469: inst = 32'h10408000;
      22470: inst = 32'hc4042fa;
      22471: inst = 32'h8220000;
      22472: inst = 32'h10408000;
      22473: inst = 32'hc4042fb;
      22474: inst = 32'h8220000;
      22475: inst = 32'h10408000;
      22476: inst = 32'hc4042fc;
      22477: inst = 32'h8220000;
      22478: inst = 32'h10408000;
      22479: inst = 32'hc4042fd;
      22480: inst = 32'h8220000;
      22481: inst = 32'h10408000;
      22482: inst = 32'hc4042fe;
      22483: inst = 32'h8220000;
      22484: inst = 32'h10408000;
      22485: inst = 32'hc4042ff;
      22486: inst = 32'h8220000;
      22487: inst = 32'h10408000;
      22488: inst = 32'hc404300;
      22489: inst = 32'h8220000;
      22490: inst = 32'h10408000;
      22491: inst = 32'hc404301;
      22492: inst = 32'h8220000;
      22493: inst = 32'h10408000;
      22494: inst = 32'hc404302;
      22495: inst = 32'h8220000;
      22496: inst = 32'h10408000;
      22497: inst = 32'hc404303;
      22498: inst = 32'h8220000;
      22499: inst = 32'h10408000;
      22500: inst = 32'hc404304;
      22501: inst = 32'h8220000;
      22502: inst = 32'h10408000;
      22503: inst = 32'hc404305;
      22504: inst = 32'h8220000;
      22505: inst = 32'h10408000;
      22506: inst = 32'hc404306;
      22507: inst = 32'h8220000;
      22508: inst = 32'h10408000;
      22509: inst = 32'hc404307;
      22510: inst = 32'h8220000;
      22511: inst = 32'h10408000;
      22512: inst = 32'hc404308;
      22513: inst = 32'h8220000;
      22514: inst = 32'h10408000;
      22515: inst = 32'hc404309;
      22516: inst = 32'h8220000;
      22517: inst = 32'h10408000;
      22518: inst = 32'hc40430a;
      22519: inst = 32'h8220000;
      22520: inst = 32'h10408000;
      22521: inst = 32'hc40430b;
      22522: inst = 32'h8220000;
      22523: inst = 32'h10408000;
      22524: inst = 32'hc40430c;
      22525: inst = 32'h8220000;
      22526: inst = 32'h10408000;
      22527: inst = 32'hc40430d;
      22528: inst = 32'h8220000;
      22529: inst = 32'h10408000;
      22530: inst = 32'hc40430e;
      22531: inst = 32'h8220000;
      22532: inst = 32'h10408000;
      22533: inst = 32'hc40430f;
      22534: inst = 32'h8220000;
      22535: inst = 32'h10408000;
      22536: inst = 32'hc404310;
      22537: inst = 32'h8220000;
      22538: inst = 32'h10408000;
      22539: inst = 32'hc404311;
      22540: inst = 32'h8220000;
      22541: inst = 32'h10408000;
      22542: inst = 32'hc404312;
      22543: inst = 32'h8220000;
      22544: inst = 32'h10408000;
      22545: inst = 32'hc404313;
      22546: inst = 32'h8220000;
      22547: inst = 32'h10408000;
      22548: inst = 32'hc404314;
      22549: inst = 32'h8220000;
      22550: inst = 32'h10408000;
      22551: inst = 32'hc404315;
      22552: inst = 32'h8220000;
      22553: inst = 32'h10408000;
      22554: inst = 32'hc404316;
      22555: inst = 32'h8220000;
      22556: inst = 32'h10408000;
      22557: inst = 32'hc404317;
      22558: inst = 32'h8220000;
      22559: inst = 32'h10408000;
      22560: inst = 32'hc404318;
      22561: inst = 32'h8220000;
      22562: inst = 32'h10408000;
      22563: inst = 32'hc404319;
      22564: inst = 32'h8220000;
      22565: inst = 32'h10408000;
      22566: inst = 32'hc40431a;
      22567: inst = 32'h8220000;
      22568: inst = 32'h10408000;
      22569: inst = 32'hc40431b;
      22570: inst = 32'h8220000;
      22571: inst = 32'h10408000;
      22572: inst = 32'hc40431c;
      22573: inst = 32'h8220000;
      22574: inst = 32'h10408000;
      22575: inst = 32'hc40431d;
      22576: inst = 32'h8220000;
      22577: inst = 32'h10408000;
      22578: inst = 32'hc40431e;
      22579: inst = 32'h8220000;
      22580: inst = 32'h10408000;
      22581: inst = 32'hc40431f;
      22582: inst = 32'h8220000;
      22583: inst = 32'h10408000;
      22584: inst = 32'hc404320;
      22585: inst = 32'h8220000;
      22586: inst = 32'h10408000;
      22587: inst = 32'hc404321;
      22588: inst = 32'h8220000;
      22589: inst = 32'h10408000;
      22590: inst = 32'hc404322;
      22591: inst = 32'h8220000;
      22592: inst = 32'h10408000;
      22593: inst = 32'hc404323;
      22594: inst = 32'h8220000;
      22595: inst = 32'h10408000;
      22596: inst = 32'hc404324;
      22597: inst = 32'h8220000;
      22598: inst = 32'h10408000;
      22599: inst = 32'hc404325;
      22600: inst = 32'h8220000;
      22601: inst = 32'h10408000;
      22602: inst = 32'hc404326;
      22603: inst = 32'h8220000;
      22604: inst = 32'h10408000;
      22605: inst = 32'hc404327;
      22606: inst = 32'h8220000;
      22607: inst = 32'h10408000;
      22608: inst = 32'hc404328;
      22609: inst = 32'h8220000;
      22610: inst = 32'h10408000;
      22611: inst = 32'hc404329;
      22612: inst = 32'h8220000;
      22613: inst = 32'h10408000;
      22614: inst = 32'hc40432a;
      22615: inst = 32'h8220000;
      22616: inst = 32'h10408000;
      22617: inst = 32'hc40432b;
      22618: inst = 32'h8220000;
      22619: inst = 32'h10408000;
      22620: inst = 32'hc40432c;
      22621: inst = 32'h8220000;
      22622: inst = 32'h10408000;
      22623: inst = 32'hc40432d;
      22624: inst = 32'h8220000;
      22625: inst = 32'h10408000;
      22626: inst = 32'hc40432e;
      22627: inst = 32'h8220000;
      22628: inst = 32'h10408000;
      22629: inst = 32'hc40432f;
      22630: inst = 32'h8220000;
      22631: inst = 32'h10408000;
      22632: inst = 32'hc404330;
      22633: inst = 32'h8220000;
      22634: inst = 32'h10408000;
      22635: inst = 32'hc404331;
      22636: inst = 32'h8220000;
      22637: inst = 32'h10408000;
      22638: inst = 32'hc404332;
      22639: inst = 32'h8220000;
      22640: inst = 32'h10408000;
      22641: inst = 32'hc404333;
      22642: inst = 32'h8220000;
      22643: inst = 32'h10408000;
      22644: inst = 32'hc404334;
      22645: inst = 32'h8220000;
      22646: inst = 32'h10408000;
      22647: inst = 32'hc404335;
      22648: inst = 32'h8220000;
      22649: inst = 32'h10408000;
      22650: inst = 32'hc404336;
      22651: inst = 32'h8220000;
      22652: inst = 32'h10408000;
      22653: inst = 32'hc405429;
      22654: inst = 32'h8220000;
      22655: inst = 32'h10408000;
      22656: inst = 32'hc40542a;
      22657: inst = 32'h8220000;
      22658: inst = 32'h10408000;
      22659: inst = 32'hc40542b;
      22660: inst = 32'h8220000;
      22661: inst = 32'h10408000;
      22662: inst = 32'hc40542c;
      22663: inst = 32'h8220000;
      22664: inst = 32'h10408000;
      22665: inst = 32'hc40542d;
      22666: inst = 32'h8220000;
      22667: inst = 32'h10408000;
      22668: inst = 32'hc40542e;
      22669: inst = 32'h8220000;
      22670: inst = 32'h10408000;
      22671: inst = 32'hc40542f;
      22672: inst = 32'h8220000;
      22673: inst = 32'h10408000;
      22674: inst = 32'hc405430;
      22675: inst = 32'h8220000;
      22676: inst = 32'h10408000;
      22677: inst = 32'hc405431;
      22678: inst = 32'h8220000;
      22679: inst = 32'h10408000;
      22680: inst = 32'hc405432;
      22681: inst = 32'h8220000;
      22682: inst = 32'h10408000;
      22683: inst = 32'hc405433;
      22684: inst = 32'h8220000;
      22685: inst = 32'h10408000;
      22686: inst = 32'hc405434;
      22687: inst = 32'h8220000;
      22688: inst = 32'h10408000;
      22689: inst = 32'hc405435;
      22690: inst = 32'h8220000;
      22691: inst = 32'h10408000;
      22692: inst = 32'hc405436;
      22693: inst = 32'h8220000;
      22694: inst = 32'h10408000;
      22695: inst = 32'hc405437;
      22696: inst = 32'h8220000;
      22697: inst = 32'h10408000;
      22698: inst = 32'hc405438;
      22699: inst = 32'h8220000;
      22700: inst = 32'h10408000;
      22701: inst = 32'hc405439;
      22702: inst = 32'h8220000;
      22703: inst = 32'h10408000;
      22704: inst = 32'hc40543a;
      22705: inst = 32'h8220000;
      22706: inst = 32'h10408000;
      22707: inst = 32'hc40543b;
      22708: inst = 32'h8220000;
      22709: inst = 32'h10408000;
      22710: inst = 32'hc40543c;
      22711: inst = 32'h8220000;
      22712: inst = 32'h10408000;
      22713: inst = 32'hc40543d;
      22714: inst = 32'h8220000;
      22715: inst = 32'h10408000;
      22716: inst = 32'hc40543e;
      22717: inst = 32'h8220000;
      22718: inst = 32'h10408000;
      22719: inst = 32'hc40543f;
      22720: inst = 32'h8220000;
      22721: inst = 32'h10408000;
      22722: inst = 32'hc405440;
      22723: inst = 32'h8220000;
      22724: inst = 32'h10408000;
      22725: inst = 32'hc405441;
      22726: inst = 32'h8220000;
      22727: inst = 32'h10408000;
      22728: inst = 32'hc405442;
      22729: inst = 32'h8220000;
      22730: inst = 32'h10408000;
      22731: inst = 32'hc405443;
      22732: inst = 32'h8220000;
      22733: inst = 32'h10408000;
      22734: inst = 32'hc405444;
      22735: inst = 32'h8220000;
      22736: inst = 32'h10408000;
      22737: inst = 32'hc405445;
      22738: inst = 32'h8220000;
      22739: inst = 32'h10408000;
      22740: inst = 32'hc405446;
      22741: inst = 32'h8220000;
      22742: inst = 32'h10408000;
      22743: inst = 32'hc405447;
      22744: inst = 32'h8220000;
      22745: inst = 32'h10408000;
      22746: inst = 32'hc405448;
      22747: inst = 32'h8220000;
      22748: inst = 32'h10408000;
      22749: inst = 32'hc405449;
      22750: inst = 32'h8220000;
      22751: inst = 32'h10408000;
      22752: inst = 32'hc40544a;
      22753: inst = 32'h8220000;
      22754: inst = 32'h10408000;
      22755: inst = 32'hc40544b;
      22756: inst = 32'h8220000;
      22757: inst = 32'h10408000;
      22758: inst = 32'hc40544c;
      22759: inst = 32'h8220000;
      22760: inst = 32'h10408000;
      22761: inst = 32'hc40544d;
      22762: inst = 32'h8220000;
      22763: inst = 32'h10408000;
      22764: inst = 32'hc40544e;
      22765: inst = 32'h8220000;
      22766: inst = 32'h10408000;
      22767: inst = 32'hc40544f;
      22768: inst = 32'h8220000;
      22769: inst = 32'h10408000;
      22770: inst = 32'hc405450;
      22771: inst = 32'h8220000;
      22772: inst = 32'h10408000;
      22773: inst = 32'hc405451;
      22774: inst = 32'h8220000;
      22775: inst = 32'h10408000;
      22776: inst = 32'hc405452;
      22777: inst = 32'h8220000;
      22778: inst = 32'h10408000;
      22779: inst = 32'hc405453;
      22780: inst = 32'h8220000;
      22781: inst = 32'h10408000;
      22782: inst = 32'hc405454;
      22783: inst = 32'h8220000;
      22784: inst = 32'h10408000;
      22785: inst = 32'hc405455;
      22786: inst = 32'h8220000;
      22787: inst = 32'h10408000;
      22788: inst = 32'hc405456;
      22789: inst = 32'h8220000;
      22790: inst = 32'h10408000;
      22791: inst = 32'hc405457;
      22792: inst = 32'h8220000;
      22793: inst = 32'h10408000;
      22794: inst = 32'hc405458;
      22795: inst = 32'h8220000;
      22796: inst = 32'h10408000;
      22797: inst = 32'hc405459;
      22798: inst = 32'h8220000;
      22799: inst = 32'h10408000;
      22800: inst = 32'hc40545a;
      22801: inst = 32'h8220000;
      22802: inst = 32'h10408000;
      22803: inst = 32'hc40545b;
      22804: inst = 32'h8220000;
      22805: inst = 32'h10408000;
      22806: inst = 32'hc40545c;
      22807: inst = 32'h8220000;
      22808: inst = 32'h10408000;
      22809: inst = 32'hc40545d;
      22810: inst = 32'h8220000;
      22811: inst = 32'h10408000;
      22812: inst = 32'hc40545e;
      22813: inst = 32'h8220000;
      22814: inst = 32'h10408000;
      22815: inst = 32'hc40545f;
      22816: inst = 32'h8220000;
      22817: inst = 32'h10408000;
      22818: inst = 32'hc405460;
      22819: inst = 32'h8220000;
      22820: inst = 32'h10408000;
      22821: inst = 32'hc405461;
      22822: inst = 32'h8220000;
      22823: inst = 32'h10408000;
      22824: inst = 32'hc405462;
      22825: inst = 32'h8220000;
      22826: inst = 32'h10408000;
      22827: inst = 32'hc405463;
      22828: inst = 32'h8220000;
      22829: inst = 32'h10408000;
      22830: inst = 32'hc405464;
      22831: inst = 32'h8220000;
      22832: inst = 32'h10408000;
      22833: inst = 32'hc405465;
      22834: inst = 32'h8220000;
      22835: inst = 32'h10408000;
      22836: inst = 32'hc405466;
      22837: inst = 32'h8220000;
      22838: inst = 32'h10408000;
      22839: inst = 32'hc405467;
      22840: inst = 32'h8220000;
      22841: inst = 32'h10408000;
      22842: inst = 32'hc405468;
      22843: inst = 32'h8220000;
      22844: inst = 32'h10408000;
      22845: inst = 32'hc405469;
      22846: inst = 32'h8220000;
      22847: inst = 32'h10408000;
      22848: inst = 32'hc40546a;
      22849: inst = 32'h8220000;
      22850: inst = 32'h10408000;
      22851: inst = 32'hc40546b;
      22852: inst = 32'h8220000;
      22853: inst = 32'h10408000;
      22854: inst = 32'hc40546c;
      22855: inst = 32'h8220000;
      22856: inst = 32'h10408000;
      22857: inst = 32'hc40546d;
      22858: inst = 32'h8220000;
      22859: inst = 32'h10408000;
      22860: inst = 32'hc40546e;
      22861: inst = 32'h8220000;
      22862: inst = 32'h10408000;
      22863: inst = 32'hc40546f;
      22864: inst = 32'h8220000;
      22865: inst = 32'h10408000;
      22866: inst = 32'hc405470;
      22867: inst = 32'h8220000;
      22868: inst = 32'h10408000;
      22869: inst = 32'hc405471;
      22870: inst = 32'h8220000;
      22871: inst = 32'h10408000;
      22872: inst = 32'hc405472;
      22873: inst = 32'h8220000;
      22874: inst = 32'h10408000;
      22875: inst = 32'hc405473;
      22876: inst = 32'h8220000;
      22877: inst = 32'h10408000;
      22878: inst = 32'hc405474;
      22879: inst = 32'h8220000;
      22880: inst = 32'h10408000;
      22881: inst = 32'hc405475;
      22882: inst = 32'h8220000;
      22883: inst = 32'h10408000;
      22884: inst = 32'hc405476;
      22885: inst = 32'h8220000;
      22886: inst = 32'hc202106;
      22887: inst = 32'h10408000;
      22888: inst = 32'hc404347;
      22889: inst = 32'h8220000;
      22890: inst = 32'h10408000;
      22891: inst = 32'hc404398;
      22892: inst = 32'h8220000;
      22893: inst = 32'h10408000;
      22894: inst = 32'hc4053c7;
      22895: inst = 32'h8220000;
      22896: inst = 32'h10408000;
      22897: inst = 32'hc405418;
      22898: inst = 32'h8220000;
      22899: inst = 32'hc2018c3;
      22900: inst = 32'h10408000;
      22901: inst = 32'hc404348;
      22902: inst = 32'h8220000;
      22903: inst = 32'h10408000;
      22904: inst = 32'hc404349;
      22905: inst = 32'h8220000;
      22906: inst = 32'h10408000;
      22907: inst = 32'hc40434a;
      22908: inst = 32'h8220000;
      22909: inst = 32'h10408000;
      22910: inst = 32'hc40434b;
      22911: inst = 32'h8220000;
      22912: inst = 32'h10408000;
      22913: inst = 32'hc40434c;
      22914: inst = 32'h8220000;
      22915: inst = 32'h10408000;
      22916: inst = 32'hc40434d;
      22917: inst = 32'h8220000;
      22918: inst = 32'h10408000;
      22919: inst = 32'hc40434e;
      22920: inst = 32'h8220000;
      22921: inst = 32'h10408000;
      22922: inst = 32'hc40434f;
      22923: inst = 32'h8220000;
      22924: inst = 32'h10408000;
      22925: inst = 32'hc404350;
      22926: inst = 32'h8220000;
      22927: inst = 32'h10408000;
      22928: inst = 32'hc404351;
      22929: inst = 32'h8220000;
      22930: inst = 32'h10408000;
      22931: inst = 32'hc404352;
      22932: inst = 32'h8220000;
      22933: inst = 32'h10408000;
      22934: inst = 32'hc404353;
      22935: inst = 32'h8220000;
      22936: inst = 32'h10408000;
      22937: inst = 32'hc404354;
      22938: inst = 32'h8220000;
      22939: inst = 32'h10408000;
      22940: inst = 32'hc404355;
      22941: inst = 32'h8220000;
      22942: inst = 32'h10408000;
      22943: inst = 32'hc404356;
      22944: inst = 32'h8220000;
      22945: inst = 32'h10408000;
      22946: inst = 32'hc404357;
      22947: inst = 32'h8220000;
      22948: inst = 32'h10408000;
      22949: inst = 32'hc404358;
      22950: inst = 32'h8220000;
      22951: inst = 32'h10408000;
      22952: inst = 32'hc404359;
      22953: inst = 32'h8220000;
      22954: inst = 32'h10408000;
      22955: inst = 32'hc40435a;
      22956: inst = 32'h8220000;
      22957: inst = 32'h10408000;
      22958: inst = 32'hc40435b;
      22959: inst = 32'h8220000;
      22960: inst = 32'h10408000;
      22961: inst = 32'hc40435c;
      22962: inst = 32'h8220000;
      22963: inst = 32'h10408000;
      22964: inst = 32'hc40435d;
      22965: inst = 32'h8220000;
      22966: inst = 32'h10408000;
      22967: inst = 32'hc40435e;
      22968: inst = 32'h8220000;
      22969: inst = 32'h10408000;
      22970: inst = 32'hc40435f;
      22971: inst = 32'h8220000;
      22972: inst = 32'h10408000;
      22973: inst = 32'hc404360;
      22974: inst = 32'h8220000;
      22975: inst = 32'h10408000;
      22976: inst = 32'hc404361;
      22977: inst = 32'h8220000;
      22978: inst = 32'h10408000;
      22979: inst = 32'hc404362;
      22980: inst = 32'h8220000;
      22981: inst = 32'h10408000;
      22982: inst = 32'hc404363;
      22983: inst = 32'h8220000;
      22984: inst = 32'h10408000;
      22985: inst = 32'hc404364;
      22986: inst = 32'h8220000;
      22987: inst = 32'h10408000;
      22988: inst = 32'hc404365;
      22989: inst = 32'h8220000;
      22990: inst = 32'h10408000;
      22991: inst = 32'hc404366;
      22992: inst = 32'h8220000;
      22993: inst = 32'h10408000;
      22994: inst = 32'hc404367;
      22995: inst = 32'h8220000;
      22996: inst = 32'h10408000;
      22997: inst = 32'hc404368;
      22998: inst = 32'h8220000;
      22999: inst = 32'h10408000;
      23000: inst = 32'hc404369;
      23001: inst = 32'h8220000;
      23002: inst = 32'h10408000;
      23003: inst = 32'hc40436a;
      23004: inst = 32'h8220000;
      23005: inst = 32'h10408000;
      23006: inst = 32'hc40436b;
      23007: inst = 32'h8220000;
      23008: inst = 32'h10408000;
      23009: inst = 32'hc40436c;
      23010: inst = 32'h8220000;
      23011: inst = 32'h10408000;
      23012: inst = 32'hc40436d;
      23013: inst = 32'h8220000;
      23014: inst = 32'h10408000;
      23015: inst = 32'hc40436e;
      23016: inst = 32'h8220000;
      23017: inst = 32'h10408000;
      23018: inst = 32'hc40436f;
      23019: inst = 32'h8220000;
      23020: inst = 32'h10408000;
      23021: inst = 32'hc404370;
      23022: inst = 32'h8220000;
      23023: inst = 32'h10408000;
      23024: inst = 32'hc404371;
      23025: inst = 32'h8220000;
      23026: inst = 32'h10408000;
      23027: inst = 32'hc404372;
      23028: inst = 32'h8220000;
      23029: inst = 32'h10408000;
      23030: inst = 32'hc404373;
      23031: inst = 32'h8220000;
      23032: inst = 32'h10408000;
      23033: inst = 32'hc404374;
      23034: inst = 32'h8220000;
      23035: inst = 32'h10408000;
      23036: inst = 32'hc404375;
      23037: inst = 32'h8220000;
      23038: inst = 32'h10408000;
      23039: inst = 32'hc404376;
      23040: inst = 32'h8220000;
      23041: inst = 32'h10408000;
      23042: inst = 32'hc404377;
      23043: inst = 32'h8220000;
      23044: inst = 32'h10408000;
      23045: inst = 32'hc404378;
      23046: inst = 32'h8220000;
      23047: inst = 32'h10408000;
      23048: inst = 32'hc404379;
      23049: inst = 32'h8220000;
      23050: inst = 32'h10408000;
      23051: inst = 32'hc40437a;
      23052: inst = 32'h8220000;
      23053: inst = 32'h10408000;
      23054: inst = 32'hc40437b;
      23055: inst = 32'h8220000;
      23056: inst = 32'h10408000;
      23057: inst = 32'hc40437c;
      23058: inst = 32'h8220000;
      23059: inst = 32'h10408000;
      23060: inst = 32'hc40437d;
      23061: inst = 32'h8220000;
      23062: inst = 32'h10408000;
      23063: inst = 32'hc40437e;
      23064: inst = 32'h8220000;
      23065: inst = 32'h10408000;
      23066: inst = 32'hc40437f;
      23067: inst = 32'h8220000;
      23068: inst = 32'h10408000;
      23069: inst = 32'hc404380;
      23070: inst = 32'h8220000;
      23071: inst = 32'h10408000;
      23072: inst = 32'hc404381;
      23073: inst = 32'h8220000;
      23074: inst = 32'h10408000;
      23075: inst = 32'hc404382;
      23076: inst = 32'h8220000;
      23077: inst = 32'h10408000;
      23078: inst = 32'hc404383;
      23079: inst = 32'h8220000;
      23080: inst = 32'h10408000;
      23081: inst = 32'hc404384;
      23082: inst = 32'h8220000;
      23083: inst = 32'h10408000;
      23084: inst = 32'hc404385;
      23085: inst = 32'h8220000;
      23086: inst = 32'h10408000;
      23087: inst = 32'hc404386;
      23088: inst = 32'h8220000;
      23089: inst = 32'h10408000;
      23090: inst = 32'hc404387;
      23091: inst = 32'h8220000;
      23092: inst = 32'h10408000;
      23093: inst = 32'hc404388;
      23094: inst = 32'h8220000;
      23095: inst = 32'h10408000;
      23096: inst = 32'hc404389;
      23097: inst = 32'h8220000;
      23098: inst = 32'h10408000;
      23099: inst = 32'hc40438a;
      23100: inst = 32'h8220000;
      23101: inst = 32'h10408000;
      23102: inst = 32'hc40438b;
      23103: inst = 32'h8220000;
      23104: inst = 32'h10408000;
      23105: inst = 32'hc40438c;
      23106: inst = 32'h8220000;
      23107: inst = 32'h10408000;
      23108: inst = 32'hc40438d;
      23109: inst = 32'h8220000;
      23110: inst = 32'h10408000;
      23111: inst = 32'hc40438e;
      23112: inst = 32'h8220000;
      23113: inst = 32'h10408000;
      23114: inst = 32'hc40438f;
      23115: inst = 32'h8220000;
      23116: inst = 32'h10408000;
      23117: inst = 32'hc404390;
      23118: inst = 32'h8220000;
      23119: inst = 32'h10408000;
      23120: inst = 32'hc404391;
      23121: inst = 32'h8220000;
      23122: inst = 32'h10408000;
      23123: inst = 32'hc404392;
      23124: inst = 32'h8220000;
      23125: inst = 32'h10408000;
      23126: inst = 32'hc404393;
      23127: inst = 32'h8220000;
      23128: inst = 32'h10408000;
      23129: inst = 32'hc404394;
      23130: inst = 32'h8220000;
      23131: inst = 32'h10408000;
      23132: inst = 32'hc404395;
      23133: inst = 32'h8220000;
      23134: inst = 32'h10408000;
      23135: inst = 32'hc404396;
      23136: inst = 32'h8220000;
      23137: inst = 32'h10408000;
      23138: inst = 32'hc404397;
      23139: inst = 32'h8220000;
      23140: inst = 32'h10408000;
      23141: inst = 32'hc4043a7;
      23142: inst = 32'h8220000;
      23143: inst = 32'h10408000;
      23144: inst = 32'hc4043a8;
      23145: inst = 32'h8220000;
      23146: inst = 32'h10408000;
      23147: inst = 32'hc4043a9;
      23148: inst = 32'h8220000;
      23149: inst = 32'h10408000;
      23150: inst = 32'hc4043aa;
      23151: inst = 32'h8220000;
      23152: inst = 32'h10408000;
      23153: inst = 32'hc4043ab;
      23154: inst = 32'h8220000;
      23155: inst = 32'h10408000;
      23156: inst = 32'hc4043ac;
      23157: inst = 32'h8220000;
      23158: inst = 32'h10408000;
      23159: inst = 32'hc4043ad;
      23160: inst = 32'h8220000;
      23161: inst = 32'h10408000;
      23162: inst = 32'hc4043ae;
      23163: inst = 32'h8220000;
      23164: inst = 32'h10408000;
      23165: inst = 32'hc4043af;
      23166: inst = 32'h8220000;
      23167: inst = 32'h10408000;
      23168: inst = 32'hc4043b0;
      23169: inst = 32'h8220000;
      23170: inst = 32'h10408000;
      23171: inst = 32'hc4043b1;
      23172: inst = 32'h8220000;
      23173: inst = 32'h10408000;
      23174: inst = 32'hc4043b2;
      23175: inst = 32'h8220000;
      23176: inst = 32'h10408000;
      23177: inst = 32'hc4043b3;
      23178: inst = 32'h8220000;
      23179: inst = 32'h10408000;
      23180: inst = 32'hc4043b4;
      23181: inst = 32'h8220000;
      23182: inst = 32'h10408000;
      23183: inst = 32'hc4043b5;
      23184: inst = 32'h8220000;
      23185: inst = 32'h10408000;
      23186: inst = 32'hc4043b6;
      23187: inst = 32'h8220000;
      23188: inst = 32'h10408000;
      23189: inst = 32'hc4043b7;
      23190: inst = 32'h8220000;
      23191: inst = 32'h10408000;
      23192: inst = 32'hc4043b8;
      23193: inst = 32'h8220000;
      23194: inst = 32'h10408000;
      23195: inst = 32'hc4043b9;
      23196: inst = 32'h8220000;
      23197: inst = 32'h10408000;
      23198: inst = 32'hc4043ba;
      23199: inst = 32'h8220000;
      23200: inst = 32'h10408000;
      23201: inst = 32'hc4043bb;
      23202: inst = 32'h8220000;
      23203: inst = 32'h10408000;
      23204: inst = 32'hc4043bc;
      23205: inst = 32'h8220000;
      23206: inst = 32'h10408000;
      23207: inst = 32'hc4043bd;
      23208: inst = 32'h8220000;
      23209: inst = 32'h10408000;
      23210: inst = 32'hc4043be;
      23211: inst = 32'h8220000;
      23212: inst = 32'h10408000;
      23213: inst = 32'hc4043bf;
      23214: inst = 32'h8220000;
      23215: inst = 32'h10408000;
      23216: inst = 32'hc4043c0;
      23217: inst = 32'h8220000;
      23218: inst = 32'h10408000;
      23219: inst = 32'hc4043c1;
      23220: inst = 32'h8220000;
      23221: inst = 32'h10408000;
      23222: inst = 32'hc4043c2;
      23223: inst = 32'h8220000;
      23224: inst = 32'h10408000;
      23225: inst = 32'hc4043c3;
      23226: inst = 32'h8220000;
      23227: inst = 32'h10408000;
      23228: inst = 32'hc4043c4;
      23229: inst = 32'h8220000;
      23230: inst = 32'h10408000;
      23231: inst = 32'hc4043c5;
      23232: inst = 32'h8220000;
      23233: inst = 32'h10408000;
      23234: inst = 32'hc4043c6;
      23235: inst = 32'h8220000;
      23236: inst = 32'h10408000;
      23237: inst = 32'hc4043c7;
      23238: inst = 32'h8220000;
      23239: inst = 32'h10408000;
      23240: inst = 32'hc4043c8;
      23241: inst = 32'h8220000;
      23242: inst = 32'h10408000;
      23243: inst = 32'hc4043c9;
      23244: inst = 32'h8220000;
      23245: inst = 32'h10408000;
      23246: inst = 32'hc4043ca;
      23247: inst = 32'h8220000;
      23248: inst = 32'h10408000;
      23249: inst = 32'hc4043cb;
      23250: inst = 32'h8220000;
      23251: inst = 32'h10408000;
      23252: inst = 32'hc4043cc;
      23253: inst = 32'h8220000;
      23254: inst = 32'h10408000;
      23255: inst = 32'hc4043cd;
      23256: inst = 32'h8220000;
      23257: inst = 32'h10408000;
      23258: inst = 32'hc4043ce;
      23259: inst = 32'h8220000;
      23260: inst = 32'h10408000;
      23261: inst = 32'hc4043cf;
      23262: inst = 32'h8220000;
      23263: inst = 32'h10408000;
      23264: inst = 32'hc4043d0;
      23265: inst = 32'h8220000;
      23266: inst = 32'h10408000;
      23267: inst = 32'hc4043d1;
      23268: inst = 32'h8220000;
      23269: inst = 32'h10408000;
      23270: inst = 32'hc4043d2;
      23271: inst = 32'h8220000;
      23272: inst = 32'h10408000;
      23273: inst = 32'hc4043d3;
      23274: inst = 32'h8220000;
      23275: inst = 32'h10408000;
      23276: inst = 32'hc4043d4;
      23277: inst = 32'h8220000;
      23278: inst = 32'h10408000;
      23279: inst = 32'hc4043d5;
      23280: inst = 32'h8220000;
      23281: inst = 32'h10408000;
      23282: inst = 32'hc4043d6;
      23283: inst = 32'h8220000;
      23284: inst = 32'h10408000;
      23285: inst = 32'hc4043d7;
      23286: inst = 32'h8220000;
      23287: inst = 32'h10408000;
      23288: inst = 32'hc4043d8;
      23289: inst = 32'h8220000;
      23290: inst = 32'h10408000;
      23291: inst = 32'hc4043d9;
      23292: inst = 32'h8220000;
      23293: inst = 32'h10408000;
      23294: inst = 32'hc4043da;
      23295: inst = 32'h8220000;
      23296: inst = 32'h10408000;
      23297: inst = 32'hc4043db;
      23298: inst = 32'h8220000;
      23299: inst = 32'h10408000;
      23300: inst = 32'hc4043dc;
      23301: inst = 32'h8220000;
      23302: inst = 32'h10408000;
      23303: inst = 32'hc4043dd;
      23304: inst = 32'h8220000;
      23305: inst = 32'h10408000;
      23306: inst = 32'hc4043de;
      23307: inst = 32'h8220000;
      23308: inst = 32'h10408000;
      23309: inst = 32'hc4043df;
      23310: inst = 32'h8220000;
      23311: inst = 32'h10408000;
      23312: inst = 32'hc4043e0;
      23313: inst = 32'h8220000;
      23314: inst = 32'h10408000;
      23315: inst = 32'hc4043e1;
      23316: inst = 32'h8220000;
      23317: inst = 32'h10408000;
      23318: inst = 32'hc4043e2;
      23319: inst = 32'h8220000;
      23320: inst = 32'h10408000;
      23321: inst = 32'hc4043e3;
      23322: inst = 32'h8220000;
      23323: inst = 32'h10408000;
      23324: inst = 32'hc4043e4;
      23325: inst = 32'h8220000;
      23326: inst = 32'h10408000;
      23327: inst = 32'hc4043e5;
      23328: inst = 32'h8220000;
      23329: inst = 32'h10408000;
      23330: inst = 32'hc4043e6;
      23331: inst = 32'h8220000;
      23332: inst = 32'h10408000;
      23333: inst = 32'hc4043e7;
      23334: inst = 32'h8220000;
      23335: inst = 32'h10408000;
      23336: inst = 32'hc4043e8;
      23337: inst = 32'h8220000;
      23338: inst = 32'h10408000;
      23339: inst = 32'hc4043e9;
      23340: inst = 32'h8220000;
      23341: inst = 32'h10408000;
      23342: inst = 32'hc4043ea;
      23343: inst = 32'h8220000;
      23344: inst = 32'h10408000;
      23345: inst = 32'hc4043eb;
      23346: inst = 32'h8220000;
      23347: inst = 32'h10408000;
      23348: inst = 32'hc4043ec;
      23349: inst = 32'h8220000;
      23350: inst = 32'h10408000;
      23351: inst = 32'hc4043ed;
      23352: inst = 32'h8220000;
      23353: inst = 32'h10408000;
      23354: inst = 32'hc4043ee;
      23355: inst = 32'h8220000;
      23356: inst = 32'h10408000;
      23357: inst = 32'hc4043ef;
      23358: inst = 32'h8220000;
      23359: inst = 32'h10408000;
      23360: inst = 32'hc4043f0;
      23361: inst = 32'h8220000;
      23362: inst = 32'h10408000;
      23363: inst = 32'hc4043f1;
      23364: inst = 32'h8220000;
      23365: inst = 32'h10408000;
      23366: inst = 32'hc4043f2;
      23367: inst = 32'h8220000;
      23368: inst = 32'h10408000;
      23369: inst = 32'hc4043f3;
      23370: inst = 32'h8220000;
      23371: inst = 32'h10408000;
      23372: inst = 32'hc4043f4;
      23373: inst = 32'h8220000;
      23374: inst = 32'h10408000;
      23375: inst = 32'hc4043f5;
      23376: inst = 32'h8220000;
      23377: inst = 32'h10408000;
      23378: inst = 32'hc4043f6;
      23379: inst = 32'h8220000;
      23380: inst = 32'h10408000;
      23381: inst = 32'hc4043f7;
      23382: inst = 32'h8220000;
      23383: inst = 32'h10408000;
      23384: inst = 32'hc4043f8;
      23385: inst = 32'h8220000;
      23386: inst = 32'h10408000;
      23387: inst = 32'hc404407;
      23388: inst = 32'h8220000;
      23389: inst = 32'h10408000;
      23390: inst = 32'hc404408;
      23391: inst = 32'h8220000;
      23392: inst = 32'h10408000;
      23393: inst = 32'hc404409;
      23394: inst = 32'h8220000;
      23395: inst = 32'h10408000;
      23396: inst = 32'hc40440a;
      23397: inst = 32'h8220000;
      23398: inst = 32'h10408000;
      23399: inst = 32'hc40440b;
      23400: inst = 32'h8220000;
      23401: inst = 32'h10408000;
      23402: inst = 32'hc40440c;
      23403: inst = 32'h8220000;
      23404: inst = 32'h10408000;
      23405: inst = 32'hc40440d;
      23406: inst = 32'h8220000;
      23407: inst = 32'h10408000;
      23408: inst = 32'hc40440e;
      23409: inst = 32'h8220000;
      23410: inst = 32'h10408000;
      23411: inst = 32'hc40440f;
      23412: inst = 32'h8220000;
      23413: inst = 32'h10408000;
      23414: inst = 32'hc404410;
      23415: inst = 32'h8220000;
      23416: inst = 32'h10408000;
      23417: inst = 32'hc404411;
      23418: inst = 32'h8220000;
      23419: inst = 32'h10408000;
      23420: inst = 32'hc404412;
      23421: inst = 32'h8220000;
      23422: inst = 32'h10408000;
      23423: inst = 32'hc404413;
      23424: inst = 32'h8220000;
      23425: inst = 32'h10408000;
      23426: inst = 32'hc404414;
      23427: inst = 32'h8220000;
      23428: inst = 32'h10408000;
      23429: inst = 32'hc404415;
      23430: inst = 32'h8220000;
      23431: inst = 32'h10408000;
      23432: inst = 32'hc404416;
      23433: inst = 32'h8220000;
      23434: inst = 32'h10408000;
      23435: inst = 32'hc404417;
      23436: inst = 32'h8220000;
      23437: inst = 32'h10408000;
      23438: inst = 32'hc404418;
      23439: inst = 32'h8220000;
      23440: inst = 32'h10408000;
      23441: inst = 32'hc404419;
      23442: inst = 32'h8220000;
      23443: inst = 32'h10408000;
      23444: inst = 32'hc40441a;
      23445: inst = 32'h8220000;
      23446: inst = 32'h10408000;
      23447: inst = 32'hc40441b;
      23448: inst = 32'h8220000;
      23449: inst = 32'h10408000;
      23450: inst = 32'hc40441c;
      23451: inst = 32'h8220000;
      23452: inst = 32'h10408000;
      23453: inst = 32'hc40441d;
      23454: inst = 32'h8220000;
      23455: inst = 32'h10408000;
      23456: inst = 32'hc40441e;
      23457: inst = 32'h8220000;
      23458: inst = 32'h10408000;
      23459: inst = 32'hc40441f;
      23460: inst = 32'h8220000;
      23461: inst = 32'h10408000;
      23462: inst = 32'hc404420;
      23463: inst = 32'h8220000;
      23464: inst = 32'h10408000;
      23465: inst = 32'hc404421;
      23466: inst = 32'h8220000;
      23467: inst = 32'h10408000;
      23468: inst = 32'hc404422;
      23469: inst = 32'h8220000;
      23470: inst = 32'h10408000;
      23471: inst = 32'hc404423;
      23472: inst = 32'h8220000;
      23473: inst = 32'h10408000;
      23474: inst = 32'hc404424;
      23475: inst = 32'h8220000;
      23476: inst = 32'h10408000;
      23477: inst = 32'hc404425;
      23478: inst = 32'h8220000;
      23479: inst = 32'h10408000;
      23480: inst = 32'hc404426;
      23481: inst = 32'h8220000;
      23482: inst = 32'h10408000;
      23483: inst = 32'hc404427;
      23484: inst = 32'h8220000;
      23485: inst = 32'h10408000;
      23486: inst = 32'hc404428;
      23487: inst = 32'h8220000;
      23488: inst = 32'h10408000;
      23489: inst = 32'hc404429;
      23490: inst = 32'h8220000;
      23491: inst = 32'h10408000;
      23492: inst = 32'hc40442a;
      23493: inst = 32'h8220000;
      23494: inst = 32'h10408000;
      23495: inst = 32'hc40442b;
      23496: inst = 32'h8220000;
      23497: inst = 32'h10408000;
      23498: inst = 32'hc40442c;
      23499: inst = 32'h8220000;
      23500: inst = 32'h10408000;
      23501: inst = 32'hc40442d;
      23502: inst = 32'h8220000;
      23503: inst = 32'h10408000;
      23504: inst = 32'hc40442e;
      23505: inst = 32'h8220000;
      23506: inst = 32'h10408000;
      23507: inst = 32'hc40442f;
      23508: inst = 32'h8220000;
      23509: inst = 32'h10408000;
      23510: inst = 32'hc404430;
      23511: inst = 32'h8220000;
      23512: inst = 32'h10408000;
      23513: inst = 32'hc404431;
      23514: inst = 32'h8220000;
      23515: inst = 32'h10408000;
      23516: inst = 32'hc404432;
      23517: inst = 32'h8220000;
      23518: inst = 32'h10408000;
      23519: inst = 32'hc404433;
      23520: inst = 32'h8220000;
      23521: inst = 32'h10408000;
      23522: inst = 32'hc404434;
      23523: inst = 32'h8220000;
      23524: inst = 32'h10408000;
      23525: inst = 32'hc404435;
      23526: inst = 32'h8220000;
      23527: inst = 32'h10408000;
      23528: inst = 32'hc404436;
      23529: inst = 32'h8220000;
      23530: inst = 32'h10408000;
      23531: inst = 32'hc404437;
      23532: inst = 32'h8220000;
      23533: inst = 32'h10408000;
      23534: inst = 32'hc404438;
      23535: inst = 32'h8220000;
      23536: inst = 32'h10408000;
      23537: inst = 32'hc404439;
      23538: inst = 32'h8220000;
      23539: inst = 32'h10408000;
      23540: inst = 32'hc40443a;
      23541: inst = 32'h8220000;
      23542: inst = 32'h10408000;
      23543: inst = 32'hc40443b;
      23544: inst = 32'h8220000;
      23545: inst = 32'h10408000;
      23546: inst = 32'hc40443c;
      23547: inst = 32'h8220000;
      23548: inst = 32'h10408000;
      23549: inst = 32'hc40443d;
      23550: inst = 32'h8220000;
      23551: inst = 32'h10408000;
      23552: inst = 32'hc40443e;
      23553: inst = 32'h8220000;
      23554: inst = 32'h10408000;
      23555: inst = 32'hc40443f;
      23556: inst = 32'h8220000;
      23557: inst = 32'h10408000;
      23558: inst = 32'hc404440;
      23559: inst = 32'h8220000;
      23560: inst = 32'h10408000;
      23561: inst = 32'hc404441;
      23562: inst = 32'h8220000;
      23563: inst = 32'h10408000;
      23564: inst = 32'hc404442;
      23565: inst = 32'h8220000;
      23566: inst = 32'h10408000;
      23567: inst = 32'hc404443;
      23568: inst = 32'h8220000;
      23569: inst = 32'h10408000;
      23570: inst = 32'hc404444;
      23571: inst = 32'h8220000;
      23572: inst = 32'h10408000;
      23573: inst = 32'hc404445;
      23574: inst = 32'h8220000;
      23575: inst = 32'h10408000;
      23576: inst = 32'hc404446;
      23577: inst = 32'h8220000;
      23578: inst = 32'h10408000;
      23579: inst = 32'hc404447;
      23580: inst = 32'h8220000;
      23581: inst = 32'h10408000;
      23582: inst = 32'hc404448;
      23583: inst = 32'h8220000;
      23584: inst = 32'h10408000;
      23585: inst = 32'hc404449;
      23586: inst = 32'h8220000;
      23587: inst = 32'h10408000;
      23588: inst = 32'hc40444a;
      23589: inst = 32'h8220000;
      23590: inst = 32'h10408000;
      23591: inst = 32'hc40444b;
      23592: inst = 32'h8220000;
      23593: inst = 32'h10408000;
      23594: inst = 32'hc40444c;
      23595: inst = 32'h8220000;
      23596: inst = 32'h10408000;
      23597: inst = 32'hc40444d;
      23598: inst = 32'h8220000;
      23599: inst = 32'h10408000;
      23600: inst = 32'hc40444e;
      23601: inst = 32'h8220000;
      23602: inst = 32'h10408000;
      23603: inst = 32'hc40444f;
      23604: inst = 32'h8220000;
      23605: inst = 32'h10408000;
      23606: inst = 32'hc404450;
      23607: inst = 32'h8220000;
      23608: inst = 32'h10408000;
      23609: inst = 32'hc404451;
      23610: inst = 32'h8220000;
      23611: inst = 32'h10408000;
      23612: inst = 32'hc404452;
      23613: inst = 32'h8220000;
      23614: inst = 32'h10408000;
      23615: inst = 32'hc404453;
      23616: inst = 32'h8220000;
      23617: inst = 32'h10408000;
      23618: inst = 32'hc404454;
      23619: inst = 32'h8220000;
      23620: inst = 32'h10408000;
      23621: inst = 32'hc404455;
      23622: inst = 32'h8220000;
      23623: inst = 32'h10408000;
      23624: inst = 32'hc404456;
      23625: inst = 32'h8220000;
      23626: inst = 32'h10408000;
      23627: inst = 32'hc404457;
      23628: inst = 32'h8220000;
      23629: inst = 32'h10408000;
      23630: inst = 32'hc404458;
      23631: inst = 32'h8220000;
      23632: inst = 32'h10408000;
      23633: inst = 32'hc404467;
      23634: inst = 32'h8220000;
      23635: inst = 32'h10408000;
      23636: inst = 32'hc404468;
      23637: inst = 32'h8220000;
      23638: inst = 32'h10408000;
      23639: inst = 32'hc404469;
      23640: inst = 32'h8220000;
      23641: inst = 32'h10408000;
      23642: inst = 32'hc40446a;
      23643: inst = 32'h8220000;
      23644: inst = 32'h10408000;
      23645: inst = 32'hc40446b;
      23646: inst = 32'h8220000;
      23647: inst = 32'h10408000;
      23648: inst = 32'hc40446c;
      23649: inst = 32'h8220000;
      23650: inst = 32'h10408000;
      23651: inst = 32'hc40446d;
      23652: inst = 32'h8220000;
      23653: inst = 32'h10408000;
      23654: inst = 32'hc40446e;
      23655: inst = 32'h8220000;
      23656: inst = 32'h10408000;
      23657: inst = 32'hc40446f;
      23658: inst = 32'h8220000;
      23659: inst = 32'h10408000;
      23660: inst = 32'hc404470;
      23661: inst = 32'h8220000;
      23662: inst = 32'h10408000;
      23663: inst = 32'hc404471;
      23664: inst = 32'h8220000;
      23665: inst = 32'h10408000;
      23666: inst = 32'hc404472;
      23667: inst = 32'h8220000;
      23668: inst = 32'h10408000;
      23669: inst = 32'hc404473;
      23670: inst = 32'h8220000;
      23671: inst = 32'h10408000;
      23672: inst = 32'hc404474;
      23673: inst = 32'h8220000;
      23674: inst = 32'h10408000;
      23675: inst = 32'hc404475;
      23676: inst = 32'h8220000;
      23677: inst = 32'h10408000;
      23678: inst = 32'hc404476;
      23679: inst = 32'h8220000;
      23680: inst = 32'h10408000;
      23681: inst = 32'hc404477;
      23682: inst = 32'h8220000;
      23683: inst = 32'h10408000;
      23684: inst = 32'hc404478;
      23685: inst = 32'h8220000;
      23686: inst = 32'h10408000;
      23687: inst = 32'hc404479;
      23688: inst = 32'h8220000;
      23689: inst = 32'h10408000;
      23690: inst = 32'hc40447a;
      23691: inst = 32'h8220000;
      23692: inst = 32'h10408000;
      23693: inst = 32'hc40447b;
      23694: inst = 32'h8220000;
      23695: inst = 32'h10408000;
      23696: inst = 32'hc40447c;
      23697: inst = 32'h8220000;
      23698: inst = 32'h10408000;
      23699: inst = 32'hc40447d;
      23700: inst = 32'h8220000;
      23701: inst = 32'h10408000;
      23702: inst = 32'hc40447e;
      23703: inst = 32'h8220000;
      23704: inst = 32'h10408000;
      23705: inst = 32'hc40447f;
      23706: inst = 32'h8220000;
      23707: inst = 32'h10408000;
      23708: inst = 32'hc404480;
      23709: inst = 32'h8220000;
      23710: inst = 32'h10408000;
      23711: inst = 32'hc404481;
      23712: inst = 32'h8220000;
      23713: inst = 32'h10408000;
      23714: inst = 32'hc404482;
      23715: inst = 32'h8220000;
      23716: inst = 32'h10408000;
      23717: inst = 32'hc404483;
      23718: inst = 32'h8220000;
      23719: inst = 32'h10408000;
      23720: inst = 32'hc404484;
      23721: inst = 32'h8220000;
      23722: inst = 32'h10408000;
      23723: inst = 32'hc404485;
      23724: inst = 32'h8220000;
      23725: inst = 32'h10408000;
      23726: inst = 32'hc404486;
      23727: inst = 32'h8220000;
      23728: inst = 32'h10408000;
      23729: inst = 32'hc404487;
      23730: inst = 32'h8220000;
      23731: inst = 32'h10408000;
      23732: inst = 32'hc404488;
      23733: inst = 32'h8220000;
      23734: inst = 32'h10408000;
      23735: inst = 32'hc404489;
      23736: inst = 32'h8220000;
      23737: inst = 32'h10408000;
      23738: inst = 32'hc40448a;
      23739: inst = 32'h8220000;
      23740: inst = 32'h10408000;
      23741: inst = 32'hc40448b;
      23742: inst = 32'h8220000;
      23743: inst = 32'h10408000;
      23744: inst = 32'hc40448c;
      23745: inst = 32'h8220000;
      23746: inst = 32'h10408000;
      23747: inst = 32'hc40448d;
      23748: inst = 32'h8220000;
      23749: inst = 32'h10408000;
      23750: inst = 32'hc40448e;
      23751: inst = 32'h8220000;
      23752: inst = 32'h10408000;
      23753: inst = 32'hc40448f;
      23754: inst = 32'h8220000;
      23755: inst = 32'h10408000;
      23756: inst = 32'hc404490;
      23757: inst = 32'h8220000;
      23758: inst = 32'h10408000;
      23759: inst = 32'hc404491;
      23760: inst = 32'h8220000;
      23761: inst = 32'h10408000;
      23762: inst = 32'hc404492;
      23763: inst = 32'h8220000;
      23764: inst = 32'h10408000;
      23765: inst = 32'hc404493;
      23766: inst = 32'h8220000;
      23767: inst = 32'h10408000;
      23768: inst = 32'hc404494;
      23769: inst = 32'h8220000;
      23770: inst = 32'h10408000;
      23771: inst = 32'hc404495;
      23772: inst = 32'h8220000;
      23773: inst = 32'h10408000;
      23774: inst = 32'hc404496;
      23775: inst = 32'h8220000;
      23776: inst = 32'h10408000;
      23777: inst = 32'hc404497;
      23778: inst = 32'h8220000;
      23779: inst = 32'h10408000;
      23780: inst = 32'hc404498;
      23781: inst = 32'h8220000;
      23782: inst = 32'h10408000;
      23783: inst = 32'hc404499;
      23784: inst = 32'h8220000;
      23785: inst = 32'h10408000;
      23786: inst = 32'hc40449a;
      23787: inst = 32'h8220000;
      23788: inst = 32'h10408000;
      23789: inst = 32'hc40449b;
      23790: inst = 32'h8220000;
      23791: inst = 32'h10408000;
      23792: inst = 32'hc40449c;
      23793: inst = 32'h8220000;
      23794: inst = 32'h10408000;
      23795: inst = 32'hc40449d;
      23796: inst = 32'h8220000;
      23797: inst = 32'h10408000;
      23798: inst = 32'hc40449e;
      23799: inst = 32'h8220000;
      23800: inst = 32'h10408000;
      23801: inst = 32'hc40449f;
      23802: inst = 32'h8220000;
      23803: inst = 32'h10408000;
      23804: inst = 32'hc4044a0;
      23805: inst = 32'h8220000;
      23806: inst = 32'h10408000;
      23807: inst = 32'hc4044a1;
      23808: inst = 32'h8220000;
      23809: inst = 32'h10408000;
      23810: inst = 32'hc4044a2;
      23811: inst = 32'h8220000;
      23812: inst = 32'h10408000;
      23813: inst = 32'hc4044a3;
      23814: inst = 32'h8220000;
      23815: inst = 32'h10408000;
      23816: inst = 32'hc4044a4;
      23817: inst = 32'h8220000;
      23818: inst = 32'h10408000;
      23819: inst = 32'hc4044a5;
      23820: inst = 32'h8220000;
      23821: inst = 32'h10408000;
      23822: inst = 32'hc4044a6;
      23823: inst = 32'h8220000;
      23824: inst = 32'h10408000;
      23825: inst = 32'hc4044a7;
      23826: inst = 32'h8220000;
      23827: inst = 32'h10408000;
      23828: inst = 32'hc4044a8;
      23829: inst = 32'h8220000;
      23830: inst = 32'h10408000;
      23831: inst = 32'hc4044a9;
      23832: inst = 32'h8220000;
      23833: inst = 32'h10408000;
      23834: inst = 32'hc4044aa;
      23835: inst = 32'h8220000;
      23836: inst = 32'h10408000;
      23837: inst = 32'hc4044ab;
      23838: inst = 32'h8220000;
      23839: inst = 32'h10408000;
      23840: inst = 32'hc4044ac;
      23841: inst = 32'h8220000;
      23842: inst = 32'h10408000;
      23843: inst = 32'hc4044ad;
      23844: inst = 32'h8220000;
      23845: inst = 32'h10408000;
      23846: inst = 32'hc4044ae;
      23847: inst = 32'h8220000;
      23848: inst = 32'h10408000;
      23849: inst = 32'hc4044af;
      23850: inst = 32'h8220000;
      23851: inst = 32'h10408000;
      23852: inst = 32'hc4044b0;
      23853: inst = 32'h8220000;
      23854: inst = 32'h10408000;
      23855: inst = 32'hc4044b1;
      23856: inst = 32'h8220000;
      23857: inst = 32'h10408000;
      23858: inst = 32'hc4044b2;
      23859: inst = 32'h8220000;
      23860: inst = 32'h10408000;
      23861: inst = 32'hc4044b3;
      23862: inst = 32'h8220000;
      23863: inst = 32'h10408000;
      23864: inst = 32'hc4044b4;
      23865: inst = 32'h8220000;
      23866: inst = 32'h10408000;
      23867: inst = 32'hc4044b5;
      23868: inst = 32'h8220000;
      23869: inst = 32'h10408000;
      23870: inst = 32'hc4044b6;
      23871: inst = 32'h8220000;
      23872: inst = 32'h10408000;
      23873: inst = 32'hc4044b7;
      23874: inst = 32'h8220000;
      23875: inst = 32'h10408000;
      23876: inst = 32'hc4044b8;
      23877: inst = 32'h8220000;
      23878: inst = 32'h10408000;
      23879: inst = 32'hc4044c7;
      23880: inst = 32'h8220000;
      23881: inst = 32'h10408000;
      23882: inst = 32'hc4044c8;
      23883: inst = 32'h8220000;
      23884: inst = 32'h10408000;
      23885: inst = 32'hc4044c9;
      23886: inst = 32'h8220000;
      23887: inst = 32'h10408000;
      23888: inst = 32'hc4044ca;
      23889: inst = 32'h8220000;
      23890: inst = 32'h10408000;
      23891: inst = 32'hc4044cb;
      23892: inst = 32'h8220000;
      23893: inst = 32'h10408000;
      23894: inst = 32'hc4044cc;
      23895: inst = 32'h8220000;
      23896: inst = 32'h10408000;
      23897: inst = 32'hc4044cd;
      23898: inst = 32'h8220000;
      23899: inst = 32'h10408000;
      23900: inst = 32'hc4044ce;
      23901: inst = 32'h8220000;
      23902: inst = 32'h10408000;
      23903: inst = 32'hc4044cf;
      23904: inst = 32'h8220000;
      23905: inst = 32'h10408000;
      23906: inst = 32'hc4044d0;
      23907: inst = 32'h8220000;
      23908: inst = 32'h10408000;
      23909: inst = 32'hc4044d1;
      23910: inst = 32'h8220000;
      23911: inst = 32'h10408000;
      23912: inst = 32'hc4044d2;
      23913: inst = 32'h8220000;
      23914: inst = 32'h10408000;
      23915: inst = 32'hc4044d3;
      23916: inst = 32'h8220000;
      23917: inst = 32'h10408000;
      23918: inst = 32'hc4044d4;
      23919: inst = 32'h8220000;
      23920: inst = 32'h10408000;
      23921: inst = 32'hc4044d5;
      23922: inst = 32'h8220000;
      23923: inst = 32'h10408000;
      23924: inst = 32'hc4044d6;
      23925: inst = 32'h8220000;
      23926: inst = 32'h10408000;
      23927: inst = 32'hc4044d7;
      23928: inst = 32'h8220000;
      23929: inst = 32'h10408000;
      23930: inst = 32'hc4044d8;
      23931: inst = 32'h8220000;
      23932: inst = 32'h10408000;
      23933: inst = 32'hc4044d9;
      23934: inst = 32'h8220000;
      23935: inst = 32'h10408000;
      23936: inst = 32'hc4044da;
      23937: inst = 32'h8220000;
      23938: inst = 32'h10408000;
      23939: inst = 32'hc4044db;
      23940: inst = 32'h8220000;
      23941: inst = 32'h10408000;
      23942: inst = 32'hc4044dc;
      23943: inst = 32'h8220000;
      23944: inst = 32'h10408000;
      23945: inst = 32'hc4044dd;
      23946: inst = 32'h8220000;
      23947: inst = 32'h10408000;
      23948: inst = 32'hc4044de;
      23949: inst = 32'h8220000;
      23950: inst = 32'h10408000;
      23951: inst = 32'hc4044df;
      23952: inst = 32'h8220000;
      23953: inst = 32'h10408000;
      23954: inst = 32'hc4044e0;
      23955: inst = 32'h8220000;
      23956: inst = 32'h10408000;
      23957: inst = 32'hc4044e1;
      23958: inst = 32'h8220000;
      23959: inst = 32'h10408000;
      23960: inst = 32'hc4044e2;
      23961: inst = 32'h8220000;
      23962: inst = 32'h10408000;
      23963: inst = 32'hc4044e3;
      23964: inst = 32'h8220000;
      23965: inst = 32'h10408000;
      23966: inst = 32'hc4044e4;
      23967: inst = 32'h8220000;
      23968: inst = 32'h10408000;
      23969: inst = 32'hc4044e5;
      23970: inst = 32'h8220000;
      23971: inst = 32'h10408000;
      23972: inst = 32'hc4044e6;
      23973: inst = 32'h8220000;
      23974: inst = 32'h10408000;
      23975: inst = 32'hc4044e7;
      23976: inst = 32'h8220000;
      23977: inst = 32'h10408000;
      23978: inst = 32'hc4044e8;
      23979: inst = 32'h8220000;
      23980: inst = 32'h10408000;
      23981: inst = 32'hc4044e9;
      23982: inst = 32'h8220000;
      23983: inst = 32'h10408000;
      23984: inst = 32'hc4044ea;
      23985: inst = 32'h8220000;
      23986: inst = 32'h10408000;
      23987: inst = 32'hc4044eb;
      23988: inst = 32'h8220000;
      23989: inst = 32'h10408000;
      23990: inst = 32'hc4044ec;
      23991: inst = 32'h8220000;
      23992: inst = 32'h10408000;
      23993: inst = 32'hc4044ed;
      23994: inst = 32'h8220000;
      23995: inst = 32'h10408000;
      23996: inst = 32'hc4044ee;
      23997: inst = 32'h8220000;
      23998: inst = 32'h10408000;
      23999: inst = 32'hc4044ef;
      24000: inst = 32'h8220000;
      24001: inst = 32'h10408000;
      24002: inst = 32'hc4044f0;
      24003: inst = 32'h8220000;
      24004: inst = 32'h10408000;
      24005: inst = 32'hc4044f1;
      24006: inst = 32'h8220000;
      24007: inst = 32'h10408000;
      24008: inst = 32'hc4044f2;
      24009: inst = 32'h8220000;
      24010: inst = 32'h10408000;
      24011: inst = 32'hc4044f3;
      24012: inst = 32'h8220000;
      24013: inst = 32'h10408000;
      24014: inst = 32'hc4044f4;
      24015: inst = 32'h8220000;
      24016: inst = 32'h10408000;
      24017: inst = 32'hc4044f5;
      24018: inst = 32'h8220000;
      24019: inst = 32'h10408000;
      24020: inst = 32'hc4044f6;
      24021: inst = 32'h8220000;
      24022: inst = 32'h10408000;
      24023: inst = 32'hc4044f7;
      24024: inst = 32'h8220000;
      24025: inst = 32'h10408000;
      24026: inst = 32'hc4044f8;
      24027: inst = 32'h8220000;
      24028: inst = 32'h10408000;
      24029: inst = 32'hc4044f9;
      24030: inst = 32'h8220000;
      24031: inst = 32'h10408000;
      24032: inst = 32'hc4044fa;
      24033: inst = 32'h8220000;
      24034: inst = 32'h10408000;
      24035: inst = 32'hc4044fb;
      24036: inst = 32'h8220000;
      24037: inst = 32'h10408000;
      24038: inst = 32'hc4044fc;
      24039: inst = 32'h8220000;
      24040: inst = 32'h10408000;
      24041: inst = 32'hc4044fd;
      24042: inst = 32'h8220000;
      24043: inst = 32'h10408000;
      24044: inst = 32'hc4044fe;
      24045: inst = 32'h8220000;
      24046: inst = 32'h10408000;
      24047: inst = 32'hc4044ff;
      24048: inst = 32'h8220000;
      24049: inst = 32'h10408000;
      24050: inst = 32'hc404500;
      24051: inst = 32'h8220000;
      24052: inst = 32'h10408000;
      24053: inst = 32'hc404501;
      24054: inst = 32'h8220000;
      24055: inst = 32'h10408000;
      24056: inst = 32'hc404502;
      24057: inst = 32'h8220000;
      24058: inst = 32'h10408000;
      24059: inst = 32'hc404503;
      24060: inst = 32'h8220000;
      24061: inst = 32'h10408000;
      24062: inst = 32'hc404504;
      24063: inst = 32'h8220000;
      24064: inst = 32'h10408000;
      24065: inst = 32'hc404505;
      24066: inst = 32'h8220000;
      24067: inst = 32'h10408000;
      24068: inst = 32'hc404506;
      24069: inst = 32'h8220000;
      24070: inst = 32'h10408000;
      24071: inst = 32'hc404507;
      24072: inst = 32'h8220000;
      24073: inst = 32'h10408000;
      24074: inst = 32'hc404508;
      24075: inst = 32'h8220000;
      24076: inst = 32'h10408000;
      24077: inst = 32'hc404509;
      24078: inst = 32'h8220000;
      24079: inst = 32'h10408000;
      24080: inst = 32'hc40450a;
      24081: inst = 32'h8220000;
      24082: inst = 32'h10408000;
      24083: inst = 32'hc40450b;
      24084: inst = 32'h8220000;
      24085: inst = 32'h10408000;
      24086: inst = 32'hc40450c;
      24087: inst = 32'h8220000;
      24088: inst = 32'h10408000;
      24089: inst = 32'hc40450d;
      24090: inst = 32'h8220000;
      24091: inst = 32'h10408000;
      24092: inst = 32'hc40450e;
      24093: inst = 32'h8220000;
      24094: inst = 32'h10408000;
      24095: inst = 32'hc40450f;
      24096: inst = 32'h8220000;
      24097: inst = 32'h10408000;
      24098: inst = 32'hc404510;
      24099: inst = 32'h8220000;
      24100: inst = 32'h10408000;
      24101: inst = 32'hc404511;
      24102: inst = 32'h8220000;
      24103: inst = 32'h10408000;
      24104: inst = 32'hc404512;
      24105: inst = 32'h8220000;
      24106: inst = 32'h10408000;
      24107: inst = 32'hc404513;
      24108: inst = 32'h8220000;
      24109: inst = 32'h10408000;
      24110: inst = 32'hc404514;
      24111: inst = 32'h8220000;
      24112: inst = 32'h10408000;
      24113: inst = 32'hc404515;
      24114: inst = 32'h8220000;
      24115: inst = 32'h10408000;
      24116: inst = 32'hc404516;
      24117: inst = 32'h8220000;
      24118: inst = 32'h10408000;
      24119: inst = 32'hc404517;
      24120: inst = 32'h8220000;
      24121: inst = 32'h10408000;
      24122: inst = 32'hc404518;
      24123: inst = 32'h8220000;
      24124: inst = 32'h10408000;
      24125: inst = 32'hc404527;
      24126: inst = 32'h8220000;
      24127: inst = 32'h10408000;
      24128: inst = 32'hc404528;
      24129: inst = 32'h8220000;
      24130: inst = 32'h10408000;
      24131: inst = 32'hc404529;
      24132: inst = 32'h8220000;
      24133: inst = 32'h10408000;
      24134: inst = 32'hc40452a;
      24135: inst = 32'h8220000;
      24136: inst = 32'h10408000;
      24137: inst = 32'hc40452b;
      24138: inst = 32'h8220000;
      24139: inst = 32'h10408000;
      24140: inst = 32'hc40452c;
      24141: inst = 32'h8220000;
      24142: inst = 32'h10408000;
      24143: inst = 32'hc40452d;
      24144: inst = 32'h8220000;
      24145: inst = 32'h10408000;
      24146: inst = 32'hc40452e;
      24147: inst = 32'h8220000;
      24148: inst = 32'h10408000;
      24149: inst = 32'hc40452f;
      24150: inst = 32'h8220000;
      24151: inst = 32'h10408000;
      24152: inst = 32'hc404530;
      24153: inst = 32'h8220000;
      24154: inst = 32'h10408000;
      24155: inst = 32'hc404531;
      24156: inst = 32'h8220000;
      24157: inst = 32'h10408000;
      24158: inst = 32'hc404532;
      24159: inst = 32'h8220000;
      24160: inst = 32'h10408000;
      24161: inst = 32'hc404533;
      24162: inst = 32'h8220000;
      24163: inst = 32'h10408000;
      24164: inst = 32'hc404534;
      24165: inst = 32'h8220000;
      24166: inst = 32'h10408000;
      24167: inst = 32'hc404535;
      24168: inst = 32'h8220000;
      24169: inst = 32'h10408000;
      24170: inst = 32'hc404536;
      24171: inst = 32'h8220000;
      24172: inst = 32'h10408000;
      24173: inst = 32'hc404537;
      24174: inst = 32'h8220000;
      24175: inst = 32'h10408000;
      24176: inst = 32'hc404538;
      24177: inst = 32'h8220000;
      24178: inst = 32'h10408000;
      24179: inst = 32'hc404539;
      24180: inst = 32'h8220000;
      24181: inst = 32'h10408000;
      24182: inst = 32'hc40453a;
      24183: inst = 32'h8220000;
      24184: inst = 32'h10408000;
      24185: inst = 32'hc40453b;
      24186: inst = 32'h8220000;
      24187: inst = 32'h10408000;
      24188: inst = 32'hc40453c;
      24189: inst = 32'h8220000;
      24190: inst = 32'h10408000;
      24191: inst = 32'hc40453d;
      24192: inst = 32'h8220000;
      24193: inst = 32'h10408000;
      24194: inst = 32'hc40453e;
      24195: inst = 32'h8220000;
      24196: inst = 32'h10408000;
      24197: inst = 32'hc40453f;
      24198: inst = 32'h8220000;
      24199: inst = 32'h10408000;
      24200: inst = 32'hc404540;
      24201: inst = 32'h8220000;
      24202: inst = 32'h10408000;
      24203: inst = 32'hc404541;
      24204: inst = 32'h8220000;
      24205: inst = 32'h10408000;
      24206: inst = 32'hc404542;
      24207: inst = 32'h8220000;
      24208: inst = 32'h10408000;
      24209: inst = 32'hc404543;
      24210: inst = 32'h8220000;
      24211: inst = 32'h10408000;
      24212: inst = 32'hc404544;
      24213: inst = 32'h8220000;
      24214: inst = 32'h10408000;
      24215: inst = 32'hc404545;
      24216: inst = 32'h8220000;
      24217: inst = 32'h10408000;
      24218: inst = 32'hc404546;
      24219: inst = 32'h8220000;
      24220: inst = 32'h10408000;
      24221: inst = 32'hc404547;
      24222: inst = 32'h8220000;
      24223: inst = 32'h10408000;
      24224: inst = 32'hc404548;
      24225: inst = 32'h8220000;
      24226: inst = 32'h10408000;
      24227: inst = 32'hc404549;
      24228: inst = 32'h8220000;
      24229: inst = 32'h10408000;
      24230: inst = 32'hc40454a;
      24231: inst = 32'h8220000;
      24232: inst = 32'h10408000;
      24233: inst = 32'hc40454b;
      24234: inst = 32'h8220000;
      24235: inst = 32'h10408000;
      24236: inst = 32'hc40454c;
      24237: inst = 32'h8220000;
      24238: inst = 32'h10408000;
      24239: inst = 32'hc40454d;
      24240: inst = 32'h8220000;
      24241: inst = 32'h10408000;
      24242: inst = 32'hc40454e;
      24243: inst = 32'h8220000;
      24244: inst = 32'h10408000;
      24245: inst = 32'hc40454f;
      24246: inst = 32'h8220000;
      24247: inst = 32'h10408000;
      24248: inst = 32'hc404550;
      24249: inst = 32'h8220000;
      24250: inst = 32'h10408000;
      24251: inst = 32'hc404551;
      24252: inst = 32'h8220000;
      24253: inst = 32'h10408000;
      24254: inst = 32'hc404552;
      24255: inst = 32'h8220000;
      24256: inst = 32'h10408000;
      24257: inst = 32'hc404553;
      24258: inst = 32'h8220000;
      24259: inst = 32'h10408000;
      24260: inst = 32'hc404554;
      24261: inst = 32'h8220000;
      24262: inst = 32'h10408000;
      24263: inst = 32'hc404555;
      24264: inst = 32'h8220000;
      24265: inst = 32'h10408000;
      24266: inst = 32'hc404556;
      24267: inst = 32'h8220000;
      24268: inst = 32'h10408000;
      24269: inst = 32'hc404557;
      24270: inst = 32'h8220000;
      24271: inst = 32'h10408000;
      24272: inst = 32'hc404558;
      24273: inst = 32'h8220000;
      24274: inst = 32'h10408000;
      24275: inst = 32'hc404559;
      24276: inst = 32'h8220000;
      24277: inst = 32'h10408000;
      24278: inst = 32'hc40455a;
      24279: inst = 32'h8220000;
      24280: inst = 32'h10408000;
      24281: inst = 32'hc40455b;
      24282: inst = 32'h8220000;
      24283: inst = 32'h10408000;
      24284: inst = 32'hc40455c;
      24285: inst = 32'h8220000;
      24286: inst = 32'h10408000;
      24287: inst = 32'hc40455d;
      24288: inst = 32'h8220000;
      24289: inst = 32'h10408000;
      24290: inst = 32'hc40455e;
      24291: inst = 32'h8220000;
      24292: inst = 32'h10408000;
      24293: inst = 32'hc40455f;
      24294: inst = 32'h8220000;
      24295: inst = 32'h10408000;
      24296: inst = 32'hc404560;
      24297: inst = 32'h8220000;
      24298: inst = 32'h10408000;
      24299: inst = 32'hc404561;
      24300: inst = 32'h8220000;
      24301: inst = 32'h10408000;
      24302: inst = 32'hc404562;
      24303: inst = 32'h8220000;
      24304: inst = 32'h10408000;
      24305: inst = 32'hc404563;
      24306: inst = 32'h8220000;
      24307: inst = 32'h10408000;
      24308: inst = 32'hc404564;
      24309: inst = 32'h8220000;
      24310: inst = 32'h10408000;
      24311: inst = 32'hc404565;
      24312: inst = 32'h8220000;
      24313: inst = 32'h10408000;
      24314: inst = 32'hc404566;
      24315: inst = 32'h8220000;
      24316: inst = 32'h10408000;
      24317: inst = 32'hc404567;
      24318: inst = 32'h8220000;
      24319: inst = 32'h10408000;
      24320: inst = 32'hc404568;
      24321: inst = 32'h8220000;
      24322: inst = 32'h10408000;
      24323: inst = 32'hc404569;
      24324: inst = 32'h8220000;
      24325: inst = 32'h10408000;
      24326: inst = 32'hc40456a;
      24327: inst = 32'h8220000;
      24328: inst = 32'h10408000;
      24329: inst = 32'hc40456b;
      24330: inst = 32'h8220000;
      24331: inst = 32'h10408000;
      24332: inst = 32'hc40456c;
      24333: inst = 32'h8220000;
      24334: inst = 32'h10408000;
      24335: inst = 32'hc40456d;
      24336: inst = 32'h8220000;
      24337: inst = 32'h10408000;
      24338: inst = 32'hc40456e;
      24339: inst = 32'h8220000;
      24340: inst = 32'h10408000;
      24341: inst = 32'hc40456f;
      24342: inst = 32'h8220000;
      24343: inst = 32'h10408000;
      24344: inst = 32'hc404570;
      24345: inst = 32'h8220000;
      24346: inst = 32'h10408000;
      24347: inst = 32'hc404571;
      24348: inst = 32'h8220000;
      24349: inst = 32'h10408000;
      24350: inst = 32'hc404572;
      24351: inst = 32'h8220000;
      24352: inst = 32'h10408000;
      24353: inst = 32'hc404573;
      24354: inst = 32'h8220000;
      24355: inst = 32'h10408000;
      24356: inst = 32'hc404574;
      24357: inst = 32'h8220000;
      24358: inst = 32'h10408000;
      24359: inst = 32'hc404575;
      24360: inst = 32'h8220000;
      24361: inst = 32'h10408000;
      24362: inst = 32'hc404576;
      24363: inst = 32'h8220000;
      24364: inst = 32'h10408000;
      24365: inst = 32'hc404577;
      24366: inst = 32'h8220000;
      24367: inst = 32'h10408000;
      24368: inst = 32'hc404578;
      24369: inst = 32'h8220000;
      24370: inst = 32'h10408000;
      24371: inst = 32'hc404587;
      24372: inst = 32'h8220000;
      24373: inst = 32'h10408000;
      24374: inst = 32'hc404588;
      24375: inst = 32'h8220000;
      24376: inst = 32'h10408000;
      24377: inst = 32'hc404589;
      24378: inst = 32'h8220000;
      24379: inst = 32'h10408000;
      24380: inst = 32'hc40458a;
      24381: inst = 32'h8220000;
      24382: inst = 32'h10408000;
      24383: inst = 32'hc40458b;
      24384: inst = 32'h8220000;
      24385: inst = 32'h10408000;
      24386: inst = 32'hc40458c;
      24387: inst = 32'h8220000;
      24388: inst = 32'h10408000;
      24389: inst = 32'hc40458d;
      24390: inst = 32'h8220000;
      24391: inst = 32'h10408000;
      24392: inst = 32'hc40458e;
      24393: inst = 32'h8220000;
      24394: inst = 32'h10408000;
      24395: inst = 32'hc40458f;
      24396: inst = 32'h8220000;
      24397: inst = 32'h10408000;
      24398: inst = 32'hc404590;
      24399: inst = 32'h8220000;
      24400: inst = 32'h10408000;
      24401: inst = 32'hc404591;
      24402: inst = 32'h8220000;
      24403: inst = 32'h10408000;
      24404: inst = 32'hc404592;
      24405: inst = 32'h8220000;
      24406: inst = 32'h10408000;
      24407: inst = 32'hc404593;
      24408: inst = 32'h8220000;
      24409: inst = 32'h10408000;
      24410: inst = 32'hc404594;
      24411: inst = 32'h8220000;
      24412: inst = 32'h10408000;
      24413: inst = 32'hc404595;
      24414: inst = 32'h8220000;
      24415: inst = 32'h10408000;
      24416: inst = 32'hc404596;
      24417: inst = 32'h8220000;
      24418: inst = 32'h10408000;
      24419: inst = 32'hc404597;
      24420: inst = 32'h8220000;
      24421: inst = 32'h10408000;
      24422: inst = 32'hc404598;
      24423: inst = 32'h8220000;
      24424: inst = 32'h10408000;
      24425: inst = 32'hc404599;
      24426: inst = 32'h8220000;
      24427: inst = 32'h10408000;
      24428: inst = 32'hc40459a;
      24429: inst = 32'h8220000;
      24430: inst = 32'h10408000;
      24431: inst = 32'hc40459b;
      24432: inst = 32'h8220000;
      24433: inst = 32'h10408000;
      24434: inst = 32'hc40459c;
      24435: inst = 32'h8220000;
      24436: inst = 32'h10408000;
      24437: inst = 32'hc40459d;
      24438: inst = 32'h8220000;
      24439: inst = 32'h10408000;
      24440: inst = 32'hc40459e;
      24441: inst = 32'h8220000;
      24442: inst = 32'h10408000;
      24443: inst = 32'hc40459f;
      24444: inst = 32'h8220000;
      24445: inst = 32'h10408000;
      24446: inst = 32'hc4045a0;
      24447: inst = 32'h8220000;
      24448: inst = 32'h10408000;
      24449: inst = 32'hc4045a1;
      24450: inst = 32'h8220000;
      24451: inst = 32'h10408000;
      24452: inst = 32'hc4045a2;
      24453: inst = 32'h8220000;
      24454: inst = 32'h10408000;
      24455: inst = 32'hc4045a3;
      24456: inst = 32'h8220000;
      24457: inst = 32'h10408000;
      24458: inst = 32'hc4045a4;
      24459: inst = 32'h8220000;
      24460: inst = 32'h10408000;
      24461: inst = 32'hc4045a5;
      24462: inst = 32'h8220000;
      24463: inst = 32'h10408000;
      24464: inst = 32'hc4045a6;
      24465: inst = 32'h8220000;
      24466: inst = 32'h10408000;
      24467: inst = 32'hc4045a7;
      24468: inst = 32'h8220000;
      24469: inst = 32'h10408000;
      24470: inst = 32'hc4045a8;
      24471: inst = 32'h8220000;
      24472: inst = 32'h10408000;
      24473: inst = 32'hc4045a9;
      24474: inst = 32'h8220000;
      24475: inst = 32'h10408000;
      24476: inst = 32'hc4045aa;
      24477: inst = 32'h8220000;
      24478: inst = 32'h10408000;
      24479: inst = 32'hc4045ab;
      24480: inst = 32'h8220000;
      24481: inst = 32'h10408000;
      24482: inst = 32'hc4045ac;
      24483: inst = 32'h8220000;
      24484: inst = 32'h10408000;
      24485: inst = 32'hc4045ad;
      24486: inst = 32'h8220000;
      24487: inst = 32'h10408000;
      24488: inst = 32'hc4045ae;
      24489: inst = 32'h8220000;
      24490: inst = 32'h10408000;
      24491: inst = 32'hc4045af;
      24492: inst = 32'h8220000;
      24493: inst = 32'h10408000;
      24494: inst = 32'hc4045b0;
      24495: inst = 32'h8220000;
      24496: inst = 32'h10408000;
      24497: inst = 32'hc4045b1;
      24498: inst = 32'h8220000;
      24499: inst = 32'h10408000;
      24500: inst = 32'hc4045b2;
      24501: inst = 32'h8220000;
      24502: inst = 32'h10408000;
      24503: inst = 32'hc4045b3;
      24504: inst = 32'h8220000;
      24505: inst = 32'h10408000;
      24506: inst = 32'hc4045b4;
      24507: inst = 32'h8220000;
      24508: inst = 32'h10408000;
      24509: inst = 32'hc4045b5;
      24510: inst = 32'h8220000;
      24511: inst = 32'h10408000;
      24512: inst = 32'hc4045b6;
      24513: inst = 32'h8220000;
      24514: inst = 32'h10408000;
      24515: inst = 32'hc4045b7;
      24516: inst = 32'h8220000;
      24517: inst = 32'h10408000;
      24518: inst = 32'hc4045b8;
      24519: inst = 32'h8220000;
      24520: inst = 32'h10408000;
      24521: inst = 32'hc4045b9;
      24522: inst = 32'h8220000;
      24523: inst = 32'h10408000;
      24524: inst = 32'hc4045ba;
      24525: inst = 32'h8220000;
      24526: inst = 32'h10408000;
      24527: inst = 32'hc4045bb;
      24528: inst = 32'h8220000;
      24529: inst = 32'h10408000;
      24530: inst = 32'hc4045bc;
      24531: inst = 32'h8220000;
      24532: inst = 32'h10408000;
      24533: inst = 32'hc4045bd;
      24534: inst = 32'h8220000;
      24535: inst = 32'h10408000;
      24536: inst = 32'hc4045be;
      24537: inst = 32'h8220000;
      24538: inst = 32'h10408000;
      24539: inst = 32'hc4045bf;
      24540: inst = 32'h8220000;
      24541: inst = 32'h10408000;
      24542: inst = 32'hc4045c0;
      24543: inst = 32'h8220000;
      24544: inst = 32'h10408000;
      24545: inst = 32'hc4045c1;
      24546: inst = 32'h8220000;
      24547: inst = 32'h10408000;
      24548: inst = 32'hc4045c2;
      24549: inst = 32'h8220000;
      24550: inst = 32'h10408000;
      24551: inst = 32'hc4045c3;
      24552: inst = 32'h8220000;
      24553: inst = 32'h10408000;
      24554: inst = 32'hc4045c4;
      24555: inst = 32'h8220000;
      24556: inst = 32'h10408000;
      24557: inst = 32'hc4045c5;
      24558: inst = 32'h8220000;
      24559: inst = 32'h10408000;
      24560: inst = 32'hc4045c6;
      24561: inst = 32'h8220000;
      24562: inst = 32'h10408000;
      24563: inst = 32'hc4045c7;
      24564: inst = 32'h8220000;
      24565: inst = 32'h10408000;
      24566: inst = 32'hc4045c8;
      24567: inst = 32'h8220000;
      24568: inst = 32'h10408000;
      24569: inst = 32'hc4045c9;
      24570: inst = 32'h8220000;
      24571: inst = 32'h10408000;
      24572: inst = 32'hc4045ca;
      24573: inst = 32'h8220000;
      24574: inst = 32'h10408000;
      24575: inst = 32'hc4045cb;
      24576: inst = 32'h8220000;
      24577: inst = 32'h10408000;
      24578: inst = 32'hc4045cc;
      24579: inst = 32'h8220000;
      24580: inst = 32'h10408000;
      24581: inst = 32'hc4045cd;
      24582: inst = 32'h8220000;
      24583: inst = 32'h10408000;
      24584: inst = 32'hc4045ce;
      24585: inst = 32'h8220000;
      24586: inst = 32'h10408000;
      24587: inst = 32'hc4045cf;
      24588: inst = 32'h8220000;
      24589: inst = 32'h10408000;
      24590: inst = 32'hc4045d0;
      24591: inst = 32'h8220000;
      24592: inst = 32'h10408000;
      24593: inst = 32'hc4045d1;
      24594: inst = 32'h8220000;
      24595: inst = 32'h10408000;
      24596: inst = 32'hc4045d2;
      24597: inst = 32'h8220000;
      24598: inst = 32'h10408000;
      24599: inst = 32'hc4045d3;
      24600: inst = 32'h8220000;
      24601: inst = 32'h10408000;
      24602: inst = 32'hc4045d4;
      24603: inst = 32'h8220000;
      24604: inst = 32'h10408000;
      24605: inst = 32'hc4045d5;
      24606: inst = 32'h8220000;
      24607: inst = 32'h10408000;
      24608: inst = 32'hc4045d6;
      24609: inst = 32'h8220000;
      24610: inst = 32'h10408000;
      24611: inst = 32'hc4045d7;
      24612: inst = 32'h8220000;
      24613: inst = 32'h10408000;
      24614: inst = 32'hc4045d8;
      24615: inst = 32'h8220000;
      24616: inst = 32'h10408000;
      24617: inst = 32'hc4045e7;
      24618: inst = 32'h8220000;
      24619: inst = 32'h10408000;
      24620: inst = 32'hc4045e8;
      24621: inst = 32'h8220000;
      24622: inst = 32'h10408000;
      24623: inst = 32'hc4045e9;
      24624: inst = 32'h8220000;
      24625: inst = 32'h10408000;
      24626: inst = 32'hc4045ea;
      24627: inst = 32'h8220000;
      24628: inst = 32'h10408000;
      24629: inst = 32'hc4045eb;
      24630: inst = 32'h8220000;
      24631: inst = 32'h10408000;
      24632: inst = 32'hc4045ec;
      24633: inst = 32'h8220000;
      24634: inst = 32'h10408000;
      24635: inst = 32'hc4045ed;
      24636: inst = 32'h8220000;
      24637: inst = 32'h10408000;
      24638: inst = 32'hc4045ee;
      24639: inst = 32'h8220000;
      24640: inst = 32'h10408000;
      24641: inst = 32'hc4045ef;
      24642: inst = 32'h8220000;
      24643: inst = 32'h10408000;
      24644: inst = 32'hc4045f0;
      24645: inst = 32'h8220000;
      24646: inst = 32'h10408000;
      24647: inst = 32'hc4045f1;
      24648: inst = 32'h8220000;
      24649: inst = 32'h10408000;
      24650: inst = 32'hc4045f2;
      24651: inst = 32'h8220000;
      24652: inst = 32'h10408000;
      24653: inst = 32'hc4045f3;
      24654: inst = 32'h8220000;
      24655: inst = 32'h10408000;
      24656: inst = 32'hc4045f4;
      24657: inst = 32'h8220000;
      24658: inst = 32'h10408000;
      24659: inst = 32'hc4045f5;
      24660: inst = 32'h8220000;
      24661: inst = 32'h10408000;
      24662: inst = 32'hc4045f6;
      24663: inst = 32'h8220000;
      24664: inst = 32'h10408000;
      24665: inst = 32'hc4045f7;
      24666: inst = 32'h8220000;
      24667: inst = 32'h10408000;
      24668: inst = 32'hc4045f8;
      24669: inst = 32'h8220000;
      24670: inst = 32'h10408000;
      24671: inst = 32'hc4045f9;
      24672: inst = 32'h8220000;
      24673: inst = 32'h10408000;
      24674: inst = 32'hc4045fa;
      24675: inst = 32'h8220000;
      24676: inst = 32'h10408000;
      24677: inst = 32'hc4045fb;
      24678: inst = 32'h8220000;
      24679: inst = 32'h10408000;
      24680: inst = 32'hc4045fc;
      24681: inst = 32'h8220000;
      24682: inst = 32'h10408000;
      24683: inst = 32'hc4045fd;
      24684: inst = 32'h8220000;
      24685: inst = 32'h10408000;
      24686: inst = 32'hc4045fe;
      24687: inst = 32'h8220000;
      24688: inst = 32'h10408000;
      24689: inst = 32'hc4045ff;
      24690: inst = 32'h8220000;
      24691: inst = 32'h10408000;
      24692: inst = 32'hc404600;
      24693: inst = 32'h8220000;
      24694: inst = 32'h10408000;
      24695: inst = 32'hc404601;
      24696: inst = 32'h8220000;
      24697: inst = 32'h10408000;
      24698: inst = 32'hc404602;
      24699: inst = 32'h8220000;
      24700: inst = 32'h10408000;
      24701: inst = 32'hc404603;
      24702: inst = 32'h8220000;
      24703: inst = 32'h10408000;
      24704: inst = 32'hc404604;
      24705: inst = 32'h8220000;
      24706: inst = 32'h10408000;
      24707: inst = 32'hc404605;
      24708: inst = 32'h8220000;
      24709: inst = 32'h10408000;
      24710: inst = 32'hc404606;
      24711: inst = 32'h8220000;
      24712: inst = 32'h10408000;
      24713: inst = 32'hc404607;
      24714: inst = 32'h8220000;
      24715: inst = 32'h10408000;
      24716: inst = 32'hc404608;
      24717: inst = 32'h8220000;
      24718: inst = 32'h10408000;
      24719: inst = 32'hc404609;
      24720: inst = 32'h8220000;
      24721: inst = 32'h10408000;
      24722: inst = 32'hc40460a;
      24723: inst = 32'h8220000;
      24724: inst = 32'h10408000;
      24725: inst = 32'hc40460b;
      24726: inst = 32'h8220000;
      24727: inst = 32'h10408000;
      24728: inst = 32'hc40460c;
      24729: inst = 32'h8220000;
      24730: inst = 32'h10408000;
      24731: inst = 32'hc40460d;
      24732: inst = 32'h8220000;
      24733: inst = 32'h10408000;
      24734: inst = 32'hc40460e;
      24735: inst = 32'h8220000;
      24736: inst = 32'h10408000;
      24737: inst = 32'hc40460f;
      24738: inst = 32'h8220000;
      24739: inst = 32'h10408000;
      24740: inst = 32'hc404610;
      24741: inst = 32'h8220000;
      24742: inst = 32'h10408000;
      24743: inst = 32'hc404611;
      24744: inst = 32'h8220000;
      24745: inst = 32'h10408000;
      24746: inst = 32'hc404612;
      24747: inst = 32'h8220000;
      24748: inst = 32'h10408000;
      24749: inst = 32'hc404613;
      24750: inst = 32'h8220000;
      24751: inst = 32'h10408000;
      24752: inst = 32'hc404614;
      24753: inst = 32'h8220000;
      24754: inst = 32'h10408000;
      24755: inst = 32'hc404615;
      24756: inst = 32'h8220000;
      24757: inst = 32'h10408000;
      24758: inst = 32'hc404616;
      24759: inst = 32'h8220000;
      24760: inst = 32'h10408000;
      24761: inst = 32'hc404617;
      24762: inst = 32'h8220000;
      24763: inst = 32'h10408000;
      24764: inst = 32'hc404618;
      24765: inst = 32'h8220000;
      24766: inst = 32'h10408000;
      24767: inst = 32'hc404619;
      24768: inst = 32'h8220000;
      24769: inst = 32'h10408000;
      24770: inst = 32'hc40461a;
      24771: inst = 32'h8220000;
      24772: inst = 32'h10408000;
      24773: inst = 32'hc40461b;
      24774: inst = 32'h8220000;
      24775: inst = 32'h10408000;
      24776: inst = 32'hc40461c;
      24777: inst = 32'h8220000;
      24778: inst = 32'h10408000;
      24779: inst = 32'hc40461d;
      24780: inst = 32'h8220000;
      24781: inst = 32'h10408000;
      24782: inst = 32'hc40461e;
      24783: inst = 32'h8220000;
      24784: inst = 32'h10408000;
      24785: inst = 32'hc40461f;
      24786: inst = 32'h8220000;
      24787: inst = 32'h10408000;
      24788: inst = 32'hc404620;
      24789: inst = 32'h8220000;
      24790: inst = 32'h10408000;
      24791: inst = 32'hc404621;
      24792: inst = 32'h8220000;
      24793: inst = 32'h10408000;
      24794: inst = 32'hc404622;
      24795: inst = 32'h8220000;
      24796: inst = 32'h10408000;
      24797: inst = 32'hc404623;
      24798: inst = 32'h8220000;
      24799: inst = 32'h10408000;
      24800: inst = 32'hc404624;
      24801: inst = 32'h8220000;
      24802: inst = 32'h10408000;
      24803: inst = 32'hc404625;
      24804: inst = 32'h8220000;
      24805: inst = 32'h10408000;
      24806: inst = 32'hc404626;
      24807: inst = 32'h8220000;
      24808: inst = 32'h10408000;
      24809: inst = 32'hc404627;
      24810: inst = 32'h8220000;
      24811: inst = 32'h10408000;
      24812: inst = 32'hc404628;
      24813: inst = 32'h8220000;
      24814: inst = 32'h10408000;
      24815: inst = 32'hc404629;
      24816: inst = 32'h8220000;
      24817: inst = 32'h10408000;
      24818: inst = 32'hc40462a;
      24819: inst = 32'h8220000;
      24820: inst = 32'h10408000;
      24821: inst = 32'hc40462b;
      24822: inst = 32'h8220000;
      24823: inst = 32'h10408000;
      24824: inst = 32'hc40462c;
      24825: inst = 32'h8220000;
      24826: inst = 32'h10408000;
      24827: inst = 32'hc40462d;
      24828: inst = 32'h8220000;
      24829: inst = 32'h10408000;
      24830: inst = 32'hc40462e;
      24831: inst = 32'h8220000;
      24832: inst = 32'h10408000;
      24833: inst = 32'hc40462f;
      24834: inst = 32'h8220000;
      24835: inst = 32'h10408000;
      24836: inst = 32'hc404630;
      24837: inst = 32'h8220000;
      24838: inst = 32'h10408000;
      24839: inst = 32'hc404631;
      24840: inst = 32'h8220000;
      24841: inst = 32'h10408000;
      24842: inst = 32'hc404632;
      24843: inst = 32'h8220000;
      24844: inst = 32'h10408000;
      24845: inst = 32'hc404633;
      24846: inst = 32'h8220000;
      24847: inst = 32'h10408000;
      24848: inst = 32'hc404634;
      24849: inst = 32'h8220000;
      24850: inst = 32'h10408000;
      24851: inst = 32'hc404635;
      24852: inst = 32'h8220000;
      24853: inst = 32'h10408000;
      24854: inst = 32'hc404636;
      24855: inst = 32'h8220000;
      24856: inst = 32'h10408000;
      24857: inst = 32'hc404637;
      24858: inst = 32'h8220000;
      24859: inst = 32'h10408000;
      24860: inst = 32'hc404638;
      24861: inst = 32'h8220000;
      24862: inst = 32'h10408000;
      24863: inst = 32'hc404647;
      24864: inst = 32'h8220000;
      24865: inst = 32'h10408000;
      24866: inst = 32'hc404648;
      24867: inst = 32'h8220000;
      24868: inst = 32'h10408000;
      24869: inst = 32'hc404649;
      24870: inst = 32'h8220000;
      24871: inst = 32'h10408000;
      24872: inst = 32'hc40464a;
      24873: inst = 32'h8220000;
      24874: inst = 32'h10408000;
      24875: inst = 32'hc40464b;
      24876: inst = 32'h8220000;
      24877: inst = 32'h10408000;
      24878: inst = 32'hc40464c;
      24879: inst = 32'h8220000;
      24880: inst = 32'h10408000;
      24881: inst = 32'hc40464d;
      24882: inst = 32'h8220000;
      24883: inst = 32'h10408000;
      24884: inst = 32'hc404651;
      24885: inst = 32'h8220000;
      24886: inst = 32'h10408000;
      24887: inst = 32'hc404652;
      24888: inst = 32'h8220000;
      24889: inst = 32'h10408000;
      24890: inst = 32'hc404653;
      24891: inst = 32'h8220000;
      24892: inst = 32'h10408000;
      24893: inst = 32'hc404654;
      24894: inst = 32'h8220000;
      24895: inst = 32'h10408000;
      24896: inst = 32'hc404655;
      24897: inst = 32'h8220000;
      24898: inst = 32'h10408000;
      24899: inst = 32'hc404656;
      24900: inst = 32'h8220000;
      24901: inst = 32'h10408000;
      24902: inst = 32'hc404657;
      24903: inst = 32'h8220000;
      24904: inst = 32'h10408000;
      24905: inst = 32'hc404658;
      24906: inst = 32'h8220000;
      24907: inst = 32'h10408000;
      24908: inst = 32'hc404659;
      24909: inst = 32'h8220000;
      24910: inst = 32'h10408000;
      24911: inst = 32'hc40465a;
      24912: inst = 32'h8220000;
      24913: inst = 32'h10408000;
      24914: inst = 32'hc40465b;
      24915: inst = 32'h8220000;
      24916: inst = 32'h10408000;
      24917: inst = 32'hc40465c;
      24918: inst = 32'h8220000;
      24919: inst = 32'h10408000;
      24920: inst = 32'hc40465d;
      24921: inst = 32'h8220000;
      24922: inst = 32'h10408000;
      24923: inst = 32'hc40465e;
      24924: inst = 32'h8220000;
      24925: inst = 32'h10408000;
      24926: inst = 32'hc40465f;
      24927: inst = 32'h8220000;
      24928: inst = 32'h10408000;
      24929: inst = 32'hc404660;
      24930: inst = 32'h8220000;
      24931: inst = 32'h10408000;
      24932: inst = 32'hc404661;
      24933: inst = 32'h8220000;
      24934: inst = 32'h10408000;
      24935: inst = 32'hc404662;
      24936: inst = 32'h8220000;
      24937: inst = 32'h10408000;
      24938: inst = 32'hc404663;
      24939: inst = 32'h8220000;
      24940: inst = 32'h10408000;
      24941: inst = 32'hc404664;
      24942: inst = 32'h8220000;
      24943: inst = 32'h10408000;
      24944: inst = 32'hc404665;
      24945: inst = 32'h8220000;
      24946: inst = 32'h10408000;
      24947: inst = 32'hc404666;
      24948: inst = 32'h8220000;
      24949: inst = 32'h10408000;
      24950: inst = 32'hc404667;
      24951: inst = 32'h8220000;
      24952: inst = 32'h10408000;
      24953: inst = 32'hc404668;
      24954: inst = 32'h8220000;
      24955: inst = 32'h10408000;
      24956: inst = 32'hc404669;
      24957: inst = 32'h8220000;
      24958: inst = 32'h10408000;
      24959: inst = 32'hc40466a;
      24960: inst = 32'h8220000;
      24961: inst = 32'h10408000;
      24962: inst = 32'hc40466b;
      24963: inst = 32'h8220000;
      24964: inst = 32'h10408000;
      24965: inst = 32'hc40466c;
      24966: inst = 32'h8220000;
      24967: inst = 32'h10408000;
      24968: inst = 32'hc40466d;
      24969: inst = 32'h8220000;
      24970: inst = 32'h10408000;
      24971: inst = 32'hc40466e;
      24972: inst = 32'h8220000;
      24973: inst = 32'h10408000;
      24974: inst = 32'hc40466f;
      24975: inst = 32'h8220000;
      24976: inst = 32'h10408000;
      24977: inst = 32'hc404670;
      24978: inst = 32'h8220000;
      24979: inst = 32'h10408000;
      24980: inst = 32'hc404671;
      24981: inst = 32'h8220000;
      24982: inst = 32'h10408000;
      24983: inst = 32'hc404672;
      24984: inst = 32'h8220000;
      24985: inst = 32'h10408000;
      24986: inst = 32'hc404673;
      24987: inst = 32'h8220000;
      24988: inst = 32'h10408000;
      24989: inst = 32'hc404674;
      24990: inst = 32'h8220000;
      24991: inst = 32'h10408000;
      24992: inst = 32'hc404675;
      24993: inst = 32'h8220000;
      24994: inst = 32'h10408000;
      24995: inst = 32'hc404676;
      24996: inst = 32'h8220000;
      24997: inst = 32'h10408000;
      24998: inst = 32'hc404677;
      24999: inst = 32'h8220000;
      25000: inst = 32'h10408000;
      25001: inst = 32'hc404678;
      25002: inst = 32'h8220000;
      25003: inst = 32'h10408000;
      25004: inst = 32'hc404679;
      25005: inst = 32'h8220000;
      25006: inst = 32'h10408000;
      25007: inst = 32'hc40467a;
      25008: inst = 32'h8220000;
      25009: inst = 32'h10408000;
      25010: inst = 32'hc40467b;
      25011: inst = 32'h8220000;
      25012: inst = 32'h10408000;
      25013: inst = 32'hc40467c;
      25014: inst = 32'h8220000;
      25015: inst = 32'h10408000;
      25016: inst = 32'hc40467d;
      25017: inst = 32'h8220000;
      25018: inst = 32'h10408000;
      25019: inst = 32'hc40467e;
      25020: inst = 32'h8220000;
      25021: inst = 32'h10408000;
      25022: inst = 32'hc40467f;
      25023: inst = 32'h8220000;
      25024: inst = 32'h10408000;
      25025: inst = 32'hc404680;
      25026: inst = 32'h8220000;
      25027: inst = 32'h10408000;
      25028: inst = 32'hc404681;
      25029: inst = 32'h8220000;
      25030: inst = 32'h10408000;
      25031: inst = 32'hc404682;
      25032: inst = 32'h8220000;
      25033: inst = 32'h10408000;
      25034: inst = 32'hc404683;
      25035: inst = 32'h8220000;
      25036: inst = 32'h10408000;
      25037: inst = 32'hc404684;
      25038: inst = 32'h8220000;
      25039: inst = 32'h10408000;
      25040: inst = 32'hc404685;
      25041: inst = 32'h8220000;
      25042: inst = 32'h10408000;
      25043: inst = 32'hc404686;
      25044: inst = 32'h8220000;
      25045: inst = 32'h10408000;
      25046: inst = 32'hc404687;
      25047: inst = 32'h8220000;
      25048: inst = 32'h10408000;
      25049: inst = 32'hc404688;
      25050: inst = 32'h8220000;
      25051: inst = 32'h10408000;
      25052: inst = 32'hc404689;
      25053: inst = 32'h8220000;
      25054: inst = 32'h10408000;
      25055: inst = 32'hc40468a;
      25056: inst = 32'h8220000;
      25057: inst = 32'h10408000;
      25058: inst = 32'hc40468b;
      25059: inst = 32'h8220000;
      25060: inst = 32'h10408000;
      25061: inst = 32'hc40468c;
      25062: inst = 32'h8220000;
      25063: inst = 32'h10408000;
      25064: inst = 32'hc40468d;
      25065: inst = 32'h8220000;
      25066: inst = 32'h10408000;
      25067: inst = 32'hc40468e;
      25068: inst = 32'h8220000;
      25069: inst = 32'h10408000;
      25070: inst = 32'hc40468f;
      25071: inst = 32'h8220000;
      25072: inst = 32'h10408000;
      25073: inst = 32'hc404693;
      25074: inst = 32'h8220000;
      25075: inst = 32'h10408000;
      25076: inst = 32'hc404694;
      25077: inst = 32'h8220000;
      25078: inst = 32'h10408000;
      25079: inst = 32'hc404695;
      25080: inst = 32'h8220000;
      25081: inst = 32'h10408000;
      25082: inst = 32'hc404696;
      25083: inst = 32'h8220000;
      25084: inst = 32'h10408000;
      25085: inst = 32'hc404697;
      25086: inst = 32'h8220000;
      25087: inst = 32'h10408000;
      25088: inst = 32'hc404698;
      25089: inst = 32'h8220000;
      25090: inst = 32'h10408000;
      25091: inst = 32'hc4046a7;
      25092: inst = 32'h8220000;
      25093: inst = 32'h10408000;
      25094: inst = 32'hc4046a8;
      25095: inst = 32'h8220000;
      25096: inst = 32'h10408000;
      25097: inst = 32'hc4046a9;
      25098: inst = 32'h8220000;
      25099: inst = 32'h10408000;
      25100: inst = 32'hc4046aa;
      25101: inst = 32'h8220000;
      25102: inst = 32'h10408000;
      25103: inst = 32'hc4046ab;
      25104: inst = 32'h8220000;
      25105: inst = 32'h10408000;
      25106: inst = 32'hc4046ac;
      25107: inst = 32'h8220000;
      25108: inst = 32'h10408000;
      25109: inst = 32'hc4046ad;
      25110: inst = 32'h8220000;
      25111: inst = 32'h10408000;
      25112: inst = 32'hc4046b1;
      25113: inst = 32'h8220000;
      25114: inst = 32'h10408000;
      25115: inst = 32'hc4046b2;
      25116: inst = 32'h8220000;
      25117: inst = 32'h10408000;
      25118: inst = 32'hc4046b3;
      25119: inst = 32'h8220000;
      25120: inst = 32'h10408000;
      25121: inst = 32'hc4046b4;
      25122: inst = 32'h8220000;
      25123: inst = 32'h10408000;
      25124: inst = 32'hc4046b5;
      25125: inst = 32'h8220000;
      25126: inst = 32'h10408000;
      25127: inst = 32'hc4046b6;
      25128: inst = 32'h8220000;
      25129: inst = 32'h10408000;
      25130: inst = 32'hc4046b7;
      25131: inst = 32'h8220000;
      25132: inst = 32'h10408000;
      25133: inst = 32'hc4046b8;
      25134: inst = 32'h8220000;
      25135: inst = 32'h10408000;
      25136: inst = 32'hc4046b9;
      25137: inst = 32'h8220000;
      25138: inst = 32'h10408000;
      25139: inst = 32'hc4046ba;
      25140: inst = 32'h8220000;
      25141: inst = 32'h10408000;
      25142: inst = 32'hc4046bb;
      25143: inst = 32'h8220000;
      25144: inst = 32'h10408000;
      25145: inst = 32'hc4046bc;
      25146: inst = 32'h8220000;
      25147: inst = 32'h10408000;
      25148: inst = 32'hc4046bd;
      25149: inst = 32'h8220000;
      25150: inst = 32'h10408000;
      25151: inst = 32'hc4046be;
      25152: inst = 32'h8220000;
      25153: inst = 32'h10408000;
      25154: inst = 32'hc4046bf;
      25155: inst = 32'h8220000;
      25156: inst = 32'h10408000;
      25157: inst = 32'hc4046c0;
      25158: inst = 32'h8220000;
      25159: inst = 32'h10408000;
      25160: inst = 32'hc4046c1;
      25161: inst = 32'h8220000;
      25162: inst = 32'h10408000;
      25163: inst = 32'hc4046c2;
      25164: inst = 32'h8220000;
      25165: inst = 32'h10408000;
      25166: inst = 32'hc4046c3;
      25167: inst = 32'h8220000;
      25168: inst = 32'h10408000;
      25169: inst = 32'hc4046c4;
      25170: inst = 32'h8220000;
      25171: inst = 32'h10408000;
      25172: inst = 32'hc4046c5;
      25173: inst = 32'h8220000;
      25174: inst = 32'h10408000;
      25175: inst = 32'hc4046c6;
      25176: inst = 32'h8220000;
      25177: inst = 32'h10408000;
      25178: inst = 32'hc4046c7;
      25179: inst = 32'h8220000;
      25180: inst = 32'h10408000;
      25181: inst = 32'hc4046c8;
      25182: inst = 32'h8220000;
      25183: inst = 32'h10408000;
      25184: inst = 32'hc4046c9;
      25185: inst = 32'h8220000;
      25186: inst = 32'h10408000;
      25187: inst = 32'hc4046ca;
      25188: inst = 32'h8220000;
      25189: inst = 32'h10408000;
      25190: inst = 32'hc4046cb;
      25191: inst = 32'h8220000;
      25192: inst = 32'h10408000;
      25193: inst = 32'hc4046cc;
      25194: inst = 32'h8220000;
      25195: inst = 32'h10408000;
      25196: inst = 32'hc4046cd;
      25197: inst = 32'h8220000;
      25198: inst = 32'h10408000;
      25199: inst = 32'hc4046ce;
      25200: inst = 32'h8220000;
      25201: inst = 32'h10408000;
      25202: inst = 32'hc4046cf;
      25203: inst = 32'h8220000;
      25204: inst = 32'h10408000;
      25205: inst = 32'hc4046d0;
      25206: inst = 32'h8220000;
      25207: inst = 32'h10408000;
      25208: inst = 32'hc4046d1;
      25209: inst = 32'h8220000;
      25210: inst = 32'h10408000;
      25211: inst = 32'hc4046d2;
      25212: inst = 32'h8220000;
      25213: inst = 32'h10408000;
      25214: inst = 32'hc4046d3;
      25215: inst = 32'h8220000;
      25216: inst = 32'h10408000;
      25217: inst = 32'hc4046d4;
      25218: inst = 32'h8220000;
      25219: inst = 32'h10408000;
      25220: inst = 32'hc4046d5;
      25221: inst = 32'h8220000;
      25222: inst = 32'h10408000;
      25223: inst = 32'hc4046d6;
      25224: inst = 32'h8220000;
      25225: inst = 32'h10408000;
      25226: inst = 32'hc4046d7;
      25227: inst = 32'h8220000;
      25228: inst = 32'h10408000;
      25229: inst = 32'hc4046d8;
      25230: inst = 32'h8220000;
      25231: inst = 32'h10408000;
      25232: inst = 32'hc4046d9;
      25233: inst = 32'h8220000;
      25234: inst = 32'h10408000;
      25235: inst = 32'hc4046da;
      25236: inst = 32'h8220000;
      25237: inst = 32'h10408000;
      25238: inst = 32'hc4046db;
      25239: inst = 32'h8220000;
      25240: inst = 32'h10408000;
      25241: inst = 32'hc4046dc;
      25242: inst = 32'h8220000;
      25243: inst = 32'h10408000;
      25244: inst = 32'hc4046dd;
      25245: inst = 32'h8220000;
      25246: inst = 32'h10408000;
      25247: inst = 32'hc4046de;
      25248: inst = 32'h8220000;
      25249: inst = 32'h10408000;
      25250: inst = 32'hc4046df;
      25251: inst = 32'h8220000;
      25252: inst = 32'h10408000;
      25253: inst = 32'hc4046e0;
      25254: inst = 32'h8220000;
      25255: inst = 32'h10408000;
      25256: inst = 32'hc4046e1;
      25257: inst = 32'h8220000;
      25258: inst = 32'h10408000;
      25259: inst = 32'hc4046e2;
      25260: inst = 32'h8220000;
      25261: inst = 32'h10408000;
      25262: inst = 32'hc4046e3;
      25263: inst = 32'h8220000;
      25264: inst = 32'h10408000;
      25265: inst = 32'hc4046e4;
      25266: inst = 32'h8220000;
      25267: inst = 32'h10408000;
      25268: inst = 32'hc4046e5;
      25269: inst = 32'h8220000;
      25270: inst = 32'h10408000;
      25271: inst = 32'hc4046e6;
      25272: inst = 32'h8220000;
      25273: inst = 32'h10408000;
      25274: inst = 32'hc4046e7;
      25275: inst = 32'h8220000;
      25276: inst = 32'h10408000;
      25277: inst = 32'hc4046e8;
      25278: inst = 32'h8220000;
      25279: inst = 32'h10408000;
      25280: inst = 32'hc4046e9;
      25281: inst = 32'h8220000;
      25282: inst = 32'h10408000;
      25283: inst = 32'hc4046ea;
      25284: inst = 32'h8220000;
      25285: inst = 32'h10408000;
      25286: inst = 32'hc4046eb;
      25287: inst = 32'h8220000;
      25288: inst = 32'h10408000;
      25289: inst = 32'hc4046ec;
      25290: inst = 32'h8220000;
      25291: inst = 32'h10408000;
      25292: inst = 32'hc4046ed;
      25293: inst = 32'h8220000;
      25294: inst = 32'h10408000;
      25295: inst = 32'hc4046ee;
      25296: inst = 32'h8220000;
      25297: inst = 32'h10408000;
      25298: inst = 32'hc4046ef;
      25299: inst = 32'h8220000;
      25300: inst = 32'h10408000;
      25301: inst = 32'hc4046f3;
      25302: inst = 32'h8220000;
      25303: inst = 32'h10408000;
      25304: inst = 32'hc4046f4;
      25305: inst = 32'h8220000;
      25306: inst = 32'h10408000;
      25307: inst = 32'hc4046f5;
      25308: inst = 32'h8220000;
      25309: inst = 32'h10408000;
      25310: inst = 32'hc4046f6;
      25311: inst = 32'h8220000;
      25312: inst = 32'h10408000;
      25313: inst = 32'hc4046f7;
      25314: inst = 32'h8220000;
      25315: inst = 32'h10408000;
      25316: inst = 32'hc4046f8;
      25317: inst = 32'h8220000;
      25318: inst = 32'h10408000;
      25319: inst = 32'hc404707;
      25320: inst = 32'h8220000;
      25321: inst = 32'h10408000;
      25322: inst = 32'hc404708;
      25323: inst = 32'h8220000;
      25324: inst = 32'h10408000;
      25325: inst = 32'hc404709;
      25326: inst = 32'h8220000;
      25327: inst = 32'h10408000;
      25328: inst = 32'hc40470a;
      25329: inst = 32'h8220000;
      25330: inst = 32'h10408000;
      25331: inst = 32'hc40470b;
      25332: inst = 32'h8220000;
      25333: inst = 32'h10408000;
      25334: inst = 32'hc40470c;
      25335: inst = 32'h8220000;
      25336: inst = 32'h10408000;
      25337: inst = 32'hc40470d;
      25338: inst = 32'h8220000;
      25339: inst = 32'h10408000;
      25340: inst = 32'hc40470e;
      25341: inst = 32'h8220000;
      25342: inst = 32'h10408000;
      25343: inst = 32'hc404711;
      25344: inst = 32'h8220000;
      25345: inst = 32'h10408000;
      25346: inst = 32'hc404712;
      25347: inst = 32'h8220000;
      25348: inst = 32'h10408000;
      25349: inst = 32'hc404713;
      25350: inst = 32'h8220000;
      25351: inst = 32'h10408000;
      25352: inst = 32'hc404714;
      25353: inst = 32'h8220000;
      25354: inst = 32'h10408000;
      25355: inst = 32'hc404717;
      25356: inst = 32'h8220000;
      25357: inst = 32'h10408000;
      25358: inst = 32'hc404718;
      25359: inst = 32'h8220000;
      25360: inst = 32'h10408000;
      25361: inst = 32'hc404719;
      25362: inst = 32'h8220000;
      25363: inst = 32'h10408000;
      25364: inst = 32'hc40471a;
      25365: inst = 32'h8220000;
      25366: inst = 32'h10408000;
      25367: inst = 32'hc40471b;
      25368: inst = 32'h8220000;
      25369: inst = 32'h10408000;
      25370: inst = 32'hc40471c;
      25371: inst = 32'h8220000;
      25372: inst = 32'h10408000;
      25373: inst = 32'hc40471d;
      25374: inst = 32'h8220000;
      25375: inst = 32'h10408000;
      25376: inst = 32'hc40471e;
      25377: inst = 32'h8220000;
      25378: inst = 32'h10408000;
      25379: inst = 32'hc40471f;
      25380: inst = 32'h8220000;
      25381: inst = 32'h10408000;
      25382: inst = 32'hc404720;
      25383: inst = 32'h8220000;
      25384: inst = 32'h10408000;
      25385: inst = 32'hc404721;
      25386: inst = 32'h8220000;
      25387: inst = 32'h10408000;
      25388: inst = 32'hc404722;
      25389: inst = 32'h8220000;
      25390: inst = 32'h10408000;
      25391: inst = 32'hc404723;
      25392: inst = 32'h8220000;
      25393: inst = 32'h10408000;
      25394: inst = 32'hc404726;
      25395: inst = 32'h8220000;
      25396: inst = 32'h10408000;
      25397: inst = 32'hc404727;
      25398: inst = 32'h8220000;
      25399: inst = 32'h10408000;
      25400: inst = 32'hc404728;
      25401: inst = 32'h8220000;
      25402: inst = 32'h10408000;
      25403: inst = 32'hc404729;
      25404: inst = 32'h8220000;
      25405: inst = 32'h10408000;
      25406: inst = 32'hc40472a;
      25407: inst = 32'h8220000;
      25408: inst = 32'h10408000;
      25409: inst = 32'hc40472b;
      25410: inst = 32'h8220000;
      25411: inst = 32'h10408000;
      25412: inst = 32'hc40472c;
      25413: inst = 32'h8220000;
      25414: inst = 32'h10408000;
      25415: inst = 32'hc40472d;
      25416: inst = 32'h8220000;
      25417: inst = 32'h10408000;
      25418: inst = 32'hc40472e;
      25419: inst = 32'h8220000;
      25420: inst = 32'h10408000;
      25421: inst = 32'hc40472f;
      25422: inst = 32'h8220000;
      25423: inst = 32'h10408000;
      25424: inst = 32'hc404730;
      25425: inst = 32'h8220000;
      25426: inst = 32'h10408000;
      25427: inst = 32'hc404731;
      25428: inst = 32'h8220000;
      25429: inst = 32'h10408000;
      25430: inst = 32'hc404732;
      25431: inst = 32'h8220000;
      25432: inst = 32'h10408000;
      25433: inst = 32'hc404733;
      25434: inst = 32'h8220000;
      25435: inst = 32'h10408000;
      25436: inst = 32'hc404734;
      25437: inst = 32'h8220000;
      25438: inst = 32'h10408000;
      25439: inst = 32'hc404735;
      25440: inst = 32'h8220000;
      25441: inst = 32'h10408000;
      25442: inst = 32'hc404736;
      25443: inst = 32'h8220000;
      25444: inst = 32'h10408000;
      25445: inst = 32'hc404737;
      25446: inst = 32'h8220000;
      25447: inst = 32'h10408000;
      25448: inst = 32'hc404738;
      25449: inst = 32'h8220000;
      25450: inst = 32'h10408000;
      25451: inst = 32'hc404739;
      25452: inst = 32'h8220000;
      25453: inst = 32'h10408000;
      25454: inst = 32'hc40473a;
      25455: inst = 32'h8220000;
      25456: inst = 32'h10408000;
      25457: inst = 32'hc40473b;
      25458: inst = 32'h8220000;
      25459: inst = 32'h10408000;
      25460: inst = 32'hc40473c;
      25461: inst = 32'h8220000;
      25462: inst = 32'h10408000;
      25463: inst = 32'hc40473d;
      25464: inst = 32'h8220000;
      25465: inst = 32'h10408000;
      25466: inst = 32'hc40473e;
      25467: inst = 32'h8220000;
      25468: inst = 32'h10408000;
      25469: inst = 32'hc40473f;
      25470: inst = 32'h8220000;
      25471: inst = 32'h10408000;
      25472: inst = 32'hc404740;
      25473: inst = 32'h8220000;
      25474: inst = 32'h10408000;
      25475: inst = 32'hc404741;
      25476: inst = 32'h8220000;
      25477: inst = 32'h10408000;
      25478: inst = 32'hc404744;
      25479: inst = 32'h8220000;
      25480: inst = 32'h10408000;
      25481: inst = 32'hc404745;
      25482: inst = 32'h8220000;
      25483: inst = 32'h10408000;
      25484: inst = 32'hc404746;
      25485: inst = 32'h8220000;
      25486: inst = 32'h10408000;
      25487: inst = 32'hc404747;
      25488: inst = 32'h8220000;
      25489: inst = 32'h10408000;
      25490: inst = 32'hc404748;
      25491: inst = 32'h8220000;
      25492: inst = 32'h10408000;
      25493: inst = 32'hc404749;
      25494: inst = 32'h8220000;
      25495: inst = 32'h10408000;
      25496: inst = 32'hc40474a;
      25497: inst = 32'h8220000;
      25498: inst = 32'h10408000;
      25499: inst = 32'hc40474b;
      25500: inst = 32'h8220000;
      25501: inst = 32'h10408000;
      25502: inst = 32'hc40474c;
      25503: inst = 32'h8220000;
      25504: inst = 32'h10408000;
      25505: inst = 32'hc40474d;
      25506: inst = 32'h8220000;
      25507: inst = 32'h10408000;
      25508: inst = 32'hc40474e;
      25509: inst = 32'h8220000;
      25510: inst = 32'h10408000;
      25511: inst = 32'hc40474f;
      25512: inst = 32'h8220000;
      25513: inst = 32'h10408000;
      25514: inst = 32'hc404750;
      25515: inst = 32'h8220000;
      25516: inst = 32'h10408000;
      25517: inst = 32'hc404753;
      25518: inst = 32'h8220000;
      25519: inst = 32'h10408000;
      25520: inst = 32'hc404754;
      25521: inst = 32'h8220000;
      25522: inst = 32'h10408000;
      25523: inst = 32'hc404755;
      25524: inst = 32'h8220000;
      25525: inst = 32'h10408000;
      25526: inst = 32'hc404756;
      25527: inst = 32'h8220000;
      25528: inst = 32'h10408000;
      25529: inst = 32'hc404757;
      25530: inst = 32'h8220000;
      25531: inst = 32'h10408000;
      25532: inst = 32'hc404758;
      25533: inst = 32'h8220000;
      25534: inst = 32'h10408000;
      25535: inst = 32'hc404767;
      25536: inst = 32'h8220000;
      25537: inst = 32'h10408000;
      25538: inst = 32'hc404768;
      25539: inst = 32'h8220000;
      25540: inst = 32'h10408000;
      25541: inst = 32'hc404769;
      25542: inst = 32'h8220000;
      25543: inst = 32'h10408000;
      25544: inst = 32'hc40476a;
      25545: inst = 32'h8220000;
      25546: inst = 32'h10408000;
      25547: inst = 32'hc40476b;
      25548: inst = 32'h8220000;
      25549: inst = 32'h10408000;
      25550: inst = 32'hc40476c;
      25551: inst = 32'h8220000;
      25552: inst = 32'h10408000;
      25553: inst = 32'hc40476d;
      25554: inst = 32'h8220000;
      25555: inst = 32'h10408000;
      25556: inst = 32'hc40476e;
      25557: inst = 32'h8220000;
      25558: inst = 32'h10408000;
      25559: inst = 32'hc404773;
      25560: inst = 32'h8220000;
      25561: inst = 32'h10408000;
      25562: inst = 32'hc404778;
      25563: inst = 32'h8220000;
      25564: inst = 32'h10408000;
      25565: inst = 32'hc40477d;
      25566: inst = 32'h8220000;
      25567: inst = 32'h10408000;
      25568: inst = 32'hc40477e;
      25569: inst = 32'h8220000;
      25570: inst = 32'h10408000;
      25571: inst = 32'hc40477f;
      25572: inst = 32'h8220000;
      25573: inst = 32'h10408000;
      25574: inst = 32'hc404780;
      25575: inst = 32'h8220000;
      25576: inst = 32'h10408000;
      25577: inst = 32'hc404781;
      25578: inst = 32'h8220000;
      25579: inst = 32'h10408000;
      25580: inst = 32'hc404782;
      25581: inst = 32'h8220000;
      25582: inst = 32'h10408000;
      25583: inst = 32'hc404787;
      25584: inst = 32'h8220000;
      25585: inst = 32'h10408000;
      25586: inst = 32'hc404788;
      25587: inst = 32'h8220000;
      25588: inst = 32'h10408000;
      25589: inst = 32'hc40478c;
      25590: inst = 32'h8220000;
      25591: inst = 32'h10408000;
      25592: inst = 32'hc40478d;
      25593: inst = 32'h8220000;
      25594: inst = 32'h10408000;
      25595: inst = 32'hc40478e;
      25596: inst = 32'h8220000;
      25597: inst = 32'h10408000;
      25598: inst = 32'hc40478f;
      25599: inst = 32'h8220000;
      25600: inst = 32'h10408000;
      25601: inst = 32'hc404790;
      25602: inst = 32'h8220000;
      25603: inst = 32'h10408000;
      25604: inst = 32'hc404791;
      25605: inst = 32'h8220000;
      25606: inst = 32'h10408000;
      25607: inst = 32'hc404792;
      25608: inst = 32'h8220000;
      25609: inst = 32'h10408000;
      25610: inst = 32'hc404796;
      25611: inst = 32'h8220000;
      25612: inst = 32'h10408000;
      25613: inst = 32'hc404797;
      25614: inst = 32'h8220000;
      25615: inst = 32'h10408000;
      25616: inst = 32'hc40479b;
      25617: inst = 32'h8220000;
      25618: inst = 32'h10408000;
      25619: inst = 32'hc4047a0;
      25620: inst = 32'h8220000;
      25621: inst = 32'h10408000;
      25622: inst = 32'hc4047a5;
      25623: inst = 32'h8220000;
      25624: inst = 32'h10408000;
      25625: inst = 32'hc4047a8;
      25626: inst = 32'h8220000;
      25627: inst = 32'h10408000;
      25628: inst = 32'hc4047ab;
      25629: inst = 32'h8220000;
      25630: inst = 32'h10408000;
      25631: inst = 32'hc4047af;
      25632: inst = 32'h8220000;
      25633: inst = 32'h10408000;
      25634: inst = 32'hc4047b0;
      25635: inst = 32'h8220000;
      25636: inst = 32'h10408000;
      25637: inst = 32'hc4047b3;
      25638: inst = 32'h8220000;
      25639: inst = 32'h10408000;
      25640: inst = 32'hc4047b4;
      25641: inst = 32'h8220000;
      25642: inst = 32'h10408000;
      25643: inst = 32'hc4047b5;
      25644: inst = 32'h8220000;
      25645: inst = 32'h10408000;
      25646: inst = 32'hc4047b6;
      25647: inst = 32'h8220000;
      25648: inst = 32'h10408000;
      25649: inst = 32'hc4047b7;
      25650: inst = 32'h8220000;
      25651: inst = 32'h10408000;
      25652: inst = 32'hc4047b8;
      25653: inst = 32'h8220000;
      25654: inst = 32'h10408000;
      25655: inst = 32'hc4047c7;
      25656: inst = 32'h8220000;
      25657: inst = 32'h10408000;
      25658: inst = 32'hc4047c8;
      25659: inst = 32'h8220000;
      25660: inst = 32'h10408000;
      25661: inst = 32'hc4047c9;
      25662: inst = 32'h8220000;
      25663: inst = 32'h10408000;
      25664: inst = 32'hc4047ca;
      25665: inst = 32'h8220000;
      25666: inst = 32'h10408000;
      25667: inst = 32'hc4047cb;
      25668: inst = 32'h8220000;
      25669: inst = 32'h10408000;
      25670: inst = 32'hc4047cc;
      25671: inst = 32'h8220000;
      25672: inst = 32'h10408000;
      25673: inst = 32'hc4047cd;
      25674: inst = 32'h8220000;
      25675: inst = 32'h10408000;
      25676: inst = 32'hc4047ce;
      25677: inst = 32'h8220000;
      25678: inst = 32'h10408000;
      25679: inst = 32'hc4047de;
      25680: inst = 32'h8220000;
      25681: inst = 32'h10408000;
      25682: inst = 32'hc4047df;
      25683: inst = 32'h8220000;
      25684: inst = 32'h10408000;
      25685: inst = 32'hc4047e0;
      25686: inst = 32'h8220000;
      25687: inst = 32'h10408000;
      25688: inst = 32'hc4047e1;
      25689: inst = 32'h8220000;
      25690: inst = 32'h10408000;
      25691: inst = 32'hc4047e2;
      25692: inst = 32'h8220000;
      25693: inst = 32'h10408000;
      25694: inst = 32'hc4047e7;
      25695: inst = 32'h8220000;
      25696: inst = 32'h10408000;
      25697: inst = 32'hc4047ed;
      25698: inst = 32'h8220000;
      25699: inst = 32'h10408000;
      25700: inst = 32'hc4047ee;
      25701: inst = 32'h8220000;
      25702: inst = 32'h10408000;
      25703: inst = 32'hc4047ef;
      25704: inst = 32'h8220000;
      25705: inst = 32'h10408000;
      25706: inst = 32'hc4047f0;
      25707: inst = 32'h8220000;
      25708: inst = 32'h10408000;
      25709: inst = 32'hc4047f1;
      25710: inst = 32'h8220000;
      25711: inst = 32'h10408000;
      25712: inst = 32'hc404810;
      25713: inst = 32'h8220000;
      25714: inst = 32'h10408000;
      25715: inst = 32'hc404813;
      25716: inst = 32'h8220000;
      25717: inst = 32'h10408000;
      25718: inst = 32'hc404814;
      25719: inst = 32'h8220000;
      25720: inst = 32'h10408000;
      25721: inst = 32'hc404815;
      25722: inst = 32'h8220000;
      25723: inst = 32'h10408000;
      25724: inst = 32'hc404816;
      25725: inst = 32'h8220000;
      25726: inst = 32'h10408000;
      25727: inst = 32'hc404817;
      25728: inst = 32'h8220000;
      25729: inst = 32'h10408000;
      25730: inst = 32'hc404818;
      25731: inst = 32'h8220000;
      25732: inst = 32'h10408000;
      25733: inst = 32'hc404827;
      25734: inst = 32'h8220000;
      25735: inst = 32'h10408000;
      25736: inst = 32'hc404828;
      25737: inst = 32'h8220000;
      25738: inst = 32'h10408000;
      25739: inst = 32'hc404829;
      25740: inst = 32'h8220000;
      25741: inst = 32'h10408000;
      25742: inst = 32'hc40482a;
      25743: inst = 32'h8220000;
      25744: inst = 32'h10408000;
      25745: inst = 32'hc40482b;
      25746: inst = 32'h8220000;
      25747: inst = 32'h10408000;
      25748: inst = 32'hc40482c;
      25749: inst = 32'h8220000;
      25750: inst = 32'h10408000;
      25751: inst = 32'hc40482d;
      25752: inst = 32'h8220000;
      25753: inst = 32'h10408000;
      25754: inst = 32'hc40482e;
      25755: inst = 32'h8220000;
      25756: inst = 32'h10408000;
      25757: inst = 32'hc404831;
      25758: inst = 32'h8220000;
      25759: inst = 32'h10408000;
      25760: inst = 32'hc404834;
      25761: inst = 32'h8220000;
      25762: inst = 32'h10408000;
      25763: inst = 32'hc404837;
      25764: inst = 32'h8220000;
      25765: inst = 32'h10408000;
      25766: inst = 32'hc404838;
      25767: inst = 32'h8220000;
      25768: inst = 32'h10408000;
      25769: inst = 32'hc40483b;
      25770: inst = 32'h8220000;
      25771: inst = 32'h10408000;
      25772: inst = 32'hc40483e;
      25773: inst = 32'h8220000;
      25774: inst = 32'h10408000;
      25775: inst = 32'hc40483f;
      25776: inst = 32'h8220000;
      25777: inst = 32'h10408000;
      25778: inst = 32'hc404840;
      25779: inst = 32'h8220000;
      25780: inst = 32'h10408000;
      25781: inst = 32'hc404841;
      25782: inst = 32'h8220000;
      25783: inst = 32'h10408000;
      25784: inst = 32'hc404842;
      25785: inst = 32'h8220000;
      25786: inst = 32'h10408000;
      25787: inst = 32'hc404843;
      25788: inst = 32'h8220000;
      25789: inst = 32'h10408000;
      25790: inst = 32'hc404846;
      25791: inst = 32'h8220000;
      25792: inst = 32'h10408000;
      25793: inst = 32'hc404849;
      25794: inst = 32'h8220000;
      25795: inst = 32'h10408000;
      25796: inst = 32'hc40484a;
      25797: inst = 32'h8220000;
      25798: inst = 32'h10408000;
      25799: inst = 32'hc40484d;
      25800: inst = 32'h8220000;
      25801: inst = 32'h10408000;
      25802: inst = 32'hc40484e;
      25803: inst = 32'h8220000;
      25804: inst = 32'h10408000;
      25805: inst = 32'hc40484f;
      25806: inst = 32'h8220000;
      25807: inst = 32'h10408000;
      25808: inst = 32'hc404850;
      25809: inst = 32'h8220000;
      25810: inst = 32'h10408000;
      25811: inst = 32'hc404851;
      25812: inst = 32'h8220000;
      25813: inst = 32'h10408000;
      25814: inst = 32'hc404854;
      25815: inst = 32'h8220000;
      25816: inst = 32'h10408000;
      25817: inst = 32'hc404858;
      25818: inst = 32'h8220000;
      25819: inst = 32'h10408000;
      25820: inst = 32'hc404859;
      25821: inst = 32'h8220000;
      25822: inst = 32'h10408000;
      25823: inst = 32'hc40485e;
      25824: inst = 32'h8220000;
      25825: inst = 32'h10408000;
      25826: inst = 32'hc404861;
      25827: inst = 32'h8220000;
      25828: inst = 32'h10408000;
      25829: inst = 32'hc404864;
      25830: inst = 32'h8220000;
      25831: inst = 32'h10408000;
      25832: inst = 32'hc404865;
      25833: inst = 32'h8220000;
      25834: inst = 32'h10408000;
      25835: inst = 32'hc404869;
      25836: inst = 32'h8220000;
      25837: inst = 32'h10408000;
      25838: inst = 32'hc40486c;
      25839: inst = 32'h8220000;
      25840: inst = 32'h10408000;
      25841: inst = 32'hc40486d;
      25842: inst = 32'h8220000;
      25843: inst = 32'h10408000;
      25844: inst = 32'hc404870;
      25845: inst = 32'h8220000;
      25846: inst = 32'h10408000;
      25847: inst = 32'hc404873;
      25848: inst = 32'h8220000;
      25849: inst = 32'h10408000;
      25850: inst = 32'hc404874;
      25851: inst = 32'h8220000;
      25852: inst = 32'h10408000;
      25853: inst = 32'hc404875;
      25854: inst = 32'h8220000;
      25855: inst = 32'h10408000;
      25856: inst = 32'hc404876;
      25857: inst = 32'h8220000;
      25858: inst = 32'h10408000;
      25859: inst = 32'hc404877;
      25860: inst = 32'h8220000;
      25861: inst = 32'h10408000;
      25862: inst = 32'hc404878;
      25863: inst = 32'h8220000;
      25864: inst = 32'h10408000;
      25865: inst = 32'hc404887;
      25866: inst = 32'h8220000;
      25867: inst = 32'h10408000;
      25868: inst = 32'hc404888;
      25869: inst = 32'h8220000;
      25870: inst = 32'h10408000;
      25871: inst = 32'hc404889;
      25872: inst = 32'h8220000;
      25873: inst = 32'h10408000;
      25874: inst = 32'hc40488a;
      25875: inst = 32'h8220000;
      25876: inst = 32'h10408000;
      25877: inst = 32'hc40488b;
      25878: inst = 32'h8220000;
      25879: inst = 32'h10408000;
      25880: inst = 32'hc40488c;
      25881: inst = 32'h8220000;
      25882: inst = 32'h10408000;
      25883: inst = 32'hc40488d;
      25884: inst = 32'h8220000;
      25885: inst = 32'h10408000;
      25886: inst = 32'hc40488e;
      25887: inst = 32'h8220000;
      25888: inst = 32'h10408000;
      25889: inst = 32'hc404891;
      25890: inst = 32'h8220000;
      25891: inst = 32'h10408000;
      25892: inst = 32'hc404894;
      25893: inst = 32'h8220000;
      25894: inst = 32'h10408000;
      25895: inst = 32'hc404897;
      25896: inst = 32'h8220000;
      25897: inst = 32'h10408000;
      25898: inst = 32'hc404898;
      25899: inst = 32'h8220000;
      25900: inst = 32'h10408000;
      25901: inst = 32'hc40489b;
      25902: inst = 32'h8220000;
      25903: inst = 32'h10408000;
      25904: inst = 32'hc40489e;
      25905: inst = 32'h8220000;
      25906: inst = 32'h10408000;
      25907: inst = 32'hc40489f;
      25908: inst = 32'h8220000;
      25909: inst = 32'h10408000;
      25910: inst = 32'hc4048a0;
      25911: inst = 32'h8220000;
      25912: inst = 32'h10408000;
      25913: inst = 32'hc4048a1;
      25914: inst = 32'h8220000;
      25915: inst = 32'h10408000;
      25916: inst = 32'hc4048a2;
      25917: inst = 32'h8220000;
      25918: inst = 32'h10408000;
      25919: inst = 32'hc4048a3;
      25920: inst = 32'h8220000;
      25921: inst = 32'h10408000;
      25922: inst = 32'hc4048a6;
      25923: inst = 32'h8220000;
      25924: inst = 32'h10408000;
      25925: inst = 32'hc4048a9;
      25926: inst = 32'h8220000;
      25927: inst = 32'h10408000;
      25928: inst = 32'hc4048aa;
      25929: inst = 32'h8220000;
      25930: inst = 32'h10408000;
      25931: inst = 32'hc4048ad;
      25932: inst = 32'h8220000;
      25933: inst = 32'h10408000;
      25934: inst = 32'hc4048ae;
      25935: inst = 32'h8220000;
      25936: inst = 32'h10408000;
      25937: inst = 32'hc4048af;
      25938: inst = 32'h8220000;
      25939: inst = 32'h10408000;
      25940: inst = 32'hc4048b0;
      25941: inst = 32'h8220000;
      25942: inst = 32'h10408000;
      25943: inst = 32'hc4048b3;
      25944: inst = 32'h8220000;
      25945: inst = 32'h10408000;
      25946: inst = 32'hc4048b4;
      25947: inst = 32'h8220000;
      25948: inst = 32'h10408000;
      25949: inst = 32'hc4048b5;
      25950: inst = 32'h8220000;
      25951: inst = 32'h10408000;
      25952: inst = 32'hc4048b8;
      25953: inst = 32'h8220000;
      25954: inst = 32'h10408000;
      25955: inst = 32'hc4048b9;
      25956: inst = 32'h8220000;
      25957: inst = 32'h10408000;
      25958: inst = 32'hc4048be;
      25959: inst = 32'h8220000;
      25960: inst = 32'h10408000;
      25961: inst = 32'hc4048c1;
      25962: inst = 32'h8220000;
      25963: inst = 32'h10408000;
      25964: inst = 32'hc4048c4;
      25965: inst = 32'h8220000;
      25966: inst = 32'h10408000;
      25967: inst = 32'hc4048c5;
      25968: inst = 32'h8220000;
      25969: inst = 32'h10408000;
      25970: inst = 32'hc4048c8;
      25971: inst = 32'h8220000;
      25972: inst = 32'h10408000;
      25973: inst = 32'hc4048c9;
      25974: inst = 32'h8220000;
      25975: inst = 32'h10408000;
      25976: inst = 32'hc4048cc;
      25977: inst = 32'h8220000;
      25978: inst = 32'h10408000;
      25979: inst = 32'hc4048cd;
      25980: inst = 32'h8220000;
      25981: inst = 32'h10408000;
      25982: inst = 32'hc4048d0;
      25983: inst = 32'h8220000;
      25984: inst = 32'h10408000;
      25985: inst = 32'hc4048d3;
      25986: inst = 32'h8220000;
      25987: inst = 32'h10408000;
      25988: inst = 32'hc4048d4;
      25989: inst = 32'h8220000;
      25990: inst = 32'h10408000;
      25991: inst = 32'hc4048d5;
      25992: inst = 32'h8220000;
      25993: inst = 32'h10408000;
      25994: inst = 32'hc4048d6;
      25995: inst = 32'h8220000;
      25996: inst = 32'h10408000;
      25997: inst = 32'hc4048d7;
      25998: inst = 32'h8220000;
      25999: inst = 32'h10408000;
      26000: inst = 32'hc4048d8;
      26001: inst = 32'h8220000;
      26002: inst = 32'h10408000;
      26003: inst = 32'hc4048e7;
      26004: inst = 32'h8220000;
      26005: inst = 32'h10408000;
      26006: inst = 32'hc4048e8;
      26007: inst = 32'h8220000;
      26008: inst = 32'h10408000;
      26009: inst = 32'hc4048e9;
      26010: inst = 32'h8220000;
      26011: inst = 32'h10408000;
      26012: inst = 32'hc4048ea;
      26013: inst = 32'h8220000;
      26014: inst = 32'h10408000;
      26015: inst = 32'hc4048eb;
      26016: inst = 32'h8220000;
      26017: inst = 32'h10408000;
      26018: inst = 32'hc4048ec;
      26019: inst = 32'h8220000;
      26020: inst = 32'h10408000;
      26021: inst = 32'hc4048ed;
      26022: inst = 32'h8220000;
      26023: inst = 32'h10408000;
      26024: inst = 32'hc4048ee;
      26025: inst = 32'h8220000;
      26026: inst = 32'h10408000;
      26027: inst = 32'hc4048f1;
      26028: inst = 32'h8220000;
      26029: inst = 32'h10408000;
      26030: inst = 32'hc4048f4;
      26031: inst = 32'h8220000;
      26032: inst = 32'h10408000;
      26033: inst = 32'hc4048f7;
      26034: inst = 32'h8220000;
      26035: inst = 32'h10408000;
      26036: inst = 32'hc4048f8;
      26037: inst = 32'h8220000;
      26038: inst = 32'h10408000;
      26039: inst = 32'hc4048fb;
      26040: inst = 32'h8220000;
      26041: inst = 32'h10408000;
      26042: inst = 32'hc4048fe;
      26043: inst = 32'h8220000;
      26044: inst = 32'h10408000;
      26045: inst = 32'hc4048ff;
      26046: inst = 32'h8220000;
      26047: inst = 32'h10408000;
      26048: inst = 32'hc404900;
      26049: inst = 32'h8220000;
      26050: inst = 32'h10408000;
      26051: inst = 32'hc404901;
      26052: inst = 32'h8220000;
      26053: inst = 32'h10408000;
      26054: inst = 32'hc404902;
      26055: inst = 32'h8220000;
      26056: inst = 32'h10408000;
      26057: inst = 32'hc404903;
      26058: inst = 32'h8220000;
      26059: inst = 32'h10408000;
      26060: inst = 32'hc404906;
      26061: inst = 32'h8220000;
      26062: inst = 32'h10408000;
      26063: inst = 32'hc404909;
      26064: inst = 32'h8220000;
      26065: inst = 32'h10408000;
      26066: inst = 32'hc40490a;
      26067: inst = 32'h8220000;
      26068: inst = 32'h10408000;
      26069: inst = 32'hc40490d;
      26070: inst = 32'h8220000;
      26071: inst = 32'h10408000;
      26072: inst = 32'hc40490e;
      26073: inst = 32'h8220000;
      26074: inst = 32'h10408000;
      26075: inst = 32'hc40490f;
      26076: inst = 32'h8220000;
      26077: inst = 32'h10408000;
      26078: inst = 32'hc404910;
      26079: inst = 32'h8220000;
      26080: inst = 32'h10408000;
      26081: inst = 32'hc404913;
      26082: inst = 32'h8220000;
      26083: inst = 32'h10408000;
      26084: inst = 32'hc404914;
      26085: inst = 32'h8220000;
      26086: inst = 32'h10408000;
      26087: inst = 32'hc404915;
      26088: inst = 32'h8220000;
      26089: inst = 32'h10408000;
      26090: inst = 32'hc404918;
      26091: inst = 32'h8220000;
      26092: inst = 32'h10408000;
      26093: inst = 32'hc404919;
      26094: inst = 32'h8220000;
      26095: inst = 32'h10408000;
      26096: inst = 32'hc40491e;
      26097: inst = 32'h8220000;
      26098: inst = 32'h10408000;
      26099: inst = 32'hc404921;
      26100: inst = 32'h8220000;
      26101: inst = 32'h10408000;
      26102: inst = 32'hc404924;
      26103: inst = 32'h8220000;
      26104: inst = 32'h10408000;
      26105: inst = 32'hc404925;
      26106: inst = 32'h8220000;
      26107: inst = 32'h10408000;
      26108: inst = 32'hc404928;
      26109: inst = 32'h8220000;
      26110: inst = 32'h10408000;
      26111: inst = 32'hc404929;
      26112: inst = 32'h8220000;
      26113: inst = 32'h10408000;
      26114: inst = 32'hc40492c;
      26115: inst = 32'h8220000;
      26116: inst = 32'h10408000;
      26117: inst = 32'hc40492d;
      26118: inst = 32'h8220000;
      26119: inst = 32'h10408000;
      26120: inst = 32'hc404930;
      26121: inst = 32'h8220000;
      26122: inst = 32'h10408000;
      26123: inst = 32'hc404933;
      26124: inst = 32'h8220000;
      26125: inst = 32'h10408000;
      26126: inst = 32'hc404934;
      26127: inst = 32'h8220000;
      26128: inst = 32'h10408000;
      26129: inst = 32'hc404935;
      26130: inst = 32'h8220000;
      26131: inst = 32'h10408000;
      26132: inst = 32'hc404936;
      26133: inst = 32'h8220000;
      26134: inst = 32'h10408000;
      26135: inst = 32'hc404937;
      26136: inst = 32'h8220000;
      26137: inst = 32'h10408000;
      26138: inst = 32'hc404938;
      26139: inst = 32'h8220000;
      26140: inst = 32'h10408000;
      26141: inst = 32'hc404947;
      26142: inst = 32'h8220000;
      26143: inst = 32'h10408000;
      26144: inst = 32'hc404948;
      26145: inst = 32'h8220000;
      26146: inst = 32'h10408000;
      26147: inst = 32'hc404949;
      26148: inst = 32'h8220000;
      26149: inst = 32'h10408000;
      26150: inst = 32'hc40494a;
      26151: inst = 32'h8220000;
      26152: inst = 32'h10408000;
      26153: inst = 32'hc40494b;
      26154: inst = 32'h8220000;
      26155: inst = 32'h10408000;
      26156: inst = 32'hc40494c;
      26157: inst = 32'h8220000;
      26158: inst = 32'h10408000;
      26159: inst = 32'hc40494d;
      26160: inst = 32'h8220000;
      26161: inst = 32'h10408000;
      26162: inst = 32'hc40494e;
      26163: inst = 32'h8220000;
      26164: inst = 32'h10408000;
      26165: inst = 32'hc404951;
      26166: inst = 32'h8220000;
      26167: inst = 32'h10408000;
      26168: inst = 32'hc404954;
      26169: inst = 32'h8220000;
      26170: inst = 32'h10408000;
      26171: inst = 32'hc404957;
      26172: inst = 32'h8220000;
      26173: inst = 32'h10408000;
      26174: inst = 32'hc40495b;
      26175: inst = 32'h8220000;
      26176: inst = 32'h10408000;
      26177: inst = 32'hc40495e;
      26178: inst = 32'h8220000;
      26179: inst = 32'h10408000;
      26180: inst = 32'hc40495f;
      26181: inst = 32'h8220000;
      26182: inst = 32'h10408000;
      26183: inst = 32'hc404960;
      26184: inst = 32'h8220000;
      26185: inst = 32'h10408000;
      26186: inst = 32'hc404961;
      26187: inst = 32'h8220000;
      26188: inst = 32'h10408000;
      26189: inst = 32'hc404962;
      26190: inst = 32'h8220000;
      26191: inst = 32'h10408000;
      26192: inst = 32'hc404963;
      26193: inst = 32'h8220000;
      26194: inst = 32'h10408000;
      26195: inst = 32'hc404966;
      26196: inst = 32'h8220000;
      26197: inst = 32'h10408000;
      26198: inst = 32'hc404969;
      26199: inst = 32'h8220000;
      26200: inst = 32'h10408000;
      26201: inst = 32'hc40496a;
      26202: inst = 32'h8220000;
      26203: inst = 32'h10408000;
      26204: inst = 32'hc40496d;
      26205: inst = 32'h8220000;
      26206: inst = 32'h10408000;
      26207: inst = 32'hc40496e;
      26208: inst = 32'h8220000;
      26209: inst = 32'h10408000;
      26210: inst = 32'hc40496f;
      26211: inst = 32'h8220000;
      26212: inst = 32'h10408000;
      26213: inst = 32'hc404970;
      26214: inst = 32'h8220000;
      26215: inst = 32'h10408000;
      26216: inst = 32'hc404974;
      26217: inst = 32'h8220000;
      26218: inst = 32'h10408000;
      26219: inst = 32'hc404975;
      26220: inst = 32'h8220000;
      26221: inst = 32'h10408000;
      26222: inst = 32'hc404978;
      26223: inst = 32'h8220000;
      26224: inst = 32'h10408000;
      26225: inst = 32'hc404979;
      26226: inst = 32'h8220000;
      26227: inst = 32'h10408000;
      26228: inst = 32'hc40497e;
      26229: inst = 32'h8220000;
      26230: inst = 32'h10408000;
      26231: inst = 32'hc404981;
      26232: inst = 32'h8220000;
      26233: inst = 32'h10408000;
      26234: inst = 32'hc404984;
      26235: inst = 32'h8220000;
      26236: inst = 32'h10408000;
      26237: inst = 32'hc404988;
      26238: inst = 32'h8220000;
      26239: inst = 32'h10408000;
      26240: inst = 32'hc404989;
      26241: inst = 32'h8220000;
      26242: inst = 32'h10408000;
      26243: inst = 32'hc40498c;
      26244: inst = 32'h8220000;
      26245: inst = 32'h10408000;
      26246: inst = 32'hc40498d;
      26247: inst = 32'h8220000;
      26248: inst = 32'h10408000;
      26249: inst = 32'hc404990;
      26250: inst = 32'h8220000;
      26251: inst = 32'h10408000;
      26252: inst = 32'hc404993;
      26253: inst = 32'h8220000;
      26254: inst = 32'h10408000;
      26255: inst = 32'hc404994;
      26256: inst = 32'h8220000;
      26257: inst = 32'h10408000;
      26258: inst = 32'hc404995;
      26259: inst = 32'h8220000;
      26260: inst = 32'h10408000;
      26261: inst = 32'hc404996;
      26262: inst = 32'h8220000;
      26263: inst = 32'h10408000;
      26264: inst = 32'hc404997;
      26265: inst = 32'h8220000;
      26266: inst = 32'h10408000;
      26267: inst = 32'hc404998;
      26268: inst = 32'h8220000;
      26269: inst = 32'h10408000;
      26270: inst = 32'hc4049a7;
      26271: inst = 32'h8220000;
      26272: inst = 32'h10408000;
      26273: inst = 32'hc4049a8;
      26274: inst = 32'h8220000;
      26275: inst = 32'h10408000;
      26276: inst = 32'hc4049a9;
      26277: inst = 32'h8220000;
      26278: inst = 32'h10408000;
      26279: inst = 32'hc4049aa;
      26280: inst = 32'h8220000;
      26281: inst = 32'h10408000;
      26282: inst = 32'hc4049ab;
      26283: inst = 32'h8220000;
      26284: inst = 32'h10408000;
      26285: inst = 32'hc4049ac;
      26286: inst = 32'h8220000;
      26287: inst = 32'h10408000;
      26288: inst = 32'hc4049ad;
      26289: inst = 32'h8220000;
      26290: inst = 32'h10408000;
      26291: inst = 32'hc4049ae;
      26292: inst = 32'h8220000;
      26293: inst = 32'h10408000;
      26294: inst = 32'hc4049b4;
      26295: inst = 32'h8220000;
      26296: inst = 32'h10408000;
      26297: inst = 32'hc4049bb;
      26298: inst = 32'h8220000;
      26299: inst = 32'h10408000;
      26300: inst = 32'hc4049be;
      26301: inst = 32'h8220000;
      26302: inst = 32'h10408000;
      26303: inst = 32'hc4049bf;
      26304: inst = 32'h8220000;
      26305: inst = 32'h10408000;
      26306: inst = 32'hc4049c0;
      26307: inst = 32'h8220000;
      26308: inst = 32'h10408000;
      26309: inst = 32'hc4049c1;
      26310: inst = 32'h8220000;
      26311: inst = 32'h10408000;
      26312: inst = 32'hc4049c2;
      26313: inst = 32'h8220000;
      26314: inst = 32'h10408000;
      26315: inst = 32'hc4049c3;
      26316: inst = 32'h8220000;
      26317: inst = 32'h10408000;
      26318: inst = 32'hc4049cd;
      26319: inst = 32'h8220000;
      26320: inst = 32'h10408000;
      26321: inst = 32'hc4049ce;
      26322: inst = 32'h8220000;
      26323: inst = 32'h10408000;
      26324: inst = 32'hc4049cf;
      26325: inst = 32'h8220000;
      26326: inst = 32'h10408000;
      26327: inst = 32'hc4049d0;
      26328: inst = 32'h8220000;
      26329: inst = 32'h10408000;
      26330: inst = 32'hc4049d1;
      26331: inst = 32'h8220000;
      26332: inst = 32'h10408000;
      26333: inst = 32'hc4049de;
      26334: inst = 32'h8220000;
      26335: inst = 32'h10408000;
      26336: inst = 32'hc4049e1;
      26337: inst = 32'h8220000;
      26338: inst = 32'h10408000;
      26339: inst = 32'hc4049ea;
      26340: inst = 32'h8220000;
      26341: inst = 32'h10408000;
      26342: inst = 32'hc4049f5;
      26343: inst = 32'h8220000;
      26344: inst = 32'h10408000;
      26345: inst = 32'hc4049f6;
      26346: inst = 32'h8220000;
      26347: inst = 32'h10408000;
      26348: inst = 32'hc4049f7;
      26349: inst = 32'h8220000;
      26350: inst = 32'h10408000;
      26351: inst = 32'hc4049f8;
      26352: inst = 32'h8220000;
      26353: inst = 32'h10408000;
      26354: inst = 32'hc404a07;
      26355: inst = 32'h8220000;
      26356: inst = 32'h10408000;
      26357: inst = 32'hc404a08;
      26358: inst = 32'h8220000;
      26359: inst = 32'h10408000;
      26360: inst = 32'hc404a09;
      26361: inst = 32'h8220000;
      26362: inst = 32'h10408000;
      26363: inst = 32'hc404a0a;
      26364: inst = 32'h8220000;
      26365: inst = 32'h10408000;
      26366: inst = 32'hc404a0b;
      26367: inst = 32'h8220000;
      26368: inst = 32'h10408000;
      26369: inst = 32'hc404a0c;
      26370: inst = 32'h8220000;
      26371: inst = 32'h10408000;
      26372: inst = 32'hc404a0d;
      26373: inst = 32'h8220000;
      26374: inst = 32'h10408000;
      26375: inst = 32'hc404a0e;
      26376: inst = 32'h8220000;
      26377: inst = 32'h10408000;
      26378: inst = 32'hc404a0f;
      26379: inst = 32'h8220000;
      26380: inst = 32'h10408000;
      26381: inst = 32'hc404a12;
      26382: inst = 32'h8220000;
      26383: inst = 32'h10408000;
      26384: inst = 32'hc404a13;
      26385: inst = 32'h8220000;
      26386: inst = 32'h10408000;
      26387: inst = 32'hc404a14;
      26388: inst = 32'h8220000;
      26389: inst = 32'h10408000;
      26390: inst = 32'hc404a15;
      26391: inst = 32'h8220000;
      26392: inst = 32'h10408000;
      26393: inst = 32'hc404a1b;
      26394: inst = 32'h8220000;
      26395: inst = 32'h10408000;
      26396: inst = 32'hc404a1e;
      26397: inst = 32'h8220000;
      26398: inst = 32'h10408000;
      26399: inst = 32'hc404a1f;
      26400: inst = 32'h8220000;
      26401: inst = 32'h10408000;
      26402: inst = 32'hc404a20;
      26403: inst = 32'h8220000;
      26404: inst = 32'h10408000;
      26405: inst = 32'hc404a21;
      26406: inst = 32'h8220000;
      26407: inst = 32'h10408000;
      26408: inst = 32'hc404a22;
      26409: inst = 32'h8220000;
      26410: inst = 32'h10408000;
      26411: inst = 32'hc404a23;
      26412: inst = 32'h8220000;
      26413: inst = 32'h10408000;
      26414: inst = 32'hc404a24;
      26415: inst = 32'h8220000;
      26416: inst = 32'h10408000;
      26417: inst = 32'hc404a27;
      26418: inst = 32'h8220000;
      26419: inst = 32'h10408000;
      26420: inst = 32'hc404a28;
      26421: inst = 32'h8220000;
      26422: inst = 32'h10408000;
      26423: inst = 32'hc404a2b;
      26424: inst = 32'h8220000;
      26425: inst = 32'h10408000;
      26426: inst = 32'hc404a2c;
      26427: inst = 32'h8220000;
      26428: inst = 32'h10408000;
      26429: inst = 32'hc404a2d;
      26430: inst = 32'h8220000;
      26431: inst = 32'h10408000;
      26432: inst = 32'hc404a2e;
      26433: inst = 32'h8220000;
      26434: inst = 32'h10408000;
      26435: inst = 32'hc404a2f;
      26436: inst = 32'h8220000;
      26437: inst = 32'h10408000;
      26438: inst = 32'hc404a30;
      26439: inst = 32'h8220000;
      26440: inst = 32'h10408000;
      26441: inst = 32'hc404a31;
      26442: inst = 32'h8220000;
      26443: inst = 32'h10408000;
      26444: inst = 32'hc404a32;
      26445: inst = 32'h8220000;
      26446: inst = 32'h10408000;
      26447: inst = 32'hc404a36;
      26448: inst = 32'h8220000;
      26449: inst = 32'h10408000;
      26450: inst = 32'hc404a37;
      26451: inst = 32'h8220000;
      26452: inst = 32'h10408000;
      26453: inst = 32'hc404a3a;
      26454: inst = 32'h8220000;
      26455: inst = 32'h10408000;
      26456: inst = 32'hc404a3e;
      26457: inst = 32'h8220000;
      26458: inst = 32'h10408000;
      26459: inst = 32'hc404a41;
      26460: inst = 32'h8220000;
      26461: inst = 32'h10408000;
      26462: inst = 32'hc404a42;
      26463: inst = 32'h8220000;
      26464: inst = 32'h10408000;
      26465: inst = 32'hc404a49;
      26466: inst = 32'h8220000;
      26467: inst = 32'h10408000;
      26468: inst = 32'hc404a4a;
      26469: inst = 32'h8220000;
      26470: inst = 32'h10408000;
      26471: inst = 32'hc404a4b;
      26472: inst = 32'h8220000;
      26473: inst = 32'h10408000;
      26474: inst = 32'hc404a4e;
      26475: inst = 32'h8220000;
      26476: inst = 32'h10408000;
      26477: inst = 32'hc404a4f;
      26478: inst = 32'h8220000;
      26479: inst = 32'h10408000;
      26480: inst = 32'hc404a54;
      26481: inst = 32'h8220000;
      26482: inst = 32'h10408000;
      26483: inst = 32'hc404a55;
      26484: inst = 32'h8220000;
      26485: inst = 32'h10408000;
      26486: inst = 32'hc404a56;
      26487: inst = 32'h8220000;
      26488: inst = 32'h10408000;
      26489: inst = 32'hc404a57;
      26490: inst = 32'h8220000;
      26491: inst = 32'h10408000;
      26492: inst = 32'hc404a58;
      26493: inst = 32'h8220000;
      26494: inst = 32'h10408000;
      26495: inst = 32'hc404a67;
      26496: inst = 32'h8220000;
      26497: inst = 32'h10408000;
      26498: inst = 32'hc404a68;
      26499: inst = 32'h8220000;
      26500: inst = 32'h10408000;
      26501: inst = 32'hc404a69;
      26502: inst = 32'h8220000;
      26503: inst = 32'h10408000;
      26504: inst = 32'hc404a6a;
      26505: inst = 32'h8220000;
      26506: inst = 32'h10408000;
      26507: inst = 32'hc404a6b;
      26508: inst = 32'h8220000;
      26509: inst = 32'h10408000;
      26510: inst = 32'hc404a6c;
      26511: inst = 32'h8220000;
      26512: inst = 32'h10408000;
      26513: inst = 32'hc404a6d;
      26514: inst = 32'h8220000;
      26515: inst = 32'h10408000;
      26516: inst = 32'hc404a6e;
      26517: inst = 32'h8220000;
      26518: inst = 32'h10408000;
      26519: inst = 32'hc404a6f;
      26520: inst = 32'h8220000;
      26521: inst = 32'h10408000;
      26522: inst = 32'hc404a70;
      26523: inst = 32'h8220000;
      26524: inst = 32'h10408000;
      26525: inst = 32'hc404a71;
      26526: inst = 32'h8220000;
      26527: inst = 32'h10408000;
      26528: inst = 32'hc404a72;
      26529: inst = 32'h8220000;
      26530: inst = 32'h10408000;
      26531: inst = 32'hc404a73;
      26532: inst = 32'h8220000;
      26533: inst = 32'h10408000;
      26534: inst = 32'hc404a74;
      26535: inst = 32'h8220000;
      26536: inst = 32'h10408000;
      26537: inst = 32'hc404a75;
      26538: inst = 32'h8220000;
      26539: inst = 32'h10408000;
      26540: inst = 32'hc404a76;
      26541: inst = 32'h8220000;
      26542: inst = 32'h10408000;
      26543: inst = 32'hc404a77;
      26544: inst = 32'h8220000;
      26545: inst = 32'h10408000;
      26546: inst = 32'hc404a78;
      26547: inst = 32'h8220000;
      26548: inst = 32'h10408000;
      26549: inst = 32'hc404a79;
      26550: inst = 32'h8220000;
      26551: inst = 32'h10408000;
      26552: inst = 32'hc404a7a;
      26553: inst = 32'h8220000;
      26554: inst = 32'h10408000;
      26555: inst = 32'hc404a7b;
      26556: inst = 32'h8220000;
      26557: inst = 32'h10408000;
      26558: inst = 32'hc404a7c;
      26559: inst = 32'h8220000;
      26560: inst = 32'h10408000;
      26561: inst = 32'hc404a7d;
      26562: inst = 32'h8220000;
      26563: inst = 32'h10408000;
      26564: inst = 32'hc404a7e;
      26565: inst = 32'h8220000;
      26566: inst = 32'h10408000;
      26567: inst = 32'hc404a7f;
      26568: inst = 32'h8220000;
      26569: inst = 32'h10408000;
      26570: inst = 32'hc404a80;
      26571: inst = 32'h8220000;
      26572: inst = 32'h10408000;
      26573: inst = 32'hc404a81;
      26574: inst = 32'h8220000;
      26575: inst = 32'h10408000;
      26576: inst = 32'hc404a82;
      26577: inst = 32'h8220000;
      26578: inst = 32'h10408000;
      26579: inst = 32'hc404a83;
      26580: inst = 32'h8220000;
      26581: inst = 32'h10408000;
      26582: inst = 32'hc404a84;
      26583: inst = 32'h8220000;
      26584: inst = 32'h10408000;
      26585: inst = 32'hc404a85;
      26586: inst = 32'h8220000;
      26587: inst = 32'h10408000;
      26588: inst = 32'hc404a86;
      26589: inst = 32'h8220000;
      26590: inst = 32'h10408000;
      26591: inst = 32'hc404a87;
      26592: inst = 32'h8220000;
      26593: inst = 32'h10408000;
      26594: inst = 32'hc404a88;
      26595: inst = 32'h8220000;
      26596: inst = 32'h10408000;
      26597: inst = 32'hc404a89;
      26598: inst = 32'h8220000;
      26599: inst = 32'h10408000;
      26600: inst = 32'hc404a8a;
      26601: inst = 32'h8220000;
      26602: inst = 32'h10408000;
      26603: inst = 32'hc404a8b;
      26604: inst = 32'h8220000;
      26605: inst = 32'h10408000;
      26606: inst = 32'hc404a8c;
      26607: inst = 32'h8220000;
      26608: inst = 32'h10408000;
      26609: inst = 32'hc404a8d;
      26610: inst = 32'h8220000;
      26611: inst = 32'h10408000;
      26612: inst = 32'hc404a8e;
      26613: inst = 32'h8220000;
      26614: inst = 32'h10408000;
      26615: inst = 32'hc404a8f;
      26616: inst = 32'h8220000;
      26617: inst = 32'h10408000;
      26618: inst = 32'hc404a90;
      26619: inst = 32'h8220000;
      26620: inst = 32'h10408000;
      26621: inst = 32'hc404a91;
      26622: inst = 32'h8220000;
      26623: inst = 32'h10408000;
      26624: inst = 32'hc404a92;
      26625: inst = 32'h8220000;
      26626: inst = 32'h10408000;
      26627: inst = 32'hc404a93;
      26628: inst = 32'h8220000;
      26629: inst = 32'h10408000;
      26630: inst = 32'hc404a94;
      26631: inst = 32'h8220000;
      26632: inst = 32'h10408000;
      26633: inst = 32'hc404a95;
      26634: inst = 32'h8220000;
      26635: inst = 32'h10408000;
      26636: inst = 32'hc404a96;
      26637: inst = 32'h8220000;
      26638: inst = 32'h10408000;
      26639: inst = 32'hc404a97;
      26640: inst = 32'h8220000;
      26641: inst = 32'h10408000;
      26642: inst = 32'hc404a98;
      26643: inst = 32'h8220000;
      26644: inst = 32'h10408000;
      26645: inst = 32'hc404a99;
      26646: inst = 32'h8220000;
      26647: inst = 32'h10408000;
      26648: inst = 32'hc404a9a;
      26649: inst = 32'h8220000;
      26650: inst = 32'h10408000;
      26651: inst = 32'hc404a9b;
      26652: inst = 32'h8220000;
      26653: inst = 32'h10408000;
      26654: inst = 32'hc404a9c;
      26655: inst = 32'h8220000;
      26656: inst = 32'h10408000;
      26657: inst = 32'hc404a9d;
      26658: inst = 32'h8220000;
      26659: inst = 32'h10408000;
      26660: inst = 32'hc404a9e;
      26661: inst = 32'h8220000;
      26662: inst = 32'h10408000;
      26663: inst = 32'hc404a9f;
      26664: inst = 32'h8220000;
      26665: inst = 32'h10408000;
      26666: inst = 32'hc404aa0;
      26667: inst = 32'h8220000;
      26668: inst = 32'h10408000;
      26669: inst = 32'hc404aa1;
      26670: inst = 32'h8220000;
      26671: inst = 32'h10408000;
      26672: inst = 32'hc404aa2;
      26673: inst = 32'h8220000;
      26674: inst = 32'h10408000;
      26675: inst = 32'hc404aa3;
      26676: inst = 32'h8220000;
      26677: inst = 32'h10408000;
      26678: inst = 32'hc404aa4;
      26679: inst = 32'h8220000;
      26680: inst = 32'h10408000;
      26681: inst = 32'hc404aa5;
      26682: inst = 32'h8220000;
      26683: inst = 32'h10408000;
      26684: inst = 32'hc404aa6;
      26685: inst = 32'h8220000;
      26686: inst = 32'h10408000;
      26687: inst = 32'hc404aa7;
      26688: inst = 32'h8220000;
      26689: inst = 32'h10408000;
      26690: inst = 32'hc404aa8;
      26691: inst = 32'h8220000;
      26692: inst = 32'h10408000;
      26693: inst = 32'hc404aa9;
      26694: inst = 32'h8220000;
      26695: inst = 32'h10408000;
      26696: inst = 32'hc404aaa;
      26697: inst = 32'h8220000;
      26698: inst = 32'h10408000;
      26699: inst = 32'hc404aab;
      26700: inst = 32'h8220000;
      26701: inst = 32'h10408000;
      26702: inst = 32'hc404aac;
      26703: inst = 32'h8220000;
      26704: inst = 32'h10408000;
      26705: inst = 32'hc404aad;
      26706: inst = 32'h8220000;
      26707: inst = 32'h10408000;
      26708: inst = 32'hc404aae;
      26709: inst = 32'h8220000;
      26710: inst = 32'h10408000;
      26711: inst = 32'hc404aaf;
      26712: inst = 32'h8220000;
      26713: inst = 32'h10408000;
      26714: inst = 32'hc404ab0;
      26715: inst = 32'h8220000;
      26716: inst = 32'h10408000;
      26717: inst = 32'hc404ab1;
      26718: inst = 32'h8220000;
      26719: inst = 32'h10408000;
      26720: inst = 32'hc404ab2;
      26721: inst = 32'h8220000;
      26722: inst = 32'h10408000;
      26723: inst = 32'hc404ab3;
      26724: inst = 32'h8220000;
      26725: inst = 32'h10408000;
      26726: inst = 32'hc404ab4;
      26727: inst = 32'h8220000;
      26728: inst = 32'h10408000;
      26729: inst = 32'hc404ab5;
      26730: inst = 32'h8220000;
      26731: inst = 32'h10408000;
      26732: inst = 32'hc404ab6;
      26733: inst = 32'h8220000;
      26734: inst = 32'h10408000;
      26735: inst = 32'hc404ab7;
      26736: inst = 32'h8220000;
      26737: inst = 32'h10408000;
      26738: inst = 32'hc404ab8;
      26739: inst = 32'h8220000;
      26740: inst = 32'h10408000;
      26741: inst = 32'hc404ac7;
      26742: inst = 32'h8220000;
      26743: inst = 32'h10408000;
      26744: inst = 32'hc404ac8;
      26745: inst = 32'h8220000;
      26746: inst = 32'h10408000;
      26747: inst = 32'hc404ac9;
      26748: inst = 32'h8220000;
      26749: inst = 32'h10408000;
      26750: inst = 32'hc404aca;
      26751: inst = 32'h8220000;
      26752: inst = 32'h10408000;
      26753: inst = 32'hc404acb;
      26754: inst = 32'h8220000;
      26755: inst = 32'h10408000;
      26756: inst = 32'hc404acc;
      26757: inst = 32'h8220000;
      26758: inst = 32'h10408000;
      26759: inst = 32'hc404acd;
      26760: inst = 32'h8220000;
      26761: inst = 32'h10408000;
      26762: inst = 32'hc404ace;
      26763: inst = 32'h8220000;
      26764: inst = 32'h10408000;
      26765: inst = 32'hc404acf;
      26766: inst = 32'h8220000;
      26767: inst = 32'h10408000;
      26768: inst = 32'hc404ad0;
      26769: inst = 32'h8220000;
      26770: inst = 32'h10408000;
      26771: inst = 32'hc404ad1;
      26772: inst = 32'h8220000;
      26773: inst = 32'h10408000;
      26774: inst = 32'hc404ad2;
      26775: inst = 32'h8220000;
      26776: inst = 32'h10408000;
      26777: inst = 32'hc404ad3;
      26778: inst = 32'h8220000;
      26779: inst = 32'h10408000;
      26780: inst = 32'hc404ad4;
      26781: inst = 32'h8220000;
      26782: inst = 32'h10408000;
      26783: inst = 32'hc404ad5;
      26784: inst = 32'h8220000;
      26785: inst = 32'h10408000;
      26786: inst = 32'hc404ad6;
      26787: inst = 32'h8220000;
      26788: inst = 32'h10408000;
      26789: inst = 32'hc404ad7;
      26790: inst = 32'h8220000;
      26791: inst = 32'h10408000;
      26792: inst = 32'hc404ad8;
      26793: inst = 32'h8220000;
      26794: inst = 32'h10408000;
      26795: inst = 32'hc404ad9;
      26796: inst = 32'h8220000;
      26797: inst = 32'h10408000;
      26798: inst = 32'hc404ada;
      26799: inst = 32'h8220000;
      26800: inst = 32'h10408000;
      26801: inst = 32'hc404adb;
      26802: inst = 32'h8220000;
      26803: inst = 32'h10408000;
      26804: inst = 32'hc404adc;
      26805: inst = 32'h8220000;
      26806: inst = 32'h10408000;
      26807: inst = 32'hc404add;
      26808: inst = 32'h8220000;
      26809: inst = 32'h10408000;
      26810: inst = 32'hc404ade;
      26811: inst = 32'h8220000;
      26812: inst = 32'h10408000;
      26813: inst = 32'hc404adf;
      26814: inst = 32'h8220000;
      26815: inst = 32'h10408000;
      26816: inst = 32'hc404ae0;
      26817: inst = 32'h8220000;
      26818: inst = 32'h10408000;
      26819: inst = 32'hc404ae1;
      26820: inst = 32'h8220000;
      26821: inst = 32'h10408000;
      26822: inst = 32'hc404ae2;
      26823: inst = 32'h8220000;
      26824: inst = 32'h10408000;
      26825: inst = 32'hc404ae3;
      26826: inst = 32'h8220000;
      26827: inst = 32'h10408000;
      26828: inst = 32'hc404ae4;
      26829: inst = 32'h8220000;
      26830: inst = 32'h10408000;
      26831: inst = 32'hc404ae5;
      26832: inst = 32'h8220000;
      26833: inst = 32'h10408000;
      26834: inst = 32'hc404ae6;
      26835: inst = 32'h8220000;
      26836: inst = 32'h10408000;
      26837: inst = 32'hc404ae7;
      26838: inst = 32'h8220000;
      26839: inst = 32'h10408000;
      26840: inst = 32'hc404ae8;
      26841: inst = 32'h8220000;
      26842: inst = 32'h10408000;
      26843: inst = 32'hc404ae9;
      26844: inst = 32'h8220000;
      26845: inst = 32'h10408000;
      26846: inst = 32'hc404aea;
      26847: inst = 32'h8220000;
      26848: inst = 32'h10408000;
      26849: inst = 32'hc404aeb;
      26850: inst = 32'h8220000;
      26851: inst = 32'h10408000;
      26852: inst = 32'hc404aec;
      26853: inst = 32'h8220000;
      26854: inst = 32'h10408000;
      26855: inst = 32'hc404aed;
      26856: inst = 32'h8220000;
      26857: inst = 32'h10408000;
      26858: inst = 32'hc404aee;
      26859: inst = 32'h8220000;
      26860: inst = 32'h10408000;
      26861: inst = 32'hc404aef;
      26862: inst = 32'h8220000;
      26863: inst = 32'h10408000;
      26864: inst = 32'hc404af0;
      26865: inst = 32'h8220000;
      26866: inst = 32'h10408000;
      26867: inst = 32'hc404af1;
      26868: inst = 32'h8220000;
      26869: inst = 32'h10408000;
      26870: inst = 32'hc404af2;
      26871: inst = 32'h8220000;
      26872: inst = 32'h10408000;
      26873: inst = 32'hc404af3;
      26874: inst = 32'h8220000;
      26875: inst = 32'h10408000;
      26876: inst = 32'hc404af4;
      26877: inst = 32'h8220000;
      26878: inst = 32'h10408000;
      26879: inst = 32'hc404af5;
      26880: inst = 32'h8220000;
      26881: inst = 32'h10408000;
      26882: inst = 32'hc404af6;
      26883: inst = 32'h8220000;
      26884: inst = 32'h10408000;
      26885: inst = 32'hc404af7;
      26886: inst = 32'h8220000;
      26887: inst = 32'h10408000;
      26888: inst = 32'hc404af8;
      26889: inst = 32'h8220000;
      26890: inst = 32'h10408000;
      26891: inst = 32'hc404af9;
      26892: inst = 32'h8220000;
      26893: inst = 32'h10408000;
      26894: inst = 32'hc404afa;
      26895: inst = 32'h8220000;
      26896: inst = 32'h10408000;
      26897: inst = 32'hc404afb;
      26898: inst = 32'h8220000;
      26899: inst = 32'h10408000;
      26900: inst = 32'hc404afc;
      26901: inst = 32'h8220000;
      26902: inst = 32'h10408000;
      26903: inst = 32'hc404afd;
      26904: inst = 32'h8220000;
      26905: inst = 32'h10408000;
      26906: inst = 32'hc404afe;
      26907: inst = 32'h8220000;
      26908: inst = 32'h10408000;
      26909: inst = 32'hc404aff;
      26910: inst = 32'h8220000;
      26911: inst = 32'h10408000;
      26912: inst = 32'hc404b00;
      26913: inst = 32'h8220000;
      26914: inst = 32'h10408000;
      26915: inst = 32'hc404b01;
      26916: inst = 32'h8220000;
      26917: inst = 32'h10408000;
      26918: inst = 32'hc404b02;
      26919: inst = 32'h8220000;
      26920: inst = 32'h10408000;
      26921: inst = 32'hc404b03;
      26922: inst = 32'h8220000;
      26923: inst = 32'h10408000;
      26924: inst = 32'hc404b04;
      26925: inst = 32'h8220000;
      26926: inst = 32'h10408000;
      26927: inst = 32'hc404b05;
      26928: inst = 32'h8220000;
      26929: inst = 32'h10408000;
      26930: inst = 32'hc404b06;
      26931: inst = 32'h8220000;
      26932: inst = 32'h10408000;
      26933: inst = 32'hc404b07;
      26934: inst = 32'h8220000;
      26935: inst = 32'h10408000;
      26936: inst = 32'hc404b08;
      26937: inst = 32'h8220000;
      26938: inst = 32'h10408000;
      26939: inst = 32'hc404b09;
      26940: inst = 32'h8220000;
      26941: inst = 32'h10408000;
      26942: inst = 32'hc404b0a;
      26943: inst = 32'h8220000;
      26944: inst = 32'h10408000;
      26945: inst = 32'hc404b0b;
      26946: inst = 32'h8220000;
      26947: inst = 32'h10408000;
      26948: inst = 32'hc404b0c;
      26949: inst = 32'h8220000;
      26950: inst = 32'h10408000;
      26951: inst = 32'hc404b0d;
      26952: inst = 32'h8220000;
      26953: inst = 32'h10408000;
      26954: inst = 32'hc404b0e;
      26955: inst = 32'h8220000;
      26956: inst = 32'h10408000;
      26957: inst = 32'hc404b0f;
      26958: inst = 32'h8220000;
      26959: inst = 32'h10408000;
      26960: inst = 32'hc404b10;
      26961: inst = 32'h8220000;
      26962: inst = 32'h10408000;
      26963: inst = 32'hc404b11;
      26964: inst = 32'h8220000;
      26965: inst = 32'h10408000;
      26966: inst = 32'hc404b12;
      26967: inst = 32'h8220000;
      26968: inst = 32'h10408000;
      26969: inst = 32'hc404b13;
      26970: inst = 32'h8220000;
      26971: inst = 32'h10408000;
      26972: inst = 32'hc404b14;
      26973: inst = 32'h8220000;
      26974: inst = 32'h10408000;
      26975: inst = 32'hc404b15;
      26976: inst = 32'h8220000;
      26977: inst = 32'h10408000;
      26978: inst = 32'hc404b16;
      26979: inst = 32'h8220000;
      26980: inst = 32'h10408000;
      26981: inst = 32'hc404b17;
      26982: inst = 32'h8220000;
      26983: inst = 32'h10408000;
      26984: inst = 32'hc404b18;
      26985: inst = 32'h8220000;
      26986: inst = 32'h10408000;
      26987: inst = 32'hc404b27;
      26988: inst = 32'h8220000;
      26989: inst = 32'h10408000;
      26990: inst = 32'hc404b28;
      26991: inst = 32'h8220000;
      26992: inst = 32'h10408000;
      26993: inst = 32'hc404b29;
      26994: inst = 32'h8220000;
      26995: inst = 32'h10408000;
      26996: inst = 32'hc404b2a;
      26997: inst = 32'h8220000;
      26998: inst = 32'h10408000;
      26999: inst = 32'hc404b2b;
      27000: inst = 32'h8220000;
      27001: inst = 32'h10408000;
      27002: inst = 32'hc404b2c;
      27003: inst = 32'h8220000;
      27004: inst = 32'h10408000;
      27005: inst = 32'hc404b2d;
      27006: inst = 32'h8220000;
      27007: inst = 32'h10408000;
      27008: inst = 32'hc404b2e;
      27009: inst = 32'h8220000;
      27010: inst = 32'h10408000;
      27011: inst = 32'hc404b2f;
      27012: inst = 32'h8220000;
      27013: inst = 32'h10408000;
      27014: inst = 32'hc404b30;
      27015: inst = 32'h8220000;
      27016: inst = 32'h10408000;
      27017: inst = 32'hc404b31;
      27018: inst = 32'h8220000;
      27019: inst = 32'h10408000;
      27020: inst = 32'hc404b32;
      27021: inst = 32'h8220000;
      27022: inst = 32'h10408000;
      27023: inst = 32'hc404b33;
      27024: inst = 32'h8220000;
      27025: inst = 32'h10408000;
      27026: inst = 32'hc404b34;
      27027: inst = 32'h8220000;
      27028: inst = 32'h10408000;
      27029: inst = 32'hc404b35;
      27030: inst = 32'h8220000;
      27031: inst = 32'h10408000;
      27032: inst = 32'hc404b36;
      27033: inst = 32'h8220000;
      27034: inst = 32'h10408000;
      27035: inst = 32'hc404b37;
      27036: inst = 32'h8220000;
      27037: inst = 32'h10408000;
      27038: inst = 32'hc404b38;
      27039: inst = 32'h8220000;
      27040: inst = 32'h10408000;
      27041: inst = 32'hc404b39;
      27042: inst = 32'h8220000;
      27043: inst = 32'h10408000;
      27044: inst = 32'hc404b3a;
      27045: inst = 32'h8220000;
      27046: inst = 32'h10408000;
      27047: inst = 32'hc404b3b;
      27048: inst = 32'h8220000;
      27049: inst = 32'h10408000;
      27050: inst = 32'hc404b3c;
      27051: inst = 32'h8220000;
      27052: inst = 32'h10408000;
      27053: inst = 32'hc404b3d;
      27054: inst = 32'h8220000;
      27055: inst = 32'h10408000;
      27056: inst = 32'hc404b3e;
      27057: inst = 32'h8220000;
      27058: inst = 32'h10408000;
      27059: inst = 32'hc404b3f;
      27060: inst = 32'h8220000;
      27061: inst = 32'h10408000;
      27062: inst = 32'hc404b40;
      27063: inst = 32'h8220000;
      27064: inst = 32'h10408000;
      27065: inst = 32'hc404b41;
      27066: inst = 32'h8220000;
      27067: inst = 32'h10408000;
      27068: inst = 32'hc404b42;
      27069: inst = 32'h8220000;
      27070: inst = 32'h10408000;
      27071: inst = 32'hc404b43;
      27072: inst = 32'h8220000;
      27073: inst = 32'h10408000;
      27074: inst = 32'hc404b44;
      27075: inst = 32'h8220000;
      27076: inst = 32'h10408000;
      27077: inst = 32'hc404b45;
      27078: inst = 32'h8220000;
      27079: inst = 32'h10408000;
      27080: inst = 32'hc404b46;
      27081: inst = 32'h8220000;
      27082: inst = 32'h10408000;
      27083: inst = 32'hc404b47;
      27084: inst = 32'h8220000;
      27085: inst = 32'h10408000;
      27086: inst = 32'hc404b48;
      27087: inst = 32'h8220000;
      27088: inst = 32'h10408000;
      27089: inst = 32'hc404b49;
      27090: inst = 32'h8220000;
      27091: inst = 32'h10408000;
      27092: inst = 32'hc404b4a;
      27093: inst = 32'h8220000;
      27094: inst = 32'h10408000;
      27095: inst = 32'hc404b4b;
      27096: inst = 32'h8220000;
      27097: inst = 32'h10408000;
      27098: inst = 32'hc404b4c;
      27099: inst = 32'h8220000;
      27100: inst = 32'h10408000;
      27101: inst = 32'hc404b4d;
      27102: inst = 32'h8220000;
      27103: inst = 32'h10408000;
      27104: inst = 32'hc404b4e;
      27105: inst = 32'h8220000;
      27106: inst = 32'h10408000;
      27107: inst = 32'hc404b4f;
      27108: inst = 32'h8220000;
      27109: inst = 32'h10408000;
      27110: inst = 32'hc404b50;
      27111: inst = 32'h8220000;
      27112: inst = 32'h10408000;
      27113: inst = 32'hc404b51;
      27114: inst = 32'h8220000;
      27115: inst = 32'h10408000;
      27116: inst = 32'hc404b52;
      27117: inst = 32'h8220000;
      27118: inst = 32'h10408000;
      27119: inst = 32'hc404b53;
      27120: inst = 32'h8220000;
      27121: inst = 32'h10408000;
      27122: inst = 32'hc404b54;
      27123: inst = 32'h8220000;
      27124: inst = 32'h10408000;
      27125: inst = 32'hc404b55;
      27126: inst = 32'h8220000;
      27127: inst = 32'h10408000;
      27128: inst = 32'hc404b56;
      27129: inst = 32'h8220000;
      27130: inst = 32'h10408000;
      27131: inst = 32'hc404b57;
      27132: inst = 32'h8220000;
      27133: inst = 32'h10408000;
      27134: inst = 32'hc404b58;
      27135: inst = 32'h8220000;
      27136: inst = 32'h10408000;
      27137: inst = 32'hc404b59;
      27138: inst = 32'h8220000;
      27139: inst = 32'h10408000;
      27140: inst = 32'hc404b5a;
      27141: inst = 32'h8220000;
      27142: inst = 32'h10408000;
      27143: inst = 32'hc404b5b;
      27144: inst = 32'h8220000;
      27145: inst = 32'h10408000;
      27146: inst = 32'hc404b5c;
      27147: inst = 32'h8220000;
      27148: inst = 32'h10408000;
      27149: inst = 32'hc404b5d;
      27150: inst = 32'h8220000;
      27151: inst = 32'h10408000;
      27152: inst = 32'hc404b5e;
      27153: inst = 32'h8220000;
      27154: inst = 32'h10408000;
      27155: inst = 32'hc404b5f;
      27156: inst = 32'h8220000;
      27157: inst = 32'h10408000;
      27158: inst = 32'hc404b60;
      27159: inst = 32'h8220000;
      27160: inst = 32'h10408000;
      27161: inst = 32'hc404b61;
      27162: inst = 32'h8220000;
      27163: inst = 32'h10408000;
      27164: inst = 32'hc404b62;
      27165: inst = 32'h8220000;
      27166: inst = 32'h10408000;
      27167: inst = 32'hc404b63;
      27168: inst = 32'h8220000;
      27169: inst = 32'h10408000;
      27170: inst = 32'hc404b64;
      27171: inst = 32'h8220000;
      27172: inst = 32'h10408000;
      27173: inst = 32'hc404b65;
      27174: inst = 32'h8220000;
      27175: inst = 32'h10408000;
      27176: inst = 32'hc404b66;
      27177: inst = 32'h8220000;
      27178: inst = 32'h10408000;
      27179: inst = 32'hc404b67;
      27180: inst = 32'h8220000;
      27181: inst = 32'h10408000;
      27182: inst = 32'hc404b68;
      27183: inst = 32'h8220000;
      27184: inst = 32'h10408000;
      27185: inst = 32'hc404b69;
      27186: inst = 32'h8220000;
      27187: inst = 32'h10408000;
      27188: inst = 32'hc404b6a;
      27189: inst = 32'h8220000;
      27190: inst = 32'h10408000;
      27191: inst = 32'hc404b6b;
      27192: inst = 32'h8220000;
      27193: inst = 32'h10408000;
      27194: inst = 32'hc404b6c;
      27195: inst = 32'h8220000;
      27196: inst = 32'h10408000;
      27197: inst = 32'hc404b6d;
      27198: inst = 32'h8220000;
      27199: inst = 32'h10408000;
      27200: inst = 32'hc404b6e;
      27201: inst = 32'h8220000;
      27202: inst = 32'h10408000;
      27203: inst = 32'hc404b6f;
      27204: inst = 32'h8220000;
      27205: inst = 32'h10408000;
      27206: inst = 32'hc404b70;
      27207: inst = 32'h8220000;
      27208: inst = 32'h10408000;
      27209: inst = 32'hc404b71;
      27210: inst = 32'h8220000;
      27211: inst = 32'h10408000;
      27212: inst = 32'hc404b72;
      27213: inst = 32'h8220000;
      27214: inst = 32'h10408000;
      27215: inst = 32'hc404b73;
      27216: inst = 32'h8220000;
      27217: inst = 32'h10408000;
      27218: inst = 32'hc404b74;
      27219: inst = 32'h8220000;
      27220: inst = 32'h10408000;
      27221: inst = 32'hc404b75;
      27222: inst = 32'h8220000;
      27223: inst = 32'h10408000;
      27224: inst = 32'hc404b76;
      27225: inst = 32'h8220000;
      27226: inst = 32'h10408000;
      27227: inst = 32'hc404b77;
      27228: inst = 32'h8220000;
      27229: inst = 32'h10408000;
      27230: inst = 32'hc404b78;
      27231: inst = 32'h8220000;
      27232: inst = 32'h10408000;
      27233: inst = 32'hc404b87;
      27234: inst = 32'h8220000;
      27235: inst = 32'h10408000;
      27236: inst = 32'hc404b88;
      27237: inst = 32'h8220000;
      27238: inst = 32'h10408000;
      27239: inst = 32'hc404b89;
      27240: inst = 32'h8220000;
      27241: inst = 32'h10408000;
      27242: inst = 32'hc404b8a;
      27243: inst = 32'h8220000;
      27244: inst = 32'h10408000;
      27245: inst = 32'hc404b8b;
      27246: inst = 32'h8220000;
      27247: inst = 32'h10408000;
      27248: inst = 32'hc404b8c;
      27249: inst = 32'h8220000;
      27250: inst = 32'h10408000;
      27251: inst = 32'hc404b8d;
      27252: inst = 32'h8220000;
      27253: inst = 32'h10408000;
      27254: inst = 32'hc404b8e;
      27255: inst = 32'h8220000;
      27256: inst = 32'h10408000;
      27257: inst = 32'hc404b8f;
      27258: inst = 32'h8220000;
      27259: inst = 32'h10408000;
      27260: inst = 32'hc404b90;
      27261: inst = 32'h8220000;
      27262: inst = 32'h10408000;
      27263: inst = 32'hc404b91;
      27264: inst = 32'h8220000;
      27265: inst = 32'h10408000;
      27266: inst = 32'hc404b92;
      27267: inst = 32'h8220000;
      27268: inst = 32'h10408000;
      27269: inst = 32'hc404b93;
      27270: inst = 32'h8220000;
      27271: inst = 32'h10408000;
      27272: inst = 32'hc404b94;
      27273: inst = 32'h8220000;
      27274: inst = 32'h10408000;
      27275: inst = 32'hc404b95;
      27276: inst = 32'h8220000;
      27277: inst = 32'h10408000;
      27278: inst = 32'hc404b96;
      27279: inst = 32'h8220000;
      27280: inst = 32'h10408000;
      27281: inst = 32'hc404b97;
      27282: inst = 32'h8220000;
      27283: inst = 32'h10408000;
      27284: inst = 32'hc404b98;
      27285: inst = 32'h8220000;
      27286: inst = 32'h10408000;
      27287: inst = 32'hc404b99;
      27288: inst = 32'h8220000;
      27289: inst = 32'h10408000;
      27290: inst = 32'hc404b9a;
      27291: inst = 32'h8220000;
      27292: inst = 32'h10408000;
      27293: inst = 32'hc404b9b;
      27294: inst = 32'h8220000;
      27295: inst = 32'h10408000;
      27296: inst = 32'hc404b9c;
      27297: inst = 32'h8220000;
      27298: inst = 32'h10408000;
      27299: inst = 32'hc404b9d;
      27300: inst = 32'h8220000;
      27301: inst = 32'h10408000;
      27302: inst = 32'hc404b9e;
      27303: inst = 32'h8220000;
      27304: inst = 32'h10408000;
      27305: inst = 32'hc404b9f;
      27306: inst = 32'h8220000;
      27307: inst = 32'h10408000;
      27308: inst = 32'hc404ba0;
      27309: inst = 32'h8220000;
      27310: inst = 32'h10408000;
      27311: inst = 32'hc404ba1;
      27312: inst = 32'h8220000;
      27313: inst = 32'h10408000;
      27314: inst = 32'hc404ba2;
      27315: inst = 32'h8220000;
      27316: inst = 32'h10408000;
      27317: inst = 32'hc404ba3;
      27318: inst = 32'h8220000;
      27319: inst = 32'h10408000;
      27320: inst = 32'hc404ba4;
      27321: inst = 32'h8220000;
      27322: inst = 32'h10408000;
      27323: inst = 32'hc404ba5;
      27324: inst = 32'h8220000;
      27325: inst = 32'h10408000;
      27326: inst = 32'hc404ba6;
      27327: inst = 32'h8220000;
      27328: inst = 32'h10408000;
      27329: inst = 32'hc404ba7;
      27330: inst = 32'h8220000;
      27331: inst = 32'h10408000;
      27332: inst = 32'hc404ba8;
      27333: inst = 32'h8220000;
      27334: inst = 32'h10408000;
      27335: inst = 32'hc404ba9;
      27336: inst = 32'h8220000;
      27337: inst = 32'h10408000;
      27338: inst = 32'hc404baa;
      27339: inst = 32'h8220000;
      27340: inst = 32'h10408000;
      27341: inst = 32'hc404bab;
      27342: inst = 32'h8220000;
      27343: inst = 32'h10408000;
      27344: inst = 32'hc404bac;
      27345: inst = 32'h8220000;
      27346: inst = 32'h10408000;
      27347: inst = 32'hc404bad;
      27348: inst = 32'h8220000;
      27349: inst = 32'h10408000;
      27350: inst = 32'hc404bae;
      27351: inst = 32'h8220000;
      27352: inst = 32'h10408000;
      27353: inst = 32'hc404baf;
      27354: inst = 32'h8220000;
      27355: inst = 32'h10408000;
      27356: inst = 32'hc404bb0;
      27357: inst = 32'h8220000;
      27358: inst = 32'h10408000;
      27359: inst = 32'hc404bb1;
      27360: inst = 32'h8220000;
      27361: inst = 32'h10408000;
      27362: inst = 32'hc404bb2;
      27363: inst = 32'h8220000;
      27364: inst = 32'h10408000;
      27365: inst = 32'hc404bb3;
      27366: inst = 32'h8220000;
      27367: inst = 32'h10408000;
      27368: inst = 32'hc404bb4;
      27369: inst = 32'h8220000;
      27370: inst = 32'h10408000;
      27371: inst = 32'hc404bb5;
      27372: inst = 32'h8220000;
      27373: inst = 32'h10408000;
      27374: inst = 32'hc404bb6;
      27375: inst = 32'h8220000;
      27376: inst = 32'h10408000;
      27377: inst = 32'hc404bb7;
      27378: inst = 32'h8220000;
      27379: inst = 32'h10408000;
      27380: inst = 32'hc404bb8;
      27381: inst = 32'h8220000;
      27382: inst = 32'h10408000;
      27383: inst = 32'hc404bb9;
      27384: inst = 32'h8220000;
      27385: inst = 32'h10408000;
      27386: inst = 32'hc404bba;
      27387: inst = 32'h8220000;
      27388: inst = 32'h10408000;
      27389: inst = 32'hc404bbb;
      27390: inst = 32'h8220000;
      27391: inst = 32'h10408000;
      27392: inst = 32'hc404bbc;
      27393: inst = 32'h8220000;
      27394: inst = 32'h10408000;
      27395: inst = 32'hc404bbd;
      27396: inst = 32'h8220000;
      27397: inst = 32'h10408000;
      27398: inst = 32'hc404bbe;
      27399: inst = 32'h8220000;
      27400: inst = 32'h10408000;
      27401: inst = 32'hc404bbf;
      27402: inst = 32'h8220000;
      27403: inst = 32'h10408000;
      27404: inst = 32'hc404bc0;
      27405: inst = 32'h8220000;
      27406: inst = 32'h10408000;
      27407: inst = 32'hc404bc1;
      27408: inst = 32'h8220000;
      27409: inst = 32'h10408000;
      27410: inst = 32'hc404bc2;
      27411: inst = 32'h8220000;
      27412: inst = 32'h10408000;
      27413: inst = 32'hc404bc3;
      27414: inst = 32'h8220000;
      27415: inst = 32'h10408000;
      27416: inst = 32'hc404bc4;
      27417: inst = 32'h8220000;
      27418: inst = 32'h10408000;
      27419: inst = 32'hc404bc5;
      27420: inst = 32'h8220000;
      27421: inst = 32'h10408000;
      27422: inst = 32'hc404bc6;
      27423: inst = 32'h8220000;
      27424: inst = 32'h10408000;
      27425: inst = 32'hc404bc7;
      27426: inst = 32'h8220000;
      27427: inst = 32'h10408000;
      27428: inst = 32'hc404bc8;
      27429: inst = 32'h8220000;
      27430: inst = 32'h10408000;
      27431: inst = 32'hc404bc9;
      27432: inst = 32'h8220000;
      27433: inst = 32'h10408000;
      27434: inst = 32'hc404bca;
      27435: inst = 32'h8220000;
      27436: inst = 32'h10408000;
      27437: inst = 32'hc404bcb;
      27438: inst = 32'h8220000;
      27439: inst = 32'h10408000;
      27440: inst = 32'hc404bcc;
      27441: inst = 32'h8220000;
      27442: inst = 32'h10408000;
      27443: inst = 32'hc404bcd;
      27444: inst = 32'h8220000;
      27445: inst = 32'h10408000;
      27446: inst = 32'hc404bce;
      27447: inst = 32'h8220000;
      27448: inst = 32'h10408000;
      27449: inst = 32'hc404bcf;
      27450: inst = 32'h8220000;
      27451: inst = 32'h10408000;
      27452: inst = 32'hc404bd0;
      27453: inst = 32'h8220000;
      27454: inst = 32'h10408000;
      27455: inst = 32'hc404bd1;
      27456: inst = 32'h8220000;
      27457: inst = 32'h10408000;
      27458: inst = 32'hc404bd2;
      27459: inst = 32'h8220000;
      27460: inst = 32'h10408000;
      27461: inst = 32'hc404bd3;
      27462: inst = 32'h8220000;
      27463: inst = 32'h10408000;
      27464: inst = 32'hc404bd4;
      27465: inst = 32'h8220000;
      27466: inst = 32'h10408000;
      27467: inst = 32'hc404bd5;
      27468: inst = 32'h8220000;
      27469: inst = 32'h10408000;
      27470: inst = 32'hc404bd6;
      27471: inst = 32'h8220000;
      27472: inst = 32'h10408000;
      27473: inst = 32'hc404bd7;
      27474: inst = 32'h8220000;
      27475: inst = 32'h10408000;
      27476: inst = 32'hc404bd8;
      27477: inst = 32'h8220000;
      27478: inst = 32'h10408000;
      27479: inst = 32'hc404be7;
      27480: inst = 32'h8220000;
      27481: inst = 32'h10408000;
      27482: inst = 32'hc404be8;
      27483: inst = 32'h8220000;
      27484: inst = 32'h10408000;
      27485: inst = 32'hc404be9;
      27486: inst = 32'h8220000;
      27487: inst = 32'h10408000;
      27488: inst = 32'hc404bea;
      27489: inst = 32'h8220000;
      27490: inst = 32'h10408000;
      27491: inst = 32'hc404beb;
      27492: inst = 32'h8220000;
      27493: inst = 32'h10408000;
      27494: inst = 32'hc404bec;
      27495: inst = 32'h8220000;
      27496: inst = 32'h10408000;
      27497: inst = 32'hc404bed;
      27498: inst = 32'h8220000;
      27499: inst = 32'h10408000;
      27500: inst = 32'hc404bee;
      27501: inst = 32'h8220000;
      27502: inst = 32'h10408000;
      27503: inst = 32'hc404bef;
      27504: inst = 32'h8220000;
      27505: inst = 32'h10408000;
      27506: inst = 32'hc404bf0;
      27507: inst = 32'h8220000;
      27508: inst = 32'h10408000;
      27509: inst = 32'hc404bf1;
      27510: inst = 32'h8220000;
      27511: inst = 32'h10408000;
      27512: inst = 32'hc404bf2;
      27513: inst = 32'h8220000;
      27514: inst = 32'h10408000;
      27515: inst = 32'hc404bf3;
      27516: inst = 32'h8220000;
      27517: inst = 32'h10408000;
      27518: inst = 32'hc404bf4;
      27519: inst = 32'h8220000;
      27520: inst = 32'h10408000;
      27521: inst = 32'hc404bf5;
      27522: inst = 32'h8220000;
      27523: inst = 32'h10408000;
      27524: inst = 32'hc404bf6;
      27525: inst = 32'h8220000;
      27526: inst = 32'h10408000;
      27527: inst = 32'hc404bf7;
      27528: inst = 32'h8220000;
      27529: inst = 32'h10408000;
      27530: inst = 32'hc404bf8;
      27531: inst = 32'h8220000;
      27532: inst = 32'h10408000;
      27533: inst = 32'hc404bf9;
      27534: inst = 32'h8220000;
      27535: inst = 32'h10408000;
      27536: inst = 32'hc404bfa;
      27537: inst = 32'h8220000;
      27538: inst = 32'h10408000;
      27539: inst = 32'hc404bfb;
      27540: inst = 32'h8220000;
      27541: inst = 32'h10408000;
      27542: inst = 32'hc404bfc;
      27543: inst = 32'h8220000;
      27544: inst = 32'h10408000;
      27545: inst = 32'hc404bfd;
      27546: inst = 32'h8220000;
      27547: inst = 32'h10408000;
      27548: inst = 32'hc404bfe;
      27549: inst = 32'h8220000;
      27550: inst = 32'h10408000;
      27551: inst = 32'hc404bff;
      27552: inst = 32'h8220000;
      27553: inst = 32'h10408000;
      27554: inst = 32'hc404c00;
      27555: inst = 32'h8220000;
      27556: inst = 32'h10408000;
      27557: inst = 32'hc404c01;
      27558: inst = 32'h8220000;
      27559: inst = 32'h10408000;
      27560: inst = 32'hc404c02;
      27561: inst = 32'h8220000;
      27562: inst = 32'h10408000;
      27563: inst = 32'hc404c03;
      27564: inst = 32'h8220000;
      27565: inst = 32'h10408000;
      27566: inst = 32'hc404c04;
      27567: inst = 32'h8220000;
      27568: inst = 32'h10408000;
      27569: inst = 32'hc404c05;
      27570: inst = 32'h8220000;
      27571: inst = 32'h10408000;
      27572: inst = 32'hc404c06;
      27573: inst = 32'h8220000;
      27574: inst = 32'h10408000;
      27575: inst = 32'hc404c07;
      27576: inst = 32'h8220000;
      27577: inst = 32'h10408000;
      27578: inst = 32'hc404c08;
      27579: inst = 32'h8220000;
      27580: inst = 32'h10408000;
      27581: inst = 32'hc404c09;
      27582: inst = 32'h8220000;
      27583: inst = 32'h10408000;
      27584: inst = 32'hc404c0a;
      27585: inst = 32'h8220000;
      27586: inst = 32'h10408000;
      27587: inst = 32'hc404c0b;
      27588: inst = 32'h8220000;
      27589: inst = 32'h10408000;
      27590: inst = 32'hc404c0c;
      27591: inst = 32'h8220000;
      27592: inst = 32'h10408000;
      27593: inst = 32'hc404c0d;
      27594: inst = 32'h8220000;
      27595: inst = 32'h10408000;
      27596: inst = 32'hc404c0e;
      27597: inst = 32'h8220000;
      27598: inst = 32'h10408000;
      27599: inst = 32'hc404c0f;
      27600: inst = 32'h8220000;
      27601: inst = 32'h10408000;
      27602: inst = 32'hc404c10;
      27603: inst = 32'h8220000;
      27604: inst = 32'h10408000;
      27605: inst = 32'hc404c11;
      27606: inst = 32'h8220000;
      27607: inst = 32'h10408000;
      27608: inst = 32'hc404c12;
      27609: inst = 32'h8220000;
      27610: inst = 32'h10408000;
      27611: inst = 32'hc404c13;
      27612: inst = 32'h8220000;
      27613: inst = 32'h10408000;
      27614: inst = 32'hc404c14;
      27615: inst = 32'h8220000;
      27616: inst = 32'h10408000;
      27617: inst = 32'hc404c15;
      27618: inst = 32'h8220000;
      27619: inst = 32'h10408000;
      27620: inst = 32'hc404c16;
      27621: inst = 32'h8220000;
      27622: inst = 32'h10408000;
      27623: inst = 32'hc404c17;
      27624: inst = 32'h8220000;
      27625: inst = 32'h10408000;
      27626: inst = 32'hc404c18;
      27627: inst = 32'h8220000;
      27628: inst = 32'h10408000;
      27629: inst = 32'hc404c19;
      27630: inst = 32'h8220000;
      27631: inst = 32'h10408000;
      27632: inst = 32'hc404c1a;
      27633: inst = 32'h8220000;
      27634: inst = 32'h10408000;
      27635: inst = 32'hc404c1b;
      27636: inst = 32'h8220000;
      27637: inst = 32'h10408000;
      27638: inst = 32'hc404c1c;
      27639: inst = 32'h8220000;
      27640: inst = 32'h10408000;
      27641: inst = 32'hc404c1d;
      27642: inst = 32'h8220000;
      27643: inst = 32'h10408000;
      27644: inst = 32'hc404c1e;
      27645: inst = 32'h8220000;
      27646: inst = 32'h10408000;
      27647: inst = 32'hc404c1f;
      27648: inst = 32'h8220000;
      27649: inst = 32'h10408000;
      27650: inst = 32'hc404c20;
      27651: inst = 32'h8220000;
      27652: inst = 32'h10408000;
      27653: inst = 32'hc404c21;
      27654: inst = 32'h8220000;
      27655: inst = 32'h10408000;
      27656: inst = 32'hc404c22;
      27657: inst = 32'h8220000;
      27658: inst = 32'h10408000;
      27659: inst = 32'hc404c23;
      27660: inst = 32'h8220000;
      27661: inst = 32'h10408000;
      27662: inst = 32'hc404c24;
      27663: inst = 32'h8220000;
      27664: inst = 32'h10408000;
      27665: inst = 32'hc404c25;
      27666: inst = 32'h8220000;
      27667: inst = 32'h10408000;
      27668: inst = 32'hc404c26;
      27669: inst = 32'h8220000;
      27670: inst = 32'h10408000;
      27671: inst = 32'hc404c27;
      27672: inst = 32'h8220000;
      27673: inst = 32'h10408000;
      27674: inst = 32'hc404c28;
      27675: inst = 32'h8220000;
      27676: inst = 32'h10408000;
      27677: inst = 32'hc404c29;
      27678: inst = 32'h8220000;
      27679: inst = 32'h10408000;
      27680: inst = 32'hc404c2a;
      27681: inst = 32'h8220000;
      27682: inst = 32'h10408000;
      27683: inst = 32'hc404c2b;
      27684: inst = 32'h8220000;
      27685: inst = 32'h10408000;
      27686: inst = 32'hc404c2c;
      27687: inst = 32'h8220000;
      27688: inst = 32'h10408000;
      27689: inst = 32'hc404c2d;
      27690: inst = 32'h8220000;
      27691: inst = 32'h10408000;
      27692: inst = 32'hc404c2e;
      27693: inst = 32'h8220000;
      27694: inst = 32'h10408000;
      27695: inst = 32'hc404c2f;
      27696: inst = 32'h8220000;
      27697: inst = 32'h10408000;
      27698: inst = 32'hc404c30;
      27699: inst = 32'h8220000;
      27700: inst = 32'h10408000;
      27701: inst = 32'hc404c31;
      27702: inst = 32'h8220000;
      27703: inst = 32'h10408000;
      27704: inst = 32'hc404c32;
      27705: inst = 32'h8220000;
      27706: inst = 32'h10408000;
      27707: inst = 32'hc404c33;
      27708: inst = 32'h8220000;
      27709: inst = 32'h10408000;
      27710: inst = 32'hc404c34;
      27711: inst = 32'h8220000;
      27712: inst = 32'h10408000;
      27713: inst = 32'hc404c35;
      27714: inst = 32'h8220000;
      27715: inst = 32'h10408000;
      27716: inst = 32'hc404c36;
      27717: inst = 32'h8220000;
      27718: inst = 32'h10408000;
      27719: inst = 32'hc404c37;
      27720: inst = 32'h8220000;
      27721: inst = 32'h10408000;
      27722: inst = 32'hc404c38;
      27723: inst = 32'h8220000;
      27724: inst = 32'h10408000;
      27725: inst = 32'hc404c47;
      27726: inst = 32'h8220000;
      27727: inst = 32'h10408000;
      27728: inst = 32'hc404c48;
      27729: inst = 32'h8220000;
      27730: inst = 32'h10408000;
      27731: inst = 32'hc404c49;
      27732: inst = 32'h8220000;
      27733: inst = 32'h10408000;
      27734: inst = 32'hc404c4a;
      27735: inst = 32'h8220000;
      27736: inst = 32'h10408000;
      27737: inst = 32'hc404c4b;
      27738: inst = 32'h8220000;
      27739: inst = 32'h10408000;
      27740: inst = 32'hc404c4c;
      27741: inst = 32'h8220000;
      27742: inst = 32'h10408000;
      27743: inst = 32'hc404c4d;
      27744: inst = 32'h8220000;
      27745: inst = 32'h10408000;
      27746: inst = 32'hc404c4e;
      27747: inst = 32'h8220000;
      27748: inst = 32'h10408000;
      27749: inst = 32'hc404c4f;
      27750: inst = 32'h8220000;
      27751: inst = 32'h10408000;
      27752: inst = 32'hc404c50;
      27753: inst = 32'h8220000;
      27754: inst = 32'h10408000;
      27755: inst = 32'hc404c51;
      27756: inst = 32'h8220000;
      27757: inst = 32'h10408000;
      27758: inst = 32'hc404c52;
      27759: inst = 32'h8220000;
      27760: inst = 32'h10408000;
      27761: inst = 32'hc404c53;
      27762: inst = 32'h8220000;
      27763: inst = 32'h10408000;
      27764: inst = 32'hc404c54;
      27765: inst = 32'h8220000;
      27766: inst = 32'h10408000;
      27767: inst = 32'hc404c55;
      27768: inst = 32'h8220000;
      27769: inst = 32'h10408000;
      27770: inst = 32'hc404c56;
      27771: inst = 32'h8220000;
      27772: inst = 32'h10408000;
      27773: inst = 32'hc404c57;
      27774: inst = 32'h8220000;
      27775: inst = 32'h10408000;
      27776: inst = 32'hc404c58;
      27777: inst = 32'h8220000;
      27778: inst = 32'h10408000;
      27779: inst = 32'hc404c59;
      27780: inst = 32'h8220000;
      27781: inst = 32'h10408000;
      27782: inst = 32'hc404c5a;
      27783: inst = 32'h8220000;
      27784: inst = 32'h10408000;
      27785: inst = 32'hc404c5b;
      27786: inst = 32'h8220000;
      27787: inst = 32'h10408000;
      27788: inst = 32'hc404c5c;
      27789: inst = 32'h8220000;
      27790: inst = 32'h10408000;
      27791: inst = 32'hc404c5d;
      27792: inst = 32'h8220000;
      27793: inst = 32'h10408000;
      27794: inst = 32'hc404c5e;
      27795: inst = 32'h8220000;
      27796: inst = 32'h10408000;
      27797: inst = 32'hc404c5f;
      27798: inst = 32'h8220000;
      27799: inst = 32'h10408000;
      27800: inst = 32'hc404c60;
      27801: inst = 32'h8220000;
      27802: inst = 32'h10408000;
      27803: inst = 32'hc404c61;
      27804: inst = 32'h8220000;
      27805: inst = 32'h10408000;
      27806: inst = 32'hc404c62;
      27807: inst = 32'h8220000;
      27808: inst = 32'h10408000;
      27809: inst = 32'hc404c63;
      27810: inst = 32'h8220000;
      27811: inst = 32'h10408000;
      27812: inst = 32'hc404c64;
      27813: inst = 32'h8220000;
      27814: inst = 32'h10408000;
      27815: inst = 32'hc404c65;
      27816: inst = 32'h8220000;
      27817: inst = 32'h10408000;
      27818: inst = 32'hc404c66;
      27819: inst = 32'h8220000;
      27820: inst = 32'h10408000;
      27821: inst = 32'hc404c67;
      27822: inst = 32'h8220000;
      27823: inst = 32'h10408000;
      27824: inst = 32'hc404c68;
      27825: inst = 32'h8220000;
      27826: inst = 32'h10408000;
      27827: inst = 32'hc404c69;
      27828: inst = 32'h8220000;
      27829: inst = 32'h10408000;
      27830: inst = 32'hc404c6a;
      27831: inst = 32'h8220000;
      27832: inst = 32'h10408000;
      27833: inst = 32'hc404c6b;
      27834: inst = 32'h8220000;
      27835: inst = 32'h10408000;
      27836: inst = 32'hc404c6c;
      27837: inst = 32'h8220000;
      27838: inst = 32'h10408000;
      27839: inst = 32'hc404c6d;
      27840: inst = 32'h8220000;
      27841: inst = 32'h10408000;
      27842: inst = 32'hc404c6e;
      27843: inst = 32'h8220000;
      27844: inst = 32'h10408000;
      27845: inst = 32'hc404c6f;
      27846: inst = 32'h8220000;
      27847: inst = 32'h10408000;
      27848: inst = 32'hc404c70;
      27849: inst = 32'h8220000;
      27850: inst = 32'h10408000;
      27851: inst = 32'hc404c71;
      27852: inst = 32'h8220000;
      27853: inst = 32'h10408000;
      27854: inst = 32'hc404c72;
      27855: inst = 32'h8220000;
      27856: inst = 32'h10408000;
      27857: inst = 32'hc404c73;
      27858: inst = 32'h8220000;
      27859: inst = 32'h10408000;
      27860: inst = 32'hc404c74;
      27861: inst = 32'h8220000;
      27862: inst = 32'h10408000;
      27863: inst = 32'hc404c75;
      27864: inst = 32'h8220000;
      27865: inst = 32'h10408000;
      27866: inst = 32'hc404c76;
      27867: inst = 32'h8220000;
      27868: inst = 32'h10408000;
      27869: inst = 32'hc404c77;
      27870: inst = 32'h8220000;
      27871: inst = 32'h10408000;
      27872: inst = 32'hc404c78;
      27873: inst = 32'h8220000;
      27874: inst = 32'h10408000;
      27875: inst = 32'hc404c79;
      27876: inst = 32'h8220000;
      27877: inst = 32'h10408000;
      27878: inst = 32'hc404c7a;
      27879: inst = 32'h8220000;
      27880: inst = 32'h10408000;
      27881: inst = 32'hc404c7b;
      27882: inst = 32'h8220000;
      27883: inst = 32'h10408000;
      27884: inst = 32'hc404c7c;
      27885: inst = 32'h8220000;
      27886: inst = 32'h10408000;
      27887: inst = 32'hc404c7d;
      27888: inst = 32'h8220000;
      27889: inst = 32'h10408000;
      27890: inst = 32'hc404c7e;
      27891: inst = 32'h8220000;
      27892: inst = 32'h10408000;
      27893: inst = 32'hc404c7f;
      27894: inst = 32'h8220000;
      27895: inst = 32'h10408000;
      27896: inst = 32'hc404c80;
      27897: inst = 32'h8220000;
      27898: inst = 32'h10408000;
      27899: inst = 32'hc404c81;
      27900: inst = 32'h8220000;
      27901: inst = 32'h10408000;
      27902: inst = 32'hc404c82;
      27903: inst = 32'h8220000;
      27904: inst = 32'h10408000;
      27905: inst = 32'hc404c83;
      27906: inst = 32'h8220000;
      27907: inst = 32'h10408000;
      27908: inst = 32'hc404c84;
      27909: inst = 32'h8220000;
      27910: inst = 32'h10408000;
      27911: inst = 32'hc404c85;
      27912: inst = 32'h8220000;
      27913: inst = 32'h10408000;
      27914: inst = 32'hc404c86;
      27915: inst = 32'h8220000;
      27916: inst = 32'h10408000;
      27917: inst = 32'hc404c87;
      27918: inst = 32'h8220000;
      27919: inst = 32'h10408000;
      27920: inst = 32'hc404c88;
      27921: inst = 32'h8220000;
      27922: inst = 32'h10408000;
      27923: inst = 32'hc404c89;
      27924: inst = 32'h8220000;
      27925: inst = 32'h10408000;
      27926: inst = 32'hc404c8a;
      27927: inst = 32'h8220000;
      27928: inst = 32'h10408000;
      27929: inst = 32'hc404c8b;
      27930: inst = 32'h8220000;
      27931: inst = 32'h10408000;
      27932: inst = 32'hc404c8c;
      27933: inst = 32'h8220000;
      27934: inst = 32'h10408000;
      27935: inst = 32'hc404c8d;
      27936: inst = 32'h8220000;
      27937: inst = 32'h10408000;
      27938: inst = 32'hc404c8e;
      27939: inst = 32'h8220000;
      27940: inst = 32'h10408000;
      27941: inst = 32'hc404c8f;
      27942: inst = 32'h8220000;
      27943: inst = 32'h10408000;
      27944: inst = 32'hc404c90;
      27945: inst = 32'h8220000;
      27946: inst = 32'h10408000;
      27947: inst = 32'hc404c91;
      27948: inst = 32'h8220000;
      27949: inst = 32'h10408000;
      27950: inst = 32'hc404c92;
      27951: inst = 32'h8220000;
      27952: inst = 32'h10408000;
      27953: inst = 32'hc404c93;
      27954: inst = 32'h8220000;
      27955: inst = 32'h10408000;
      27956: inst = 32'hc404c94;
      27957: inst = 32'h8220000;
      27958: inst = 32'h10408000;
      27959: inst = 32'hc404c95;
      27960: inst = 32'h8220000;
      27961: inst = 32'h10408000;
      27962: inst = 32'hc404c96;
      27963: inst = 32'h8220000;
      27964: inst = 32'h10408000;
      27965: inst = 32'hc404c97;
      27966: inst = 32'h8220000;
      27967: inst = 32'h10408000;
      27968: inst = 32'hc404c98;
      27969: inst = 32'h8220000;
      27970: inst = 32'h10408000;
      27971: inst = 32'hc404ca7;
      27972: inst = 32'h8220000;
      27973: inst = 32'h10408000;
      27974: inst = 32'hc404ca8;
      27975: inst = 32'h8220000;
      27976: inst = 32'h10408000;
      27977: inst = 32'hc404ca9;
      27978: inst = 32'h8220000;
      27979: inst = 32'h10408000;
      27980: inst = 32'hc404caa;
      27981: inst = 32'h8220000;
      27982: inst = 32'h10408000;
      27983: inst = 32'hc404cab;
      27984: inst = 32'h8220000;
      27985: inst = 32'h10408000;
      27986: inst = 32'hc404cac;
      27987: inst = 32'h8220000;
      27988: inst = 32'h10408000;
      27989: inst = 32'hc404cad;
      27990: inst = 32'h8220000;
      27991: inst = 32'h10408000;
      27992: inst = 32'hc404cae;
      27993: inst = 32'h8220000;
      27994: inst = 32'h10408000;
      27995: inst = 32'hc404cb2;
      27996: inst = 32'h8220000;
      27997: inst = 32'h10408000;
      27998: inst = 32'hc404cb3;
      27999: inst = 32'h8220000;
      28000: inst = 32'h10408000;
      28001: inst = 32'hc404cb4;
      28002: inst = 32'h8220000;
      28003: inst = 32'h10408000;
      28004: inst = 32'hc404cb5;
      28005: inst = 32'h8220000;
      28006: inst = 32'h10408000;
      28007: inst = 32'hc404cb6;
      28008: inst = 32'h8220000;
      28009: inst = 32'h10408000;
      28010: inst = 32'hc404cb7;
      28011: inst = 32'h8220000;
      28012: inst = 32'h10408000;
      28013: inst = 32'hc404cb8;
      28014: inst = 32'h8220000;
      28015: inst = 32'h10408000;
      28016: inst = 32'hc404cb9;
      28017: inst = 32'h8220000;
      28018: inst = 32'h10408000;
      28019: inst = 32'hc404cba;
      28020: inst = 32'h8220000;
      28021: inst = 32'h10408000;
      28022: inst = 32'hc404cbb;
      28023: inst = 32'h8220000;
      28024: inst = 32'h10408000;
      28025: inst = 32'hc404cbc;
      28026: inst = 32'h8220000;
      28027: inst = 32'h10408000;
      28028: inst = 32'hc404cbd;
      28029: inst = 32'h8220000;
      28030: inst = 32'h10408000;
      28031: inst = 32'hc404cbe;
      28032: inst = 32'h8220000;
      28033: inst = 32'h10408000;
      28034: inst = 32'hc404cbf;
      28035: inst = 32'h8220000;
      28036: inst = 32'h10408000;
      28037: inst = 32'hc404cc0;
      28038: inst = 32'h8220000;
      28039: inst = 32'h10408000;
      28040: inst = 32'hc404cc1;
      28041: inst = 32'h8220000;
      28042: inst = 32'h10408000;
      28043: inst = 32'hc404cc2;
      28044: inst = 32'h8220000;
      28045: inst = 32'h10408000;
      28046: inst = 32'hc404cc3;
      28047: inst = 32'h8220000;
      28048: inst = 32'h10408000;
      28049: inst = 32'hc404cc4;
      28050: inst = 32'h8220000;
      28051: inst = 32'h10408000;
      28052: inst = 32'hc404cc5;
      28053: inst = 32'h8220000;
      28054: inst = 32'h10408000;
      28055: inst = 32'hc404cc6;
      28056: inst = 32'h8220000;
      28057: inst = 32'h10408000;
      28058: inst = 32'hc404cc7;
      28059: inst = 32'h8220000;
      28060: inst = 32'h10408000;
      28061: inst = 32'hc404cc8;
      28062: inst = 32'h8220000;
      28063: inst = 32'h10408000;
      28064: inst = 32'hc404cc9;
      28065: inst = 32'h8220000;
      28066: inst = 32'h10408000;
      28067: inst = 32'hc404cca;
      28068: inst = 32'h8220000;
      28069: inst = 32'h10408000;
      28070: inst = 32'hc404ccb;
      28071: inst = 32'h8220000;
      28072: inst = 32'h10408000;
      28073: inst = 32'hc404ccc;
      28074: inst = 32'h8220000;
      28075: inst = 32'h10408000;
      28076: inst = 32'hc404ccd;
      28077: inst = 32'h8220000;
      28078: inst = 32'h10408000;
      28079: inst = 32'hc404cce;
      28080: inst = 32'h8220000;
      28081: inst = 32'h10408000;
      28082: inst = 32'hc404ccf;
      28083: inst = 32'h8220000;
      28084: inst = 32'h10408000;
      28085: inst = 32'hc404cd0;
      28086: inst = 32'h8220000;
      28087: inst = 32'h10408000;
      28088: inst = 32'hc404cd1;
      28089: inst = 32'h8220000;
      28090: inst = 32'h10408000;
      28091: inst = 32'hc404cd2;
      28092: inst = 32'h8220000;
      28093: inst = 32'h10408000;
      28094: inst = 32'hc404cd3;
      28095: inst = 32'h8220000;
      28096: inst = 32'h10408000;
      28097: inst = 32'hc404cd4;
      28098: inst = 32'h8220000;
      28099: inst = 32'h10408000;
      28100: inst = 32'hc404cd5;
      28101: inst = 32'h8220000;
      28102: inst = 32'h10408000;
      28103: inst = 32'hc404cd6;
      28104: inst = 32'h8220000;
      28105: inst = 32'h10408000;
      28106: inst = 32'hc404cd7;
      28107: inst = 32'h8220000;
      28108: inst = 32'h10408000;
      28109: inst = 32'hc404cd8;
      28110: inst = 32'h8220000;
      28111: inst = 32'h10408000;
      28112: inst = 32'hc404cd9;
      28113: inst = 32'h8220000;
      28114: inst = 32'h10408000;
      28115: inst = 32'hc404cda;
      28116: inst = 32'h8220000;
      28117: inst = 32'h10408000;
      28118: inst = 32'hc404cdb;
      28119: inst = 32'h8220000;
      28120: inst = 32'h10408000;
      28121: inst = 32'hc404cdc;
      28122: inst = 32'h8220000;
      28123: inst = 32'h10408000;
      28124: inst = 32'hc404cdd;
      28125: inst = 32'h8220000;
      28126: inst = 32'h10408000;
      28127: inst = 32'hc404cde;
      28128: inst = 32'h8220000;
      28129: inst = 32'h10408000;
      28130: inst = 32'hc404cdf;
      28131: inst = 32'h8220000;
      28132: inst = 32'h10408000;
      28133: inst = 32'hc404ce0;
      28134: inst = 32'h8220000;
      28135: inst = 32'h10408000;
      28136: inst = 32'hc404ce1;
      28137: inst = 32'h8220000;
      28138: inst = 32'h10408000;
      28139: inst = 32'hc404ce2;
      28140: inst = 32'h8220000;
      28141: inst = 32'h10408000;
      28142: inst = 32'hc404ce3;
      28143: inst = 32'h8220000;
      28144: inst = 32'h10408000;
      28145: inst = 32'hc404ce4;
      28146: inst = 32'h8220000;
      28147: inst = 32'h10408000;
      28148: inst = 32'hc404ce5;
      28149: inst = 32'h8220000;
      28150: inst = 32'h10408000;
      28151: inst = 32'hc404ce6;
      28152: inst = 32'h8220000;
      28153: inst = 32'h10408000;
      28154: inst = 32'hc404ce7;
      28155: inst = 32'h8220000;
      28156: inst = 32'h10408000;
      28157: inst = 32'hc404ce8;
      28158: inst = 32'h8220000;
      28159: inst = 32'h10408000;
      28160: inst = 32'hc404ce9;
      28161: inst = 32'h8220000;
      28162: inst = 32'h10408000;
      28163: inst = 32'hc404cea;
      28164: inst = 32'h8220000;
      28165: inst = 32'h10408000;
      28166: inst = 32'hc404ceb;
      28167: inst = 32'h8220000;
      28168: inst = 32'h10408000;
      28169: inst = 32'hc404cec;
      28170: inst = 32'h8220000;
      28171: inst = 32'h10408000;
      28172: inst = 32'hc404ced;
      28173: inst = 32'h8220000;
      28174: inst = 32'h10408000;
      28175: inst = 32'hc404cee;
      28176: inst = 32'h8220000;
      28177: inst = 32'h10408000;
      28178: inst = 32'hc404cef;
      28179: inst = 32'h8220000;
      28180: inst = 32'h10408000;
      28181: inst = 32'hc404cf3;
      28182: inst = 32'h8220000;
      28183: inst = 32'h10408000;
      28184: inst = 32'hc404cf4;
      28185: inst = 32'h8220000;
      28186: inst = 32'h10408000;
      28187: inst = 32'hc404cf5;
      28188: inst = 32'h8220000;
      28189: inst = 32'h10408000;
      28190: inst = 32'hc404cf6;
      28191: inst = 32'h8220000;
      28192: inst = 32'h10408000;
      28193: inst = 32'hc404cf7;
      28194: inst = 32'h8220000;
      28195: inst = 32'h10408000;
      28196: inst = 32'hc404cf8;
      28197: inst = 32'h8220000;
      28198: inst = 32'h10408000;
      28199: inst = 32'hc404d07;
      28200: inst = 32'h8220000;
      28201: inst = 32'h10408000;
      28202: inst = 32'hc404d08;
      28203: inst = 32'h8220000;
      28204: inst = 32'h10408000;
      28205: inst = 32'hc404d09;
      28206: inst = 32'h8220000;
      28207: inst = 32'h10408000;
      28208: inst = 32'hc404d0a;
      28209: inst = 32'h8220000;
      28210: inst = 32'h10408000;
      28211: inst = 32'hc404d0b;
      28212: inst = 32'h8220000;
      28213: inst = 32'h10408000;
      28214: inst = 32'hc404d0c;
      28215: inst = 32'h8220000;
      28216: inst = 32'h10408000;
      28217: inst = 32'hc404d0d;
      28218: inst = 32'h8220000;
      28219: inst = 32'h10408000;
      28220: inst = 32'hc404d0e;
      28221: inst = 32'h8220000;
      28222: inst = 32'h10408000;
      28223: inst = 32'hc404d12;
      28224: inst = 32'h8220000;
      28225: inst = 32'h10408000;
      28226: inst = 32'hc404d13;
      28227: inst = 32'h8220000;
      28228: inst = 32'h10408000;
      28229: inst = 32'hc404d14;
      28230: inst = 32'h8220000;
      28231: inst = 32'h10408000;
      28232: inst = 32'hc404d15;
      28233: inst = 32'h8220000;
      28234: inst = 32'h10408000;
      28235: inst = 32'hc404d16;
      28236: inst = 32'h8220000;
      28237: inst = 32'h10408000;
      28238: inst = 32'hc404d17;
      28239: inst = 32'h8220000;
      28240: inst = 32'h10408000;
      28241: inst = 32'hc404d18;
      28242: inst = 32'h8220000;
      28243: inst = 32'h10408000;
      28244: inst = 32'hc404d19;
      28245: inst = 32'h8220000;
      28246: inst = 32'h10408000;
      28247: inst = 32'hc404d1a;
      28248: inst = 32'h8220000;
      28249: inst = 32'h10408000;
      28250: inst = 32'hc404d1b;
      28251: inst = 32'h8220000;
      28252: inst = 32'h10408000;
      28253: inst = 32'hc404d1c;
      28254: inst = 32'h8220000;
      28255: inst = 32'h10408000;
      28256: inst = 32'hc404d1d;
      28257: inst = 32'h8220000;
      28258: inst = 32'h10408000;
      28259: inst = 32'hc404d1e;
      28260: inst = 32'h8220000;
      28261: inst = 32'h10408000;
      28262: inst = 32'hc404d1f;
      28263: inst = 32'h8220000;
      28264: inst = 32'h10408000;
      28265: inst = 32'hc404d20;
      28266: inst = 32'h8220000;
      28267: inst = 32'h10408000;
      28268: inst = 32'hc404d22;
      28269: inst = 32'h8220000;
      28270: inst = 32'h10408000;
      28271: inst = 32'hc404d23;
      28272: inst = 32'h8220000;
      28273: inst = 32'h10408000;
      28274: inst = 32'hc404d24;
      28275: inst = 32'h8220000;
      28276: inst = 32'h10408000;
      28277: inst = 32'hc404d25;
      28278: inst = 32'h8220000;
      28279: inst = 32'h10408000;
      28280: inst = 32'hc404d26;
      28281: inst = 32'h8220000;
      28282: inst = 32'h10408000;
      28283: inst = 32'hc404d27;
      28284: inst = 32'h8220000;
      28285: inst = 32'h10408000;
      28286: inst = 32'hc404d28;
      28287: inst = 32'h8220000;
      28288: inst = 32'h10408000;
      28289: inst = 32'hc404d29;
      28290: inst = 32'h8220000;
      28291: inst = 32'h10408000;
      28292: inst = 32'hc404d2a;
      28293: inst = 32'h8220000;
      28294: inst = 32'h10408000;
      28295: inst = 32'hc404d2c;
      28296: inst = 32'h8220000;
      28297: inst = 32'h10408000;
      28298: inst = 32'hc404d2d;
      28299: inst = 32'h8220000;
      28300: inst = 32'h10408000;
      28301: inst = 32'hc404d2e;
      28302: inst = 32'h8220000;
      28303: inst = 32'h10408000;
      28304: inst = 32'hc404d2f;
      28305: inst = 32'h8220000;
      28306: inst = 32'h10408000;
      28307: inst = 32'hc404d30;
      28308: inst = 32'h8220000;
      28309: inst = 32'h10408000;
      28310: inst = 32'hc404d31;
      28311: inst = 32'h8220000;
      28312: inst = 32'h10408000;
      28313: inst = 32'hc404d32;
      28314: inst = 32'h8220000;
      28315: inst = 32'h10408000;
      28316: inst = 32'hc404d33;
      28317: inst = 32'h8220000;
      28318: inst = 32'h10408000;
      28319: inst = 32'hc404d34;
      28320: inst = 32'h8220000;
      28321: inst = 32'h10408000;
      28322: inst = 32'hc404d35;
      28323: inst = 32'h8220000;
      28324: inst = 32'h10408000;
      28325: inst = 32'hc404d36;
      28326: inst = 32'h8220000;
      28327: inst = 32'h10408000;
      28328: inst = 32'hc404d37;
      28329: inst = 32'h8220000;
      28330: inst = 32'h10408000;
      28331: inst = 32'hc404d38;
      28332: inst = 32'h8220000;
      28333: inst = 32'h10408000;
      28334: inst = 32'hc404d39;
      28335: inst = 32'h8220000;
      28336: inst = 32'h10408000;
      28337: inst = 32'hc404d3a;
      28338: inst = 32'h8220000;
      28339: inst = 32'h10408000;
      28340: inst = 32'hc404d3b;
      28341: inst = 32'h8220000;
      28342: inst = 32'h10408000;
      28343: inst = 32'hc404d3c;
      28344: inst = 32'h8220000;
      28345: inst = 32'h10408000;
      28346: inst = 32'hc404d3d;
      28347: inst = 32'h8220000;
      28348: inst = 32'h10408000;
      28349: inst = 32'hc404d3e;
      28350: inst = 32'h8220000;
      28351: inst = 32'h10408000;
      28352: inst = 32'hc404d40;
      28353: inst = 32'h8220000;
      28354: inst = 32'h10408000;
      28355: inst = 32'hc404d41;
      28356: inst = 32'h8220000;
      28357: inst = 32'h10408000;
      28358: inst = 32'hc404d42;
      28359: inst = 32'h8220000;
      28360: inst = 32'h10408000;
      28361: inst = 32'hc404d43;
      28362: inst = 32'h8220000;
      28363: inst = 32'h10408000;
      28364: inst = 32'hc404d45;
      28365: inst = 32'h8220000;
      28366: inst = 32'h10408000;
      28367: inst = 32'hc404d46;
      28368: inst = 32'h8220000;
      28369: inst = 32'h10408000;
      28370: inst = 32'hc404d47;
      28371: inst = 32'h8220000;
      28372: inst = 32'h10408000;
      28373: inst = 32'hc404d48;
      28374: inst = 32'h8220000;
      28375: inst = 32'h10408000;
      28376: inst = 32'hc404d49;
      28377: inst = 32'h8220000;
      28378: inst = 32'h10408000;
      28379: inst = 32'hc404d4a;
      28380: inst = 32'h8220000;
      28381: inst = 32'h10408000;
      28382: inst = 32'hc404d4b;
      28383: inst = 32'h8220000;
      28384: inst = 32'h10408000;
      28385: inst = 32'hc404d4c;
      28386: inst = 32'h8220000;
      28387: inst = 32'h10408000;
      28388: inst = 32'hc404d4d;
      28389: inst = 32'h8220000;
      28390: inst = 32'h10408000;
      28391: inst = 32'hc404d4e;
      28392: inst = 32'h8220000;
      28393: inst = 32'h10408000;
      28394: inst = 32'hc404d4f;
      28395: inst = 32'h8220000;
      28396: inst = 32'h10408000;
      28397: inst = 32'hc404d53;
      28398: inst = 32'h8220000;
      28399: inst = 32'h10408000;
      28400: inst = 32'hc404d54;
      28401: inst = 32'h8220000;
      28402: inst = 32'h10408000;
      28403: inst = 32'hc404d55;
      28404: inst = 32'h8220000;
      28405: inst = 32'h10408000;
      28406: inst = 32'hc404d56;
      28407: inst = 32'h8220000;
      28408: inst = 32'h10408000;
      28409: inst = 32'hc404d57;
      28410: inst = 32'h8220000;
      28411: inst = 32'h10408000;
      28412: inst = 32'hc404d58;
      28413: inst = 32'h8220000;
      28414: inst = 32'h10408000;
      28415: inst = 32'hc404d67;
      28416: inst = 32'h8220000;
      28417: inst = 32'h10408000;
      28418: inst = 32'hc404d68;
      28419: inst = 32'h8220000;
      28420: inst = 32'h10408000;
      28421: inst = 32'hc404d69;
      28422: inst = 32'h8220000;
      28423: inst = 32'h10408000;
      28424: inst = 32'hc404d6a;
      28425: inst = 32'h8220000;
      28426: inst = 32'h10408000;
      28427: inst = 32'hc404d6b;
      28428: inst = 32'h8220000;
      28429: inst = 32'h10408000;
      28430: inst = 32'hc404d6c;
      28431: inst = 32'h8220000;
      28432: inst = 32'h10408000;
      28433: inst = 32'hc404d6d;
      28434: inst = 32'h8220000;
      28435: inst = 32'h10408000;
      28436: inst = 32'hc404d6e;
      28437: inst = 32'h8220000;
      28438: inst = 32'h10408000;
      28439: inst = 32'hc404d6f;
      28440: inst = 32'h8220000;
      28441: inst = 32'h10408000;
      28442: inst = 32'hc404d72;
      28443: inst = 32'h8220000;
      28444: inst = 32'h10408000;
      28445: inst = 32'hc404d73;
      28446: inst = 32'h8220000;
      28447: inst = 32'h10408000;
      28448: inst = 32'hc404d74;
      28449: inst = 32'h8220000;
      28450: inst = 32'h10408000;
      28451: inst = 32'hc404d75;
      28452: inst = 32'h8220000;
      28453: inst = 32'h10408000;
      28454: inst = 32'hc404d76;
      28455: inst = 32'h8220000;
      28456: inst = 32'h10408000;
      28457: inst = 32'hc404d77;
      28458: inst = 32'h8220000;
      28459: inst = 32'h10408000;
      28460: inst = 32'hc404d78;
      28461: inst = 32'h8220000;
      28462: inst = 32'h10408000;
      28463: inst = 32'hc404d79;
      28464: inst = 32'h8220000;
      28465: inst = 32'h10408000;
      28466: inst = 32'hc404d7a;
      28467: inst = 32'h8220000;
      28468: inst = 32'h10408000;
      28469: inst = 32'hc404d7b;
      28470: inst = 32'h8220000;
      28471: inst = 32'h10408000;
      28472: inst = 32'hc404d7c;
      28473: inst = 32'h8220000;
      28474: inst = 32'h10408000;
      28475: inst = 32'hc404d7d;
      28476: inst = 32'h8220000;
      28477: inst = 32'h10408000;
      28478: inst = 32'hc404d7e;
      28479: inst = 32'h8220000;
      28480: inst = 32'h10408000;
      28481: inst = 32'hc404d7f;
      28482: inst = 32'h8220000;
      28483: inst = 32'h10408000;
      28484: inst = 32'hc404d82;
      28485: inst = 32'h8220000;
      28486: inst = 32'h10408000;
      28487: inst = 32'hc404d83;
      28488: inst = 32'h8220000;
      28489: inst = 32'h10408000;
      28490: inst = 32'hc404d84;
      28491: inst = 32'h8220000;
      28492: inst = 32'h10408000;
      28493: inst = 32'hc404d85;
      28494: inst = 32'h8220000;
      28495: inst = 32'h10408000;
      28496: inst = 32'hc404d86;
      28497: inst = 32'h8220000;
      28498: inst = 32'h10408000;
      28499: inst = 32'hc404d87;
      28500: inst = 32'h8220000;
      28501: inst = 32'h10408000;
      28502: inst = 32'hc404d88;
      28503: inst = 32'h8220000;
      28504: inst = 32'h10408000;
      28505: inst = 32'hc404d89;
      28506: inst = 32'h8220000;
      28507: inst = 32'h10408000;
      28508: inst = 32'hc404d8c;
      28509: inst = 32'h8220000;
      28510: inst = 32'h10408000;
      28511: inst = 32'hc404d8d;
      28512: inst = 32'h8220000;
      28513: inst = 32'h10408000;
      28514: inst = 32'hc404d8e;
      28515: inst = 32'h8220000;
      28516: inst = 32'h10408000;
      28517: inst = 32'hc404d8f;
      28518: inst = 32'h8220000;
      28519: inst = 32'h10408000;
      28520: inst = 32'hc404d90;
      28521: inst = 32'h8220000;
      28522: inst = 32'h10408000;
      28523: inst = 32'hc404d91;
      28524: inst = 32'h8220000;
      28525: inst = 32'h10408000;
      28526: inst = 32'hc404d92;
      28527: inst = 32'h8220000;
      28528: inst = 32'h10408000;
      28529: inst = 32'hc404d93;
      28530: inst = 32'h8220000;
      28531: inst = 32'h10408000;
      28532: inst = 32'hc404d94;
      28533: inst = 32'h8220000;
      28534: inst = 32'h10408000;
      28535: inst = 32'hc404d95;
      28536: inst = 32'h8220000;
      28537: inst = 32'h10408000;
      28538: inst = 32'hc404d96;
      28539: inst = 32'h8220000;
      28540: inst = 32'h10408000;
      28541: inst = 32'hc404d97;
      28542: inst = 32'h8220000;
      28543: inst = 32'h10408000;
      28544: inst = 32'hc404d98;
      28545: inst = 32'h8220000;
      28546: inst = 32'h10408000;
      28547: inst = 32'hc404d99;
      28548: inst = 32'h8220000;
      28549: inst = 32'h10408000;
      28550: inst = 32'hc404d9a;
      28551: inst = 32'h8220000;
      28552: inst = 32'h10408000;
      28553: inst = 32'hc404d9b;
      28554: inst = 32'h8220000;
      28555: inst = 32'h10408000;
      28556: inst = 32'hc404d9c;
      28557: inst = 32'h8220000;
      28558: inst = 32'h10408000;
      28559: inst = 32'hc404d9d;
      28560: inst = 32'h8220000;
      28561: inst = 32'h10408000;
      28562: inst = 32'hc404da0;
      28563: inst = 32'h8220000;
      28564: inst = 32'h10408000;
      28565: inst = 32'hc404da1;
      28566: inst = 32'h8220000;
      28567: inst = 32'h10408000;
      28568: inst = 32'hc404da2;
      28569: inst = 32'h8220000;
      28570: inst = 32'h10408000;
      28571: inst = 32'hc404da5;
      28572: inst = 32'h8220000;
      28573: inst = 32'h10408000;
      28574: inst = 32'hc404da6;
      28575: inst = 32'h8220000;
      28576: inst = 32'h10408000;
      28577: inst = 32'hc404da7;
      28578: inst = 32'h8220000;
      28579: inst = 32'h10408000;
      28580: inst = 32'hc404da8;
      28581: inst = 32'h8220000;
      28582: inst = 32'h10408000;
      28583: inst = 32'hc404da9;
      28584: inst = 32'h8220000;
      28585: inst = 32'h10408000;
      28586: inst = 32'hc404daa;
      28587: inst = 32'h8220000;
      28588: inst = 32'h10408000;
      28589: inst = 32'hc404dab;
      28590: inst = 32'h8220000;
      28591: inst = 32'h10408000;
      28592: inst = 32'hc404dac;
      28593: inst = 32'h8220000;
      28594: inst = 32'h10408000;
      28595: inst = 32'hc404dad;
      28596: inst = 32'h8220000;
      28597: inst = 32'h10408000;
      28598: inst = 32'hc404dae;
      28599: inst = 32'h8220000;
      28600: inst = 32'h10408000;
      28601: inst = 32'hc404daf;
      28602: inst = 32'h8220000;
      28603: inst = 32'h10408000;
      28604: inst = 32'hc404db0;
      28605: inst = 32'h8220000;
      28606: inst = 32'h10408000;
      28607: inst = 32'hc404db3;
      28608: inst = 32'h8220000;
      28609: inst = 32'h10408000;
      28610: inst = 32'hc404db4;
      28611: inst = 32'h8220000;
      28612: inst = 32'h10408000;
      28613: inst = 32'hc404db5;
      28614: inst = 32'h8220000;
      28615: inst = 32'h10408000;
      28616: inst = 32'hc404db6;
      28617: inst = 32'h8220000;
      28618: inst = 32'h10408000;
      28619: inst = 32'hc404db7;
      28620: inst = 32'h8220000;
      28621: inst = 32'h10408000;
      28622: inst = 32'hc404db8;
      28623: inst = 32'h8220000;
      28624: inst = 32'h10408000;
      28625: inst = 32'hc404dc7;
      28626: inst = 32'h8220000;
      28627: inst = 32'h10408000;
      28628: inst = 32'hc404dc8;
      28629: inst = 32'h8220000;
      28630: inst = 32'h10408000;
      28631: inst = 32'hc404dc9;
      28632: inst = 32'h8220000;
      28633: inst = 32'h10408000;
      28634: inst = 32'hc404dca;
      28635: inst = 32'h8220000;
      28636: inst = 32'h10408000;
      28637: inst = 32'hc404dcb;
      28638: inst = 32'h8220000;
      28639: inst = 32'h10408000;
      28640: inst = 32'hc404dd4;
      28641: inst = 32'h8220000;
      28642: inst = 32'h10408000;
      28643: inst = 32'hc404dd5;
      28644: inst = 32'h8220000;
      28645: inst = 32'h10408000;
      28646: inst = 32'hc404dd9;
      28647: inst = 32'h8220000;
      28648: inst = 32'h10408000;
      28649: inst = 32'hc404ddc;
      28650: inst = 32'h8220000;
      28651: inst = 32'h10408000;
      28652: inst = 32'hc404de3;
      28653: inst = 32'h8220000;
      28654: inst = 32'h10408000;
      28655: inst = 32'hc404de4;
      28656: inst = 32'h8220000;
      28657: inst = 32'h10408000;
      28658: inst = 32'hc404de5;
      28659: inst = 32'h8220000;
      28660: inst = 32'h10408000;
      28661: inst = 32'hc404de6;
      28662: inst = 32'h8220000;
      28663: inst = 32'h10408000;
      28664: inst = 32'hc404de7;
      28665: inst = 32'h8220000;
      28666: inst = 32'h10408000;
      28667: inst = 32'hc404de8;
      28668: inst = 32'h8220000;
      28669: inst = 32'h10408000;
      28670: inst = 32'hc404ded;
      28671: inst = 32'h8220000;
      28672: inst = 32'h10408000;
      28673: inst = 32'hc404dee;
      28674: inst = 32'h8220000;
      28675: inst = 32'h10408000;
      28676: inst = 32'hc404df2;
      28677: inst = 32'h8220000;
      28678: inst = 32'h10408000;
      28679: inst = 32'hc404df3;
      28680: inst = 32'h8220000;
      28681: inst = 32'h10408000;
      28682: inst = 32'hc404df4;
      28683: inst = 32'h8220000;
      28684: inst = 32'h10408000;
      28685: inst = 32'hc404df5;
      28686: inst = 32'h8220000;
      28687: inst = 32'h10408000;
      28688: inst = 32'hc404df6;
      28689: inst = 32'h8220000;
      28690: inst = 32'h10408000;
      28691: inst = 32'hc404df7;
      28692: inst = 32'h8220000;
      28693: inst = 32'h10408000;
      28694: inst = 32'hc404df8;
      28695: inst = 32'h8220000;
      28696: inst = 32'h10408000;
      28697: inst = 32'hc404dfc;
      28698: inst = 32'h8220000;
      28699: inst = 32'h10408000;
      28700: inst = 32'hc404e01;
      28701: inst = 32'h8220000;
      28702: inst = 32'h10408000;
      28703: inst = 32'hc404e06;
      28704: inst = 32'h8220000;
      28705: inst = 32'h10408000;
      28706: inst = 32'hc404e07;
      28707: inst = 32'h8220000;
      28708: inst = 32'h10408000;
      28709: inst = 32'hc404e0b;
      28710: inst = 32'h8220000;
      28711: inst = 32'h10408000;
      28712: inst = 32'hc404e0c;
      28713: inst = 32'h8220000;
      28714: inst = 32'h10408000;
      28715: inst = 32'hc404e0d;
      28716: inst = 32'h8220000;
      28717: inst = 32'h10408000;
      28718: inst = 32'hc404e10;
      28719: inst = 32'h8220000;
      28720: inst = 32'h10408000;
      28721: inst = 32'hc404e13;
      28722: inst = 32'h8220000;
      28723: inst = 32'h10408000;
      28724: inst = 32'hc404e16;
      28725: inst = 32'h8220000;
      28726: inst = 32'h10408000;
      28727: inst = 32'hc404e17;
      28728: inst = 32'h8220000;
      28729: inst = 32'h10408000;
      28730: inst = 32'hc404e18;
      28731: inst = 32'h8220000;
      28732: inst = 32'h10408000;
      28733: inst = 32'hc404e27;
      28734: inst = 32'h8220000;
      28735: inst = 32'h10408000;
      28736: inst = 32'hc404e28;
      28737: inst = 32'h8220000;
      28738: inst = 32'h10408000;
      28739: inst = 32'hc404e29;
      28740: inst = 32'h8220000;
      28741: inst = 32'h10408000;
      28742: inst = 32'hc404e2a;
      28743: inst = 32'h8220000;
      28744: inst = 32'h10408000;
      28745: inst = 32'hc404e3c;
      28746: inst = 32'h8220000;
      28747: inst = 32'h10408000;
      28748: inst = 32'hc404e44;
      28749: inst = 32'h8220000;
      28750: inst = 32'h10408000;
      28751: inst = 32'hc404e45;
      28752: inst = 32'h8220000;
      28753: inst = 32'h10408000;
      28754: inst = 32'hc404e46;
      28755: inst = 32'h8220000;
      28756: inst = 32'h10408000;
      28757: inst = 32'hc404e47;
      28758: inst = 32'h8220000;
      28759: inst = 32'h10408000;
      28760: inst = 32'hc404e48;
      28761: inst = 32'h8220000;
      28762: inst = 32'h10408000;
      28763: inst = 32'hc404e53;
      28764: inst = 32'h8220000;
      28765: inst = 32'h10408000;
      28766: inst = 32'hc404e54;
      28767: inst = 32'h8220000;
      28768: inst = 32'h10408000;
      28769: inst = 32'hc404e55;
      28770: inst = 32'h8220000;
      28771: inst = 32'h10408000;
      28772: inst = 32'hc404e56;
      28773: inst = 32'h8220000;
      28774: inst = 32'h10408000;
      28775: inst = 32'hc404e57;
      28776: inst = 32'h8220000;
      28777: inst = 32'h10408000;
      28778: inst = 32'hc404e76;
      28779: inst = 32'h8220000;
      28780: inst = 32'h10408000;
      28781: inst = 32'hc404e77;
      28782: inst = 32'h8220000;
      28783: inst = 32'h10408000;
      28784: inst = 32'hc404e78;
      28785: inst = 32'h8220000;
      28786: inst = 32'h10408000;
      28787: inst = 32'hc404e87;
      28788: inst = 32'h8220000;
      28789: inst = 32'h10408000;
      28790: inst = 32'hc404e88;
      28791: inst = 32'h8220000;
      28792: inst = 32'h10408000;
      28793: inst = 32'hc404e89;
      28794: inst = 32'h8220000;
      28795: inst = 32'h10408000;
      28796: inst = 32'hc404e8a;
      28797: inst = 32'h8220000;
      28798: inst = 32'h10408000;
      28799: inst = 32'hc404e8d;
      28800: inst = 32'h8220000;
      28801: inst = 32'h10408000;
      28802: inst = 32'hc404e8e;
      28803: inst = 32'h8220000;
      28804: inst = 32'h10408000;
      28805: inst = 32'hc404e92;
      28806: inst = 32'h8220000;
      28807: inst = 32'h10408000;
      28808: inst = 32'hc404e97;
      28809: inst = 32'h8220000;
      28810: inst = 32'h10408000;
      28811: inst = 32'hc404e9c;
      28812: inst = 32'h8220000;
      28813: inst = 32'h10408000;
      28814: inst = 32'hc404e9f;
      28815: inst = 32'h8220000;
      28816: inst = 32'h10408000;
      28817: inst = 32'hc404ea2;
      28818: inst = 32'h8220000;
      28819: inst = 32'h10408000;
      28820: inst = 32'hc404ea3;
      28821: inst = 32'h8220000;
      28822: inst = 32'h10408000;
      28823: inst = 32'hc404ea4;
      28824: inst = 32'h8220000;
      28825: inst = 32'h10408000;
      28826: inst = 32'hc404ea5;
      28827: inst = 32'h8220000;
      28828: inst = 32'h10408000;
      28829: inst = 32'hc404ea6;
      28830: inst = 32'h8220000;
      28831: inst = 32'h10408000;
      28832: inst = 32'hc404ea7;
      28833: inst = 32'h8220000;
      28834: inst = 32'h10408000;
      28835: inst = 32'hc404ea8;
      28836: inst = 32'h8220000;
      28837: inst = 32'h10408000;
      28838: inst = 32'hc404ea9;
      28839: inst = 32'h8220000;
      28840: inst = 32'h10408000;
      28841: inst = 32'hc404eac;
      28842: inst = 32'h8220000;
      28843: inst = 32'h10408000;
      28844: inst = 32'hc404ead;
      28845: inst = 32'h8220000;
      28846: inst = 32'h10408000;
      28847: inst = 32'hc404eb0;
      28848: inst = 32'h8220000;
      28849: inst = 32'h10408000;
      28850: inst = 32'hc404eb3;
      28851: inst = 32'h8220000;
      28852: inst = 32'h10408000;
      28853: inst = 32'hc404eb4;
      28854: inst = 32'h8220000;
      28855: inst = 32'h10408000;
      28856: inst = 32'hc404eb5;
      28857: inst = 32'h8220000;
      28858: inst = 32'h10408000;
      28859: inst = 32'hc404eb6;
      28860: inst = 32'h8220000;
      28861: inst = 32'h10408000;
      28862: inst = 32'hc404eb7;
      28863: inst = 32'h8220000;
      28864: inst = 32'h10408000;
      28865: inst = 32'hc404eba;
      28866: inst = 32'h8220000;
      28867: inst = 32'h10408000;
      28868: inst = 32'hc404ebd;
      28869: inst = 32'h8220000;
      28870: inst = 32'h10408000;
      28871: inst = 32'hc404ec0;
      28872: inst = 32'h8220000;
      28873: inst = 32'h10408000;
      28874: inst = 32'hc404ec1;
      28875: inst = 32'h8220000;
      28876: inst = 32'h10408000;
      28877: inst = 32'hc404ec2;
      28878: inst = 32'h8220000;
      28879: inst = 32'h10408000;
      28880: inst = 32'hc404ec5;
      28881: inst = 32'h8220000;
      28882: inst = 32'h10408000;
      28883: inst = 32'hc404ec6;
      28884: inst = 32'h8220000;
      28885: inst = 32'h10408000;
      28886: inst = 32'hc404ec9;
      28887: inst = 32'h8220000;
      28888: inst = 32'h10408000;
      28889: inst = 32'hc404ece;
      28890: inst = 32'h8220000;
      28891: inst = 32'h10408000;
      28892: inst = 32'hc404ed5;
      28893: inst = 32'h8220000;
      28894: inst = 32'h10408000;
      28895: inst = 32'hc404ed6;
      28896: inst = 32'h8220000;
      28897: inst = 32'h10408000;
      28898: inst = 32'hc404ed7;
      28899: inst = 32'h8220000;
      28900: inst = 32'h10408000;
      28901: inst = 32'hc404ed8;
      28902: inst = 32'h8220000;
      28903: inst = 32'h10408000;
      28904: inst = 32'hc404ee7;
      28905: inst = 32'h8220000;
      28906: inst = 32'h10408000;
      28907: inst = 32'hc404ee8;
      28908: inst = 32'h8220000;
      28909: inst = 32'h10408000;
      28910: inst = 32'hc404ee9;
      28911: inst = 32'h8220000;
      28912: inst = 32'h10408000;
      28913: inst = 32'hc404eea;
      28914: inst = 32'h8220000;
      28915: inst = 32'h10408000;
      28916: inst = 32'hc404eef;
      28917: inst = 32'h8220000;
      28918: inst = 32'h10408000;
      28919: inst = 32'hc404ef2;
      28920: inst = 32'h8220000;
      28921: inst = 32'h10408000;
      28922: inst = 32'hc404ef6;
      28923: inst = 32'h8220000;
      28924: inst = 32'h10408000;
      28925: inst = 32'hc404ef7;
      28926: inst = 32'h8220000;
      28927: inst = 32'h10408000;
      28928: inst = 32'hc404ef8;
      28929: inst = 32'h8220000;
      28930: inst = 32'h10408000;
      28931: inst = 32'hc404efc;
      28932: inst = 32'h8220000;
      28933: inst = 32'h10408000;
      28934: inst = 32'hc404eff;
      28935: inst = 32'h8220000;
      28936: inst = 32'h10408000;
      28937: inst = 32'hc404f02;
      28938: inst = 32'h8220000;
      28939: inst = 32'h10408000;
      28940: inst = 32'hc404f03;
      28941: inst = 32'h8220000;
      28942: inst = 32'h10408000;
      28943: inst = 32'hc404f04;
      28944: inst = 32'h8220000;
      28945: inst = 32'h10408000;
      28946: inst = 32'hc404f05;
      28947: inst = 32'h8220000;
      28948: inst = 32'h10408000;
      28949: inst = 32'hc404f06;
      28950: inst = 32'h8220000;
      28951: inst = 32'h10408000;
      28952: inst = 32'hc404f07;
      28953: inst = 32'h8220000;
      28954: inst = 32'h10408000;
      28955: inst = 32'hc404f08;
      28956: inst = 32'h8220000;
      28957: inst = 32'h10408000;
      28958: inst = 32'hc404f09;
      28959: inst = 32'h8220000;
      28960: inst = 32'h10408000;
      28961: inst = 32'hc404f0c;
      28962: inst = 32'h8220000;
      28963: inst = 32'h10408000;
      28964: inst = 32'hc404f0f;
      28965: inst = 32'h8220000;
      28966: inst = 32'h10408000;
      28967: inst = 32'hc404f10;
      28968: inst = 32'h8220000;
      28969: inst = 32'h10408000;
      28970: inst = 32'hc404f11;
      28971: inst = 32'h8220000;
      28972: inst = 32'h10408000;
      28973: inst = 32'hc404f14;
      28974: inst = 32'h8220000;
      28975: inst = 32'h10408000;
      28976: inst = 32'hc404f15;
      28977: inst = 32'h8220000;
      28978: inst = 32'h10408000;
      28979: inst = 32'hc404f16;
      28980: inst = 32'h8220000;
      28981: inst = 32'h10408000;
      28982: inst = 32'hc404f17;
      28983: inst = 32'h8220000;
      28984: inst = 32'h10408000;
      28985: inst = 32'hc404f1d;
      28986: inst = 32'h8220000;
      28987: inst = 32'h10408000;
      28988: inst = 32'hc404f20;
      28989: inst = 32'h8220000;
      28990: inst = 32'h10408000;
      28991: inst = 32'hc404f21;
      28992: inst = 32'h8220000;
      28993: inst = 32'h10408000;
      28994: inst = 32'hc404f22;
      28995: inst = 32'h8220000;
      28996: inst = 32'h10408000;
      28997: inst = 32'hc404f25;
      28998: inst = 32'h8220000;
      28999: inst = 32'h10408000;
      29000: inst = 32'hc404f26;
      29001: inst = 32'h8220000;
      29002: inst = 32'h10408000;
      29003: inst = 32'hc404f2e;
      29004: inst = 32'h8220000;
      29005: inst = 32'h10408000;
      29006: inst = 32'hc404f2f;
      29007: inst = 32'h8220000;
      29008: inst = 32'h10408000;
      29009: inst = 32'hc404f30;
      29010: inst = 32'h8220000;
      29011: inst = 32'h10408000;
      29012: inst = 32'hc404f35;
      29013: inst = 32'h8220000;
      29014: inst = 32'h10408000;
      29015: inst = 32'hc404f36;
      29016: inst = 32'h8220000;
      29017: inst = 32'h10408000;
      29018: inst = 32'hc404f37;
      29019: inst = 32'h8220000;
      29020: inst = 32'h10408000;
      29021: inst = 32'hc404f38;
      29022: inst = 32'h8220000;
      29023: inst = 32'h10408000;
      29024: inst = 32'hc404f47;
      29025: inst = 32'h8220000;
      29026: inst = 32'h10408000;
      29027: inst = 32'hc404f48;
      29028: inst = 32'h8220000;
      29029: inst = 32'h10408000;
      29030: inst = 32'hc404f49;
      29031: inst = 32'h8220000;
      29032: inst = 32'h10408000;
      29033: inst = 32'hc404f4a;
      29034: inst = 32'h8220000;
      29035: inst = 32'h10408000;
      29036: inst = 32'hc404f4b;
      29037: inst = 32'h8220000;
      29038: inst = 32'h10408000;
      29039: inst = 32'hc404f4c;
      29040: inst = 32'h8220000;
      29041: inst = 32'h10408000;
      29042: inst = 32'hc404f52;
      29043: inst = 32'h8220000;
      29044: inst = 32'h10408000;
      29045: inst = 32'hc404f56;
      29046: inst = 32'h8220000;
      29047: inst = 32'h10408000;
      29048: inst = 32'hc404f57;
      29049: inst = 32'h8220000;
      29050: inst = 32'h10408000;
      29051: inst = 32'hc404f58;
      29052: inst = 32'h8220000;
      29053: inst = 32'h10408000;
      29054: inst = 32'hc404f5c;
      29055: inst = 32'h8220000;
      29056: inst = 32'h10408000;
      29057: inst = 32'hc404f5f;
      29058: inst = 32'h8220000;
      29059: inst = 32'h10408000;
      29060: inst = 32'hc404f62;
      29061: inst = 32'h8220000;
      29062: inst = 32'h10408000;
      29063: inst = 32'hc404f63;
      29064: inst = 32'h8220000;
      29065: inst = 32'h10408000;
      29066: inst = 32'hc404f64;
      29067: inst = 32'h8220000;
      29068: inst = 32'h10408000;
      29069: inst = 32'hc404f65;
      29070: inst = 32'h8220000;
      29071: inst = 32'h10408000;
      29072: inst = 32'hc404f66;
      29073: inst = 32'h8220000;
      29074: inst = 32'h10408000;
      29075: inst = 32'hc404f67;
      29076: inst = 32'h8220000;
      29077: inst = 32'h10408000;
      29078: inst = 32'hc404f68;
      29079: inst = 32'h8220000;
      29080: inst = 32'h10408000;
      29081: inst = 32'hc404f69;
      29082: inst = 32'h8220000;
      29083: inst = 32'h10408000;
      29084: inst = 32'hc404f6c;
      29085: inst = 32'h8220000;
      29086: inst = 32'h10408000;
      29087: inst = 32'hc404f6f;
      29088: inst = 32'h8220000;
      29089: inst = 32'h10408000;
      29090: inst = 32'hc404f70;
      29091: inst = 32'h8220000;
      29092: inst = 32'h10408000;
      29093: inst = 32'hc404f71;
      29094: inst = 32'h8220000;
      29095: inst = 32'h10408000;
      29096: inst = 32'hc404f74;
      29097: inst = 32'h8220000;
      29098: inst = 32'h10408000;
      29099: inst = 32'hc404f75;
      29100: inst = 32'h8220000;
      29101: inst = 32'h10408000;
      29102: inst = 32'hc404f76;
      29103: inst = 32'h8220000;
      29104: inst = 32'h10408000;
      29105: inst = 32'hc404f77;
      29106: inst = 32'h8220000;
      29107: inst = 32'h10408000;
      29108: inst = 32'hc404f7a;
      29109: inst = 32'h8220000;
      29110: inst = 32'h10408000;
      29111: inst = 32'hc404f7d;
      29112: inst = 32'h8220000;
      29113: inst = 32'h10408000;
      29114: inst = 32'hc404f80;
      29115: inst = 32'h8220000;
      29116: inst = 32'h10408000;
      29117: inst = 32'hc404f81;
      29118: inst = 32'h8220000;
      29119: inst = 32'h10408000;
      29120: inst = 32'hc404f82;
      29121: inst = 32'h8220000;
      29122: inst = 32'h10408000;
      29123: inst = 32'hc404f85;
      29124: inst = 32'h8220000;
      29125: inst = 32'h10408000;
      29126: inst = 32'hc404f86;
      29127: inst = 32'h8220000;
      29128: inst = 32'h10408000;
      29129: inst = 32'hc404f89;
      29130: inst = 32'h8220000;
      29131: inst = 32'h10408000;
      29132: inst = 32'hc404f8e;
      29133: inst = 32'h8220000;
      29134: inst = 32'h10408000;
      29135: inst = 32'hc404f8f;
      29136: inst = 32'h8220000;
      29137: inst = 32'h10408000;
      29138: inst = 32'hc404f90;
      29139: inst = 32'h8220000;
      29140: inst = 32'h10408000;
      29141: inst = 32'hc404f95;
      29142: inst = 32'h8220000;
      29143: inst = 32'h10408000;
      29144: inst = 32'hc404f96;
      29145: inst = 32'h8220000;
      29146: inst = 32'h10408000;
      29147: inst = 32'hc404f97;
      29148: inst = 32'h8220000;
      29149: inst = 32'h10408000;
      29150: inst = 32'hc404f98;
      29151: inst = 32'h8220000;
      29152: inst = 32'h10408000;
      29153: inst = 32'hc404fa7;
      29154: inst = 32'h8220000;
      29155: inst = 32'h10408000;
      29156: inst = 32'hc404fa8;
      29157: inst = 32'h8220000;
      29158: inst = 32'h10408000;
      29159: inst = 32'hc404fa9;
      29160: inst = 32'h8220000;
      29161: inst = 32'h10408000;
      29162: inst = 32'hc404faa;
      29163: inst = 32'h8220000;
      29164: inst = 32'h10408000;
      29165: inst = 32'hc404fad;
      29166: inst = 32'h8220000;
      29167: inst = 32'h10408000;
      29168: inst = 32'hc404fae;
      29169: inst = 32'h8220000;
      29170: inst = 32'h10408000;
      29171: inst = 32'hc404fb2;
      29172: inst = 32'h8220000;
      29173: inst = 32'h10408000;
      29174: inst = 32'hc404fb7;
      29175: inst = 32'h8220000;
      29176: inst = 32'h10408000;
      29177: inst = 32'hc404fbc;
      29178: inst = 32'h8220000;
      29179: inst = 32'h10408000;
      29180: inst = 32'hc404fbf;
      29181: inst = 32'h8220000;
      29182: inst = 32'h10408000;
      29183: inst = 32'hc404fc2;
      29184: inst = 32'h8220000;
      29185: inst = 32'h10408000;
      29186: inst = 32'hc404fc4;
      29187: inst = 32'h8220000;
      29188: inst = 32'h10408000;
      29189: inst = 32'hc404fc5;
      29190: inst = 32'h8220000;
      29191: inst = 32'h10408000;
      29192: inst = 32'hc404fc6;
      29193: inst = 32'h8220000;
      29194: inst = 32'h10408000;
      29195: inst = 32'hc404fc7;
      29196: inst = 32'h8220000;
      29197: inst = 32'h10408000;
      29198: inst = 32'hc404fc8;
      29199: inst = 32'h8220000;
      29200: inst = 32'h10408000;
      29201: inst = 32'hc404fc9;
      29202: inst = 32'h8220000;
      29203: inst = 32'h10408000;
      29204: inst = 32'hc404fcc;
      29205: inst = 32'h8220000;
      29206: inst = 32'h10408000;
      29207: inst = 32'hc404fd0;
      29208: inst = 32'h8220000;
      29209: inst = 32'h10408000;
      29210: inst = 32'hc404fd4;
      29211: inst = 32'h8220000;
      29212: inst = 32'h10408000;
      29213: inst = 32'hc404fd5;
      29214: inst = 32'h8220000;
      29215: inst = 32'h10408000;
      29216: inst = 32'hc404fd6;
      29217: inst = 32'h8220000;
      29218: inst = 32'h10408000;
      29219: inst = 32'hc404fd9;
      29220: inst = 32'h8220000;
      29221: inst = 32'h10408000;
      29222: inst = 32'hc404fda;
      29223: inst = 32'h8220000;
      29224: inst = 32'h10408000;
      29225: inst = 32'hc404fe0;
      29226: inst = 32'h8220000;
      29227: inst = 32'h10408000;
      29228: inst = 32'hc404fe2;
      29229: inst = 32'h8220000;
      29230: inst = 32'h10408000;
      29231: inst = 32'hc404fe5;
      29232: inst = 32'h8220000;
      29233: inst = 32'h10408000;
      29234: inst = 32'hc404fe8;
      29235: inst = 32'h8220000;
      29236: inst = 32'h10408000;
      29237: inst = 32'hc404fe9;
      29238: inst = 32'h8220000;
      29239: inst = 32'h10408000;
      29240: inst = 32'hc404fee;
      29241: inst = 32'h8220000;
      29242: inst = 32'h10408000;
      29243: inst = 32'hc404fef;
      29244: inst = 32'h8220000;
      29245: inst = 32'h10408000;
      29246: inst = 32'hc404ff3;
      29247: inst = 32'h8220000;
      29248: inst = 32'h10408000;
      29249: inst = 32'hc404ff6;
      29250: inst = 32'h8220000;
      29251: inst = 32'h10408000;
      29252: inst = 32'hc404ff7;
      29253: inst = 32'h8220000;
      29254: inst = 32'h10408000;
      29255: inst = 32'hc404ff8;
      29256: inst = 32'h8220000;
      29257: inst = 32'h10408000;
      29258: inst = 32'hc405007;
      29259: inst = 32'h8220000;
      29260: inst = 32'h10408000;
      29261: inst = 32'hc405008;
      29262: inst = 32'h8220000;
      29263: inst = 32'h10408000;
      29264: inst = 32'hc405009;
      29265: inst = 32'h8220000;
      29266: inst = 32'h10408000;
      29267: inst = 32'hc40500a;
      29268: inst = 32'h8220000;
      29269: inst = 32'h10408000;
      29270: inst = 32'hc405012;
      29271: inst = 32'h8220000;
      29272: inst = 32'h10408000;
      29273: inst = 32'hc405024;
      29274: inst = 32'h8220000;
      29275: inst = 32'h10408000;
      29276: inst = 32'hc405025;
      29277: inst = 32'h8220000;
      29278: inst = 32'h10408000;
      29279: inst = 32'hc405026;
      29280: inst = 32'h8220000;
      29281: inst = 32'h10408000;
      29282: inst = 32'hc405027;
      29283: inst = 32'h8220000;
      29284: inst = 32'h10408000;
      29285: inst = 32'hc405028;
      29286: inst = 32'h8220000;
      29287: inst = 32'h10408000;
      29288: inst = 32'hc405029;
      29289: inst = 32'h8220000;
      29290: inst = 32'h10408000;
      29291: inst = 32'hc405033;
      29292: inst = 32'h8220000;
      29293: inst = 32'h10408000;
      29294: inst = 32'hc405034;
      29295: inst = 32'h8220000;
      29296: inst = 32'h10408000;
      29297: inst = 32'hc405035;
      29298: inst = 32'h8220000;
      29299: inst = 32'h10408000;
      29300: inst = 32'hc405036;
      29301: inst = 32'h8220000;
      29302: inst = 32'h10408000;
      29303: inst = 32'hc405037;
      29304: inst = 32'h8220000;
      29305: inst = 32'h10408000;
      29306: inst = 32'hc405042;
      29307: inst = 32'h8220000;
      29308: inst = 32'h10408000;
      29309: inst = 32'hc405053;
      29310: inst = 32'h8220000;
      29311: inst = 32'h10408000;
      29312: inst = 32'hc405057;
      29313: inst = 32'h8220000;
      29314: inst = 32'h10408000;
      29315: inst = 32'hc405058;
      29316: inst = 32'h8220000;
      29317: inst = 32'h10408000;
      29318: inst = 32'hc405067;
      29319: inst = 32'h8220000;
      29320: inst = 32'h10408000;
      29321: inst = 32'hc405068;
      29322: inst = 32'h8220000;
      29323: inst = 32'h10408000;
      29324: inst = 32'hc405069;
      29325: inst = 32'h8220000;
      29326: inst = 32'h10408000;
      29327: inst = 32'hc40506a;
      29328: inst = 32'h8220000;
      29329: inst = 32'h10408000;
      29330: inst = 32'hc40506c;
      29331: inst = 32'h8220000;
      29332: inst = 32'h10408000;
      29333: inst = 32'hc40506f;
      29334: inst = 32'h8220000;
      29335: inst = 32'h10408000;
      29336: inst = 32'hc405072;
      29337: inst = 32'h8220000;
      29338: inst = 32'h10408000;
      29339: inst = 32'hc405075;
      29340: inst = 32'h8220000;
      29341: inst = 32'h10408000;
      29342: inst = 32'hc405079;
      29343: inst = 32'h8220000;
      29344: inst = 32'h10408000;
      29345: inst = 32'hc40507a;
      29346: inst = 32'h8220000;
      29347: inst = 32'h10408000;
      29348: inst = 32'hc40507d;
      29349: inst = 32'h8220000;
      29350: inst = 32'h10408000;
      29351: inst = 32'hc40507e;
      29352: inst = 32'h8220000;
      29353: inst = 32'h10408000;
      29354: inst = 32'hc40507f;
      29355: inst = 32'h8220000;
      29356: inst = 32'h10408000;
      29357: inst = 32'hc405080;
      29358: inst = 32'h8220000;
      29359: inst = 32'h10408000;
      29360: inst = 32'hc405083;
      29361: inst = 32'h8220000;
      29362: inst = 32'h10408000;
      29363: inst = 32'hc405084;
      29364: inst = 32'h8220000;
      29365: inst = 32'h10408000;
      29366: inst = 32'hc405085;
      29367: inst = 32'h8220000;
      29368: inst = 32'h10408000;
      29369: inst = 32'hc405086;
      29370: inst = 32'h8220000;
      29371: inst = 32'h10408000;
      29372: inst = 32'hc405087;
      29373: inst = 32'h8220000;
      29374: inst = 32'h10408000;
      29375: inst = 32'hc405088;
      29376: inst = 32'h8220000;
      29377: inst = 32'h10408000;
      29378: inst = 32'hc405089;
      29379: inst = 32'h8220000;
      29380: inst = 32'h10408000;
      29381: inst = 32'hc40508a;
      29382: inst = 32'h8220000;
      29383: inst = 32'h10408000;
      29384: inst = 32'hc40508d;
      29385: inst = 32'h8220000;
      29386: inst = 32'h10408000;
      29387: inst = 32'hc40508e;
      29388: inst = 32'h8220000;
      29389: inst = 32'h10408000;
      29390: inst = 32'hc405092;
      29391: inst = 32'h8220000;
      29392: inst = 32'h10408000;
      29393: inst = 32'hc405093;
      29394: inst = 32'h8220000;
      29395: inst = 32'h10408000;
      29396: inst = 32'hc405094;
      29397: inst = 32'h8220000;
      29398: inst = 32'h10408000;
      29399: inst = 32'hc405095;
      29400: inst = 32'h8220000;
      29401: inst = 32'h10408000;
      29402: inst = 32'hc405096;
      29403: inst = 32'h8220000;
      29404: inst = 32'h10408000;
      29405: inst = 32'hc405097;
      29406: inst = 32'h8220000;
      29407: inst = 32'h10408000;
      29408: inst = 32'hc405098;
      29409: inst = 32'h8220000;
      29410: inst = 32'h10408000;
      29411: inst = 32'hc40509b;
      29412: inst = 32'h8220000;
      29413: inst = 32'h10408000;
      29414: inst = 32'hc40509d;
      29415: inst = 32'h8220000;
      29416: inst = 32'h10408000;
      29417: inst = 32'hc40509e;
      29418: inst = 32'h8220000;
      29419: inst = 32'h10408000;
      29420: inst = 32'hc4050a1;
      29421: inst = 32'h8220000;
      29422: inst = 32'h10408000;
      29423: inst = 32'hc4050a2;
      29424: inst = 32'h8220000;
      29425: inst = 32'h10408000;
      29426: inst = 32'hc4050a3;
      29427: inst = 32'h8220000;
      29428: inst = 32'h10408000;
      29429: inst = 32'hc4050a6;
      29430: inst = 32'h8220000;
      29431: inst = 32'h10408000;
      29432: inst = 32'hc4050a7;
      29433: inst = 32'h8220000;
      29434: inst = 32'h10408000;
      29435: inst = 32'hc4050aa;
      29436: inst = 32'h8220000;
      29437: inst = 32'h10408000;
      29438: inst = 32'hc4050ac;
      29439: inst = 32'h8220000;
      29440: inst = 32'h10408000;
      29441: inst = 32'hc4050b0;
      29442: inst = 32'h8220000;
      29443: inst = 32'h10408000;
      29444: inst = 32'hc4050b3;
      29445: inst = 32'h8220000;
      29446: inst = 32'h10408000;
      29447: inst = 32'hc4050b6;
      29448: inst = 32'h8220000;
      29449: inst = 32'h10408000;
      29450: inst = 32'hc4050b7;
      29451: inst = 32'h8220000;
      29452: inst = 32'h10408000;
      29453: inst = 32'hc4050b8;
      29454: inst = 32'h8220000;
      29455: inst = 32'h10408000;
      29456: inst = 32'hc4050c7;
      29457: inst = 32'h8220000;
      29458: inst = 32'h10408000;
      29459: inst = 32'hc4050c8;
      29460: inst = 32'h8220000;
      29461: inst = 32'h10408000;
      29462: inst = 32'hc4050c9;
      29463: inst = 32'h8220000;
      29464: inst = 32'h10408000;
      29465: inst = 32'hc4050ca;
      29466: inst = 32'h8220000;
      29467: inst = 32'h10408000;
      29468: inst = 32'hc4050cb;
      29469: inst = 32'h8220000;
      29470: inst = 32'h10408000;
      29471: inst = 32'hc4050cc;
      29472: inst = 32'h8220000;
      29473: inst = 32'h10408000;
      29474: inst = 32'hc4050cd;
      29475: inst = 32'h8220000;
      29476: inst = 32'h10408000;
      29477: inst = 32'hc4050ce;
      29478: inst = 32'h8220000;
      29479: inst = 32'h10408000;
      29480: inst = 32'hc4050cf;
      29481: inst = 32'h8220000;
      29482: inst = 32'h10408000;
      29483: inst = 32'hc4050d0;
      29484: inst = 32'h8220000;
      29485: inst = 32'h10408000;
      29486: inst = 32'hc4050d1;
      29487: inst = 32'h8220000;
      29488: inst = 32'h10408000;
      29489: inst = 32'hc4050d2;
      29490: inst = 32'h8220000;
      29491: inst = 32'h10408000;
      29492: inst = 32'hc4050d3;
      29493: inst = 32'h8220000;
      29494: inst = 32'h10408000;
      29495: inst = 32'hc4050d4;
      29496: inst = 32'h8220000;
      29497: inst = 32'h10408000;
      29498: inst = 32'hc4050d5;
      29499: inst = 32'h8220000;
      29500: inst = 32'h10408000;
      29501: inst = 32'hc4050d6;
      29502: inst = 32'h8220000;
      29503: inst = 32'h10408000;
      29504: inst = 32'hc4050d7;
      29505: inst = 32'h8220000;
      29506: inst = 32'h10408000;
      29507: inst = 32'hc4050d8;
      29508: inst = 32'h8220000;
      29509: inst = 32'h10408000;
      29510: inst = 32'hc4050d9;
      29511: inst = 32'h8220000;
      29512: inst = 32'h10408000;
      29513: inst = 32'hc4050da;
      29514: inst = 32'h8220000;
      29515: inst = 32'h10408000;
      29516: inst = 32'hc4050db;
      29517: inst = 32'h8220000;
      29518: inst = 32'h10408000;
      29519: inst = 32'hc4050dc;
      29520: inst = 32'h8220000;
      29521: inst = 32'h10408000;
      29522: inst = 32'hc4050dd;
      29523: inst = 32'h8220000;
      29524: inst = 32'h10408000;
      29525: inst = 32'hc4050de;
      29526: inst = 32'h8220000;
      29527: inst = 32'h10408000;
      29528: inst = 32'hc4050df;
      29529: inst = 32'h8220000;
      29530: inst = 32'h10408000;
      29531: inst = 32'hc4050e0;
      29532: inst = 32'h8220000;
      29533: inst = 32'h10408000;
      29534: inst = 32'hc4050e1;
      29535: inst = 32'h8220000;
      29536: inst = 32'h10408000;
      29537: inst = 32'hc4050e2;
      29538: inst = 32'h8220000;
      29539: inst = 32'h10408000;
      29540: inst = 32'hc4050e3;
      29541: inst = 32'h8220000;
      29542: inst = 32'h10408000;
      29543: inst = 32'hc4050e4;
      29544: inst = 32'h8220000;
      29545: inst = 32'h10408000;
      29546: inst = 32'hc4050e5;
      29547: inst = 32'h8220000;
      29548: inst = 32'h10408000;
      29549: inst = 32'hc4050e6;
      29550: inst = 32'h8220000;
      29551: inst = 32'h10408000;
      29552: inst = 32'hc4050e7;
      29553: inst = 32'h8220000;
      29554: inst = 32'h10408000;
      29555: inst = 32'hc4050e8;
      29556: inst = 32'h8220000;
      29557: inst = 32'h10408000;
      29558: inst = 32'hc4050e9;
      29559: inst = 32'h8220000;
      29560: inst = 32'h10408000;
      29561: inst = 32'hc4050ea;
      29562: inst = 32'h8220000;
      29563: inst = 32'h10408000;
      29564: inst = 32'hc4050eb;
      29565: inst = 32'h8220000;
      29566: inst = 32'h10408000;
      29567: inst = 32'hc4050ec;
      29568: inst = 32'h8220000;
      29569: inst = 32'h10408000;
      29570: inst = 32'hc4050ed;
      29571: inst = 32'h8220000;
      29572: inst = 32'h10408000;
      29573: inst = 32'hc4050ee;
      29574: inst = 32'h8220000;
      29575: inst = 32'h10408000;
      29576: inst = 32'hc4050ef;
      29577: inst = 32'h8220000;
      29578: inst = 32'h10408000;
      29579: inst = 32'hc4050f0;
      29580: inst = 32'h8220000;
      29581: inst = 32'h10408000;
      29582: inst = 32'hc4050f1;
      29583: inst = 32'h8220000;
      29584: inst = 32'h10408000;
      29585: inst = 32'hc4050f2;
      29586: inst = 32'h8220000;
      29587: inst = 32'h10408000;
      29588: inst = 32'hc4050f3;
      29589: inst = 32'h8220000;
      29590: inst = 32'h10408000;
      29591: inst = 32'hc4050f4;
      29592: inst = 32'h8220000;
      29593: inst = 32'h10408000;
      29594: inst = 32'hc4050f5;
      29595: inst = 32'h8220000;
      29596: inst = 32'h10408000;
      29597: inst = 32'hc4050f6;
      29598: inst = 32'h8220000;
      29599: inst = 32'h10408000;
      29600: inst = 32'hc4050f7;
      29601: inst = 32'h8220000;
      29602: inst = 32'h10408000;
      29603: inst = 32'hc4050f8;
      29604: inst = 32'h8220000;
      29605: inst = 32'h10408000;
      29606: inst = 32'hc4050f9;
      29607: inst = 32'h8220000;
      29608: inst = 32'h10408000;
      29609: inst = 32'hc4050fa;
      29610: inst = 32'h8220000;
      29611: inst = 32'h10408000;
      29612: inst = 32'hc4050fb;
      29613: inst = 32'h8220000;
      29614: inst = 32'h10408000;
      29615: inst = 32'hc4050fc;
      29616: inst = 32'h8220000;
      29617: inst = 32'h10408000;
      29618: inst = 32'hc4050fd;
      29619: inst = 32'h8220000;
      29620: inst = 32'h10408000;
      29621: inst = 32'hc4050fe;
      29622: inst = 32'h8220000;
      29623: inst = 32'h10408000;
      29624: inst = 32'hc4050ff;
      29625: inst = 32'h8220000;
      29626: inst = 32'h10408000;
      29627: inst = 32'hc405100;
      29628: inst = 32'h8220000;
      29629: inst = 32'h10408000;
      29630: inst = 32'hc405101;
      29631: inst = 32'h8220000;
      29632: inst = 32'h10408000;
      29633: inst = 32'hc405102;
      29634: inst = 32'h8220000;
      29635: inst = 32'h10408000;
      29636: inst = 32'hc405103;
      29637: inst = 32'h8220000;
      29638: inst = 32'h10408000;
      29639: inst = 32'hc405104;
      29640: inst = 32'h8220000;
      29641: inst = 32'h10408000;
      29642: inst = 32'hc405105;
      29643: inst = 32'h8220000;
      29644: inst = 32'h10408000;
      29645: inst = 32'hc405106;
      29646: inst = 32'h8220000;
      29647: inst = 32'h10408000;
      29648: inst = 32'hc405107;
      29649: inst = 32'h8220000;
      29650: inst = 32'h10408000;
      29651: inst = 32'hc405108;
      29652: inst = 32'h8220000;
      29653: inst = 32'h10408000;
      29654: inst = 32'hc405109;
      29655: inst = 32'h8220000;
      29656: inst = 32'h10408000;
      29657: inst = 32'hc40510a;
      29658: inst = 32'h8220000;
      29659: inst = 32'h10408000;
      29660: inst = 32'hc40510b;
      29661: inst = 32'h8220000;
      29662: inst = 32'h10408000;
      29663: inst = 32'hc40510c;
      29664: inst = 32'h8220000;
      29665: inst = 32'h10408000;
      29666: inst = 32'hc40510d;
      29667: inst = 32'h8220000;
      29668: inst = 32'h10408000;
      29669: inst = 32'hc40510e;
      29670: inst = 32'h8220000;
      29671: inst = 32'h10408000;
      29672: inst = 32'hc40510f;
      29673: inst = 32'h8220000;
      29674: inst = 32'h10408000;
      29675: inst = 32'hc405110;
      29676: inst = 32'h8220000;
      29677: inst = 32'h10408000;
      29678: inst = 32'hc405111;
      29679: inst = 32'h8220000;
      29680: inst = 32'h10408000;
      29681: inst = 32'hc405112;
      29682: inst = 32'h8220000;
      29683: inst = 32'h10408000;
      29684: inst = 32'hc405113;
      29685: inst = 32'h8220000;
      29686: inst = 32'h10408000;
      29687: inst = 32'hc405114;
      29688: inst = 32'h8220000;
      29689: inst = 32'h10408000;
      29690: inst = 32'hc405115;
      29691: inst = 32'h8220000;
      29692: inst = 32'h10408000;
      29693: inst = 32'hc405116;
      29694: inst = 32'h8220000;
      29695: inst = 32'h10408000;
      29696: inst = 32'hc405117;
      29697: inst = 32'h8220000;
      29698: inst = 32'h10408000;
      29699: inst = 32'hc405118;
      29700: inst = 32'h8220000;
      29701: inst = 32'h10408000;
      29702: inst = 32'hc405127;
      29703: inst = 32'h8220000;
      29704: inst = 32'h10408000;
      29705: inst = 32'hc405128;
      29706: inst = 32'h8220000;
      29707: inst = 32'h10408000;
      29708: inst = 32'hc405129;
      29709: inst = 32'h8220000;
      29710: inst = 32'h10408000;
      29711: inst = 32'hc40512a;
      29712: inst = 32'h8220000;
      29713: inst = 32'h10408000;
      29714: inst = 32'hc40512b;
      29715: inst = 32'h8220000;
      29716: inst = 32'h10408000;
      29717: inst = 32'hc40512c;
      29718: inst = 32'h8220000;
      29719: inst = 32'h10408000;
      29720: inst = 32'hc40512d;
      29721: inst = 32'h8220000;
      29722: inst = 32'h10408000;
      29723: inst = 32'hc40512e;
      29724: inst = 32'h8220000;
      29725: inst = 32'h10408000;
      29726: inst = 32'hc40512f;
      29727: inst = 32'h8220000;
      29728: inst = 32'h10408000;
      29729: inst = 32'hc405130;
      29730: inst = 32'h8220000;
      29731: inst = 32'h10408000;
      29732: inst = 32'hc405131;
      29733: inst = 32'h8220000;
      29734: inst = 32'h10408000;
      29735: inst = 32'hc405132;
      29736: inst = 32'h8220000;
      29737: inst = 32'h10408000;
      29738: inst = 32'hc405133;
      29739: inst = 32'h8220000;
      29740: inst = 32'h10408000;
      29741: inst = 32'hc405134;
      29742: inst = 32'h8220000;
      29743: inst = 32'h10408000;
      29744: inst = 32'hc405135;
      29745: inst = 32'h8220000;
      29746: inst = 32'h10408000;
      29747: inst = 32'hc405136;
      29748: inst = 32'h8220000;
      29749: inst = 32'h10408000;
      29750: inst = 32'hc405137;
      29751: inst = 32'h8220000;
      29752: inst = 32'h10408000;
      29753: inst = 32'hc405138;
      29754: inst = 32'h8220000;
      29755: inst = 32'h10408000;
      29756: inst = 32'hc405139;
      29757: inst = 32'h8220000;
      29758: inst = 32'h10408000;
      29759: inst = 32'hc40513a;
      29760: inst = 32'h8220000;
      29761: inst = 32'h10408000;
      29762: inst = 32'hc40513b;
      29763: inst = 32'h8220000;
      29764: inst = 32'h10408000;
      29765: inst = 32'hc40513c;
      29766: inst = 32'h8220000;
      29767: inst = 32'h10408000;
      29768: inst = 32'hc40513d;
      29769: inst = 32'h8220000;
      29770: inst = 32'h10408000;
      29771: inst = 32'hc40513e;
      29772: inst = 32'h8220000;
      29773: inst = 32'h10408000;
      29774: inst = 32'hc40513f;
      29775: inst = 32'h8220000;
      29776: inst = 32'h10408000;
      29777: inst = 32'hc405140;
      29778: inst = 32'h8220000;
      29779: inst = 32'h10408000;
      29780: inst = 32'hc405141;
      29781: inst = 32'h8220000;
      29782: inst = 32'h10408000;
      29783: inst = 32'hc405142;
      29784: inst = 32'h8220000;
      29785: inst = 32'h10408000;
      29786: inst = 32'hc405143;
      29787: inst = 32'h8220000;
      29788: inst = 32'h10408000;
      29789: inst = 32'hc405144;
      29790: inst = 32'h8220000;
      29791: inst = 32'h10408000;
      29792: inst = 32'hc405145;
      29793: inst = 32'h8220000;
      29794: inst = 32'h10408000;
      29795: inst = 32'hc405146;
      29796: inst = 32'h8220000;
      29797: inst = 32'h10408000;
      29798: inst = 32'hc405147;
      29799: inst = 32'h8220000;
      29800: inst = 32'h10408000;
      29801: inst = 32'hc405148;
      29802: inst = 32'h8220000;
      29803: inst = 32'h10408000;
      29804: inst = 32'hc405149;
      29805: inst = 32'h8220000;
      29806: inst = 32'h10408000;
      29807: inst = 32'hc40514a;
      29808: inst = 32'h8220000;
      29809: inst = 32'h10408000;
      29810: inst = 32'hc40514b;
      29811: inst = 32'h8220000;
      29812: inst = 32'h10408000;
      29813: inst = 32'hc40514c;
      29814: inst = 32'h8220000;
      29815: inst = 32'h10408000;
      29816: inst = 32'hc40514d;
      29817: inst = 32'h8220000;
      29818: inst = 32'h10408000;
      29819: inst = 32'hc40514e;
      29820: inst = 32'h8220000;
      29821: inst = 32'h10408000;
      29822: inst = 32'hc40514f;
      29823: inst = 32'h8220000;
      29824: inst = 32'h10408000;
      29825: inst = 32'hc405150;
      29826: inst = 32'h8220000;
      29827: inst = 32'h10408000;
      29828: inst = 32'hc405151;
      29829: inst = 32'h8220000;
      29830: inst = 32'h10408000;
      29831: inst = 32'hc405152;
      29832: inst = 32'h8220000;
      29833: inst = 32'h10408000;
      29834: inst = 32'hc405153;
      29835: inst = 32'h8220000;
      29836: inst = 32'h10408000;
      29837: inst = 32'hc405154;
      29838: inst = 32'h8220000;
      29839: inst = 32'h10408000;
      29840: inst = 32'hc405155;
      29841: inst = 32'h8220000;
      29842: inst = 32'h10408000;
      29843: inst = 32'hc405156;
      29844: inst = 32'h8220000;
      29845: inst = 32'h10408000;
      29846: inst = 32'hc405157;
      29847: inst = 32'h8220000;
      29848: inst = 32'h10408000;
      29849: inst = 32'hc405158;
      29850: inst = 32'h8220000;
      29851: inst = 32'h10408000;
      29852: inst = 32'hc405159;
      29853: inst = 32'h8220000;
      29854: inst = 32'h10408000;
      29855: inst = 32'hc40515a;
      29856: inst = 32'h8220000;
      29857: inst = 32'h10408000;
      29858: inst = 32'hc40515b;
      29859: inst = 32'h8220000;
      29860: inst = 32'h10408000;
      29861: inst = 32'hc40515c;
      29862: inst = 32'h8220000;
      29863: inst = 32'h10408000;
      29864: inst = 32'hc40515d;
      29865: inst = 32'h8220000;
      29866: inst = 32'h10408000;
      29867: inst = 32'hc40515e;
      29868: inst = 32'h8220000;
      29869: inst = 32'h10408000;
      29870: inst = 32'hc40515f;
      29871: inst = 32'h8220000;
      29872: inst = 32'h10408000;
      29873: inst = 32'hc405160;
      29874: inst = 32'h8220000;
      29875: inst = 32'h10408000;
      29876: inst = 32'hc405161;
      29877: inst = 32'h8220000;
      29878: inst = 32'h10408000;
      29879: inst = 32'hc405162;
      29880: inst = 32'h8220000;
      29881: inst = 32'h10408000;
      29882: inst = 32'hc405163;
      29883: inst = 32'h8220000;
      29884: inst = 32'h10408000;
      29885: inst = 32'hc405164;
      29886: inst = 32'h8220000;
      29887: inst = 32'h10408000;
      29888: inst = 32'hc405165;
      29889: inst = 32'h8220000;
      29890: inst = 32'h10408000;
      29891: inst = 32'hc405166;
      29892: inst = 32'h8220000;
      29893: inst = 32'h10408000;
      29894: inst = 32'hc405167;
      29895: inst = 32'h8220000;
      29896: inst = 32'h10408000;
      29897: inst = 32'hc405168;
      29898: inst = 32'h8220000;
      29899: inst = 32'h10408000;
      29900: inst = 32'hc405169;
      29901: inst = 32'h8220000;
      29902: inst = 32'h10408000;
      29903: inst = 32'hc40516a;
      29904: inst = 32'h8220000;
      29905: inst = 32'h10408000;
      29906: inst = 32'hc40516b;
      29907: inst = 32'h8220000;
      29908: inst = 32'h10408000;
      29909: inst = 32'hc40516c;
      29910: inst = 32'h8220000;
      29911: inst = 32'h10408000;
      29912: inst = 32'hc40516d;
      29913: inst = 32'h8220000;
      29914: inst = 32'h10408000;
      29915: inst = 32'hc40516e;
      29916: inst = 32'h8220000;
      29917: inst = 32'h10408000;
      29918: inst = 32'hc40516f;
      29919: inst = 32'h8220000;
      29920: inst = 32'h10408000;
      29921: inst = 32'hc405170;
      29922: inst = 32'h8220000;
      29923: inst = 32'h10408000;
      29924: inst = 32'hc405171;
      29925: inst = 32'h8220000;
      29926: inst = 32'h10408000;
      29927: inst = 32'hc405172;
      29928: inst = 32'h8220000;
      29929: inst = 32'h10408000;
      29930: inst = 32'hc405173;
      29931: inst = 32'h8220000;
      29932: inst = 32'h10408000;
      29933: inst = 32'hc405174;
      29934: inst = 32'h8220000;
      29935: inst = 32'h10408000;
      29936: inst = 32'hc405175;
      29937: inst = 32'h8220000;
      29938: inst = 32'h10408000;
      29939: inst = 32'hc405176;
      29940: inst = 32'h8220000;
      29941: inst = 32'h10408000;
      29942: inst = 32'hc405177;
      29943: inst = 32'h8220000;
      29944: inst = 32'h10408000;
      29945: inst = 32'hc405178;
      29946: inst = 32'h8220000;
      29947: inst = 32'h10408000;
      29948: inst = 32'hc405187;
      29949: inst = 32'h8220000;
      29950: inst = 32'h10408000;
      29951: inst = 32'hc405188;
      29952: inst = 32'h8220000;
      29953: inst = 32'h10408000;
      29954: inst = 32'hc405189;
      29955: inst = 32'h8220000;
      29956: inst = 32'h10408000;
      29957: inst = 32'hc40518a;
      29958: inst = 32'h8220000;
      29959: inst = 32'h10408000;
      29960: inst = 32'hc40518b;
      29961: inst = 32'h8220000;
      29962: inst = 32'h10408000;
      29963: inst = 32'hc40518c;
      29964: inst = 32'h8220000;
      29965: inst = 32'h10408000;
      29966: inst = 32'hc40518d;
      29967: inst = 32'h8220000;
      29968: inst = 32'h10408000;
      29969: inst = 32'hc40518e;
      29970: inst = 32'h8220000;
      29971: inst = 32'h10408000;
      29972: inst = 32'hc40518f;
      29973: inst = 32'h8220000;
      29974: inst = 32'h10408000;
      29975: inst = 32'hc405190;
      29976: inst = 32'h8220000;
      29977: inst = 32'h10408000;
      29978: inst = 32'hc405191;
      29979: inst = 32'h8220000;
      29980: inst = 32'h10408000;
      29981: inst = 32'hc405192;
      29982: inst = 32'h8220000;
      29983: inst = 32'h10408000;
      29984: inst = 32'hc405193;
      29985: inst = 32'h8220000;
      29986: inst = 32'h10408000;
      29987: inst = 32'hc405194;
      29988: inst = 32'h8220000;
      29989: inst = 32'h10408000;
      29990: inst = 32'hc405195;
      29991: inst = 32'h8220000;
      29992: inst = 32'h10408000;
      29993: inst = 32'hc405196;
      29994: inst = 32'h8220000;
      29995: inst = 32'h10408000;
      29996: inst = 32'hc405197;
      29997: inst = 32'h8220000;
      29998: inst = 32'h10408000;
      29999: inst = 32'hc405198;
      30000: inst = 32'h8220000;
      30001: inst = 32'h10408000;
      30002: inst = 32'hc405199;
      30003: inst = 32'h8220000;
      30004: inst = 32'h10408000;
      30005: inst = 32'hc40519a;
      30006: inst = 32'h8220000;
      30007: inst = 32'h10408000;
      30008: inst = 32'hc40519b;
      30009: inst = 32'h8220000;
      30010: inst = 32'h10408000;
      30011: inst = 32'hc40519c;
      30012: inst = 32'h8220000;
      30013: inst = 32'h10408000;
      30014: inst = 32'hc40519d;
      30015: inst = 32'h8220000;
      30016: inst = 32'h10408000;
      30017: inst = 32'hc40519e;
      30018: inst = 32'h8220000;
      30019: inst = 32'h10408000;
      30020: inst = 32'hc40519f;
      30021: inst = 32'h8220000;
      30022: inst = 32'h10408000;
      30023: inst = 32'hc4051a0;
      30024: inst = 32'h8220000;
      30025: inst = 32'h10408000;
      30026: inst = 32'hc4051a1;
      30027: inst = 32'h8220000;
      30028: inst = 32'h10408000;
      30029: inst = 32'hc4051a2;
      30030: inst = 32'h8220000;
      30031: inst = 32'h10408000;
      30032: inst = 32'hc4051a3;
      30033: inst = 32'h8220000;
      30034: inst = 32'h10408000;
      30035: inst = 32'hc4051a4;
      30036: inst = 32'h8220000;
      30037: inst = 32'h10408000;
      30038: inst = 32'hc4051a5;
      30039: inst = 32'h8220000;
      30040: inst = 32'h10408000;
      30041: inst = 32'hc4051a6;
      30042: inst = 32'h8220000;
      30043: inst = 32'h10408000;
      30044: inst = 32'hc4051a7;
      30045: inst = 32'h8220000;
      30046: inst = 32'h10408000;
      30047: inst = 32'hc4051a8;
      30048: inst = 32'h8220000;
      30049: inst = 32'h10408000;
      30050: inst = 32'hc4051a9;
      30051: inst = 32'h8220000;
      30052: inst = 32'h10408000;
      30053: inst = 32'hc4051aa;
      30054: inst = 32'h8220000;
      30055: inst = 32'h10408000;
      30056: inst = 32'hc4051ab;
      30057: inst = 32'h8220000;
      30058: inst = 32'h10408000;
      30059: inst = 32'hc4051ac;
      30060: inst = 32'h8220000;
      30061: inst = 32'h10408000;
      30062: inst = 32'hc4051ad;
      30063: inst = 32'h8220000;
      30064: inst = 32'h10408000;
      30065: inst = 32'hc4051ae;
      30066: inst = 32'h8220000;
      30067: inst = 32'h10408000;
      30068: inst = 32'hc4051af;
      30069: inst = 32'h8220000;
      30070: inst = 32'h10408000;
      30071: inst = 32'hc4051b0;
      30072: inst = 32'h8220000;
      30073: inst = 32'h10408000;
      30074: inst = 32'hc4051b1;
      30075: inst = 32'h8220000;
      30076: inst = 32'h10408000;
      30077: inst = 32'hc4051b2;
      30078: inst = 32'h8220000;
      30079: inst = 32'h10408000;
      30080: inst = 32'hc4051b3;
      30081: inst = 32'h8220000;
      30082: inst = 32'h10408000;
      30083: inst = 32'hc4051b4;
      30084: inst = 32'h8220000;
      30085: inst = 32'h10408000;
      30086: inst = 32'hc4051b5;
      30087: inst = 32'h8220000;
      30088: inst = 32'h10408000;
      30089: inst = 32'hc4051b6;
      30090: inst = 32'h8220000;
      30091: inst = 32'h10408000;
      30092: inst = 32'hc4051b7;
      30093: inst = 32'h8220000;
      30094: inst = 32'h10408000;
      30095: inst = 32'hc4051b8;
      30096: inst = 32'h8220000;
      30097: inst = 32'h10408000;
      30098: inst = 32'hc4051b9;
      30099: inst = 32'h8220000;
      30100: inst = 32'h10408000;
      30101: inst = 32'hc4051ba;
      30102: inst = 32'h8220000;
      30103: inst = 32'h10408000;
      30104: inst = 32'hc4051bb;
      30105: inst = 32'h8220000;
      30106: inst = 32'h10408000;
      30107: inst = 32'hc4051bc;
      30108: inst = 32'h8220000;
      30109: inst = 32'h10408000;
      30110: inst = 32'hc4051bd;
      30111: inst = 32'h8220000;
      30112: inst = 32'h10408000;
      30113: inst = 32'hc4051be;
      30114: inst = 32'h8220000;
      30115: inst = 32'h10408000;
      30116: inst = 32'hc4051bf;
      30117: inst = 32'h8220000;
      30118: inst = 32'h10408000;
      30119: inst = 32'hc4051c0;
      30120: inst = 32'h8220000;
      30121: inst = 32'h10408000;
      30122: inst = 32'hc4051c1;
      30123: inst = 32'h8220000;
      30124: inst = 32'h10408000;
      30125: inst = 32'hc4051c2;
      30126: inst = 32'h8220000;
      30127: inst = 32'h10408000;
      30128: inst = 32'hc4051c3;
      30129: inst = 32'h8220000;
      30130: inst = 32'h10408000;
      30131: inst = 32'hc4051c4;
      30132: inst = 32'h8220000;
      30133: inst = 32'h10408000;
      30134: inst = 32'hc4051c5;
      30135: inst = 32'h8220000;
      30136: inst = 32'h10408000;
      30137: inst = 32'hc4051c6;
      30138: inst = 32'h8220000;
      30139: inst = 32'h10408000;
      30140: inst = 32'hc4051c7;
      30141: inst = 32'h8220000;
      30142: inst = 32'h10408000;
      30143: inst = 32'hc4051c8;
      30144: inst = 32'h8220000;
      30145: inst = 32'h10408000;
      30146: inst = 32'hc4051c9;
      30147: inst = 32'h8220000;
      30148: inst = 32'h10408000;
      30149: inst = 32'hc4051ca;
      30150: inst = 32'h8220000;
      30151: inst = 32'h10408000;
      30152: inst = 32'hc4051cb;
      30153: inst = 32'h8220000;
      30154: inst = 32'h10408000;
      30155: inst = 32'hc4051cc;
      30156: inst = 32'h8220000;
      30157: inst = 32'h10408000;
      30158: inst = 32'hc4051cd;
      30159: inst = 32'h8220000;
      30160: inst = 32'h10408000;
      30161: inst = 32'hc4051ce;
      30162: inst = 32'h8220000;
      30163: inst = 32'h10408000;
      30164: inst = 32'hc4051cf;
      30165: inst = 32'h8220000;
      30166: inst = 32'h10408000;
      30167: inst = 32'hc4051d0;
      30168: inst = 32'h8220000;
      30169: inst = 32'h10408000;
      30170: inst = 32'hc4051d1;
      30171: inst = 32'h8220000;
      30172: inst = 32'h10408000;
      30173: inst = 32'hc4051d2;
      30174: inst = 32'h8220000;
      30175: inst = 32'h10408000;
      30176: inst = 32'hc4051d3;
      30177: inst = 32'h8220000;
      30178: inst = 32'h10408000;
      30179: inst = 32'hc4051d4;
      30180: inst = 32'h8220000;
      30181: inst = 32'h10408000;
      30182: inst = 32'hc4051d5;
      30183: inst = 32'h8220000;
      30184: inst = 32'h10408000;
      30185: inst = 32'hc4051d6;
      30186: inst = 32'h8220000;
      30187: inst = 32'h10408000;
      30188: inst = 32'hc4051d7;
      30189: inst = 32'h8220000;
      30190: inst = 32'h10408000;
      30191: inst = 32'hc4051d8;
      30192: inst = 32'h8220000;
      30193: inst = 32'h10408000;
      30194: inst = 32'hc4051e7;
      30195: inst = 32'h8220000;
      30196: inst = 32'h10408000;
      30197: inst = 32'hc4051e8;
      30198: inst = 32'h8220000;
      30199: inst = 32'h10408000;
      30200: inst = 32'hc4051e9;
      30201: inst = 32'h8220000;
      30202: inst = 32'h10408000;
      30203: inst = 32'hc4051ea;
      30204: inst = 32'h8220000;
      30205: inst = 32'h10408000;
      30206: inst = 32'hc4051eb;
      30207: inst = 32'h8220000;
      30208: inst = 32'h10408000;
      30209: inst = 32'hc4051ec;
      30210: inst = 32'h8220000;
      30211: inst = 32'h10408000;
      30212: inst = 32'hc4051ed;
      30213: inst = 32'h8220000;
      30214: inst = 32'h10408000;
      30215: inst = 32'hc4051ee;
      30216: inst = 32'h8220000;
      30217: inst = 32'h10408000;
      30218: inst = 32'hc4051ef;
      30219: inst = 32'h8220000;
      30220: inst = 32'h10408000;
      30221: inst = 32'hc4051f0;
      30222: inst = 32'h8220000;
      30223: inst = 32'h10408000;
      30224: inst = 32'hc4051f1;
      30225: inst = 32'h8220000;
      30226: inst = 32'h10408000;
      30227: inst = 32'hc4051f2;
      30228: inst = 32'h8220000;
      30229: inst = 32'h10408000;
      30230: inst = 32'hc4051f3;
      30231: inst = 32'h8220000;
      30232: inst = 32'h10408000;
      30233: inst = 32'hc4051f4;
      30234: inst = 32'h8220000;
      30235: inst = 32'h10408000;
      30236: inst = 32'hc4051f5;
      30237: inst = 32'h8220000;
      30238: inst = 32'h10408000;
      30239: inst = 32'hc4051f6;
      30240: inst = 32'h8220000;
      30241: inst = 32'h10408000;
      30242: inst = 32'hc4051f7;
      30243: inst = 32'h8220000;
      30244: inst = 32'h10408000;
      30245: inst = 32'hc4051f8;
      30246: inst = 32'h8220000;
      30247: inst = 32'h10408000;
      30248: inst = 32'hc4051f9;
      30249: inst = 32'h8220000;
      30250: inst = 32'h10408000;
      30251: inst = 32'hc4051fa;
      30252: inst = 32'h8220000;
      30253: inst = 32'h10408000;
      30254: inst = 32'hc4051fb;
      30255: inst = 32'h8220000;
      30256: inst = 32'h10408000;
      30257: inst = 32'hc4051fc;
      30258: inst = 32'h8220000;
      30259: inst = 32'h10408000;
      30260: inst = 32'hc4051fd;
      30261: inst = 32'h8220000;
      30262: inst = 32'h10408000;
      30263: inst = 32'hc4051fe;
      30264: inst = 32'h8220000;
      30265: inst = 32'h10408000;
      30266: inst = 32'hc4051ff;
      30267: inst = 32'h8220000;
      30268: inst = 32'h10408000;
      30269: inst = 32'hc405200;
      30270: inst = 32'h8220000;
      30271: inst = 32'h10408000;
      30272: inst = 32'hc405201;
      30273: inst = 32'h8220000;
      30274: inst = 32'h10408000;
      30275: inst = 32'hc405202;
      30276: inst = 32'h8220000;
      30277: inst = 32'h10408000;
      30278: inst = 32'hc405203;
      30279: inst = 32'h8220000;
      30280: inst = 32'h10408000;
      30281: inst = 32'hc405204;
      30282: inst = 32'h8220000;
      30283: inst = 32'h10408000;
      30284: inst = 32'hc405205;
      30285: inst = 32'h8220000;
      30286: inst = 32'h10408000;
      30287: inst = 32'hc405206;
      30288: inst = 32'h8220000;
      30289: inst = 32'h10408000;
      30290: inst = 32'hc405207;
      30291: inst = 32'h8220000;
      30292: inst = 32'h10408000;
      30293: inst = 32'hc405208;
      30294: inst = 32'h8220000;
      30295: inst = 32'h10408000;
      30296: inst = 32'hc405209;
      30297: inst = 32'h8220000;
      30298: inst = 32'h10408000;
      30299: inst = 32'hc40520a;
      30300: inst = 32'h8220000;
      30301: inst = 32'h10408000;
      30302: inst = 32'hc40520b;
      30303: inst = 32'h8220000;
      30304: inst = 32'h10408000;
      30305: inst = 32'hc40520c;
      30306: inst = 32'h8220000;
      30307: inst = 32'h10408000;
      30308: inst = 32'hc40520d;
      30309: inst = 32'h8220000;
      30310: inst = 32'h10408000;
      30311: inst = 32'hc40520e;
      30312: inst = 32'h8220000;
      30313: inst = 32'h10408000;
      30314: inst = 32'hc40520f;
      30315: inst = 32'h8220000;
      30316: inst = 32'h10408000;
      30317: inst = 32'hc405210;
      30318: inst = 32'h8220000;
      30319: inst = 32'h10408000;
      30320: inst = 32'hc405211;
      30321: inst = 32'h8220000;
      30322: inst = 32'h10408000;
      30323: inst = 32'hc405212;
      30324: inst = 32'h8220000;
      30325: inst = 32'h10408000;
      30326: inst = 32'hc405213;
      30327: inst = 32'h8220000;
      30328: inst = 32'h10408000;
      30329: inst = 32'hc405214;
      30330: inst = 32'h8220000;
      30331: inst = 32'h10408000;
      30332: inst = 32'hc405215;
      30333: inst = 32'h8220000;
      30334: inst = 32'h10408000;
      30335: inst = 32'hc405216;
      30336: inst = 32'h8220000;
      30337: inst = 32'h10408000;
      30338: inst = 32'hc405217;
      30339: inst = 32'h8220000;
      30340: inst = 32'h10408000;
      30341: inst = 32'hc405218;
      30342: inst = 32'h8220000;
      30343: inst = 32'h10408000;
      30344: inst = 32'hc405219;
      30345: inst = 32'h8220000;
      30346: inst = 32'h10408000;
      30347: inst = 32'hc40521a;
      30348: inst = 32'h8220000;
      30349: inst = 32'h10408000;
      30350: inst = 32'hc40521b;
      30351: inst = 32'h8220000;
      30352: inst = 32'h10408000;
      30353: inst = 32'hc40521c;
      30354: inst = 32'h8220000;
      30355: inst = 32'h10408000;
      30356: inst = 32'hc40521d;
      30357: inst = 32'h8220000;
      30358: inst = 32'h10408000;
      30359: inst = 32'hc40521e;
      30360: inst = 32'h8220000;
      30361: inst = 32'h10408000;
      30362: inst = 32'hc40521f;
      30363: inst = 32'h8220000;
      30364: inst = 32'h10408000;
      30365: inst = 32'hc405220;
      30366: inst = 32'h8220000;
      30367: inst = 32'h10408000;
      30368: inst = 32'hc405221;
      30369: inst = 32'h8220000;
      30370: inst = 32'h10408000;
      30371: inst = 32'hc405222;
      30372: inst = 32'h8220000;
      30373: inst = 32'h10408000;
      30374: inst = 32'hc405223;
      30375: inst = 32'h8220000;
      30376: inst = 32'h10408000;
      30377: inst = 32'hc405224;
      30378: inst = 32'h8220000;
      30379: inst = 32'h10408000;
      30380: inst = 32'hc405225;
      30381: inst = 32'h8220000;
      30382: inst = 32'h10408000;
      30383: inst = 32'hc405226;
      30384: inst = 32'h8220000;
      30385: inst = 32'h10408000;
      30386: inst = 32'hc405227;
      30387: inst = 32'h8220000;
      30388: inst = 32'h10408000;
      30389: inst = 32'hc405228;
      30390: inst = 32'h8220000;
      30391: inst = 32'h10408000;
      30392: inst = 32'hc405229;
      30393: inst = 32'h8220000;
      30394: inst = 32'h10408000;
      30395: inst = 32'hc40522a;
      30396: inst = 32'h8220000;
      30397: inst = 32'h10408000;
      30398: inst = 32'hc40522b;
      30399: inst = 32'h8220000;
      30400: inst = 32'h10408000;
      30401: inst = 32'hc40522c;
      30402: inst = 32'h8220000;
      30403: inst = 32'h10408000;
      30404: inst = 32'hc40522d;
      30405: inst = 32'h8220000;
      30406: inst = 32'h10408000;
      30407: inst = 32'hc40522e;
      30408: inst = 32'h8220000;
      30409: inst = 32'h10408000;
      30410: inst = 32'hc40522f;
      30411: inst = 32'h8220000;
      30412: inst = 32'h10408000;
      30413: inst = 32'hc405230;
      30414: inst = 32'h8220000;
      30415: inst = 32'h10408000;
      30416: inst = 32'hc405231;
      30417: inst = 32'h8220000;
      30418: inst = 32'h10408000;
      30419: inst = 32'hc405232;
      30420: inst = 32'h8220000;
      30421: inst = 32'h10408000;
      30422: inst = 32'hc405233;
      30423: inst = 32'h8220000;
      30424: inst = 32'h10408000;
      30425: inst = 32'hc405234;
      30426: inst = 32'h8220000;
      30427: inst = 32'h10408000;
      30428: inst = 32'hc405235;
      30429: inst = 32'h8220000;
      30430: inst = 32'h10408000;
      30431: inst = 32'hc405236;
      30432: inst = 32'h8220000;
      30433: inst = 32'h10408000;
      30434: inst = 32'hc405237;
      30435: inst = 32'h8220000;
      30436: inst = 32'h10408000;
      30437: inst = 32'hc405238;
      30438: inst = 32'h8220000;
      30439: inst = 32'h10408000;
      30440: inst = 32'hc405247;
      30441: inst = 32'h8220000;
      30442: inst = 32'h10408000;
      30443: inst = 32'hc405248;
      30444: inst = 32'h8220000;
      30445: inst = 32'h10408000;
      30446: inst = 32'hc405249;
      30447: inst = 32'h8220000;
      30448: inst = 32'h10408000;
      30449: inst = 32'hc40524a;
      30450: inst = 32'h8220000;
      30451: inst = 32'h10408000;
      30452: inst = 32'hc40524b;
      30453: inst = 32'h8220000;
      30454: inst = 32'h10408000;
      30455: inst = 32'hc40524c;
      30456: inst = 32'h8220000;
      30457: inst = 32'h10408000;
      30458: inst = 32'hc40524d;
      30459: inst = 32'h8220000;
      30460: inst = 32'h10408000;
      30461: inst = 32'hc40524e;
      30462: inst = 32'h8220000;
      30463: inst = 32'h10408000;
      30464: inst = 32'hc40524f;
      30465: inst = 32'h8220000;
      30466: inst = 32'h10408000;
      30467: inst = 32'hc405250;
      30468: inst = 32'h8220000;
      30469: inst = 32'h10408000;
      30470: inst = 32'hc405251;
      30471: inst = 32'h8220000;
      30472: inst = 32'h10408000;
      30473: inst = 32'hc405252;
      30474: inst = 32'h8220000;
      30475: inst = 32'h10408000;
      30476: inst = 32'hc405253;
      30477: inst = 32'h8220000;
      30478: inst = 32'h10408000;
      30479: inst = 32'hc405254;
      30480: inst = 32'h8220000;
      30481: inst = 32'h10408000;
      30482: inst = 32'hc405255;
      30483: inst = 32'h8220000;
      30484: inst = 32'h10408000;
      30485: inst = 32'hc405256;
      30486: inst = 32'h8220000;
      30487: inst = 32'h10408000;
      30488: inst = 32'hc405257;
      30489: inst = 32'h8220000;
      30490: inst = 32'h10408000;
      30491: inst = 32'hc405258;
      30492: inst = 32'h8220000;
      30493: inst = 32'h10408000;
      30494: inst = 32'hc405259;
      30495: inst = 32'h8220000;
      30496: inst = 32'h10408000;
      30497: inst = 32'hc40525a;
      30498: inst = 32'h8220000;
      30499: inst = 32'h10408000;
      30500: inst = 32'hc40525b;
      30501: inst = 32'h8220000;
      30502: inst = 32'h10408000;
      30503: inst = 32'hc40525c;
      30504: inst = 32'h8220000;
      30505: inst = 32'h10408000;
      30506: inst = 32'hc40525d;
      30507: inst = 32'h8220000;
      30508: inst = 32'h10408000;
      30509: inst = 32'hc40525e;
      30510: inst = 32'h8220000;
      30511: inst = 32'h10408000;
      30512: inst = 32'hc40525f;
      30513: inst = 32'h8220000;
      30514: inst = 32'h10408000;
      30515: inst = 32'hc405260;
      30516: inst = 32'h8220000;
      30517: inst = 32'h10408000;
      30518: inst = 32'hc405261;
      30519: inst = 32'h8220000;
      30520: inst = 32'h10408000;
      30521: inst = 32'hc405262;
      30522: inst = 32'h8220000;
      30523: inst = 32'h10408000;
      30524: inst = 32'hc405263;
      30525: inst = 32'h8220000;
      30526: inst = 32'h10408000;
      30527: inst = 32'hc405264;
      30528: inst = 32'h8220000;
      30529: inst = 32'h10408000;
      30530: inst = 32'hc405265;
      30531: inst = 32'h8220000;
      30532: inst = 32'h10408000;
      30533: inst = 32'hc405266;
      30534: inst = 32'h8220000;
      30535: inst = 32'h10408000;
      30536: inst = 32'hc405267;
      30537: inst = 32'h8220000;
      30538: inst = 32'h10408000;
      30539: inst = 32'hc405268;
      30540: inst = 32'h8220000;
      30541: inst = 32'h10408000;
      30542: inst = 32'hc405269;
      30543: inst = 32'h8220000;
      30544: inst = 32'h10408000;
      30545: inst = 32'hc40526a;
      30546: inst = 32'h8220000;
      30547: inst = 32'h10408000;
      30548: inst = 32'hc40526b;
      30549: inst = 32'h8220000;
      30550: inst = 32'h10408000;
      30551: inst = 32'hc40526c;
      30552: inst = 32'h8220000;
      30553: inst = 32'h10408000;
      30554: inst = 32'hc40526d;
      30555: inst = 32'h8220000;
      30556: inst = 32'h10408000;
      30557: inst = 32'hc40526e;
      30558: inst = 32'h8220000;
      30559: inst = 32'h10408000;
      30560: inst = 32'hc40526f;
      30561: inst = 32'h8220000;
      30562: inst = 32'h10408000;
      30563: inst = 32'hc405270;
      30564: inst = 32'h8220000;
      30565: inst = 32'h10408000;
      30566: inst = 32'hc405271;
      30567: inst = 32'h8220000;
      30568: inst = 32'h10408000;
      30569: inst = 32'hc405272;
      30570: inst = 32'h8220000;
      30571: inst = 32'h10408000;
      30572: inst = 32'hc405273;
      30573: inst = 32'h8220000;
      30574: inst = 32'h10408000;
      30575: inst = 32'hc405274;
      30576: inst = 32'h8220000;
      30577: inst = 32'h10408000;
      30578: inst = 32'hc405275;
      30579: inst = 32'h8220000;
      30580: inst = 32'h10408000;
      30581: inst = 32'hc405276;
      30582: inst = 32'h8220000;
      30583: inst = 32'h10408000;
      30584: inst = 32'hc405277;
      30585: inst = 32'h8220000;
      30586: inst = 32'h10408000;
      30587: inst = 32'hc405278;
      30588: inst = 32'h8220000;
      30589: inst = 32'h10408000;
      30590: inst = 32'hc405279;
      30591: inst = 32'h8220000;
      30592: inst = 32'h10408000;
      30593: inst = 32'hc40527a;
      30594: inst = 32'h8220000;
      30595: inst = 32'h10408000;
      30596: inst = 32'hc40527b;
      30597: inst = 32'h8220000;
      30598: inst = 32'h10408000;
      30599: inst = 32'hc40527c;
      30600: inst = 32'h8220000;
      30601: inst = 32'h10408000;
      30602: inst = 32'hc40527d;
      30603: inst = 32'h8220000;
      30604: inst = 32'h10408000;
      30605: inst = 32'hc40527e;
      30606: inst = 32'h8220000;
      30607: inst = 32'h10408000;
      30608: inst = 32'hc40527f;
      30609: inst = 32'h8220000;
      30610: inst = 32'h10408000;
      30611: inst = 32'hc405280;
      30612: inst = 32'h8220000;
      30613: inst = 32'h10408000;
      30614: inst = 32'hc405281;
      30615: inst = 32'h8220000;
      30616: inst = 32'h10408000;
      30617: inst = 32'hc405282;
      30618: inst = 32'h8220000;
      30619: inst = 32'h10408000;
      30620: inst = 32'hc405283;
      30621: inst = 32'h8220000;
      30622: inst = 32'h10408000;
      30623: inst = 32'hc405284;
      30624: inst = 32'h8220000;
      30625: inst = 32'h10408000;
      30626: inst = 32'hc405285;
      30627: inst = 32'h8220000;
      30628: inst = 32'h10408000;
      30629: inst = 32'hc405286;
      30630: inst = 32'h8220000;
      30631: inst = 32'h10408000;
      30632: inst = 32'hc405287;
      30633: inst = 32'h8220000;
      30634: inst = 32'h10408000;
      30635: inst = 32'hc405288;
      30636: inst = 32'h8220000;
      30637: inst = 32'h10408000;
      30638: inst = 32'hc405289;
      30639: inst = 32'h8220000;
      30640: inst = 32'h10408000;
      30641: inst = 32'hc40528a;
      30642: inst = 32'h8220000;
      30643: inst = 32'h10408000;
      30644: inst = 32'hc40528b;
      30645: inst = 32'h8220000;
      30646: inst = 32'h10408000;
      30647: inst = 32'hc40528c;
      30648: inst = 32'h8220000;
      30649: inst = 32'h10408000;
      30650: inst = 32'hc40528d;
      30651: inst = 32'h8220000;
      30652: inst = 32'h10408000;
      30653: inst = 32'hc40528e;
      30654: inst = 32'h8220000;
      30655: inst = 32'h10408000;
      30656: inst = 32'hc40528f;
      30657: inst = 32'h8220000;
      30658: inst = 32'h10408000;
      30659: inst = 32'hc405290;
      30660: inst = 32'h8220000;
      30661: inst = 32'h10408000;
      30662: inst = 32'hc405291;
      30663: inst = 32'h8220000;
      30664: inst = 32'h10408000;
      30665: inst = 32'hc405292;
      30666: inst = 32'h8220000;
      30667: inst = 32'h10408000;
      30668: inst = 32'hc405293;
      30669: inst = 32'h8220000;
      30670: inst = 32'h10408000;
      30671: inst = 32'hc405294;
      30672: inst = 32'h8220000;
      30673: inst = 32'h10408000;
      30674: inst = 32'hc405295;
      30675: inst = 32'h8220000;
      30676: inst = 32'h10408000;
      30677: inst = 32'hc405296;
      30678: inst = 32'h8220000;
      30679: inst = 32'h10408000;
      30680: inst = 32'hc405297;
      30681: inst = 32'h8220000;
      30682: inst = 32'h10408000;
      30683: inst = 32'hc405298;
      30684: inst = 32'h8220000;
      30685: inst = 32'h10408000;
      30686: inst = 32'hc4052a7;
      30687: inst = 32'h8220000;
      30688: inst = 32'h10408000;
      30689: inst = 32'hc4052a8;
      30690: inst = 32'h8220000;
      30691: inst = 32'h10408000;
      30692: inst = 32'hc4052a9;
      30693: inst = 32'h8220000;
      30694: inst = 32'h10408000;
      30695: inst = 32'hc4052aa;
      30696: inst = 32'h8220000;
      30697: inst = 32'h10408000;
      30698: inst = 32'hc4052ab;
      30699: inst = 32'h8220000;
      30700: inst = 32'h10408000;
      30701: inst = 32'hc4052ac;
      30702: inst = 32'h8220000;
      30703: inst = 32'h10408000;
      30704: inst = 32'hc4052ad;
      30705: inst = 32'h8220000;
      30706: inst = 32'h10408000;
      30707: inst = 32'hc4052ae;
      30708: inst = 32'h8220000;
      30709: inst = 32'h10408000;
      30710: inst = 32'hc4052af;
      30711: inst = 32'h8220000;
      30712: inst = 32'h10408000;
      30713: inst = 32'hc4052b0;
      30714: inst = 32'h8220000;
      30715: inst = 32'h10408000;
      30716: inst = 32'hc4052b1;
      30717: inst = 32'h8220000;
      30718: inst = 32'h10408000;
      30719: inst = 32'hc4052b2;
      30720: inst = 32'h8220000;
      30721: inst = 32'h10408000;
      30722: inst = 32'hc4052b3;
      30723: inst = 32'h8220000;
      30724: inst = 32'h10408000;
      30725: inst = 32'hc4052b4;
      30726: inst = 32'h8220000;
      30727: inst = 32'h10408000;
      30728: inst = 32'hc4052b5;
      30729: inst = 32'h8220000;
      30730: inst = 32'h10408000;
      30731: inst = 32'hc4052b6;
      30732: inst = 32'h8220000;
      30733: inst = 32'h10408000;
      30734: inst = 32'hc4052b7;
      30735: inst = 32'h8220000;
      30736: inst = 32'h10408000;
      30737: inst = 32'hc4052b8;
      30738: inst = 32'h8220000;
      30739: inst = 32'h10408000;
      30740: inst = 32'hc4052b9;
      30741: inst = 32'h8220000;
      30742: inst = 32'h10408000;
      30743: inst = 32'hc4052ba;
      30744: inst = 32'h8220000;
      30745: inst = 32'h10408000;
      30746: inst = 32'hc4052bb;
      30747: inst = 32'h8220000;
      30748: inst = 32'h10408000;
      30749: inst = 32'hc4052bc;
      30750: inst = 32'h8220000;
      30751: inst = 32'h10408000;
      30752: inst = 32'hc4052bd;
      30753: inst = 32'h8220000;
      30754: inst = 32'h10408000;
      30755: inst = 32'hc4052be;
      30756: inst = 32'h8220000;
      30757: inst = 32'h10408000;
      30758: inst = 32'hc4052bf;
      30759: inst = 32'h8220000;
      30760: inst = 32'h10408000;
      30761: inst = 32'hc4052c0;
      30762: inst = 32'h8220000;
      30763: inst = 32'h10408000;
      30764: inst = 32'hc4052c1;
      30765: inst = 32'h8220000;
      30766: inst = 32'h10408000;
      30767: inst = 32'hc4052c2;
      30768: inst = 32'h8220000;
      30769: inst = 32'h10408000;
      30770: inst = 32'hc4052c3;
      30771: inst = 32'h8220000;
      30772: inst = 32'h10408000;
      30773: inst = 32'hc4052c4;
      30774: inst = 32'h8220000;
      30775: inst = 32'h10408000;
      30776: inst = 32'hc4052c5;
      30777: inst = 32'h8220000;
      30778: inst = 32'h10408000;
      30779: inst = 32'hc4052c6;
      30780: inst = 32'h8220000;
      30781: inst = 32'h10408000;
      30782: inst = 32'hc4052c7;
      30783: inst = 32'h8220000;
      30784: inst = 32'h10408000;
      30785: inst = 32'hc4052c8;
      30786: inst = 32'h8220000;
      30787: inst = 32'h10408000;
      30788: inst = 32'hc4052c9;
      30789: inst = 32'h8220000;
      30790: inst = 32'h10408000;
      30791: inst = 32'hc4052ca;
      30792: inst = 32'h8220000;
      30793: inst = 32'h10408000;
      30794: inst = 32'hc4052cb;
      30795: inst = 32'h8220000;
      30796: inst = 32'h10408000;
      30797: inst = 32'hc4052cc;
      30798: inst = 32'h8220000;
      30799: inst = 32'h10408000;
      30800: inst = 32'hc4052cd;
      30801: inst = 32'h8220000;
      30802: inst = 32'h10408000;
      30803: inst = 32'hc4052ce;
      30804: inst = 32'h8220000;
      30805: inst = 32'h10408000;
      30806: inst = 32'hc4052cf;
      30807: inst = 32'h8220000;
      30808: inst = 32'h10408000;
      30809: inst = 32'hc4052d0;
      30810: inst = 32'h8220000;
      30811: inst = 32'h10408000;
      30812: inst = 32'hc4052d1;
      30813: inst = 32'h8220000;
      30814: inst = 32'h10408000;
      30815: inst = 32'hc4052d2;
      30816: inst = 32'h8220000;
      30817: inst = 32'h10408000;
      30818: inst = 32'hc4052d3;
      30819: inst = 32'h8220000;
      30820: inst = 32'h10408000;
      30821: inst = 32'hc4052d4;
      30822: inst = 32'h8220000;
      30823: inst = 32'h10408000;
      30824: inst = 32'hc4052d5;
      30825: inst = 32'h8220000;
      30826: inst = 32'h10408000;
      30827: inst = 32'hc4052d6;
      30828: inst = 32'h8220000;
      30829: inst = 32'h10408000;
      30830: inst = 32'hc4052d7;
      30831: inst = 32'h8220000;
      30832: inst = 32'h10408000;
      30833: inst = 32'hc4052d8;
      30834: inst = 32'h8220000;
      30835: inst = 32'h10408000;
      30836: inst = 32'hc4052d9;
      30837: inst = 32'h8220000;
      30838: inst = 32'h10408000;
      30839: inst = 32'hc4052da;
      30840: inst = 32'h8220000;
      30841: inst = 32'h10408000;
      30842: inst = 32'hc4052db;
      30843: inst = 32'h8220000;
      30844: inst = 32'h10408000;
      30845: inst = 32'hc4052dc;
      30846: inst = 32'h8220000;
      30847: inst = 32'h10408000;
      30848: inst = 32'hc4052dd;
      30849: inst = 32'h8220000;
      30850: inst = 32'h10408000;
      30851: inst = 32'hc4052de;
      30852: inst = 32'h8220000;
      30853: inst = 32'h10408000;
      30854: inst = 32'hc4052df;
      30855: inst = 32'h8220000;
      30856: inst = 32'h10408000;
      30857: inst = 32'hc4052e0;
      30858: inst = 32'h8220000;
      30859: inst = 32'h10408000;
      30860: inst = 32'hc4052e1;
      30861: inst = 32'h8220000;
      30862: inst = 32'h10408000;
      30863: inst = 32'hc4052e2;
      30864: inst = 32'h8220000;
      30865: inst = 32'h10408000;
      30866: inst = 32'hc4052e3;
      30867: inst = 32'h8220000;
      30868: inst = 32'h10408000;
      30869: inst = 32'hc4052e4;
      30870: inst = 32'h8220000;
      30871: inst = 32'h10408000;
      30872: inst = 32'hc4052e5;
      30873: inst = 32'h8220000;
      30874: inst = 32'h10408000;
      30875: inst = 32'hc4052e6;
      30876: inst = 32'h8220000;
      30877: inst = 32'h10408000;
      30878: inst = 32'hc4052e7;
      30879: inst = 32'h8220000;
      30880: inst = 32'h10408000;
      30881: inst = 32'hc4052e8;
      30882: inst = 32'h8220000;
      30883: inst = 32'h10408000;
      30884: inst = 32'hc4052e9;
      30885: inst = 32'h8220000;
      30886: inst = 32'h10408000;
      30887: inst = 32'hc4052ea;
      30888: inst = 32'h8220000;
      30889: inst = 32'h10408000;
      30890: inst = 32'hc4052eb;
      30891: inst = 32'h8220000;
      30892: inst = 32'h10408000;
      30893: inst = 32'hc4052ec;
      30894: inst = 32'h8220000;
      30895: inst = 32'h10408000;
      30896: inst = 32'hc4052ed;
      30897: inst = 32'h8220000;
      30898: inst = 32'h10408000;
      30899: inst = 32'hc4052ee;
      30900: inst = 32'h8220000;
      30901: inst = 32'h10408000;
      30902: inst = 32'hc4052ef;
      30903: inst = 32'h8220000;
      30904: inst = 32'h10408000;
      30905: inst = 32'hc4052f0;
      30906: inst = 32'h8220000;
      30907: inst = 32'h10408000;
      30908: inst = 32'hc4052f1;
      30909: inst = 32'h8220000;
      30910: inst = 32'h10408000;
      30911: inst = 32'hc4052f2;
      30912: inst = 32'h8220000;
      30913: inst = 32'h10408000;
      30914: inst = 32'hc4052f3;
      30915: inst = 32'h8220000;
      30916: inst = 32'h10408000;
      30917: inst = 32'hc4052f4;
      30918: inst = 32'h8220000;
      30919: inst = 32'h10408000;
      30920: inst = 32'hc4052f5;
      30921: inst = 32'h8220000;
      30922: inst = 32'h10408000;
      30923: inst = 32'hc4052f6;
      30924: inst = 32'h8220000;
      30925: inst = 32'h10408000;
      30926: inst = 32'hc4052f7;
      30927: inst = 32'h8220000;
      30928: inst = 32'h10408000;
      30929: inst = 32'hc4052f8;
      30930: inst = 32'h8220000;
      30931: inst = 32'h10408000;
      30932: inst = 32'hc405307;
      30933: inst = 32'h8220000;
      30934: inst = 32'h10408000;
      30935: inst = 32'hc405308;
      30936: inst = 32'h8220000;
      30937: inst = 32'h10408000;
      30938: inst = 32'hc405309;
      30939: inst = 32'h8220000;
      30940: inst = 32'h10408000;
      30941: inst = 32'hc40530a;
      30942: inst = 32'h8220000;
      30943: inst = 32'h10408000;
      30944: inst = 32'hc40530b;
      30945: inst = 32'h8220000;
      30946: inst = 32'h10408000;
      30947: inst = 32'hc40530c;
      30948: inst = 32'h8220000;
      30949: inst = 32'h10408000;
      30950: inst = 32'hc40530d;
      30951: inst = 32'h8220000;
      30952: inst = 32'h10408000;
      30953: inst = 32'hc40530e;
      30954: inst = 32'h8220000;
      30955: inst = 32'h10408000;
      30956: inst = 32'hc40530f;
      30957: inst = 32'h8220000;
      30958: inst = 32'h10408000;
      30959: inst = 32'hc405310;
      30960: inst = 32'h8220000;
      30961: inst = 32'h10408000;
      30962: inst = 32'hc405311;
      30963: inst = 32'h8220000;
      30964: inst = 32'h10408000;
      30965: inst = 32'hc405312;
      30966: inst = 32'h8220000;
      30967: inst = 32'h10408000;
      30968: inst = 32'hc405313;
      30969: inst = 32'h8220000;
      30970: inst = 32'h10408000;
      30971: inst = 32'hc405314;
      30972: inst = 32'h8220000;
      30973: inst = 32'h10408000;
      30974: inst = 32'hc405315;
      30975: inst = 32'h8220000;
      30976: inst = 32'h10408000;
      30977: inst = 32'hc405316;
      30978: inst = 32'h8220000;
      30979: inst = 32'h10408000;
      30980: inst = 32'hc405317;
      30981: inst = 32'h8220000;
      30982: inst = 32'h10408000;
      30983: inst = 32'hc405318;
      30984: inst = 32'h8220000;
      30985: inst = 32'h10408000;
      30986: inst = 32'hc405319;
      30987: inst = 32'h8220000;
      30988: inst = 32'h10408000;
      30989: inst = 32'hc40531a;
      30990: inst = 32'h8220000;
      30991: inst = 32'h10408000;
      30992: inst = 32'hc40531b;
      30993: inst = 32'h8220000;
      30994: inst = 32'h10408000;
      30995: inst = 32'hc40531c;
      30996: inst = 32'h8220000;
      30997: inst = 32'h10408000;
      30998: inst = 32'hc40531d;
      30999: inst = 32'h8220000;
      31000: inst = 32'h10408000;
      31001: inst = 32'hc40531e;
      31002: inst = 32'h8220000;
      31003: inst = 32'h10408000;
      31004: inst = 32'hc40531f;
      31005: inst = 32'h8220000;
      31006: inst = 32'h10408000;
      31007: inst = 32'hc405320;
      31008: inst = 32'h8220000;
      31009: inst = 32'h10408000;
      31010: inst = 32'hc405321;
      31011: inst = 32'h8220000;
      31012: inst = 32'h10408000;
      31013: inst = 32'hc405322;
      31014: inst = 32'h8220000;
      31015: inst = 32'h10408000;
      31016: inst = 32'hc405323;
      31017: inst = 32'h8220000;
      31018: inst = 32'h10408000;
      31019: inst = 32'hc405324;
      31020: inst = 32'h8220000;
      31021: inst = 32'h10408000;
      31022: inst = 32'hc405325;
      31023: inst = 32'h8220000;
      31024: inst = 32'h10408000;
      31025: inst = 32'hc405326;
      31026: inst = 32'h8220000;
      31027: inst = 32'h10408000;
      31028: inst = 32'hc405327;
      31029: inst = 32'h8220000;
      31030: inst = 32'h10408000;
      31031: inst = 32'hc405328;
      31032: inst = 32'h8220000;
      31033: inst = 32'h10408000;
      31034: inst = 32'hc405329;
      31035: inst = 32'h8220000;
      31036: inst = 32'h10408000;
      31037: inst = 32'hc40532a;
      31038: inst = 32'h8220000;
      31039: inst = 32'h10408000;
      31040: inst = 32'hc40532b;
      31041: inst = 32'h8220000;
      31042: inst = 32'h10408000;
      31043: inst = 32'hc40532c;
      31044: inst = 32'h8220000;
      31045: inst = 32'h10408000;
      31046: inst = 32'hc40532d;
      31047: inst = 32'h8220000;
      31048: inst = 32'h10408000;
      31049: inst = 32'hc40532e;
      31050: inst = 32'h8220000;
      31051: inst = 32'h10408000;
      31052: inst = 32'hc40532f;
      31053: inst = 32'h8220000;
      31054: inst = 32'h10408000;
      31055: inst = 32'hc405330;
      31056: inst = 32'h8220000;
      31057: inst = 32'h10408000;
      31058: inst = 32'hc405331;
      31059: inst = 32'h8220000;
      31060: inst = 32'h10408000;
      31061: inst = 32'hc405332;
      31062: inst = 32'h8220000;
      31063: inst = 32'h10408000;
      31064: inst = 32'hc405333;
      31065: inst = 32'h8220000;
      31066: inst = 32'h10408000;
      31067: inst = 32'hc405334;
      31068: inst = 32'h8220000;
      31069: inst = 32'h10408000;
      31070: inst = 32'hc405335;
      31071: inst = 32'h8220000;
      31072: inst = 32'h10408000;
      31073: inst = 32'hc405336;
      31074: inst = 32'h8220000;
      31075: inst = 32'h10408000;
      31076: inst = 32'hc405337;
      31077: inst = 32'h8220000;
      31078: inst = 32'h10408000;
      31079: inst = 32'hc405338;
      31080: inst = 32'h8220000;
      31081: inst = 32'h10408000;
      31082: inst = 32'hc405339;
      31083: inst = 32'h8220000;
      31084: inst = 32'h10408000;
      31085: inst = 32'hc40533a;
      31086: inst = 32'h8220000;
      31087: inst = 32'h10408000;
      31088: inst = 32'hc40533b;
      31089: inst = 32'h8220000;
      31090: inst = 32'h10408000;
      31091: inst = 32'hc40533c;
      31092: inst = 32'h8220000;
      31093: inst = 32'h10408000;
      31094: inst = 32'hc40533d;
      31095: inst = 32'h8220000;
      31096: inst = 32'h10408000;
      31097: inst = 32'hc40533e;
      31098: inst = 32'h8220000;
      31099: inst = 32'h10408000;
      31100: inst = 32'hc40533f;
      31101: inst = 32'h8220000;
      31102: inst = 32'h10408000;
      31103: inst = 32'hc405340;
      31104: inst = 32'h8220000;
      31105: inst = 32'h10408000;
      31106: inst = 32'hc405341;
      31107: inst = 32'h8220000;
      31108: inst = 32'h10408000;
      31109: inst = 32'hc405342;
      31110: inst = 32'h8220000;
      31111: inst = 32'h10408000;
      31112: inst = 32'hc405343;
      31113: inst = 32'h8220000;
      31114: inst = 32'h10408000;
      31115: inst = 32'hc405344;
      31116: inst = 32'h8220000;
      31117: inst = 32'h10408000;
      31118: inst = 32'hc405345;
      31119: inst = 32'h8220000;
      31120: inst = 32'h10408000;
      31121: inst = 32'hc405346;
      31122: inst = 32'h8220000;
      31123: inst = 32'h10408000;
      31124: inst = 32'hc405347;
      31125: inst = 32'h8220000;
      31126: inst = 32'h10408000;
      31127: inst = 32'hc405348;
      31128: inst = 32'h8220000;
      31129: inst = 32'h10408000;
      31130: inst = 32'hc405349;
      31131: inst = 32'h8220000;
      31132: inst = 32'h10408000;
      31133: inst = 32'hc40534a;
      31134: inst = 32'h8220000;
      31135: inst = 32'h10408000;
      31136: inst = 32'hc40534b;
      31137: inst = 32'h8220000;
      31138: inst = 32'h10408000;
      31139: inst = 32'hc40534c;
      31140: inst = 32'h8220000;
      31141: inst = 32'h10408000;
      31142: inst = 32'hc40534d;
      31143: inst = 32'h8220000;
      31144: inst = 32'h10408000;
      31145: inst = 32'hc40534e;
      31146: inst = 32'h8220000;
      31147: inst = 32'h10408000;
      31148: inst = 32'hc40534f;
      31149: inst = 32'h8220000;
      31150: inst = 32'h10408000;
      31151: inst = 32'hc405350;
      31152: inst = 32'h8220000;
      31153: inst = 32'h10408000;
      31154: inst = 32'hc405351;
      31155: inst = 32'h8220000;
      31156: inst = 32'h10408000;
      31157: inst = 32'hc405352;
      31158: inst = 32'h8220000;
      31159: inst = 32'h10408000;
      31160: inst = 32'hc405353;
      31161: inst = 32'h8220000;
      31162: inst = 32'h10408000;
      31163: inst = 32'hc405354;
      31164: inst = 32'h8220000;
      31165: inst = 32'h10408000;
      31166: inst = 32'hc405355;
      31167: inst = 32'h8220000;
      31168: inst = 32'h10408000;
      31169: inst = 32'hc405356;
      31170: inst = 32'h8220000;
      31171: inst = 32'h10408000;
      31172: inst = 32'hc405357;
      31173: inst = 32'h8220000;
      31174: inst = 32'h10408000;
      31175: inst = 32'hc405358;
      31176: inst = 32'h8220000;
      31177: inst = 32'h10408000;
      31178: inst = 32'hc405367;
      31179: inst = 32'h8220000;
      31180: inst = 32'h10408000;
      31181: inst = 32'hc405368;
      31182: inst = 32'h8220000;
      31183: inst = 32'h10408000;
      31184: inst = 32'hc405369;
      31185: inst = 32'h8220000;
      31186: inst = 32'h10408000;
      31187: inst = 32'hc40536a;
      31188: inst = 32'h8220000;
      31189: inst = 32'h10408000;
      31190: inst = 32'hc40536b;
      31191: inst = 32'h8220000;
      31192: inst = 32'h10408000;
      31193: inst = 32'hc40536c;
      31194: inst = 32'h8220000;
      31195: inst = 32'h10408000;
      31196: inst = 32'hc40536d;
      31197: inst = 32'h8220000;
      31198: inst = 32'h10408000;
      31199: inst = 32'hc40536e;
      31200: inst = 32'h8220000;
      31201: inst = 32'h10408000;
      31202: inst = 32'hc40536f;
      31203: inst = 32'h8220000;
      31204: inst = 32'h10408000;
      31205: inst = 32'hc405370;
      31206: inst = 32'h8220000;
      31207: inst = 32'h10408000;
      31208: inst = 32'hc405371;
      31209: inst = 32'h8220000;
      31210: inst = 32'h10408000;
      31211: inst = 32'hc405372;
      31212: inst = 32'h8220000;
      31213: inst = 32'h10408000;
      31214: inst = 32'hc405373;
      31215: inst = 32'h8220000;
      31216: inst = 32'h10408000;
      31217: inst = 32'hc405374;
      31218: inst = 32'h8220000;
      31219: inst = 32'h10408000;
      31220: inst = 32'hc405375;
      31221: inst = 32'h8220000;
      31222: inst = 32'h10408000;
      31223: inst = 32'hc405376;
      31224: inst = 32'h8220000;
      31225: inst = 32'h10408000;
      31226: inst = 32'hc405377;
      31227: inst = 32'h8220000;
      31228: inst = 32'h10408000;
      31229: inst = 32'hc405378;
      31230: inst = 32'h8220000;
      31231: inst = 32'h10408000;
      31232: inst = 32'hc405379;
      31233: inst = 32'h8220000;
      31234: inst = 32'h10408000;
      31235: inst = 32'hc40537a;
      31236: inst = 32'h8220000;
      31237: inst = 32'h10408000;
      31238: inst = 32'hc40537b;
      31239: inst = 32'h8220000;
      31240: inst = 32'h10408000;
      31241: inst = 32'hc40537c;
      31242: inst = 32'h8220000;
      31243: inst = 32'h10408000;
      31244: inst = 32'hc40537d;
      31245: inst = 32'h8220000;
      31246: inst = 32'h10408000;
      31247: inst = 32'hc40537e;
      31248: inst = 32'h8220000;
      31249: inst = 32'h10408000;
      31250: inst = 32'hc40537f;
      31251: inst = 32'h8220000;
      31252: inst = 32'h10408000;
      31253: inst = 32'hc405380;
      31254: inst = 32'h8220000;
      31255: inst = 32'h10408000;
      31256: inst = 32'hc405381;
      31257: inst = 32'h8220000;
      31258: inst = 32'h10408000;
      31259: inst = 32'hc405382;
      31260: inst = 32'h8220000;
      31261: inst = 32'h10408000;
      31262: inst = 32'hc405383;
      31263: inst = 32'h8220000;
      31264: inst = 32'h10408000;
      31265: inst = 32'hc405384;
      31266: inst = 32'h8220000;
      31267: inst = 32'h10408000;
      31268: inst = 32'hc405385;
      31269: inst = 32'h8220000;
      31270: inst = 32'h10408000;
      31271: inst = 32'hc405386;
      31272: inst = 32'h8220000;
      31273: inst = 32'h10408000;
      31274: inst = 32'hc405387;
      31275: inst = 32'h8220000;
      31276: inst = 32'h10408000;
      31277: inst = 32'hc405388;
      31278: inst = 32'h8220000;
      31279: inst = 32'h10408000;
      31280: inst = 32'hc405389;
      31281: inst = 32'h8220000;
      31282: inst = 32'h10408000;
      31283: inst = 32'hc40538a;
      31284: inst = 32'h8220000;
      31285: inst = 32'h10408000;
      31286: inst = 32'hc40538b;
      31287: inst = 32'h8220000;
      31288: inst = 32'h10408000;
      31289: inst = 32'hc40538c;
      31290: inst = 32'h8220000;
      31291: inst = 32'h10408000;
      31292: inst = 32'hc40538d;
      31293: inst = 32'h8220000;
      31294: inst = 32'h10408000;
      31295: inst = 32'hc40538e;
      31296: inst = 32'h8220000;
      31297: inst = 32'h10408000;
      31298: inst = 32'hc40538f;
      31299: inst = 32'h8220000;
      31300: inst = 32'h10408000;
      31301: inst = 32'hc405390;
      31302: inst = 32'h8220000;
      31303: inst = 32'h10408000;
      31304: inst = 32'hc405391;
      31305: inst = 32'h8220000;
      31306: inst = 32'h10408000;
      31307: inst = 32'hc405392;
      31308: inst = 32'h8220000;
      31309: inst = 32'h10408000;
      31310: inst = 32'hc405393;
      31311: inst = 32'h8220000;
      31312: inst = 32'h10408000;
      31313: inst = 32'hc405394;
      31314: inst = 32'h8220000;
      31315: inst = 32'h10408000;
      31316: inst = 32'hc405395;
      31317: inst = 32'h8220000;
      31318: inst = 32'h10408000;
      31319: inst = 32'hc405396;
      31320: inst = 32'h8220000;
      31321: inst = 32'h10408000;
      31322: inst = 32'hc405397;
      31323: inst = 32'h8220000;
      31324: inst = 32'h10408000;
      31325: inst = 32'hc405398;
      31326: inst = 32'h8220000;
      31327: inst = 32'h10408000;
      31328: inst = 32'hc405399;
      31329: inst = 32'h8220000;
      31330: inst = 32'h10408000;
      31331: inst = 32'hc40539a;
      31332: inst = 32'h8220000;
      31333: inst = 32'h10408000;
      31334: inst = 32'hc40539b;
      31335: inst = 32'h8220000;
      31336: inst = 32'h10408000;
      31337: inst = 32'hc40539c;
      31338: inst = 32'h8220000;
      31339: inst = 32'h10408000;
      31340: inst = 32'hc40539d;
      31341: inst = 32'h8220000;
      31342: inst = 32'h10408000;
      31343: inst = 32'hc40539e;
      31344: inst = 32'h8220000;
      31345: inst = 32'h10408000;
      31346: inst = 32'hc40539f;
      31347: inst = 32'h8220000;
      31348: inst = 32'h10408000;
      31349: inst = 32'hc4053a0;
      31350: inst = 32'h8220000;
      31351: inst = 32'h10408000;
      31352: inst = 32'hc4053a1;
      31353: inst = 32'h8220000;
      31354: inst = 32'h10408000;
      31355: inst = 32'hc4053a2;
      31356: inst = 32'h8220000;
      31357: inst = 32'h10408000;
      31358: inst = 32'hc4053a3;
      31359: inst = 32'h8220000;
      31360: inst = 32'h10408000;
      31361: inst = 32'hc4053a4;
      31362: inst = 32'h8220000;
      31363: inst = 32'h10408000;
      31364: inst = 32'hc4053a5;
      31365: inst = 32'h8220000;
      31366: inst = 32'h10408000;
      31367: inst = 32'hc4053a6;
      31368: inst = 32'h8220000;
      31369: inst = 32'h10408000;
      31370: inst = 32'hc4053a7;
      31371: inst = 32'h8220000;
      31372: inst = 32'h10408000;
      31373: inst = 32'hc4053a8;
      31374: inst = 32'h8220000;
      31375: inst = 32'h10408000;
      31376: inst = 32'hc4053a9;
      31377: inst = 32'h8220000;
      31378: inst = 32'h10408000;
      31379: inst = 32'hc4053aa;
      31380: inst = 32'h8220000;
      31381: inst = 32'h10408000;
      31382: inst = 32'hc4053ab;
      31383: inst = 32'h8220000;
      31384: inst = 32'h10408000;
      31385: inst = 32'hc4053ac;
      31386: inst = 32'h8220000;
      31387: inst = 32'h10408000;
      31388: inst = 32'hc4053ad;
      31389: inst = 32'h8220000;
      31390: inst = 32'h10408000;
      31391: inst = 32'hc4053ae;
      31392: inst = 32'h8220000;
      31393: inst = 32'h10408000;
      31394: inst = 32'hc4053af;
      31395: inst = 32'h8220000;
      31396: inst = 32'h10408000;
      31397: inst = 32'hc4053b0;
      31398: inst = 32'h8220000;
      31399: inst = 32'h10408000;
      31400: inst = 32'hc4053b1;
      31401: inst = 32'h8220000;
      31402: inst = 32'h10408000;
      31403: inst = 32'hc4053b2;
      31404: inst = 32'h8220000;
      31405: inst = 32'h10408000;
      31406: inst = 32'hc4053b3;
      31407: inst = 32'h8220000;
      31408: inst = 32'h10408000;
      31409: inst = 32'hc4053b4;
      31410: inst = 32'h8220000;
      31411: inst = 32'h10408000;
      31412: inst = 32'hc4053b5;
      31413: inst = 32'h8220000;
      31414: inst = 32'h10408000;
      31415: inst = 32'hc4053b6;
      31416: inst = 32'h8220000;
      31417: inst = 32'h10408000;
      31418: inst = 32'hc4053b7;
      31419: inst = 32'h8220000;
      31420: inst = 32'h10408000;
      31421: inst = 32'hc4053b8;
      31422: inst = 32'h8220000;
      31423: inst = 32'h10408000;
      31424: inst = 32'hc4053c8;
      31425: inst = 32'h8220000;
      31426: inst = 32'h10408000;
      31427: inst = 32'hc4053c9;
      31428: inst = 32'h8220000;
      31429: inst = 32'h10408000;
      31430: inst = 32'hc4053ca;
      31431: inst = 32'h8220000;
      31432: inst = 32'h10408000;
      31433: inst = 32'hc4053cb;
      31434: inst = 32'h8220000;
      31435: inst = 32'h10408000;
      31436: inst = 32'hc4053cc;
      31437: inst = 32'h8220000;
      31438: inst = 32'h10408000;
      31439: inst = 32'hc4053cd;
      31440: inst = 32'h8220000;
      31441: inst = 32'h10408000;
      31442: inst = 32'hc4053ce;
      31443: inst = 32'h8220000;
      31444: inst = 32'h10408000;
      31445: inst = 32'hc4053cf;
      31446: inst = 32'h8220000;
      31447: inst = 32'h10408000;
      31448: inst = 32'hc4053d0;
      31449: inst = 32'h8220000;
      31450: inst = 32'h10408000;
      31451: inst = 32'hc4053d1;
      31452: inst = 32'h8220000;
      31453: inst = 32'h10408000;
      31454: inst = 32'hc4053d2;
      31455: inst = 32'h8220000;
      31456: inst = 32'h10408000;
      31457: inst = 32'hc4053d3;
      31458: inst = 32'h8220000;
      31459: inst = 32'h10408000;
      31460: inst = 32'hc4053d4;
      31461: inst = 32'h8220000;
      31462: inst = 32'h10408000;
      31463: inst = 32'hc4053d5;
      31464: inst = 32'h8220000;
      31465: inst = 32'h10408000;
      31466: inst = 32'hc4053d6;
      31467: inst = 32'h8220000;
      31468: inst = 32'h10408000;
      31469: inst = 32'hc4053d7;
      31470: inst = 32'h8220000;
      31471: inst = 32'h10408000;
      31472: inst = 32'hc4053d8;
      31473: inst = 32'h8220000;
      31474: inst = 32'h10408000;
      31475: inst = 32'hc4053d9;
      31476: inst = 32'h8220000;
      31477: inst = 32'h10408000;
      31478: inst = 32'hc4053da;
      31479: inst = 32'h8220000;
      31480: inst = 32'h10408000;
      31481: inst = 32'hc4053db;
      31482: inst = 32'h8220000;
      31483: inst = 32'h10408000;
      31484: inst = 32'hc4053dc;
      31485: inst = 32'h8220000;
      31486: inst = 32'h10408000;
      31487: inst = 32'hc4053dd;
      31488: inst = 32'h8220000;
      31489: inst = 32'h10408000;
      31490: inst = 32'hc4053de;
      31491: inst = 32'h8220000;
      31492: inst = 32'h10408000;
      31493: inst = 32'hc4053df;
      31494: inst = 32'h8220000;
      31495: inst = 32'h10408000;
      31496: inst = 32'hc4053e0;
      31497: inst = 32'h8220000;
      31498: inst = 32'h10408000;
      31499: inst = 32'hc4053e1;
      31500: inst = 32'h8220000;
      31501: inst = 32'h10408000;
      31502: inst = 32'hc4053e2;
      31503: inst = 32'h8220000;
      31504: inst = 32'h10408000;
      31505: inst = 32'hc4053e3;
      31506: inst = 32'h8220000;
      31507: inst = 32'h10408000;
      31508: inst = 32'hc4053e4;
      31509: inst = 32'h8220000;
      31510: inst = 32'h10408000;
      31511: inst = 32'hc4053e5;
      31512: inst = 32'h8220000;
      31513: inst = 32'h10408000;
      31514: inst = 32'hc4053e6;
      31515: inst = 32'h8220000;
      31516: inst = 32'h10408000;
      31517: inst = 32'hc4053e7;
      31518: inst = 32'h8220000;
      31519: inst = 32'h10408000;
      31520: inst = 32'hc4053e8;
      31521: inst = 32'h8220000;
      31522: inst = 32'h10408000;
      31523: inst = 32'hc4053e9;
      31524: inst = 32'h8220000;
      31525: inst = 32'h10408000;
      31526: inst = 32'hc4053ea;
      31527: inst = 32'h8220000;
      31528: inst = 32'h10408000;
      31529: inst = 32'hc4053eb;
      31530: inst = 32'h8220000;
      31531: inst = 32'h10408000;
      31532: inst = 32'hc4053ec;
      31533: inst = 32'h8220000;
      31534: inst = 32'h10408000;
      31535: inst = 32'hc4053ed;
      31536: inst = 32'h8220000;
      31537: inst = 32'h10408000;
      31538: inst = 32'hc4053ee;
      31539: inst = 32'h8220000;
      31540: inst = 32'h10408000;
      31541: inst = 32'hc4053ef;
      31542: inst = 32'h8220000;
      31543: inst = 32'h10408000;
      31544: inst = 32'hc4053f0;
      31545: inst = 32'h8220000;
      31546: inst = 32'h10408000;
      31547: inst = 32'hc4053f1;
      31548: inst = 32'h8220000;
      31549: inst = 32'h10408000;
      31550: inst = 32'hc4053f2;
      31551: inst = 32'h8220000;
      31552: inst = 32'h10408000;
      31553: inst = 32'hc4053f3;
      31554: inst = 32'h8220000;
      31555: inst = 32'h10408000;
      31556: inst = 32'hc4053f4;
      31557: inst = 32'h8220000;
      31558: inst = 32'h10408000;
      31559: inst = 32'hc4053f5;
      31560: inst = 32'h8220000;
      31561: inst = 32'h10408000;
      31562: inst = 32'hc4053f6;
      31563: inst = 32'h8220000;
      31564: inst = 32'h10408000;
      31565: inst = 32'hc4053f7;
      31566: inst = 32'h8220000;
      31567: inst = 32'h10408000;
      31568: inst = 32'hc4053f8;
      31569: inst = 32'h8220000;
      31570: inst = 32'h10408000;
      31571: inst = 32'hc4053f9;
      31572: inst = 32'h8220000;
      31573: inst = 32'h10408000;
      31574: inst = 32'hc4053fa;
      31575: inst = 32'h8220000;
      31576: inst = 32'h10408000;
      31577: inst = 32'hc4053fb;
      31578: inst = 32'h8220000;
      31579: inst = 32'h10408000;
      31580: inst = 32'hc4053fc;
      31581: inst = 32'h8220000;
      31582: inst = 32'h10408000;
      31583: inst = 32'hc4053fd;
      31584: inst = 32'h8220000;
      31585: inst = 32'h10408000;
      31586: inst = 32'hc4053fe;
      31587: inst = 32'h8220000;
      31588: inst = 32'h10408000;
      31589: inst = 32'hc4053ff;
      31590: inst = 32'h8220000;
      31591: inst = 32'h10408000;
      31592: inst = 32'hc405400;
      31593: inst = 32'h8220000;
      31594: inst = 32'h10408000;
      31595: inst = 32'hc405401;
      31596: inst = 32'h8220000;
      31597: inst = 32'h10408000;
      31598: inst = 32'hc405402;
      31599: inst = 32'h8220000;
      31600: inst = 32'h10408000;
      31601: inst = 32'hc405403;
      31602: inst = 32'h8220000;
      31603: inst = 32'h10408000;
      31604: inst = 32'hc405404;
      31605: inst = 32'h8220000;
      31606: inst = 32'h10408000;
      31607: inst = 32'hc405405;
      31608: inst = 32'h8220000;
      31609: inst = 32'h10408000;
      31610: inst = 32'hc405406;
      31611: inst = 32'h8220000;
      31612: inst = 32'h10408000;
      31613: inst = 32'hc405407;
      31614: inst = 32'h8220000;
      31615: inst = 32'h10408000;
      31616: inst = 32'hc405408;
      31617: inst = 32'h8220000;
      31618: inst = 32'h10408000;
      31619: inst = 32'hc405409;
      31620: inst = 32'h8220000;
      31621: inst = 32'h10408000;
      31622: inst = 32'hc40540a;
      31623: inst = 32'h8220000;
      31624: inst = 32'h10408000;
      31625: inst = 32'hc40540b;
      31626: inst = 32'h8220000;
      31627: inst = 32'h10408000;
      31628: inst = 32'hc40540c;
      31629: inst = 32'h8220000;
      31630: inst = 32'h10408000;
      31631: inst = 32'hc40540d;
      31632: inst = 32'h8220000;
      31633: inst = 32'h10408000;
      31634: inst = 32'hc40540e;
      31635: inst = 32'h8220000;
      31636: inst = 32'h10408000;
      31637: inst = 32'hc40540f;
      31638: inst = 32'h8220000;
      31639: inst = 32'h10408000;
      31640: inst = 32'hc405410;
      31641: inst = 32'h8220000;
      31642: inst = 32'h10408000;
      31643: inst = 32'hc405411;
      31644: inst = 32'h8220000;
      31645: inst = 32'h10408000;
      31646: inst = 32'hc405412;
      31647: inst = 32'h8220000;
      31648: inst = 32'h10408000;
      31649: inst = 32'hc405413;
      31650: inst = 32'h8220000;
      31651: inst = 32'h10408000;
      31652: inst = 32'hc405414;
      31653: inst = 32'h8220000;
      31654: inst = 32'h10408000;
      31655: inst = 32'hc405415;
      31656: inst = 32'h8220000;
      31657: inst = 32'h10408000;
      31658: inst = 32'hc405416;
      31659: inst = 32'h8220000;
      31660: inst = 32'h10408000;
      31661: inst = 32'hc405417;
      31662: inst = 32'h8220000;
      31663: inst = 32'hc20296c;
      31664: inst = 32'h10408000;
      31665: inst = 32'hc404406;
      31666: inst = 32'h8220000;
      31667: inst = 32'h10408000;
      31668: inst = 32'hc404459;
      31669: inst = 32'h8220000;
      31670: inst = 32'h10408000;
      31671: inst = 32'hc404466;
      31672: inst = 32'h8220000;
      31673: inst = 32'h10408000;
      31674: inst = 32'hc4044b9;
      31675: inst = 32'h8220000;
      31676: inst = 32'h10408000;
      31677: inst = 32'hc4044c6;
      31678: inst = 32'h8220000;
      31679: inst = 32'h10408000;
      31680: inst = 32'hc404519;
      31681: inst = 32'h8220000;
      31682: inst = 32'h10408000;
      31683: inst = 32'hc404526;
      31684: inst = 32'h8220000;
      31685: inst = 32'h10408000;
      31686: inst = 32'hc404579;
      31687: inst = 32'h8220000;
      31688: inst = 32'h10408000;
      31689: inst = 32'hc404586;
      31690: inst = 32'h8220000;
      31691: inst = 32'h10408000;
      31692: inst = 32'hc4045d9;
      31693: inst = 32'h8220000;
      31694: inst = 32'h10408000;
      31695: inst = 32'hc4045e6;
      31696: inst = 32'h8220000;
      31697: inst = 32'h10408000;
      31698: inst = 32'hc404639;
      31699: inst = 32'h8220000;
      31700: inst = 32'h10408000;
      31701: inst = 32'hc404646;
      31702: inst = 32'h8220000;
      31703: inst = 32'h10408000;
      31704: inst = 32'hc404699;
      31705: inst = 32'h8220000;
      31706: inst = 32'h10408000;
      31707: inst = 32'hc4046a6;
      31708: inst = 32'h8220000;
      31709: inst = 32'h10408000;
      31710: inst = 32'hc4046f9;
      31711: inst = 32'h8220000;
      31712: inst = 32'h10408000;
      31713: inst = 32'hc404706;
      31714: inst = 32'h8220000;
      31715: inst = 32'h10408000;
      31716: inst = 32'hc404759;
      31717: inst = 32'h8220000;
      31718: inst = 32'h10408000;
      31719: inst = 32'hc404766;
      31720: inst = 32'h8220000;
      31721: inst = 32'h10408000;
      31722: inst = 32'hc4047b9;
      31723: inst = 32'h8220000;
      31724: inst = 32'h10408000;
      31725: inst = 32'hc4047c6;
      31726: inst = 32'h8220000;
      31727: inst = 32'h10408000;
      31728: inst = 32'hc404819;
      31729: inst = 32'h8220000;
      31730: inst = 32'h10408000;
      31731: inst = 32'hc404826;
      31732: inst = 32'h8220000;
      31733: inst = 32'h10408000;
      31734: inst = 32'hc404879;
      31735: inst = 32'h8220000;
      31736: inst = 32'h10408000;
      31737: inst = 32'hc404886;
      31738: inst = 32'h8220000;
      31739: inst = 32'h10408000;
      31740: inst = 32'hc4048d9;
      31741: inst = 32'h8220000;
      31742: inst = 32'h10408000;
      31743: inst = 32'hc4048e6;
      31744: inst = 32'h8220000;
      31745: inst = 32'h10408000;
      31746: inst = 32'hc404939;
      31747: inst = 32'h8220000;
      31748: inst = 32'h10408000;
      31749: inst = 32'hc404946;
      31750: inst = 32'h8220000;
      31751: inst = 32'h10408000;
      31752: inst = 32'hc404999;
      31753: inst = 32'h8220000;
      31754: inst = 32'h10408000;
      31755: inst = 32'hc4049a6;
      31756: inst = 32'h8220000;
      31757: inst = 32'h10408000;
      31758: inst = 32'hc4049f9;
      31759: inst = 32'h8220000;
      31760: inst = 32'h10408000;
      31761: inst = 32'hc404a06;
      31762: inst = 32'h8220000;
      31763: inst = 32'h10408000;
      31764: inst = 32'hc404a59;
      31765: inst = 32'h8220000;
      31766: inst = 32'h10408000;
      31767: inst = 32'hc404a66;
      31768: inst = 32'h8220000;
      31769: inst = 32'h10408000;
      31770: inst = 32'hc404ab9;
      31771: inst = 32'h8220000;
      31772: inst = 32'h10408000;
      31773: inst = 32'hc404ac6;
      31774: inst = 32'h8220000;
      31775: inst = 32'h10408000;
      31776: inst = 32'hc404b19;
      31777: inst = 32'h8220000;
      31778: inst = 32'h10408000;
      31779: inst = 32'hc404b26;
      31780: inst = 32'h8220000;
      31781: inst = 32'h10408000;
      31782: inst = 32'hc404b79;
      31783: inst = 32'h8220000;
      31784: inst = 32'h10408000;
      31785: inst = 32'hc404b86;
      31786: inst = 32'h8220000;
      31787: inst = 32'h10408000;
      31788: inst = 32'hc404bd9;
      31789: inst = 32'h8220000;
      31790: inst = 32'h10408000;
      31791: inst = 32'hc404be6;
      31792: inst = 32'h8220000;
      31793: inst = 32'h10408000;
      31794: inst = 32'hc404c39;
      31795: inst = 32'h8220000;
      31796: inst = 32'h10408000;
      31797: inst = 32'hc404c46;
      31798: inst = 32'h8220000;
      31799: inst = 32'h10408000;
      31800: inst = 32'hc404c99;
      31801: inst = 32'h8220000;
      31802: inst = 32'h10408000;
      31803: inst = 32'hc404ca6;
      31804: inst = 32'h8220000;
      31805: inst = 32'h10408000;
      31806: inst = 32'hc404cf9;
      31807: inst = 32'h8220000;
      31808: inst = 32'h10408000;
      31809: inst = 32'hc404d06;
      31810: inst = 32'h8220000;
      31811: inst = 32'h10408000;
      31812: inst = 32'hc404d59;
      31813: inst = 32'h8220000;
      31814: inst = 32'h10408000;
      31815: inst = 32'hc404d66;
      31816: inst = 32'h8220000;
      31817: inst = 32'h10408000;
      31818: inst = 32'hc404db9;
      31819: inst = 32'h8220000;
      31820: inst = 32'h10408000;
      31821: inst = 32'hc404dc6;
      31822: inst = 32'h8220000;
      31823: inst = 32'h10408000;
      31824: inst = 32'hc404e19;
      31825: inst = 32'h8220000;
      31826: inst = 32'h10408000;
      31827: inst = 32'hc404e26;
      31828: inst = 32'h8220000;
      31829: inst = 32'h10408000;
      31830: inst = 32'hc404e79;
      31831: inst = 32'h8220000;
      31832: inst = 32'h10408000;
      31833: inst = 32'hc404e86;
      31834: inst = 32'h8220000;
      31835: inst = 32'h10408000;
      31836: inst = 32'hc404ed9;
      31837: inst = 32'h8220000;
      31838: inst = 32'h10408000;
      31839: inst = 32'hc404ee6;
      31840: inst = 32'h8220000;
      31841: inst = 32'h10408000;
      31842: inst = 32'hc404f39;
      31843: inst = 32'h8220000;
      31844: inst = 32'h10408000;
      31845: inst = 32'hc404f46;
      31846: inst = 32'h8220000;
      31847: inst = 32'h10408000;
      31848: inst = 32'hc404f99;
      31849: inst = 32'h8220000;
      31850: inst = 32'h10408000;
      31851: inst = 32'hc404fa6;
      31852: inst = 32'h8220000;
      31853: inst = 32'h10408000;
      31854: inst = 32'hc404ff9;
      31855: inst = 32'h8220000;
      31856: inst = 32'h10408000;
      31857: inst = 32'hc405006;
      31858: inst = 32'h8220000;
      31859: inst = 32'h10408000;
      31860: inst = 32'hc405059;
      31861: inst = 32'h8220000;
      31862: inst = 32'h10408000;
      31863: inst = 32'hc405066;
      31864: inst = 32'h8220000;
      31865: inst = 32'h10408000;
      31866: inst = 32'hc4050b9;
      31867: inst = 32'h8220000;
      31868: inst = 32'h10408000;
      31869: inst = 32'hc4050c6;
      31870: inst = 32'h8220000;
      31871: inst = 32'h10408000;
      31872: inst = 32'hc405119;
      31873: inst = 32'h8220000;
      31874: inst = 32'h10408000;
      31875: inst = 32'hc405126;
      31876: inst = 32'h8220000;
      31877: inst = 32'h10408000;
      31878: inst = 32'hc405179;
      31879: inst = 32'h8220000;
      31880: inst = 32'h10408000;
      31881: inst = 32'hc405186;
      31882: inst = 32'h8220000;
      31883: inst = 32'h10408000;
      31884: inst = 32'hc4051d9;
      31885: inst = 32'h8220000;
      31886: inst = 32'h10408000;
      31887: inst = 32'hc4051e6;
      31888: inst = 32'h8220000;
      31889: inst = 32'h10408000;
      31890: inst = 32'hc405239;
      31891: inst = 32'h8220000;
      31892: inst = 32'h10408000;
      31893: inst = 32'hc405246;
      31894: inst = 32'h8220000;
      31895: inst = 32'h10408000;
      31896: inst = 32'hc405299;
      31897: inst = 32'h8220000;
      31898: inst = 32'h10408000;
      31899: inst = 32'hc4052a6;
      31900: inst = 32'h8220000;
      31901: inst = 32'h10408000;
      31902: inst = 32'hc4052f9;
      31903: inst = 32'h8220000;
      31904: inst = 32'h10408000;
      31905: inst = 32'hc405306;
      31906: inst = 32'h8220000;
      31907: inst = 32'h10408000;
      31908: inst = 32'hc405359;
      31909: inst = 32'h8220000;
      31910: inst = 32'hc20738e;
      31911: inst = 32'h10408000;
      31912: inst = 32'hc40464e;
      31913: inst = 32'h8220000;
      31914: inst = 32'h10408000;
      31915: inst = 32'hc404690;
      31916: inst = 32'h8220000;
      31917: inst = 32'h10408000;
      31918: inst = 32'hc4046ae;
      31919: inst = 32'h8220000;
      31920: inst = 32'h10408000;
      31921: inst = 32'hc4046f0;
      31922: inst = 32'h8220000;
      31923: inst = 32'h10408000;
      31924: inst = 32'hc4047d3;
      31925: inst = 32'h8220000;
      31926: inst = 32'h10408000;
      31927: inst = 32'hc4047dd;
      31928: inst = 32'h8220000;
      31929: inst = 32'h10408000;
      31930: inst = 32'hc404800;
      31931: inst = 32'h8220000;
      31932: inst = 32'h10408000;
      31933: inst = 32'hc40483a;
      31934: inst = 32'h8220000;
      31935: inst = 32'h10408000;
      31936: inst = 32'hc40485d;
      31937: inst = 32'h8220000;
      31938: inst = 32'h10408000;
      31939: inst = 32'hc4049b8;
      31940: inst = 32'h8220000;
      31941: inst = 32'h10408000;
      31942: inst = 32'hc4049c7;
      31943: inst = 32'h8220000;
      31944: inst = 32'h10408000;
      31945: inst = 32'hc4049e5;
      31946: inst = 32'h8220000;
      31947: inst = 32'h10408000;
      31948: inst = 32'hc4049f0;
      31949: inst = 32'h8220000;
      31950: inst = 32'h10408000;
      31951: inst = 32'hc404cb1;
      31952: inst = 32'h8220000;
      31953: inst = 32'h10408000;
      31954: inst = 32'hc404cf2;
      31955: inst = 32'h8220000;
      31956: inst = 32'h10408000;
      31957: inst = 32'hc404dda;
      31958: inst = 32'h8220000;
      31959: inst = 32'h10408000;
      31960: inst = 32'hc404e5c;
      31961: inst = 32'h8220000;
      31962: inst = 32'h10408000;
      31963: inst = 32'hc404e6b;
      31964: inst = 32'h8220000;
      31965: inst = 32'h10408000;
      31966: inst = 32'hc404e96;
      31967: inst = 32'h8220000;
      31968: inst = 32'h10408000;
      31969: inst = 32'hc404eaf;
      31970: inst = 32'h8220000;
      31971: inst = 32'h10408000;
      31972: inst = 32'hc404fb6;
      31973: inst = 32'h8220000;
      31974: inst = 32'h10408000;
      31975: inst = 32'hc404fcf;
      31976: inst = 32'h8220000;
      31977: inst = 32'h10408000;
      31978: inst = 32'hc40501a;
      31979: inst = 32'h8220000;
      31980: inst = 32'hc20ad75;
      31981: inst = 32'h10408000;
      31982: inst = 32'hc40464f;
      31983: inst = 32'h8220000;
      31984: inst = 32'h10408000;
      31985: inst = 32'hc404692;
      31986: inst = 32'h8220000;
      31987: inst = 32'h10408000;
      31988: inst = 32'hc404809;
      31989: inst = 32'h8220000;
      31990: inst = 32'h10408000;
      31991: inst = 32'hc40483d;
      31992: inst = 32'h8220000;
      31993: inst = 32'h10408000;
      31994: inst = 32'hc404860;
      31995: inst = 32'h8220000;
      31996: inst = 32'h10408000;
      31997: inst = 32'hc404e58;
      31998: inst = 32'h8220000;
      31999: inst = 32'h10408000;
      32000: inst = 32'hc404e59;
      32001: inst = 32'h8220000;
      32002: inst = 32'h10408000;
      32003: inst = 32'hc404e67;
      32004: inst = 32'h8220000;
      32005: inst = 32'h10408000;
      32006: inst = 32'hc404e68;
      32007: inst = 32'h8220000;
      32008: inst = 32'h10408000;
      32009: inst = 32'hc404f19;
      32010: inst = 32'h8220000;
      32011: inst = 32'h10408000;
      32012: inst = 32'hc404f28;
      32013: inst = 32'h8220000;
      32014: inst = 32'h10408000;
      32015: inst = 32'hc404f4f;
      32016: inst = 32'h8220000;
      32017: inst = 32'h10408000;
      32018: inst = 32'hc404fc3;
      32019: inst = 32'h8220000;
      32020: inst = 32'h10408000;
      32021: inst = 32'hc404fcd;
      32022: inst = 32'h8220000;
      32023: inst = 32'h10408000;
      32024: inst = 32'hc404fe1;
      32025: inst = 32'h8220000;
      32026: inst = 32'h10408000;
      32027: inst = 32'hc404ff0;
      32028: inst = 32'h8220000;
      32029: inst = 32'h10408000;
      32030: inst = 32'hc40500e;
      32031: inst = 32'h8220000;
      32032: inst = 32'h10408000;
      32033: inst = 32'hc405054;
      32034: inst = 32'h8220000;
      32035: inst = 32'hc2031a6;
      32036: inst = 32'h10408000;
      32037: inst = 32'hc404650;
      32038: inst = 32'h8220000;
      32039: inst = 32'h10408000;
      32040: inst = 32'hc404772;
      32041: inst = 32'h8220000;
      32042: inst = 32'h10408000;
      32043: inst = 32'hc40477a;
      32044: inst = 32'h8220000;
      32045: inst = 32'h10408000;
      32046: inst = 32'hc40478b;
      32047: inst = 32'h8220000;
      32048: inst = 32'h10408000;
      32049: inst = 32'hc404793;
      32050: inst = 32'h8220000;
      32051: inst = 32'h10408000;
      32052: inst = 32'hc404795;
      32053: inst = 32'h8220000;
      32054: inst = 32'h10408000;
      32055: inst = 32'hc40479a;
      32056: inst = 32'h8220000;
      32057: inst = 32'h10408000;
      32058: inst = 32'hc40479d;
      32059: inst = 32'h8220000;
      32060: inst = 32'h10408000;
      32061: inst = 32'hc4047ae;
      32062: inst = 32'h8220000;
      32063: inst = 32'h10408000;
      32064: inst = 32'hc404847;
      32065: inst = 32'h8220000;
      32066: inst = 32'h10408000;
      32067: inst = 32'hc404971;
      32068: inst = 32'h8220000;
      32069: inst = 32'h10408000;
      32070: inst = 32'hc40498a;
      32071: inst = 32'h8220000;
      32072: inst = 32'h10408000;
      32073: inst = 32'hc404a10;
      32074: inst = 32'h8220000;
      32075: inst = 32'h10408000;
      32076: inst = 32'hc404a18;
      32077: inst = 32'h8220000;
      32078: inst = 32'h10408000;
      32079: inst = 32'hc404a35;
      32080: inst = 32'h8220000;
      32081: inst = 32'h10408000;
      32082: inst = 32'hc404a3b;
      32083: inst = 32'h8220000;
      32084: inst = 32'h10408000;
      32085: inst = 32'hc404a45;
      32086: inst = 32'h8220000;
      32087: inst = 32'h10408000;
      32088: inst = 32'hc404a50;
      32089: inst = 32'h8220000;
      32090: inst = 32'h10408000;
      32091: inst = 32'hc404d21;
      32092: inst = 32'h8220000;
      32093: inst = 32'h10408000;
      32094: inst = 32'hc404d2b;
      32095: inst = 32'h8220000;
      32096: inst = 32'h10408000;
      32097: inst = 32'hc404d3f;
      32098: inst = 32'h8220000;
      32099: inst = 32'h10408000;
      32100: inst = 32'hc404d44;
      32101: inst = 32'h8220000;
      32102: inst = 32'h10408000;
      32103: inst = 32'hc404dcc;
      32104: inst = 32'h8220000;
      32105: inst = 32'h10408000;
      32106: inst = 32'hc404dcf;
      32107: inst = 32'h8220000;
      32108: inst = 32'h10408000;
      32109: inst = 32'hc404dd6;
      32110: inst = 32'h8220000;
      32111: inst = 32'h10408000;
      32112: inst = 32'hc404def;
      32113: inst = 32'h8220000;
      32114: inst = 32'h10408000;
      32115: inst = 32'hc404e98;
      32116: inst = 32'h8220000;
      32117: inst = 32'h10408000;
      32118: inst = 32'hc404eb1;
      32119: inst = 32'h8220000;
      32120: inst = 32'h10408000;
      32121: inst = 32'hc404fac;
      32122: inst = 32'h8220000;
      32123: inst = 32'h10408000;
      32124: inst = 32'hc404fb8;
      32125: inst = 32'h8220000;
      32126: inst = 32'h10408000;
      32127: inst = 32'hc404fd1;
      32128: inst = 32'h8220000;
      32129: inst = 32'h10408000;
      32130: inst = 32'hc404fd3;
      32131: inst = 32'h8220000;
      32132: inst = 32'h10408000;
      32133: inst = 32'hc40506b;
      32134: inst = 32'h8220000;
      32135: inst = 32'h10408000;
      32136: inst = 32'hc405076;
      32137: inst = 32'h8220000;
      32138: inst = 32'h10408000;
      32139: inst = 32'hc405078;
      32140: inst = 32'h8220000;
      32141: inst = 32'h10408000;
      32142: inst = 32'hc405081;
      32143: inst = 32'h8220000;
      32144: inst = 32'h10408000;
      32145: inst = 32'hc40508b;
      32146: inst = 32'h8220000;
      32147: inst = 32'h10408000;
      32148: inst = 32'hc40508f;
      32149: inst = 32'h8220000;
      32150: inst = 32'h10408000;
      32151: inst = 32'hc405091;
      32152: inst = 32'h8220000;
      32153: inst = 32'h10408000;
      32154: inst = 32'hc40509f;
      32155: inst = 32'h8220000;
      32156: inst = 32'h10408000;
      32157: inst = 32'hc4050a4;
      32158: inst = 32'h8220000;
      32159: inst = 32'h10408000;
      32160: inst = 32'hc4050ad;
      32161: inst = 32'h8220000;
      32162: inst = 32'hc20a514;
      32163: inst = 32'h10408000;
      32164: inst = 32'hc404691;
      32165: inst = 32'h8220000;
      32166: inst = 32'h10408000;
      32167: inst = 32'hc4046f1;
      32168: inst = 32'h8220000;
      32169: inst = 32'h10408000;
      32170: inst = 32'hc404715;
      32171: inst = 32'h8220000;
      32172: inst = 32'h10408000;
      32173: inst = 32'hc404716;
      32174: inst = 32'h8220000;
      32175: inst = 32'h10408000;
      32176: inst = 32'hc404724;
      32177: inst = 32'h8220000;
      32178: inst = 32'h10408000;
      32179: inst = 32'hc404725;
      32180: inst = 32'h8220000;
      32181: inst = 32'h10408000;
      32182: inst = 32'hc404742;
      32183: inst = 32'h8220000;
      32184: inst = 32'h10408000;
      32185: inst = 32'hc404743;
      32186: inst = 32'h8220000;
      32187: inst = 32'h10408000;
      32188: inst = 32'hc404776;
      32189: inst = 32'h8220000;
      32190: inst = 32'h10408000;
      32191: inst = 32'hc404785;
      32192: inst = 32'h8220000;
      32193: inst = 32'h10408000;
      32194: inst = 32'hc4047a3;
      32195: inst = 32'h8220000;
      32196: inst = 32'h10408000;
      32197: inst = 32'hc4047d4;
      32198: inst = 32'h8220000;
      32199: inst = 32'h10408000;
      32200: inst = 32'hc4047d7;
      32201: inst = 32'h8220000;
      32202: inst = 32'h10408000;
      32203: inst = 32'hc4047db;
      32204: inst = 32'h8220000;
      32205: inst = 32'h10408000;
      32206: inst = 32'hc4047e3;
      32207: inst = 32'h8220000;
      32208: inst = 32'h10408000;
      32209: inst = 32'hc4047e6;
      32210: inst = 32'h8220000;
      32211: inst = 32'h10408000;
      32212: inst = 32'hc4047ea;
      32213: inst = 32'h8220000;
      32214: inst = 32'h10408000;
      32215: inst = 32'hc4047f4;
      32216: inst = 32'h8220000;
      32217: inst = 32'h10408000;
      32218: inst = 32'hc4047f9;
      32219: inst = 32'h8220000;
      32220: inst = 32'h10408000;
      32221: inst = 32'hc4047fe;
      32222: inst = 32'h8220000;
      32223: inst = 32'h10408000;
      32224: inst = 32'hc404801;
      32225: inst = 32'h8220000;
      32226: inst = 32'h10408000;
      32227: inst = 32'hc404804;
      32228: inst = 32'h8220000;
      32229: inst = 32'h10408000;
      32230: inst = 32'hc404806;
      32231: inst = 32'h8220000;
      32232: inst = 32'h10408000;
      32233: inst = 32'hc404808;
      32234: inst = 32'h8220000;
      32235: inst = 32'h10408000;
      32236: inst = 32'hc40480d;
      32237: inst = 32'h8220000;
      32238: inst = 32'h10408000;
      32239: inst = 32'hc404836;
      32240: inst = 32'h8220000;
      32241: inst = 32'h10408000;
      32242: inst = 32'hc40483c;
      32243: inst = 32'h8220000;
      32244: inst = 32'h10408000;
      32245: inst = 32'hc404845;
      32246: inst = 32'h8220000;
      32247: inst = 32'h10408000;
      32248: inst = 32'hc404856;
      32249: inst = 32'h8220000;
      32250: inst = 32'h10408000;
      32251: inst = 32'hc40485f;
      32252: inst = 32'h8220000;
      32253: inst = 32'h10408000;
      32254: inst = 32'hc404863;
      32255: inst = 32'h8220000;
      32256: inst = 32'h10408000;
      32257: inst = 32'hc40486a;
      32258: inst = 32'h8220000;
      32259: inst = 32'h10408000;
      32260: inst = 32'hc404896;
      32261: inst = 32'h8220000;
      32262: inst = 32'h10408000;
      32263: inst = 32'hc40489c;
      32264: inst = 32'h8220000;
      32265: inst = 32'h10408000;
      32266: inst = 32'hc4048a5;
      32267: inst = 32'h8220000;
      32268: inst = 32'h10408000;
      32269: inst = 32'hc4048bf;
      32270: inst = 32'h8220000;
      32271: inst = 32'h10408000;
      32272: inst = 32'hc4048c3;
      32273: inst = 32'h8220000;
      32274: inst = 32'h10408000;
      32275: inst = 32'hc4048f6;
      32276: inst = 32'h8220000;
      32277: inst = 32'h10408000;
      32278: inst = 32'hc4048fc;
      32279: inst = 32'h8220000;
      32280: inst = 32'h10408000;
      32281: inst = 32'hc404905;
      32282: inst = 32'h8220000;
      32283: inst = 32'h10408000;
      32284: inst = 32'hc40491f;
      32285: inst = 32'h8220000;
      32286: inst = 32'h10408000;
      32287: inst = 32'hc404923;
      32288: inst = 32'h8220000;
      32289: inst = 32'h10408000;
      32290: inst = 32'hc404956;
      32291: inst = 32'h8220000;
      32292: inst = 32'h10408000;
      32293: inst = 32'hc404958;
      32294: inst = 32'h8220000;
      32295: inst = 32'h10408000;
      32296: inst = 32'hc40495c;
      32297: inst = 32'h8220000;
      32298: inst = 32'h10408000;
      32299: inst = 32'hc404965;
      32300: inst = 32'h8220000;
      32301: inst = 32'h10408000;
      32302: inst = 32'hc404967;
      32303: inst = 32'h8220000;
      32304: inst = 32'h10408000;
      32305: inst = 32'hc404976;
      32306: inst = 32'h8220000;
      32307: inst = 32'h10408000;
      32308: inst = 32'hc40497f;
      32309: inst = 32'h8220000;
      32310: inst = 32'h10408000;
      32311: inst = 32'hc404983;
      32312: inst = 32'h8220000;
      32313: inst = 32'h10408000;
      32314: inst = 32'hc404985;
      32315: inst = 32'h8220000;
      32316: inst = 32'h10408000;
      32317: inst = 32'hc4049b1;
      32318: inst = 32'h8220000;
      32319: inst = 32'h10408000;
      32320: inst = 32'hc4049b5;
      32321: inst = 32'h8220000;
      32322: inst = 32'h10408000;
      32323: inst = 32'hc4049ba;
      32324: inst = 32'h8220000;
      32325: inst = 32'h10408000;
      32326: inst = 32'hc4049c4;
      32327: inst = 32'h8220000;
      32328: inst = 32'h10408000;
      32329: inst = 32'hc4049ca;
      32330: inst = 32'h8220000;
      32331: inst = 32'h10408000;
      32332: inst = 32'hc4049d4;
      32333: inst = 32'h8220000;
      32334: inst = 32'h10408000;
      32335: inst = 32'hc4049d9;
      32336: inst = 32'h8220000;
      32337: inst = 32'h10408000;
      32338: inst = 32'hc4049dd;
      32339: inst = 32'h8220000;
      32340: inst = 32'h10408000;
      32341: inst = 32'hc4049e2;
      32342: inst = 32'h8220000;
      32343: inst = 32'h10408000;
      32344: inst = 32'hc4049e6;
      32345: inst = 32'h8220000;
      32346: inst = 32'h10408000;
      32347: inst = 32'hc4049e8;
      32348: inst = 32'h8220000;
      32349: inst = 32'h10408000;
      32350: inst = 32'hc4049ed;
      32351: inst = 32'h8220000;
      32352: inst = 32'h10408000;
      32353: inst = 32'hc4049f1;
      32354: inst = 32'h8220000;
      32355: inst = 32'h10408000;
      32356: inst = 32'hc4049f3;
      32357: inst = 32'h8220000;
      32358: inst = 32'h10408000;
      32359: inst = 32'hc404cb0;
      32360: inst = 32'h8220000;
      32361: inst = 32'h10408000;
      32362: inst = 32'hc404cf1;
      32363: inst = 32'h8220000;
      32364: inst = 32'h10408000;
      32365: inst = 32'hc404d11;
      32366: inst = 32'h8220000;
      32367: inst = 32'h10408000;
      32368: inst = 32'hc404d52;
      32369: inst = 32'h8220000;
      32370: inst = 32'h10408000;
      32371: inst = 32'hc404d71;
      32372: inst = 32'h8220000;
      32373: inst = 32'h10408000;
      32374: inst = 32'hc404db2;
      32375: inst = 32'h8220000;
      32376: inst = 32'h10408000;
      32377: inst = 32'hc404dd1;
      32378: inst = 32'h8220000;
      32379: inst = 32'h10408000;
      32380: inst = 32'hc404e12;
      32381: inst = 32'h8220000;
      32382: inst = 32'h10408000;
      32383: inst = 32'hc404e2d;
      32384: inst = 32'h8220000;
      32385: inst = 32'h10408000;
      32386: inst = 32'hc404e34;
      32387: inst = 32'h8220000;
      32388: inst = 32'h10408000;
      32389: inst = 32'hc404e37;
      32390: inst = 32'h8220000;
      32391: inst = 32'h10408000;
      32392: inst = 32'hc404e39;
      32393: inst = 32'h8220000;
      32394: inst = 32'h10408000;
      32395: inst = 32'hc404e3b;
      32396: inst = 32'h8220000;
      32397: inst = 32'h10408000;
      32398: inst = 32'hc404e3d;
      32399: inst = 32'h8220000;
      32400: inst = 32'h10408000;
      32401: inst = 32'hc404e42;
      32402: inst = 32'h8220000;
      32403: inst = 32'h10408000;
      32404: inst = 32'hc404e4c;
      32405: inst = 32'h8220000;
      32406: inst = 32'h10408000;
      32407: inst = 32'hc404e50;
      32408: inst = 32'h8220000;
      32409: inst = 32'h10408000;
      32410: inst = 32'hc404e5a;
      32411: inst = 32'h8220000;
      32412: inst = 32'h10408000;
      32413: inst = 32'hc404e60;
      32414: inst = 32'h8220000;
      32415: inst = 32'h10408000;
      32416: inst = 32'hc404e65;
      32417: inst = 32'h8220000;
      32418: inst = 32'h10408000;
      32419: inst = 32'hc404e69;
      32420: inst = 32'h8220000;
      32421: inst = 32'h10408000;
      32422: inst = 32'hc404e6e;
      32423: inst = 32'h8220000;
      32424: inst = 32'h10408000;
      32425: inst = 32'hc404e70;
      32426: inst = 32'h8220000;
      32427: inst = 32'h10408000;
      32428: inst = 32'hc404e72;
      32429: inst = 32'h8220000;
      32430: inst = 32'h10408000;
      32431: inst = 32'hc404e75;
      32432: inst = 32'h8220000;
      32433: inst = 32'h10408000;
      32434: inst = 32'hc404e8b;
      32435: inst = 32'h8220000;
      32436: inst = 32'h10408000;
      32437: inst = 32'hc404e8c;
      32438: inst = 32'h8220000;
      32439: inst = 32'h10408000;
      32440: inst = 32'hc404e91;
      32441: inst = 32'h8220000;
      32442: inst = 32'h10408000;
      32443: inst = 32'hc404e9b;
      32444: inst = 32'h8220000;
      32445: inst = 32'h10408000;
      32446: inst = 32'hc404ea0;
      32447: inst = 32'h8220000;
      32448: inst = 32'h10408000;
      32449: inst = 32'hc404eaa;
      32450: inst = 32'h8220000;
      32451: inst = 32'h10408000;
      32452: inst = 32'hc404ebb;
      32453: inst = 32'h8220000;
      32454: inst = 32'h10408000;
      32455: inst = 32'hc404ebe;
      32456: inst = 32'h8220000;
      32457: inst = 32'h10408000;
      32458: inst = 32'hc404ec3;
      32459: inst = 32'h8220000;
      32460: inst = 32'h10408000;
      32461: inst = 32'hc404eca;
      32462: inst = 32'h8220000;
      32463: inst = 32'h10408000;
      32464: inst = 32'hc404ecd;
      32465: inst = 32'h8220000;
      32466: inst = 32'h10408000;
      32467: inst = 32'hc404ed2;
      32468: inst = 32'h8220000;
      32469: inst = 32'h10408000;
      32470: inst = 32'hc404ed3;
      32471: inst = 32'h8220000;
      32472: inst = 32'h10408000;
      32473: inst = 32'hc404ed4;
      32474: inst = 32'h8220000;
      32475: inst = 32'h10408000;
      32476: inst = 32'hc404ef1;
      32477: inst = 32'h8220000;
      32478: inst = 32'h10408000;
      32479: inst = 32'hc404efb;
      32480: inst = 32'h8220000;
      32481: inst = 32'h10408000;
      32482: inst = 32'hc404f00;
      32483: inst = 32'h8220000;
      32484: inst = 32'h10408000;
      32485: inst = 32'hc404f0a;
      32486: inst = 32'h8220000;
      32487: inst = 32'h10408000;
      32488: inst = 32'hc404f1e;
      32489: inst = 32'h8220000;
      32490: inst = 32'h10408000;
      32491: inst = 32'hc404f23;
      32492: inst = 32'h8220000;
      32493: inst = 32'h10408000;
      32494: inst = 32'hc404f4d;
      32495: inst = 32'h8220000;
      32496: inst = 32'h10408000;
      32497: inst = 32'hc404f51;
      32498: inst = 32'h8220000;
      32499: inst = 32'h10408000;
      32500: inst = 32'hc404f5b;
      32501: inst = 32'h8220000;
      32502: inst = 32'h10408000;
      32503: inst = 32'hc404f60;
      32504: inst = 32'h8220000;
      32505: inst = 32'h10408000;
      32506: inst = 32'hc404f6a;
      32507: inst = 32'h8220000;
      32508: inst = 32'h10408000;
      32509: inst = 32'hc404f7b;
      32510: inst = 32'h8220000;
      32511: inst = 32'h10408000;
      32512: inst = 32'hc404f7e;
      32513: inst = 32'h8220000;
      32514: inst = 32'h10408000;
      32515: inst = 32'hc404f83;
      32516: inst = 32'h8220000;
      32517: inst = 32'h10408000;
      32518: inst = 32'hc404f8a;
      32519: inst = 32'h8220000;
      32520: inst = 32'h10408000;
      32521: inst = 32'hc404f93;
      32522: inst = 32'h8220000;
      32523: inst = 32'h10408000;
      32524: inst = 32'hc404fb1;
      32525: inst = 32'h8220000;
      32526: inst = 32'h10408000;
      32527: inst = 32'hc404fbb;
      32528: inst = 32'h8220000;
      32529: inst = 32'h10408000;
      32530: inst = 32'hc404fbd;
      32531: inst = 32'h8220000;
      32532: inst = 32'h10408000;
      32533: inst = 32'hc404fc0;
      32534: inst = 32'h8220000;
      32535: inst = 32'h10408000;
      32536: inst = 32'hc404fca;
      32537: inst = 32'h8220000;
      32538: inst = 32'h10408000;
      32539: inst = 32'hc404fdb;
      32540: inst = 32'h8220000;
      32541: inst = 32'h10408000;
      32542: inst = 32'hc404fde;
      32543: inst = 32'h8220000;
      32544: inst = 32'h10408000;
      32545: inst = 32'hc404fe3;
      32546: inst = 32'h8220000;
      32547: inst = 32'h10408000;
      32548: inst = 32'hc404fea;
      32549: inst = 32'h8220000;
      32550: inst = 32'h10408000;
      32551: inst = 32'hc404ff2;
      32552: inst = 32'h8220000;
      32553: inst = 32'h10408000;
      32554: inst = 32'hc40500d;
      32555: inst = 32'h8220000;
      32556: inst = 32'h10408000;
      32557: inst = 32'hc40500f;
      32558: inst = 32'h8220000;
      32559: inst = 32'h10408000;
      32560: inst = 32'hc405013;
      32561: inst = 32'h8220000;
      32562: inst = 32'h10408000;
      32563: inst = 32'hc405017;
      32564: inst = 32'h8220000;
      32565: inst = 32'h10408000;
      32566: inst = 32'hc405023;
      32567: inst = 32'h8220000;
      32568: inst = 32'h10408000;
      32569: inst = 32'hc40502d;
      32570: inst = 32'h8220000;
      32571: inst = 32'h10408000;
      32572: inst = 32'hc405030;
      32573: inst = 32'h8220000;
      32574: inst = 32'h10408000;
      32575: inst = 32'hc40503a;
      32576: inst = 32'h8220000;
      32577: inst = 32'h10408000;
      32578: inst = 32'hc40503d;
      32579: inst = 32'h8220000;
      32580: inst = 32'h10408000;
      32581: inst = 32'hc405041;
      32582: inst = 32'h8220000;
      32583: inst = 32'h10408000;
      32584: inst = 32'hc405046;
      32585: inst = 32'h8220000;
      32586: inst = 32'h10408000;
      32587: inst = 32'hc405049;
      32588: inst = 32'h8220000;
      32589: inst = 32'h10408000;
      32590: inst = 32'hc40504c;
      32591: inst = 32'h8220000;
      32592: inst = 32'h10408000;
      32593: inst = 32'hc40504e;
      32594: inst = 32'h8220000;
      32595: inst = 32'hc20f7be;
      32596: inst = 32'h10408000;
      32597: inst = 32'hc4046af;
      32598: inst = 32'h8220000;
      32599: inst = 32'h10408000;
      32600: inst = 32'hc4046f2;
      32601: inst = 32'h8220000;
      32602: inst = 32'h10408000;
      32603: inst = 32'hc40470f;
      32604: inst = 32'h8220000;
      32605: inst = 32'h10408000;
      32606: inst = 32'hc404752;
      32607: inst = 32'h8220000;
      32608: inst = 32'h10408000;
      32609: inst = 32'hc40476f;
      32610: inst = 32'h8220000;
      32611: inst = 32'h10408000;
      32612: inst = 32'hc4047b2;
      32613: inst = 32'h8220000;
      32614: inst = 32'h10408000;
      32615: inst = 32'hc4047cf;
      32616: inst = 32'h8220000;
      32617: inst = 32'h10408000;
      32618: inst = 32'hc4047d9;
      32619: inst = 32'h8220000;
      32620: inst = 32'h10408000;
      32621: inst = 32'hc4047fc;
      32622: inst = 32'h8220000;
      32623: inst = 32'h10408000;
      32624: inst = 32'hc404807;
      32625: inst = 32'h8220000;
      32626: inst = 32'h10408000;
      32627: inst = 32'hc40480a;
      32628: inst = 32'h8220000;
      32629: inst = 32'h10408000;
      32630: inst = 32'hc404812;
      32631: inst = 32'h8220000;
      32632: inst = 32'h10408000;
      32633: inst = 32'hc40482f;
      32634: inst = 32'h8220000;
      32635: inst = 32'h10408000;
      32636: inst = 32'hc404839;
      32637: inst = 32'h8220000;
      32638: inst = 32'h10408000;
      32639: inst = 32'hc40485c;
      32640: inst = 32'h8220000;
      32641: inst = 32'h10408000;
      32642: inst = 32'hc404867;
      32643: inst = 32'h8220000;
      32644: inst = 32'h10408000;
      32645: inst = 32'hc404872;
      32646: inst = 32'h8220000;
      32647: inst = 32'h10408000;
      32648: inst = 32'hc40488f;
      32649: inst = 32'h8220000;
      32650: inst = 32'h10408000;
      32651: inst = 32'hc404893;
      32652: inst = 32'h8220000;
      32653: inst = 32'h10408000;
      32654: inst = 32'hc404899;
      32655: inst = 32'h8220000;
      32656: inst = 32'h10408000;
      32657: inst = 32'hc4048ac;
      32658: inst = 32'h8220000;
      32659: inst = 32'h10408000;
      32660: inst = 32'hc4048b2;
      32661: inst = 32'h8220000;
      32662: inst = 32'h10408000;
      32663: inst = 32'hc4048bb;
      32664: inst = 32'h8220000;
      32665: inst = 32'h10408000;
      32666: inst = 32'hc4048bc;
      32667: inst = 32'h8220000;
      32668: inst = 32'h10408000;
      32669: inst = 32'hc4048c7;
      32670: inst = 32'h8220000;
      32671: inst = 32'h10408000;
      32672: inst = 32'hc4048cf;
      32673: inst = 32'h8220000;
      32674: inst = 32'h10408000;
      32675: inst = 32'hc4048d2;
      32676: inst = 32'h8220000;
      32677: inst = 32'h10408000;
      32678: inst = 32'hc4048ef;
      32679: inst = 32'h8220000;
      32680: inst = 32'h10408000;
      32681: inst = 32'hc4048f3;
      32682: inst = 32'h8220000;
      32683: inst = 32'h10408000;
      32684: inst = 32'hc4048f9;
      32685: inst = 32'h8220000;
      32686: inst = 32'h10408000;
      32687: inst = 32'hc40490c;
      32688: inst = 32'h8220000;
      32689: inst = 32'h10408000;
      32690: inst = 32'hc404912;
      32691: inst = 32'h8220000;
      32692: inst = 32'h10408000;
      32693: inst = 32'hc40491b;
      32694: inst = 32'h8220000;
      32695: inst = 32'h10408000;
      32696: inst = 32'hc40491c;
      32697: inst = 32'h8220000;
      32698: inst = 32'h10408000;
      32699: inst = 32'hc404927;
      32700: inst = 32'h8220000;
      32701: inst = 32'h10408000;
      32702: inst = 32'hc40492f;
      32703: inst = 32'h8220000;
      32704: inst = 32'h10408000;
      32705: inst = 32'hc404932;
      32706: inst = 32'h8220000;
      32707: inst = 32'h10408000;
      32708: inst = 32'hc40494f;
      32709: inst = 32'h8220000;
      32710: inst = 32'h10408000;
      32711: inst = 32'hc404959;
      32712: inst = 32'h8220000;
      32713: inst = 32'h10408000;
      32714: inst = 32'hc404972;
      32715: inst = 32'h8220000;
      32716: inst = 32'h10408000;
      32717: inst = 32'hc40497c;
      32718: inst = 32'h8220000;
      32719: inst = 32'h10408000;
      32720: inst = 32'hc404987;
      32721: inst = 32'h8220000;
      32722: inst = 32'h10408000;
      32723: inst = 32'hc404992;
      32724: inst = 32'h8220000;
      32725: inst = 32'h10408000;
      32726: inst = 32'hc4049b9;
      32727: inst = 32'h8220000;
      32728: inst = 32'h10408000;
      32729: inst = 32'hc4049dc;
      32730: inst = 32'h8220000;
      32731: inst = 32'h10408000;
      32732: inst = 32'hc4049e7;
      32733: inst = 32'h8220000;
      32734: inst = 32'h10408000;
      32735: inst = 32'hc4049f2;
      32736: inst = 32'h8220000;
      32737: inst = 32'h10408000;
      32738: inst = 32'hc404e74;
      32739: inst = 32'h8220000;
      32740: inst = 32'h10408000;
      32741: inst = 32'hc404ef4;
      32742: inst = 32'h8220000;
      32743: inst = 32'h10408000;
      32744: inst = 32'hc404ef5;
      32745: inst = 32'h8220000;
      32746: inst = 32'h10408000;
      32747: inst = 32'hc404ef9;
      32748: inst = 32'h8220000;
      32749: inst = 32'h10408000;
      32750: inst = 32'hc404f0e;
      32751: inst = 32'h8220000;
      32752: inst = 32'h10408000;
      32753: inst = 32'hc404f12;
      32754: inst = 32'h8220000;
      32755: inst = 32'h10408000;
      32756: inst = 32'hc404f2c;
      32757: inst = 32'h8220000;
      32758: inst = 32'h10408000;
      32759: inst = 32'hc404f33;
      32760: inst = 32'h8220000;
      32761: inst = 32'h10408000;
      32762: inst = 32'hc404f54;
      32763: inst = 32'h8220000;
      32764: inst = 32'h10408000;
      32765: inst = 32'hc404f59;
      32766: inst = 32'h8220000;
      32767: inst = 32'h10408000;
      32768: inst = 32'hc404f72;
      32769: inst = 32'h8220000;
      32770: inst = 32'h10408000;
      32771: inst = 32'hc404f8c;
      32772: inst = 32'h8220000;
      32773: inst = 32'h10408000;
      32774: inst = 32'hc404fb4;
      32775: inst = 32'h8220000;
      32776: inst = 32'h10408000;
      32777: inst = 32'hc404fb9;
      32778: inst = 32'h8220000;
      32779: inst = 32'h10408000;
      32780: inst = 32'hc404fd2;
      32781: inst = 32'h8220000;
      32782: inst = 32'h10408000;
      32783: inst = 32'hc404fd8;
      32784: inst = 32'h8220000;
      32785: inst = 32'h10408000;
      32786: inst = 32'hc404fe7;
      32787: inst = 32'h8220000;
      32788: inst = 32'h10408000;
      32789: inst = 32'hc405014;
      32790: inst = 32'h8220000;
      32791: inst = 32'hc20630c;
      32792: inst = 32'h10408000;
      32793: inst = 32'hc4046b0;
      32794: inst = 32'h8220000;
      32795: inst = 32'h10408000;
      32796: inst = 32'hc404710;
      32797: inst = 32'h8220000;
      32798: inst = 32'h10408000;
      32799: inst = 32'hc404751;
      32800: inst = 32'h8220000;
      32801: inst = 32'h10408000;
      32802: inst = 32'hc404770;
      32803: inst = 32'h8220000;
      32804: inst = 32'h10408000;
      32805: inst = 32'hc404771;
      32806: inst = 32'h8220000;
      32807: inst = 32'h10408000;
      32808: inst = 32'hc404774;
      32809: inst = 32'h8220000;
      32810: inst = 32'h10408000;
      32811: inst = 32'hc404777;
      32812: inst = 32'h8220000;
      32813: inst = 32'h10408000;
      32814: inst = 32'hc40477b;
      32815: inst = 32'h8220000;
      32816: inst = 32'h10408000;
      32817: inst = 32'hc404783;
      32818: inst = 32'h8220000;
      32819: inst = 32'h10408000;
      32820: inst = 32'hc404786;
      32821: inst = 32'h8220000;
      32822: inst = 32'h10408000;
      32823: inst = 32'hc40478a;
      32824: inst = 32'h8220000;
      32825: inst = 32'h10408000;
      32826: inst = 32'hc404794;
      32827: inst = 32'h8220000;
      32828: inst = 32'h10408000;
      32829: inst = 32'hc404799;
      32830: inst = 32'h8220000;
      32831: inst = 32'h10408000;
      32832: inst = 32'hc40479e;
      32833: inst = 32'h8220000;
      32834: inst = 32'h10408000;
      32835: inst = 32'hc4047a1;
      32836: inst = 32'h8220000;
      32837: inst = 32'h10408000;
      32838: inst = 32'hc4047a4;
      32839: inst = 32'h8220000;
      32840: inst = 32'h10408000;
      32841: inst = 32'hc4047a6;
      32842: inst = 32'h8220000;
      32843: inst = 32'h10408000;
      32844: inst = 32'hc4047a9;
      32845: inst = 32'h8220000;
      32846: inst = 32'h10408000;
      32847: inst = 32'hc4047ad;
      32848: inst = 32'h8220000;
      32849: inst = 32'h10408000;
      32850: inst = 32'hc4047b1;
      32851: inst = 32'h8220000;
      32852: inst = 32'h10408000;
      32853: inst = 32'hc4047f6;
      32854: inst = 32'h8220000;
      32855: inst = 32'h10408000;
      32856: inst = 32'hc404811;
      32857: inst = 32'h8220000;
      32858: inst = 32'h10408000;
      32859: inst = 32'hc404853;
      32860: inst = 32'h8220000;
      32861: inst = 32'h10408000;
      32862: inst = 32'hc404866;
      32863: inst = 32'h8220000;
      32864: inst = 32'h10408000;
      32865: inst = 32'hc404871;
      32866: inst = 32'h8220000;
      32867: inst = 32'h10408000;
      32868: inst = 32'hc404890;
      32869: inst = 32'h8220000;
      32870: inst = 32'h10408000;
      32871: inst = 32'hc404892;
      32872: inst = 32'h8220000;
      32873: inst = 32'h10408000;
      32874: inst = 32'hc40489a;
      32875: inst = 32'h8220000;
      32876: inst = 32'h10408000;
      32877: inst = 32'hc4048ab;
      32878: inst = 32'h8220000;
      32879: inst = 32'h10408000;
      32880: inst = 32'hc4048b1;
      32881: inst = 32'h8220000;
      32882: inst = 32'h10408000;
      32883: inst = 32'hc4048ba;
      32884: inst = 32'h8220000;
      32885: inst = 32'h10408000;
      32886: inst = 32'hc4048bd;
      32887: inst = 32'h8220000;
      32888: inst = 32'h10408000;
      32889: inst = 32'hc4048c6;
      32890: inst = 32'h8220000;
      32891: inst = 32'h10408000;
      32892: inst = 32'hc4048ce;
      32893: inst = 32'h8220000;
      32894: inst = 32'h10408000;
      32895: inst = 32'hc4048d1;
      32896: inst = 32'h8220000;
      32897: inst = 32'h10408000;
      32898: inst = 32'hc4048f0;
      32899: inst = 32'h8220000;
      32900: inst = 32'h10408000;
      32901: inst = 32'hc4048f2;
      32902: inst = 32'h8220000;
      32903: inst = 32'h10408000;
      32904: inst = 32'hc4048fa;
      32905: inst = 32'h8220000;
      32906: inst = 32'h10408000;
      32907: inst = 32'hc40490b;
      32908: inst = 32'h8220000;
      32909: inst = 32'h10408000;
      32910: inst = 32'hc404911;
      32911: inst = 32'h8220000;
      32912: inst = 32'h10408000;
      32913: inst = 32'hc40491a;
      32914: inst = 32'h8220000;
      32915: inst = 32'h10408000;
      32916: inst = 32'hc40491d;
      32917: inst = 32'h8220000;
      32918: inst = 32'h10408000;
      32919: inst = 32'hc404926;
      32920: inst = 32'h8220000;
      32921: inst = 32'h10408000;
      32922: inst = 32'hc40492e;
      32923: inst = 32'h8220000;
      32924: inst = 32'h10408000;
      32925: inst = 32'hc404931;
      32926: inst = 32'h8220000;
      32927: inst = 32'h10408000;
      32928: inst = 32'hc404950;
      32929: inst = 32'h8220000;
      32930: inst = 32'h10408000;
      32931: inst = 32'hc40495a;
      32932: inst = 32'h8220000;
      32933: inst = 32'h10408000;
      32934: inst = 32'hc40497d;
      32935: inst = 32'h8220000;
      32936: inst = 32'h10408000;
      32937: inst = 32'hc404986;
      32938: inst = 32'h8220000;
      32939: inst = 32'h10408000;
      32940: inst = 32'hc404991;
      32941: inst = 32'h8220000;
      32942: inst = 32'h10408000;
      32943: inst = 32'hc404a11;
      32944: inst = 32'h8220000;
      32945: inst = 32'h10408000;
      32946: inst = 32'hc404a19;
      32947: inst = 32'h8220000;
      32948: inst = 32'h10408000;
      32949: inst = 32'hc404a1c;
      32950: inst = 32'h8220000;
      32951: inst = 32'h10408000;
      32952: inst = 32'hc404a1d;
      32953: inst = 32'h8220000;
      32954: inst = 32'h10408000;
      32955: inst = 32'hc404a2a;
      32956: inst = 32'h8220000;
      32957: inst = 32'h10408000;
      32958: inst = 32'hc404a34;
      32959: inst = 32'h8220000;
      32960: inst = 32'h10408000;
      32961: inst = 32'hc404a39;
      32962: inst = 32'h8220000;
      32963: inst = 32'h10408000;
      32964: inst = 32'hc404a3c;
      32965: inst = 32'h8220000;
      32966: inst = 32'h10408000;
      32967: inst = 32'hc404a3f;
      32968: inst = 32'h8220000;
      32969: inst = 32'h10408000;
      32970: inst = 32'hc404a40;
      32971: inst = 32'h8220000;
      32972: inst = 32'h10408000;
      32973: inst = 32'hc404a46;
      32974: inst = 32'h8220000;
      32975: inst = 32'h10408000;
      32976: inst = 32'hc404a47;
      32977: inst = 32'h8220000;
      32978: inst = 32'h10408000;
      32979: inst = 32'hc404a48;
      32980: inst = 32'h8220000;
      32981: inst = 32'h10408000;
      32982: inst = 32'hc404a4d;
      32983: inst = 32'h8220000;
      32984: inst = 32'h10408000;
      32985: inst = 32'hc404a51;
      32986: inst = 32'h8220000;
      32987: inst = 32'h10408000;
      32988: inst = 32'hc404a52;
      32989: inst = 32'h8220000;
      32990: inst = 32'h10408000;
      32991: inst = 32'hc404a53;
      32992: inst = 32'h8220000;
      32993: inst = 32'h10408000;
      32994: inst = 32'hc404d80;
      32995: inst = 32'h8220000;
      32996: inst = 32'h10408000;
      32997: inst = 32'hc404d8a;
      32998: inst = 32'h8220000;
      32999: inst = 32'h10408000;
      33000: inst = 32'hc404d9e;
      33001: inst = 32'h8220000;
      33002: inst = 32'h10408000;
      33003: inst = 32'hc404da3;
      33004: inst = 32'h8220000;
      33005: inst = 32'h10408000;
      33006: inst = 32'hc404dcd;
      33007: inst = 32'h8220000;
      33008: inst = 32'h10408000;
      33009: inst = 32'hc404dd2;
      33010: inst = 32'h8220000;
      33011: inst = 32'h10408000;
      33012: inst = 32'hc404dd3;
      33013: inst = 32'h8220000;
      33014: inst = 32'h10408000;
      33015: inst = 32'hc404dd7;
      33016: inst = 32'h8220000;
      33017: inst = 32'h10408000;
      33018: inst = 32'hc404dde;
      33019: inst = 32'h8220000;
      33020: inst = 32'h10408000;
      33021: inst = 32'hc404de2;
      33022: inst = 32'h8220000;
      33023: inst = 32'h10408000;
      33024: inst = 32'hc404dec;
      33025: inst = 32'h8220000;
      33026: inst = 32'h10408000;
      33027: inst = 32'hc404df0;
      33028: inst = 32'h8220000;
      33029: inst = 32'h10408000;
      33030: inst = 32'hc404dfa;
      33031: inst = 32'h8220000;
      33032: inst = 32'h10408000;
      33033: inst = 32'hc404e00;
      33034: inst = 32'h8220000;
      33035: inst = 32'h10408000;
      33036: inst = 32'hc404e05;
      33037: inst = 32'h8220000;
      33038: inst = 32'h10408000;
      33039: inst = 32'hc404e09;
      33040: inst = 32'h8220000;
      33041: inst = 32'h10408000;
      33042: inst = 32'hc404e0e;
      33043: inst = 32'h8220000;
      33044: inst = 32'h10408000;
      33045: inst = 32'hc404e14;
      33046: inst = 32'h8220000;
      33047: inst = 32'h10408000;
      33048: inst = 32'hc404e15;
      33049: inst = 32'h8220000;
      33050: inst = 32'h10408000;
      33051: inst = 32'hc404e93;
      33052: inst = 32'h8220000;
      33053: inst = 32'h10408000;
      33054: inst = 32'hc404e9d;
      33055: inst = 32'h8220000;
      33056: inst = 32'h10408000;
      33057: inst = 32'hc404eb9;
      33058: inst = 32'h8220000;
      33059: inst = 32'h10408000;
      33060: inst = 32'hc404ec8;
      33061: inst = 32'h8220000;
      33062: inst = 32'h10408000;
      33063: inst = 32'hc404ef3;
      33064: inst = 32'h8220000;
      33065: inst = 32'h10408000;
      33066: inst = 32'hc404efd;
      33067: inst = 32'h8220000;
      33068: inst = 32'h10408000;
      33069: inst = 32'hc404f13;
      33070: inst = 32'h8220000;
      33071: inst = 32'h10408000;
      33072: inst = 32'hc404f2d;
      33073: inst = 32'h8220000;
      33074: inst = 32'h10408000;
      33075: inst = 32'hc404f53;
      33076: inst = 32'h8220000;
      33077: inst = 32'h10408000;
      33078: inst = 32'hc404f5d;
      33079: inst = 32'h8220000;
      33080: inst = 32'h10408000;
      33081: inst = 32'hc404f73;
      33082: inst = 32'h8220000;
      33083: inst = 32'h10408000;
      33084: inst = 32'hc404f8d;
      33085: inst = 32'h8220000;
      33086: inst = 32'h10408000;
      33087: inst = 32'hc404fb3;
      33088: inst = 32'h8220000;
      33089: inst = 32'h10408000;
      33090: inst = 32'hc404fd7;
      33091: inst = 32'h8220000;
      33092: inst = 32'h10408000;
      33093: inst = 32'hc404fdd;
      33094: inst = 32'h8220000;
      33095: inst = 32'h10408000;
      33096: inst = 32'hc405020;
      33097: inst = 32'h8220000;
      33098: inst = 32'h10408000;
      33099: inst = 32'hc40502a;
      33100: inst = 32'h8220000;
      33101: inst = 32'h10408000;
      33102: inst = 32'hc40503e;
      33103: inst = 32'h8220000;
      33104: inst = 32'h10408000;
      33105: inst = 32'hc405043;
      33106: inst = 32'h8220000;
      33107: inst = 32'h10408000;
      33108: inst = 32'hc40506d;
      33109: inst = 32'h8220000;
      33110: inst = 32'h10408000;
      33111: inst = 32'hc405070;
      33112: inst = 32'h8220000;
      33113: inst = 32'h10408000;
      33114: inst = 32'hc405071;
      33115: inst = 32'h8220000;
      33116: inst = 32'h10408000;
      33117: inst = 32'hc405074;
      33118: inst = 32'h8220000;
      33119: inst = 32'h10408000;
      33120: inst = 32'hc405077;
      33121: inst = 32'h8220000;
      33122: inst = 32'h10408000;
      33123: inst = 32'hc40507c;
      33124: inst = 32'h8220000;
      33125: inst = 32'h10408000;
      33126: inst = 32'hc405082;
      33127: inst = 32'h8220000;
      33128: inst = 32'h10408000;
      33129: inst = 32'hc40508c;
      33130: inst = 32'h8220000;
      33131: inst = 32'h10408000;
      33132: inst = 32'hc405090;
      33133: inst = 32'h8220000;
      33134: inst = 32'h10408000;
      33135: inst = 32'hc405099;
      33136: inst = 32'h8220000;
      33137: inst = 32'h10408000;
      33138: inst = 32'hc40509c;
      33139: inst = 32'h8220000;
      33140: inst = 32'h10408000;
      33141: inst = 32'hc4050a0;
      33142: inst = 32'h8220000;
      33143: inst = 32'h10408000;
      33144: inst = 32'hc4050a5;
      33145: inst = 32'h8220000;
      33146: inst = 32'h10408000;
      33147: inst = 32'hc4050a8;
      33148: inst = 32'h8220000;
      33149: inst = 32'h10408000;
      33150: inst = 32'hc4050ab;
      33151: inst = 32'h8220000;
      33152: inst = 32'h10408000;
      33153: inst = 32'hc4050ae;
      33154: inst = 32'h8220000;
      33155: inst = 32'h10408000;
      33156: inst = 32'hc4050b1;
      33157: inst = 32'h8220000;
      33158: inst = 32'h10408000;
      33159: inst = 32'hc4050b2;
      33160: inst = 32'h8220000;
      33161: inst = 32'h10408000;
      33162: inst = 32'hc4050b5;
      33163: inst = 32'h8220000;
      33164: inst = 32'hc20defb;
      33165: inst = 32'h10408000;
      33166: inst = 32'hc404775;
      33167: inst = 32'h8220000;
      33168: inst = 32'h10408000;
      33169: inst = 32'hc404784;
      33170: inst = 32'h8220000;
      33171: inst = 32'h10408000;
      33172: inst = 32'hc4047a2;
      33173: inst = 32'h8220000;
      33174: inst = 32'h10408000;
      33175: inst = 32'hc4047d2;
      33176: inst = 32'h8220000;
      33177: inst = 32'h10408000;
      33178: inst = 32'hc4047d5;
      33179: inst = 32'h8220000;
      33180: inst = 32'h10408000;
      33181: inst = 32'hc4047e4;
      33182: inst = 32'h8220000;
      33183: inst = 32'h10408000;
      33184: inst = 32'hc4047eb;
      33185: inst = 32'h8220000;
      33186: inst = 32'h10408000;
      33187: inst = 32'hc4047fa;
      33188: inst = 32'h8220000;
      33189: inst = 32'h10408000;
      33190: inst = 32'hc404802;
      33191: inst = 32'h8220000;
      33192: inst = 32'h10408000;
      33193: inst = 32'hc40480e;
      33194: inst = 32'h8220000;
      33195: inst = 32'h10408000;
      33196: inst = 32'hc404833;
      33197: inst = 32'h8220000;
      33198: inst = 32'h10408000;
      33199: inst = 32'hc40496c;
      33200: inst = 32'h8220000;
      33201: inst = 32'h10408000;
      33202: inst = 32'hc40497b;
      33203: inst = 32'h8220000;
      33204: inst = 32'h10408000;
      33205: inst = 32'hc40498f;
      33206: inst = 32'h8220000;
      33207: inst = 32'h10408000;
      33208: inst = 32'hc4049af;
      33209: inst = 32'h8220000;
      33210: inst = 32'h10408000;
      33211: inst = 32'hc4049b6;
      33212: inst = 32'h8220000;
      33213: inst = 32'h10408000;
      33214: inst = 32'hc4049bd;
      33215: inst = 32'h8220000;
      33216: inst = 32'h10408000;
      33217: inst = 32'hc4049c5;
      33218: inst = 32'h8220000;
      33219: inst = 32'h10408000;
      33220: inst = 32'hc4049d3;
      33221: inst = 32'h8220000;
      33222: inst = 32'h10408000;
      33223: inst = 32'hc4049e0;
      33224: inst = 32'h8220000;
      33225: inst = 32'h10408000;
      33226: inst = 32'hc4049e3;
      33227: inst = 32'h8220000;
      33228: inst = 32'h10408000;
      33229: inst = 32'hc404d10;
      33230: inst = 32'h8220000;
      33231: inst = 32'h10408000;
      33232: inst = 32'hc404d51;
      33233: inst = 32'h8220000;
      33234: inst = 32'h10408000;
      33235: inst = 32'hc404e31;
      33236: inst = 32'h8220000;
      33237: inst = 32'h10408000;
      33238: inst = 32'hc404e3a;
      33239: inst = 32'h8220000;
      33240: inst = 32'h10408000;
      33241: inst = 32'hc404e41;
      33242: inst = 32'h8220000;
      33243: inst = 32'h10408000;
      33244: inst = 32'hc404e4b;
      33245: inst = 32'h8220000;
      33246: inst = 32'h10408000;
      33247: inst = 32'hc404e5f;
      33248: inst = 32'h8220000;
      33249: inst = 32'h10408000;
      33250: inst = 32'hc404e64;
      33251: inst = 32'h8220000;
      33252: inst = 32'h10408000;
      33253: inst = 32'hc404e94;
      33254: inst = 32'h8220000;
      33255: inst = 32'h10408000;
      33256: inst = 32'hc404e95;
      33257: inst = 32'h8220000;
      33258: inst = 32'h10408000;
      33259: inst = 32'hc404e99;
      33260: inst = 32'h8220000;
      33261: inst = 32'h10408000;
      33262: inst = 32'hc404eae;
      33263: inst = 32'h8220000;
      33264: inst = 32'h10408000;
      33265: inst = 32'hc404eb2;
      33266: inst = 32'h8220000;
      33267: inst = 32'h10408000;
      33268: inst = 32'hc404f4e;
      33269: inst = 32'h8220000;
      33270: inst = 32'h10408000;
      33271: inst = 32'hc404fb5;
      33272: inst = 32'h8220000;
      33273: inst = 32'h10408000;
      33274: inst = 32'hc404fce;
      33275: inst = 32'h8220000;
      33276: inst = 32'h10408000;
      33277: inst = 32'hc405010;
      33278: inst = 32'h8220000;
      33279: inst = 32'h10408000;
      33280: inst = 32'hc40504d;
      33281: inst = 32'h8220000;
      33282: inst = 32'h10408000;
      33283: inst = 32'hc405051;
      33284: inst = 32'h8220000;
      33285: inst = 32'hc208410;
      33286: inst = 32'h10408000;
      33287: inst = 32'hc404779;
      33288: inst = 32'h8220000;
      33289: inst = 32'h10408000;
      33290: inst = 32'hc40479c;
      33291: inst = 32'h8220000;
      33292: inst = 32'h10408000;
      33293: inst = 32'hc4047e8;
      33294: inst = 32'h8220000;
      33295: inst = 32'h10408000;
      33296: inst = 32'hc4047f2;
      33297: inst = 32'h8220000;
      33298: inst = 32'h10408000;
      33299: inst = 32'hc4047f7;
      33300: inst = 32'h8220000;
      33301: inst = 32'h10408000;
      33302: inst = 32'hc40480b;
      33303: inst = 32'h8220000;
      33304: inst = 32'h10408000;
      33305: inst = 32'hc404830;
      33306: inst = 32'h8220000;
      33307: inst = 32'h10408000;
      33308: inst = 32'hc40484b;
      33309: inst = 32'h8220000;
      33310: inst = 32'h10408000;
      33311: inst = 32'hc40485a;
      33312: inst = 32'h8220000;
      33313: inst = 32'h10408000;
      33314: inst = 32'hc40486e;
      33315: inst = 32'h8220000;
      33316: inst = 32'h10408000;
      33317: inst = 32'hc40496b;
      33318: inst = 32'h8220000;
      33319: inst = 32'h10408000;
      33320: inst = 32'hc40497a;
      33321: inst = 32'h8220000;
      33322: inst = 32'h10408000;
      33323: inst = 32'hc40498e;
      33324: inst = 32'h8220000;
      33325: inst = 32'h10408000;
      33326: inst = 32'hc4049c8;
      33327: inst = 32'h8220000;
      33328: inst = 32'h10408000;
      33329: inst = 32'hc4049d2;
      33330: inst = 32'h8220000;
      33331: inst = 32'h10408000;
      33332: inst = 32'hc4049d7;
      33333: inst = 32'h8220000;
      33334: inst = 32'h10408000;
      33335: inst = 32'hc4049eb;
      33336: inst = 32'h8220000;
      33337: inst = 32'h10408000;
      33338: inst = 32'hc404e52;
      33339: inst = 32'h8220000;
      33340: inst = 32'h10408000;
      33341: inst = 32'hc404eee;
      33342: inst = 32'h8220000;
      33343: inst = 32'h10408000;
      33344: inst = 32'hc404ff5;
      33345: inst = 32'h8220000;
      33346: inst = 32'h10408000;
      33347: inst = 32'hc405019;
      33348: inst = 32'h8220000;
      33349: inst = 32'h10408000;
      33350: inst = 32'hc40501f;
      33351: inst = 32'h8220000;
      33352: inst = 32'h10408000;
      33353: inst = 32'hc405032;
      33354: inst = 32'h8220000;
      33355: inst = 32'h10408000;
      33356: inst = 32'hc405050;
      33357: inst = 32'h8220000;
      33358: inst = 32'hc204a69;
      33359: inst = 32'h10408000;
      33360: inst = 32'hc40477c;
      33361: inst = 32'h8220000;
      33362: inst = 32'h10408000;
      33363: inst = 32'hc404789;
      33364: inst = 32'h8220000;
      33365: inst = 32'h10408000;
      33366: inst = 32'hc404798;
      33367: inst = 32'h8220000;
      33368: inst = 32'h10408000;
      33369: inst = 32'hc40479f;
      33370: inst = 32'h8220000;
      33371: inst = 32'h10408000;
      33372: inst = 32'hc4047aa;
      33373: inst = 32'h8220000;
      33374: inst = 32'h10408000;
      33375: inst = 32'hc4047ac;
      33376: inst = 32'h8220000;
      33377: inst = 32'h10408000;
      33378: inst = 32'hc4047d8;
      33379: inst = 32'h8220000;
      33380: inst = 32'h10408000;
      33381: inst = 32'hc4047ec;
      33382: inst = 32'h8220000;
      33383: inst = 32'h10408000;
      33384: inst = 32'hc4047fb;
      33385: inst = 32'h8220000;
      33386: inst = 32'h10408000;
      33387: inst = 32'hc404805;
      33388: inst = 32'h8220000;
      33389: inst = 32'h10408000;
      33390: inst = 32'hc40480f;
      33391: inst = 32'h8220000;
      33392: inst = 32'h10408000;
      33393: inst = 32'hc404973;
      33394: inst = 32'h8220000;
      33395: inst = 32'h10408000;
      33396: inst = 32'hc4049b3;
      33397: inst = 32'h8220000;
      33398: inst = 32'h10408000;
      33399: inst = 32'hc4049cc;
      33400: inst = 32'h8220000;
      33401: inst = 32'h10408000;
      33402: inst = 32'hc4049d6;
      33403: inst = 32'h8220000;
      33404: inst = 32'h10408000;
      33405: inst = 32'hc4049e9;
      33406: inst = 32'h8220000;
      33407: inst = 32'h10408000;
      33408: inst = 32'hc4049ef;
      33409: inst = 32'h8220000;
      33410: inst = 32'h10408000;
      33411: inst = 32'hc4049f4;
      33412: inst = 32'h8220000;
      33413: inst = 32'h10408000;
      33414: inst = 32'hc404a16;
      33415: inst = 32'h8220000;
      33416: inst = 32'h10408000;
      33417: inst = 32'hc404a17;
      33418: inst = 32'h8220000;
      33419: inst = 32'h10408000;
      33420: inst = 32'hc404a1a;
      33421: inst = 32'h8220000;
      33422: inst = 32'h10408000;
      33423: inst = 32'hc404a25;
      33424: inst = 32'h8220000;
      33425: inst = 32'h10408000;
      33426: inst = 32'hc404a26;
      33427: inst = 32'h8220000;
      33428: inst = 32'h10408000;
      33429: inst = 32'hc404a29;
      33430: inst = 32'h8220000;
      33431: inst = 32'h10408000;
      33432: inst = 32'hc404a33;
      33433: inst = 32'h8220000;
      33434: inst = 32'h10408000;
      33435: inst = 32'hc404a38;
      33436: inst = 32'h8220000;
      33437: inst = 32'h10408000;
      33438: inst = 32'hc404a3d;
      33439: inst = 32'h8220000;
      33440: inst = 32'h10408000;
      33441: inst = 32'hc404a43;
      33442: inst = 32'h8220000;
      33443: inst = 32'h10408000;
      33444: inst = 32'hc404a44;
      33445: inst = 32'h8220000;
      33446: inst = 32'h10408000;
      33447: inst = 32'hc404a4c;
      33448: inst = 32'h8220000;
      33449: inst = 32'h10408000;
      33450: inst = 32'hc404caf;
      33451: inst = 32'h8220000;
      33452: inst = 32'h10408000;
      33453: inst = 32'hc404cf0;
      33454: inst = 32'h8220000;
      33455: inst = 32'h10408000;
      33456: inst = 32'hc404d0f;
      33457: inst = 32'h8220000;
      33458: inst = 32'h10408000;
      33459: inst = 32'hc404d50;
      33460: inst = 32'h8220000;
      33461: inst = 32'h10408000;
      33462: inst = 32'hc404dce;
      33463: inst = 32'h8220000;
      33464: inst = 32'h10408000;
      33465: inst = 32'hc404dd8;
      33466: inst = 32'h8220000;
      33467: inst = 32'h10408000;
      33468: inst = 32'hc404ddb;
      33469: inst = 32'h8220000;
      33470: inst = 32'h10408000;
      33471: inst = 32'hc404ddd;
      33472: inst = 32'h8220000;
      33473: inst = 32'h10408000;
      33474: inst = 32'hc404ddf;
      33475: inst = 32'h8220000;
      33476: inst = 32'h10408000;
      33477: inst = 32'hc404de9;
      33478: inst = 32'h8220000;
      33479: inst = 32'h10408000;
      33480: inst = 32'hc404df1;
      33481: inst = 32'h8220000;
      33482: inst = 32'h10408000;
      33483: inst = 32'hc404df9;
      33484: inst = 32'h8220000;
      33485: inst = 32'h10408000;
      33486: inst = 32'hc404dfb;
      33487: inst = 32'h8220000;
      33488: inst = 32'h10408000;
      33489: inst = 32'hc404dfd;
      33490: inst = 32'h8220000;
      33491: inst = 32'h10408000;
      33492: inst = 32'hc404e02;
      33493: inst = 32'h8220000;
      33494: inst = 32'h10408000;
      33495: inst = 32'hc404e08;
      33496: inst = 32'h8220000;
      33497: inst = 32'h10408000;
      33498: inst = 32'hc404e0a;
      33499: inst = 32'h8220000;
      33500: inst = 32'h10408000;
      33501: inst = 32'hc404e0f;
      33502: inst = 32'h8220000;
      33503: inst = 32'h10408000;
      33504: inst = 32'hc404e2b;
      33505: inst = 32'h8220000;
      33506: inst = 32'h10408000;
      33507: inst = 32'hc404e35;
      33508: inst = 32'h8220000;
      33509: inst = 32'h10408000;
      33510: inst = 32'hc404e43;
      33511: inst = 32'h8220000;
      33512: inst = 32'h10408000;
      33513: inst = 32'hc404e4d;
      33514: inst = 32'h8220000;
      33515: inst = 32'h10408000;
      33516: inst = 32'hc404e4e;
      33517: inst = 32'h8220000;
      33518: inst = 32'h10408000;
      33519: inst = 32'hc404e61;
      33520: inst = 32'h8220000;
      33521: inst = 32'h10408000;
      33522: inst = 32'hc404e66;
      33523: inst = 32'h8220000;
      33524: inst = 32'h10408000;
      33525: inst = 32'hc404e6c;
      33526: inst = 32'h8220000;
      33527: inst = 32'h10408000;
      33528: inst = 32'hc404e73;
      33529: inst = 32'h8220000;
      33530: inst = 32'h10408000;
      33531: inst = 32'hc404eeb;
      33532: inst = 32'h8220000;
      33533: inst = 32'h10408000;
      33534: inst = 32'hc404f0d;
      33535: inst = 32'h8220000;
      33536: inst = 32'h10408000;
      33537: inst = 32'hc404f18;
      33538: inst = 32'h8220000;
      33539: inst = 32'h10408000;
      33540: inst = 32'hc404f27;
      33541: inst = 32'h8220000;
      33542: inst = 32'h10408000;
      33543: inst = 32'hc404f34;
      33544: inst = 32'h8220000;
      33545: inst = 32'h10408000;
      33546: inst = 32'hc404f6d;
      33547: inst = 32'h8220000;
      33548: inst = 32'h10408000;
      33549: inst = 32'hc405015;
      33550: inst = 32'h8220000;
      33551: inst = 32'h10408000;
      33552: inst = 32'hc40502e;
      33553: inst = 32'h8220000;
      33554: inst = 32'h10408000;
      33555: inst = 32'hc405056;
      33556: inst = 32'h8220000;
      33557: inst = 32'h10408000;
      33558: inst = 32'hc40506e;
      33559: inst = 32'h8220000;
      33560: inst = 32'h10408000;
      33561: inst = 32'hc405073;
      33562: inst = 32'h8220000;
      33563: inst = 32'h10408000;
      33564: inst = 32'hc40507b;
      33565: inst = 32'h8220000;
      33566: inst = 32'h10408000;
      33567: inst = 32'hc40509a;
      33568: inst = 32'h8220000;
      33569: inst = 32'h10408000;
      33570: inst = 32'hc4050a9;
      33571: inst = 32'h8220000;
      33572: inst = 32'h10408000;
      33573: inst = 32'hc4050af;
      33574: inst = 32'h8220000;
      33575: inst = 32'h10408000;
      33576: inst = 32'hc4050b4;
      33577: inst = 32'h8220000;
      33578: inst = 32'hc209492;
      33579: inst = 32'h10408000;
      33580: inst = 32'hc4047a7;
      33581: inst = 32'h8220000;
      33582: inst = 32'h10408000;
      33583: inst = 32'hc404832;
      33584: inst = 32'h8220000;
      33585: inst = 32'h10408000;
      33586: inst = 32'hc404868;
      33587: inst = 32'h8220000;
      33588: inst = 32'h10408000;
      33589: inst = 32'hc4048a7;
      33590: inst = 32'h8220000;
      33591: inst = 32'h10408000;
      33592: inst = 32'hc4048b6;
      33593: inst = 32'h8220000;
      33594: inst = 32'h10408000;
      33595: inst = 32'hc4048ca;
      33596: inst = 32'h8220000;
      33597: inst = 32'h10408000;
      33598: inst = 32'hc404907;
      33599: inst = 32'h8220000;
      33600: inst = 32'h10408000;
      33601: inst = 32'hc404916;
      33602: inst = 32'h8220000;
      33603: inst = 32'h10408000;
      33604: inst = 32'hc40492a;
      33605: inst = 32'h8220000;
      33606: inst = 32'h10408000;
      33607: inst = 32'hc404952;
      33608: inst = 32'h8220000;
      33609: inst = 32'h10408000;
      33610: inst = 32'hc4049db;
      33611: inst = 32'h8220000;
      33612: inst = 32'h10408000;
      33613: inst = 32'hc404e3f;
      33614: inst = 32'h8220000;
      33615: inst = 32'h10408000;
      33616: inst = 32'hc404e49;
      33617: inst = 32'h8220000;
      33618: inst = 32'h10408000;
      33619: inst = 32'hc404e5d;
      33620: inst = 32'h8220000;
      33621: inst = 32'h10408000;
      33622: inst = 32'hc404e62;
      33623: inst = 32'h8220000;
      33624: inst = 32'h10408000;
      33625: inst = 32'hc404ecf;
      33626: inst = 32'h8220000;
      33627: inst = 32'h10408000;
      33628: inst = 32'hc404f79;
      33629: inst = 32'h8220000;
      33630: inst = 32'h10408000;
      33631: inst = 32'hc404f88;
      33632: inst = 32'h8220000;
      33633: inst = 32'h10408000;
      33634: inst = 32'hc404fed;
      33635: inst = 32'h8220000;
      33636: inst = 32'hc20d69a;
      33637: inst = 32'h10408000;
      33638: inst = 32'hc4047d0;
      33639: inst = 32'h8220000;
      33640: inst = 32'h10408000;
      33641: inst = 32'hc4047da;
      33642: inst = 32'h8220000;
      33643: inst = 32'h10408000;
      33644: inst = 32'hc4047f5;
      33645: inst = 32'h8220000;
      33646: inst = 32'h10408000;
      33647: inst = 32'hc4047fd;
      33648: inst = 32'h8220000;
      33649: inst = 32'h10408000;
      33650: inst = 32'hc4048a8;
      33651: inst = 32'h8220000;
      33652: inst = 32'h10408000;
      33653: inst = 32'hc4048b7;
      33654: inst = 32'h8220000;
      33655: inst = 32'h10408000;
      33656: inst = 32'hc4048cb;
      33657: inst = 32'h8220000;
      33658: inst = 32'h10408000;
      33659: inst = 32'hc404953;
      33660: inst = 32'h8220000;
      33661: inst = 32'h10408000;
      33662: inst = 32'hc4049b2;
      33663: inst = 32'h8220000;
      33664: inst = 32'h10408000;
      33665: inst = 32'hc4049cb;
      33666: inst = 32'h8220000;
      33667: inst = 32'h10408000;
      33668: inst = 32'hc4049da;
      33669: inst = 32'h8220000;
      33670: inst = 32'h10408000;
      33671: inst = 32'hc4049ee;
      33672: inst = 32'h8220000;
      33673: inst = 32'h10408000;
      33674: inst = 32'hc404e33;
      33675: inst = 32'h8220000;
      33676: inst = 32'h10408000;
      33677: inst = 32'hc404e36;
      33678: inst = 32'h8220000;
      33679: inst = 32'h10408000;
      33680: inst = 32'hc404e38;
      33681: inst = 32'h8220000;
      33682: inst = 32'h10408000;
      33683: inst = 32'hc404e4f;
      33684: inst = 32'h8220000;
      33685: inst = 32'h10408000;
      33686: inst = 32'hc404e51;
      33687: inst = 32'h8220000;
      33688: inst = 32'h10408000;
      33689: inst = 32'hc404e5b;
      33690: inst = 32'h8220000;
      33691: inst = 32'h10408000;
      33692: inst = 32'hc404e6a;
      33693: inst = 32'h8220000;
      33694: inst = 32'h10408000;
      33695: inst = 32'hc404e6d;
      33696: inst = 32'h8220000;
      33697: inst = 32'h10408000;
      33698: inst = 32'hc404eed;
      33699: inst = 32'h8220000;
      33700: inst = 32'h10408000;
      33701: inst = 32'hc404efa;
      33702: inst = 32'h8220000;
      33703: inst = 32'h10408000;
      33704: inst = 32'hc404f1a;
      33705: inst = 32'h8220000;
      33706: inst = 32'h10408000;
      33707: inst = 32'hc404f1b;
      33708: inst = 32'h8220000;
      33709: inst = 32'h10408000;
      33710: inst = 32'hc404f29;
      33711: inst = 32'h8220000;
      33712: inst = 32'h10408000;
      33713: inst = 32'hc404f2a;
      33714: inst = 32'h8220000;
      33715: inst = 32'h10408000;
      33716: inst = 32'hc404f5a;
      33717: inst = 32'h8220000;
      33718: inst = 32'h10408000;
      33719: inst = 32'hc404fba;
      33720: inst = 32'h8220000;
      33721: inst = 32'h10408000;
      33722: inst = 32'hc404fe6;
      33723: inst = 32'h8220000;
      33724: inst = 32'h10408000;
      33725: inst = 32'hc40500c;
      33726: inst = 32'h8220000;
      33727: inst = 32'h10408000;
      33728: inst = 32'hc405038;
      33729: inst = 32'h8220000;
      33730: inst = 32'h10408000;
      33731: inst = 32'hc40503b;
      33732: inst = 32'h8220000;
      33733: inst = 32'h10408000;
      33734: inst = 32'hc405047;
      33735: inst = 32'h8220000;
      33736: inst = 32'h10408000;
      33737: inst = 32'hc40504a;
      33738: inst = 32'h8220000;
      33739: inst = 32'hc20bdd7;
      33740: inst = 32'h10408000;
      33741: inst = 32'hc4047d1;
      33742: inst = 32'h8220000;
      33743: inst = 32'h10408000;
      33744: inst = 32'hc4047d6;
      33745: inst = 32'h8220000;
      33746: inst = 32'h10408000;
      33747: inst = 32'hc4047e5;
      33748: inst = 32'h8220000;
      33749: inst = 32'h10408000;
      33750: inst = 32'hc404803;
      33751: inst = 32'h8220000;
      33752: inst = 32'h10408000;
      33753: inst = 32'hc404855;
      33754: inst = 32'h8220000;
      33755: inst = 32'h10408000;
      33756: inst = 32'hc4049c9;
      33757: inst = 32'h8220000;
      33758: inst = 32'h10408000;
      33759: inst = 32'hc4049d8;
      33760: inst = 32'h8220000;
      33761: inst = 32'h10408000;
      33762: inst = 32'hc4049ec;
      33763: inst = 32'h8220000;
      33764: inst = 32'h10408000;
      33765: inst = 32'hc404de0;
      33766: inst = 32'h8220000;
      33767: inst = 32'h10408000;
      33768: inst = 32'hc404dea;
      33769: inst = 32'h8220000;
      33770: inst = 32'h10408000;
      33771: inst = 32'hc404dfe;
      33772: inst = 32'h8220000;
      33773: inst = 32'h10408000;
      33774: inst = 32'hc404e03;
      33775: inst = 32'h8220000;
      33776: inst = 32'h10408000;
      33777: inst = 32'hc404e2c;
      33778: inst = 32'h8220000;
      33779: inst = 32'h10408000;
      33780: inst = 32'hc404e2e;
      33781: inst = 32'h8220000;
      33782: inst = 32'h10408000;
      33783: inst = 32'hc404e32;
      33784: inst = 32'h8220000;
      33785: inst = 32'h10408000;
      33786: inst = 32'hc404e40;
      33787: inst = 32'h8220000;
      33788: inst = 32'h10408000;
      33789: inst = 32'hc404e4a;
      33790: inst = 32'h8220000;
      33791: inst = 32'h10408000;
      33792: inst = 32'hc404e5e;
      33793: inst = 32'h8220000;
      33794: inst = 32'h10408000;
      33795: inst = 32'hc404e63;
      33796: inst = 32'h8220000;
      33797: inst = 32'h10408000;
      33798: inst = 32'hc404e6f;
      33799: inst = 32'h8220000;
      33800: inst = 32'h10408000;
      33801: inst = 32'hc404e8f;
      33802: inst = 32'h8220000;
      33803: inst = 32'h10408000;
      33804: inst = 32'hc404ed0;
      33805: inst = 32'h8220000;
      33806: inst = 32'h10408000;
      33807: inst = 32'hc404fab;
      33808: inst = 32'h8220000;
      33809: inst = 32'h10408000;
      33810: inst = 32'hc405039;
      33811: inst = 32'h8220000;
      33812: inst = 32'h10408000;
      33813: inst = 32'hc405048;
      33814: inst = 32'h8220000;
      33815: inst = 32'h10408000;
      33816: inst = 32'hc40504f;
      33817: inst = 32'h8220000;
      33818: inst = 32'hc20ef5d;
      33819: inst = 32'h10408000;
      33820: inst = 32'hc4047dc;
      33821: inst = 32'h8220000;
      33822: inst = 32'h10408000;
      33823: inst = 32'hc4047ff;
      33824: inst = 32'h8220000;
      33825: inst = 32'h10408000;
      33826: inst = 32'hc404848;
      33827: inst = 32'h8220000;
      33828: inst = 32'h10408000;
      33829: inst = 32'hc404852;
      33830: inst = 32'h8220000;
      33831: inst = 32'h10408000;
      33832: inst = 32'hc404857;
      33833: inst = 32'h8220000;
      33834: inst = 32'h10408000;
      33835: inst = 32'hc40486b;
      33836: inst = 32'h8220000;
      33837: inst = 32'h10408000;
      33838: inst = 32'hc404968;
      33839: inst = 32'h8220000;
      33840: inst = 32'h10408000;
      33841: inst = 32'hc404977;
      33842: inst = 32'h8220000;
      33843: inst = 32'h10408000;
      33844: inst = 32'hc40498b;
      33845: inst = 32'h8220000;
      33846: inst = 32'h10408000;
      33847: inst = 32'hc404eec;
      33848: inst = 32'h8220000;
      33849: inst = 32'h10408000;
      33850: inst = 32'hc404f55;
      33851: inst = 32'h8220000;
      33852: inst = 32'h10408000;
      33853: inst = 32'hc404f6e;
      33854: inst = 32'h8220000;
      33855: inst = 32'h10408000;
      33856: inst = 32'hc404f78;
      33857: inst = 32'h8220000;
      33858: inst = 32'h10408000;
      33859: inst = 32'hc404f87;
      33860: inst = 32'h8220000;
      33861: inst = 32'h10408000;
      33862: inst = 32'hc404faf;
      33863: inst = 32'h8220000;
      33864: inst = 32'h10408000;
      33865: inst = 32'hc404ff4;
      33866: inst = 32'h8220000;
      33867: inst = 32'h10408000;
      33868: inst = 32'hc40501b;
      33869: inst = 32'h8220000;
      33870: inst = 32'h10408000;
      33871: inst = 32'hc40501e;
      33872: inst = 32'h8220000;
      33873: inst = 32'h10408000;
      33874: inst = 32'hc405021;
      33875: inst = 32'h8220000;
      33876: inst = 32'h10408000;
      33877: inst = 32'hc40502b;
      33878: inst = 32'h8220000;
      33879: inst = 32'h10408000;
      33880: inst = 32'hc40503c;
      33881: inst = 32'h8220000;
      33882: inst = 32'h10408000;
      33883: inst = 32'hc40503f;
      33884: inst = 32'h8220000;
      33885: inst = 32'h10408000;
      33886: inst = 32'hc405044;
      33887: inst = 32'h8220000;
      33888: inst = 32'h10408000;
      33889: inst = 32'hc40504b;
      33890: inst = 32'h8220000;
      33891: inst = 32'h10408000;
      33892: inst = 32'hc405055;
      33893: inst = 32'h8220000;
      33894: inst = 32'hc20c638;
      33895: inst = 32'h10408000;
      33896: inst = 32'hc4047e9;
      33897: inst = 32'h8220000;
      33898: inst = 32'h10408000;
      33899: inst = 32'hc4047f3;
      33900: inst = 32'h8220000;
      33901: inst = 32'h10408000;
      33902: inst = 32'hc4047f8;
      33903: inst = 32'h8220000;
      33904: inst = 32'h10408000;
      33905: inst = 32'hc40480c;
      33906: inst = 32'h8220000;
      33907: inst = 32'h10408000;
      33908: inst = 32'hc404835;
      33909: inst = 32'h8220000;
      33910: inst = 32'h10408000;
      33911: inst = 32'hc404844;
      33912: inst = 32'h8220000;
      33913: inst = 32'h10408000;
      33914: inst = 32'hc40484c;
      33915: inst = 32'h8220000;
      33916: inst = 32'h10408000;
      33917: inst = 32'hc40485b;
      33918: inst = 32'h8220000;
      33919: inst = 32'h10408000;
      33920: inst = 32'hc404862;
      33921: inst = 32'h8220000;
      33922: inst = 32'h10408000;
      33923: inst = 32'hc40486f;
      33924: inst = 32'h8220000;
      33925: inst = 32'h10408000;
      33926: inst = 32'hc404895;
      33927: inst = 32'h8220000;
      33928: inst = 32'h10408000;
      33929: inst = 32'hc40489d;
      33930: inst = 32'h8220000;
      33931: inst = 32'h10408000;
      33932: inst = 32'hc4048a4;
      33933: inst = 32'h8220000;
      33934: inst = 32'h10408000;
      33935: inst = 32'hc4048c0;
      33936: inst = 32'h8220000;
      33937: inst = 32'h10408000;
      33938: inst = 32'hc4048c2;
      33939: inst = 32'h8220000;
      33940: inst = 32'h10408000;
      33941: inst = 32'hc4048f5;
      33942: inst = 32'h8220000;
      33943: inst = 32'h10408000;
      33944: inst = 32'hc4048fd;
      33945: inst = 32'h8220000;
      33946: inst = 32'h10408000;
      33947: inst = 32'hc404904;
      33948: inst = 32'h8220000;
      33949: inst = 32'h10408000;
      33950: inst = 32'hc404908;
      33951: inst = 32'h8220000;
      33952: inst = 32'h10408000;
      33953: inst = 32'hc404917;
      33954: inst = 32'h8220000;
      33955: inst = 32'h10408000;
      33956: inst = 32'hc404920;
      33957: inst = 32'h8220000;
      33958: inst = 32'h10408000;
      33959: inst = 32'hc404922;
      33960: inst = 32'h8220000;
      33961: inst = 32'h10408000;
      33962: inst = 32'hc40492b;
      33963: inst = 32'h8220000;
      33964: inst = 32'h10408000;
      33965: inst = 32'hc404955;
      33966: inst = 32'h8220000;
      33967: inst = 32'h10408000;
      33968: inst = 32'hc40495d;
      33969: inst = 32'h8220000;
      33970: inst = 32'h10408000;
      33971: inst = 32'hc404964;
      33972: inst = 32'h8220000;
      33973: inst = 32'h10408000;
      33974: inst = 32'hc404980;
      33975: inst = 32'h8220000;
      33976: inst = 32'h10408000;
      33977: inst = 32'hc404982;
      33978: inst = 32'h8220000;
      33979: inst = 32'h10408000;
      33980: inst = 32'hc4049b0;
      33981: inst = 32'h8220000;
      33982: inst = 32'h10408000;
      33983: inst = 32'hc4049b7;
      33984: inst = 32'h8220000;
      33985: inst = 32'h10408000;
      33986: inst = 32'hc4049bc;
      33987: inst = 32'h8220000;
      33988: inst = 32'h10408000;
      33989: inst = 32'hc4049c6;
      33990: inst = 32'h8220000;
      33991: inst = 32'h10408000;
      33992: inst = 32'hc4049d5;
      33993: inst = 32'h8220000;
      33994: inst = 32'h10408000;
      33995: inst = 32'hc4049df;
      33996: inst = 32'h8220000;
      33997: inst = 32'h10408000;
      33998: inst = 32'hc4049e4;
      33999: inst = 32'h8220000;
      34000: inst = 32'h10408000;
      34001: inst = 32'hc404d70;
      34002: inst = 32'h8220000;
      34003: inst = 32'h10408000;
      34004: inst = 32'hc404d81;
      34005: inst = 32'h8220000;
      34006: inst = 32'h10408000;
      34007: inst = 32'hc404d8b;
      34008: inst = 32'h8220000;
      34009: inst = 32'h10408000;
      34010: inst = 32'hc404d9f;
      34011: inst = 32'h8220000;
      34012: inst = 32'h10408000;
      34013: inst = 32'hc404da4;
      34014: inst = 32'h8220000;
      34015: inst = 32'h10408000;
      34016: inst = 32'hc404db1;
      34017: inst = 32'h8220000;
      34018: inst = 32'h10408000;
      34019: inst = 32'hc404dd0;
      34020: inst = 32'h8220000;
      34021: inst = 32'h10408000;
      34022: inst = 32'hc404de1;
      34023: inst = 32'h8220000;
      34024: inst = 32'h10408000;
      34025: inst = 32'hc404deb;
      34026: inst = 32'h8220000;
      34027: inst = 32'h10408000;
      34028: inst = 32'hc404dff;
      34029: inst = 32'h8220000;
      34030: inst = 32'h10408000;
      34031: inst = 32'hc404e04;
      34032: inst = 32'h8220000;
      34033: inst = 32'h10408000;
      34034: inst = 32'hc404e11;
      34035: inst = 32'h8220000;
      34036: inst = 32'h10408000;
      34037: inst = 32'hc404e2f;
      34038: inst = 32'h8220000;
      34039: inst = 32'h10408000;
      34040: inst = 32'hc404e30;
      34041: inst = 32'h8220000;
      34042: inst = 32'h10408000;
      34043: inst = 32'hc404e3e;
      34044: inst = 32'h8220000;
      34045: inst = 32'h10408000;
      34046: inst = 32'hc404e71;
      34047: inst = 32'h8220000;
      34048: inst = 32'h10408000;
      34049: inst = 32'hc404e90;
      34050: inst = 32'h8220000;
      34051: inst = 32'h10408000;
      34052: inst = 32'hc404e9a;
      34053: inst = 32'h8220000;
      34054: inst = 32'h10408000;
      34055: inst = 32'hc404e9e;
      34056: inst = 32'h8220000;
      34057: inst = 32'h10408000;
      34058: inst = 32'hc404ea1;
      34059: inst = 32'h8220000;
      34060: inst = 32'h10408000;
      34061: inst = 32'hc404eab;
      34062: inst = 32'h8220000;
      34063: inst = 32'h10408000;
      34064: inst = 32'hc404eb8;
      34065: inst = 32'h8220000;
      34066: inst = 32'h10408000;
      34067: inst = 32'hc404ebc;
      34068: inst = 32'h8220000;
      34069: inst = 32'h10408000;
      34070: inst = 32'hc404ebf;
      34071: inst = 32'h8220000;
      34072: inst = 32'h10408000;
      34073: inst = 32'hc404ec4;
      34074: inst = 32'h8220000;
      34075: inst = 32'h10408000;
      34076: inst = 32'hc404ec7;
      34077: inst = 32'h8220000;
      34078: inst = 32'h10408000;
      34079: inst = 32'hc404ecb;
      34080: inst = 32'h8220000;
      34081: inst = 32'h10408000;
      34082: inst = 32'hc404ecc;
      34083: inst = 32'h8220000;
      34084: inst = 32'h10408000;
      34085: inst = 32'hc404ed1;
      34086: inst = 32'h8220000;
      34087: inst = 32'h10408000;
      34088: inst = 32'hc404ef0;
      34089: inst = 32'h8220000;
      34090: inst = 32'h10408000;
      34091: inst = 32'hc404efe;
      34092: inst = 32'h8220000;
      34093: inst = 32'h10408000;
      34094: inst = 32'hc404f01;
      34095: inst = 32'h8220000;
      34096: inst = 32'h10408000;
      34097: inst = 32'hc404f0b;
      34098: inst = 32'h8220000;
      34099: inst = 32'h10408000;
      34100: inst = 32'hc404f1c;
      34101: inst = 32'h8220000;
      34102: inst = 32'h10408000;
      34103: inst = 32'hc404f1f;
      34104: inst = 32'h8220000;
      34105: inst = 32'h10408000;
      34106: inst = 32'hc404f24;
      34107: inst = 32'h8220000;
      34108: inst = 32'h10408000;
      34109: inst = 32'hc404f2b;
      34110: inst = 32'h8220000;
      34111: inst = 32'h10408000;
      34112: inst = 32'hc404f31;
      34113: inst = 32'h8220000;
      34114: inst = 32'h10408000;
      34115: inst = 32'hc404f32;
      34116: inst = 32'h8220000;
      34117: inst = 32'h10408000;
      34118: inst = 32'hc404f50;
      34119: inst = 32'h8220000;
      34120: inst = 32'h10408000;
      34121: inst = 32'hc404f5e;
      34122: inst = 32'h8220000;
      34123: inst = 32'h10408000;
      34124: inst = 32'hc404f61;
      34125: inst = 32'h8220000;
      34126: inst = 32'h10408000;
      34127: inst = 32'hc404f6b;
      34128: inst = 32'h8220000;
      34129: inst = 32'h10408000;
      34130: inst = 32'hc404f7c;
      34131: inst = 32'h8220000;
      34132: inst = 32'h10408000;
      34133: inst = 32'hc404f7f;
      34134: inst = 32'h8220000;
      34135: inst = 32'h10408000;
      34136: inst = 32'hc404f84;
      34137: inst = 32'h8220000;
      34138: inst = 32'h10408000;
      34139: inst = 32'hc404f8b;
      34140: inst = 32'h8220000;
      34141: inst = 32'h10408000;
      34142: inst = 32'hc404f91;
      34143: inst = 32'h8220000;
      34144: inst = 32'h10408000;
      34145: inst = 32'hc404f92;
      34146: inst = 32'h8220000;
      34147: inst = 32'h10408000;
      34148: inst = 32'hc404f94;
      34149: inst = 32'h8220000;
      34150: inst = 32'h10408000;
      34151: inst = 32'hc404fb0;
      34152: inst = 32'h8220000;
      34153: inst = 32'h10408000;
      34154: inst = 32'hc404fbe;
      34155: inst = 32'h8220000;
      34156: inst = 32'h10408000;
      34157: inst = 32'hc404fc1;
      34158: inst = 32'h8220000;
      34159: inst = 32'h10408000;
      34160: inst = 32'hc404fcb;
      34161: inst = 32'h8220000;
      34162: inst = 32'h10408000;
      34163: inst = 32'hc404fdc;
      34164: inst = 32'h8220000;
      34165: inst = 32'h10408000;
      34166: inst = 32'hc404fdf;
      34167: inst = 32'h8220000;
      34168: inst = 32'h10408000;
      34169: inst = 32'hc404fe4;
      34170: inst = 32'h8220000;
      34171: inst = 32'h10408000;
      34172: inst = 32'hc404feb;
      34173: inst = 32'h8220000;
      34174: inst = 32'h10408000;
      34175: inst = 32'hc404ff1;
      34176: inst = 32'h8220000;
      34177: inst = 32'h10408000;
      34178: inst = 32'hc40500b;
      34179: inst = 32'h8220000;
      34180: inst = 32'h10408000;
      34181: inst = 32'hc405011;
      34182: inst = 32'h8220000;
      34183: inst = 32'h10408000;
      34184: inst = 32'hc405016;
      34185: inst = 32'h8220000;
      34186: inst = 32'h10408000;
      34187: inst = 32'hc405018;
      34188: inst = 32'h8220000;
      34189: inst = 32'h10408000;
      34190: inst = 32'hc40501c;
      34191: inst = 32'h8220000;
      34192: inst = 32'h10408000;
      34193: inst = 32'hc40501d;
      34194: inst = 32'h8220000;
      34195: inst = 32'h10408000;
      34196: inst = 32'hc405022;
      34197: inst = 32'h8220000;
      34198: inst = 32'h10408000;
      34199: inst = 32'hc40502c;
      34200: inst = 32'h8220000;
      34201: inst = 32'h10408000;
      34202: inst = 32'hc40502f;
      34203: inst = 32'h8220000;
      34204: inst = 32'h10408000;
      34205: inst = 32'hc405031;
      34206: inst = 32'h8220000;
      34207: inst = 32'h10408000;
      34208: inst = 32'hc405040;
      34209: inst = 32'h8220000;
      34210: inst = 32'h10408000;
      34211: inst = 32'hc405045;
      34212: inst = 32'h8220000;
      34213: inst = 32'h10408000;
      34214: inst = 32'hc405052;
      34215: inst = 32'h8220000;
      34216: inst = 32'hc20ffff;
      34217: inst = 32'h10408000;
      34218: inst = 32'hc404fec;
      34219: inst = 32'h8220000;
      34220: inst = 32'h58000000;
      34221: inst = 32'h13e0ffff;
      34222: inst = 32'h13e00000;
      34223: inst = 32'hfe085c4;
      34224: inst = 32'h5be00000;
      34225: inst = 32'h13e0ffff;
      34226: inst = 32'h13e00000;
      34227: inst = 32'hfe0882f;
      34228: inst = 32'h5be00000;
      34229: inst = 32'h13e0ffff;
      34230: inst = 32'h13e00000;
      34231: inst = 32'hfe0882f;
      34232: inst = 32'h5be00000;
      34233: inst = 32'h13e0ffff;
      34234: inst = 32'h13e00000;
      34235: inst = 32'hfe086ff;
      34236: inst = 32'h5be00000;
      34237: inst = 32'h13e0ffff;
      34238: inst = 32'h13e00000;
      34239: inst = 32'hfe086ff;
      34240: inst = 32'h5be00000;
      34241: inst = 32'h13e00000;
      34242: inst = 32'hfe085c4;
      34243: inst = 32'h5be00000;
      34244: inst = 32'hc6018c3;
      34245: inst = 32'h10408000;
      34246: inst = 32'hc40496b;
      34247: inst = 32'h8620000;
      34248: inst = 32'h10408000;
      34249: inst = 32'hc40496c;
      34250: inst = 32'h8620000;
      34251: inst = 32'h10408000;
      34252: inst = 32'hc40496d;
      34253: inst = 32'h8620000;
      34254: inst = 32'h10408000;
      34255: inst = 32'hc40496e;
      34256: inst = 32'h8620000;
      34257: inst = 32'h10408000;
      34258: inst = 32'hc40496f;
      34259: inst = 32'h8620000;
      34260: inst = 32'h10408000;
      34261: inst = 32'hc404970;
      34262: inst = 32'h8620000;
      34263: inst = 32'h10408000;
      34264: inst = 32'hc404971;
      34265: inst = 32'h8620000;
      34266: inst = 32'h10408000;
      34267: inst = 32'hc404972;
      34268: inst = 32'h8620000;
      34269: inst = 32'h10408000;
      34270: inst = 32'hc404973;
      34271: inst = 32'h8620000;
      34272: inst = 32'h10408000;
      34273: inst = 32'hc404974;
      34274: inst = 32'h8620000;
      34275: inst = 32'h10408000;
      34276: inst = 32'hc4049cb;
      34277: inst = 32'h8620000;
      34278: inst = 32'h10408000;
      34279: inst = 32'hc4049cc;
      34280: inst = 32'h8620000;
      34281: inst = 32'h10408000;
      34282: inst = 32'hc4049cd;
      34283: inst = 32'h8620000;
      34284: inst = 32'h10408000;
      34285: inst = 32'hc4049ce;
      34286: inst = 32'h8620000;
      34287: inst = 32'h10408000;
      34288: inst = 32'hc4049cf;
      34289: inst = 32'h8620000;
      34290: inst = 32'h10408000;
      34291: inst = 32'hc4049d0;
      34292: inst = 32'h8620000;
      34293: inst = 32'h10408000;
      34294: inst = 32'hc4049d1;
      34295: inst = 32'h8620000;
      34296: inst = 32'h10408000;
      34297: inst = 32'hc4049d2;
      34298: inst = 32'h8620000;
      34299: inst = 32'h10408000;
      34300: inst = 32'hc4049d3;
      34301: inst = 32'h8620000;
      34302: inst = 32'h10408000;
      34303: inst = 32'hc4049d4;
      34304: inst = 32'h8620000;
      34305: inst = 32'h10408000;
      34306: inst = 32'hc404a2b;
      34307: inst = 32'h8620000;
      34308: inst = 32'h10408000;
      34309: inst = 32'hc404a34;
      34310: inst = 32'h8620000;
      34311: inst = 32'h10408000;
      34312: inst = 32'hc404a8b;
      34313: inst = 32'h8620000;
      34314: inst = 32'h10408000;
      34315: inst = 32'hc404a8d;
      34316: inst = 32'h8620000;
      34317: inst = 32'h10408000;
      34318: inst = 32'hc404a92;
      34319: inst = 32'h8620000;
      34320: inst = 32'h10408000;
      34321: inst = 32'hc404a94;
      34322: inst = 32'h8620000;
      34323: inst = 32'h10408000;
      34324: inst = 32'hc404aeb;
      34325: inst = 32'h8620000;
      34326: inst = 32'h10408000;
      34327: inst = 32'hc404aed;
      34328: inst = 32'h8620000;
      34329: inst = 32'h10408000;
      34330: inst = 32'hc404af2;
      34331: inst = 32'h8620000;
      34332: inst = 32'h10408000;
      34333: inst = 32'hc404af4;
      34334: inst = 32'h8620000;
      34335: inst = 32'h10408000;
      34336: inst = 32'hc404b4b;
      34337: inst = 32'h8620000;
      34338: inst = 32'h10408000;
      34339: inst = 32'hc404b54;
      34340: inst = 32'h8620000;
      34341: inst = 32'h10408000;
      34342: inst = 32'hc404bab;
      34343: inst = 32'h8620000;
      34344: inst = 32'h10408000;
      34345: inst = 32'hc404bb4;
      34346: inst = 32'h8620000;
      34347: inst = 32'hc60f4ce;
      34348: inst = 32'h10408000;
      34349: inst = 32'hc404a2c;
      34350: inst = 32'h8620000;
      34351: inst = 32'h10408000;
      34352: inst = 32'hc404a2d;
      34353: inst = 32'h8620000;
      34354: inst = 32'h10408000;
      34355: inst = 32'hc404a2e;
      34356: inst = 32'h8620000;
      34357: inst = 32'h10408000;
      34358: inst = 32'hc404a2f;
      34359: inst = 32'h8620000;
      34360: inst = 32'h10408000;
      34361: inst = 32'hc404a30;
      34362: inst = 32'h8620000;
      34363: inst = 32'h10408000;
      34364: inst = 32'hc404a31;
      34365: inst = 32'h8620000;
      34366: inst = 32'h10408000;
      34367: inst = 32'hc404a32;
      34368: inst = 32'h8620000;
      34369: inst = 32'h10408000;
      34370: inst = 32'hc404a33;
      34371: inst = 32'h8620000;
      34372: inst = 32'h10408000;
      34373: inst = 32'hc404a8c;
      34374: inst = 32'h8620000;
      34375: inst = 32'h10408000;
      34376: inst = 32'hc404a8e;
      34377: inst = 32'h8620000;
      34378: inst = 32'h10408000;
      34379: inst = 32'hc404a8f;
      34380: inst = 32'h8620000;
      34381: inst = 32'h10408000;
      34382: inst = 32'hc404a90;
      34383: inst = 32'h8620000;
      34384: inst = 32'h10408000;
      34385: inst = 32'hc404a91;
      34386: inst = 32'h8620000;
      34387: inst = 32'h10408000;
      34388: inst = 32'hc404a93;
      34389: inst = 32'h8620000;
      34390: inst = 32'h10408000;
      34391: inst = 32'hc404aec;
      34392: inst = 32'h8620000;
      34393: inst = 32'h10408000;
      34394: inst = 32'hc404aee;
      34395: inst = 32'h8620000;
      34396: inst = 32'h10408000;
      34397: inst = 32'hc404aef;
      34398: inst = 32'h8620000;
      34399: inst = 32'h10408000;
      34400: inst = 32'hc404af0;
      34401: inst = 32'h8620000;
      34402: inst = 32'h10408000;
      34403: inst = 32'hc404af1;
      34404: inst = 32'h8620000;
      34405: inst = 32'h10408000;
      34406: inst = 32'hc404af3;
      34407: inst = 32'h8620000;
      34408: inst = 32'h10408000;
      34409: inst = 32'hc404b4c;
      34410: inst = 32'h8620000;
      34411: inst = 32'h10408000;
      34412: inst = 32'hc404b4d;
      34413: inst = 32'h8620000;
      34414: inst = 32'h10408000;
      34415: inst = 32'hc404b4e;
      34416: inst = 32'h8620000;
      34417: inst = 32'h10408000;
      34418: inst = 32'hc404b4f;
      34419: inst = 32'h8620000;
      34420: inst = 32'h10408000;
      34421: inst = 32'hc404b50;
      34422: inst = 32'h8620000;
      34423: inst = 32'h10408000;
      34424: inst = 32'hc404b51;
      34425: inst = 32'h8620000;
      34426: inst = 32'h10408000;
      34427: inst = 32'hc404b52;
      34428: inst = 32'h8620000;
      34429: inst = 32'h10408000;
      34430: inst = 32'hc404b53;
      34431: inst = 32'h8620000;
      34432: inst = 32'h10408000;
      34433: inst = 32'hc404bac;
      34434: inst = 32'h8620000;
      34435: inst = 32'h10408000;
      34436: inst = 32'hc404bad;
      34437: inst = 32'h8620000;
      34438: inst = 32'h10408000;
      34439: inst = 32'hc404bae;
      34440: inst = 32'h8620000;
      34441: inst = 32'h10408000;
      34442: inst = 32'hc404baf;
      34443: inst = 32'h8620000;
      34444: inst = 32'h10408000;
      34445: inst = 32'hc404bb0;
      34446: inst = 32'h8620000;
      34447: inst = 32'h10408000;
      34448: inst = 32'hc404bb1;
      34449: inst = 32'h8620000;
      34450: inst = 32'h10408000;
      34451: inst = 32'hc404bb2;
      34452: inst = 32'h8620000;
      34453: inst = 32'h10408000;
      34454: inst = 32'hc404bb3;
      34455: inst = 32'h8620000;
      34456: inst = 32'h10408000;
      34457: inst = 32'hc404c6b;
      34458: inst = 32'h8620000;
      34459: inst = 32'h10408000;
      34460: inst = 32'hc404c6c;
      34461: inst = 32'h8620000;
      34462: inst = 32'h10408000;
      34463: inst = 32'hc404c73;
      34464: inst = 32'h8620000;
      34465: inst = 32'h10408000;
      34466: inst = 32'hc404c74;
      34467: inst = 32'h8620000;
      34468: inst = 32'h10408000;
      34469: inst = 32'hc404dee;
      34470: inst = 32'h8620000;
      34471: inst = 32'h10408000;
      34472: inst = 32'hc404df1;
      34473: inst = 32'h8620000;
      34474: inst = 32'hc607800;
      34475: inst = 32'h10408000;
      34476: inst = 32'hc404c0d;
      34477: inst = 32'h8620000;
      34478: inst = 32'h10408000;
      34479: inst = 32'hc404c0e;
      34480: inst = 32'h8620000;
      34481: inst = 32'h10408000;
      34482: inst = 32'hc404c11;
      34483: inst = 32'h8620000;
      34484: inst = 32'h10408000;
      34485: inst = 32'hc404c12;
      34486: inst = 32'h8620000;
      34487: inst = 32'hc60a000;
      34488: inst = 32'h10408000;
      34489: inst = 32'hc404c0f;
      34490: inst = 32'h8620000;
      34491: inst = 32'h10408000;
      34492: inst = 32'hc404c10;
      34493: inst = 32'h8620000;
      34494: inst = 32'h10408000;
      34495: inst = 32'hc404c6d;
      34496: inst = 32'h8620000;
      34497: inst = 32'h10408000;
      34498: inst = 32'hc404c6e;
      34499: inst = 32'h8620000;
      34500: inst = 32'h10408000;
      34501: inst = 32'hc404c6f;
      34502: inst = 32'h8620000;
      34503: inst = 32'h10408000;
      34504: inst = 32'hc404c70;
      34505: inst = 32'h8620000;
      34506: inst = 32'h10408000;
      34507: inst = 32'hc404c71;
      34508: inst = 32'h8620000;
      34509: inst = 32'h10408000;
      34510: inst = 32'hc404c72;
      34511: inst = 32'h8620000;
      34512: inst = 32'h10408000;
      34513: inst = 32'hc404ccd;
      34514: inst = 32'h8620000;
      34515: inst = 32'h10408000;
      34516: inst = 32'hc404cce;
      34517: inst = 32'h8620000;
      34518: inst = 32'h10408000;
      34519: inst = 32'hc404ccf;
      34520: inst = 32'h8620000;
      34521: inst = 32'h10408000;
      34522: inst = 32'hc404cd0;
      34523: inst = 32'h8620000;
      34524: inst = 32'h10408000;
      34525: inst = 32'hc404cd1;
      34526: inst = 32'h8620000;
      34527: inst = 32'h10408000;
      34528: inst = 32'hc404cd2;
      34529: inst = 32'h8620000;
      34530: inst = 32'hc6010ac;
      34531: inst = 32'h10408000;
      34532: inst = 32'hc404d2d;
      34533: inst = 32'h8620000;
      34534: inst = 32'h10408000;
      34535: inst = 32'hc404d2e;
      34536: inst = 32'h8620000;
      34537: inst = 32'h10408000;
      34538: inst = 32'hc404d2f;
      34539: inst = 32'h8620000;
      34540: inst = 32'h10408000;
      34541: inst = 32'hc404d30;
      34542: inst = 32'h8620000;
      34543: inst = 32'h10408000;
      34544: inst = 32'hc404d31;
      34545: inst = 32'h8620000;
      34546: inst = 32'h10408000;
      34547: inst = 32'hc404d32;
      34548: inst = 32'h8620000;
      34549: inst = 32'hc60d42c;
      34550: inst = 32'h10408000;
      34551: inst = 32'hc404d8e;
      34552: inst = 32'h8620000;
      34553: inst = 32'h10408000;
      34554: inst = 32'hc404d91;
      34555: inst = 32'h8620000;
      34556: inst = 32'h13e00000;
      34557: inst = 32'hfe0895f;
      34558: inst = 32'h5be00000;
      34559: inst = 32'hc6018c3;
      34560: inst = 32'h10408000;
      34561: inst = 32'hc40496b;
      34562: inst = 32'h8620000;
      34563: inst = 32'h10408000;
      34564: inst = 32'hc40496c;
      34565: inst = 32'h8620000;
      34566: inst = 32'h10408000;
      34567: inst = 32'hc40496d;
      34568: inst = 32'h8620000;
      34569: inst = 32'h10408000;
      34570: inst = 32'hc40496e;
      34571: inst = 32'h8620000;
      34572: inst = 32'h10408000;
      34573: inst = 32'hc40496f;
      34574: inst = 32'h8620000;
      34575: inst = 32'h10408000;
      34576: inst = 32'hc404970;
      34577: inst = 32'h8620000;
      34578: inst = 32'h10408000;
      34579: inst = 32'hc404971;
      34580: inst = 32'h8620000;
      34581: inst = 32'h10408000;
      34582: inst = 32'hc404972;
      34583: inst = 32'h8620000;
      34584: inst = 32'h10408000;
      34585: inst = 32'hc404973;
      34586: inst = 32'h8620000;
      34587: inst = 32'h10408000;
      34588: inst = 32'hc404974;
      34589: inst = 32'h8620000;
      34590: inst = 32'h10408000;
      34591: inst = 32'hc4049cb;
      34592: inst = 32'h8620000;
      34593: inst = 32'h10408000;
      34594: inst = 32'hc4049cc;
      34595: inst = 32'h8620000;
      34596: inst = 32'h10408000;
      34597: inst = 32'hc4049cd;
      34598: inst = 32'h8620000;
      34599: inst = 32'h10408000;
      34600: inst = 32'hc4049ce;
      34601: inst = 32'h8620000;
      34602: inst = 32'h10408000;
      34603: inst = 32'hc4049cf;
      34604: inst = 32'h8620000;
      34605: inst = 32'h10408000;
      34606: inst = 32'hc4049d0;
      34607: inst = 32'h8620000;
      34608: inst = 32'h10408000;
      34609: inst = 32'hc4049d1;
      34610: inst = 32'h8620000;
      34611: inst = 32'h10408000;
      34612: inst = 32'hc4049d2;
      34613: inst = 32'h8620000;
      34614: inst = 32'h10408000;
      34615: inst = 32'hc4049d3;
      34616: inst = 32'h8620000;
      34617: inst = 32'h10408000;
      34618: inst = 32'hc4049d4;
      34619: inst = 32'h8620000;
      34620: inst = 32'h10408000;
      34621: inst = 32'hc404a2b;
      34622: inst = 32'h8620000;
      34623: inst = 32'h10408000;
      34624: inst = 32'hc404a2c;
      34625: inst = 32'h8620000;
      34626: inst = 32'h10408000;
      34627: inst = 32'hc404a8b;
      34628: inst = 32'h8620000;
      34629: inst = 32'h10408000;
      34630: inst = 32'hc404a93;
      34631: inst = 32'h8620000;
      34632: inst = 32'h10408000;
      34633: inst = 32'hc404aeb;
      34634: inst = 32'h8620000;
      34635: inst = 32'h10408000;
      34636: inst = 32'hc404af3;
      34637: inst = 32'h8620000;
      34638: inst = 32'h10408000;
      34639: inst = 32'hc404b4b;
      34640: inst = 32'h8620000;
      34641: inst = 32'h10408000;
      34642: inst = 32'hc404b4c;
      34643: inst = 32'h8620000;
      34644: inst = 32'h10408000;
      34645: inst = 32'hc404bab;
      34646: inst = 32'h8620000;
      34647: inst = 32'h10408000;
      34648: inst = 32'hc404bac;
      34649: inst = 32'h8620000;
      34650: inst = 32'hc60d42c;
      34651: inst = 32'h10408000;
      34652: inst = 32'hc404a2d;
      34653: inst = 32'h8620000;
      34654: inst = 32'h10408000;
      34655: inst = 32'hc404a2e;
      34656: inst = 32'h8620000;
      34657: inst = 32'h10408000;
      34658: inst = 32'hc404a2f;
      34659: inst = 32'h8620000;
      34660: inst = 32'h10408000;
      34661: inst = 32'hc404a30;
      34662: inst = 32'h8620000;
      34663: inst = 32'h10408000;
      34664: inst = 32'hc404a31;
      34665: inst = 32'h8620000;
      34666: inst = 32'h10408000;
      34667: inst = 32'hc404a32;
      34668: inst = 32'h8620000;
      34669: inst = 32'h10408000;
      34670: inst = 32'hc404a33;
      34671: inst = 32'h8620000;
      34672: inst = 32'h10408000;
      34673: inst = 32'hc404a34;
      34674: inst = 32'h8620000;
      34675: inst = 32'h10408000;
      34676: inst = 32'hc404b4d;
      34677: inst = 32'h8620000;
      34678: inst = 32'h10408000;
      34679: inst = 32'hc404bad;
      34680: inst = 32'h8620000;
      34681: inst = 32'h10408000;
      34682: inst = 32'hc404d8e;
      34683: inst = 32'h8620000;
      34684: inst = 32'h10408000;
      34685: inst = 32'hc404d91;
      34686: inst = 32'h8620000;
      34687: inst = 32'hc60f4ce;
      34688: inst = 32'h10408000;
      34689: inst = 32'hc404a8c;
      34690: inst = 32'h8620000;
      34691: inst = 32'h10408000;
      34692: inst = 32'hc404a8d;
      34693: inst = 32'h8620000;
      34694: inst = 32'h10408000;
      34695: inst = 32'hc404a8e;
      34696: inst = 32'h8620000;
      34697: inst = 32'h10408000;
      34698: inst = 32'hc404a8f;
      34699: inst = 32'h8620000;
      34700: inst = 32'h10408000;
      34701: inst = 32'hc404a90;
      34702: inst = 32'h8620000;
      34703: inst = 32'h10408000;
      34704: inst = 32'hc404a91;
      34705: inst = 32'h8620000;
      34706: inst = 32'h10408000;
      34707: inst = 32'hc404a92;
      34708: inst = 32'h8620000;
      34709: inst = 32'h10408000;
      34710: inst = 32'hc404a94;
      34711: inst = 32'h8620000;
      34712: inst = 32'h10408000;
      34713: inst = 32'hc404aec;
      34714: inst = 32'h8620000;
      34715: inst = 32'h10408000;
      34716: inst = 32'hc404aed;
      34717: inst = 32'h8620000;
      34718: inst = 32'h10408000;
      34719: inst = 32'hc404aee;
      34720: inst = 32'h8620000;
      34721: inst = 32'h10408000;
      34722: inst = 32'hc404aef;
      34723: inst = 32'h8620000;
      34724: inst = 32'h10408000;
      34725: inst = 32'hc404af0;
      34726: inst = 32'h8620000;
      34727: inst = 32'h10408000;
      34728: inst = 32'hc404af1;
      34729: inst = 32'h8620000;
      34730: inst = 32'h10408000;
      34731: inst = 32'hc404af2;
      34732: inst = 32'h8620000;
      34733: inst = 32'h10408000;
      34734: inst = 32'hc404af4;
      34735: inst = 32'h8620000;
      34736: inst = 32'h10408000;
      34737: inst = 32'hc404b4e;
      34738: inst = 32'h8620000;
      34739: inst = 32'h10408000;
      34740: inst = 32'hc404b4f;
      34741: inst = 32'h8620000;
      34742: inst = 32'h10408000;
      34743: inst = 32'hc404b50;
      34744: inst = 32'h8620000;
      34745: inst = 32'h10408000;
      34746: inst = 32'hc404b51;
      34747: inst = 32'h8620000;
      34748: inst = 32'h10408000;
      34749: inst = 32'hc404b52;
      34750: inst = 32'h8620000;
      34751: inst = 32'h10408000;
      34752: inst = 32'hc404b53;
      34753: inst = 32'h8620000;
      34754: inst = 32'h10408000;
      34755: inst = 32'hc404b54;
      34756: inst = 32'h8620000;
      34757: inst = 32'h10408000;
      34758: inst = 32'hc404bae;
      34759: inst = 32'h8620000;
      34760: inst = 32'h10408000;
      34761: inst = 32'hc404baf;
      34762: inst = 32'h8620000;
      34763: inst = 32'h10408000;
      34764: inst = 32'hc404bb0;
      34765: inst = 32'h8620000;
      34766: inst = 32'h10408000;
      34767: inst = 32'hc404bb1;
      34768: inst = 32'h8620000;
      34769: inst = 32'h10408000;
      34770: inst = 32'hc404bb2;
      34771: inst = 32'h8620000;
      34772: inst = 32'h10408000;
      34773: inst = 32'hc404bb3;
      34774: inst = 32'h8620000;
      34775: inst = 32'h10408000;
      34776: inst = 32'hc404bb4;
      34777: inst = 32'h8620000;
      34778: inst = 32'h10408000;
      34779: inst = 32'hc404c6f;
      34780: inst = 32'h8620000;
      34781: inst = 32'hc607841;
      34782: inst = 32'h10408000;
      34783: inst = 32'hc404c0d;
      34784: inst = 32'h8620000;
      34785: inst = 32'h10408000;
      34786: inst = 32'hc404c6d;
      34787: inst = 32'h8620000;
      34788: inst = 32'hc60a000;
      34789: inst = 32'h10408000;
      34790: inst = 32'hc404c0e;
      34791: inst = 32'h8620000;
      34792: inst = 32'h10408000;
      34793: inst = 32'hc404c0f;
      34794: inst = 32'h8620000;
      34795: inst = 32'h10408000;
      34796: inst = 32'hc404c10;
      34797: inst = 32'h8620000;
      34798: inst = 32'h10408000;
      34799: inst = 32'hc404c11;
      34800: inst = 32'h8620000;
      34801: inst = 32'h10408000;
      34802: inst = 32'hc404c12;
      34803: inst = 32'h8620000;
      34804: inst = 32'h10408000;
      34805: inst = 32'hc404c6e;
      34806: inst = 32'h8620000;
      34807: inst = 32'h10408000;
      34808: inst = 32'hc404c70;
      34809: inst = 32'h8620000;
      34810: inst = 32'h10408000;
      34811: inst = 32'hc404c71;
      34812: inst = 32'h8620000;
      34813: inst = 32'h10408000;
      34814: inst = 32'hc404c72;
      34815: inst = 32'h8620000;
      34816: inst = 32'h10408000;
      34817: inst = 32'hc404ccd;
      34818: inst = 32'h8620000;
      34819: inst = 32'h10408000;
      34820: inst = 32'hc404cce;
      34821: inst = 32'h8620000;
      34822: inst = 32'h10408000;
      34823: inst = 32'hc404ccf;
      34824: inst = 32'h8620000;
      34825: inst = 32'h10408000;
      34826: inst = 32'hc404cd0;
      34827: inst = 32'h8620000;
      34828: inst = 32'h10408000;
      34829: inst = 32'hc404cd1;
      34830: inst = 32'h8620000;
      34831: inst = 32'h10408000;
      34832: inst = 32'hc404cd2;
      34833: inst = 32'h8620000;
      34834: inst = 32'hc6010ac;
      34835: inst = 32'h10408000;
      34836: inst = 32'hc404d2d;
      34837: inst = 32'h8620000;
      34838: inst = 32'h10408000;
      34839: inst = 32'hc404d2e;
      34840: inst = 32'h8620000;
      34841: inst = 32'h10408000;
      34842: inst = 32'hc404d2f;
      34843: inst = 32'h8620000;
      34844: inst = 32'h10408000;
      34845: inst = 32'hc404d30;
      34846: inst = 32'h8620000;
      34847: inst = 32'h10408000;
      34848: inst = 32'hc404d31;
      34849: inst = 32'h8620000;
      34850: inst = 32'h10408000;
      34851: inst = 32'hc404d32;
      34852: inst = 32'h8620000;
      34853: inst = 32'h13e0ffff;
      34854: inst = 32'h13e00000;
      34855: inst = 32'hfe0882c;
      34856: inst = 32'h5be00000;
      34857: inst = 32'h13e00000;
      34858: inst = 32'hfe0895f;
      34859: inst = 32'h5be00000;
      34860: inst = 32'h13e00000;
      34861: inst = 32'hfe0895f;
      34862: inst = 32'h5be00000;
      34863: inst = 32'hc6018c3;
      34864: inst = 32'h10408000;
      34865: inst = 32'hc4049cb;
      34866: inst = 32'h8620000;
      34867: inst = 32'h10408000;
      34868: inst = 32'hc4049ca;
      34869: inst = 32'h8620000;
      34870: inst = 32'h10408000;
      34871: inst = 32'hc4049c9;
      34872: inst = 32'h8620000;
      34873: inst = 32'h10408000;
      34874: inst = 32'hc4049c8;
      34875: inst = 32'h8620000;
      34876: inst = 32'h10408000;
      34877: inst = 32'hc4049c7;
      34878: inst = 32'h8620000;
      34879: inst = 32'h10408000;
      34880: inst = 32'hc4049c6;
      34881: inst = 32'h8620000;
      34882: inst = 32'h10408000;
      34883: inst = 32'hc4049c5;
      34884: inst = 32'h8620000;
      34885: inst = 32'h10408000;
      34886: inst = 32'hc4049c4;
      34887: inst = 32'h8620000;
      34888: inst = 32'h10408000;
      34889: inst = 32'hc4049c3;
      34890: inst = 32'h8620000;
      34891: inst = 32'h10408000;
      34892: inst = 32'hc4049c2;
      34893: inst = 32'h8620000;
      34894: inst = 32'h10408000;
      34895: inst = 32'hc404a2b;
      34896: inst = 32'h8620000;
      34897: inst = 32'h10408000;
      34898: inst = 32'hc404a2a;
      34899: inst = 32'h8620000;
      34900: inst = 32'h10408000;
      34901: inst = 32'hc404a29;
      34902: inst = 32'h8620000;
      34903: inst = 32'h10408000;
      34904: inst = 32'hc404a28;
      34905: inst = 32'h8620000;
      34906: inst = 32'h10408000;
      34907: inst = 32'hc404a27;
      34908: inst = 32'h8620000;
      34909: inst = 32'h10408000;
      34910: inst = 32'hc404a26;
      34911: inst = 32'h8620000;
      34912: inst = 32'h10408000;
      34913: inst = 32'hc404a25;
      34914: inst = 32'h8620000;
      34915: inst = 32'h10408000;
      34916: inst = 32'hc404a24;
      34917: inst = 32'h8620000;
      34918: inst = 32'h10408000;
      34919: inst = 32'hc404a23;
      34920: inst = 32'h8620000;
      34921: inst = 32'h10408000;
      34922: inst = 32'hc404a22;
      34923: inst = 32'h8620000;
      34924: inst = 32'h10408000;
      34925: inst = 32'hc404a8b;
      34926: inst = 32'h8620000;
      34927: inst = 32'h10408000;
      34928: inst = 32'hc404a8a;
      34929: inst = 32'h8620000;
      34930: inst = 32'h10408000;
      34931: inst = 32'hc404aeb;
      34932: inst = 32'h8620000;
      34933: inst = 32'h10408000;
      34934: inst = 32'hc404ae3;
      34935: inst = 32'h8620000;
      34936: inst = 32'h10408000;
      34937: inst = 32'hc404b4b;
      34938: inst = 32'h8620000;
      34939: inst = 32'h10408000;
      34940: inst = 32'hc404b43;
      34941: inst = 32'h8620000;
      34942: inst = 32'h10408000;
      34943: inst = 32'hc404bab;
      34944: inst = 32'h8620000;
      34945: inst = 32'h10408000;
      34946: inst = 32'hc404baa;
      34947: inst = 32'h8620000;
      34948: inst = 32'h10408000;
      34949: inst = 32'hc404c0b;
      34950: inst = 32'h8620000;
      34951: inst = 32'h10408000;
      34952: inst = 32'hc404c0a;
      34953: inst = 32'h8620000;
      34954: inst = 32'hc60d42c;
      34955: inst = 32'h10408000;
      34956: inst = 32'hc404a89;
      34957: inst = 32'h8620000;
      34958: inst = 32'h10408000;
      34959: inst = 32'hc404a88;
      34960: inst = 32'h8620000;
      34961: inst = 32'h10408000;
      34962: inst = 32'hc404a87;
      34963: inst = 32'h8620000;
      34964: inst = 32'h10408000;
      34965: inst = 32'hc404a86;
      34966: inst = 32'h8620000;
      34967: inst = 32'h10408000;
      34968: inst = 32'hc404a85;
      34969: inst = 32'h8620000;
      34970: inst = 32'h10408000;
      34971: inst = 32'hc404a84;
      34972: inst = 32'h8620000;
      34973: inst = 32'h10408000;
      34974: inst = 32'hc404a83;
      34975: inst = 32'h8620000;
      34976: inst = 32'h10408000;
      34977: inst = 32'hc404a82;
      34978: inst = 32'h8620000;
      34979: inst = 32'h10408000;
      34980: inst = 32'hc404ba9;
      34981: inst = 32'h8620000;
      34982: inst = 32'h10408000;
      34983: inst = 32'hc404c09;
      34984: inst = 32'h8620000;
      34985: inst = 32'h10408000;
      34986: inst = 32'hc404de8;
      34987: inst = 32'h8620000;
      34988: inst = 32'h10408000;
      34989: inst = 32'hc404de5;
      34990: inst = 32'h8620000;
      34991: inst = 32'hc60f4ce;
      34992: inst = 32'h10408000;
      34993: inst = 32'hc404aea;
      34994: inst = 32'h8620000;
      34995: inst = 32'h10408000;
      34996: inst = 32'hc404ae9;
      34997: inst = 32'h8620000;
      34998: inst = 32'h10408000;
      34999: inst = 32'hc404ae8;
      35000: inst = 32'h8620000;
      35001: inst = 32'h10408000;
      35002: inst = 32'hc404ae7;
      35003: inst = 32'h8620000;
      35004: inst = 32'h10408000;
      35005: inst = 32'hc404ae6;
      35006: inst = 32'h8620000;
      35007: inst = 32'h10408000;
      35008: inst = 32'hc404ae5;
      35009: inst = 32'h8620000;
      35010: inst = 32'h10408000;
      35011: inst = 32'hc404ae4;
      35012: inst = 32'h8620000;
      35013: inst = 32'h10408000;
      35014: inst = 32'hc404ae2;
      35015: inst = 32'h8620000;
      35016: inst = 32'h10408000;
      35017: inst = 32'hc404b4a;
      35018: inst = 32'h8620000;
      35019: inst = 32'h10408000;
      35020: inst = 32'hc404b49;
      35021: inst = 32'h8620000;
      35022: inst = 32'h10408000;
      35023: inst = 32'hc404b48;
      35024: inst = 32'h8620000;
      35025: inst = 32'h10408000;
      35026: inst = 32'hc404b47;
      35027: inst = 32'h8620000;
      35028: inst = 32'h10408000;
      35029: inst = 32'hc404b46;
      35030: inst = 32'h8620000;
      35031: inst = 32'h10408000;
      35032: inst = 32'hc404b45;
      35033: inst = 32'h8620000;
      35034: inst = 32'h10408000;
      35035: inst = 32'hc404b44;
      35036: inst = 32'h8620000;
      35037: inst = 32'h10408000;
      35038: inst = 32'hc404b42;
      35039: inst = 32'h8620000;
      35040: inst = 32'h10408000;
      35041: inst = 32'hc404ba8;
      35042: inst = 32'h8620000;
      35043: inst = 32'h10408000;
      35044: inst = 32'hc404ba7;
      35045: inst = 32'h8620000;
      35046: inst = 32'h10408000;
      35047: inst = 32'hc404ba6;
      35048: inst = 32'h8620000;
      35049: inst = 32'h10408000;
      35050: inst = 32'hc404ba5;
      35051: inst = 32'h8620000;
      35052: inst = 32'h10408000;
      35053: inst = 32'hc404ba4;
      35054: inst = 32'h8620000;
      35055: inst = 32'h10408000;
      35056: inst = 32'hc404ba3;
      35057: inst = 32'h8620000;
      35058: inst = 32'h10408000;
      35059: inst = 32'hc404ba2;
      35060: inst = 32'h8620000;
      35061: inst = 32'h10408000;
      35062: inst = 32'hc404c08;
      35063: inst = 32'h8620000;
      35064: inst = 32'h10408000;
      35065: inst = 32'hc404c07;
      35066: inst = 32'h8620000;
      35067: inst = 32'h10408000;
      35068: inst = 32'hc404c06;
      35069: inst = 32'h8620000;
      35070: inst = 32'h10408000;
      35071: inst = 32'hc404c05;
      35072: inst = 32'h8620000;
      35073: inst = 32'h10408000;
      35074: inst = 32'hc404c04;
      35075: inst = 32'h8620000;
      35076: inst = 32'h10408000;
      35077: inst = 32'hc404c03;
      35078: inst = 32'h8620000;
      35079: inst = 32'h10408000;
      35080: inst = 32'hc404c02;
      35081: inst = 32'h8620000;
      35082: inst = 32'h10408000;
      35083: inst = 32'hc404cc7;
      35084: inst = 32'h8620000;
      35085: inst = 32'hc607841;
      35086: inst = 32'h10408000;
      35087: inst = 32'hc404c69;
      35088: inst = 32'h8620000;
      35089: inst = 32'h10408000;
      35090: inst = 32'hc404cc9;
      35091: inst = 32'h8620000;
      35092: inst = 32'hc60a000;
      35093: inst = 32'h10408000;
      35094: inst = 32'hc404c68;
      35095: inst = 32'h8620000;
      35096: inst = 32'h10408000;
      35097: inst = 32'hc404c67;
      35098: inst = 32'h8620000;
      35099: inst = 32'h10408000;
      35100: inst = 32'hc404c66;
      35101: inst = 32'h8620000;
      35102: inst = 32'h10408000;
      35103: inst = 32'hc404c65;
      35104: inst = 32'h8620000;
      35105: inst = 32'h10408000;
      35106: inst = 32'hc404c64;
      35107: inst = 32'h8620000;
      35108: inst = 32'h10408000;
      35109: inst = 32'hc404cc8;
      35110: inst = 32'h8620000;
      35111: inst = 32'h10408000;
      35112: inst = 32'hc404cc6;
      35113: inst = 32'h8620000;
      35114: inst = 32'h10408000;
      35115: inst = 32'hc404cc5;
      35116: inst = 32'h8620000;
      35117: inst = 32'h10408000;
      35118: inst = 32'hc404cc4;
      35119: inst = 32'h8620000;
      35120: inst = 32'h10408000;
      35121: inst = 32'hc404d29;
      35122: inst = 32'h8620000;
      35123: inst = 32'h10408000;
      35124: inst = 32'hc404d28;
      35125: inst = 32'h8620000;
      35126: inst = 32'h10408000;
      35127: inst = 32'hc404d27;
      35128: inst = 32'h8620000;
      35129: inst = 32'h10408000;
      35130: inst = 32'hc404d26;
      35131: inst = 32'h8620000;
      35132: inst = 32'h10408000;
      35133: inst = 32'hc404d25;
      35134: inst = 32'h8620000;
      35135: inst = 32'h10408000;
      35136: inst = 32'hc404d24;
      35137: inst = 32'h8620000;
      35138: inst = 32'hc6010ac;
      35139: inst = 32'h10408000;
      35140: inst = 32'hc404d89;
      35141: inst = 32'h8620000;
      35142: inst = 32'h10408000;
      35143: inst = 32'hc404d88;
      35144: inst = 32'h8620000;
      35145: inst = 32'h10408000;
      35146: inst = 32'hc404d87;
      35147: inst = 32'h8620000;
      35148: inst = 32'h10408000;
      35149: inst = 32'hc404d86;
      35150: inst = 32'h8620000;
      35151: inst = 32'h10408000;
      35152: inst = 32'hc404d85;
      35153: inst = 32'h8620000;
      35154: inst = 32'h10408000;
      35155: inst = 32'hc404d84;
      35156: inst = 32'h8620000;
      35157: inst = 32'h13e0ffff;
      35158: inst = 32'h13e00000;
      35159: inst = 32'hfe0895c;
      35160: inst = 32'h5be00000;
      35161: inst = 32'h13e00000;
      35162: inst = 32'hfe0895f;
      35163: inst = 32'h5be00000;
      35164: inst = 32'h13e00000;
      35165: inst = 32'hfe0895f;
      35166: inst = 32'h5be00000;
      35167: inst = 32'h58000000;
      35168: inst = 32'h10408000;
      35169: inst = 32'hc400002;
      35170: inst = 32'h4420000;
      35171: inst = 32'h10600000;
      35172: inst = 32'hc600010;
      35173: inst = 32'h38421800;
      35174: inst = 32'h4042000f;
      35175: inst = 32'h1c40000f;
      35176: inst = 32'h58000000;
      35177: inst = 32'h58200000;
      35178: inst = 32'h11400000;
      35179: inst = 32'hd400000;
      35180: inst = 32'h11600000;
      35181: inst = 32'hd600060;
      35182: inst = 32'h11200000;
      35183: inst = 32'hd208973;
      35184: inst = 32'h13e00000;
      35185: inst = 32'hfe08f6a;
      35186: inst = 32'h5be00000;
      35187: inst = 32'h29ec0000;
      35188: inst = 32'h12000000;
      35189: inst = 32'he000001;
      35190: inst = 32'h3a0b8000;
      35191: inst = 32'h2def8000;
      35192: inst = 32'h11200000;
      35193: inst = 32'hd20897d;
      35194: inst = 32'h13e00000;
      35195: inst = 32'hfe08f5e;
      35196: inst = 32'h5be00000;
      35197: inst = 32'h2a0c0000;
      35198: inst = 32'h12200000;
      35199: inst = 32'he200040;
      35200: inst = 32'h12400000;
      35201: inst = 32'he400001;
      35202: inst = 32'h3a319000;
      35203: inst = 32'h2e108800;
      35204: inst = 32'h294a0001;
      35205: inst = 32'h24617800;
      35206: inst = 32'h24828000;
      35207: inst = 32'h10a00000;
      35208: inst = 32'hca00004;
      35209: inst = 32'h38632800;
      35210: inst = 32'h38842800;
      35211: inst = 32'h10a00000;
      35212: inst = 32'hca08990;
      35213: inst = 32'h13e00000;
      35214: inst = 32'hfe08998;
      35215: inst = 32'h5be00000;
      35216: inst = 32'h10a08000;
      35217: inst = 32'hca04061;
      35218: inst = 32'h8c50000;
      35219: inst = 32'h13e00000;
      35220: inst = 32'hfe0896c;
      35221: inst = 32'h1d401800;
      35222: inst = 32'h5be00000;
      35223: inst = 32'h58000000;
      35224: inst = 32'h13e0ffff;
      35225: inst = 32'h13e00000;
      35226: inst = 32'hfe089ff;
      35227: inst = 32'h5be00000;
      35228: inst = 32'h13e0ffff;
      35229: inst = 32'h13e00000;
      35230: inst = 32'hfe08a36;
      35231: inst = 32'h5be00000;
      35232: inst = 32'h13e0ffff;
      35233: inst = 32'h13e00000;
      35234: inst = 32'hfe08a6d;
      35235: inst = 32'h5be00000;
      35236: inst = 32'h13e0ffff;
      35237: inst = 32'h13e00000;
      35238: inst = 32'hfe08aa4;
      35239: inst = 32'h5be00000;
      35240: inst = 32'h13e0ffff;
      35241: inst = 32'h13e00000;
      35242: inst = 32'hfe08adb;
      35243: inst = 32'h5be00000;
      35244: inst = 32'h13e0ffff;
      35245: inst = 32'h13e00000;
      35246: inst = 32'hfe08b12;
      35247: inst = 32'h5be00000;
      35248: inst = 32'h13e0ffff;
      35249: inst = 32'h13e00000;
      35250: inst = 32'hfe08b49;
      35251: inst = 32'h5be00000;
      35252: inst = 32'h13e0ffff;
      35253: inst = 32'h13e00000;
      35254: inst = 32'hfe08b80;
      35255: inst = 32'h5be00000;
      35256: inst = 32'h13e0ffff;
      35257: inst = 32'h13e00000;
      35258: inst = 32'hfe08bb7;
      35259: inst = 32'h5be00000;
      35260: inst = 32'h13e0ffff;
      35261: inst = 32'h13e00000;
      35262: inst = 32'hfe08bee;
      35263: inst = 32'h5be00000;
      35264: inst = 32'h13e0ffff;
      35265: inst = 32'h13e00000;
      35266: inst = 32'hfe08c25;
      35267: inst = 32'h5be00000;
      35268: inst = 32'h13e0ffff;
      35269: inst = 32'h13e00000;
      35270: inst = 32'hfe08c5c;
      35271: inst = 32'h5be00000;
      35272: inst = 32'h13e0ffff;
      35273: inst = 32'h13e00000;
      35274: inst = 32'hfe08c93;
      35275: inst = 32'h5be00000;
      35276: inst = 32'h13e0ffff;
      35277: inst = 32'h13e00000;
      35278: inst = 32'hfe08cca;
      35279: inst = 32'h5be00000;
      35280: inst = 32'h13e0ffff;
      35281: inst = 32'h13e00000;
      35282: inst = 32'hfe08d01;
      35283: inst = 32'h5be00000;
      35284: inst = 32'h13e0ffff;
      35285: inst = 32'h13e00000;
      35286: inst = 32'hfe08d38;
      35287: inst = 32'h5be00000;
      35288: inst = 32'h13e0ffff;
      35289: inst = 32'h13e00000;
      35290: inst = 32'hfe08d6f;
      35291: inst = 32'h5be00000;
      35292: inst = 32'h13e0ffff;
      35293: inst = 32'h13e00000;
      35294: inst = 32'hfe08da6;
      35295: inst = 32'h5be00000;
      35296: inst = 32'h13e0ffff;
      35297: inst = 32'h13e00000;
      35298: inst = 32'hfe08ddd;
      35299: inst = 32'h5be00000;
      35300: inst = 32'h13e0ffff;
      35301: inst = 32'h13e00000;
      35302: inst = 32'hfe08e14;
      35303: inst = 32'h5be00000;
      35304: inst = 32'h13e0ffff;
      35305: inst = 32'h13e00000;
      35306: inst = 32'hfe08e4b;
      35307: inst = 32'h5be00000;
      35308: inst = 32'h13e0ffff;
      35309: inst = 32'h13e00000;
      35310: inst = 32'hfe08e82;
      35311: inst = 32'h5be00000;
      35312: inst = 32'h13e0ffff;
      35313: inst = 32'h13e00000;
      35314: inst = 32'hfe08eb9;
      35315: inst = 32'h5be00000;
      35316: inst = 32'h13e0ffff;
      35317: inst = 32'h13e00000;
      35318: inst = 32'hfe08ef0;
      35319: inst = 32'h5be00000;
      35320: inst = 32'h13e0ffff;
      35321: inst = 32'h13e00000;
      35322: inst = 32'hfe08f27;
      35323: inst = 32'h5be00000;
      35324: inst = 32'h10c00000;
      35325: inst = 32'hcc00000;
      35326: inst = 32'h58a00000;
      35327: inst = 32'h20800000;
      35328: inst = 32'h10c00000;
      35329: inst = 32'hcc06b50;
      35330: inst = 32'h20800001;
      35331: inst = 32'h10c00000;
      35332: inst = 32'hcc06b50;
      35333: inst = 32'h20800002;
      35334: inst = 32'h10c00000;
      35335: inst = 32'hcc06b50;
      35336: inst = 32'h20800003;
      35337: inst = 32'h10c00000;
      35338: inst = 32'hcc06b50;
      35339: inst = 32'h20800004;
      35340: inst = 32'h10c00000;
      35341: inst = 32'hcc06b50;
      35342: inst = 32'h20800005;
      35343: inst = 32'h10c00000;
      35344: inst = 32'hcc06b50;
      35345: inst = 32'h20800006;
      35346: inst = 32'h10c00000;
      35347: inst = 32'hcc06b50;
      35348: inst = 32'h20800007;
      35349: inst = 32'h10c00000;
      35350: inst = 32'hcc06b50;
      35351: inst = 32'h20800008;
      35352: inst = 32'h10c00000;
      35353: inst = 32'hcc06b50;
      35354: inst = 32'h20800009;
      35355: inst = 32'h10c00000;
      35356: inst = 32'hcc06b50;
      35357: inst = 32'h2080000a;
      35358: inst = 32'h10c00000;
      35359: inst = 32'hcc06b50;
      35360: inst = 32'h2080000b;
      35361: inst = 32'h10c00000;
      35362: inst = 32'hcc06b50;
      35363: inst = 32'h2080000c;
      35364: inst = 32'h10c00000;
      35365: inst = 32'hcc06b50;
      35366: inst = 32'h2080000d;
      35367: inst = 32'h10c00000;
      35368: inst = 32'hcc06b50;
      35369: inst = 32'h2080000e;
      35370: inst = 32'h10c00000;
      35371: inst = 32'hcc06b50;
      35372: inst = 32'h2080000f;
      35373: inst = 32'h10c00000;
      35374: inst = 32'hcc06b50;
      35375: inst = 32'h20800010;
      35376: inst = 32'h10c00000;
      35377: inst = 32'hcc06b50;
      35378: inst = 32'h20800011;
      35379: inst = 32'h10c00000;
      35380: inst = 32'hcc06b50;
      35381: inst = 32'h58a00000;
      35382: inst = 32'h20800000;
      35383: inst = 32'h10c00000;
      35384: inst = 32'hcc06b50;
      35385: inst = 32'h20800001;
      35386: inst = 32'h10c00000;
      35387: inst = 32'hcc06b50;
      35388: inst = 32'h20800002;
      35389: inst = 32'h10c00000;
      35390: inst = 32'hcc06b50;
      35391: inst = 32'h20800003;
      35392: inst = 32'h10c00000;
      35393: inst = 32'hcc06b50;
      35394: inst = 32'h20800004;
      35395: inst = 32'h10c00000;
      35396: inst = 32'hcc06b50;
      35397: inst = 32'h20800005;
      35398: inst = 32'h10c00000;
      35399: inst = 32'hcc06b50;
      35400: inst = 32'h20800006;
      35401: inst = 32'h10c00000;
      35402: inst = 32'hcc06b50;
      35403: inst = 32'h20800007;
      35404: inst = 32'h10c00000;
      35405: inst = 32'hcc06b50;
      35406: inst = 32'h20800008;
      35407: inst = 32'h10c00000;
      35408: inst = 32'hcc06b50;
      35409: inst = 32'h20800009;
      35410: inst = 32'h10c00000;
      35411: inst = 32'hcc06b50;
      35412: inst = 32'h2080000a;
      35413: inst = 32'h10c00000;
      35414: inst = 32'hcc06b50;
      35415: inst = 32'h2080000b;
      35416: inst = 32'h10c00000;
      35417: inst = 32'hcc06b50;
      35418: inst = 32'h2080000c;
      35419: inst = 32'h10c00000;
      35420: inst = 32'hcc06b50;
      35421: inst = 32'h2080000d;
      35422: inst = 32'h10c00000;
      35423: inst = 32'hcc06b50;
      35424: inst = 32'h2080000e;
      35425: inst = 32'h10c00000;
      35426: inst = 32'hcc06b50;
      35427: inst = 32'h2080000f;
      35428: inst = 32'h10c00000;
      35429: inst = 32'hcc06b50;
      35430: inst = 32'h20800010;
      35431: inst = 32'h10c00000;
      35432: inst = 32'hcc06b50;
      35433: inst = 32'h20800011;
      35434: inst = 32'h10c00000;
      35435: inst = 32'hcc06b50;
      35436: inst = 32'h58a00000;
      35437: inst = 32'h20800000;
      35438: inst = 32'h10c00000;
      35439: inst = 32'hcc06b50;
      35440: inst = 32'h20800001;
      35441: inst = 32'h10c00000;
      35442: inst = 32'hcc06b50;
      35443: inst = 32'h20800002;
      35444: inst = 32'h10c00000;
      35445: inst = 32'hcc06b50;
      35446: inst = 32'h20800003;
      35447: inst = 32'h10c00000;
      35448: inst = 32'hcc06b50;
      35449: inst = 32'h20800004;
      35450: inst = 32'h10c00000;
      35451: inst = 32'hcc06b50;
      35452: inst = 32'h20800005;
      35453: inst = 32'h10c00000;
      35454: inst = 32'hcc06b50;
      35455: inst = 32'h20800006;
      35456: inst = 32'h10c00000;
      35457: inst = 32'hcc06b50;
      35458: inst = 32'h20800007;
      35459: inst = 32'h10c00000;
      35460: inst = 32'hcc06b50;
      35461: inst = 32'h20800008;
      35462: inst = 32'h10c00000;
      35463: inst = 32'hcc06b50;
      35464: inst = 32'h20800009;
      35465: inst = 32'h10c00000;
      35466: inst = 32'hcc06b50;
      35467: inst = 32'h2080000a;
      35468: inst = 32'h10c00000;
      35469: inst = 32'hcc06b50;
      35470: inst = 32'h2080000b;
      35471: inst = 32'h10c00000;
      35472: inst = 32'hcc06b50;
      35473: inst = 32'h2080000c;
      35474: inst = 32'h10c00000;
      35475: inst = 32'hcc06b50;
      35476: inst = 32'h2080000d;
      35477: inst = 32'h10c00000;
      35478: inst = 32'hcc06b50;
      35479: inst = 32'h2080000e;
      35480: inst = 32'h10c00000;
      35481: inst = 32'hcc06b50;
      35482: inst = 32'h2080000f;
      35483: inst = 32'h10c00000;
      35484: inst = 32'hcc06b50;
      35485: inst = 32'h20800010;
      35486: inst = 32'h10c00000;
      35487: inst = 32'hcc06b50;
      35488: inst = 32'h20800011;
      35489: inst = 32'h10c00000;
      35490: inst = 32'hcc06b50;
      35491: inst = 32'h58a00000;
      35492: inst = 32'h20800000;
      35493: inst = 32'h10c00000;
      35494: inst = 32'hcc06b50;
      35495: inst = 32'h20800001;
      35496: inst = 32'h10c00000;
      35497: inst = 32'hcc06b50;
      35498: inst = 32'h20800002;
      35499: inst = 32'h10c00000;
      35500: inst = 32'hcc06b50;
      35501: inst = 32'h20800003;
      35502: inst = 32'h10c00000;
      35503: inst = 32'hcc06b50;
      35504: inst = 32'h20800004;
      35505: inst = 32'h10c00000;
      35506: inst = 32'hcc06b50;
      35507: inst = 32'h20800005;
      35508: inst = 32'h10c00000;
      35509: inst = 32'hcc06b50;
      35510: inst = 32'h20800006;
      35511: inst = 32'h10c00000;
      35512: inst = 32'hcc06b50;
      35513: inst = 32'h20800007;
      35514: inst = 32'h10c00000;
      35515: inst = 32'hcc06b50;
      35516: inst = 32'h20800008;
      35517: inst = 32'h10c00000;
      35518: inst = 32'hcc06b50;
      35519: inst = 32'h20800009;
      35520: inst = 32'h10c00000;
      35521: inst = 32'hcc06b50;
      35522: inst = 32'h2080000a;
      35523: inst = 32'h10c00000;
      35524: inst = 32'hcc06b50;
      35525: inst = 32'h2080000b;
      35526: inst = 32'h10c00000;
      35527: inst = 32'hcc06b50;
      35528: inst = 32'h2080000c;
      35529: inst = 32'h10c00000;
      35530: inst = 32'hcc06b50;
      35531: inst = 32'h2080000d;
      35532: inst = 32'h10c00000;
      35533: inst = 32'hcc06b50;
      35534: inst = 32'h2080000e;
      35535: inst = 32'h10c00000;
      35536: inst = 32'hcc06b50;
      35537: inst = 32'h2080000f;
      35538: inst = 32'h10c00000;
      35539: inst = 32'hcc06b50;
      35540: inst = 32'h20800010;
      35541: inst = 32'h10c00000;
      35542: inst = 32'hcc06b50;
      35543: inst = 32'h20800011;
      35544: inst = 32'h10c00000;
      35545: inst = 32'hcc06b50;
      35546: inst = 32'h58a00000;
      35547: inst = 32'h20800000;
      35548: inst = 32'h10c00000;
      35549: inst = 32'hcc06b50;
      35550: inst = 32'h20800001;
      35551: inst = 32'h10c00000;
      35552: inst = 32'hcc06b50;
      35553: inst = 32'h20800002;
      35554: inst = 32'h10c00000;
      35555: inst = 32'hcc06b50;
      35556: inst = 32'h20800003;
      35557: inst = 32'h10c00000;
      35558: inst = 32'hcc06b50;
      35559: inst = 32'h20800004;
      35560: inst = 32'h10c00000;
      35561: inst = 32'hcc06b50;
      35562: inst = 32'h20800005;
      35563: inst = 32'h10c00000;
      35564: inst = 32'hcc06b50;
      35565: inst = 32'h20800006;
      35566: inst = 32'h10c00000;
      35567: inst = 32'hcc06b50;
      35568: inst = 32'h20800007;
      35569: inst = 32'h10c00000;
      35570: inst = 32'hcc06b50;
      35571: inst = 32'h20800008;
      35572: inst = 32'h10c00000;
      35573: inst = 32'hcc06b50;
      35574: inst = 32'h20800009;
      35575: inst = 32'h10c00000;
      35576: inst = 32'hcc06b50;
      35577: inst = 32'h2080000a;
      35578: inst = 32'h10c00000;
      35579: inst = 32'hcc0eeb6;
      35580: inst = 32'h2080000b;
      35581: inst = 32'h10c00000;
      35582: inst = 32'hcc0eeb6;
      35583: inst = 32'h2080000c;
      35584: inst = 32'h10c00000;
      35585: inst = 32'hcc0eeb6;
      35586: inst = 32'h2080000d;
      35587: inst = 32'h10c00000;
      35588: inst = 32'hcc06b50;
      35589: inst = 32'h2080000e;
      35590: inst = 32'h10c00000;
      35591: inst = 32'hcc06b50;
      35592: inst = 32'h2080000f;
      35593: inst = 32'h10c00000;
      35594: inst = 32'hcc06b50;
      35595: inst = 32'h20800010;
      35596: inst = 32'h10c00000;
      35597: inst = 32'hcc06b50;
      35598: inst = 32'h20800011;
      35599: inst = 32'h10c00000;
      35600: inst = 32'hcc06b50;
      35601: inst = 32'h58a00000;
      35602: inst = 32'h20800000;
      35603: inst = 32'h10c00000;
      35604: inst = 32'hcc06b50;
      35605: inst = 32'h20800001;
      35606: inst = 32'h10c00000;
      35607: inst = 32'hcc06b50;
      35608: inst = 32'h20800002;
      35609: inst = 32'h10c00000;
      35610: inst = 32'hcc06b50;
      35611: inst = 32'h20800003;
      35612: inst = 32'h10c00000;
      35613: inst = 32'hcc06b50;
      35614: inst = 32'h20800004;
      35615: inst = 32'h10c00000;
      35616: inst = 32'hcc06b50;
      35617: inst = 32'h20800005;
      35618: inst = 32'h10c00000;
      35619: inst = 32'hcc06b50;
      35620: inst = 32'h20800006;
      35621: inst = 32'h10c00000;
      35622: inst = 32'hcc06b50;
      35623: inst = 32'h20800007;
      35624: inst = 32'h10c00000;
      35625: inst = 32'hcc06b50;
      35626: inst = 32'h20800008;
      35627: inst = 32'h10c00000;
      35628: inst = 32'hcc06b50;
      35629: inst = 32'h20800009;
      35630: inst = 32'h10c00000;
      35631: inst = 32'hcc06b50;
      35632: inst = 32'h2080000a;
      35633: inst = 32'h10c00000;
      35634: inst = 32'hcc0eeb6;
      35635: inst = 32'h2080000b;
      35636: inst = 32'h10c00000;
      35637: inst = 32'hcc0eeb6;
      35638: inst = 32'h2080000c;
      35639: inst = 32'h10c00000;
      35640: inst = 32'hcc0eeb6;
      35641: inst = 32'h2080000d;
      35642: inst = 32'h10c00000;
      35643: inst = 32'hcc06b50;
      35644: inst = 32'h2080000e;
      35645: inst = 32'h10c00000;
      35646: inst = 32'hcc06b50;
      35647: inst = 32'h2080000f;
      35648: inst = 32'h10c00000;
      35649: inst = 32'hcc06b50;
      35650: inst = 32'h20800010;
      35651: inst = 32'h10c00000;
      35652: inst = 32'hcc06b50;
      35653: inst = 32'h20800011;
      35654: inst = 32'h10c00000;
      35655: inst = 32'hcc06b50;
      35656: inst = 32'h58a00000;
      35657: inst = 32'h20800000;
      35658: inst = 32'h10c00000;
      35659: inst = 32'hcc06b50;
      35660: inst = 32'h20800001;
      35661: inst = 32'h10c00000;
      35662: inst = 32'hcc06b50;
      35663: inst = 32'h20800002;
      35664: inst = 32'h10c00000;
      35665: inst = 32'hcc06b50;
      35666: inst = 32'h20800003;
      35667: inst = 32'h10c00000;
      35668: inst = 32'hcc06b50;
      35669: inst = 32'h20800004;
      35670: inst = 32'h10c00000;
      35671: inst = 32'hcc06b50;
      35672: inst = 32'h20800005;
      35673: inst = 32'h10c00000;
      35674: inst = 32'hcc0eeb6;
      35675: inst = 32'h20800006;
      35676: inst = 32'h10c00000;
      35677: inst = 32'hcc0eeb6;
      35678: inst = 32'h20800007;
      35679: inst = 32'h10c00000;
      35680: inst = 32'hcc0eeb6;
      35681: inst = 32'h20800008;
      35682: inst = 32'h10c00000;
      35683: inst = 32'hcc06b50;
      35684: inst = 32'h20800009;
      35685: inst = 32'h10c00000;
      35686: inst = 32'hcc06b50;
      35687: inst = 32'h2080000a;
      35688: inst = 32'h10c00000;
      35689: inst = 32'hcc0eeb6;
      35690: inst = 32'h2080000b;
      35691: inst = 32'h10c00000;
      35692: inst = 32'hcc0eeb6;
      35693: inst = 32'h2080000c;
      35694: inst = 32'h10c00000;
      35695: inst = 32'hcc0eeb6;
      35696: inst = 32'h2080000d;
      35697: inst = 32'h10c00000;
      35698: inst = 32'hcc06b50;
      35699: inst = 32'h2080000e;
      35700: inst = 32'h10c00000;
      35701: inst = 32'hcc06b50;
      35702: inst = 32'h2080000f;
      35703: inst = 32'h10c00000;
      35704: inst = 32'hcc06b50;
      35705: inst = 32'h20800010;
      35706: inst = 32'h10c00000;
      35707: inst = 32'hcc06b50;
      35708: inst = 32'h20800011;
      35709: inst = 32'h10c00000;
      35710: inst = 32'hcc06b50;
      35711: inst = 32'h58a00000;
      35712: inst = 32'h20800000;
      35713: inst = 32'h10c00000;
      35714: inst = 32'hcc06b50;
      35715: inst = 32'h20800001;
      35716: inst = 32'h10c00000;
      35717: inst = 32'hcc06b50;
      35718: inst = 32'h20800002;
      35719: inst = 32'h10c00000;
      35720: inst = 32'hcc06b50;
      35721: inst = 32'h20800003;
      35722: inst = 32'h10c00000;
      35723: inst = 32'hcc06b50;
      35724: inst = 32'h20800004;
      35725: inst = 32'h10c00000;
      35726: inst = 32'hcc06b50;
      35727: inst = 32'h20800005;
      35728: inst = 32'h10c00000;
      35729: inst = 32'hcc0eeb6;
      35730: inst = 32'h20800006;
      35731: inst = 32'h10c00000;
      35732: inst = 32'hcc0eeb6;
      35733: inst = 32'h20800007;
      35734: inst = 32'h10c00000;
      35735: inst = 32'hcc0eeb6;
      35736: inst = 32'h20800008;
      35737: inst = 32'h10c00000;
      35738: inst = 32'hcc06b50;
      35739: inst = 32'h20800009;
      35740: inst = 32'h10c00000;
      35741: inst = 32'hcc06b50;
      35742: inst = 32'h2080000a;
      35743: inst = 32'h10c00000;
      35744: inst = 32'hcc0eeb6;
      35745: inst = 32'h2080000b;
      35746: inst = 32'h10c00000;
      35747: inst = 32'hcc0eeb6;
      35748: inst = 32'h2080000c;
      35749: inst = 32'h10c00000;
      35750: inst = 32'hcc06b50;
      35751: inst = 32'h2080000d;
      35752: inst = 32'h10c00000;
      35753: inst = 32'hcc06b50;
      35754: inst = 32'h2080000e;
      35755: inst = 32'h10c00000;
      35756: inst = 32'hcc06b50;
      35757: inst = 32'h2080000f;
      35758: inst = 32'h10c00000;
      35759: inst = 32'hcc06b50;
      35760: inst = 32'h20800010;
      35761: inst = 32'h10c00000;
      35762: inst = 32'hcc06b50;
      35763: inst = 32'h20800011;
      35764: inst = 32'h10c00000;
      35765: inst = 32'hcc06b50;
      35766: inst = 32'h58a00000;
      35767: inst = 32'h20800000;
      35768: inst = 32'h10c00000;
      35769: inst = 32'hcc06b50;
      35770: inst = 32'h20800001;
      35771: inst = 32'h10c00000;
      35772: inst = 32'hcc06b50;
      35773: inst = 32'h20800002;
      35774: inst = 32'h10c00000;
      35775: inst = 32'hcc06b50;
      35776: inst = 32'h20800003;
      35777: inst = 32'h10c00000;
      35778: inst = 32'hcc06b50;
      35779: inst = 32'h20800004;
      35780: inst = 32'h10c00000;
      35781: inst = 32'hcc06b50;
      35782: inst = 32'h20800005;
      35783: inst = 32'h10c00000;
      35784: inst = 32'hcc0eeb6;
      35785: inst = 32'h20800006;
      35786: inst = 32'h10c00000;
      35787: inst = 32'hcc0eeb6;
      35788: inst = 32'h20800007;
      35789: inst = 32'h10c00000;
      35790: inst = 32'hcc0eeb6;
      35791: inst = 32'h20800008;
      35792: inst = 32'h10c00000;
      35793: inst = 32'hcc0eeb6;
      35794: inst = 32'h20800009;
      35795: inst = 32'h10c00000;
      35796: inst = 32'hcc06b50;
      35797: inst = 32'h2080000a;
      35798: inst = 32'h10c00000;
      35799: inst = 32'hcc0eeb6;
      35800: inst = 32'h2080000b;
      35801: inst = 32'h10c00000;
      35802: inst = 32'hcc0eeb6;
      35803: inst = 32'h2080000c;
      35804: inst = 32'h10c00000;
      35805: inst = 32'hcc06b50;
      35806: inst = 32'h2080000d;
      35807: inst = 32'h10c00000;
      35808: inst = 32'hcc06b50;
      35809: inst = 32'h2080000e;
      35810: inst = 32'h10c00000;
      35811: inst = 32'hcc06b50;
      35812: inst = 32'h2080000f;
      35813: inst = 32'h10c00000;
      35814: inst = 32'hcc06b50;
      35815: inst = 32'h20800010;
      35816: inst = 32'h10c00000;
      35817: inst = 32'hcc06b50;
      35818: inst = 32'h20800011;
      35819: inst = 32'h10c00000;
      35820: inst = 32'hcc06b50;
      35821: inst = 32'h58a00000;
      35822: inst = 32'h20800000;
      35823: inst = 32'h10c00000;
      35824: inst = 32'hcc06b50;
      35825: inst = 32'h20800001;
      35826: inst = 32'h10c00000;
      35827: inst = 32'hcc06b50;
      35828: inst = 32'h20800002;
      35829: inst = 32'h10c00000;
      35830: inst = 32'hcc06b50;
      35831: inst = 32'h20800003;
      35832: inst = 32'h10c00000;
      35833: inst = 32'hcc06b50;
      35834: inst = 32'h20800004;
      35835: inst = 32'h10c00000;
      35836: inst = 32'hcc06b50;
      35837: inst = 32'h20800005;
      35838: inst = 32'h10c00000;
      35839: inst = 32'hcc0eeb6;
      35840: inst = 32'h20800006;
      35841: inst = 32'h10c00000;
      35842: inst = 32'hcc0eeb6;
      35843: inst = 32'h20800007;
      35844: inst = 32'h10c00000;
      35845: inst = 32'hcc06b50;
      35846: inst = 32'h20800008;
      35847: inst = 32'h10c00000;
      35848: inst = 32'hcc0eeb6;
      35849: inst = 32'h20800009;
      35850: inst = 32'h10c00000;
      35851: inst = 32'hcc06b50;
      35852: inst = 32'h2080000a;
      35853: inst = 32'h10c00000;
      35854: inst = 32'hcc0eeb6;
      35855: inst = 32'h2080000b;
      35856: inst = 32'h10c00000;
      35857: inst = 32'hcc0eeb6;
      35858: inst = 32'h2080000c;
      35859: inst = 32'h10c00000;
      35860: inst = 32'hcc06b50;
      35861: inst = 32'h2080000d;
      35862: inst = 32'h10c00000;
      35863: inst = 32'hcc06b50;
      35864: inst = 32'h2080000e;
      35865: inst = 32'h10c00000;
      35866: inst = 32'hcc06b50;
      35867: inst = 32'h2080000f;
      35868: inst = 32'h10c00000;
      35869: inst = 32'hcc06b50;
      35870: inst = 32'h20800010;
      35871: inst = 32'h10c00000;
      35872: inst = 32'hcc06b50;
      35873: inst = 32'h20800011;
      35874: inst = 32'h10c00000;
      35875: inst = 32'hcc06b50;
      35876: inst = 32'h58a00000;
      35877: inst = 32'h20800000;
      35878: inst = 32'h10c00000;
      35879: inst = 32'hcc06b50;
      35880: inst = 32'h20800001;
      35881: inst = 32'h10c00000;
      35882: inst = 32'hcc06b50;
      35883: inst = 32'h20800002;
      35884: inst = 32'h10c00000;
      35885: inst = 32'hcc06b50;
      35886: inst = 32'h20800003;
      35887: inst = 32'h10c00000;
      35888: inst = 32'hcc06b50;
      35889: inst = 32'h20800004;
      35890: inst = 32'h10c00000;
      35891: inst = 32'hcc06b50;
      35892: inst = 32'h20800005;
      35893: inst = 32'h10c00000;
      35894: inst = 32'hcc06b50;
      35895: inst = 32'h20800006;
      35896: inst = 32'h10c00000;
      35897: inst = 32'hcc0eeb6;
      35898: inst = 32'h20800007;
      35899: inst = 32'h10c00000;
      35900: inst = 32'hcc06b50;
      35901: inst = 32'h20800008;
      35902: inst = 32'h10c00000;
      35903: inst = 32'hcc0eeb6;
      35904: inst = 32'h20800009;
      35905: inst = 32'h10c00000;
      35906: inst = 32'hcc0eeb6;
      35907: inst = 32'h2080000a;
      35908: inst = 32'h10c00000;
      35909: inst = 32'hcc0eeb6;
      35910: inst = 32'h2080000b;
      35911: inst = 32'h10c00000;
      35912: inst = 32'hcc0eeb6;
      35913: inst = 32'h2080000c;
      35914: inst = 32'h10c00000;
      35915: inst = 32'hcc0eeb6;
      35916: inst = 32'h2080000d;
      35917: inst = 32'h10c00000;
      35918: inst = 32'hcc06b50;
      35919: inst = 32'h2080000e;
      35920: inst = 32'h10c00000;
      35921: inst = 32'hcc06b50;
      35922: inst = 32'h2080000f;
      35923: inst = 32'h10c00000;
      35924: inst = 32'hcc06b50;
      35925: inst = 32'h20800010;
      35926: inst = 32'h10c00000;
      35927: inst = 32'hcc06b50;
      35928: inst = 32'h20800011;
      35929: inst = 32'h10c00000;
      35930: inst = 32'hcc06b50;
      35931: inst = 32'h58a00000;
      35932: inst = 32'h20800000;
      35933: inst = 32'h10c00000;
      35934: inst = 32'hcc06b50;
      35935: inst = 32'h20800001;
      35936: inst = 32'h10c00000;
      35937: inst = 32'hcc06b50;
      35938: inst = 32'h20800002;
      35939: inst = 32'h10c00000;
      35940: inst = 32'hcc06b50;
      35941: inst = 32'h20800003;
      35942: inst = 32'h10c00000;
      35943: inst = 32'hcc06b50;
      35944: inst = 32'h20800004;
      35945: inst = 32'h10c00000;
      35946: inst = 32'hcc06b50;
      35947: inst = 32'h20800005;
      35948: inst = 32'h10c00000;
      35949: inst = 32'hcc06b50;
      35950: inst = 32'h20800006;
      35951: inst = 32'h10c00000;
      35952: inst = 32'hcc0eeb6;
      35953: inst = 32'h20800007;
      35954: inst = 32'h10c00000;
      35955: inst = 32'hcc06b50;
      35956: inst = 32'h20800008;
      35957: inst = 32'h10c00000;
      35958: inst = 32'hcc0eeb6;
      35959: inst = 32'h20800009;
      35960: inst = 32'h10c00000;
      35961: inst = 32'hcc0eeb6;
      35962: inst = 32'h2080000a;
      35963: inst = 32'h10c00000;
      35964: inst = 32'hcc06b50;
      35965: inst = 32'h2080000b;
      35966: inst = 32'h10c00000;
      35967: inst = 32'hcc0eeb6;
      35968: inst = 32'h2080000c;
      35969: inst = 32'h10c00000;
      35970: inst = 32'hcc0eeb6;
      35971: inst = 32'h2080000d;
      35972: inst = 32'h10c00000;
      35973: inst = 32'hcc06b50;
      35974: inst = 32'h2080000e;
      35975: inst = 32'h10c00000;
      35976: inst = 32'hcc06b50;
      35977: inst = 32'h2080000f;
      35978: inst = 32'h10c00000;
      35979: inst = 32'hcc06b50;
      35980: inst = 32'h20800010;
      35981: inst = 32'h10c00000;
      35982: inst = 32'hcc06b50;
      35983: inst = 32'h20800011;
      35984: inst = 32'h10c00000;
      35985: inst = 32'hcc06b50;
      35986: inst = 32'h58a00000;
      35987: inst = 32'h20800000;
      35988: inst = 32'h10c00000;
      35989: inst = 32'hcc06b50;
      35990: inst = 32'h20800001;
      35991: inst = 32'h10c00000;
      35992: inst = 32'hcc06b50;
      35993: inst = 32'h20800002;
      35994: inst = 32'h10c00000;
      35995: inst = 32'hcc06b50;
      35996: inst = 32'h20800003;
      35997: inst = 32'h10c00000;
      35998: inst = 32'hcc06b50;
      35999: inst = 32'h20800004;
      36000: inst = 32'h10c00000;
      36001: inst = 32'hcc06b50;
      36002: inst = 32'h20800005;
      36003: inst = 32'h10c00000;
      36004: inst = 32'hcc06b50;
      36005: inst = 32'h20800006;
      36006: inst = 32'h10c00000;
      36007: inst = 32'hcc0eeb6;
      36008: inst = 32'h20800007;
      36009: inst = 32'h10c00000;
      36010: inst = 32'hcc06b50;
      36011: inst = 32'h20800008;
      36012: inst = 32'h10c00000;
      36013: inst = 32'hcc0eeb6;
      36014: inst = 32'h20800009;
      36015: inst = 32'h10c00000;
      36016: inst = 32'hcc0eeb6;
      36017: inst = 32'h2080000a;
      36018: inst = 32'h10c00000;
      36019: inst = 32'hcc06b50;
      36020: inst = 32'h2080000b;
      36021: inst = 32'h10c00000;
      36022: inst = 32'hcc0eeb6;
      36023: inst = 32'h2080000c;
      36024: inst = 32'h10c00000;
      36025: inst = 32'hcc0eeb6;
      36026: inst = 32'h2080000d;
      36027: inst = 32'h10c00000;
      36028: inst = 32'hcc06b50;
      36029: inst = 32'h2080000e;
      36030: inst = 32'h10c00000;
      36031: inst = 32'hcc06b50;
      36032: inst = 32'h2080000f;
      36033: inst = 32'h10c00000;
      36034: inst = 32'hcc06b50;
      36035: inst = 32'h20800010;
      36036: inst = 32'h10c00000;
      36037: inst = 32'hcc06b50;
      36038: inst = 32'h20800011;
      36039: inst = 32'h10c00000;
      36040: inst = 32'hcc06b50;
      36041: inst = 32'h58a00000;
      36042: inst = 32'h20800000;
      36043: inst = 32'h10c00000;
      36044: inst = 32'hcc06b50;
      36045: inst = 32'h20800001;
      36046: inst = 32'h10c00000;
      36047: inst = 32'hcc06b50;
      36048: inst = 32'h20800002;
      36049: inst = 32'h10c00000;
      36050: inst = 32'hcc06b50;
      36051: inst = 32'h20800003;
      36052: inst = 32'h10c00000;
      36053: inst = 32'hcc06b50;
      36054: inst = 32'h20800004;
      36055: inst = 32'h10c00000;
      36056: inst = 32'hcc06b50;
      36057: inst = 32'h20800005;
      36058: inst = 32'h10c00000;
      36059: inst = 32'hcc06b50;
      36060: inst = 32'h20800006;
      36061: inst = 32'h10c00000;
      36062: inst = 32'hcc0eeb6;
      36063: inst = 32'h20800007;
      36064: inst = 32'h10c00000;
      36065: inst = 32'hcc06b50;
      36066: inst = 32'h20800008;
      36067: inst = 32'h10c00000;
      36068: inst = 32'hcc0eeb6;
      36069: inst = 32'h20800009;
      36070: inst = 32'h10c00000;
      36071: inst = 32'hcc0eeb6;
      36072: inst = 32'h2080000a;
      36073: inst = 32'h10c00000;
      36074: inst = 32'hcc06b50;
      36075: inst = 32'h2080000b;
      36076: inst = 32'h10c00000;
      36077: inst = 32'hcc0eeb6;
      36078: inst = 32'h2080000c;
      36079: inst = 32'h10c00000;
      36080: inst = 32'hcc06b50;
      36081: inst = 32'h2080000d;
      36082: inst = 32'h10c00000;
      36083: inst = 32'hcc06b50;
      36084: inst = 32'h2080000e;
      36085: inst = 32'h10c00000;
      36086: inst = 32'hcc06b50;
      36087: inst = 32'h2080000f;
      36088: inst = 32'h10c00000;
      36089: inst = 32'hcc06b50;
      36090: inst = 32'h20800010;
      36091: inst = 32'h10c00000;
      36092: inst = 32'hcc06b50;
      36093: inst = 32'h20800011;
      36094: inst = 32'h10c00000;
      36095: inst = 32'hcc06b50;
      36096: inst = 32'h58a00000;
      36097: inst = 32'h20800000;
      36098: inst = 32'h10c00000;
      36099: inst = 32'hcc06b50;
      36100: inst = 32'h20800001;
      36101: inst = 32'h10c00000;
      36102: inst = 32'hcc06b50;
      36103: inst = 32'h20800002;
      36104: inst = 32'h10c00000;
      36105: inst = 32'hcc06b50;
      36106: inst = 32'h20800003;
      36107: inst = 32'h10c00000;
      36108: inst = 32'hcc06b50;
      36109: inst = 32'h20800004;
      36110: inst = 32'h10c00000;
      36111: inst = 32'hcc06b50;
      36112: inst = 32'h20800005;
      36113: inst = 32'h10c00000;
      36114: inst = 32'hcc06b50;
      36115: inst = 32'h20800006;
      36116: inst = 32'h10c00000;
      36117: inst = 32'hcc0eeb6;
      36118: inst = 32'h20800007;
      36119: inst = 32'h10c00000;
      36120: inst = 32'hcc06b50;
      36121: inst = 32'h20800008;
      36122: inst = 32'h10c00000;
      36123: inst = 32'hcc0eeb6;
      36124: inst = 32'h20800009;
      36125: inst = 32'h10c00000;
      36126: inst = 32'hcc0eeb6;
      36127: inst = 32'h2080000a;
      36128: inst = 32'h10c00000;
      36129: inst = 32'hcc06b50;
      36130: inst = 32'h2080000b;
      36131: inst = 32'h10c00000;
      36132: inst = 32'hcc0eeb6;
      36133: inst = 32'h2080000c;
      36134: inst = 32'h10c00000;
      36135: inst = 32'hcc06b50;
      36136: inst = 32'h2080000d;
      36137: inst = 32'h10c00000;
      36138: inst = 32'hcc06b50;
      36139: inst = 32'h2080000e;
      36140: inst = 32'h10c00000;
      36141: inst = 32'hcc06b50;
      36142: inst = 32'h2080000f;
      36143: inst = 32'h10c00000;
      36144: inst = 32'hcc06b50;
      36145: inst = 32'h20800010;
      36146: inst = 32'h10c00000;
      36147: inst = 32'hcc06b50;
      36148: inst = 32'h20800011;
      36149: inst = 32'h10c00000;
      36150: inst = 32'hcc06b50;
      36151: inst = 32'h58a00000;
      36152: inst = 32'h20800000;
      36153: inst = 32'h10c00000;
      36154: inst = 32'hcc06b50;
      36155: inst = 32'h20800001;
      36156: inst = 32'h10c00000;
      36157: inst = 32'hcc06b50;
      36158: inst = 32'h20800002;
      36159: inst = 32'h10c00000;
      36160: inst = 32'hcc06b50;
      36161: inst = 32'h20800003;
      36162: inst = 32'h10c00000;
      36163: inst = 32'hcc06b50;
      36164: inst = 32'h20800004;
      36165: inst = 32'h10c00000;
      36166: inst = 32'hcc06b50;
      36167: inst = 32'h20800005;
      36168: inst = 32'h10c00000;
      36169: inst = 32'hcc0eeb6;
      36170: inst = 32'h20800006;
      36171: inst = 32'h10c00000;
      36172: inst = 32'hcc0eeb6;
      36173: inst = 32'h20800007;
      36174: inst = 32'h10c00000;
      36175: inst = 32'hcc06b50;
      36176: inst = 32'h20800008;
      36177: inst = 32'h10c00000;
      36178: inst = 32'hcc0eeb6;
      36179: inst = 32'h20800009;
      36180: inst = 32'h10c00000;
      36181: inst = 32'hcc0eeb6;
      36182: inst = 32'h2080000a;
      36183: inst = 32'h10c00000;
      36184: inst = 32'hcc0eeb6;
      36185: inst = 32'h2080000b;
      36186: inst = 32'h10c00000;
      36187: inst = 32'hcc0eeb6;
      36188: inst = 32'h2080000c;
      36189: inst = 32'h10c00000;
      36190: inst = 32'hcc06b50;
      36191: inst = 32'h2080000d;
      36192: inst = 32'h10c00000;
      36193: inst = 32'hcc06b50;
      36194: inst = 32'h2080000e;
      36195: inst = 32'h10c00000;
      36196: inst = 32'hcc06b50;
      36197: inst = 32'h2080000f;
      36198: inst = 32'h10c00000;
      36199: inst = 32'hcc06b50;
      36200: inst = 32'h20800010;
      36201: inst = 32'h10c00000;
      36202: inst = 32'hcc06b50;
      36203: inst = 32'h20800011;
      36204: inst = 32'h10c00000;
      36205: inst = 32'hcc06b50;
      36206: inst = 32'h58a00000;
      36207: inst = 32'h20800000;
      36208: inst = 32'h10c00000;
      36209: inst = 32'hcc06b50;
      36210: inst = 32'h20800001;
      36211: inst = 32'h10c00000;
      36212: inst = 32'hcc06b50;
      36213: inst = 32'h20800002;
      36214: inst = 32'h10c00000;
      36215: inst = 32'hcc06b50;
      36216: inst = 32'h20800003;
      36217: inst = 32'h10c00000;
      36218: inst = 32'hcc06b50;
      36219: inst = 32'h20800004;
      36220: inst = 32'h10c00000;
      36221: inst = 32'hcc06b50;
      36222: inst = 32'h20800005;
      36223: inst = 32'h10c00000;
      36224: inst = 32'hcc0eeb6;
      36225: inst = 32'h20800006;
      36226: inst = 32'h10c00000;
      36227: inst = 32'hcc0eeb6;
      36228: inst = 32'h20800007;
      36229: inst = 32'h10c00000;
      36230: inst = 32'hcc0eeb6;
      36231: inst = 32'h20800008;
      36232: inst = 32'h10c00000;
      36233: inst = 32'hcc0eeb6;
      36234: inst = 32'h20800009;
      36235: inst = 32'h10c00000;
      36236: inst = 32'hcc0eeb6;
      36237: inst = 32'h2080000a;
      36238: inst = 32'h10c00000;
      36239: inst = 32'hcc0eeb6;
      36240: inst = 32'h2080000b;
      36241: inst = 32'h10c00000;
      36242: inst = 32'hcc06b50;
      36243: inst = 32'h2080000c;
      36244: inst = 32'h10c00000;
      36245: inst = 32'hcc06b50;
      36246: inst = 32'h2080000d;
      36247: inst = 32'h10c00000;
      36248: inst = 32'hcc06b50;
      36249: inst = 32'h2080000e;
      36250: inst = 32'h10c00000;
      36251: inst = 32'hcc06b50;
      36252: inst = 32'h2080000f;
      36253: inst = 32'h10c00000;
      36254: inst = 32'hcc06b50;
      36255: inst = 32'h20800010;
      36256: inst = 32'h10c00000;
      36257: inst = 32'hcc06b50;
      36258: inst = 32'h20800011;
      36259: inst = 32'h10c00000;
      36260: inst = 32'hcc06b50;
      36261: inst = 32'h58a00000;
      36262: inst = 32'h20800000;
      36263: inst = 32'h10c00000;
      36264: inst = 32'hcc06b50;
      36265: inst = 32'h20800001;
      36266: inst = 32'h10c00000;
      36267: inst = 32'hcc06b50;
      36268: inst = 32'h20800002;
      36269: inst = 32'h10c00000;
      36270: inst = 32'hcc06b50;
      36271: inst = 32'h20800003;
      36272: inst = 32'h10c00000;
      36273: inst = 32'hcc06b50;
      36274: inst = 32'h20800004;
      36275: inst = 32'h10c00000;
      36276: inst = 32'hcc06b50;
      36277: inst = 32'h20800005;
      36278: inst = 32'h10c00000;
      36279: inst = 32'hcc0eeb6;
      36280: inst = 32'h20800006;
      36281: inst = 32'h10c00000;
      36282: inst = 32'hcc0eeb6;
      36283: inst = 32'h20800007;
      36284: inst = 32'h10c00000;
      36285: inst = 32'hcc06b50;
      36286: inst = 32'h20800008;
      36287: inst = 32'h10c00000;
      36288: inst = 32'hcc0eeb6;
      36289: inst = 32'h20800009;
      36290: inst = 32'h10c00000;
      36291: inst = 32'hcc0eeb6;
      36292: inst = 32'h2080000a;
      36293: inst = 32'h10c00000;
      36294: inst = 32'hcc0eeb6;
      36295: inst = 32'h2080000b;
      36296: inst = 32'h10c00000;
      36297: inst = 32'hcc06b50;
      36298: inst = 32'h2080000c;
      36299: inst = 32'h10c00000;
      36300: inst = 32'hcc06b50;
      36301: inst = 32'h2080000d;
      36302: inst = 32'h10c00000;
      36303: inst = 32'hcc06b50;
      36304: inst = 32'h2080000e;
      36305: inst = 32'h10c00000;
      36306: inst = 32'hcc06b50;
      36307: inst = 32'h2080000f;
      36308: inst = 32'h10c00000;
      36309: inst = 32'hcc06b50;
      36310: inst = 32'h20800010;
      36311: inst = 32'h10c00000;
      36312: inst = 32'hcc06b50;
      36313: inst = 32'h20800011;
      36314: inst = 32'h10c00000;
      36315: inst = 32'hcc06b50;
      36316: inst = 32'h58a00000;
      36317: inst = 32'h20800000;
      36318: inst = 32'h10c00000;
      36319: inst = 32'hcc06b50;
      36320: inst = 32'h20800001;
      36321: inst = 32'h10c00000;
      36322: inst = 32'hcc06b50;
      36323: inst = 32'h20800002;
      36324: inst = 32'h10c00000;
      36325: inst = 32'hcc06b50;
      36326: inst = 32'h20800003;
      36327: inst = 32'h10c00000;
      36328: inst = 32'hcc06b50;
      36329: inst = 32'h20800004;
      36330: inst = 32'h10c00000;
      36331: inst = 32'hcc06b50;
      36332: inst = 32'h20800005;
      36333: inst = 32'h10c00000;
      36334: inst = 32'hcc0eeb6;
      36335: inst = 32'h20800006;
      36336: inst = 32'h10c00000;
      36337: inst = 32'hcc0eeb6;
      36338: inst = 32'h20800007;
      36339: inst = 32'h10c00000;
      36340: inst = 32'hcc06b50;
      36341: inst = 32'h20800008;
      36342: inst = 32'h10c00000;
      36343: inst = 32'hcc0eeb6;
      36344: inst = 32'h20800009;
      36345: inst = 32'h10c00000;
      36346: inst = 32'hcc0eeb6;
      36347: inst = 32'h2080000a;
      36348: inst = 32'h10c00000;
      36349: inst = 32'hcc0eeb6;
      36350: inst = 32'h2080000b;
      36351: inst = 32'h10c00000;
      36352: inst = 32'hcc06b50;
      36353: inst = 32'h2080000c;
      36354: inst = 32'h10c00000;
      36355: inst = 32'hcc06b50;
      36356: inst = 32'h2080000d;
      36357: inst = 32'h10c00000;
      36358: inst = 32'hcc06b50;
      36359: inst = 32'h2080000e;
      36360: inst = 32'h10c00000;
      36361: inst = 32'hcc06b50;
      36362: inst = 32'h2080000f;
      36363: inst = 32'h10c00000;
      36364: inst = 32'hcc06b50;
      36365: inst = 32'h20800010;
      36366: inst = 32'h10c00000;
      36367: inst = 32'hcc06b50;
      36368: inst = 32'h20800011;
      36369: inst = 32'h10c00000;
      36370: inst = 32'hcc06b50;
      36371: inst = 32'h58a00000;
      36372: inst = 32'h20800000;
      36373: inst = 32'h10c00000;
      36374: inst = 32'hcc06b50;
      36375: inst = 32'h20800001;
      36376: inst = 32'h10c00000;
      36377: inst = 32'hcc06b50;
      36378: inst = 32'h20800002;
      36379: inst = 32'h10c00000;
      36380: inst = 32'hcc06b50;
      36381: inst = 32'h20800003;
      36382: inst = 32'h10c00000;
      36383: inst = 32'hcc06b50;
      36384: inst = 32'h20800004;
      36385: inst = 32'h10c00000;
      36386: inst = 32'hcc06b50;
      36387: inst = 32'h20800005;
      36388: inst = 32'h10c00000;
      36389: inst = 32'hcc0eeb6;
      36390: inst = 32'h20800006;
      36391: inst = 32'h10c00000;
      36392: inst = 32'hcc0eeb6;
      36393: inst = 32'h20800007;
      36394: inst = 32'h10c00000;
      36395: inst = 32'hcc06b50;
      36396: inst = 32'h20800008;
      36397: inst = 32'h10c00000;
      36398: inst = 32'hcc0eeb6;
      36399: inst = 32'h20800009;
      36400: inst = 32'h10c00000;
      36401: inst = 32'hcc0eeb6;
      36402: inst = 32'h2080000a;
      36403: inst = 32'h10c00000;
      36404: inst = 32'hcc0eeb6;
      36405: inst = 32'h2080000b;
      36406: inst = 32'h10c00000;
      36407: inst = 32'hcc06b50;
      36408: inst = 32'h2080000c;
      36409: inst = 32'h10c00000;
      36410: inst = 32'hcc06b50;
      36411: inst = 32'h2080000d;
      36412: inst = 32'h10c00000;
      36413: inst = 32'hcc06b50;
      36414: inst = 32'h2080000e;
      36415: inst = 32'h10c00000;
      36416: inst = 32'hcc06b50;
      36417: inst = 32'h2080000f;
      36418: inst = 32'h10c00000;
      36419: inst = 32'hcc06b50;
      36420: inst = 32'h20800010;
      36421: inst = 32'h10c00000;
      36422: inst = 32'hcc06b50;
      36423: inst = 32'h20800011;
      36424: inst = 32'h10c00000;
      36425: inst = 32'hcc06b50;
      36426: inst = 32'h58a00000;
      36427: inst = 32'h20800000;
      36428: inst = 32'h10c00000;
      36429: inst = 32'hcc06b50;
      36430: inst = 32'h20800001;
      36431: inst = 32'h10c00000;
      36432: inst = 32'hcc06b50;
      36433: inst = 32'h20800002;
      36434: inst = 32'h10c00000;
      36435: inst = 32'hcc06b50;
      36436: inst = 32'h20800003;
      36437: inst = 32'h10c00000;
      36438: inst = 32'hcc06b50;
      36439: inst = 32'h20800004;
      36440: inst = 32'h10c00000;
      36441: inst = 32'hcc06b50;
      36442: inst = 32'h20800005;
      36443: inst = 32'h10c00000;
      36444: inst = 32'hcc0eeb6;
      36445: inst = 32'h20800006;
      36446: inst = 32'h10c00000;
      36447: inst = 32'hcc0eeb6;
      36448: inst = 32'h20800007;
      36449: inst = 32'h10c00000;
      36450: inst = 32'hcc06b50;
      36451: inst = 32'h20800008;
      36452: inst = 32'h10c00000;
      36453: inst = 32'hcc0eeb6;
      36454: inst = 32'h20800009;
      36455: inst = 32'h10c00000;
      36456: inst = 32'hcc0eeb6;
      36457: inst = 32'h2080000a;
      36458: inst = 32'h10c00000;
      36459: inst = 32'hcc0eeb6;
      36460: inst = 32'h2080000b;
      36461: inst = 32'h10c00000;
      36462: inst = 32'hcc06b50;
      36463: inst = 32'h2080000c;
      36464: inst = 32'h10c00000;
      36465: inst = 32'hcc06b50;
      36466: inst = 32'h2080000d;
      36467: inst = 32'h10c00000;
      36468: inst = 32'hcc06b50;
      36469: inst = 32'h2080000e;
      36470: inst = 32'h10c00000;
      36471: inst = 32'hcc06b50;
      36472: inst = 32'h2080000f;
      36473: inst = 32'h10c00000;
      36474: inst = 32'hcc06b50;
      36475: inst = 32'h20800010;
      36476: inst = 32'h10c00000;
      36477: inst = 32'hcc06b50;
      36478: inst = 32'h20800011;
      36479: inst = 32'h10c00000;
      36480: inst = 32'hcc06b50;
      36481: inst = 32'h58a00000;
      36482: inst = 32'h20800000;
      36483: inst = 32'h10c00000;
      36484: inst = 32'hcc06b50;
      36485: inst = 32'h20800001;
      36486: inst = 32'h10c00000;
      36487: inst = 32'hcc06b50;
      36488: inst = 32'h20800002;
      36489: inst = 32'h10c00000;
      36490: inst = 32'hcc06b50;
      36491: inst = 32'h20800003;
      36492: inst = 32'h10c00000;
      36493: inst = 32'hcc06b50;
      36494: inst = 32'h20800004;
      36495: inst = 32'h10c00000;
      36496: inst = 32'hcc06b50;
      36497: inst = 32'h20800005;
      36498: inst = 32'h10c00000;
      36499: inst = 32'hcc06b50;
      36500: inst = 32'h20800006;
      36501: inst = 32'h10c00000;
      36502: inst = 32'hcc06b50;
      36503: inst = 32'h20800007;
      36504: inst = 32'h10c00000;
      36505: inst = 32'hcc06b50;
      36506: inst = 32'h20800008;
      36507: inst = 32'h10c00000;
      36508: inst = 32'hcc06b50;
      36509: inst = 32'h20800009;
      36510: inst = 32'h10c00000;
      36511: inst = 32'hcc06b50;
      36512: inst = 32'h2080000a;
      36513: inst = 32'h10c00000;
      36514: inst = 32'hcc06b50;
      36515: inst = 32'h2080000b;
      36516: inst = 32'h10c00000;
      36517: inst = 32'hcc06b50;
      36518: inst = 32'h2080000c;
      36519: inst = 32'h10c00000;
      36520: inst = 32'hcc06b50;
      36521: inst = 32'h2080000d;
      36522: inst = 32'h10c00000;
      36523: inst = 32'hcc06b50;
      36524: inst = 32'h2080000e;
      36525: inst = 32'h10c00000;
      36526: inst = 32'hcc06b50;
      36527: inst = 32'h2080000f;
      36528: inst = 32'h10c00000;
      36529: inst = 32'hcc06b50;
      36530: inst = 32'h20800010;
      36531: inst = 32'h10c00000;
      36532: inst = 32'hcc06b50;
      36533: inst = 32'h20800011;
      36534: inst = 32'h10c00000;
      36535: inst = 32'hcc06b50;
      36536: inst = 32'h58a00000;
      36537: inst = 32'h20800000;
      36538: inst = 32'h10c00000;
      36539: inst = 32'hcc06b50;
      36540: inst = 32'h20800001;
      36541: inst = 32'h10c00000;
      36542: inst = 32'hcc06b50;
      36543: inst = 32'h20800002;
      36544: inst = 32'h10c00000;
      36545: inst = 32'hcc06b50;
      36546: inst = 32'h20800003;
      36547: inst = 32'h10c00000;
      36548: inst = 32'hcc06b50;
      36549: inst = 32'h20800004;
      36550: inst = 32'h10c00000;
      36551: inst = 32'hcc06b50;
      36552: inst = 32'h20800005;
      36553: inst = 32'h10c00000;
      36554: inst = 32'hcc06b50;
      36555: inst = 32'h20800006;
      36556: inst = 32'h10c00000;
      36557: inst = 32'hcc06b50;
      36558: inst = 32'h20800007;
      36559: inst = 32'h10c00000;
      36560: inst = 32'hcc06b50;
      36561: inst = 32'h20800008;
      36562: inst = 32'h10c00000;
      36563: inst = 32'hcc06b50;
      36564: inst = 32'h20800009;
      36565: inst = 32'h10c00000;
      36566: inst = 32'hcc06b50;
      36567: inst = 32'h2080000a;
      36568: inst = 32'h10c00000;
      36569: inst = 32'hcc06b50;
      36570: inst = 32'h2080000b;
      36571: inst = 32'h10c00000;
      36572: inst = 32'hcc06b50;
      36573: inst = 32'h2080000c;
      36574: inst = 32'h10c00000;
      36575: inst = 32'hcc06b50;
      36576: inst = 32'h2080000d;
      36577: inst = 32'h10c00000;
      36578: inst = 32'hcc06b50;
      36579: inst = 32'h2080000e;
      36580: inst = 32'h10c00000;
      36581: inst = 32'hcc06b50;
      36582: inst = 32'h2080000f;
      36583: inst = 32'h10c00000;
      36584: inst = 32'hcc06b50;
      36585: inst = 32'h20800010;
      36586: inst = 32'h10c00000;
      36587: inst = 32'hcc06b50;
      36588: inst = 32'h20800011;
      36589: inst = 32'h10c00000;
      36590: inst = 32'hcc06b50;
      36591: inst = 32'h58a00000;
      36592: inst = 32'h20800000;
      36593: inst = 32'h10c00000;
      36594: inst = 32'hcc06b50;
      36595: inst = 32'h20800001;
      36596: inst = 32'h10c00000;
      36597: inst = 32'hcc06b50;
      36598: inst = 32'h20800002;
      36599: inst = 32'h10c00000;
      36600: inst = 32'hcc06b50;
      36601: inst = 32'h20800003;
      36602: inst = 32'h10c00000;
      36603: inst = 32'hcc06b50;
      36604: inst = 32'h20800004;
      36605: inst = 32'h10c00000;
      36606: inst = 32'hcc06b50;
      36607: inst = 32'h20800005;
      36608: inst = 32'h10c00000;
      36609: inst = 32'hcc06b50;
      36610: inst = 32'h20800006;
      36611: inst = 32'h10c00000;
      36612: inst = 32'hcc06b50;
      36613: inst = 32'h20800007;
      36614: inst = 32'h10c00000;
      36615: inst = 32'hcc06b50;
      36616: inst = 32'h20800008;
      36617: inst = 32'h10c00000;
      36618: inst = 32'hcc06b50;
      36619: inst = 32'h20800009;
      36620: inst = 32'h10c00000;
      36621: inst = 32'hcc06b50;
      36622: inst = 32'h2080000a;
      36623: inst = 32'h10c00000;
      36624: inst = 32'hcc06b50;
      36625: inst = 32'h2080000b;
      36626: inst = 32'h10c00000;
      36627: inst = 32'hcc06b50;
      36628: inst = 32'h2080000c;
      36629: inst = 32'h10c00000;
      36630: inst = 32'hcc06b50;
      36631: inst = 32'h2080000d;
      36632: inst = 32'h10c00000;
      36633: inst = 32'hcc06b50;
      36634: inst = 32'h2080000e;
      36635: inst = 32'h10c00000;
      36636: inst = 32'hcc06b50;
      36637: inst = 32'h2080000f;
      36638: inst = 32'h10c00000;
      36639: inst = 32'hcc06b50;
      36640: inst = 32'h20800010;
      36641: inst = 32'h10c00000;
      36642: inst = 32'hcc06b50;
      36643: inst = 32'h20800011;
      36644: inst = 32'h10c00000;
      36645: inst = 32'hcc06b50;
      36646: inst = 32'h58a00000;
      36647: inst = 32'h20800000;
      36648: inst = 32'h10c00000;
      36649: inst = 32'hcc06b50;
      36650: inst = 32'h20800001;
      36651: inst = 32'h10c00000;
      36652: inst = 32'hcc06b50;
      36653: inst = 32'h20800002;
      36654: inst = 32'h10c00000;
      36655: inst = 32'hcc06b50;
      36656: inst = 32'h20800003;
      36657: inst = 32'h10c00000;
      36658: inst = 32'hcc06b50;
      36659: inst = 32'h20800004;
      36660: inst = 32'h10c00000;
      36661: inst = 32'hcc06b50;
      36662: inst = 32'h20800005;
      36663: inst = 32'h10c00000;
      36664: inst = 32'hcc06b50;
      36665: inst = 32'h20800006;
      36666: inst = 32'h10c00000;
      36667: inst = 32'hcc06b50;
      36668: inst = 32'h20800007;
      36669: inst = 32'h10c00000;
      36670: inst = 32'hcc06b50;
      36671: inst = 32'h20800008;
      36672: inst = 32'h10c00000;
      36673: inst = 32'hcc06b50;
      36674: inst = 32'h20800009;
      36675: inst = 32'h10c00000;
      36676: inst = 32'hcc06b50;
      36677: inst = 32'h2080000a;
      36678: inst = 32'h10c00000;
      36679: inst = 32'hcc06b50;
      36680: inst = 32'h2080000b;
      36681: inst = 32'h10c00000;
      36682: inst = 32'hcc06b50;
      36683: inst = 32'h2080000c;
      36684: inst = 32'h10c00000;
      36685: inst = 32'hcc06b50;
      36686: inst = 32'h2080000d;
      36687: inst = 32'h10c00000;
      36688: inst = 32'hcc06b50;
      36689: inst = 32'h2080000e;
      36690: inst = 32'h10c00000;
      36691: inst = 32'hcc06b50;
      36692: inst = 32'h2080000f;
      36693: inst = 32'h10c00000;
      36694: inst = 32'hcc06b50;
      36695: inst = 32'h20800010;
      36696: inst = 32'h10c00000;
      36697: inst = 32'hcc06b50;
      36698: inst = 32'h20800011;
      36699: inst = 32'h10c00000;
      36700: inst = 32'hcc06b50;
      36701: inst = 32'h58a00000;
      36702: inst = 32'h11800000;
      36703: inst = 32'hd800000;
      36704: inst = 32'h11a00000;
      36705: inst = 32'hda00000;
      36706: inst = 32'h25ad5800;
      36707: inst = 32'h15ca6800;
      36708: inst = 32'h21c00001;
      36709: inst = 32'h59200000;
      36710: inst = 32'h298c0001;
      36711: inst = 32'h13e00000;
      36712: inst = 32'hfe08f62;
      36713: inst = 32'h5be00000;
      36714: inst = 32'h11800000;
      36715: inst = 32'hd800000;
      36716: inst = 32'h258c5800;
      36717: inst = 32'h15aa6000;
      36718: inst = 32'h13e0ffff;
      36719: inst = 32'h13e00000;
      36720: inst = 32'hfe08f75;
      36721: inst = 32'h5be00000;
      36722: inst = 32'h13e00000;
      36723: inst = 32'hfe08f6c;
      36724: inst = 32'h5be00000;
      36725: inst = 32'h2d8c5800;
      36726: inst = 32'h2d8a6000;
      36727: inst = 32'h59200000;
    endcase
  end
endmodule
