`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: lirc572
// Engineer: lirc572
// 
// Create Date: 
// Design Name: NECPU
// Module Name: InstMem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module instMem (
    input  [31:0]  address,
    output reg [31:0] inst
  );
  always @ (address) begin
    inst = 32'd0;
    case (address)
      0: inst = 32'h10000000;
      1: inst = 32'hc000005;
      2: inst = 32'h13e00000;
      3: inst = 32'hfe00098;
      4: inst = 32'h5be00000;
      5: inst = 32'h1020007f;
      6: inst = 32'hc202815;
      7: inst = 32'h30210001;
      8: inst = 32'h13e00000;
      9: inst = 32'hfe00007;
      10: inst = 32'h1c200000;
      11: inst = 32'h5be00000;
      12: inst = 32'h10000000;
      13: inst = 32'hc000011;
      14: inst = 32'h13e00000;
      15: inst = 32'hfe048f0;
      16: inst = 32'h5be00000;
      17: inst = 32'h1020007f;
      18: inst = 32'hc202815;
      19: inst = 32'h30210001;
      20: inst = 32'h13e00000;
      21: inst = 32'hfe00013;
      22: inst = 32'h1c200000;
      23: inst = 32'h5be00000;
      24: inst = 32'h10000000;
      25: inst = 32'hc000000;
      26: inst = 32'h10200000;
      27: inst = 32'hc20001f;
      28: inst = 32'h13e00000;
      29: inst = 32'hfe06109;
      30: inst = 32'h5be00000;
      31: inst = 32'h10000000;
      32: inst = 32'hc000024;
      33: inst = 32'h13a00000;
      34: inst = 32'hfa00000;
      35: inst = 32'h13600000;
      36: inst = 32'hf600000;
      37: inst = 32'h13800000;
      38: inst = 32'hf800000;
      39: inst = 32'h12800000;
      40: inst = 32'he800045;
      41: inst = 32'h12a00000;
      42: inst = 32'hea0002b;
      43: inst = 32'h1734d800;
      44: inst = 32'h1755e000;
      45: inst = 32'h13e00000;
      46: inst = 32'hfe00038;
      47: inst = 32'h1f200001;
      48: inst = 32'h5be00000;
      49: inst = 32'h13e00000;
      50: inst = 32'hfe00038;
      51: inst = 32'h1f400001;
      52: inst = 32'h5be00000;
      53: inst = 32'h13e00000;
      54: inst = 32'hfe00095;
      55: inst = 32'h5be00000;
      56: inst = 32'h10208000;
      57: inst = 32'hc200001;
      58: inst = 32'h4210000;
      59: inst = 32'h10400000;
      60: inst = 32'hc40001b;
      61: inst = 32'h34211000;
      62: inst = 32'h38211000;
      63: inst = 32'h13e00000;
      64: inst = 32'hfe00052;
      65: inst = 32'h20200010;
      66: inst = 32'h5be00000;
      67: inst = 32'h13e00000;
      68: inst = 32'hfe0005c;
      69: inst = 32'h20200008;
      70: inst = 32'h5be00000;
      71: inst = 32'h13e00000;
      72: inst = 32'hfe00066;
      73: inst = 32'h20200004;
      74: inst = 32'h5be00000;
      75: inst = 32'h13e00000;
      76: inst = 32'hfe00070;
      77: inst = 32'h20200002;
      78: inst = 32'h5be00000;
      79: inst = 32'h13e00000;
      80: inst = 32'hfe0007a;
      81: inst = 32'h5be00000;
      82: inst = 32'h339c0001;
      83: inst = 32'h13a00000;
      84: inst = 32'hfa00000;
      85: inst = 32'hca00001;
      86: inst = 32'h10c08000;
      87: inst = 32'hcc00000;
      88: inst = 32'h8a60000;
      89: inst = 32'h13e00000;
      90: inst = 32'hfe0007e;
      91: inst = 32'h5be00000;
      92: inst = 32'h2b7b0001;
      93: inst = 32'h13a00000;
      94: inst = 32'hfa00003;
      95: inst = 32'hca00002;
      96: inst = 32'h10c08000;
      97: inst = 32'hcc00000;
      98: inst = 32'h8a60000;
      99: inst = 32'h13e00000;
      100: inst = 32'hfe0007e;
      101: inst = 32'h5be00000;
      102: inst = 32'h337b0001;
      103: inst = 32'h13a00000;
      104: inst = 32'hfa00001;
      105: inst = 32'hca00004;
      106: inst = 32'h10c08000;
      107: inst = 32'hcc00000;
      108: inst = 32'h8a60000;
      109: inst = 32'h13e00000;
      110: inst = 32'hfe0007e;
      111: inst = 32'h5be00000;
      112: inst = 32'h2b9c0001;
      113: inst = 32'h13a00000;
      114: inst = 32'hfa00005;
      115: inst = 32'hca00008;
      116: inst = 32'h10c08000;
      117: inst = 32'hcc00000;
      118: inst = 32'h8a60000;
      119: inst = 32'h13e00000;
      120: inst = 32'hfe0007e;
      121: inst = 32'h5be00000;
      122: inst = 32'hca00010;
      123: inst = 32'h10c08000;
      124: inst = 32'hcc00000;
      125: inst = 32'h8a60000;
      126: inst = 32'h10000000;
      127: inst = 32'hc000083;
      128: inst = 32'h13e00000;
      129: inst = 32'hfe06113;
      130: inst = 32'h5be00000;
      131: inst = 32'h283d0000;
      132: inst = 32'h285b0000;
      133: inst = 32'h287c0000;
      134: inst = 32'h10000000;
      135: inst = 32'hc00008b;
      136: inst = 32'h13e00000;
      137: inst = 32'hfe05141;
      138: inst = 32'h5be00000;
      139: inst = 32'h10200002;
      140: inst = 32'hc208b0a;
      141: inst = 32'h30210001;
      142: inst = 32'h13e00000;
      143: inst = 32'hfe0008d;
      144: inst = 32'h1c200000;
      145: inst = 32'h5be00000;
      146: inst = 32'h13e00000;
      147: inst = 32'hfe00027;
      148: inst = 32'h5be00000;
      149: inst = 32'h13e00000;
      150: inst = 32'hfe0aa05;
      151: inst = 32'h5be00000;
      152: inst = 32'hc20eeb6;
      153: inst = 32'h10408000;
      154: inst = 32'hc403fe0;
      155: inst = 32'h8220000;
      156: inst = 32'h10408000;
      157: inst = 32'hc403fe1;
      158: inst = 32'h8220000;
      159: inst = 32'h10408000;
      160: inst = 32'hc403fe2;
      161: inst = 32'h8220000;
      162: inst = 32'h10408000;
      163: inst = 32'hc403fe3;
      164: inst = 32'h8220000;
      165: inst = 32'h10408000;
      166: inst = 32'hc403fe4;
      167: inst = 32'h8220000;
      168: inst = 32'h10408000;
      169: inst = 32'hc403fe5;
      170: inst = 32'h8220000;
      171: inst = 32'h10408000;
      172: inst = 32'hc403fe6;
      173: inst = 32'h8220000;
      174: inst = 32'h10408000;
      175: inst = 32'hc403fe7;
      176: inst = 32'h8220000;
      177: inst = 32'h10408000;
      178: inst = 32'hc403fe8;
      179: inst = 32'h8220000;
      180: inst = 32'h10408000;
      181: inst = 32'hc403fe9;
      182: inst = 32'h8220000;
      183: inst = 32'h10408000;
      184: inst = 32'hc403fea;
      185: inst = 32'h8220000;
      186: inst = 32'h10408000;
      187: inst = 32'hc403fec;
      188: inst = 32'h8220000;
      189: inst = 32'h10408000;
      190: inst = 32'hc403fed;
      191: inst = 32'h8220000;
      192: inst = 32'h10408000;
      193: inst = 32'hc403fee;
      194: inst = 32'h8220000;
      195: inst = 32'h10408000;
      196: inst = 32'hc403fef;
      197: inst = 32'h8220000;
      198: inst = 32'h10408000;
      199: inst = 32'hc403ff0;
      200: inst = 32'h8220000;
      201: inst = 32'h10408000;
      202: inst = 32'hc403ff1;
      203: inst = 32'h8220000;
      204: inst = 32'h10408000;
      205: inst = 32'hc403ff2;
      206: inst = 32'h8220000;
      207: inst = 32'h10408000;
      208: inst = 32'hc403ff3;
      209: inst = 32'h8220000;
      210: inst = 32'h10408000;
      211: inst = 32'hc403ff4;
      212: inst = 32'h8220000;
      213: inst = 32'h10408000;
      214: inst = 32'hc403ff5;
      215: inst = 32'h8220000;
      216: inst = 32'h10408000;
      217: inst = 32'hc403ff6;
      218: inst = 32'h8220000;
      219: inst = 32'h10408000;
      220: inst = 32'hc403ff7;
      221: inst = 32'h8220000;
      222: inst = 32'h10408000;
      223: inst = 32'hc403ff8;
      224: inst = 32'h8220000;
      225: inst = 32'h10408000;
      226: inst = 32'hc403ff9;
      227: inst = 32'h8220000;
      228: inst = 32'h10408000;
      229: inst = 32'hc403ffa;
      230: inst = 32'h8220000;
      231: inst = 32'h10408000;
      232: inst = 32'hc403ffb;
      233: inst = 32'h8220000;
      234: inst = 32'h10408000;
      235: inst = 32'hc403ffc;
      236: inst = 32'h8220000;
      237: inst = 32'h10408000;
      238: inst = 32'hc403ffd;
      239: inst = 32'h8220000;
      240: inst = 32'h10408000;
      241: inst = 32'hc403ffe;
      242: inst = 32'h8220000;
      243: inst = 32'h10408000;
      244: inst = 32'hc403fff;
      245: inst = 32'h8220000;
      246: inst = 32'h10408000;
      247: inst = 32'hc404000;
      248: inst = 32'h8220000;
      249: inst = 32'h10408000;
      250: inst = 32'hc404001;
      251: inst = 32'h8220000;
      252: inst = 32'h10408000;
      253: inst = 32'hc404002;
      254: inst = 32'h8220000;
      255: inst = 32'h10408000;
      256: inst = 32'hc404003;
      257: inst = 32'h8220000;
      258: inst = 32'h10408000;
      259: inst = 32'hc404004;
      260: inst = 32'h8220000;
      261: inst = 32'h10408000;
      262: inst = 32'hc404005;
      263: inst = 32'h8220000;
      264: inst = 32'h10408000;
      265: inst = 32'hc404006;
      266: inst = 32'h8220000;
      267: inst = 32'h10408000;
      268: inst = 32'hc404007;
      269: inst = 32'h8220000;
      270: inst = 32'h10408000;
      271: inst = 32'hc404008;
      272: inst = 32'h8220000;
      273: inst = 32'h10408000;
      274: inst = 32'hc404009;
      275: inst = 32'h8220000;
      276: inst = 32'h10408000;
      277: inst = 32'hc40400a;
      278: inst = 32'h8220000;
      279: inst = 32'h10408000;
      280: inst = 32'hc40400b;
      281: inst = 32'h8220000;
      282: inst = 32'h10408000;
      283: inst = 32'hc40400c;
      284: inst = 32'h8220000;
      285: inst = 32'h10408000;
      286: inst = 32'hc40400d;
      287: inst = 32'h8220000;
      288: inst = 32'h10408000;
      289: inst = 32'hc40400e;
      290: inst = 32'h8220000;
      291: inst = 32'h10408000;
      292: inst = 32'hc40400f;
      293: inst = 32'h8220000;
      294: inst = 32'h10408000;
      295: inst = 32'hc404010;
      296: inst = 32'h8220000;
      297: inst = 32'h10408000;
      298: inst = 32'hc404011;
      299: inst = 32'h8220000;
      300: inst = 32'h10408000;
      301: inst = 32'hc404012;
      302: inst = 32'h8220000;
      303: inst = 32'h10408000;
      304: inst = 32'hc404013;
      305: inst = 32'h8220000;
      306: inst = 32'h10408000;
      307: inst = 32'hc404014;
      308: inst = 32'h8220000;
      309: inst = 32'h10408000;
      310: inst = 32'hc404015;
      311: inst = 32'h8220000;
      312: inst = 32'h10408000;
      313: inst = 32'hc404016;
      314: inst = 32'h8220000;
      315: inst = 32'h10408000;
      316: inst = 32'hc404017;
      317: inst = 32'h8220000;
      318: inst = 32'h10408000;
      319: inst = 32'hc404018;
      320: inst = 32'h8220000;
      321: inst = 32'h10408000;
      322: inst = 32'hc404019;
      323: inst = 32'h8220000;
      324: inst = 32'h10408000;
      325: inst = 32'hc40401a;
      326: inst = 32'h8220000;
      327: inst = 32'h10408000;
      328: inst = 32'hc40401b;
      329: inst = 32'h8220000;
      330: inst = 32'h10408000;
      331: inst = 32'hc40401c;
      332: inst = 32'h8220000;
      333: inst = 32'h10408000;
      334: inst = 32'hc40401d;
      335: inst = 32'h8220000;
      336: inst = 32'h10408000;
      337: inst = 32'hc40401e;
      338: inst = 32'h8220000;
      339: inst = 32'h10408000;
      340: inst = 32'hc40401f;
      341: inst = 32'h8220000;
      342: inst = 32'h10408000;
      343: inst = 32'hc404020;
      344: inst = 32'h8220000;
      345: inst = 32'h10408000;
      346: inst = 32'hc404021;
      347: inst = 32'h8220000;
      348: inst = 32'h10408000;
      349: inst = 32'hc404022;
      350: inst = 32'h8220000;
      351: inst = 32'h10408000;
      352: inst = 32'hc404023;
      353: inst = 32'h8220000;
      354: inst = 32'h10408000;
      355: inst = 32'hc404024;
      356: inst = 32'h8220000;
      357: inst = 32'h10408000;
      358: inst = 32'hc404025;
      359: inst = 32'h8220000;
      360: inst = 32'h10408000;
      361: inst = 32'hc404026;
      362: inst = 32'h8220000;
      363: inst = 32'h10408000;
      364: inst = 32'hc404027;
      365: inst = 32'h8220000;
      366: inst = 32'h10408000;
      367: inst = 32'hc404028;
      368: inst = 32'h8220000;
      369: inst = 32'h10408000;
      370: inst = 32'hc404029;
      371: inst = 32'h8220000;
      372: inst = 32'h10408000;
      373: inst = 32'hc40402a;
      374: inst = 32'h8220000;
      375: inst = 32'h10408000;
      376: inst = 32'hc40402b;
      377: inst = 32'h8220000;
      378: inst = 32'h10408000;
      379: inst = 32'hc40402c;
      380: inst = 32'h8220000;
      381: inst = 32'h10408000;
      382: inst = 32'hc40402d;
      383: inst = 32'h8220000;
      384: inst = 32'h10408000;
      385: inst = 32'hc40402e;
      386: inst = 32'h8220000;
      387: inst = 32'h10408000;
      388: inst = 32'hc40402f;
      389: inst = 32'h8220000;
      390: inst = 32'h10408000;
      391: inst = 32'hc404030;
      392: inst = 32'h8220000;
      393: inst = 32'h10408000;
      394: inst = 32'hc404031;
      395: inst = 32'h8220000;
      396: inst = 32'h10408000;
      397: inst = 32'hc404032;
      398: inst = 32'h8220000;
      399: inst = 32'h10408000;
      400: inst = 32'hc404033;
      401: inst = 32'h8220000;
      402: inst = 32'h10408000;
      403: inst = 32'hc404034;
      404: inst = 32'h8220000;
      405: inst = 32'h10408000;
      406: inst = 32'hc404035;
      407: inst = 32'h8220000;
      408: inst = 32'h10408000;
      409: inst = 32'hc404036;
      410: inst = 32'h8220000;
      411: inst = 32'h10408000;
      412: inst = 32'hc404037;
      413: inst = 32'h8220000;
      414: inst = 32'h10408000;
      415: inst = 32'hc404038;
      416: inst = 32'h8220000;
      417: inst = 32'h10408000;
      418: inst = 32'hc404039;
      419: inst = 32'h8220000;
      420: inst = 32'h10408000;
      421: inst = 32'hc40403a;
      422: inst = 32'h8220000;
      423: inst = 32'h10408000;
      424: inst = 32'hc40403b;
      425: inst = 32'h8220000;
      426: inst = 32'h10408000;
      427: inst = 32'hc40403c;
      428: inst = 32'h8220000;
      429: inst = 32'h10408000;
      430: inst = 32'hc40403d;
      431: inst = 32'h8220000;
      432: inst = 32'h10408000;
      433: inst = 32'hc40403e;
      434: inst = 32'h8220000;
      435: inst = 32'h10408000;
      436: inst = 32'hc40403f;
      437: inst = 32'h8220000;
      438: inst = 32'h10408000;
      439: inst = 32'hc404040;
      440: inst = 32'h8220000;
      441: inst = 32'h10408000;
      442: inst = 32'hc404041;
      443: inst = 32'h8220000;
      444: inst = 32'h10408000;
      445: inst = 32'hc404042;
      446: inst = 32'h8220000;
      447: inst = 32'h10408000;
      448: inst = 32'hc404043;
      449: inst = 32'h8220000;
      450: inst = 32'h10408000;
      451: inst = 32'hc404044;
      452: inst = 32'h8220000;
      453: inst = 32'h10408000;
      454: inst = 32'hc404045;
      455: inst = 32'h8220000;
      456: inst = 32'h10408000;
      457: inst = 32'hc404046;
      458: inst = 32'h8220000;
      459: inst = 32'h10408000;
      460: inst = 32'hc404047;
      461: inst = 32'h8220000;
      462: inst = 32'h10408000;
      463: inst = 32'hc404048;
      464: inst = 32'h8220000;
      465: inst = 32'h10408000;
      466: inst = 32'hc404049;
      467: inst = 32'h8220000;
      468: inst = 32'h10408000;
      469: inst = 32'hc40404a;
      470: inst = 32'h8220000;
      471: inst = 32'h10408000;
      472: inst = 32'hc40404c;
      473: inst = 32'h8220000;
      474: inst = 32'h10408000;
      475: inst = 32'hc40404d;
      476: inst = 32'h8220000;
      477: inst = 32'h10408000;
      478: inst = 32'hc40404e;
      479: inst = 32'h8220000;
      480: inst = 32'h10408000;
      481: inst = 32'hc40404f;
      482: inst = 32'h8220000;
      483: inst = 32'h10408000;
      484: inst = 32'hc404050;
      485: inst = 32'h8220000;
      486: inst = 32'h10408000;
      487: inst = 32'hc404051;
      488: inst = 32'h8220000;
      489: inst = 32'h10408000;
      490: inst = 32'hc404052;
      491: inst = 32'h8220000;
      492: inst = 32'h10408000;
      493: inst = 32'hc404053;
      494: inst = 32'h8220000;
      495: inst = 32'h10408000;
      496: inst = 32'hc404054;
      497: inst = 32'h8220000;
      498: inst = 32'h10408000;
      499: inst = 32'hc404055;
      500: inst = 32'h8220000;
      501: inst = 32'h10408000;
      502: inst = 32'hc404056;
      503: inst = 32'h8220000;
      504: inst = 32'h10408000;
      505: inst = 32'hc404057;
      506: inst = 32'h8220000;
      507: inst = 32'h10408000;
      508: inst = 32'hc404058;
      509: inst = 32'h8220000;
      510: inst = 32'h10408000;
      511: inst = 32'hc404059;
      512: inst = 32'h8220000;
      513: inst = 32'h10408000;
      514: inst = 32'hc40405a;
      515: inst = 32'h8220000;
      516: inst = 32'h10408000;
      517: inst = 32'hc40405b;
      518: inst = 32'h8220000;
      519: inst = 32'h10408000;
      520: inst = 32'hc40405c;
      521: inst = 32'h8220000;
      522: inst = 32'h10408000;
      523: inst = 32'hc40405d;
      524: inst = 32'h8220000;
      525: inst = 32'h10408000;
      526: inst = 32'hc40405e;
      527: inst = 32'h8220000;
      528: inst = 32'h10408000;
      529: inst = 32'hc40405f;
      530: inst = 32'h8220000;
      531: inst = 32'h10408000;
      532: inst = 32'hc404060;
      533: inst = 32'h8220000;
      534: inst = 32'h10408000;
      535: inst = 32'hc404061;
      536: inst = 32'h8220000;
      537: inst = 32'h10408000;
      538: inst = 32'hc404062;
      539: inst = 32'h8220000;
      540: inst = 32'h10408000;
      541: inst = 32'hc404063;
      542: inst = 32'h8220000;
      543: inst = 32'h10408000;
      544: inst = 32'hc404064;
      545: inst = 32'h8220000;
      546: inst = 32'h10408000;
      547: inst = 32'hc404065;
      548: inst = 32'h8220000;
      549: inst = 32'h10408000;
      550: inst = 32'hc404066;
      551: inst = 32'h8220000;
      552: inst = 32'h10408000;
      553: inst = 32'hc404067;
      554: inst = 32'h8220000;
      555: inst = 32'h10408000;
      556: inst = 32'hc404068;
      557: inst = 32'h8220000;
      558: inst = 32'h10408000;
      559: inst = 32'hc404069;
      560: inst = 32'h8220000;
      561: inst = 32'h10408000;
      562: inst = 32'hc40406a;
      563: inst = 32'h8220000;
      564: inst = 32'h10408000;
      565: inst = 32'hc40406b;
      566: inst = 32'h8220000;
      567: inst = 32'h10408000;
      568: inst = 32'hc40406c;
      569: inst = 32'h8220000;
      570: inst = 32'h10408000;
      571: inst = 32'hc40406d;
      572: inst = 32'h8220000;
      573: inst = 32'h10408000;
      574: inst = 32'hc40406e;
      575: inst = 32'h8220000;
      576: inst = 32'h10408000;
      577: inst = 32'hc40406f;
      578: inst = 32'h8220000;
      579: inst = 32'h10408000;
      580: inst = 32'hc404070;
      581: inst = 32'h8220000;
      582: inst = 32'h10408000;
      583: inst = 32'hc404071;
      584: inst = 32'h8220000;
      585: inst = 32'h10408000;
      586: inst = 32'hc404072;
      587: inst = 32'h8220000;
      588: inst = 32'h10408000;
      589: inst = 32'hc404073;
      590: inst = 32'h8220000;
      591: inst = 32'h10408000;
      592: inst = 32'hc404074;
      593: inst = 32'h8220000;
      594: inst = 32'h10408000;
      595: inst = 32'hc404075;
      596: inst = 32'h8220000;
      597: inst = 32'h10408000;
      598: inst = 32'hc404076;
      599: inst = 32'h8220000;
      600: inst = 32'h10408000;
      601: inst = 32'hc404077;
      602: inst = 32'h8220000;
      603: inst = 32'h10408000;
      604: inst = 32'hc404078;
      605: inst = 32'h8220000;
      606: inst = 32'h10408000;
      607: inst = 32'hc404079;
      608: inst = 32'h8220000;
      609: inst = 32'h10408000;
      610: inst = 32'hc40407a;
      611: inst = 32'h8220000;
      612: inst = 32'h10408000;
      613: inst = 32'hc40407b;
      614: inst = 32'h8220000;
      615: inst = 32'h10408000;
      616: inst = 32'hc40407c;
      617: inst = 32'h8220000;
      618: inst = 32'h10408000;
      619: inst = 32'hc40407d;
      620: inst = 32'h8220000;
      621: inst = 32'h10408000;
      622: inst = 32'hc40407e;
      623: inst = 32'h8220000;
      624: inst = 32'h10408000;
      625: inst = 32'hc40407f;
      626: inst = 32'h8220000;
      627: inst = 32'h10408000;
      628: inst = 32'hc404080;
      629: inst = 32'h8220000;
      630: inst = 32'h10408000;
      631: inst = 32'hc404081;
      632: inst = 32'h8220000;
      633: inst = 32'h10408000;
      634: inst = 32'hc404082;
      635: inst = 32'h8220000;
      636: inst = 32'h10408000;
      637: inst = 32'hc404083;
      638: inst = 32'h8220000;
      639: inst = 32'h10408000;
      640: inst = 32'hc404084;
      641: inst = 32'h8220000;
      642: inst = 32'h10408000;
      643: inst = 32'hc404085;
      644: inst = 32'h8220000;
      645: inst = 32'h10408000;
      646: inst = 32'hc404086;
      647: inst = 32'h8220000;
      648: inst = 32'h10408000;
      649: inst = 32'hc404087;
      650: inst = 32'h8220000;
      651: inst = 32'h10408000;
      652: inst = 32'hc404088;
      653: inst = 32'h8220000;
      654: inst = 32'h10408000;
      655: inst = 32'hc404089;
      656: inst = 32'h8220000;
      657: inst = 32'h10408000;
      658: inst = 32'hc40408a;
      659: inst = 32'h8220000;
      660: inst = 32'h10408000;
      661: inst = 32'hc40408b;
      662: inst = 32'h8220000;
      663: inst = 32'h10408000;
      664: inst = 32'hc40408c;
      665: inst = 32'h8220000;
      666: inst = 32'h10408000;
      667: inst = 32'hc40408d;
      668: inst = 32'h8220000;
      669: inst = 32'h10408000;
      670: inst = 32'hc40408e;
      671: inst = 32'h8220000;
      672: inst = 32'h10408000;
      673: inst = 32'hc40408f;
      674: inst = 32'h8220000;
      675: inst = 32'h10408000;
      676: inst = 32'hc404090;
      677: inst = 32'h8220000;
      678: inst = 32'h10408000;
      679: inst = 32'hc404091;
      680: inst = 32'h8220000;
      681: inst = 32'h10408000;
      682: inst = 32'hc404092;
      683: inst = 32'h8220000;
      684: inst = 32'h10408000;
      685: inst = 32'hc404093;
      686: inst = 32'h8220000;
      687: inst = 32'h10408000;
      688: inst = 32'hc404094;
      689: inst = 32'h8220000;
      690: inst = 32'h10408000;
      691: inst = 32'hc404095;
      692: inst = 32'h8220000;
      693: inst = 32'h10408000;
      694: inst = 32'hc404096;
      695: inst = 32'h8220000;
      696: inst = 32'h10408000;
      697: inst = 32'hc404097;
      698: inst = 32'h8220000;
      699: inst = 32'h10408000;
      700: inst = 32'hc404098;
      701: inst = 32'h8220000;
      702: inst = 32'h10408000;
      703: inst = 32'hc404099;
      704: inst = 32'h8220000;
      705: inst = 32'h10408000;
      706: inst = 32'hc40409a;
      707: inst = 32'h8220000;
      708: inst = 32'h10408000;
      709: inst = 32'hc40409b;
      710: inst = 32'h8220000;
      711: inst = 32'h10408000;
      712: inst = 32'hc40409c;
      713: inst = 32'h8220000;
      714: inst = 32'h10408000;
      715: inst = 32'hc40409d;
      716: inst = 32'h8220000;
      717: inst = 32'h10408000;
      718: inst = 32'hc40409e;
      719: inst = 32'h8220000;
      720: inst = 32'h10408000;
      721: inst = 32'hc40409f;
      722: inst = 32'h8220000;
      723: inst = 32'h10408000;
      724: inst = 32'hc4040a0;
      725: inst = 32'h8220000;
      726: inst = 32'h10408000;
      727: inst = 32'hc4040a1;
      728: inst = 32'h8220000;
      729: inst = 32'h10408000;
      730: inst = 32'hc4040a2;
      731: inst = 32'h8220000;
      732: inst = 32'h10408000;
      733: inst = 32'hc4040a3;
      734: inst = 32'h8220000;
      735: inst = 32'h10408000;
      736: inst = 32'hc4040a4;
      737: inst = 32'h8220000;
      738: inst = 32'h10408000;
      739: inst = 32'hc4040a5;
      740: inst = 32'h8220000;
      741: inst = 32'h10408000;
      742: inst = 32'hc4040a6;
      743: inst = 32'h8220000;
      744: inst = 32'h10408000;
      745: inst = 32'hc4040a7;
      746: inst = 32'h8220000;
      747: inst = 32'h10408000;
      748: inst = 32'hc4040a8;
      749: inst = 32'h8220000;
      750: inst = 32'h10408000;
      751: inst = 32'hc4040a9;
      752: inst = 32'h8220000;
      753: inst = 32'h10408000;
      754: inst = 32'hc4040aa;
      755: inst = 32'h8220000;
      756: inst = 32'h10408000;
      757: inst = 32'hc4040ac;
      758: inst = 32'h8220000;
      759: inst = 32'h10408000;
      760: inst = 32'hc4040ad;
      761: inst = 32'h8220000;
      762: inst = 32'h10408000;
      763: inst = 32'hc4040ae;
      764: inst = 32'h8220000;
      765: inst = 32'h10408000;
      766: inst = 32'hc4040af;
      767: inst = 32'h8220000;
      768: inst = 32'h10408000;
      769: inst = 32'hc4040b0;
      770: inst = 32'h8220000;
      771: inst = 32'h10408000;
      772: inst = 32'hc4040b1;
      773: inst = 32'h8220000;
      774: inst = 32'h10408000;
      775: inst = 32'hc4040b2;
      776: inst = 32'h8220000;
      777: inst = 32'h10408000;
      778: inst = 32'hc4040b3;
      779: inst = 32'h8220000;
      780: inst = 32'h10408000;
      781: inst = 32'hc4040b4;
      782: inst = 32'h8220000;
      783: inst = 32'h10408000;
      784: inst = 32'hc4040b5;
      785: inst = 32'h8220000;
      786: inst = 32'h10408000;
      787: inst = 32'hc4040b6;
      788: inst = 32'h8220000;
      789: inst = 32'h10408000;
      790: inst = 32'hc4040b7;
      791: inst = 32'h8220000;
      792: inst = 32'h10408000;
      793: inst = 32'hc4040b8;
      794: inst = 32'h8220000;
      795: inst = 32'h10408000;
      796: inst = 32'hc4040b9;
      797: inst = 32'h8220000;
      798: inst = 32'h10408000;
      799: inst = 32'hc4040ba;
      800: inst = 32'h8220000;
      801: inst = 32'h10408000;
      802: inst = 32'hc4040bb;
      803: inst = 32'h8220000;
      804: inst = 32'h10408000;
      805: inst = 32'hc4040bc;
      806: inst = 32'h8220000;
      807: inst = 32'h10408000;
      808: inst = 32'hc4040bd;
      809: inst = 32'h8220000;
      810: inst = 32'h10408000;
      811: inst = 32'hc4040be;
      812: inst = 32'h8220000;
      813: inst = 32'h10408000;
      814: inst = 32'hc4040bf;
      815: inst = 32'h8220000;
      816: inst = 32'h10408000;
      817: inst = 32'hc4040c0;
      818: inst = 32'h8220000;
      819: inst = 32'h10408000;
      820: inst = 32'hc4040c1;
      821: inst = 32'h8220000;
      822: inst = 32'h10408000;
      823: inst = 32'hc4040c2;
      824: inst = 32'h8220000;
      825: inst = 32'h10408000;
      826: inst = 32'hc4040c3;
      827: inst = 32'h8220000;
      828: inst = 32'h10408000;
      829: inst = 32'hc4040c4;
      830: inst = 32'h8220000;
      831: inst = 32'h10408000;
      832: inst = 32'hc4040c5;
      833: inst = 32'h8220000;
      834: inst = 32'h10408000;
      835: inst = 32'hc4040c6;
      836: inst = 32'h8220000;
      837: inst = 32'h10408000;
      838: inst = 32'hc4040c7;
      839: inst = 32'h8220000;
      840: inst = 32'h10408000;
      841: inst = 32'hc4040c8;
      842: inst = 32'h8220000;
      843: inst = 32'h10408000;
      844: inst = 32'hc4040c9;
      845: inst = 32'h8220000;
      846: inst = 32'h10408000;
      847: inst = 32'hc4040ca;
      848: inst = 32'h8220000;
      849: inst = 32'h10408000;
      850: inst = 32'hc4040cb;
      851: inst = 32'h8220000;
      852: inst = 32'h10408000;
      853: inst = 32'hc4040cc;
      854: inst = 32'h8220000;
      855: inst = 32'h10408000;
      856: inst = 32'hc4040cd;
      857: inst = 32'h8220000;
      858: inst = 32'h10408000;
      859: inst = 32'hc4040ce;
      860: inst = 32'h8220000;
      861: inst = 32'h10408000;
      862: inst = 32'hc4040cf;
      863: inst = 32'h8220000;
      864: inst = 32'h10408000;
      865: inst = 32'hc4040d0;
      866: inst = 32'h8220000;
      867: inst = 32'h10408000;
      868: inst = 32'hc4040d1;
      869: inst = 32'h8220000;
      870: inst = 32'h10408000;
      871: inst = 32'hc4040d2;
      872: inst = 32'h8220000;
      873: inst = 32'h10408000;
      874: inst = 32'hc4040d3;
      875: inst = 32'h8220000;
      876: inst = 32'h10408000;
      877: inst = 32'hc4040d4;
      878: inst = 32'h8220000;
      879: inst = 32'h10408000;
      880: inst = 32'hc4040d5;
      881: inst = 32'h8220000;
      882: inst = 32'h10408000;
      883: inst = 32'hc4040d6;
      884: inst = 32'h8220000;
      885: inst = 32'h10408000;
      886: inst = 32'hc4040d7;
      887: inst = 32'h8220000;
      888: inst = 32'h10408000;
      889: inst = 32'hc4040d8;
      890: inst = 32'h8220000;
      891: inst = 32'h10408000;
      892: inst = 32'hc4040d9;
      893: inst = 32'h8220000;
      894: inst = 32'h10408000;
      895: inst = 32'hc4040da;
      896: inst = 32'h8220000;
      897: inst = 32'h10408000;
      898: inst = 32'hc4040db;
      899: inst = 32'h8220000;
      900: inst = 32'h10408000;
      901: inst = 32'hc4040dc;
      902: inst = 32'h8220000;
      903: inst = 32'h10408000;
      904: inst = 32'hc4040dd;
      905: inst = 32'h8220000;
      906: inst = 32'h10408000;
      907: inst = 32'hc4040de;
      908: inst = 32'h8220000;
      909: inst = 32'h10408000;
      910: inst = 32'hc4040df;
      911: inst = 32'h8220000;
      912: inst = 32'h10408000;
      913: inst = 32'hc4040e0;
      914: inst = 32'h8220000;
      915: inst = 32'h10408000;
      916: inst = 32'hc4040e1;
      917: inst = 32'h8220000;
      918: inst = 32'h10408000;
      919: inst = 32'hc4040e2;
      920: inst = 32'h8220000;
      921: inst = 32'h10408000;
      922: inst = 32'hc4040e3;
      923: inst = 32'h8220000;
      924: inst = 32'h10408000;
      925: inst = 32'hc4040e4;
      926: inst = 32'h8220000;
      927: inst = 32'h10408000;
      928: inst = 32'hc4040e5;
      929: inst = 32'h8220000;
      930: inst = 32'h10408000;
      931: inst = 32'hc4040e6;
      932: inst = 32'h8220000;
      933: inst = 32'h10408000;
      934: inst = 32'hc4040e7;
      935: inst = 32'h8220000;
      936: inst = 32'h10408000;
      937: inst = 32'hc4040e8;
      938: inst = 32'h8220000;
      939: inst = 32'h10408000;
      940: inst = 32'hc4040e9;
      941: inst = 32'h8220000;
      942: inst = 32'h10408000;
      943: inst = 32'hc4040ea;
      944: inst = 32'h8220000;
      945: inst = 32'h10408000;
      946: inst = 32'hc4040eb;
      947: inst = 32'h8220000;
      948: inst = 32'h10408000;
      949: inst = 32'hc4040ec;
      950: inst = 32'h8220000;
      951: inst = 32'h10408000;
      952: inst = 32'hc4040ed;
      953: inst = 32'h8220000;
      954: inst = 32'h10408000;
      955: inst = 32'hc4040ee;
      956: inst = 32'h8220000;
      957: inst = 32'h10408000;
      958: inst = 32'hc4040ef;
      959: inst = 32'h8220000;
      960: inst = 32'h10408000;
      961: inst = 32'hc4040f0;
      962: inst = 32'h8220000;
      963: inst = 32'h10408000;
      964: inst = 32'hc4040f1;
      965: inst = 32'h8220000;
      966: inst = 32'h10408000;
      967: inst = 32'hc4040f2;
      968: inst = 32'h8220000;
      969: inst = 32'h10408000;
      970: inst = 32'hc4040f3;
      971: inst = 32'h8220000;
      972: inst = 32'h10408000;
      973: inst = 32'hc4040f4;
      974: inst = 32'h8220000;
      975: inst = 32'h10408000;
      976: inst = 32'hc4040f5;
      977: inst = 32'h8220000;
      978: inst = 32'h10408000;
      979: inst = 32'hc4040f6;
      980: inst = 32'h8220000;
      981: inst = 32'h10408000;
      982: inst = 32'hc4040f7;
      983: inst = 32'h8220000;
      984: inst = 32'h10408000;
      985: inst = 32'hc4040f8;
      986: inst = 32'h8220000;
      987: inst = 32'h10408000;
      988: inst = 32'hc4040f9;
      989: inst = 32'h8220000;
      990: inst = 32'h10408000;
      991: inst = 32'hc4040fa;
      992: inst = 32'h8220000;
      993: inst = 32'h10408000;
      994: inst = 32'hc4040fb;
      995: inst = 32'h8220000;
      996: inst = 32'h10408000;
      997: inst = 32'hc4040fc;
      998: inst = 32'h8220000;
      999: inst = 32'h10408000;
      1000: inst = 32'hc4040fd;
      1001: inst = 32'h8220000;
      1002: inst = 32'h10408000;
      1003: inst = 32'hc4040fe;
      1004: inst = 32'h8220000;
      1005: inst = 32'h10408000;
      1006: inst = 32'hc4040ff;
      1007: inst = 32'h8220000;
      1008: inst = 32'h10408000;
      1009: inst = 32'hc404100;
      1010: inst = 32'h8220000;
      1011: inst = 32'h10408000;
      1012: inst = 32'hc404101;
      1013: inst = 32'h8220000;
      1014: inst = 32'h10408000;
      1015: inst = 32'hc404102;
      1016: inst = 32'h8220000;
      1017: inst = 32'h10408000;
      1018: inst = 32'hc404103;
      1019: inst = 32'h8220000;
      1020: inst = 32'h10408000;
      1021: inst = 32'hc404104;
      1022: inst = 32'h8220000;
      1023: inst = 32'h10408000;
      1024: inst = 32'hc404105;
      1025: inst = 32'h8220000;
      1026: inst = 32'h10408000;
      1027: inst = 32'hc404106;
      1028: inst = 32'h8220000;
      1029: inst = 32'h10408000;
      1030: inst = 32'hc404107;
      1031: inst = 32'h8220000;
      1032: inst = 32'h10408000;
      1033: inst = 32'hc404108;
      1034: inst = 32'h8220000;
      1035: inst = 32'h10408000;
      1036: inst = 32'hc404109;
      1037: inst = 32'h8220000;
      1038: inst = 32'h10408000;
      1039: inst = 32'hc40410a;
      1040: inst = 32'h8220000;
      1041: inst = 32'h10408000;
      1042: inst = 32'hc40410c;
      1043: inst = 32'h8220000;
      1044: inst = 32'h10408000;
      1045: inst = 32'hc40410d;
      1046: inst = 32'h8220000;
      1047: inst = 32'h10408000;
      1048: inst = 32'hc40410e;
      1049: inst = 32'h8220000;
      1050: inst = 32'h10408000;
      1051: inst = 32'hc40410f;
      1052: inst = 32'h8220000;
      1053: inst = 32'h10408000;
      1054: inst = 32'hc404110;
      1055: inst = 32'h8220000;
      1056: inst = 32'h10408000;
      1057: inst = 32'hc404111;
      1058: inst = 32'h8220000;
      1059: inst = 32'h10408000;
      1060: inst = 32'hc404112;
      1061: inst = 32'h8220000;
      1062: inst = 32'h10408000;
      1063: inst = 32'hc404113;
      1064: inst = 32'h8220000;
      1065: inst = 32'h10408000;
      1066: inst = 32'hc404114;
      1067: inst = 32'h8220000;
      1068: inst = 32'h10408000;
      1069: inst = 32'hc404115;
      1070: inst = 32'h8220000;
      1071: inst = 32'h10408000;
      1072: inst = 32'hc404116;
      1073: inst = 32'h8220000;
      1074: inst = 32'h10408000;
      1075: inst = 32'hc404117;
      1076: inst = 32'h8220000;
      1077: inst = 32'h10408000;
      1078: inst = 32'hc404118;
      1079: inst = 32'h8220000;
      1080: inst = 32'h10408000;
      1081: inst = 32'hc404119;
      1082: inst = 32'h8220000;
      1083: inst = 32'h10408000;
      1084: inst = 32'hc40411a;
      1085: inst = 32'h8220000;
      1086: inst = 32'h10408000;
      1087: inst = 32'hc40411b;
      1088: inst = 32'h8220000;
      1089: inst = 32'h10408000;
      1090: inst = 32'hc40411c;
      1091: inst = 32'h8220000;
      1092: inst = 32'h10408000;
      1093: inst = 32'hc40411d;
      1094: inst = 32'h8220000;
      1095: inst = 32'h10408000;
      1096: inst = 32'hc40411e;
      1097: inst = 32'h8220000;
      1098: inst = 32'h10408000;
      1099: inst = 32'hc40411f;
      1100: inst = 32'h8220000;
      1101: inst = 32'h10408000;
      1102: inst = 32'hc404120;
      1103: inst = 32'h8220000;
      1104: inst = 32'h10408000;
      1105: inst = 32'hc404121;
      1106: inst = 32'h8220000;
      1107: inst = 32'h10408000;
      1108: inst = 32'hc404122;
      1109: inst = 32'h8220000;
      1110: inst = 32'h10408000;
      1111: inst = 32'hc404123;
      1112: inst = 32'h8220000;
      1113: inst = 32'h10408000;
      1114: inst = 32'hc404124;
      1115: inst = 32'h8220000;
      1116: inst = 32'h10408000;
      1117: inst = 32'hc404125;
      1118: inst = 32'h8220000;
      1119: inst = 32'h10408000;
      1120: inst = 32'hc404126;
      1121: inst = 32'h8220000;
      1122: inst = 32'h10408000;
      1123: inst = 32'hc404127;
      1124: inst = 32'h8220000;
      1125: inst = 32'h10408000;
      1126: inst = 32'hc404128;
      1127: inst = 32'h8220000;
      1128: inst = 32'h10408000;
      1129: inst = 32'hc404129;
      1130: inst = 32'h8220000;
      1131: inst = 32'h10408000;
      1132: inst = 32'hc40412a;
      1133: inst = 32'h8220000;
      1134: inst = 32'h10408000;
      1135: inst = 32'hc40412b;
      1136: inst = 32'h8220000;
      1137: inst = 32'h10408000;
      1138: inst = 32'hc40412c;
      1139: inst = 32'h8220000;
      1140: inst = 32'h10408000;
      1141: inst = 32'hc40412d;
      1142: inst = 32'h8220000;
      1143: inst = 32'h10408000;
      1144: inst = 32'hc40412e;
      1145: inst = 32'h8220000;
      1146: inst = 32'h10408000;
      1147: inst = 32'hc40412f;
      1148: inst = 32'h8220000;
      1149: inst = 32'h10408000;
      1150: inst = 32'hc404130;
      1151: inst = 32'h8220000;
      1152: inst = 32'h10408000;
      1153: inst = 32'hc404131;
      1154: inst = 32'h8220000;
      1155: inst = 32'h10408000;
      1156: inst = 32'hc404132;
      1157: inst = 32'h8220000;
      1158: inst = 32'h10408000;
      1159: inst = 32'hc404133;
      1160: inst = 32'h8220000;
      1161: inst = 32'h10408000;
      1162: inst = 32'hc404134;
      1163: inst = 32'h8220000;
      1164: inst = 32'h10408000;
      1165: inst = 32'hc404135;
      1166: inst = 32'h8220000;
      1167: inst = 32'h10408000;
      1168: inst = 32'hc404136;
      1169: inst = 32'h8220000;
      1170: inst = 32'h10408000;
      1171: inst = 32'hc404137;
      1172: inst = 32'h8220000;
      1173: inst = 32'h10408000;
      1174: inst = 32'hc404138;
      1175: inst = 32'h8220000;
      1176: inst = 32'h10408000;
      1177: inst = 32'hc404139;
      1178: inst = 32'h8220000;
      1179: inst = 32'h10408000;
      1180: inst = 32'hc40413a;
      1181: inst = 32'h8220000;
      1182: inst = 32'h10408000;
      1183: inst = 32'hc40413b;
      1184: inst = 32'h8220000;
      1185: inst = 32'h10408000;
      1186: inst = 32'hc40413c;
      1187: inst = 32'h8220000;
      1188: inst = 32'h10408000;
      1189: inst = 32'hc40413d;
      1190: inst = 32'h8220000;
      1191: inst = 32'h10408000;
      1192: inst = 32'hc40413e;
      1193: inst = 32'h8220000;
      1194: inst = 32'h10408000;
      1195: inst = 32'hc40413f;
      1196: inst = 32'h8220000;
      1197: inst = 32'h10408000;
      1198: inst = 32'hc404140;
      1199: inst = 32'h8220000;
      1200: inst = 32'h10408000;
      1201: inst = 32'hc404141;
      1202: inst = 32'h8220000;
      1203: inst = 32'h10408000;
      1204: inst = 32'hc404142;
      1205: inst = 32'h8220000;
      1206: inst = 32'h10408000;
      1207: inst = 32'hc404143;
      1208: inst = 32'h8220000;
      1209: inst = 32'h10408000;
      1210: inst = 32'hc404144;
      1211: inst = 32'h8220000;
      1212: inst = 32'h10408000;
      1213: inst = 32'hc404145;
      1214: inst = 32'h8220000;
      1215: inst = 32'h10408000;
      1216: inst = 32'hc404146;
      1217: inst = 32'h8220000;
      1218: inst = 32'h10408000;
      1219: inst = 32'hc404147;
      1220: inst = 32'h8220000;
      1221: inst = 32'h10408000;
      1222: inst = 32'hc404148;
      1223: inst = 32'h8220000;
      1224: inst = 32'h10408000;
      1225: inst = 32'hc404149;
      1226: inst = 32'h8220000;
      1227: inst = 32'h10408000;
      1228: inst = 32'hc40414a;
      1229: inst = 32'h8220000;
      1230: inst = 32'h10408000;
      1231: inst = 32'hc40414b;
      1232: inst = 32'h8220000;
      1233: inst = 32'h10408000;
      1234: inst = 32'hc40414c;
      1235: inst = 32'h8220000;
      1236: inst = 32'h10408000;
      1237: inst = 32'hc40414d;
      1238: inst = 32'h8220000;
      1239: inst = 32'h10408000;
      1240: inst = 32'hc40414e;
      1241: inst = 32'h8220000;
      1242: inst = 32'h10408000;
      1243: inst = 32'hc40414f;
      1244: inst = 32'h8220000;
      1245: inst = 32'h10408000;
      1246: inst = 32'hc404150;
      1247: inst = 32'h8220000;
      1248: inst = 32'h10408000;
      1249: inst = 32'hc404151;
      1250: inst = 32'h8220000;
      1251: inst = 32'h10408000;
      1252: inst = 32'hc404152;
      1253: inst = 32'h8220000;
      1254: inst = 32'h10408000;
      1255: inst = 32'hc404153;
      1256: inst = 32'h8220000;
      1257: inst = 32'h10408000;
      1258: inst = 32'hc404154;
      1259: inst = 32'h8220000;
      1260: inst = 32'h10408000;
      1261: inst = 32'hc404155;
      1262: inst = 32'h8220000;
      1263: inst = 32'h10408000;
      1264: inst = 32'hc404156;
      1265: inst = 32'h8220000;
      1266: inst = 32'h10408000;
      1267: inst = 32'hc404157;
      1268: inst = 32'h8220000;
      1269: inst = 32'h10408000;
      1270: inst = 32'hc404158;
      1271: inst = 32'h8220000;
      1272: inst = 32'h10408000;
      1273: inst = 32'hc404159;
      1274: inst = 32'h8220000;
      1275: inst = 32'h10408000;
      1276: inst = 32'hc40415a;
      1277: inst = 32'h8220000;
      1278: inst = 32'h10408000;
      1279: inst = 32'hc40415b;
      1280: inst = 32'h8220000;
      1281: inst = 32'h10408000;
      1282: inst = 32'hc40415c;
      1283: inst = 32'h8220000;
      1284: inst = 32'h10408000;
      1285: inst = 32'hc40415d;
      1286: inst = 32'h8220000;
      1287: inst = 32'h10408000;
      1288: inst = 32'hc40415e;
      1289: inst = 32'h8220000;
      1290: inst = 32'h10408000;
      1291: inst = 32'hc40415f;
      1292: inst = 32'h8220000;
      1293: inst = 32'h10408000;
      1294: inst = 32'hc404160;
      1295: inst = 32'h8220000;
      1296: inst = 32'h10408000;
      1297: inst = 32'hc404161;
      1298: inst = 32'h8220000;
      1299: inst = 32'h10408000;
      1300: inst = 32'hc404162;
      1301: inst = 32'h8220000;
      1302: inst = 32'h10408000;
      1303: inst = 32'hc404163;
      1304: inst = 32'h8220000;
      1305: inst = 32'h10408000;
      1306: inst = 32'hc404164;
      1307: inst = 32'h8220000;
      1308: inst = 32'h10408000;
      1309: inst = 32'hc404165;
      1310: inst = 32'h8220000;
      1311: inst = 32'h10408000;
      1312: inst = 32'hc404166;
      1313: inst = 32'h8220000;
      1314: inst = 32'h10408000;
      1315: inst = 32'hc404167;
      1316: inst = 32'h8220000;
      1317: inst = 32'h10408000;
      1318: inst = 32'hc404168;
      1319: inst = 32'h8220000;
      1320: inst = 32'h10408000;
      1321: inst = 32'hc404169;
      1322: inst = 32'h8220000;
      1323: inst = 32'h10408000;
      1324: inst = 32'hc40416a;
      1325: inst = 32'h8220000;
      1326: inst = 32'h10408000;
      1327: inst = 32'hc40416c;
      1328: inst = 32'h8220000;
      1329: inst = 32'h10408000;
      1330: inst = 32'hc40416d;
      1331: inst = 32'h8220000;
      1332: inst = 32'h10408000;
      1333: inst = 32'hc40416e;
      1334: inst = 32'h8220000;
      1335: inst = 32'h10408000;
      1336: inst = 32'hc40416f;
      1337: inst = 32'h8220000;
      1338: inst = 32'h10408000;
      1339: inst = 32'hc404170;
      1340: inst = 32'h8220000;
      1341: inst = 32'h10408000;
      1342: inst = 32'hc404171;
      1343: inst = 32'h8220000;
      1344: inst = 32'h10408000;
      1345: inst = 32'hc404172;
      1346: inst = 32'h8220000;
      1347: inst = 32'h10408000;
      1348: inst = 32'hc404173;
      1349: inst = 32'h8220000;
      1350: inst = 32'h10408000;
      1351: inst = 32'hc404174;
      1352: inst = 32'h8220000;
      1353: inst = 32'h10408000;
      1354: inst = 32'hc404175;
      1355: inst = 32'h8220000;
      1356: inst = 32'h10408000;
      1357: inst = 32'hc404176;
      1358: inst = 32'h8220000;
      1359: inst = 32'h10408000;
      1360: inst = 32'hc404177;
      1361: inst = 32'h8220000;
      1362: inst = 32'h10408000;
      1363: inst = 32'hc404178;
      1364: inst = 32'h8220000;
      1365: inst = 32'h10408000;
      1366: inst = 32'hc404179;
      1367: inst = 32'h8220000;
      1368: inst = 32'h10408000;
      1369: inst = 32'hc40417a;
      1370: inst = 32'h8220000;
      1371: inst = 32'h10408000;
      1372: inst = 32'hc40417b;
      1373: inst = 32'h8220000;
      1374: inst = 32'h10408000;
      1375: inst = 32'hc40417c;
      1376: inst = 32'h8220000;
      1377: inst = 32'h10408000;
      1378: inst = 32'hc40417d;
      1379: inst = 32'h8220000;
      1380: inst = 32'h10408000;
      1381: inst = 32'hc40417e;
      1382: inst = 32'h8220000;
      1383: inst = 32'h10408000;
      1384: inst = 32'hc40417f;
      1385: inst = 32'h8220000;
      1386: inst = 32'h10408000;
      1387: inst = 32'hc404180;
      1388: inst = 32'h8220000;
      1389: inst = 32'h10408000;
      1390: inst = 32'hc404181;
      1391: inst = 32'h8220000;
      1392: inst = 32'h10408000;
      1393: inst = 32'hc404182;
      1394: inst = 32'h8220000;
      1395: inst = 32'h10408000;
      1396: inst = 32'hc404183;
      1397: inst = 32'h8220000;
      1398: inst = 32'h10408000;
      1399: inst = 32'hc404184;
      1400: inst = 32'h8220000;
      1401: inst = 32'h10408000;
      1402: inst = 32'hc404185;
      1403: inst = 32'h8220000;
      1404: inst = 32'h10408000;
      1405: inst = 32'hc404186;
      1406: inst = 32'h8220000;
      1407: inst = 32'h10408000;
      1408: inst = 32'hc404187;
      1409: inst = 32'h8220000;
      1410: inst = 32'h10408000;
      1411: inst = 32'hc404188;
      1412: inst = 32'h8220000;
      1413: inst = 32'h10408000;
      1414: inst = 32'hc404189;
      1415: inst = 32'h8220000;
      1416: inst = 32'h10408000;
      1417: inst = 32'hc40418a;
      1418: inst = 32'h8220000;
      1419: inst = 32'h10408000;
      1420: inst = 32'hc40418b;
      1421: inst = 32'h8220000;
      1422: inst = 32'h10408000;
      1423: inst = 32'hc40418c;
      1424: inst = 32'h8220000;
      1425: inst = 32'h10408000;
      1426: inst = 32'hc40418d;
      1427: inst = 32'h8220000;
      1428: inst = 32'h10408000;
      1429: inst = 32'hc40418e;
      1430: inst = 32'h8220000;
      1431: inst = 32'h10408000;
      1432: inst = 32'hc40418f;
      1433: inst = 32'h8220000;
      1434: inst = 32'h10408000;
      1435: inst = 32'hc404190;
      1436: inst = 32'h8220000;
      1437: inst = 32'h10408000;
      1438: inst = 32'hc404191;
      1439: inst = 32'h8220000;
      1440: inst = 32'h10408000;
      1441: inst = 32'hc404192;
      1442: inst = 32'h8220000;
      1443: inst = 32'h10408000;
      1444: inst = 32'hc404193;
      1445: inst = 32'h8220000;
      1446: inst = 32'h10408000;
      1447: inst = 32'hc404194;
      1448: inst = 32'h8220000;
      1449: inst = 32'h10408000;
      1450: inst = 32'hc404195;
      1451: inst = 32'h8220000;
      1452: inst = 32'h10408000;
      1453: inst = 32'hc404196;
      1454: inst = 32'h8220000;
      1455: inst = 32'h10408000;
      1456: inst = 32'hc404197;
      1457: inst = 32'h8220000;
      1458: inst = 32'h10408000;
      1459: inst = 32'hc404198;
      1460: inst = 32'h8220000;
      1461: inst = 32'h10408000;
      1462: inst = 32'hc404199;
      1463: inst = 32'h8220000;
      1464: inst = 32'h10408000;
      1465: inst = 32'hc40419a;
      1466: inst = 32'h8220000;
      1467: inst = 32'h10408000;
      1468: inst = 32'hc40419b;
      1469: inst = 32'h8220000;
      1470: inst = 32'h10408000;
      1471: inst = 32'hc40419c;
      1472: inst = 32'h8220000;
      1473: inst = 32'h10408000;
      1474: inst = 32'hc40419d;
      1475: inst = 32'h8220000;
      1476: inst = 32'h10408000;
      1477: inst = 32'hc40419e;
      1478: inst = 32'h8220000;
      1479: inst = 32'h10408000;
      1480: inst = 32'hc40419f;
      1481: inst = 32'h8220000;
      1482: inst = 32'h10408000;
      1483: inst = 32'hc4041a0;
      1484: inst = 32'h8220000;
      1485: inst = 32'h10408000;
      1486: inst = 32'hc4041a1;
      1487: inst = 32'h8220000;
      1488: inst = 32'h10408000;
      1489: inst = 32'hc4041a2;
      1490: inst = 32'h8220000;
      1491: inst = 32'h10408000;
      1492: inst = 32'hc4041a3;
      1493: inst = 32'h8220000;
      1494: inst = 32'h10408000;
      1495: inst = 32'hc4041a4;
      1496: inst = 32'h8220000;
      1497: inst = 32'h10408000;
      1498: inst = 32'hc4041a5;
      1499: inst = 32'h8220000;
      1500: inst = 32'h10408000;
      1501: inst = 32'hc4041a6;
      1502: inst = 32'h8220000;
      1503: inst = 32'h10408000;
      1504: inst = 32'hc4041a7;
      1505: inst = 32'h8220000;
      1506: inst = 32'h10408000;
      1507: inst = 32'hc4041a8;
      1508: inst = 32'h8220000;
      1509: inst = 32'h10408000;
      1510: inst = 32'hc4041a9;
      1511: inst = 32'h8220000;
      1512: inst = 32'h10408000;
      1513: inst = 32'hc4041aa;
      1514: inst = 32'h8220000;
      1515: inst = 32'h10408000;
      1516: inst = 32'hc4041ab;
      1517: inst = 32'h8220000;
      1518: inst = 32'h10408000;
      1519: inst = 32'hc4041ac;
      1520: inst = 32'h8220000;
      1521: inst = 32'h10408000;
      1522: inst = 32'hc4041ad;
      1523: inst = 32'h8220000;
      1524: inst = 32'h10408000;
      1525: inst = 32'hc4041ae;
      1526: inst = 32'h8220000;
      1527: inst = 32'h10408000;
      1528: inst = 32'hc4041af;
      1529: inst = 32'h8220000;
      1530: inst = 32'h10408000;
      1531: inst = 32'hc4041b0;
      1532: inst = 32'h8220000;
      1533: inst = 32'h10408000;
      1534: inst = 32'hc4041b1;
      1535: inst = 32'h8220000;
      1536: inst = 32'h10408000;
      1537: inst = 32'hc4041b2;
      1538: inst = 32'h8220000;
      1539: inst = 32'h10408000;
      1540: inst = 32'hc4041b3;
      1541: inst = 32'h8220000;
      1542: inst = 32'h10408000;
      1543: inst = 32'hc4041b4;
      1544: inst = 32'h8220000;
      1545: inst = 32'h10408000;
      1546: inst = 32'hc4041b5;
      1547: inst = 32'h8220000;
      1548: inst = 32'h10408000;
      1549: inst = 32'hc4041b6;
      1550: inst = 32'h8220000;
      1551: inst = 32'h10408000;
      1552: inst = 32'hc4041b7;
      1553: inst = 32'h8220000;
      1554: inst = 32'h10408000;
      1555: inst = 32'hc4041b8;
      1556: inst = 32'h8220000;
      1557: inst = 32'h10408000;
      1558: inst = 32'hc4041b9;
      1559: inst = 32'h8220000;
      1560: inst = 32'h10408000;
      1561: inst = 32'hc4041ba;
      1562: inst = 32'h8220000;
      1563: inst = 32'h10408000;
      1564: inst = 32'hc4041bb;
      1565: inst = 32'h8220000;
      1566: inst = 32'h10408000;
      1567: inst = 32'hc4041bc;
      1568: inst = 32'h8220000;
      1569: inst = 32'h10408000;
      1570: inst = 32'hc4041bd;
      1571: inst = 32'h8220000;
      1572: inst = 32'h10408000;
      1573: inst = 32'hc4041be;
      1574: inst = 32'h8220000;
      1575: inst = 32'h10408000;
      1576: inst = 32'hc4041bf;
      1577: inst = 32'h8220000;
      1578: inst = 32'h10408000;
      1579: inst = 32'hc4041c0;
      1580: inst = 32'h8220000;
      1581: inst = 32'h10408000;
      1582: inst = 32'hc4041c1;
      1583: inst = 32'h8220000;
      1584: inst = 32'h10408000;
      1585: inst = 32'hc4041c2;
      1586: inst = 32'h8220000;
      1587: inst = 32'h10408000;
      1588: inst = 32'hc4041c3;
      1589: inst = 32'h8220000;
      1590: inst = 32'h10408000;
      1591: inst = 32'hc4041c4;
      1592: inst = 32'h8220000;
      1593: inst = 32'h10408000;
      1594: inst = 32'hc4041c5;
      1595: inst = 32'h8220000;
      1596: inst = 32'h10408000;
      1597: inst = 32'hc4041c6;
      1598: inst = 32'h8220000;
      1599: inst = 32'h10408000;
      1600: inst = 32'hc4041c7;
      1601: inst = 32'h8220000;
      1602: inst = 32'h10408000;
      1603: inst = 32'hc4041c8;
      1604: inst = 32'h8220000;
      1605: inst = 32'h10408000;
      1606: inst = 32'hc4041c9;
      1607: inst = 32'h8220000;
      1608: inst = 32'h10408000;
      1609: inst = 32'hc4041ca;
      1610: inst = 32'h8220000;
      1611: inst = 32'h10408000;
      1612: inst = 32'hc4041cc;
      1613: inst = 32'h8220000;
      1614: inst = 32'h10408000;
      1615: inst = 32'hc4041cd;
      1616: inst = 32'h8220000;
      1617: inst = 32'h10408000;
      1618: inst = 32'hc4041ce;
      1619: inst = 32'h8220000;
      1620: inst = 32'h10408000;
      1621: inst = 32'hc4041cf;
      1622: inst = 32'h8220000;
      1623: inst = 32'h10408000;
      1624: inst = 32'hc4041d0;
      1625: inst = 32'h8220000;
      1626: inst = 32'h10408000;
      1627: inst = 32'hc4041d1;
      1628: inst = 32'h8220000;
      1629: inst = 32'h10408000;
      1630: inst = 32'hc4041d2;
      1631: inst = 32'h8220000;
      1632: inst = 32'h10408000;
      1633: inst = 32'hc4041d3;
      1634: inst = 32'h8220000;
      1635: inst = 32'h10408000;
      1636: inst = 32'hc4041d4;
      1637: inst = 32'h8220000;
      1638: inst = 32'h10408000;
      1639: inst = 32'hc4041d5;
      1640: inst = 32'h8220000;
      1641: inst = 32'h10408000;
      1642: inst = 32'hc4041d6;
      1643: inst = 32'h8220000;
      1644: inst = 32'h10408000;
      1645: inst = 32'hc4041d7;
      1646: inst = 32'h8220000;
      1647: inst = 32'h10408000;
      1648: inst = 32'hc4041d8;
      1649: inst = 32'h8220000;
      1650: inst = 32'h10408000;
      1651: inst = 32'hc4041d9;
      1652: inst = 32'h8220000;
      1653: inst = 32'h10408000;
      1654: inst = 32'hc404206;
      1655: inst = 32'h8220000;
      1656: inst = 32'h10408000;
      1657: inst = 32'hc404207;
      1658: inst = 32'h8220000;
      1659: inst = 32'h10408000;
      1660: inst = 32'hc404208;
      1661: inst = 32'h8220000;
      1662: inst = 32'h10408000;
      1663: inst = 32'hc404209;
      1664: inst = 32'h8220000;
      1665: inst = 32'h10408000;
      1666: inst = 32'hc40420a;
      1667: inst = 32'h8220000;
      1668: inst = 32'h10408000;
      1669: inst = 32'hc40420b;
      1670: inst = 32'h8220000;
      1671: inst = 32'h10408000;
      1672: inst = 32'hc40420c;
      1673: inst = 32'h8220000;
      1674: inst = 32'h10408000;
      1675: inst = 32'hc40420d;
      1676: inst = 32'h8220000;
      1677: inst = 32'h10408000;
      1678: inst = 32'hc40420e;
      1679: inst = 32'h8220000;
      1680: inst = 32'h10408000;
      1681: inst = 32'hc40420f;
      1682: inst = 32'h8220000;
      1683: inst = 32'h10408000;
      1684: inst = 32'hc404210;
      1685: inst = 32'h8220000;
      1686: inst = 32'h10408000;
      1687: inst = 32'hc404211;
      1688: inst = 32'h8220000;
      1689: inst = 32'h10408000;
      1690: inst = 32'hc404212;
      1691: inst = 32'h8220000;
      1692: inst = 32'h10408000;
      1693: inst = 32'hc404213;
      1694: inst = 32'h8220000;
      1695: inst = 32'h10408000;
      1696: inst = 32'hc404214;
      1697: inst = 32'h8220000;
      1698: inst = 32'h10408000;
      1699: inst = 32'hc404215;
      1700: inst = 32'h8220000;
      1701: inst = 32'h10408000;
      1702: inst = 32'hc404216;
      1703: inst = 32'h8220000;
      1704: inst = 32'h10408000;
      1705: inst = 32'hc404217;
      1706: inst = 32'h8220000;
      1707: inst = 32'h10408000;
      1708: inst = 32'hc404218;
      1709: inst = 32'h8220000;
      1710: inst = 32'h10408000;
      1711: inst = 32'hc404219;
      1712: inst = 32'h8220000;
      1713: inst = 32'h10408000;
      1714: inst = 32'hc40421a;
      1715: inst = 32'h8220000;
      1716: inst = 32'h10408000;
      1717: inst = 32'hc40421b;
      1718: inst = 32'h8220000;
      1719: inst = 32'h10408000;
      1720: inst = 32'hc40421c;
      1721: inst = 32'h8220000;
      1722: inst = 32'h10408000;
      1723: inst = 32'hc40421d;
      1724: inst = 32'h8220000;
      1725: inst = 32'h10408000;
      1726: inst = 32'hc40421e;
      1727: inst = 32'h8220000;
      1728: inst = 32'h10408000;
      1729: inst = 32'hc40421f;
      1730: inst = 32'h8220000;
      1731: inst = 32'h10408000;
      1732: inst = 32'hc404220;
      1733: inst = 32'h8220000;
      1734: inst = 32'h10408000;
      1735: inst = 32'hc404221;
      1736: inst = 32'h8220000;
      1737: inst = 32'h10408000;
      1738: inst = 32'hc404222;
      1739: inst = 32'h8220000;
      1740: inst = 32'h10408000;
      1741: inst = 32'hc404223;
      1742: inst = 32'h8220000;
      1743: inst = 32'h10408000;
      1744: inst = 32'hc404224;
      1745: inst = 32'h8220000;
      1746: inst = 32'h10408000;
      1747: inst = 32'hc404225;
      1748: inst = 32'h8220000;
      1749: inst = 32'h10408000;
      1750: inst = 32'hc404226;
      1751: inst = 32'h8220000;
      1752: inst = 32'h10408000;
      1753: inst = 32'hc404227;
      1754: inst = 32'h8220000;
      1755: inst = 32'h10408000;
      1756: inst = 32'hc404228;
      1757: inst = 32'h8220000;
      1758: inst = 32'h10408000;
      1759: inst = 32'hc404229;
      1760: inst = 32'h8220000;
      1761: inst = 32'h10408000;
      1762: inst = 32'hc40422a;
      1763: inst = 32'h8220000;
      1764: inst = 32'h10408000;
      1765: inst = 32'hc40422c;
      1766: inst = 32'h8220000;
      1767: inst = 32'h10408000;
      1768: inst = 32'hc40422d;
      1769: inst = 32'h8220000;
      1770: inst = 32'h10408000;
      1771: inst = 32'hc40422e;
      1772: inst = 32'h8220000;
      1773: inst = 32'h10408000;
      1774: inst = 32'hc40422f;
      1775: inst = 32'h8220000;
      1776: inst = 32'h10408000;
      1777: inst = 32'hc404230;
      1778: inst = 32'h8220000;
      1779: inst = 32'h10408000;
      1780: inst = 32'hc404231;
      1781: inst = 32'h8220000;
      1782: inst = 32'h10408000;
      1783: inst = 32'hc404232;
      1784: inst = 32'h8220000;
      1785: inst = 32'h10408000;
      1786: inst = 32'hc404233;
      1787: inst = 32'h8220000;
      1788: inst = 32'h10408000;
      1789: inst = 32'hc404234;
      1790: inst = 32'h8220000;
      1791: inst = 32'h10408000;
      1792: inst = 32'hc404235;
      1793: inst = 32'h8220000;
      1794: inst = 32'h10408000;
      1795: inst = 32'hc404236;
      1796: inst = 32'h8220000;
      1797: inst = 32'h10408000;
      1798: inst = 32'hc404237;
      1799: inst = 32'h8220000;
      1800: inst = 32'h10408000;
      1801: inst = 32'hc404238;
      1802: inst = 32'h8220000;
      1803: inst = 32'h10408000;
      1804: inst = 32'hc404239;
      1805: inst = 32'h8220000;
      1806: inst = 32'h10408000;
      1807: inst = 32'hc40423a;
      1808: inst = 32'h8220000;
      1809: inst = 32'h10408000;
      1810: inst = 32'hc40423b;
      1811: inst = 32'h8220000;
      1812: inst = 32'h10408000;
      1813: inst = 32'hc404264;
      1814: inst = 32'h8220000;
      1815: inst = 32'h10408000;
      1816: inst = 32'hc404265;
      1817: inst = 32'h8220000;
      1818: inst = 32'h10408000;
      1819: inst = 32'hc404266;
      1820: inst = 32'h8220000;
      1821: inst = 32'h10408000;
      1822: inst = 32'hc404267;
      1823: inst = 32'h8220000;
      1824: inst = 32'h10408000;
      1825: inst = 32'hc404268;
      1826: inst = 32'h8220000;
      1827: inst = 32'h10408000;
      1828: inst = 32'hc404269;
      1829: inst = 32'h8220000;
      1830: inst = 32'h10408000;
      1831: inst = 32'hc40426a;
      1832: inst = 32'h8220000;
      1833: inst = 32'h10408000;
      1834: inst = 32'hc40426b;
      1835: inst = 32'h8220000;
      1836: inst = 32'h10408000;
      1837: inst = 32'hc40426c;
      1838: inst = 32'h8220000;
      1839: inst = 32'h10408000;
      1840: inst = 32'hc40426d;
      1841: inst = 32'h8220000;
      1842: inst = 32'h10408000;
      1843: inst = 32'hc40426e;
      1844: inst = 32'h8220000;
      1845: inst = 32'h10408000;
      1846: inst = 32'hc40426f;
      1847: inst = 32'h8220000;
      1848: inst = 32'h10408000;
      1849: inst = 32'hc404270;
      1850: inst = 32'h8220000;
      1851: inst = 32'h10408000;
      1852: inst = 32'hc404271;
      1853: inst = 32'h8220000;
      1854: inst = 32'h10408000;
      1855: inst = 32'hc404272;
      1856: inst = 32'h8220000;
      1857: inst = 32'h10408000;
      1858: inst = 32'hc404273;
      1859: inst = 32'h8220000;
      1860: inst = 32'h10408000;
      1861: inst = 32'hc404274;
      1862: inst = 32'h8220000;
      1863: inst = 32'h10408000;
      1864: inst = 32'hc404275;
      1865: inst = 32'h8220000;
      1866: inst = 32'h10408000;
      1867: inst = 32'hc404276;
      1868: inst = 32'h8220000;
      1869: inst = 32'h10408000;
      1870: inst = 32'hc404277;
      1871: inst = 32'h8220000;
      1872: inst = 32'h10408000;
      1873: inst = 32'hc404278;
      1874: inst = 32'h8220000;
      1875: inst = 32'h10408000;
      1876: inst = 32'hc404279;
      1877: inst = 32'h8220000;
      1878: inst = 32'h10408000;
      1879: inst = 32'hc40427a;
      1880: inst = 32'h8220000;
      1881: inst = 32'h10408000;
      1882: inst = 32'hc40427b;
      1883: inst = 32'h8220000;
      1884: inst = 32'h10408000;
      1885: inst = 32'hc40427c;
      1886: inst = 32'h8220000;
      1887: inst = 32'h10408000;
      1888: inst = 32'hc40427d;
      1889: inst = 32'h8220000;
      1890: inst = 32'h10408000;
      1891: inst = 32'hc40427e;
      1892: inst = 32'h8220000;
      1893: inst = 32'h10408000;
      1894: inst = 32'hc40427f;
      1895: inst = 32'h8220000;
      1896: inst = 32'h10408000;
      1897: inst = 32'hc404280;
      1898: inst = 32'h8220000;
      1899: inst = 32'h10408000;
      1900: inst = 32'hc404281;
      1901: inst = 32'h8220000;
      1902: inst = 32'h10408000;
      1903: inst = 32'hc404282;
      1904: inst = 32'h8220000;
      1905: inst = 32'h10408000;
      1906: inst = 32'hc404283;
      1907: inst = 32'h8220000;
      1908: inst = 32'h10408000;
      1909: inst = 32'hc404284;
      1910: inst = 32'h8220000;
      1911: inst = 32'h10408000;
      1912: inst = 32'hc404285;
      1913: inst = 32'h8220000;
      1914: inst = 32'h10408000;
      1915: inst = 32'hc404286;
      1916: inst = 32'h8220000;
      1917: inst = 32'h10408000;
      1918: inst = 32'hc404287;
      1919: inst = 32'h8220000;
      1920: inst = 32'h10408000;
      1921: inst = 32'hc404288;
      1922: inst = 32'h8220000;
      1923: inst = 32'h10408000;
      1924: inst = 32'hc404289;
      1925: inst = 32'h8220000;
      1926: inst = 32'h10408000;
      1927: inst = 32'hc40428a;
      1928: inst = 32'h8220000;
      1929: inst = 32'h10408000;
      1930: inst = 32'hc40428c;
      1931: inst = 32'h8220000;
      1932: inst = 32'h10408000;
      1933: inst = 32'hc40428d;
      1934: inst = 32'h8220000;
      1935: inst = 32'h10408000;
      1936: inst = 32'hc40428e;
      1937: inst = 32'h8220000;
      1938: inst = 32'h10408000;
      1939: inst = 32'hc40428f;
      1940: inst = 32'h8220000;
      1941: inst = 32'h10408000;
      1942: inst = 32'hc404290;
      1943: inst = 32'h8220000;
      1944: inst = 32'h10408000;
      1945: inst = 32'hc404291;
      1946: inst = 32'h8220000;
      1947: inst = 32'h10408000;
      1948: inst = 32'hc404292;
      1949: inst = 32'h8220000;
      1950: inst = 32'h10408000;
      1951: inst = 32'hc404293;
      1952: inst = 32'h8220000;
      1953: inst = 32'h10408000;
      1954: inst = 32'hc404294;
      1955: inst = 32'h8220000;
      1956: inst = 32'h10408000;
      1957: inst = 32'hc404295;
      1958: inst = 32'h8220000;
      1959: inst = 32'h10408000;
      1960: inst = 32'hc404296;
      1961: inst = 32'h8220000;
      1962: inst = 32'h10408000;
      1963: inst = 32'hc404297;
      1964: inst = 32'h8220000;
      1965: inst = 32'h10408000;
      1966: inst = 32'hc404298;
      1967: inst = 32'h8220000;
      1968: inst = 32'h10408000;
      1969: inst = 32'hc404299;
      1970: inst = 32'h8220000;
      1971: inst = 32'h10408000;
      1972: inst = 32'hc40429a;
      1973: inst = 32'h8220000;
      1974: inst = 32'h10408000;
      1975: inst = 32'hc40429b;
      1976: inst = 32'h8220000;
      1977: inst = 32'h10408000;
      1978: inst = 32'hc4042c4;
      1979: inst = 32'h8220000;
      1980: inst = 32'h10408000;
      1981: inst = 32'hc4042c5;
      1982: inst = 32'h8220000;
      1983: inst = 32'h10408000;
      1984: inst = 32'hc4042c6;
      1985: inst = 32'h8220000;
      1986: inst = 32'h10408000;
      1987: inst = 32'hc4042c7;
      1988: inst = 32'h8220000;
      1989: inst = 32'h10408000;
      1990: inst = 32'hc4042c8;
      1991: inst = 32'h8220000;
      1992: inst = 32'h10408000;
      1993: inst = 32'hc4042c9;
      1994: inst = 32'h8220000;
      1995: inst = 32'h10408000;
      1996: inst = 32'hc4042ca;
      1997: inst = 32'h8220000;
      1998: inst = 32'h10408000;
      1999: inst = 32'hc4042cb;
      2000: inst = 32'h8220000;
      2001: inst = 32'h10408000;
      2002: inst = 32'hc4042cc;
      2003: inst = 32'h8220000;
      2004: inst = 32'h10408000;
      2005: inst = 32'hc4042cd;
      2006: inst = 32'h8220000;
      2007: inst = 32'h10408000;
      2008: inst = 32'hc4042ce;
      2009: inst = 32'h8220000;
      2010: inst = 32'h10408000;
      2011: inst = 32'hc4042cf;
      2012: inst = 32'h8220000;
      2013: inst = 32'h10408000;
      2014: inst = 32'hc4042d0;
      2015: inst = 32'h8220000;
      2016: inst = 32'h10408000;
      2017: inst = 32'hc4042d1;
      2018: inst = 32'h8220000;
      2019: inst = 32'h10408000;
      2020: inst = 32'hc4042d2;
      2021: inst = 32'h8220000;
      2022: inst = 32'h10408000;
      2023: inst = 32'hc4042d3;
      2024: inst = 32'h8220000;
      2025: inst = 32'h10408000;
      2026: inst = 32'hc4042d4;
      2027: inst = 32'h8220000;
      2028: inst = 32'h10408000;
      2029: inst = 32'hc4042d5;
      2030: inst = 32'h8220000;
      2031: inst = 32'h10408000;
      2032: inst = 32'hc4042d6;
      2033: inst = 32'h8220000;
      2034: inst = 32'h10408000;
      2035: inst = 32'hc4042d7;
      2036: inst = 32'h8220000;
      2037: inst = 32'h10408000;
      2038: inst = 32'hc4042d8;
      2039: inst = 32'h8220000;
      2040: inst = 32'h10408000;
      2041: inst = 32'hc4042d9;
      2042: inst = 32'h8220000;
      2043: inst = 32'h10408000;
      2044: inst = 32'hc4042da;
      2045: inst = 32'h8220000;
      2046: inst = 32'h10408000;
      2047: inst = 32'hc4042db;
      2048: inst = 32'h8220000;
      2049: inst = 32'h10408000;
      2050: inst = 32'hc4042dc;
      2051: inst = 32'h8220000;
      2052: inst = 32'h10408000;
      2053: inst = 32'hc4042dd;
      2054: inst = 32'h8220000;
      2055: inst = 32'h10408000;
      2056: inst = 32'hc4042de;
      2057: inst = 32'h8220000;
      2058: inst = 32'h10408000;
      2059: inst = 32'hc4042df;
      2060: inst = 32'h8220000;
      2061: inst = 32'h10408000;
      2062: inst = 32'hc4042e0;
      2063: inst = 32'h8220000;
      2064: inst = 32'h10408000;
      2065: inst = 32'hc4042e1;
      2066: inst = 32'h8220000;
      2067: inst = 32'h10408000;
      2068: inst = 32'hc4042e2;
      2069: inst = 32'h8220000;
      2070: inst = 32'h10408000;
      2071: inst = 32'hc4042e3;
      2072: inst = 32'h8220000;
      2073: inst = 32'h10408000;
      2074: inst = 32'hc4042e4;
      2075: inst = 32'h8220000;
      2076: inst = 32'h10408000;
      2077: inst = 32'hc4042e5;
      2078: inst = 32'h8220000;
      2079: inst = 32'h10408000;
      2080: inst = 32'hc4042e6;
      2081: inst = 32'h8220000;
      2082: inst = 32'h10408000;
      2083: inst = 32'hc4042e7;
      2084: inst = 32'h8220000;
      2085: inst = 32'h10408000;
      2086: inst = 32'hc4042e8;
      2087: inst = 32'h8220000;
      2088: inst = 32'h10408000;
      2089: inst = 32'hc4042e9;
      2090: inst = 32'h8220000;
      2091: inst = 32'h10408000;
      2092: inst = 32'hc4042ee;
      2093: inst = 32'h8220000;
      2094: inst = 32'h10408000;
      2095: inst = 32'hc4042ef;
      2096: inst = 32'h8220000;
      2097: inst = 32'h10408000;
      2098: inst = 32'hc4042f0;
      2099: inst = 32'h8220000;
      2100: inst = 32'h10408000;
      2101: inst = 32'hc4042f1;
      2102: inst = 32'h8220000;
      2103: inst = 32'h10408000;
      2104: inst = 32'hc4042f2;
      2105: inst = 32'h8220000;
      2106: inst = 32'h10408000;
      2107: inst = 32'hc4042f3;
      2108: inst = 32'h8220000;
      2109: inst = 32'h10408000;
      2110: inst = 32'hc4042f4;
      2111: inst = 32'h8220000;
      2112: inst = 32'h10408000;
      2113: inst = 32'hc4042f5;
      2114: inst = 32'h8220000;
      2115: inst = 32'h10408000;
      2116: inst = 32'hc4042f6;
      2117: inst = 32'h8220000;
      2118: inst = 32'h10408000;
      2119: inst = 32'hc4042f7;
      2120: inst = 32'h8220000;
      2121: inst = 32'h10408000;
      2122: inst = 32'hc4042f8;
      2123: inst = 32'h8220000;
      2124: inst = 32'h10408000;
      2125: inst = 32'hc4042f9;
      2126: inst = 32'h8220000;
      2127: inst = 32'h10408000;
      2128: inst = 32'hc4042fa;
      2129: inst = 32'h8220000;
      2130: inst = 32'h10408000;
      2131: inst = 32'hc4042fb;
      2132: inst = 32'h8220000;
      2133: inst = 32'h10408000;
      2134: inst = 32'hc404324;
      2135: inst = 32'h8220000;
      2136: inst = 32'h10408000;
      2137: inst = 32'hc404325;
      2138: inst = 32'h8220000;
      2139: inst = 32'h10408000;
      2140: inst = 32'hc404326;
      2141: inst = 32'h8220000;
      2142: inst = 32'h10408000;
      2143: inst = 32'hc404327;
      2144: inst = 32'h8220000;
      2145: inst = 32'h10408000;
      2146: inst = 32'hc404328;
      2147: inst = 32'h8220000;
      2148: inst = 32'h10408000;
      2149: inst = 32'hc404329;
      2150: inst = 32'h8220000;
      2151: inst = 32'h10408000;
      2152: inst = 32'hc40432a;
      2153: inst = 32'h8220000;
      2154: inst = 32'h10408000;
      2155: inst = 32'hc40432b;
      2156: inst = 32'h8220000;
      2157: inst = 32'h10408000;
      2158: inst = 32'hc40432c;
      2159: inst = 32'h8220000;
      2160: inst = 32'h10408000;
      2161: inst = 32'hc40432d;
      2162: inst = 32'h8220000;
      2163: inst = 32'h10408000;
      2164: inst = 32'hc40432e;
      2165: inst = 32'h8220000;
      2166: inst = 32'h10408000;
      2167: inst = 32'hc40432f;
      2168: inst = 32'h8220000;
      2169: inst = 32'h10408000;
      2170: inst = 32'hc404330;
      2171: inst = 32'h8220000;
      2172: inst = 32'h10408000;
      2173: inst = 32'hc404331;
      2174: inst = 32'h8220000;
      2175: inst = 32'h10408000;
      2176: inst = 32'hc404332;
      2177: inst = 32'h8220000;
      2178: inst = 32'h10408000;
      2179: inst = 32'hc404333;
      2180: inst = 32'h8220000;
      2181: inst = 32'h10408000;
      2182: inst = 32'hc404334;
      2183: inst = 32'h8220000;
      2184: inst = 32'h10408000;
      2185: inst = 32'hc404335;
      2186: inst = 32'h8220000;
      2187: inst = 32'h10408000;
      2188: inst = 32'hc404336;
      2189: inst = 32'h8220000;
      2190: inst = 32'h10408000;
      2191: inst = 32'hc404337;
      2192: inst = 32'h8220000;
      2193: inst = 32'h10408000;
      2194: inst = 32'hc404338;
      2195: inst = 32'h8220000;
      2196: inst = 32'h10408000;
      2197: inst = 32'hc404339;
      2198: inst = 32'h8220000;
      2199: inst = 32'h10408000;
      2200: inst = 32'hc40433a;
      2201: inst = 32'h8220000;
      2202: inst = 32'h10408000;
      2203: inst = 32'hc40433b;
      2204: inst = 32'h8220000;
      2205: inst = 32'h10408000;
      2206: inst = 32'hc40433c;
      2207: inst = 32'h8220000;
      2208: inst = 32'h10408000;
      2209: inst = 32'hc40433d;
      2210: inst = 32'h8220000;
      2211: inst = 32'h10408000;
      2212: inst = 32'hc40433e;
      2213: inst = 32'h8220000;
      2214: inst = 32'h10408000;
      2215: inst = 32'hc40433f;
      2216: inst = 32'h8220000;
      2217: inst = 32'h10408000;
      2218: inst = 32'hc404340;
      2219: inst = 32'h8220000;
      2220: inst = 32'h10408000;
      2221: inst = 32'hc404341;
      2222: inst = 32'h8220000;
      2223: inst = 32'h10408000;
      2224: inst = 32'hc404342;
      2225: inst = 32'h8220000;
      2226: inst = 32'h10408000;
      2227: inst = 32'hc404343;
      2228: inst = 32'h8220000;
      2229: inst = 32'h10408000;
      2230: inst = 32'hc404344;
      2231: inst = 32'h8220000;
      2232: inst = 32'h10408000;
      2233: inst = 32'hc404345;
      2234: inst = 32'h8220000;
      2235: inst = 32'h10408000;
      2236: inst = 32'hc404346;
      2237: inst = 32'h8220000;
      2238: inst = 32'h10408000;
      2239: inst = 32'hc404347;
      2240: inst = 32'h8220000;
      2241: inst = 32'h10408000;
      2242: inst = 32'hc404348;
      2243: inst = 32'h8220000;
      2244: inst = 32'h10408000;
      2245: inst = 32'hc40434f;
      2246: inst = 32'h8220000;
      2247: inst = 32'h10408000;
      2248: inst = 32'hc404350;
      2249: inst = 32'h8220000;
      2250: inst = 32'h10408000;
      2251: inst = 32'hc404351;
      2252: inst = 32'h8220000;
      2253: inst = 32'h10408000;
      2254: inst = 32'hc404352;
      2255: inst = 32'h8220000;
      2256: inst = 32'h10408000;
      2257: inst = 32'hc404353;
      2258: inst = 32'h8220000;
      2259: inst = 32'h10408000;
      2260: inst = 32'hc404354;
      2261: inst = 32'h8220000;
      2262: inst = 32'h10408000;
      2263: inst = 32'hc404355;
      2264: inst = 32'h8220000;
      2265: inst = 32'h10408000;
      2266: inst = 32'hc404356;
      2267: inst = 32'h8220000;
      2268: inst = 32'h10408000;
      2269: inst = 32'hc404357;
      2270: inst = 32'h8220000;
      2271: inst = 32'h10408000;
      2272: inst = 32'hc404358;
      2273: inst = 32'h8220000;
      2274: inst = 32'h10408000;
      2275: inst = 32'hc404359;
      2276: inst = 32'h8220000;
      2277: inst = 32'h10408000;
      2278: inst = 32'hc40435a;
      2279: inst = 32'h8220000;
      2280: inst = 32'h10408000;
      2281: inst = 32'hc40435b;
      2282: inst = 32'h8220000;
      2283: inst = 32'h10408000;
      2284: inst = 32'hc404384;
      2285: inst = 32'h8220000;
      2286: inst = 32'h10408000;
      2287: inst = 32'hc404385;
      2288: inst = 32'h8220000;
      2289: inst = 32'h10408000;
      2290: inst = 32'hc404386;
      2291: inst = 32'h8220000;
      2292: inst = 32'h10408000;
      2293: inst = 32'hc404387;
      2294: inst = 32'h8220000;
      2295: inst = 32'h10408000;
      2296: inst = 32'hc404388;
      2297: inst = 32'h8220000;
      2298: inst = 32'h10408000;
      2299: inst = 32'hc404389;
      2300: inst = 32'h8220000;
      2301: inst = 32'h10408000;
      2302: inst = 32'hc40438a;
      2303: inst = 32'h8220000;
      2304: inst = 32'h10408000;
      2305: inst = 32'hc40438b;
      2306: inst = 32'h8220000;
      2307: inst = 32'h10408000;
      2308: inst = 32'hc40438c;
      2309: inst = 32'h8220000;
      2310: inst = 32'h10408000;
      2311: inst = 32'hc40438d;
      2312: inst = 32'h8220000;
      2313: inst = 32'h10408000;
      2314: inst = 32'hc40438e;
      2315: inst = 32'h8220000;
      2316: inst = 32'h10408000;
      2317: inst = 32'hc40438f;
      2318: inst = 32'h8220000;
      2319: inst = 32'h10408000;
      2320: inst = 32'hc404390;
      2321: inst = 32'h8220000;
      2322: inst = 32'h10408000;
      2323: inst = 32'hc404391;
      2324: inst = 32'h8220000;
      2325: inst = 32'h10408000;
      2326: inst = 32'hc404392;
      2327: inst = 32'h8220000;
      2328: inst = 32'h10408000;
      2329: inst = 32'hc404393;
      2330: inst = 32'h8220000;
      2331: inst = 32'h10408000;
      2332: inst = 32'hc404394;
      2333: inst = 32'h8220000;
      2334: inst = 32'h10408000;
      2335: inst = 32'hc404395;
      2336: inst = 32'h8220000;
      2337: inst = 32'h10408000;
      2338: inst = 32'hc404396;
      2339: inst = 32'h8220000;
      2340: inst = 32'h10408000;
      2341: inst = 32'hc404397;
      2342: inst = 32'h8220000;
      2343: inst = 32'h10408000;
      2344: inst = 32'hc404398;
      2345: inst = 32'h8220000;
      2346: inst = 32'h10408000;
      2347: inst = 32'hc404399;
      2348: inst = 32'h8220000;
      2349: inst = 32'h10408000;
      2350: inst = 32'hc40439a;
      2351: inst = 32'h8220000;
      2352: inst = 32'h10408000;
      2353: inst = 32'hc40439b;
      2354: inst = 32'h8220000;
      2355: inst = 32'h10408000;
      2356: inst = 32'hc40439c;
      2357: inst = 32'h8220000;
      2358: inst = 32'h10408000;
      2359: inst = 32'hc40439d;
      2360: inst = 32'h8220000;
      2361: inst = 32'h10408000;
      2362: inst = 32'hc40439e;
      2363: inst = 32'h8220000;
      2364: inst = 32'h10408000;
      2365: inst = 32'hc40439f;
      2366: inst = 32'h8220000;
      2367: inst = 32'h10408000;
      2368: inst = 32'hc4043a0;
      2369: inst = 32'h8220000;
      2370: inst = 32'h10408000;
      2371: inst = 32'hc4043a1;
      2372: inst = 32'h8220000;
      2373: inst = 32'h10408000;
      2374: inst = 32'hc4043a2;
      2375: inst = 32'h8220000;
      2376: inst = 32'h10408000;
      2377: inst = 32'hc4043a3;
      2378: inst = 32'h8220000;
      2379: inst = 32'h10408000;
      2380: inst = 32'hc4043a4;
      2381: inst = 32'h8220000;
      2382: inst = 32'h10408000;
      2383: inst = 32'hc4043a5;
      2384: inst = 32'h8220000;
      2385: inst = 32'h10408000;
      2386: inst = 32'hc4043a6;
      2387: inst = 32'h8220000;
      2388: inst = 32'h10408000;
      2389: inst = 32'hc4043b1;
      2390: inst = 32'h8220000;
      2391: inst = 32'h10408000;
      2392: inst = 32'hc4043b2;
      2393: inst = 32'h8220000;
      2394: inst = 32'h10408000;
      2395: inst = 32'hc4043b3;
      2396: inst = 32'h8220000;
      2397: inst = 32'h10408000;
      2398: inst = 32'hc4043b4;
      2399: inst = 32'h8220000;
      2400: inst = 32'h10408000;
      2401: inst = 32'hc4043b5;
      2402: inst = 32'h8220000;
      2403: inst = 32'h10408000;
      2404: inst = 32'hc4043b6;
      2405: inst = 32'h8220000;
      2406: inst = 32'h10408000;
      2407: inst = 32'hc4043b7;
      2408: inst = 32'h8220000;
      2409: inst = 32'h10408000;
      2410: inst = 32'hc4043b8;
      2411: inst = 32'h8220000;
      2412: inst = 32'h10408000;
      2413: inst = 32'hc4043b9;
      2414: inst = 32'h8220000;
      2415: inst = 32'h10408000;
      2416: inst = 32'hc4043ba;
      2417: inst = 32'h8220000;
      2418: inst = 32'h10408000;
      2419: inst = 32'hc4043bb;
      2420: inst = 32'h8220000;
      2421: inst = 32'h10408000;
      2422: inst = 32'hc4043e4;
      2423: inst = 32'h8220000;
      2424: inst = 32'h10408000;
      2425: inst = 32'hc4043e5;
      2426: inst = 32'h8220000;
      2427: inst = 32'h10408000;
      2428: inst = 32'hc4043e6;
      2429: inst = 32'h8220000;
      2430: inst = 32'h10408000;
      2431: inst = 32'hc4043e7;
      2432: inst = 32'h8220000;
      2433: inst = 32'h10408000;
      2434: inst = 32'hc4043e8;
      2435: inst = 32'h8220000;
      2436: inst = 32'h10408000;
      2437: inst = 32'hc4043e9;
      2438: inst = 32'h8220000;
      2439: inst = 32'h10408000;
      2440: inst = 32'hc4043ea;
      2441: inst = 32'h8220000;
      2442: inst = 32'h10408000;
      2443: inst = 32'hc4043eb;
      2444: inst = 32'h8220000;
      2445: inst = 32'h10408000;
      2446: inst = 32'hc4043ec;
      2447: inst = 32'h8220000;
      2448: inst = 32'h10408000;
      2449: inst = 32'hc4043ed;
      2450: inst = 32'h8220000;
      2451: inst = 32'h10408000;
      2452: inst = 32'hc4043ee;
      2453: inst = 32'h8220000;
      2454: inst = 32'h10408000;
      2455: inst = 32'hc4043ef;
      2456: inst = 32'h8220000;
      2457: inst = 32'h10408000;
      2458: inst = 32'hc4043f0;
      2459: inst = 32'h8220000;
      2460: inst = 32'h10408000;
      2461: inst = 32'hc4043f1;
      2462: inst = 32'h8220000;
      2463: inst = 32'h10408000;
      2464: inst = 32'hc4043f2;
      2465: inst = 32'h8220000;
      2466: inst = 32'h10408000;
      2467: inst = 32'hc4043f3;
      2468: inst = 32'h8220000;
      2469: inst = 32'h10408000;
      2470: inst = 32'hc4043f4;
      2471: inst = 32'h8220000;
      2472: inst = 32'h10408000;
      2473: inst = 32'hc4043f5;
      2474: inst = 32'h8220000;
      2475: inst = 32'h10408000;
      2476: inst = 32'hc4043f6;
      2477: inst = 32'h8220000;
      2478: inst = 32'h10408000;
      2479: inst = 32'hc4043f7;
      2480: inst = 32'h8220000;
      2481: inst = 32'h10408000;
      2482: inst = 32'hc4043f8;
      2483: inst = 32'h8220000;
      2484: inst = 32'h10408000;
      2485: inst = 32'hc4043f9;
      2486: inst = 32'h8220000;
      2487: inst = 32'h10408000;
      2488: inst = 32'hc4043fa;
      2489: inst = 32'h8220000;
      2490: inst = 32'h10408000;
      2491: inst = 32'hc4043fb;
      2492: inst = 32'h8220000;
      2493: inst = 32'h10408000;
      2494: inst = 32'hc4043fc;
      2495: inst = 32'h8220000;
      2496: inst = 32'h10408000;
      2497: inst = 32'hc4043fd;
      2498: inst = 32'h8220000;
      2499: inst = 32'h10408000;
      2500: inst = 32'hc4043fe;
      2501: inst = 32'h8220000;
      2502: inst = 32'h10408000;
      2503: inst = 32'hc4043ff;
      2504: inst = 32'h8220000;
      2505: inst = 32'h10408000;
      2506: inst = 32'hc404400;
      2507: inst = 32'h8220000;
      2508: inst = 32'h10408000;
      2509: inst = 32'hc404401;
      2510: inst = 32'h8220000;
      2511: inst = 32'h10408000;
      2512: inst = 32'hc404402;
      2513: inst = 32'h8220000;
      2514: inst = 32'h10408000;
      2515: inst = 32'hc404403;
      2516: inst = 32'h8220000;
      2517: inst = 32'h10408000;
      2518: inst = 32'hc404404;
      2519: inst = 32'h8220000;
      2520: inst = 32'h10408000;
      2521: inst = 32'hc404405;
      2522: inst = 32'h8220000;
      2523: inst = 32'h10408000;
      2524: inst = 32'hc404412;
      2525: inst = 32'h8220000;
      2526: inst = 32'h10408000;
      2527: inst = 32'hc404413;
      2528: inst = 32'h8220000;
      2529: inst = 32'h10408000;
      2530: inst = 32'hc404414;
      2531: inst = 32'h8220000;
      2532: inst = 32'h10408000;
      2533: inst = 32'hc404415;
      2534: inst = 32'h8220000;
      2535: inst = 32'h10408000;
      2536: inst = 32'hc404416;
      2537: inst = 32'h8220000;
      2538: inst = 32'h10408000;
      2539: inst = 32'hc404417;
      2540: inst = 32'h8220000;
      2541: inst = 32'h10408000;
      2542: inst = 32'hc404418;
      2543: inst = 32'h8220000;
      2544: inst = 32'h10408000;
      2545: inst = 32'hc404419;
      2546: inst = 32'h8220000;
      2547: inst = 32'h10408000;
      2548: inst = 32'hc40441a;
      2549: inst = 32'h8220000;
      2550: inst = 32'h10408000;
      2551: inst = 32'hc40441b;
      2552: inst = 32'h8220000;
      2553: inst = 32'h10408000;
      2554: inst = 32'hc404444;
      2555: inst = 32'h8220000;
      2556: inst = 32'h10408000;
      2557: inst = 32'hc404445;
      2558: inst = 32'h8220000;
      2559: inst = 32'h10408000;
      2560: inst = 32'hc404446;
      2561: inst = 32'h8220000;
      2562: inst = 32'h10408000;
      2563: inst = 32'hc404447;
      2564: inst = 32'h8220000;
      2565: inst = 32'h10408000;
      2566: inst = 32'hc404448;
      2567: inst = 32'h8220000;
      2568: inst = 32'h10408000;
      2569: inst = 32'hc404449;
      2570: inst = 32'h8220000;
      2571: inst = 32'h10408000;
      2572: inst = 32'hc40444a;
      2573: inst = 32'h8220000;
      2574: inst = 32'h10408000;
      2575: inst = 32'hc40444b;
      2576: inst = 32'h8220000;
      2577: inst = 32'h10408000;
      2578: inst = 32'hc40444c;
      2579: inst = 32'h8220000;
      2580: inst = 32'h10408000;
      2581: inst = 32'hc40444d;
      2582: inst = 32'h8220000;
      2583: inst = 32'h10408000;
      2584: inst = 32'hc40444e;
      2585: inst = 32'h8220000;
      2586: inst = 32'h10408000;
      2587: inst = 32'hc40444f;
      2588: inst = 32'h8220000;
      2589: inst = 32'h10408000;
      2590: inst = 32'hc404450;
      2591: inst = 32'h8220000;
      2592: inst = 32'h10408000;
      2593: inst = 32'hc404451;
      2594: inst = 32'h8220000;
      2595: inst = 32'h10408000;
      2596: inst = 32'hc404452;
      2597: inst = 32'h8220000;
      2598: inst = 32'h10408000;
      2599: inst = 32'hc404453;
      2600: inst = 32'h8220000;
      2601: inst = 32'h10408000;
      2602: inst = 32'hc404454;
      2603: inst = 32'h8220000;
      2604: inst = 32'h10408000;
      2605: inst = 32'hc404455;
      2606: inst = 32'h8220000;
      2607: inst = 32'h10408000;
      2608: inst = 32'hc404456;
      2609: inst = 32'h8220000;
      2610: inst = 32'h10408000;
      2611: inst = 32'hc404457;
      2612: inst = 32'h8220000;
      2613: inst = 32'h10408000;
      2614: inst = 32'hc404458;
      2615: inst = 32'h8220000;
      2616: inst = 32'h10408000;
      2617: inst = 32'hc404459;
      2618: inst = 32'h8220000;
      2619: inst = 32'h10408000;
      2620: inst = 32'hc40445a;
      2621: inst = 32'h8220000;
      2622: inst = 32'h10408000;
      2623: inst = 32'hc40445b;
      2624: inst = 32'h8220000;
      2625: inst = 32'h10408000;
      2626: inst = 32'hc40445c;
      2627: inst = 32'h8220000;
      2628: inst = 32'h10408000;
      2629: inst = 32'hc40445d;
      2630: inst = 32'h8220000;
      2631: inst = 32'h10408000;
      2632: inst = 32'hc40445e;
      2633: inst = 32'h8220000;
      2634: inst = 32'h10408000;
      2635: inst = 32'hc40445f;
      2636: inst = 32'h8220000;
      2637: inst = 32'h10408000;
      2638: inst = 32'hc404460;
      2639: inst = 32'h8220000;
      2640: inst = 32'h10408000;
      2641: inst = 32'hc404461;
      2642: inst = 32'h8220000;
      2643: inst = 32'h10408000;
      2644: inst = 32'hc404462;
      2645: inst = 32'h8220000;
      2646: inst = 32'h10408000;
      2647: inst = 32'hc404463;
      2648: inst = 32'h8220000;
      2649: inst = 32'h10408000;
      2650: inst = 32'hc404464;
      2651: inst = 32'h8220000;
      2652: inst = 32'h10408000;
      2653: inst = 32'hc404465;
      2654: inst = 32'h8220000;
      2655: inst = 32'h10408000;
      2656: inst = 32'hc404466;
      2657: inst = 32'h8220000;
      2658: inst = 32'h10408000;
      2659: inst = 32'hc404467;
      2660: inst = 32'h8220000;
      2661: inst = 32'h10408000;
      2662: inst = 32'hc404468;
      2663: inst = 32'h8220000;
      2664: inst = 32'h10408000;
      2665: inst = 32'hc404469;
      2666: inst = 32'h8220000;
      2667: inst = 32'h10408000;
      2668: inst = 32'hc40446e;
      2669: inst = 32'h8220000;
      2670: inst = 32'h10408000;
      2671: inst = 32'hc40446f;
      2672: inst = 32'h8220000;
      2673: inst = 32'h10408000;
      2674: inst = 32'hc404470;
      2675: inst = 32'h8220000;
      2676: inst = 32'h10408000;
      2677: inst = 32'hc404471;
      2678: inst = 32'h8220000;
      2679: inst = 32'h10408000;
      2680: inst = 32'hc404472;
      2681: inst = 32'h8220000;
      2682: inst = 32'h10408000;
      2683: inst = 32'hc404473;
      2684: inst = 32'h8220000;
      2685: inst = 32'h10408000;
      2686: inst = 32'hc404474;
      2687: inst = 32'h8220000;
      2688: inst = 32'h10408000;
      2689: inst = 32'hc404475;
      2690: inst = 32'h8220000;
      2691: inst = 32'h10408000;
      2692: inst = 32'hc404476;
      2693: inst = 32'h8220000;
      2694: inst = 32'h10408000;
      2695: inst = 32'hc404477;
      2696: inst = 32'h8220000;
      2697: inst = 32'h10408000;
      2698: inst = 32'hc404478;
      2699: inst = 32'h8220000;
      2700: inst = 32'h10408000;
      2701: inst = 32'hc404479;
      2702: inst = 32'h8220000;
      2703: inst = 32'h10408000;
      2704: inst = 32'hc40447a;
      2705: inst = 32'h8220000;
      2706: inst = 32'h10408000;
      2707: inst = 32'hc40447b;
      2708: inst = 32'h8220000;
      2709: inst = 32'h10408000;
      2710: inst = 32'hc4044a4;
      2711: inst = 32'h8220000;
      2712: inst = 32'h10408000;
      2713: inst = 32'hc4044a5;
      2714: inst = 32'h8220000;
      2715: inst = 32'h10408000;
      2716: inst = 32'hc4044a6;
      2717: inst = 32'h8220000;
      2718: inst = 32'h10408000;
      2719: inst = 32'hc4044a7;
      2720: inst = 32'h8220000;
      2721: inst = 32'h10408000;
      2722: inst = 32'hc4044a8;
      2723: inst = 32'h8220000;
      2724: inst = 32'h10408000;
      2725: inst = 32'hc4044a9;
      2726: inst = 32'h8220000;
      2727: inst = 32'h10408000;
      2728: inst = 32'hc4044aa;
      2729: inst = 32'h8220000;
      2730: inst = 32'h10408000;
      2731: inst = 32'hc4044ab;
      2732: inst = 32'h8220000;
      2733: inst = 32'h10408000;
      2734: inst = 32'hc4044ac;
      2735: inst = 32'h8220000;
      2736: inst = 32'h10408000;
      2737: inst = 32'hc4044ad;
      2738: inst = 32'h8220000;
      2739: inst = 32'h10408000;
      2740: inst = 32'hc4044ae;
      2741: inst = 32'h8220000;
      2742: inst = 32'h10408000;
      2743: inst = 32'hc4044af;
      2744: inst = 32'h8220000;
      2745: inst = 32'h10408000;
      2746: inst = 32'hc4044b0;
      2747: inst = 32'h8220000;
      2748: inst = 32'h10408000;
      2749: inst = 32'hc4044b1;
      2750: inst = 32'h8220000;
      2751: inst = 32'h10408000;
      2752: inst = 32'hc4044b6;
      2753: inst = 32'h8220000;
      2754: inst = 32'h10408000;
      2755: inst = 32'hc4044b7;
      2756: inst = 32'h8220000;
      2757: inst = 32'h10408000;
      2758: inst = 32'hc4044b8;
      2759: inst = 32'h8220000;
      2760: inst = 32'h10408000;
      2761: inst = 32'hc4044b9;
      2762: inst = 32'h8220000;
      2763: inst = 32'h10408000;
      2764: inst = 32'hc4044ba;
      2765: inst = 32'h8220000;
      2766: inst = 32'h10408000;
      2767: inst = 32'hc4044bb;
      2768: inst = 32'h8220000;
      2769: inst = 32'h10408000;
      2770: inst = 32'hc4044bc;
      2771: inst = 32'h8220000;
      2772: inst = 32'h10408000;
      2773: inst = 32'hc4044bd;
      2774: inst = 32'h8220000;
      2775: inst = 32'h10408000;
      2776: inst = 32'hc4044be;
      2777: inst = 32'h8220000;
      2778: inst = 32'h10408000;
      2779: inst = 32'hc4044bf;
      2780: inst = 32'h8220000;
      2781: inst = 32'h10408000;
      2782: inst = 32'hc4044c0;
      2783: inst = 32'h8220000;
      2784: inst = 32'h10408000;
      2785: inst = 32'hc4044c1;
      2786: inst = 32'h8220000;
      2787: inst = 32'h10408000;
      2788: inst = 32'hc4044c2;
      2789: inst = 32'h8220000;
      2790: inst = 32'h10408000;
      2791: inst = 32'hc4044c3;
      2792: inst = 32'h8220000;
      2793: inst = 32'h10408000;
      2794: inst = 32'hc4044c4;
      2795: inst = 32'h8220000;
      2796: inst = 32'h10408000;
      2797: inst = 32'hc4044c5;
      2798: inst = 32'h8220000;
      2799: inst = 32'h10408000;
      2800: inst = 32'hc4044c6;
      2801: inst = 32'h8220000;
      2802: inst = 32'h10408000;
      2803: inst = 32'hc4044c7;
      2804: inst = 32'h8220000;
      2805: inst = 32'h10408000;
      2806: inst = 32'hc4044c8;
      2807: inst = 32'h8220000;
      2808: inst = 32'h10408000;
      2809: inst = 32'hc4044c9;
      2810: inst = 32'h8220000;
      2811: inst = 32'h10408000;
      2812: inst = 32'hc4044ca;
      2813: inst = 32'h8220000;
      2814: inst = 32'h10408000;
      2815: inst = 32'hc4044cd;
      2816: inst = 32'h8220000;
      2817: inst = 32'h10408000;
      2818: inst = 32'hc4044ce;
      2819: inst = 32'h8220000;
      2820: inst = 32'h10408000;
      2821: inst = 32'hc4044cf;
      2822: inst = 32'h8220000;
      2823: inst = 32'h10408000;
      2824: inst = 32'hc4044d0;
      2825: inst = 32'h8220000;
      2826: inst = 32'h10408000;
      2827: inst = 32'hc4044d1;
      2828: inst = 32'h8220000;
      2829: inst = 32'h10408000;
      2830: inst = 32'hc4044d2;
      2831: inst = 32'h8220000;
      2832: inst = 32'h10408000;
      2833: inst = 32'hc4044d3;
      2834: inst = 32'h8220000;
      2835: inst = 32'h10408000;
      2836: inst = 32'hc4044d4;
      2837: inst = 32'h8220000;
      2838: inst = 32'h10408000;
      2839: inst = 32'hc4044d5;
      2840: inst = 32'h8220000;
      2841: inst = 32'h10408000;
      2842: inst = 32'hc4044d6;
      2843: inst = 32'h8220000;
      2844: inst = 32'h10408000;
      2845: inst = 32'hc4044d7;
      2846: inst = 32'h8220000;
      2847: inst = 32'h10408000;
      2848: inst = 32'hc4044d8;
      2849: inst = 32'h8220000;
      2850: inst = 32'h10408000;
      2851: inst = 32'hc4044d9;
      2852: inst = 32'h8220000;
      2853: inst = 32'h10408000;
      2854: inst = 32'hc4044da;
      2855: inst = 32'h8220000;
      2856: inst = 32'h10408000;
      2857: inst = 32'hc4044db;
      2858: inst = 32'h8220000;
      2859: inst = 32'h10408000;
      2860: inst = 32'hc404504;
      2861: inst = 32'h8220000;
      2862: inst = 32'h10408000;
      2863: inst = 32'hc404505;
      2864: inst = 32'h8220000;
      2865: inst = 32'h10408000;
      2866: inst = 32'hc404506;
      2867: inst = 32'h8220000;
      2868: inst = 32'h10408000;
      2869: inst = 32'hc404507;
      2870: inst = 32'h8220000;
      2871: inst = 32'h10408000;
      2872: inst = 32'hc404508;
      2873: inst = 32'h8220000;
      2874: inst = 32'h10408000;
      2875: inst = 32'hc404509;
      2876: inst = 32'h8220000;
      2877: inst = 32'h10408000;
      2878: inst = 32'hc40450a;
      2879: inst = 32'h8220000;
      2880: inst = 32'h10408000;
      2881: inst = 32'hc40450b;
      2882: inst = 32'h8220000;
      2883: inst = 32'h10408000;
      2884: inst = 32'hc40450c;
      2885: inst = 32'h8220000;
      2886: inst = 32'h10408000;
      2887: inst = 32'hc40450d;
      2888: inst = 32'h8220000;
      2889: inst = 32'h10408000;
      2890: inst = 32'hc40450e;
      2891: inst = 32'h8220000;
      2892: inst = 32'h10408000;
      2893: inst = 32'hc40450f;
      2894: inst = 32'h8220000;
      2895: inst = 32'h10408000;
      2896: inst = 32'hc404510;
      2897: inst = 32'h8220000;
      2898: inst = 32'h10408000;
      2899: inst = 32'hc404511;
      2900: inst = 32'h8220000;
      2901: inst = 32'h10408000;
      2902: inst = 32'hc404512;
      2903: inst = 32'h8220000;
      2904: inst = 32'h10408000;
      2905: inst = 32'hc404515;
      2906: inst = 32'h8220000;
      2907: inst = 32'h10408000;
      2908: inst = 32'hc404516;
      2909: inst = 32'h8220000;
      2910: inst = 32'h10408000;
      2911: inst = 32'hc404517;
      2912: inst = 32'h8220000;
      2913: inst = 32'h10408000;
      2914: inst = 32'hc404518;
      2915: inst = 32'h8220000;
      2916: inst = 32'h10408000;
      2917: inst = 32'hc404519;
      2918: inst = 32'h8220000;
      2919: inst = 32'h10408000;
      2920: inst = 32'hc40451a;
      2921: inst = 32'h8220000;
      2922: inst = 32'h10408000;
      2923: inst = 32'hc40451b;
      2924: inst = 32'h8220000;
      2925: inst = 32'h10408000;
      2926: inst = 32'hc40451c;
      2927: inst = 32'h8220000;
      2928: inst = 32'h10408000;
      2929: inst = 32'hc40451d;
      2930: inst = 32'h8220000;
      2931: inst = 32'h10408000;
      2932: inst = 32'hc40451e;
      2933: inst = 32'h8220000;
      2934: inst = 32'h10408000;
      2935: inst = 32'hc40451f;
      2936: inst = 32'h8220000;
      2937: inst = 32'h10408000;
      2938: inst = 32'hc404520;
      2939: inst = 32'h8220000;
      2940: inst = 32'h10408000;
      2941: inst = 32'hc404521;
      2942: inst = 32'h8220000;
      2943: inst = 32'h10408000;
      2944: inst = 32'hc404522;
      2945: inst = 32'h8220000;
      2946: inst = 32'h10408000;
      2947: inst = 32'hc404523;
      2948: inst = 32'h8220000;
      2949: inst = 32'h10408000;
      2950: inst = 32'hc404524;
      2951: inst = 32'h8220000;
      2952: inst = 32'h10408000;
      2953: inst = 32'hc404525;
      2954: inst = 32'h8220000;
      2955: inst = 32'h10408000;
      2956: inst = 32'hc404526;
      2957: inst = 32'h8220000;
      2958: inst = 32'h10408000;
      2959: inst = 32'hc404527;
      2960: inst = 32'h8220000;
      2961: inst = 32'h10408000;
      2962: inst = 32'hc404528;
      2963: inst = 32'h8220000;
      2964: inst = 32'h10408000;
      2965: inst = 32'hc404529;
      2966: inst = 32'h8220000;
      2967: inst = 32'h10408000;
      2968: inst = 32'hc40452a;
      2969: inst = 32'h8220000;
      2970: inst = 32'h10408000;
      2971: inst = 32'hc40452b;
      2972: inst = 32'h8220000;
      2973: inst = 32'h10408000;
      2974: inst = 32'hc40452c;
      2975: inst = 32'h8220000;
      2976: inst = 32'h10408000;
      2977: inst = 32'hc40452d;
      2978: inst = 32'h8220000;
      2979: inst = 32'h10408000;
      2980: inst = 32'hc40452e;
      2981: inst = 32'h8220000;
      2982: inst = 32'h10408000;
      2983: inst = 32'hc40452f;
      2984: inst = 32'h8220000;
      2985: inst = 32'h10408000;
      2986: inst = 32'hc404530;
      2987: inst = 32'h8220000;
      2988: inst = 32'h10408000;
      2989: inst = 32'hc404531;
      2990: inst = 32'h8220000;
      2991: inst = 32'h10408000;
      2992: inst = 32'hc404532;
      2993: inst = 32'h8220000;
      2994: inst = 32'h10408000;
      2995: inst = 32'hc404533;
      2996: inst = 32'h8220000;
      2997: inst = 32'h10408000;
      2998: inst = 32'hc404534;
      2999: inst = 32'h8220000;
      3000: inst = 32'h10408000;
      3001: inst = 32'hc404535;
      3002: inst = 32'h8220000;
      3003: inst = 32'h10408000;
      3004: inst = 32'hc404536;
      3005: inst = 32'h8220000;
      3006: inst = 32'h10408000;
      3007: inst = 32'hc404537;
      3008: inst = 32'h8220000;
      3009: inst = 32'h10408000;
      3010: inst = 32'hc404538;
      3011: inst = 32'h8220000;
      3012: inst = 32'h10408000;
      3013: inst = 32'hc404539;
      3014: inst = 32'h8220000;
      3015: inst = 32'h10408000;
      3016: inst = 32'hc40453a;
      3017: inst = 32'h8220000;
      3018: inst = 32'h10408000;
      3019: inst = 32'hc40453b;
      3020: inst = 32'h8220000;
      3021: inst = 32'h10408000;
      3022: inst = 32'hc404564;
      3023: inst = 32'h8220000;
      3024: inst = 32'h10408000;
      3025: inst = 32'hc404565;
      3026: inst = 32'h8220000;
      3027: inst = 32'h10408000;
      3028: inst = 32'hc404566;
      3029: inst = 32'h8220000;
      3030: inst = 32'h10408000;
      3031: inst = 32'hc404567;
      3032: inst = 32'h8220000;
      3033: inst = 32'h10408000;
      3034: inst = 32'hc404568;
      3035: inst = 32'h8220000;
      3036: inst = 32'h10408000;
      3037: inst = 32'hc404569;
      3038: inst = 32'h8220000;
      3039: inst = 32'h10408000;
      3040: inst = 32'hc40456a;
      3041: inst = 32'h8220000;
      3042: inst = 32'h10408000;
      3043: inst = 32'hc40456b;
      3044: inst = 32'h8220000;
      3045: inst = 32'h10408000;
      3046: inst = 32'hc40456c;
      3047: inst = 32'h8220000;
      3048: inst = 32'h10408000;
      3049: inst = 32'hc40456d;
      3050: inst = 32'h8220000;
      3051: inst = 32'h10408000;
      3052: inst = 32'hc40456e;
      3053: inst = 32'h8220000;
      3054: inst = 32'h10408000;
      3055: inst = 32'hc40456f;
      3056: inst = 32'h8220000;
      3057: inst = 32'h10408000;
      3058: inst = 32'hc404570;
      3059: inst = 32'h8220000;
      3060: inst = 32'h10408000;
      3061: inst = 32'hc404571;
      3062: inst = 32'h8220000;
      3063: inst = 32'h10408000;
      3064: inst = 32'hc404572;
      3065: inst = 32'h8220000;
      3066: inst = 32'h10408000;
      3067: inst = 32'hc404573;
      3068: inst = 32'h8220000;
      3069: inst = 32'h10408000;
      3070: inst = 32'hc404574;
      3071: inst = 32'h8220000;
      3072: inst = 32'h10408000;
      3073: inst = 32'hc404575;
      3074: inst = 32'h8220000;
      3075: inst = 32'h10408000;
      3076: inst = 32'hc404576;
      3077: inst = 32'h8220000;
      3078: inst = 32'h10408000;
      3079: inst = 32'hc404577;
      3080: inst = 32'h8220000;
      3081: inst = 32'h10408000;
      3082: inst = 32'hc404578;
      3083: inst = 32'h8220000;
      3084: inst = 32'h10408000;
      3085: inst = 32'hc404579;
      3086: inst = 32'h8220000;
      3087: inst = 32'h10408000;
      3088: inst = 32'hc40457a;
      3089: inst = 32'h8220000;
      3090: inst = 32'h10408000;
      3091: inst = 32'hc40457b;
      3092: inst = 32'h8220000;
      3093: inst = 32'h10408000;
      3094: inst = 32'hc40457c;
      3095: inst = 32'h8220000;
      3096: inst = 32'h10408000;
      3097: inst = 32'hc40457d;
      3098: inst = 32'h8220000;
      3099: inst = 32'h10408000;
      3100: inst = 32'hc40457e;
      3101: inst = 32'h8220000;
      3102: inst = 32'h10408000;
      3103: inst = 32'hc40457f;
      3104: inst = 32'h8220000;
      3105: inst = 32'h10408000;
      3106: inst = 32'hc404580;
      3107: inst = 32'h8220000;
      3108: inst = 32'h10408000;
      3109: inst = 32'hc404581;
      3110: inst = 32'h8220000;
      3111: inst = 32'h10408000;
      3112: inst = 32'hc404582;
      3113: inst = 32'h8220000;
      3114: inst = 32'h10408000;
      3115: inst = 32'hc404583;
      3116: inst = 32'h8220000;
      3117: inst = 32'h10408000;
      3118: inst = 32'hc404584;
      3119: inst = 32'h8220000;
      3120: inst = 32'h10408000;
      3121: inst = 32'hc404585;
      3122: inst = 32'h8220000;
      3123: inst = 32'h10408000;
      3124: inst = 32'hc404586;
      3125: inst = 32'h8220000;
      3126: inst = 32'h10408000;
      3127: inst = 32'hc404587;
      3128: inst = 32'h8220000;
      3129: inst = 32'h10408000;
      3130: inst = 32'hc404588;
      3131: inst = 32'h8220000;
      3132: inst = 32'h10408000;
      3133: inst = 32'hc404589;
      3134: inst = 32'h8220000;
      3135: inst = 32'h10408000;
      3136: inst = 32'hc40458a;
      3137: inst = 32'h8220000;
      3138: inst = 32'h10408000;
      3139: inst = 32'hc40458b;
      3140: inst = 32'h8220000;
      3141: inst = 32'h10408000;
      3142: inst = 32'hc40458c;
      3143: inst = 32'h8220000;
      3144: inst = 32'h10408000;
      3145: inst = 32'hc40458d;
      3146: inst = 32'h8220000;
      3147: inst = 32'h10408000;
      3148: inst = 32'hc40458e;
      3149: inst = 32'h8220000;
      3150: inst = 32'h10408000;
      3151: inst = 32'hc40458f;
      3152: inst = 32'h8220000;
      3153: inst = 32'h10408000;
      3154: inst = 32'hc404590;
      3155: inst = 32'h8220000;
      3156: inst = 32'h10408000;
      3157: inst = 32'hc404591;
      3158: inst = 32'h8220000;
      3159: inst = 32'h10408000;
      3160: inst = 32'hc404592;
      3161: inst = 32'h8220000;
      3162: inst = 32'h10408000;
      3163: inst = 32'hc404593;
      3164: inst = 32'h8220000;
      3165: inst = 32'h10408000;
      3166: inst = 32'hc404594;
      3167: inst = 32'h8220000;
      3168: inst = 32'h10408000;
      3169: inst = 32'hc404595;
      3170: inst = 32'h8220000;
      3171: inst = 32'h10408000;
      3172: inst = 32'hc404596;
      3173: inst = 32'h8220000;
      3174: inst = 32'h10408000;
      3175: inst = 32'hc404597;
      3176: inst = 32'h8220000;
      3177: inst = 32'h10408000;
      3178: inst = 32'hc404598;
      3179: inst = 32'h8220000;
      3180: inst = 32'h10408000;
      3181: inst = 32'hc404599;
      3182: inst = 32'h8220000;
      3183: inst = 32'h10408000;
      3184: inst = 32'hc40459a;
      3185: inst = 32'h8220000;
      3186: inst = 32'h10408000;
      3187: inst = 32'hc40459b;
      3188: inst = 32'h8220000;
      3189: inst = 32'h10408000;
      3190: inst = 32'hc4045c4;
      3191: inst = 32'h8220000;
      3192: inst = 32'h10408000;
      3193: inst = 32'hc4045c5;
      3194: inst = 32'h8220000;
      3195: inst = 32'h10408000;
      3196: inst = 32'hc4045c6;
      3197: inst = 32'h8220000;
      3198: inst = 32'h10408000;
      3199: inst = 32'hc4045c7;
      3200: inst = 32'h8220000;
      3201: inst = 32'h10408000;
      3202: inst = 32'hc4045c8;
      3203: inst = 32'h8220000;
      3204: inst = 32'h10408000;
      3205: inst = 32'hc4045c9;
      3206: inst = 32'h8220000;
      3207: inst = 32'h10408000;
      3208: inst = 32'hc4045ca;
      3209: inst = 32'h8220000;
      3210: inst = 32'h10408000;
      3211: inst = 32'hc4045cb;
      3212: inst = 32'h8220000;
      3213: inst = 32'h10408000;
      3214: inst = 32'hc4045cc;
      3215: inst = 32'h8220000;
      3216: inst = 32'h10408000;
      3217: inst = 32'hc4045cd;
      3218: inst = 32'h8220000;
      3219: inst = 32'h10408000;
      3220: inst = 32'hc4045ce;
      3221: inst = 32'h8220000;
      3222: inst = 32'h10408000;
      3223: inst = 32'hc4045cf;
      3224: inst = 32'h8220000;
      3225: inst = 32'h10408000;
      3226: inst = 32'hc4045d0;
      3227: inst = 32'h8220000;
      3228: inst = 32'h10408000;
      3229: inst = 32'hc4045d1;
      3230: inst = 32'h8220000;
      3231: inst = 32'h10408000;
      3232: inst = 32'hc4045d2;
      3233: inst = 32'h8220000;
      3234: inst = 32'h10408000;
      3235: inst = 32'hc4045d3;
      3236: inst = 32'h8220000;
      3237: inst = 32'h10408000;
      3238: inst = 32'hc4045d4;
      3239: inst = 32'h8220000;
      3240: inst = 32'h10408000;
      3241: inst = 32'hc4045d5;
      3242: inst = 32'h8220000;
      3243: inst = 32'h10408000;
      3244: inst = 32'hc4045d6;
      3245: inst = 32'h8220000;
      3246: inst = 32'h10408000;
      3247: inst = 32'hc4045d7;
      3248: inst = 32'h8220000;
      3249: inst = 32'h10408000;
      3250: inst = 32'hc4045d8;
      3251: inst = 32'h8220000;
      3252: inst = 32'h10408000;
      3253: inst = 32'hc4045d9;
      3254: inst = 32'h8220000;
      3255: inst = 32'h10408000;
      3256: inst = 32'hc4045da;
      3257: inst = 32'h8220000;
      3258: inst = 32'h10408000;
      3259: inst = 32'hc4045db;
      3260: inst = 32'h8220000;
      3261: inst = 32'h10408000;
      3262: inst = 32'hc4045dc;
      3263: inst = 32'h8220000;
      3264: inst = 32'h10408000;
      3265: inst = 32'hc4045dd;
      3266: inst = 32'h8220000;
      3267: inst = 32'h10408000;
      3268: inst = 32'hc4045de;
      3269: inst = 32'h8220000;
      3270: inst = 32'h10408000;
      3271: inst = 32'hc4045df;
      3272: inst = 32'h8220000;
      3273: inst = 32'h10408000;
      3274: inst = 32'hc4045e0;
      3275: inst = 32'h8220000;
      3276: inst = 32'h10408000;
      3277: inst = 32'hc4045e1;
      3278: inst = 32'h8220000;
      3279: inst = 32'h10408000;
      3280: inst = 32'hc4045e2;
      3281: inst = 32'h8220000;
      3282: inst = 32'h10408000;
      3283: inst = 32'hc4045e3;
      3284: inst = 32'h8220000;
      3285: inst = 32'h10408000;
      3286: inst = 32'hc4045e4;
      3287: inst = 32'h8220000;
      3288: inst = 32'h10408000;
      3289: inst = 32'hc4045e5;
      3290: inst = 32'h8220000;
      3291: inst = 32'h10408000;
      3292: inst = 32'hc4045e6;
      3293: inst = 32'h8220000;
      3294: inst = 32'h10408000;
      3295: inst = 32'hc4045e7;
      3296: inst = 32'h8220000;
      3297: inst = 32'h10408000;
      3298: inst = 32'hc4045e8;
      3299: inst = 32'h8220000;
      3300: inst = 32'h10408000;
      3301: inst = 32'hc4045e9;
      3302: inst = 32'h8220000;
      3303: inst = 32'h10408000;
      3304: inst = 32'hc4045ea;
      3305: inst = 32'h8220000;
      3306: inst = 32'h10408000;
      3307: inst = 32'hc4045eb;
      3308: inst = 32'h8220000;
      3309: inst = 32'h10408000;
      3310: inst = 32'hc4045ec;
      3311: inst = 32'h8220000;
      3312: inst = 32'h10408000;
      3313: inst = 32'hc4045ed;
      3314: inst = 32'h8220000;
      3315: inst = 32'h10408000;
      3316: inst = 32'hc4045ee;
      3317: inst = 32'h8220000;
      3318: inst = 32'h10408000;
      3319: inst = 32'hc4045ef;
      3320: inst = 32'h8220000;
      3321: inst = 32'h10408000;
      3322: inst = 32'hc4045f0;
      3323: inst = 32'h8220000;
      3324: inst = 32'h10408000;
      3325: inst = 32'hc4045f1;
      3326: inst = 32'h8220000;
      3327: inst = 32'h10408000;
      3328: inst = 32'hc4045f2;
      3329: inst = 32'h8220000;
      3330: inst = 32'h10408000;
      3331: inst = 32'hc4045f3;
      3332: inst = 32'h8220000;
      3333: inst = 32'h10408000;
      3334: inst = 32'hc4045f4;
      3335: inst = 32'h8220000;
      3336: inst = 32'h10408000;
      3337: inst = 32'hc4045f5;
      3338: inst = 32'h8220000;
      3339: inst = 32'h10408000;
      3340: inst = 32'hc4045f6;
      3341: inst = 32'h8220000;
      3342: inst = 32'h10408000;
      3343: inst = 32'hc4045f7;
      3344: inst = 32'h8220000;
      3345: inst = 32'h10408000;
      3346: inst = 32'hc4045f8;
      3347: inst = 32'h8220000;
      3348: inst = 32'h10408000;
      3349: inst = 32'hc4045f9;
      3350: inst = 32'h8220000;
      3351: inst = 32'h10408000;
      3352: inst = 32'hc4045fa;
      3353: inst = 32'h8220000;
      3354: inst = 32'h10408000;
      3355: inst = 32'hc4045fb;
      3356: inst = 32'h8220000;
      3357: inst = 32'h10408000;
      3358: inst = 32'hc404624;
      3359: inst = 32'h8220000;
      3360: inst = 32'h10408000;
      3361: inst = 32'hc404625;
      3362: inst = 32'h8220000;
      3363: inst = 32'h10408000;
      3364: inst = 32'hc404626;
      3365: inst = 32'h8220000;
      3366: inst = 32'h10408000;
      3367: inst = 32'hc404627;
      3368: inst = 32'h8220000;
      3369: inst = 32'h10408000;
      3370: inst = 32'hc404628;
      3371: inst = 32'h8220000;
      3372: inst = 32'h10408000;
      3373: inst = 32'hc404629;
      3374: inst = 32'h8220000;
      3375: inst = 32'h10408000;
      3376: inst = 32'hc40462a;
      3377: inst = 32'h8220000;
      3378: inst = 32'h10408000;
      3379: inst = 32'hc40462b;
      3380: inst = 32'h8220000;
      3381: inst = 32'h10408000;
      3382: inst = 32'hc40462c;
      3383: inst = 32'h8220000;
      3384: inst = 32'h10408000;
      3385: inst = 32'hc40462d;
      3386: inst = 32'h8220000;
      3387: inst = 32'h10408000;
      3388: inst = 32'hc40462e;
      3389: inst = 32'h8220000;
      3390: inst = 32'h10408000;
      3391: inst = 32'hc40462f;
      3392: inst = 32'h8220000;
      3393: inst = 32'h10408000;
      3394: inst = 32'hc404630;
      3395: inst = 32'h8220000;
      3396: inst = 32'h10408000;
      3397: inst = 32'hc404631;
      3398: inst = 32'h8220000;
      3399: inst = 32'h10408000;
      3400: inst = 32'hc404632;
      3401: inst = 32'h8220000;
      3402: inst = 32'h10408000;
      3403: inst = 32'hc404633;
      3404: inst = 32'h8220000;
      3405: inst = 32'h10408000;
      3406: inst = 32'hc404634;
      3407: inst = 32'h8220000;
      3408: inst = 32'h10408000;
      3409: inst = 32'hc404635;
      3410: inst = 32'h8220000;
      3411: inst = 32'h10408000;
      3412: inst = 32'hc404636;
      3413: inst = 32'h8220000;
      3414: inst = 32'h10408000;
      3415: inst = 32'hc404637;
      3416: inst = 32'h8220000;
      3417: inst = 32'h10408000;
      3418: inst = 32'hc404638;
      3419: inst = 32'h8220000;
      3420: inst = 32'h10408000;
      3421: inst = 32'hc404639;
      3422: inst = 32'h8220000;
      3423: inst = 32'h10408000;
      3424: inst = 32'hc40463a;
      3425: inst = 32'h8220000;
      3426: inst = 32'h10408000;
      3427: inst = 32'hc40463b;
      3428: inst = 32'h8220000;
      3429: inst = 32'h10408000;
      3430: inst = 32'hc40463c;
      3431: inst = 32'h8220000;
      3432: inst = 32'h10408000;
      3433: inst = 32'hc40463d;
      3434: inst = 32'h8220000;
      3435: inst = 32'h10408000;
      3436: inst = 32'hc40463e;
      3437: inst = 32'h8220000;
      3438: inst = 32'h10408000;
      3439: inst = 32'hc40463f;
      3440: inst = 32'h8220000;
      3441: inst = 32'h10408000;
      3442: inst = 32'hc404640;
      3443: inst = 32'h8220000;
      3444: inst = 32'h10408000;
      3445: inst = 32'hc404641;
      3446: inst = 32'h8220000;
      3447: inst = 32'h10408000;
      3448: inst = 32'hc404642;
      3449: inst = 32'h8220000;
      3450: inst = 32'h10408000;
      3451: inst = 32'hc404643;
      3452: inst = 32'h8220000;
      3453: inst = 32'h10408000;
      3454: inst = 32'hc404644;
      3455: inst = 32'h8220000;
      3456: inst = 32'h10408000;
      3457: inst = 32'hc404645;
      3458: inst = 32'h8220000;
      3459: inst = 32'h10408000;
      3460: inst = 32'hc404646;
      3461: inst = 32'h8220000;
      3462: inst = 32'h10408000;
      3463: inst = 32'hc404647;
      3464: inst = 32'h8220000;
      3465: inst = 32'h10408000;
      3466: inst = 32'hc404648;
      3467: inst = 32'h8220000;
      3468: inst = 32'h10408000;
      3469: inst = 32'hc404649;
      3470: inst = 32'h8220000;
      3471: inst = 32'h10408000;
      3472: inst = 32'hc40464a;
      3473: inst = 32'h8220000;
      3474: inst = 32'h10408000;
      3475: inst = 32'hc40464b;
      3476: inst = 32'h8220000;
      3477: inst = 32'h10408000;
      3478: inst = 32'hc40464c;
      3479: inst = 32'h8220000;
      3480: inst = 32'h10408000;
      3481: inst = 32'hc40464d;
      3482: inst = 32'h8220000;
      3483: inst = 32'h10408000;
      3484: inst = 32'hc40464e;
      3485: inst = 32'h8220000;
      3486: inst = 32'h10408000;
      3487: inst = 32'hc40464f;
      3488: inst = 32'h8220000;
      3489: inst = 32'h10408000;
      3490: inst = 32'hc404650;
      3491: inst = 32'h8220000;
      3492: inst = 32'h10408000;
      3493: inst = 32'hc404651;
      3494: inst = 32'h8220000;
      3495: inst = 32'h10408000;
      3496: inst = 32'hc404652;
      3497: inst = 32'h8220000;
      3498: inst = 32'h10408000;
      3499: inst = 32'hc404653;
      3500: inst = 32'h8220000;
      3501: inst = 32'h10408000;
      3502: inst = 32'hc404654;
      3503: inst = 32'h8220000;
      3504: inst = 32'h10408000;
      3505: inst = 32'hc404655;
      3506: inst = 32'h8220000;
      3507: inst = 32'h10408000;
      3508: inst = 32'hc404656;
      3509: inst = 32'h8220000;
      3510: inst = 32'h10408000;
      3511: inst = 32'hc404657;
      3512: inst = 32'h8220000;
      3513: inst = 32'h10408000;
      3514: inst = 32'hc404658;
      3515: inst = 32'h8220000;
      3516: inst = 32'h10408000;
      3517: inst = 32'hc404659;
      3518: inst = 32'h8220000;
      3519: inst = 32'h10408000;
      3520: inst = 32'hc40465a;
      3521: inst = 32'h8220000;
      3522: inst = 32'h10408000;
      3523: inst = 32'hc40465b;
      3524: inst = 32'h8220000;
      3525: inst = 32'h10408000;
      3526: inst = 32'hc404684;
      3527: inst = 32'h8220000;
      3528: inst = 32'h10408000;
      3529: inst = 32'hc404685;
      3530: inst = 32'h8220000;
      3531: inst = 32'h10408000;
      3532: inst = 32'hc404686;
      3533: inst = 32'h8220000;
      3534: inst = 32'h10408000;
      3535: inst = 32'hc404687;
      3536: inst = 32'h8220000;
      3537: inst = 32'h10408000;
      3538: inst = 32'hc404688;
      3539: inst = 32'h8220000;
      3540: inst = 32'h10408000;
      3541: inst = 32'hc404689;
      3542: inst = 32'h8220000;
      3543: inst = 32'h10408000;
      3544: inst = 32'hc40468a;
      3545: inst = 32'h8220000;
      3546: inst = 32'h10408000;
      3547: inst = 32'hc40468b;
      3548: inst = 32'h8220000;
      3549: inst = 32'h10408000;
      3550: inst = 32'hc40468c;
      3551: inst = 32'h8220000;
      3552: inst = 32'h10408000;
      3553: inst = 32'hc40468d;
      3554: inst = 32'h8220000;
      3555: inst = 32'h10408000;
      3556: inst = 32'hc40468e;
      3557: inst = 32'h8220000;
      3558: inst = 32'h10408000;
      3559: inst = 32'hc40468f;
      3560: inst = 32'h8220000;
      3561: inst = 32'h10408000;
      3562: inst = 32'hc404690;
      3563: inst = 32'h8220000;
      3564: inst = 32'h10408000;
      3565: inst = 32'hc404691;
      3566: inst = 32'h8220000;
      3567: inst = 32'h10408000;
      3568: inst = 32'hc404692;
      3569: inst = 32'h8220000;
      3570: inst = 32'h10408000;
      3571: inst = 32'hc404693;
      3572: inst = 32'h8220000;
      3573: inst = 32'h10408000;
      3574: inst = 32'hc404694;
      3575: inst = 32'h8220000;
      3576: inst = 32'h10408000;
      3577: inst = 32'hc404695;
      3578: inst = 32'h8220000;
      3579: inst = 32'h10408000;
      3580: inst = 32'hc404696;
      3581: inst = 32'h8220000;
      3582: inst = 32'h10408000;
      3583: inst = 32'hc404697;
      3584: inst = 32'h8220000;
      3585: inst = 32'h10408000;
      3586: inst = 32'hc404698;
      3587: inst = 32'h8220000;
      3588: inst = 32'h10408000;
      3589: inst = 32'hc404699;
      3590: inst = 32'h8220000;
      3591: inst = 32'h10408000;
      3592: inst = 32'hc40469a;
      3593: inst = 32'h8220000;
      3594: inst = 32'h10408000;
      3595: inst = 32'hc40469b;
      3596: inst = 32'h8220000;
      3597: inst = 32'h10408000;
      3598: inst = 32'hc40469c;
      3599: inst = 32'h8220000;
      3600: inst = 32'h10408000;
      3601: inst = 32'hc40469d;
      3602: inst = 32'h8220000;
      3603: inst = 32'h10408000;
      3604: inst = 32'hc40469e;
      3605: inst = 32'h8220000;
      3606: inst = 32'h10408000;
      3607: inst = 32'hc40469f;
      3608: inst = 32'h8220000;
      3609: inst = 32'h10408000;
      3610: inst = 32'hc4046a0;
      3611: inst = 32'h8220000;
      3612: inst = 32'h10408000;
      3613: inst = 32'hc4046a1;
      3614: inst = 32'h8220000;
      3615: inst = 32'h10408000;
      3616: inst = 32'hc4046a2;
      3617: inst = 32'h8220000;
      3618: inst = 32'h10408000;
      3619: inst = 32'hc4046a3;
      3620: inst = 32'h8220000;
      3621: inst = 32'h10408000;
      3622: inst = 32'hc4046a4;
      3623: inst = 32'h8220000;
      3624: inst = 32'h10408000;
      3625: inst = 32'hc4046a5;
      3626: inst = 32'h8220000;
      3627: inst = 32'h10408000;
      3628: inst = 32'hc4046a6;
      3629: inst = 32'h8220000;
      3630: inst = 32'h10408000;
      3631: inst = 32'hc4046a7;
      3632: inst = 32'h8220000;
      3633: inst = 32'h10408000;
      3634: inst = 32'hc4046a8;
      3635: inst = 32'h8220000;
      3636: inst = 32'h10408000;
      3637: inst = 32'hc4046a9;
      3638: inst = 32'h8220000;
      3639: inst = 32'h10408000;
      3640: inst = 32'hc4046aa;
      3641: inst = 32'h8220000;
      3642: inst = 32'h10408000;
      3643: inst = 32'hc4046ab;
      3644: inst = 32'h8220000;
      3645: inst = 32'h10408000;
      3646: inst = 32'hc4046ac;
      3647: inst = 32'h8220000;
      3648: inst = 32'h10408000;
      3649: inst = 32'hc4046ad;
      3650: inst = 32'h8220000;
      3651: inst = 32'h10408000;
      3652: inst = 32'hc4046ae;
      3653: inst = 32'h8220000;
      3654: inst = 32'h10408000;
      3655: inst = 32'hc4046af;
      3656: inst = 32'h8220000;
      3657: inst = 32'h10408000;
      3658: inst = 32'hc4046b0;
      3659: inst = 32'h8220000;
      3660: inst = 32'h10408000;
      3661: inst = 32'hc4046b1;
      3662: inst = 32'h8220000;
      3663: inst = 32'h10408000;
      3664: inst = 32'hc4046b2;
      3665: inst = 32'h8220000;
      3666: inst = 32'h10408000;
      3667: inst = 32'hc4046b3;
      3668: inst = 32'h8220000;
      3669: inst = 32'h10408000;
      3670: inst = 32'hc4046b4;
      3671: inst = 32'h8220000;
      3672: inst = 32'h10408000;
      3673: inst = 32'hc4046b5;
      3674: inst = 32'h8220000;
      3675: inst = 32'h10408000;
      3676: inst = 32'hc4046b6;
      3677: inst = 32'h8220000;
      3678: inst = 32'h10408000;
      3679: inst = 32'hc4046b7;
      3680: inst = 32'h8220000;
      3681: inst = 32'h10408000;
      3682: inst = 32'hc4046b8;
      3683: inst = 32'h8220000;
      3684: inst = 32'h10408000;
      3685: inst = 32'hc4046b9;
      3686: inst = 32'h8220000;
      3687: inst = 32'h10408000;
      3688: inst = 32'hc4046ba;
      3689: inst = 32'h8220000;
      3690: inst = 32'h10408000;
      3691: inst = 32'hc4046bb;
      3692: inst = 32'h8220000;
      3693: inst = 32'h10408000;
      3694: inst = 32'hc4046e4;
      3695: inst = 32'h8220000;
      3696: inst = 32'h10408000;
      3697: inst = 32'hc4046e5;
      3698: inst = 32'h8220000;
      3699: inst = 32'h10408000;
      3700: inst = 32'hc4046e6;
      3701: inst = 32'h8220000;
      3702: inst = 32'h10408000;
      3703: inst = 32'hc4046e7;
      3704: inst = 32'h8220000;
      3705: inst = 32'h10408000;
      3706: inst = 32'hc4046e8;
      3707: inst = 32'h8220000;
      3708: inst = 32'h10408000;
      3709: inst = 32'hc4046e9;
      3710: inst = 32'h8220000;
      3711: inst = 32'h10408000;
      3712: inst = 32'hc4046ea;
      3713: inst = 32'h8220000;
      3714: inst = 32'h10408000;
      3715: inst = 32'hc4046eb;
      3716: inst = 32'h8220000;
      3717: inst = 32'h10408000;
      3718: inst = 32'hc4046ec;
      3719: inst = 32'h8220000;
      3720: inst = 32'h10408000;
      3721: inst = 32'hc4046ed;
      3722: inst = 32'h8220000;
      3723: inst = 32'h10408000;
      3724: inst = 32'hc4046ee;
      3725: inst = 32'h8220000;
      3726: inst = 32'h10408000;
      3727: inst = 32'hc404700;
      3728: inst = 32'h8220000;
      3729: inst = 32'h10408000;
      3730: inst = 32'hc404701;
      3731: inst = 32'h8220000;
      3732: inst = 32'h10408000;
      3733: inst = 32'hc404702;
      3734: inst = 32'h8220000;
      3735: inst = 32'h10408000;
      3736: inst = 32'hc404703;
      3737: inst = 32'h8220000;
      3738: inst = 32'h10408000;
      3739: inst = 32'hc404704;
      3740: inst = 32'h8220000;
      3741: inst = 32'h10408000;
      3742: inst = 32'hc404705;
      3743: inst = 32'h8220000;
      3744: inst = 32'h10408000;
      3745: inst = 32'hc404706;
      3746: inst = 32'h8220000;
      3747: inst = 32'h10408000;
      3748: inst = 32'hc404707;
      3749: inst = 32'h8220000;
      3750: inst = 32'h10408000;
      3751: inst = 32'hc404708;
      3752: inst = 32'h8220000;
      3753: inst = 32'h10408000;
      3754: inst = 32'hc404709;
      3755: inst = 32'h8220000;
      3756: inst = 32'h10408000;
      3757: inst = 32'hc40470a;
      3758: inst = 32'h8220000;
      3759: inst = 32'h10408000;
      3760: inst = 32'hc40470b;
      3761: inst = 32'h8220000;
      3762: inst = 32'h10408000;
      3763: inst = 32'hc40470c;
      3764: inst = 32'h8220000;
      3765: inst = 32'h10408000;
      3766: inst = 32'hc40470d;
      3767: inst = 32'h8220000;
      3768: inst = 32'h10408000;
      3769: inst = 32'hc40470e;
      3770: inst = 32'h8220000;
      3771: inst = 32'h10408000;
      3772: inst = 32'hc40470f;
      3773: inst = 32'h8220000;
      3774: inst = 32'h10408000;
      3775: inst = 32'hc404710;
      3776: inst = 32'h8220000;
      3777: inst = 32'h10408000;
      3778: inst = 32'hc404711;
      3779: inst = 32'h8220000;
      3780: inst = 32'h10408000;
      3781: inst = 32'hc404712;
      3782: inst = 32'h8220000;
      3783: inst = 32'h10408000;
      3784: inst = 32'hc404713;
      3785: inst = 32'h8220000;
      3786: inst = 32'h10408000;
      3787: inst = 32'hc404714;
      3788: inst = 32'h8220000;
      3789: inst = 32'h10408000;
      3790: inst = 32'hc404715;
      3791: inst = 32'h8220000;
      3792: inst = 32'h10408000;
      3793: inst = 32'hc404716;
      3794: inst = 32'h8220000;
      3795: inst = 32'h10408000;
      3796: inst = 32'hc404717;
      3797: inst = 32'h8220000;
      3798: inst = 32'h10408000;
      3799: inst = 32'hc404718;
      3800: inst = 32'h8220000;
      3801: inst = 32'h10408000;
      3802: inst = 32'hc404719;
      3803: inst = 32'h8220000;
      3804: inst = 32'h10408000;
      3805: inst = 32'hc40471a;
      3806: inst = 32'h8220000;
      3807: inst = 32'h10408000;
      3808: inst = 32'hc40471b;
      3809: inst = 32'h8220000;
      3810: inst = 32'h10408000;
      3811: inst = 32'hc404744;
      3812: inst = 32'h8220000;
      3813: inst = 32'h10408000;
      3814: inst = 32'hc404745;
      3815: inst = 32'h8220000;
      3816: inst = 32'h10408000;
      3817: inst = 32'hc404746;
      3818: inst = 32'h8220000;
      3819: inst = 32'h10408000;
      3820: inst = 32'hc404747;
      3821: inst = 32'h8220000;
      3822: inst = 32'h10408000;
      3823: inst = 32'hc404748;
      3824: inst = 32'h8220000;
      3825: inst = 32'h10408000;
      3826: inst = 32'hc404749;
      3827: inst = 32'h8220000;
      3828: inst = 32'h10408000;
      3829: inst = 32'hc40474a;
      3830: inst = 32'h8220000;
      3831: inst = 32'h10408000;
      3832: inst = 32'hc40474b;
      3833: inst = 32'h8220000;
      3834: inst = 32'h10408000;
      3835: inst = 32'hc40474c;
      3836: inst = 32'h8220000;
      3837: inst = 32'h10408000;
      3838: inst = 32'hc40474d;
      3839: inst = 32'h8220000;
      3840: inst = 32'h10408000;
      3841: inst = 32'hc40474e;
      3842: inst = 32'h8220000;
      3843: inst = 32'h10408000;
      3844: inst = 32'hc404760;
      3845: inst = 32'h8220000;
      3846: inst = 32'h10408000;
      3847: inst = 32'hc404761;
      3848: inst = 32'h8220000;
      3849: inst = 32'h10408000;
      3850: inst = 32'hc404762;
      3851: inst = 32'h8220000;
      3852: inst = 32'h10408000;
      3853: inst = 32'hc404763;
      3854: inst = 32'h8220000;
      3855: inst = 32'h10408000;
      3856: inst = 32'hc404764;
      3857: inst = 32'h8220000;
      3858: inst = 32'h10408000;
      3859: inst = 32'hc404765;
      3860: inst = 32'h8220000;
      3861: inst = 32'h10408000;
      3862: inst = 32'hc404766;
      3863: inst = 32'h8220000;
      3864: inst = 32'h10408000;
      3865: inst = 32'hc404767;
      3866: inst = 32'h8220000;
      3867: inst = 32'h10408000;
      3868: inst = 32'hc404768;
      3869: inst = 32'h8220000;
      3870: inst = 32'h10408000;
      3871: inst = 32'hc404769;
      3872: inst = 32'h8220000;
      3873: inst = 32'h10408000;
      3874: inst = 32'hc40476a;
      3875: inst = 32'h8220000;
      3876: inst = 32'h10408000;
      3877: inst = 32'hc40476b;
      3878: inst = 32'h8220000;
      3879: inst = 32'h10408000;
      3880: inst = 32'hc40476c;
      3881: inst = 32'h8220000;
      3882: inst = 32'h10408000;
      3883: inst = 32'hc40476d;
      3884: inst = 32'h8220000;
      3885: inst = 32'h10408000;
      3886: inst = 32'hc40476e;
      3887: inst = 32'h8220000;
      3888: inst = 32'h10408000;
      3889: inst = 32'hc40476f;
      3890: inst = 32'h8220000;
      3891: inst = 32'h10408000;
      3892: inst = 32'hc404770;
      3893: inst = 32'h8220000;
      3894: inst = 32'h10408000;
      3895: inst = 32'hc404771;
      3896: inst = 32'h8220000;
      3897: inst = 32'h10408000;
      3898: inst = 32'hc404772;
      3899: inst = 32'h8220000;
      3900: inst = 32'h10408000;
      3901: inst = 32'hc404773;
      3902: inst = 32'h8220000;
      3903: inst = 32'h10408000;
      3904: inst = 32'hc404774;
      3905: inst = 32'h8220000;
      3906: inst = 32'h10408000;
      3907: inst = 32'hc404775;
      3908: inst = 32'h8220000;
      3909: inst = 32'h10408000;
      3910: inst = 32'hc404776;
      3911: inst = 32'h8220000;
      3912: inst = 32'h10408000;
      3913: inst = 32'hc404777;
      3914: inst = 32'h8220000;
      3915: inst = 32'h10408000;
      3916: inst = 32'hc404778;
      3917: inst = 32'h8220000;
      3918: inst = 32'h10408000;
      3919: inst = 32'hc404779;
      3920: inst = 32'h8220000;
      3921: inst = 32'h10408000;
      3922: inst = 32'hc40477a;
      3923: inst = 32'h8220000;
      3924: inst = 32'h10408000;
      3925: inst = 32'hc40477b;
      3926: inst = 32'h8220000;
      3927: inst = 32'h10408000;
      3928: inst = 32'hc4047a4;
      3929: inst = 32'h8220000;
      3930: inst = 32'h10408000;
      3931: inst = 32'hc4047a5;
      3932: inst = 32'h8220000;
      3933: inst = 32'h10408000;
      3934: inst = 32'hc4047a6;
      3935: inst = 32'h8220000;
      3936: inst = 32'h10408000;
      3937: inst = 32'hc4047a7;
      3938: inst = 32'h8220000;
      3939: inst = 32'h10408000;
      3940: inst = 32'hc4047a8;
      3941: inst = 32'h8220000;
      3942: inst = 32'h10408000;
      3943: inst = 32'hc4047a9;
      3944: inst = 32'h8220000;
      3945: inst = 32'h10408000;
      3946: inst = 32'hc4047aa;
      3947: inst = 32'h8220000;
      3948: inst = 32'h10408000;
      3949: inst = 32'hc4047ab;
      3950: inst = 32'h8220000;
      3951: inst = 32'h10408000;
      3952: inst = 32'hc4047ac;
      3953: inst = 32'h8220000;
      3954: inst = 32'h10408000;
      3955: inst = 32'hc4047ad;
      3956: inst = 32'h8220000;
      3957: inst = 32'h10408000;
      3958: inst = 32'hc4047ae;
      3959: inst = 32'h8220000;
      3960: inst = 32'h10408000;
      3961: inst = 32'hc4047c0;
      3962: inst = 32'h8220000;
      3963: inst = 32'h10408000;
      3964: inst = 32'hc4047c1;
      3965: inst = 32'h8220000;
      3966: inst = 32'h10408000;
      3967: inst = 32'hc4047c2;
      3968: inst = 32'h8220000;
      3969: inst = 32'h10408000;
      3970: inst = 32'hc4047c3;
      3971: inst = 32'h8220000;
      3972: inst = 32'h10408000;
      3973: inst = 32'hc4047c4;
      3974: inst = 32'h8220000;
      3975: inst = 32'h10408000;
      3976: inst = 32'hc4047c5;
      3977: inst = 32'h8220000;
      3978: inst = 32'h10408000;
      3979: inst = 32'hc4047c6;
      3980: inst = 32'h8220000;
      3981: inst = 32'h10408000;
      3982: inst = 32'hc4047c7;
      3983: inst = 32'h8220000;
      3984: inst = 32'h10408000;
      3985: inst = 32'hc4047c8;
      3986: inst = 32'h8220000;
      3987: inst = 32'h10408000;
      3988: inst = 32'hc4047c9;
      3989: inst = 32'h8220000;
      3990: inst = 32'h10408000;
      3991: inst = 32'hc4047ca;
      3992: inst = 32'h8220000;
      3993: inst = 32'h10408000;
      3994: inst = 32'hc4047cb;
      3995: inst = 32'h8220000;
      3996: inst = 32'h10408000;
      3997: inst = 32'hc4047cc;
      3998: inst = 32'h8220000;
      3999: inst = 32'h10408000;
      4000: inst = 32'hc4047cd;
      4001: inst = 32'h8220000;
      4002: inst = 32'h10408000;
      4003: inst = 32'hc4047ce;
      4004: inst = 32'h8220000;
      4005: inst = 32'h10408000;
      4006: inst = 32'hc4047cf;
      4007: inst = 32'h8220000;
      4008: inst = 32'h10408000;
      4009: inst = 32'hc4047d0;
      4010: inst = 32'h8220000;
      4011: inst = 32'h10408000;
      4012: inst = 32'hc4047d1;
      4013: inst = 32'h8220000;
      4014: inst = 32'h10408000;
      4015: inst = 32'hc4047d2;
      4016: inst = 32'h8220000;
      4017: inst = 32'h10408000;
      4018: inst = 32'hc4047d3;
      4019: inst = 32'h8220000;
      4020: inst = 32'h10408000;
      4021: inst = 32'hc4047d4;
      4022: inst = 32'h8220000;
      4023: inst = 32'h10408000;
      4024: inst = 32'hc4047d5;
      4025: inst = 32'h8220000;
      4026: inst = 32'h10408000;
      4027: inst = 32'hc4047d6;
      4028: inst = 32'h8220000;
      4029: inst = 32'h10408000;
      4030: inst = 32'hc4047d7;
      4031: inst = 32'h8220000;
      4032: inst = 32'h10408000;
      4033: inst = 32'hc4047d8;
      4034: inst = 32'h8220000;
      4035: inst = 32'h10408000;
      4036: inst = 32'hc4047d9;
      4037: inst = 32'h8220000;
      4038: inst = 32'h10408000;
      4039: inst = 32'hc4047da;
      4040: inst = 32'h8220000;
      4041: inst = 32'h10408000;
      4042: inst = 32'hc4047db;
      4043: inst = 32'h8220000;
      4044: inst = 32'h10408000;
      4045: inst = 32'hc404804;
      4046: inst = 32'h8220000;
      4047: inst = 32'h10408000;
      4048: inst = 32'hc404805;
      4049: inst = 32'h8220000;
      4050: inst = 32'h10408000;
      4051: inst = 32'hc404806;
      4052: inst = 32'h8220000;
      4053: inst = 32'h10408000;
      4054: inst = 32'hc404807;
      4055: inst = 32'h8220000;
      4056: inst = 32'h10408000;
      4057: inst = 32'hc404808;
      4058: inst = 32'h8220000;
      4059: inst = 32'h10408000;
      4060: inst = 32'hc404809;
      4061: inst = 32'h8220000;
      4062: inst = 32'h10408000;
      4063: inst = 32'hc40480a;
      4064: inst = 32'h8220000;
      4065: inst = 32'h10408000;
      4066: inst = 32'hc40480b;
      4067: inst = 32'h8220000;
      4068: inst = 32'h10408000;
      4069: inst = 32'hc40480c;
      4070: inst = 32'h8220000;
      4071: inst = 32'h10408000;
      4072: inst = 32'hc40480d;
      4073: inst = 32'h8220000;
      4074: inst = 32'h10408000;
      4075: inst = 32'hc40480e;
      4076: inst = 32'h8220000;
      4077: inst = 32'h10408000;
      4078: inst = 32'hc404820;
      4079: inst = 32'h8220000;
      4080: inst = 32'h10408000;
      4081: inst = 32'hc404821;
      4082: inst = 32'h8220000;
      4083: inst = 32'h10408000;
      4084: inst = 32'hc404822;
      4085: inst = 32'h8220000;
      4086: inst = 32'h10408000;
      4087: inst = 32'hc404823;
      4088: inst = 32'h8220000;
      4089: inst = 32'h10408000;
      4090: inst = 32'hc404824;
      4091: inst = 32'h8220000;
      4092: inst = 32'h10408000;
      4093: inst = 32'hc404825;
      4094: inst = 32'h8220000;
      4095: inst = 32'h10408000;
      4096: inst = 32'hc404826;
      4097: inst = 32'h8220000;
      4098: inst = 32'h10408000;
      4099: inst = 32'hc404827;
      4100: inst = 32'h8220000;
      4101: inst = 32'h10408000;
      4102: inst = 32'hc404828;
      4103: inst = 32'h8220000;
      4104: inst = 32'h10408000;
      4105: inst = 32'hc404829;
      4106: inst = 32'h8220000;
      4107: inst = 32'h10408000;
      4108: inst = 32'hc40482a;
      4109: inst = 32'h8220000;
      4110: inst = 32'h10408000;
      4111: inst = 32'hc40482b;
      4112: inst = 32'h8220000;
      4113: inst = 32'h10408000;
      4114: inst = 32'hc40482c;
      4115: inst = 32'h8220000;
      4116: inst = 32'h10408000;
      4117: inst = 32'hc40482d;
      4118: inst = 32'h8220000;
      4119: inst = 32'h10408000;
      4120: inst = 32'hc40482e;
      4121: inst = 32'h8220000;
      4122: inst = 32'h10408000;
      4123: inst = 32'hc40482f;
      4124: inst = 32'h8220000;
      4125: inst = 32'h10408000;
      4126: inst = 32'hc404830;
      4127: inst = 32'h8220000;
      4128: inst = 32'h10408000;
      4129: inst = 32'hc404831;
      4130: inst = 32'h8220000;
      4131: inst = 32'h10408000;
      4132: inst = 32'hc404832;
      4133: inst = 32'h8220000;
      4134: inst = 32'h10408000;
      4135: inst = 32'hc404833;
      4136: inst = 32'h8220000;
      4137: inst = 32'h10408000;
      4138: inst = 32'hc404834;
      4139: inst = 32'h8220000;
      4140: inst = 32'h10408000;
      4141: inst = 32'hc404835;
      4142: inst = 32'h8220000;
      4143: inst = 32'h10408000;
      4144: inst = 32'hc404836;
      4145: inst = 32'h8220000;
      4146: inst = 32'h10408000;
      4147: inst = 32'hc404837;
      4148: inst = 32'h8220000;
      4149: inst = 32'h10408000;
      4150: inst = 32'hc404838;
      4151: inst = 32'h8220000;
      4152: inst = 32'h10408000;
      4153: inst = 32'hc404839;
      4154: inst = 32'h8220000;
      4155: inst = 32'h10408000;
      4156: inst = 32'hc40483a;
      4157: inst = 32'h8220000;
      4158: inst = 32'h10408000;
      4159: inst = 32'hc40483b;
      4160: inst = 32'h8220000;
      4161: inst = 32'h10408000;
      4162: inst = 32'hc404864;
      4163: inst = 32'h8220000;
      4164: inst = 32'h10408000;
      4165: inst = 32'hc404865;
      4166: inst = 32'h8220000;
      4167: inst = 32'h10408000;
      4168: inst = 32'hc404866;
      4169: inst = 32'h8220000;
      4170: inst = 32'h10408000;
      4171: inst = 32'hc404867;
      4172: inst = 32'h8220000;
      4173: inst = 32'h10408000;
      4174: inst = 32'hc404868;
      4175: inst = 32'h8220000;
      4176: inst = 32'h10408000;
      4177: inst = 32'hc404869;
      4178: inst = 32'h8220000;
      4179: inst = 32'h10408000;
      4180: inst = 32'hc40486a;
      4181: inst = 32'h8220000;
      4182: inst = 32'h10408000;
      4183: inst = 32'hc40486b;
      4184: inst = 32'h8220000;
      4185: inst = 32'h10408000;
      4186: inst = 32'hc40486c;
      4187: inst = 32'h8220000;
      4188: inst = 32'h10408000;
      4189: inst = 32'hc40486d;
      4190: inst = 32'h8220000;
      4191: inst = 32'h10408000;
      4192: inst = 32'hc40486e;
      4193: inst = 32'h8220000;
      4194: inst = 32'h10408000;
      4195: inst = 32'hc404880;
      4196: inst = 32'h8220000;
      4197: inst = 32'h10408000;
      4198: inst = 32'hc404881;
      4199: inst = 32'h8220000;
      4200: inst = 32'h10408000;
      4201: inst = 32'hc404882;
      4202: inst = 32'h8220000;
      4203: inst = 32'h10408000;
      4204: inst = 32'hc404883;
      4205: inst = 32'h8220000;
      4206: inst = 32'h10408000;
      4207: inst = 32'hc404884;
      4208: inst = 32'h8220000;
      4209: inst = 32'h10408000;
      4210: inst = 32'hc404885;
      4211: inst = 32'h8220000;
      4212: inst = 32'h10408000;
      4213: inst = 32'hc404886;
      4214: inst = 32'h8220000;
      4215: inst = 32'h10408000;
      4216: inst = 32'hc404887;
      4217: inst = 32'h8220000;
      4218: inst = 32'h10408000;
      4219: inst = 32'hc404888;
      4220: inst = 32'h8220000;
      4221: inst = 32'h10408000;
      4222: inst = 32'hc404889;
      4223: inst = 32'h8220000;
      4224: inst = 32'h10408000;
      4225: inst = 32'hc40488a;
      4226: inst = 32'h8220000;
      4227: inst = 32'h10408000;
      4228: inst = 32'hc40488b;
      4229: inst = 32'h8220000;
      4230: inst = 32'h10408000;
      4231: inst = 32'hc40488c;
      4232: inst = 32'h8220000;
      4233: inst = 32'h10408000;
      4234: inst = 32'hc40488d;
      4235: inst = 32'h8220000;
      4236: inst = 32'h10408000;
      4237: inst = 32'hc40488e;
      4238: inst = 32'h8220000;
      4239: inst = 32'h10408000;
      4240: inst = 32'hc40488f;
      4241: inst = 32'h8220000;
      4242: inst = 32'h10408000;
      4243: inst = 32'hc404890;
      4244: inst = 32'h8220000;
      4245: inst = 32'h10408000;
      4246: inst = 32'hc404891;
      4247: inst = 32'h8220000;
      4248: inst = 32'h10408000;
      4249: inst = 32'hc404892;
      4250: inst = 32'h8220000;
      4251: inst = 32'h10408000;
      4252: inst = 32'hc404893;
      4253: inst = 32'h8220000;
      4254: inst = 32'h10408000;
      4255: inst = 32'hc404894;
      4256: inst = 32'h8220000;
      4257: inst = 32'h10408000;
      4258: inst = 32'hc404895;
      4259: inst = 32'h8220000;
      4260: inst = 32'h10408000;
      4261: inst = 32'hc404896;
      4262: inst = 32'h8220000;
      4263: inst = 32'h10408000;
      4264: inst = 32'hc404897;
      4265: inst = 32'h8220000;
      4266: inst = 32'h10408000;
      4267: inst = 32'hc404898;
      4268: inst = 32'h8220000;
      4269: inst = 32'h10408000;
      4270: inst = 32'hc404899;
      4271: inst = 32'h8220000;
      4272: inst = 32'h10408000;
      4273: inst = 32'hc40489a;
      4274: inst = 32'h8220000;
      4275: inst = 32'h10408000;
      4276: inst = 32'hc40489b;
      4277: inst = 32'h8220000;
      4278: inst = 32'h10408000;
      4279: inst = 32'hc4048c4;
      4280: inst = 32'h8220000;
      4281: inst = 32'h10408000;
      4282: inst = 32'hc4048c5;
      4283: inst = 32'h8220000;
      4284: inst = 32'h10408000;
      4285: inst = 32'hc4048c6;
      4286: inst = 32'h8220000;
      4287: inst = 32'h10408000;
      4288: inst = 32'hc4048c7;
      4289: inst = 32'h8220000;
      4290: inst = 32'h10408000;
      4291: inst = 32'hc4048c8;
      4292: inst = 32'h8220000;
      4293: inst = 32'h10408000;
      4294: inst = 32'hc4048c9;
      4295: inst = 32'h8220000;
      4296: inst = 32'h10408000;
      4297: inst = 32'hc4048ca;
      4298: inst = 32'h8220000;
      4299: inst = 32'h10408000;
      4300: inst = 32'hc4048cb;
      4301: inst = 32'h8220000;
      4302: inst = 32'h10408000;
      4303: inst = 32'hc4048cc;
      4304: inst = 32'h8220000;
      4305: inst = 32'h10408000;
      4306: inst = 32'hc4048cd;
      4307: inst = 32'h8220000;
      4308: inst = 32'h10408000;
      4309: inst = 32'hc4048ce;
      4310: inst = 32'h8220000;
      4311: inst = 32'h10408000;
      4312: inst = 32'hc4048e0;
      4313: inst = 32'h8220000;
      4314: inst = 32'h10408000;
      4315: inst = 32'hc4048e1;
      4316: inst = 32'h8220000;
      4317: inst = 32'h10408000;
      4318: inst = 32'hc4048e2;
      4319: inst = 32'h8220000;
      4320: inst = 32'h10408000;
      4321: inst = 32'hc4048e3;
      4322: inst = 32'h8220000;
      4323: inst = 32'h10408000;
      4324: inst = 32'hc4048e4;
      4325: inst = 32'h8220000;
      4326: inst = 32'h10408000;
      4327: inst = 32'hc4048e5;
      4328: inst = 32'h8220000;
      4329: inst = 32'h10408000;
      4330: inst = 32'hc4048e6;
      4331: inst = 32'h8220000;
      4332: inst = 32'h10408000;
      4333: inst = 32'hc4048e7;
      4334: inst = 32'h8220000;
      4335: inst = 32'h10408000;
      4336: inst = 32'hc4048e8;
      4337: inst = 32'h8220000;
      4338: inst = 32'h10408000;
      4339: inst = 32'hc4048e9;
      4340: inst = 32'h8220000;
      4341: inst = 32'h10408000;
      4342: inst = 32'hc4048ea;
      4343: inst = 32'h8220000;
      4344: inst = 32'h10408000;
      4345: inst = 32'hc4048eb;
      4346: inst = 32'h8220000;
      4347: inst = 32'h10408000;
      4348: inst = 32'hc4048ec;
      4349: inst = 32'h8220000;
      4350: inst = 32'h10408000;
      4351: inst = 32'hc4048ed;
      4352: inst = 32'h8220000;
      4353: inst = 32'h10408000;
      4354: inst = 32'hc4048ee;
      4355: inst = 32'h8220000;
      4356: inst = 32'h10408000;
      4357: inst = 32'hc4048ef;
      4358: inst = 32'h8220000;
      4359: inst = 32'h10408000;
      4360: inst = 32'hc4048f0;
      4361: inst = 32'h8220000;
      4362: inst = 32'h10408000;
      4363: inst = 32'hc4048f1;
      4364: inst = 32'h8220000;
      4365: inst = 32'h10408000;
      4366: inst = 32'hc4048f2;
      4367: inst = 32'h8220000;
      4368: inst = 32'h10408000;
      4369: inst = 32'hc4048f3;
      4370: inst = 32'h8220000;
      4371: inst = 32'h10408000;
      4372: inst = 32'hc4048f4;
      4373: inst = 32'h8220000;
      4374: inst = 32'h10408000;
      4375: inst = 32'hc4048f5;
      4376: inst = 32'h8220000;
      4377: inst = 32'h10408000;
      4378: inst = 32'hc4048f6;
      4379: inst = 32'h8220000;
      4380: inst = 32'h10408000;
      4381: inst = 32'hc4048f7;
      4382: inst = 32'h8220000;
      4383: inst = 32'h10408000;
      4384: inst = 32'hc4048f8;
      4385: inst = 32'h8220000;
      4386: inst = 32'h10408000;
      4387: inst = 32'hc4048f9;
      4388: inst = 32'h8220000;
      4389: inst = 32'h10408000;
      4390: inst = 32'hc4048fa;
      4391: inst = 32'h8220000;
      4392: inst = 32'h10408000;
      4393: inst = 32'hc4048fb;
      4394: inst = 32'h8220000;
      4395: inst = 32'h10408000;
      4396: inst = 32'hc404924;
      4397: inst = 32'h8220000;
      4398: inst = 32'h10408000;
      4399: inst = 32'hc404925;
      4400: inst = 32'h8220000;
      4401: inst = 32'h10408000;
      4402: inst = 32'hc404926;
      4403: inst = 32'h8220000;
      4404: inst = 32'h10408000;
      4405: inst = 32'hc404927;
      4406: inst = 32'h8220000;
      4407: inst = 32'h10408000;
      4408: inst = 32'hc404928;
      4409: inst = 32'h8220000;
      4410: inst = 32'h10408000;
      4411: inst = 32'hc404929;
      4412: inst = 32'h8220000;
      4413: inst = 32'h10408000;
      4414: inst = 32'hc40492a;
      4415: inst = 32'h8220000;
      4416: inst = 32'h10408000;
      4417: inst = 32'hc40492b;
      4418: inst = 32'h8220000;
      4419: inst = 32'h10408000;
      4420: inst = 32'hc40492c;
      4421: inst = 32'h8220000;
      4422: inst = 32'h10408000;
      4423: inst = 32'hc40492d;
      4424: inst = 32'h8220000;
      4425: inst = 32'h10408000;
      4426: inst = 32'hc40492e;
      4427: inst = 32'h8220000;
      4428: inst = 32'h10408000;
      4429: inst = 32'hc404940;
      4430: inst = 32'h8220000;
      4431: inst = 32'h10408000;
      4432: inst = 32'hc404941;
      4433: inst = 32'h8220000;
      4434: inst = 32'h10408000;
      4435: inst = 32'hc404942;
      4436: inst = 32'h8220000;
      4437: inst = 32'h10408000;
      4438: inst = 32'hc404943;
      4439: inst = 32'h8220000;
      4440: inst = 32'h10408000;
      4441: inst = 32'hc404944;
      4442: inst = 32'h8220000;
      4443: inst = 32'h10408000;
      4444: inst = 32'hc404945;
      4445: inst = 32'h8220000;
      4446: inst = 32'h10408000;
      4447: inst = 32'hc404946;
      4448: inst = 32'h8220000;
      4449: inst = 32'h10408000;
      4450: inst = 32'hc404947;
      4451: inst = 32'h8220000;
      4452: inst = 32'h10408000;
      4453: inst = 32'hc404948;
      4454: inst = 32'h8220000;
      4455: inst = 32'h10408000;
      4456: inst = 32'hc404949;
      4457: inst = 32'h8220000;
      4458: inst = 32'h10408000;
      4459: inst = 32'hc40494a;
      4460: inst = 32'h8220000;
      4461: inst = 32'h10408000;
      4462: inst = 32'hc40494b;
      4463: inst = 32'h8220000;
      4464: inst = 32'h10408000;
      4465: inst = 32'hc40494c;
      4466: inst = 32'h8220000;
      4467: inst = 32'h10408000;
      4468: inst = 32'hc40494d;
      4469: inst = 32'h8220000;
      4470: inst = 32'h10408000;
      4471: inst = 32'hc40494e;
      4472: inst = 32'h8220000;
      4473: inst = 32'h10408000;
      4474: inst = 32'hc40494f;
      4475: inst = 32'h8220000;
      4476: inst = 32'h10408000;
      4477: inst = 32'hc404950;
      4478: inst = 32'h8220000;
      4479: inst = 32'h10408000;
      4480: inst = 32'hc404951;
      4481: inst = 32'h8220000;
      4482: inst = 32'h10408000;
      4483: inst = 32'hc404952;
      4484: inst = 32'h8220000;
      4485: inst = 32'h10408000;
      4486: inst = 32'hc404953;
      4487: inst = 32'h8220000;
      4488: inst = 32'h10408000;
      4489: inst = 32'hc404954;
      4490: inst = 32'h8220000;
      4491: inst = 32'h10408000;
      4492: inst = 32'hc404955;
      4493: inst = 32'h8220000;
      4494: inst = 32'h10408000;
      4495: inst = 32'hc404956;
      4496: inst = 32'h8220000;
      4497: inst = 32'h10408000;
      4498: inst = 32'hc404957;
      4499: inst = 32'h8220000;
      4500: inst = 32'h10408000;
      4501: inst = 32'hc404958;
      4502: inst = 32'h8220000;
      4503: inst = 32'h10408000;
      4504: inst = 32'hc404959;
      4505: inst = 32'h8220000;
      4506: inst = 32'h10408000;
      4507: inst = 32'hc40495a;
      4508: inst = 32'h8220000;
      4509: inst = 32'h10408000;
      4510: inst = 32'hc40495b;
      4511: inst = 32'h8220000;
      4512: inst = 32'h10408000;
      4513: inst = 32'hc404984;
      4514: inst = 32'h8220000;
      4515: inst = 32'h10408000;
      4516: inst = 32'hc404985;
      4517: inst = 32'h8220000;
      4518: inst = 32'h10408000;
      4519: inst = 32'hc404986;
      4520: inst = 32'h8220000;
      4521: inst = 32'h10408000;
      4522: inst = 32'hc404987;
      4523: inst = 32'h8220000;
      4524: inst = 32'h10408000;
      4525: inst = 32'hc404988;
      4526: inst = 32'h8220000;
      4527: inst = 32'h10408000;
      4528: inst = 32'hc404989;
      4529: inst = 32'h8220000;
      4530: inst = 32'h10408000;
      4531: inst = 32'hc40498a;
      4532: inst = 32'h8220000;
      4533: inst = 32'h10408000;
      4534: inst = 32'hc40498b;
      4535: inst = 32'h8220000;
      4536: inst = 32'h10408000;
      4537: inst = 32'hc40498c;
      4538: inst = 32'h8220000;
      4539: inst = 32'h10408000;
      4540: inst = 32'hc40498d;
      4541: inst = 32'h8220000;
      4542: inst = 32'h10408000;
      4543: inst = 32'hc40498e;
      4544: inst = 32'h8220000;
      4545: inst = 32'h10408000;
      4546: inst = 32'hc4049a0;
      4547: inst = 32'h8220000;
      4548: inst = 32'h10408000;
      4549: inst = 32'hc4049a1;
      4550: inst = 32'h8220000;
      4551: inst = 32'h10408000;
      4552: inst = 32'hc4049a2;
      4553: inst = 32'h8220000;
      4554: inst = 32'h10408000;
      4555: inst = 32'hc4049a3;
      4556: inst = 32'h8220000;
      4557: inst = 32'h10408000;
      4558: inst = 32'hc4049a4;
      4559: inst = 32'h8220000;
      4560: inst = 32'h10408000;
      4561: inst = 32'hc4049a5;
      4562: inst = 32'h8220000;
      4563: inst = 32'h10408000;
      4564: inst = 32'hc4049a6;
      4565: inst = 32'h8220000;
      4566: inst = 32'h10408000;
      4567: inst = 32'hc4049a7;
      4568: inst = 32'h8220000;
      4569: inst = 32'h10408000;
      4570: inst = 32'hc4049a8;
      4571: inst = 32'h8220000;
      4572: inst = 32'h10408000;
      4573: inst = 32'hc4049a9;
      4574: inst = 32'h8220000;
      4575: inst = 32'h10408000;
      4576: inst = 32'hc4049aa;
      4577: inst = 32'h8220000;
      4578: inst = 32'h10408000;
      4579: inst = 32'hc4049ab;
      4580: inst = 32'h8220000;
      4581: inst = 32'h10408000;
      4582: inst = 32'hc4049ac;
      4583: inst = 32'h8220000;
      4584: inst = 32'h10408000;
      4585: inst = 32'hc4049ad;
      4586: inst = 32'h8220000;
      4587: inst = 32'h10408000;
      4588: inst = 32'hc4049ae;
      4589: inst = 32'h8220000;
      4590: inst = 32'h10408000;
      4591: inst = 32'hc4049af;
      4592: inst = 32'h8220000;
      4593: inst = 32'h10408000;
      4594: inst = 32'hc4049b0;
      4595: inst = 32'h8220000;
      4596: inst = 32'h10408000;
      4597: inst = 32'hc4049b1;
      4598: inst = 32'h8220000;
      4599: inst = 32'h10408000;
      4600: inst = 32'hc4049b2;
      4601: inst = 32'h8220000;
      4602: inst = 32'h10408000;
      4603: inst = 32'hc4049b3;
      4604: inst = 32'h8220000;
      4605: inst = 32'h10408000;
      4606: inst = 32'hc4049b4;
      4607: inst = 32'h8220000;
      4608: inst = 32'h10408000;
      4609: inst = 32'hc4049b5;
      4610: inst = 32'h8220000;
      4611: inst = 32'h10408000;
      4612: inst = 32'hc4049b6;
      4613: inst = 32'h8220000;
      4614: inst = 32'h10408000;
      4615: inst = 32'hc4049b7;
      4616: inst = 32'h8220000;
      4617: inst = 32'h10408000;
      4618: inst = 32'hc4049b8;
      4619: inst = 32'h8220000;
      4620: inst = 32'h10408000;
      4621: inst = 32'hc4049b9;
      4622: inst = 32'h8220000;
      4623: inst = 32'h10408000;
      4624: inst = 32'hc4049ba;
      4625: inst = 32'h8220000;
      4626: inst = 32'h10408000;
      4627: inst = 32'hc4049bb;
      4628: inst = 32'h8220000;
      4629: inst = 32'h10408000;
      4630: inst = 32'hc4049e4;
      4631: inst = 32'h8220000;
      4632: inst = 32'h10408000;
      4633: inst = 32'hc4049e5;
      4634: inst = 32'h8220000;
      4635: inst = 32'h10408000;
      4636: inst = 32'hc4049e6;
      4637: inst = 32'h8220000;
      4638: inst = 32'h10408000;
      4639: inst = 32'hc4049e7;
      4640: inst = 32'h8220000;
      4641: inst = 32'h10408000;
      4642: inst = 32'hc4049e8;
      4643: inst = 32'h8220000;
      4644: inst = 32'h10408000;
      4645: inst = 32'hc4049e9;
      4646: inst = 32'h8220000;
      4647: inst = 32'h10408000;
      4648: inst = 32'hc4049ea;
      4649: inst = 32'h8220000;
      4650: inst = 32'h10408000;
      4651: inst = 32'hc4049eb;
      4652: inst = 32'h8220000;
      4653: inst = 32'h10408000;
      4654: inst = 32'hc4049ec;
      4655: inst = 32'h8220000;
      4656: inst = 32'h10408000;
      4657: inst = 32'hc4049ed;
      4658: inst = 32'h8220000;
      4659: inst = 32'h10408000;
      4660: inst = 32'hc4049ee;
      4661: inst = 32'h8220000;
      4662: inst = 32'h10408000;
      4663: inst = 32'hc404a00;
      4664: inst = 32'h8220000;
      4665: inst = 32'h10408000;
      4666: inst = 32'hc404a01;
      4667: inst = 32'h8220000;
      4668: inst = 32'h10408000;
      4669: inst = 32'hc404a02;
      4670: inst = 32'h8220000;
      4671: inst = 32'h10408000;
      4672: inst = 32'hc404a03;
      4673: inst = 32'h8220000;
      4674: inst = 32'h10408000;
      4675: inst = 32'hc404a04;
      4676: inst = 32'h8220000;
      4677: inst = 32'h10408000;
      4678: inst = 32'hc404a05;
      4679: inst = 32'h8220000;
      4680: inst = 32'h10408000;
      4681: inst = 32'hc404a06;
      4682: inst = 32'h8220000;
      4683: inst = 32'h10408000;
      4684: inst = 32'hc404a07;
      4685: inst = 32'h8220000;
      4686: inst = 32'h10408000;
      4687: inst = 32'hc404a0f;
      4688: inst = 32'h8220000;
      4689: inst = 32'h10408000;
      4690: inst = 32'hc404a10;
      4691: inst = 32'h8220000;
      4692: inst = 32'h10408000;
      4693: inst = 32'hc404a11;
      4694: inst = 32'h8220000;
      4695: inst = 32'h10408000;
      4696: inst = 32'hc404a12;
      4697: inst = 32'h8220000;
      4698: inst = 32'h10408000;
      4699: inst = 32'hc404a13;
      4700: inst = 32'h8220000;
      4701: inst = 32'h10408000;
      4702: inst = 32'hc404a14;
      4703: inst = 32'h8220000;
      4704: inst = 32'h10408000;
      4705: inst = 32'hc404a15;
      4706: inst = 32'h8220000;
      4707: inst = 32'h10408000;
      4708: inst = 32'hc404a16;
      4709: inst = 32'h8220000;
      4710: inst = 32'h10408000;
      4711: inst = 32'hc404a17;
      4712: inst = 32'h8220000;
      4713: inst = 32'h10408000;
      4714: inst = 32'hc404a18;
      4715: inst = 32'h8220000;
      4716: inst = 32'h10408000;
      4717: inst = 32'hc404a19;
      4718: inst = 32'h8220000;
      4719: inst = 32'h10408000;
      4720: inst = 32'hc404a1a;
      4721: inst = 32'h8220000;
      4722: inst = 32'h10408000;
      4723: inst = 32'hc404a1b;
      4724: inst = 32'h8220000;
      4725: inst = 32'h10408000;
      4726: inst = 32'hc404a44;
      4727: inst = 32'h8220000;
      4728: inst = 32'h10408000;
      4729: inst = 32'hc404a45;
      4730: inst = 32'h8220000;
      4731: inst = 32'h10408000;
      4732: inst = 32'hc404a46;
      4733: inst = 32'h8220000;
      4734: inst = 32'h10408000;
      4735: inst = 32'hc404a47;
      4736: inst = 32'h8220000;
      4737: inst = 32'h10408000;
      4738: inst = 32'hc404a48;
      4739: inst = 32'h8220000;
      4740: inst = 32'h10408000;
      4741: inst = 32'hc404a49;
      4742: inst = 32'h8220000;
      4743: inst = 32'h10408000;
      4744: inst = 32'hc404a4a;
      4745: inst = 32'h8220000;
      4746: inst = 32'h10408000;
      4747: inst = 32'hc404a4b;
      4748: inst = 32'h8220000;
      4749: inst = 32'h10408000;
      4750: inst = 32'hc404a4c;
      4751: inst = 32'h8220000;
      4752: inst = 32'h10408000;
      4753: inst = 32'hc404a4d;
      4754: inst = 32'h8220000;
      4755: inst = 32'h10408000;
      4756: inst = 32'hc404a4e;
      4757: inst = 32'h8220000;
      4758: inst = 32'h10408000;
      4759: inst = 32'hc404a60;
      4760: inst = 32'h8220000;
      4761: inst = 32'h10408000;
      4762: inst = 32'hc404a61;
      4763: inst = 32'h8220000;
      4764: inst = 32'h10408000;
      4765: inst = 32'hc404a62;
      4766: inst = 32'h8220000;
      4767: inst = 32'h10408000;
      4768: inst = 32'hc404a63;
      4769: inst = 32'h8220000;
      4770: inst = 32'h10408000;
      4771: inst = 32'hc404a64;
      4772: inst = 32'h8220000;
      4773: inst = 32'h10408000;
      4774: inst = 32'hc404a65;
      4775: inst = 32'h8220000;
      4776: inst = 32'h10408000;
      4777: inst = 32'hc404a66;
      4778: inst = 32'h8220000;
      4779: inst = 32'h10408000;
      4780: inst = 32'hc404a70;
      4781: inst = 32'h8220000;
      4782: inst = 32'h10408000;
      4783: inst = 32'hc404a71;
      4784: inst = 32'h8220000;
      4785: inst = 32'h10408000;
      4786: inst = 32'hc404a72;
      4787: inst = 32'h8220000;
      4788: inst = 32'h10408000;
      4789: inst = 32'hc404a73;
      4790: inst = 32'h8220000;
      4791: inst = 32'h10408000;
      4792: inst = 32'hc404a74;
      4793: inst = 32'h8220000;
      4794: inst = 32'h10408000;
      4795: inst = 32'hc404a75;
      4796: inst = 32'h8220000;
      4797: inst = 32'h10408000;
      4798: inst = 32'hc404a76;
      4799: inst = 32'h8220000;
      4800: inst = 32'h10408000;
      4801: inst = 32'hc404a77;
      4802: inst = 32'h8220000;
      4803: inst = 32'h10408000;
      4804: inst = 32'hc404a78;
      4805: inst = 32'h8220000;
      4806: inst = 32'h10408000;
      4807: inst = 32'hc404a79;
      4808: inst = 32'h8220000;
      4809: inst = 32'h10408000;
      4810: inst = 32'hc404a7a;
      4811: inst = 32'h8220000;
      4812: inst = 32'h10408000;
      4813: inst = 32'hc404a7b;
      4814: inst = 32'h8220000;
      4815: inst = 32'h10408000;
      4816: inst = 32'hc404aa4;
      4817: inst = 32'h8220000;
      4818: inst = 32'h10408000;
      4819: inst = 32'hc404aa5;
      4820: inst = 32'h8220000;
      4821: inst = 32'h10408000;
      4822: inst = 32'hc404aa6;
      4823: inst = 32'h8220000;
      4824: inst = 32'h10408000;
      4825: inst = 32'hc404aa7;
      4826: inst = 32'h8220000;
      4827: inst = 32'h10408000;
      4828: inst = 32'hc404aa8;
      4829: inst = 32'h8220000;
      4830: inst = 32'h10408000;
      4831: inst = 32'hc404aa9;
      4832: inst = 32'h8220000;
      4833: inst = 32'h10408000;
      4834: inst = 32'hc404aaa;
      4835: inst = 32'h8220000;
      4836: inst = 32'h10408000;
      4837: inst = 32'hc404aab;
      4838: inst = 32'h8220000;
      4839: inst = 32'h10408000;
      4840: inst = 32'hc404aac;
      4841: inst = 32'h8220000;
      4842: inst = 32'h10408000;
      4843: inst = 32'hc404aad;
      4844: inst = 32'h8220000;
      4845: inst = 32'h10408000;
      4846: inst = 32'hc404aae;
      4847: inst = 32'h8220000;
      4848: inst = 32'h10408000;
      4849: inst = 32'hc404ac0;
      4850: inst = 32'h8220000;
      4851: inst = 32'h10408000;
      4852: inst = 32'hc404ac1;
      4853: inst = 32'h8220000;
      4854: inst = 32'h10408000;
      4855: inst = 32'hc404ac2;
      4856: inst = 32'h8220000;
      4857: inst = 32'h10408000;
      4858: inst = 32'hc404ac3;
      4859: inst = 32'h8220000;
      4860: inst = 32'h10408000;
      4861: inst = 32'hc404ac4;
      4862: inst = 32'h8220000;
      4863: inst = 32'h10408000;
      4864: inst = 32'hc404ac5;
      4865: inst = 32'h8220000;
      4866: inst = 32'h10408000;
      4867: inst = 32'hc404ac6;
      4868: inst = 32'h8220000;
      4869: inst = 32'h10408000;
      4870: inst = 32'hc404ad0;
      4871: inst = 32'h8220000;
      4872: inst = 32'h10408000;
      4873: inst = 32'hc404ad1;
      4874: inst = 32'h8220000;
      4875: inst = 32'h10408000;
      4876: inst = 32'hc404ad2;
      4877: inst = 32'h8220000;
      4878: inst = 32'h10408000;
      4879: inst = 32'hc404ad3;
      4880: inst = 32'h8220000;
      4881: inst = 32'h10408000;
      4882: inst = 32'hc404ad4;
      4883: inst = 32'h8220000;
      4884: inst = 32'h10408000;
      4885: inst = 32'hc404ad5;
      4886: inst = 32'h8220000;
      4887: inst = 32'h10408000;
      4888: inst = 32'hc404ad6;
      4889: inst = 32'h8220000;
      4890: inst = 32'h10408000;
      4891: inst = 32'hc404ad7;
      4892: inst = 32'h8220000;
      4893: inst = 32'h10408000;
      4894: inst = 32'hc404ad8;
      4895: inst = 32'h8220000;
      4896: inst = 32'h10408000;
      4897: inst = 32'hc404ad9;
      4898: inst = 32'h8220000;
      4899: inst = 32'h10408000;
      4900: inst = 32'hc404ada;
      4901: inst = 32'h8220000;
      4902: inst = 32'h10408000;
      4903: inst = 32'hc404adb;
      4904: inst = 32'h8220000;
      4905: inst = 32'h10408000;
      4906: inst = 32'hc404b04;
      4907: inst = 32'h8220000;
      4908: inst = 32'h10408000;
      4909: inst = 32'hc404b05;
      4910: inst = 32'h8220000;
      4911: inst = 32'h10408000;
      4912: inst = 32'hc404b06;
      4913: inst = 32'h8220000;
      4914: inst = 32'h10408000;
      4915: inst = 32'hc404b07;
      4916: inst = 32'h8220000;
      4917: inst = 32'h10408000;
      4918: inst = 32'hc404b08;
      4919: inst = 32'h8220000;
      4920: inst = 32'h10408000;
      4921: inst = 32'hc404b09;
      4922: inst = 32'h8220000;
      4923: inst = 32'h10408000;
      4924: inst = 32'hc404b0a;
      4925: inst = 32'h8220000;
      4926: inst = 32'h10408000;
      4927: inst = 32'hc404b0b;
      4928: inst = 32'h8220000;
      4929: inst = 32'h10408000;
      4930: inst = 32'hc404b0c;
      4931: inst = 32'h8220000;
      4932: inst = 32'h10408000;
      4933: inst = 32'hc404b0d;
      4934: inst = 32'h8220000;
      4935: inst = 32'h10408000;
      4936: inst = 32'hc404b0e;
      4937: inst = 32'h8220000;
      4938: inst = 32'h10408000;
      4939: inst = 32'hc404b20;
      4940: inst = 32'h8220000;
      4941: inst = 32'h10408000;
      4942: inst = 32'hc404b21;
      4943: inst = 32'h8220000;
      4944: inst = 32'h10408000;
      4945: inst = 32'hc404b22;
      4946: inst = 32'h8220000;
      4947: inst = 32'h10408000;
      4948: inst = 32'hc404b23;
      4949: inst = 32'h8220000;
      4950: inst = 32'h10408000;
      4951: inst = 32'hc404b24;
      4952: inst = 32'h8220000;
      4953: inst = 32'h10408000;
      4954: inst = 32'hc404b25;
      4955: inst = 32'h8220000;
      4956: inst = 32'h10408000;
      4957: inst = 32'hc404b26;
      4958: inst = 32'h8220000;
      4959: inst = 32'h10408000;
      4960: inst = 32'hc404b30;
      4961: inst = 32'h8220000;
      4962: inst = 32'h10408000;
      4963: inst = 32'hc404b31;
      4964: inst = 32'h8220000;
      4965: inst = 32'h10408000;
      4966: inst = 32'hc404b32;
      4967: inst = 32'h8220000;
      4968: inst = 32'h10408000;
      4969: inst = 32'hc404b33;
      4970: inst = 32'h8220000;
      4971: inst = 32'h10408000;
      4972: inst = 32'hc404b34;
      4973: inst = 32'h8220000;
      4974: inst = 32'h10408000;
      4975: inst = 32'hc404b35;
      4976: inst = 32'h8220000;
      4977: inst = 32'h10408000;
      4978: inst = 32'hc404b36;
      4979: inst = 32'h8220000;
      4980: inst = 32'h10408000;
      4981: inst = 32'hc404b37;
      4982: inst = 32'h8220000;
      4983: inst = 32'h10408000;
      4984: inst = 32'hc404b38;
      4985: inst = 32'h8220000;
      4986: inst = 32'h10408000;
      4987: inst = 32'hc404b39;
      4988: inst = 32'h8220000;
      4989: inst = 32'h10408000;
      4990: inst = 32'hc404b3a;
      4991: inst = 32'h8220000;
      4992: inst = 32'h10408000;
      4993: inst = 32'hc404b3b;
      4994: inst = 32'h8220000;
      4995: inst = 32'h10408000;
      4996: inst = 32'hc404b64;
      4997: inst = 32'h8220000;
      4998: inst = 32'h10408000;
      4999: inst = 32'hc404b65;
      5000: inst = 32'h8220000;
      5001: inst = 32'h10408000;
      5002: inst = 32'hc404b66;
      5003: inst = 32'h8220000;
      5004: inst = 32'h10408000;
      5005: inst = 32'hc404b67;
      5006: inst = 32'h8220000;
      5007: inst = 32'h10408000;
      5008: inst = 32'hc404b68;
      5009: inst = 32'h8220000;
      5010: inst = 32'h10408000;
      5011: inst = 32'hc404b69;
      5012: inst = 32'h8220000;
      5013: inst = 32'h10408000;
      5014: inst = 32'hc404b6a;
      5015: inst = 32'h8220000;
      5016: inst = 32'h10408000;
      5017: inst = 32'hc404b6b;
      5018: inst = 32'h8220000;
      5019: inst = 32'h10408000;
      5020: inst = 32'hc404b6c;
      5021: inst = 32'h8220000;
      5022: inst = 32'h10408000;
      5023: inst = 32'hc404b6d;
      5024: inst = 32'h8220000;
      5025: inst = 32'h10408000;
      5026: inst = 32'hc404b6e;
      5027: inst = 32'h8220000;
      5028: inst = 32'h10408000;
      5029: inst = 32'hc404b80;
      5030: inst = 32'h8220000;
      5031: inst = 32'h10408000;
      5032: inst = 32'hc404b81;
      5033: inst = 32'h8220000;
      5034: inst = 32'h10408000;
      5035: inst = 32'hc404b82;
      5036: inst = 32'h8220000;
      5037: inst = 32'h10408000;
      5038: inst = 32'hc404b83;
      5039: inst = 32'h8220000;
      5040: inst = 32'h10408000;
      5041: inst = 32'hc404b84;
      5042: inst = 32'h8220000;
      5043: inst = 32'h10408000;
      5044: inst = 32'hc404b85;
      5045: inst = 32'h8220000;
      5046: inst = 32'h10408000;
      5047: inst = 32'hc404b86;
      5048: inst = 32'h8220000;
      5049: inst = 32'h10408000;
      5050: inst = 32'hc404b90;
      5051: inst = 32'h8220000;
      5052: inst = 32'h10408000;
      5053: inst = 32'hc404b91;
      5054: inst = 32'h8220000;
      5055: inst = 32'h10408000;
      5056: inst = 32'hc404b92;
      5057: inst = 32'h8220000;
      5058: inst = 32'h10408000;
      5059: inst = 32'hc404b93;
      5060: inst = 32'h8220000;
      5061: inst = 32'h10408000;
      5062: inst = 32'hc404b94;
      5063: inst = 32'h8220000;
      5064: inst = 32'h10408000;
      5065: inst = 32'hc404b95;
      5066: inst = 32'h8220000;
      5067: inst = 32'h10408000;
      5068: inst = 32'hc404b96;
      5069: inst = 32'h8220000;
      5070: inst = 32'h10408000;
      5071: inst = 32'hc404b97;
      5072: inst = 32'h8220000;
      5073: inst = 32'h10408000;
      5074: inst = 32'hc404b98;
      5075: inst = 32'h8220000;
      5076: inst = 32'h10408000;
      5077: inst = 32'hc404b99;
      5078: inst = 32'h8220000;
      5079: inst = 32'h10408000;
      5080: inst = 32'hc404b9a;
      5081: inst = 32'h8220000;
      5082: inst = 32'h10408000;
      5083: inst = 32'hc404b9b;
      5084: inst = 32'h8220000;
      5085: inst = 32'h10408000;
      5086: inst = 32'hc404bc4;
      5087: inst = 32'h8220000;
      5088: inst = 32'h10408000;
      5089: inst = 32'hc404bc5;
      5090: inst = 32'h8220000;
      5091: inst = 32'h10408000;
      5092: inst = 32'hc404bc6;
      5093: inst = 32'h8220000;
      5094: inst = 32'h10408000;
      5095: inst = 32'hc404bc7;
      5096: inst = 32'h8220000;
      5097: inst = 32'h10408000;
      5098: inst = 32'hc404bc8;
      5099: inst = 32'h8220000;
      5100: inst = 32'h10408000;
      5101: inst = 32'hc404bc9;
      5102: inst = 32'h8220000;
      5103: inst = 32'h10408000;
      5104: inst = 32'hc404bca;
      5105: inst = 32'h8220000;
      5106: inst = 32'h10408000;
      5107: inst = 32'hc404bcb;
      5108: inst = 32'h8220000;
      5109: inst = 32'h10408000;
      5110: inst = 32'hc404bcc;
      5111: inst = 32'h8220000;
      5112: inst = 32'h10408000;
      5113: inst = 32'hc404bcd;
      5114: inst = 32'h8220000;
      5115: inst = 32'h10408000;
      5116: inst = 32'hc404bce;
      5117: inst = 32'h8220000;
      5118: inst = 32'h10408000;
      5119: inst = 32'hc404be0;
      5120: inst = 32'h8220000;
      5121: inst = 32'h10408000;
      5122: inst = 32'hc404be1;
      5123: inst = 32'h8220000;
      5124: inst = 32'h10408000;
      5125: inst = 32'hc404be2;
      5126: inst = 32'h8220000;
      5127: inst = 32'h10408000;
      5128: inst = 32'hc404be3;
      5129: inst = 32'h8220000;
      5130: inst = 32'h10408000;
      5131: inst = 32'hc404be4;
      5132: inst = 32'h8220000;
      5133: inst = 32'h10408000;
      5134: inst = 32'hc404be5;
      5135: inst = 32'h8220000;
      5136: inst = 32'h10408000;
      5137: inst = 32'hc404be6;
      5138: inst = 32'h8220000;
      5139: inst = 32'h10408000;
      5140: inst = 32'hc404bf0;
      5141: inst = 32'h8220000;
      5142: inst = 32'h10408000;
      5143: inst = 32'hc404bf1;
      5144: inst = 32'h8220000;
      5145: inst = 32'h10408000;
      5146: inst = 32'hc404bf2;
      5147: inst = 32'h8220000;
      5148: inst = 32'h10408000;
      5149: inst = 32'hc404bf3;
      5150: inst = 32'h8220000;
      5151: inst = 32'h10408000;
      5152: inst = 32'hc404bf4;
      5153: inst = 32'h8220000;
      5154: inst = 32'h10408000;
      5155: inst = 32'hc404bf5;
      5156: inst = 32'h8220000;
      5157: inst = 32'h10408000;
      5158: inst = 32'hc404bf6;
      5159: inst = 32'h8220000;
      5160: inst = 32'h10408000;
      5161: inst = 32'hc404bf7;
      5162: inst = 32'h8220000;
      5163: inst = 32'h10408000;
      5164: inst = 32'hc404bf8;
      5165: inst = 32'h8220000;
      5166: inst = 32'h10408000;
      5167: inst = 32'hc404bf9;
      5168: inst = 32'h8220000;
      5169: inst = 32'h10408000;
      5170: inst = 32'hc404c26;
      5171: inst = 32'h8220000;
      5172: inst = 32'h10408000;
      5173: inst = 32'hc404c27;
      5174: inst = 32'h8220000;
      5175: inst = 32'h10408000;
      5176: inst = 32'hc404c28;
      5177: inst = 32'h8220000;
      5178: inst = 32'h10408000;
      5179: inst = 32'hc404c29;
      5180: inst = 32'h8220000;
      5181: inst = 32'h10408000;
      5182: inst = 32'hc404c2a;
      5183: inst = 32'h8220000;
      5184: inst = 32'h10408000;
      5185: inst = 32'hc404c2b;
      5186: inst = 32'h8220000;
      5187: inst = 32'h10408000;
      5188: inst = 32'hc404c2c;
      5189: inst = 32'h8220000;
      5190: inst = 32'h10408000;
      5191: inst = 32'hc404c2d;
      5192: inst = 32'h8220000;
      5193: inst = 32'h10408000;
      5194: inst = 32'hc404c2e;
      5195: inst = 32'h8220000;
      5196: inst = 32'h10408000;
      5197: inst = 32'hc404c40;
      5198: inst = 32'h8220000;
      5199: inst = 32'h10408000;
      5200: inst = 32'hc404c41;
      5201: inst = 32'h8220000;
      5202: inst = 32'h10408000;
      5203: inst = 32'hc404c42;
      5204: inst = 32'h8220000;
      5205: inst = 32'h10408000;
      5206: inst = 32'hc404c43;
      5207: inst = 32'h8220000;
      5208: inst = 32'h10408000;
      5209: inst = 32'hc404c44;
      5210: inst = 32'h8220000;
      5211: inst = 32'h10408000;
      5212: inst = 32'hc404c45;
      5213: inst = 32'h8220000;
      5214: inst = 32'h10408000;
      5215: inst = 32'hc404c46;
      5216: inst = 32'h8220000;
      5217: inst = 32'h10408000;
      5218: inst = 32'hc404c4f;
      5219: inst = 32'h8220000;
      5220: inst = 32'h10408000;
      5221: inst = 32'hc404c50;
      5222: inst = 32'h8220000;
      5223: inst = 32'h10408000;
      5224: inst = 32'hc404c51;
      5225: inst = 32'h8220000;
      5226: inst = 32'h10408000;
      5227: inst = 32'hc404c52;
      5228: inst = 32'h8220000;
      5229: inst = 32'h10408000;
      5230: inst = 32'hc404c53;
      5231: inst = 32'h8220000;
      5232: inst = 32'h10408000;
      5233: inst = 32'hc404c54;
      5234: inst = 32'h8220000;
      5235: inst = 32'h10408000;
      5236: inst = 32'hc404c55;
      5237: inst = 32'h8220000;
      5238: inst = 32'h10408000;
      5239: inst = 32'hc404c56;
      5240: inst = 32'h8220000;
      5241: inst = 32'h10408000;
      5242: inst = 32'hc404c57;
      5243: inst = 32'h8220000;
      5244: inst = 32'h10408000;
      5245: inst = 32'hc404c58;
      5246: inst = 32'h8220000;
      5247: inst = 32'h10408000;
      5248: inst = 32'hc404c59;
      5249: inst = 32'h8220000;
      5250: inst = 32'h10408000;
      5251: inst = 32'hc404c5a;
      5252: inst = 32'h8220000;
      5253: inst = 32'h10408000;
      5254: inst = 32'hc404c5b;
      5255: inst = 32'h8220000;
      5256: inst = 32'h10408000;
      5257: inst = 32'hc404c5c;
      5258: inst = 32'h8220000;
      5259: inst = 32'h10408000;
      5260: inst = 32'hc404c5d;
      5261: inst = 32'h8220000;
      5262: inst = 32'h10408000;
      5263: inst = 32'hc404c5e;
      5264: inst = 32'h8220000;
      5265: inst = 32'h10408000;
      5266: inst = 32'hc404c5f;
      5267: inst = 32'h8220000;
      5268: inst = 32'h10408000;
      5269: inst = 32'hc404c60;
      5270: inst = 32'h8220000;
      5271: inst = 32'h10408000;
      5272: inst = 32'hc404c61;
      5273: inst = 32'h8220000;
      5274: inst = 32'h10408000;
      5275: inst = 32'hc404c62;
      5276: inst = 32'h8220000;
      5277: inst = 32'h10408000;
      5278: inst = 32'hc404c63;
      5279: inst = 32'h8220000;
      5280: inst = 32'h10408000;
      5281: inst = 32'hc404c64;
      5282: inst = 32'h8220000;
      5283: inst = 32'h10408000;
      5284: inst = 32'hc404c65;
      5285: inst = 32'h8220000;
      5286: inst = 32'h10408000;
      5287: inst = 32'hc404c66;
      5288: inst = 32'h8220000;
      5289: inst = 32'h10408000;
      5290: inst = 32'hc404c67;
      5291: inst = 32'h8220000;
      5292: inst = 32'h10408000;
      5293: inst = 32'hc404c68;
      5294: inst = 32'h8220000;
      5295: inst = 32'h10408000;
      5296: inst = 32'hc404c69;
      5297: inst = 32'h8220000;
      5298: inst = 32'h10408000;
      5299: inst = 32'hc404c6a;
      5300: inst = 32'h8220000;
      5301: inst = 32'h10408000;
      5302: inst = 32'hc404c6b;
      5303: inst = 32'h8220000;
      5304: inst = 32'h10408000;
      5305: inst = 32'hc404c6c;
      5306: inst = 32'h8220000;
      5307: inst = 32'h10408000;
      5308: inst = 32'hc404c6d;
      5309: inst = 32'h8220000;
      5310: inst = 32'h10408000;
      5311: inst = 32'hc404c6e;
      5312: inst = 32'h8220000;
      5313: inst = 32'h10408000;
      5314: inst = 32'hc404c6f;
      5315: inst = 32'h8220000;
      5316: inst = 32'h10408000;
      5317: inst = 32'hc404c70;
      5318: inst = 32'h8220000;
      5319: inst = 32'h10408000;
      5320: inst = 32'hc404c71;
      5321: inst = 32'h8220000;
      5322: inst = 32'h10408000;
      5323: inst = 32'hc404c72;
      5324: inst = 32'h8220000;
      5325: inst = 32'h10408000;
      5326: inst = 32'hc404c73;
      5327: inst = 32'h8220000;
      5328: inst = 32'h10408000;
      5329: inst = 32'hc404c74;
      5330: inst = 32'h8220000;
      5331: inst = 32'h10408000;
      5332: inst = 32'hc404c75;
      5333: inst = 32'h8220000;
      5334: inst = 32'h10408000;
      5335: inst = 32'hc404c76;
      5336: inst = 32'h8220000;
      5337: inst = 32'h10408000;
      5338: inst = 32'hc404c77;
      5339: inst = 32'h8220000;
      5340: inst = 32'h10408000;
      5341: inst = 32'hc404c78;
      5342: inst = 32'h8220000;
      5343: inst = 32'h10408000;
      5344: inst = 32'hc404c79;
      5345: inst = 32'h8220000;
      5346: inst = 32'h10408000;
      5347: inst = 32'hc404c7a;
      5348: inst = 32'h8220000;
      5349: inst = 32'h10408000;
      5350: inst = 32'hc404c7b;
      5351: inst = 32'h8220000;
      5352: inst = 32'h10408000;
      5353: inst = 32'hc404c7c;
      5354: inst = 32'h8220000;
      5355: inst = 32'h10408000;
      5356: inst = 32'hc404c7d;
      5357: inst = 32'h8220000;
      5358: inst = 32'h10408000;
      5359: inst = 32'hc404c7e;
      5360: inst = 32'h8220000;
      5361: inst = 32'h10408000;
      5362: inst = 32'hc404c7f;
      5363: inst = 32'h8220000;
      5364: inst = 32'h10408000;
      5365: inst = 32'hc404c80;
      5366: inst = 32'h8220000;
      5367: inst = 32'h10408000;
      5368: inst = 32'hc404c81;
      5369: inst = 32'h8220000;
      5370: inst = 32'h10408000;
      5371: inst = 32'hc404c82;
      5372: inst = 32'h8220000;
      5373: inst = 32'h10408000;
      5374: inst = 32'hc404c83;
      5375: inst = 32'h8220000;
      5376: inst = 32'h10408000;
      5377: inst = 32'hc404c84;
      5378: inst = 32'h8220000;
      5379: inst = 32'h10408000;
      5380: inst = 32'hc404c85;
      5381: inst = 32'h8220000;
      5382: inst = 32'h10408000;
      5383: inst = 32'hc404c86;
      5384: inst = 32'h8220000;
      5385: inst = 32'h10408000;
      5386: inst = 32'hc404c87;
      5387: inst = 32'h8220000;
      5388: inst = 32'h10408000;
      5389: inst = 32'hc404c88;
      5390: inst = 32'h8220000;
      5391: inst = 32'h10408000;
      5392: inst = 32'hc404c89;
      5393: inst = 32'h8220000;
      5394: inst = 32'h10408000;
      5395: inst = 32'hc404c8a;
      5396: inst = 32'h8220000;
      5397: inst = 32'h10408000;
      5398: inst = 32'hc404c8b;
      5399: inst = 32'h8220000;
      5400: inst = 32'h10408000;
      5401: inst = 32'hc404c8c;
      5402: inst = 32'h8220000;
      5403: inst = 32'h10408000;
      5404: inst = 32'hc404c8d;
      5405: inst = 32'h8220000;
      5406: inst = 32'h10408000;
      5407: inst = 32'hc404c8e;
      5408: inst = 32'h8220000;
      5409: inst = 32'h10408000;
      5410: inst = 32'hc404ca0;
      5411: inst = 32'h8220000;
      5412: inst = 32'h10408000;
      5413: inst = 32'hc404ca1;
      5414: inst = 32'h8220000;
      5415: inst = 32'h10408000;
      5416: inst = 32'hc404cb7;
      5417: inst = 32'h8220000;
      5418: inst = 32'h10408000;
      5419: inst = 32'hc404cb8;
      5420: inst = 32'h8220000;
      5421: inst = 32'h10408000;
      5422: inst = 32'hc404cb9;
      5423: inst = 32'h8220000;
      5424: inst = 32'h10408000;
      5425: inst = 32'hc404cba;
      5426: inst = 32'h8220000;
      5427: inst = 32'h10408000;
      5428: inst = 32'hc404cbb;
      5429: inst = 32'h8220000;
      5430: inst = 32'h10408000;
      5431: inst = 32'hc404cbc;
      5432: inst = 32'h8220000;
      5433: inst = 32'h10408000;
      5434: inst = 32'hc404cbd;
      5435: inst = 32'h8220000;
      5436: inst = 32'h10408000;
      5437: inst = 32'hc404cbe;
      5438: inst = 32'h8220000;
      5439: inst = 32'h10408000;
      5440: inst = 32'hc404cbf;
      5441: inst = 32'h8220000;
      5442: inst = 32'h10408000;
      5443: inst = 32'hc404cc0;
      5444: inst = 32'h8220000;
      5445: inst = 32'h10408000;
      5446: inst = 32'hc404cc1;
      5447: inst = 32'h8220000;
      5448: inst = 32'h10408000;
      5449: inst = 32'hc404cc2;
      5450: inst = 32'h8220000;
      5451: inst = 32'h10408000;
      5452: inst = 32'hc404cc3;
      5453: inst = 32'h8220000;
      5454: inst = 32'h10408000;
      5455: inst = 32'hc404cc4;
      5456: inst = 32'h8220000;
      5457: inst = 32'h10408000;
      5458: inst = 32'hc404cc5;
      5459: inst = 32'h8220000;
      5460: inst = 32'h10408000;
      5461: inst = 32'hc404cc6;
      5462: inst = 32'h8220000;
      5463: inst = 32'h10408000;
      5464: inst = 32'hc404cc7;
      5465: inst = 32'h8220000;
      5466: inst = 32'h10408000;
      5467: inst = 32'hc404cc8;
      5468: inst = 32'h8220000;
      5469: inst = 32'h10408000;
      5470: inst = 32'hc404cc9;
      5471: inst = 32'h8220000;
      5472: inst = 32'h10408000;
      5473: inst = 32'hc404cca;
      5474: inst = 32'h8220000;
      5475: inst = 32'h10408000;
      5476: inst = 32'hc404ccb;
      5477: inst = 32'h8220000;
      5478: inst = 32'h10408000;
      5479: inst = 32'hc404ccc;
      5480: inst = 32'h8220000;
      5481: inst = 32'h10408000;
      5482: inst = 32'hc404ccd;
      5483: inst = 32'h8220000;
      5484: inst = 32'h10408000;
      5485: inst = 32'hc404cce;
      5486: inst = 32'h8220000;
      5487: inst = 32'h10408000;
      5488: inst = 32'hc404ccf;
      5489: inst = 32'h8220000;
      5490: inst = 32'h10408000;
      5491: inst = 32'hc404cd0;
      5492: inst = 32'h8220000;
      5493: inst = 32'h10408000;
      5494: inst = 32'hc404cd1;
      5495: inst = 32'h8220000;
      5496: inst = 32'h10408000;
      5497: inst = 32'hc404cd2;
      5498: inst = 32'h8220000;
      5499: inst = 32'h10408000;
      5500: inst = 32'hc404cd3;
      5501: inst = 32'h8220000;
      5502: inst = 32'h10408000;
      5503: inst = 32'hc404cd4;
      5504: inst = 32'h8220000;
      5505: inst = 32'h10408000;
      5506: inst = 32'hc404cd5;
      5507: inst = 32'h8220000;
      5508: inst = 32'h10408000;
      5509: inst = 32'hc404cd6;
      5510: inst = 32'h8220000;
      5511: inst = 32'h10408000;
      5512: inst = 32'hc404cd7;
      5513: inst = 32'h8220000;
      5514: inst = 32'h10408000;
      5515: inst = 32'hc404cd8;
      5516: inst = 32'h8220000;
      5517: inst = 32'h10408000;
      5518: inst = 32'hc404cd9;
      5519: inst = 32'h8220000;
      5520: inst = 32'h10408000;
      5521: inst = 32'hc404cda;
      5522: inst = 32'h8220000;
      5523: inst = 32'h10408000;
      5524: inst = 32'hc404cdb;
      5525: inst = 32'h8220000;
      5526: inst = 32'h10408000;
      5527: inst = 32'hc404cdc;
      5528: inst = 32'h8220000;
      5529: inst = 32'h10408000;
      5530: inst = 32'hc404cdd;
      5531: inst = 32'h8220000;
      5532: inst = 32'h10408000;
      5533: inst = 32'hc404cde;
      5534: inst = 32'h8220000;
      5535: inst = 32'h10408000;
      5536: inst = 32'hc404cdf;
      5537: inst = 32'h8220000;
      5538: inst = 32'h10408000;
      5539: inst = 32'hc404ce0;
      5540: inst = 32'h8220000;
      5541: inst = 32'h10408000;
      5542: inst = 32'hc404ce1;
      5543: inst = 32'h8220000;
      5544: inst = 32'h10408000;
      5545: inst = 32'hc404ce2;
      5546: inst = 32'h8220000;
      5547: inst = 32'h10408000;
      5548: inst = 32'hc404ce3;
      5549: inst = 32'h8220000;
      5550: inst = 32'h10408000;
      5551: inst = 32'hc404ce4;
      5552: inst = 32'h8220000;
      5553: inst = 32'h10408000;
      5554: inst = 32'hc404ce5;
      5555: inst = 32'h8220000;
      5556: inst = 32'h10408000;
      5557: inst = 32'hc404ce6;
      5558: inst = 32'h8220000;
      5559: inst = 32'h10408000;
      5560: inst = 32'hc404ce7;
      5561: inst = 32'h8220000;
      5562: inst = 32'h10408000;
      5563: inst = 32'hc404ce8;
      5564: inst = 32'h8220000;
      5565: inst = 32'h10408000;
      5566: inst = 32'hc404ce9;
      5567: inst = 32'h8220000;
      5568: inst = 32'h10408000;
      5569: inst = 32'hc404cea;
      5570: inst = 32'h8220000;
      5571: inst = 32'h10408000;
      5572: inst = 32'hc404ceb;
      5573: inst = 32'h8220000;
      5574: inst = 32'h10408000;
      5575: inst = 32'hc404cec;
      5576: inst = 32'h8220000;
      5577: inst = 32'h10408000;
      5578: inst = 32'hc404ced;
      5579: inst = 32'h8220000;
      5580: inst = 32'h10408000;
      5581: inst = 32'hc404cee;
      5582: inst = 32'h8220000;
      5583: inst = 32'h10408000;
      5584: inst = 32'hc404d17;
      5585: inst = 32'h8220000;
      5586: inst = 32'h10408000;
      5587: inst = 32'hc404d18;
      5588: inst = 32'h8220000;
      5589: inst = 32'h10408000;
      5590: inst = 32'hc404d19;
      5591: inst = 32'h8220000;
      5592: inst = 32'h10408000;
      5593: inst = 32'hc404d1a;
      5594: inst = 32'h8220000;
      5595: inst = 32'h10408000;
      5596: inst = 32'hc404d1b;
      5597: inst = 32'h8220000;
      5598: inst = 32'h10408000;
      5599: inst = 32'hc404d1c;
      5600: inst = 32'h8220000;
      5601: inst = 32'h10408000;
      5602: inst = 32'hc404d1d;
      5603: inst = 32'h8220000;
      5604: inst = 32'h10408000;
      5605: inst = 32'hc404d1e;
      5606: inst = 32'h8220000;
      5607: inst = 32'h10408000;
      5608: inst = 32'hc404d1f;
      5609: inst = 32'h8220000;
      5610: inst = 32'h10408000;
      5611: inst = 32'hc404d20;
      5612: inst = 32'h8220000;
      5613: inst = 32'h10408000;
      5614: inst = 32'hc404d21;
      5615: inst = 32'h8220000;
      5616: inst = 32'h10408000;
      5617: inst = 32'hc404d22;
      5618: inst = 32'h8220000;
      5619: inst = 32'h10408000;
      5620: inst = 32'hc404d23;
      5621: inst = 32'h8220000;
      5622: inst = 32'h10408000;
      5623: inst = 32'hc404d24;
      5624: inst = 32'h8220000;
      5625: inst = 32'h10408000;
      5626: inst = 32'hc404d25;
      5627: inst = 32'h8220000;
      5628: inst = 32'h10408000;
      5629: inst = 32'hc404d26;
      5630: inst = 32'h8220000;
      5631: inst = 32'h10408000;
      5632: inst = 32'hc404d27;
      5633: inst = 32'h8220000;
      5634: inst = 32'h10408000;
      5635: inst = 32'hc404d28;
      5636: inst = 32'h8220000;
      5637: inst = 32'h10408000;
      5638: inst = 32'hc404d29;
      5639: inst = 32'h8220000;
      5640: inst = 32'h10408000;
      5641: inst = 32'hc404d2a;
      5642: inst = 32'h8220000;
      5643: inst = 32'h10408000;
      5644: inst = 32'hc404d2b;
      5645: inst = 32'h8220000;
      5646: inst = 32'h10408000;
      5647: inst = 32'hc404d2c;
      5648: inst = 32'h8220000;
      5649: inst = 32'h10408000;
      5650: inst = 32'hc404d2d;
      5651: inst = 32'h8220000;
      5652: inst = 32'h10408000;
      5653: inst = 32'hc404d2e;
      5654: inst = 32'h8220000;
      5655: inst = 32'h10408000;
      5656: inst = 32'hc404d2f;
      5657: inst = 32'h8220000;
      5658: inst = 32'h10408000;
      5659: inst = 32'hc404d30;
      5660: inst = 32'h8220000;
      5661: inst = 32'h10408000;
      5662: inst = 32'hc404d31;
      5663: inst = 32'h8220000;
      5664: inst = 32'h10408000;
      5665: inst = 32'hc404d32;
      5666: inst = 32'h8220000;
      5667: inst = 32'h10408000;
      5668: inst = 32'hc404d33;
      5669: inst = 32'h8220000;
      5670: inst = 32'h10408000;
      5671: inst = 32'hc404d34;
      5672: inst = 32'h8220000;
      5673: inst = 32'h10408000;
      5674: inst = 32'hc404d35;
      5675: inst = 32'h8220000;
      5676: inst = 32'h10408000;
      5677: inst = 32'hc404d36;
      5678: inst = 32'h8220000;
      5679: inst = 32'h10408000;
      5680: inst = 32'hc404d37;
      5681: inst = 32'h8220000;
      5682: inst = 32'h10408000;
      5683: inst = 32'hc404d38;
      5684: inst = 32'h8220000;
      5685: inst = 32'h10408000;
      5686: inst = 32'hc404d39;
      5687: inst = 32'h8220000;
      5688: inst = 32'h10408000;
      5689: inst = 32'hc404d3a;
      5690: inst = 32'h8220000;
      5691: inst = 32'h10408000;
      5692: inst = 32'hc404d3b;
      5693: inst = 32'h8220000;
      5694: inst = 32'h10408000;
      5695: inst = 32'hc404d3c;
      5696: inst = 32'h8220000;
      5697: inst = 32'h10408000;
      5698: inst = 32'hc404d3d;
      5699: inst = 32'h8220000;
      5700: inst = 32'h10408000;
      5701: inst = 32'hc404d3e;
      5702: inst = 32'h8220000;
      5703: inst = 32'h10408000;
      5704: inst = 32'hc404d3f;
      5705: inst = 32'h8220000;
      5706: inst = 32'h10408000;
      5707: inst = 32'hc404d40;
      5708: inst = 32'h8220000;
      5709: inst = 32'h10408000;
      5710: inst = 32'hc404d41;
      5711: inst = 32'h8220000;
      5712: inst = 32'h10408000;
      5713: inst = 32'hc404d42;
      5714: inst = 32'h8220000;
      5715: inst = 32'h10408000;
      5716: inst = 32'hc404d43;
      5717: inst = 32'h8220000;
      5718: inst = 32'h10408000;
      5719: inst = 32'hc404d44;
      5720: inst = 32'h8220000;
      5721: inst = 32'h10408000;
      5722: inst = 32'hc404d45;
      5723: inst = 32'h8220000;
      5724: inst = 32'h10408000;
      5725: inst = 32'hc404d46;
      5726: inst = 32'h8220000;
      5727: inst = 32'h10408000;
      5728: inst = 32'hc404d47;
      5729: inst = 32'h8220000;
      5730: inst = 32'h10408000;
      5731: inst = 32'hc404d48;
      5732: inst = 32'h8220000;
      5733: inst = 32'h10408000;
      5734: inst = 32'hc404d49;
      5735: inst = 32'h8220000;
      5736: inst = 32'h10408000;
      5737: inst = 32'hc404d4a;
      5738: inst = 32'h8220000;
      5739: inst = 32'h10408000;
      5740: inst = 32'hc404d4b;
      5741: inst = 32'h8220000;
      5742: inst = 32'h10408000;
      5743: inst = 32'hc404d4c;
      5744: inst = 32'h8220000;
      5745: inst = 32'h10408000;
      5746: inst = 32'hc404d4d;
      5747: inst = 32'h8220000;
      5748: inst = 32'h10408000;
      5749: inst = 32'hc404d4e;
      5750: inst = 32'h8220000;
      5751: inst = 32'h10408000;
      5752: inst = 32'hc404d77;
      5753: inst = 32'h8220000;
      5754: inst = 32'h10408000;
      5755: inst = 32'hc404d78;
      5756: inst = 32'h8220000;
      5757: inst = 32'h10408000;
      5758: inst = 32'hc404d79;
      5759: inst = 32'h8220000;
      5760: inst = 32'h10408000;
      5761: inst = 32'hc404d7a;
      5762: inst = 32'h8220000;
      5763: inst = 32'h10408000;
      5764: inst = 32'hc404d7b;
      5765: inst = 32'h8220000;
      5766: inst = 32'h10408000;
      5767: inst = 32'hc404d7c;
      5768: inst = 32'h8220000;
      5769: inst = 32'h10408000;
      5770: inst = 32'hc404d7d;
      5771: inst = 32'h8220000;
      5772: inst = 32'h10408000;
      5773: inst = 32'hc404d7e;
      5774: inst = 32'h8220000;
      5775: inst = 32'h10408000;
      5776: inst = 32'hc404d7f;
      5777: inst = 32'h8220000;
      5778: inst = 32'h10408000;
      5779: inst = 32'hc404d80;
      5780: inst = 32'h8220000;
      5781: inst = 32'h10408000;
      5782: inst = 32'hc404d81;
      5783: inst = 32'h8220000;
      5784: inst = 32'h10408000;
      5785: inst = 32'hc404d82;
      5786: inst = 32'h8220000;
      5787: inst = 32'h10408000;
      5788: inst = 32'hc404d83;
      5789: inst = 32'h8220000;
      5790: inst = 32'h10408000;
      5791: inst = 32'hc404d84;
      5792: inst = 32'h8220000;
      5793: inst = 32'h10408000;
      5794: inst = 32'hc404d85;
      5795: inst = 32'h8220000;
      5796: inst = 32'h10408000;
      5797: inst = 32'hc404d86;
      5798: inst = 32'h8220000;
      5799: inst = 32'h10408000;
      5800: inst = 32'hc404d87;
      5801: inst = 32'h8220000;
      5802: inst = 32'h10408000;
      5803: inst = 32'hc404d88;
      5804: inst = 32'h8220000;
      5805: inst = 32'h10408000;
      5806: inst = 32'hc404d89;
      5807: inst = 32'h8220000;
      5808: inst = 32'h10408000;
      5809: inst = 32'hc404d8a;
      5810: inst = 32'h8220000;
      5811: inst = 32'h10408000;
      5812: inst = 32'hc404d8b;
      5813: inst = 32'h8220000;
      5814: inst = 32'h10408000;
      5815: inst = 32'hc404d8c;
      5816: inst = 32'h8220000;
      5817: inst = 32'h10408000;
      5818: inst = 32'hc404d8d;
      5819: inst = 32'h8220000;
      5820: inst = 32'h10408000;
      5821: inst = 32'hc404d8e;
      5822: inst = 32'h8220000;
      5823: inst = 32'h10408000;
      5824: inst = 32'hc404d8f;
      5825: inst = 32'h8220000;
      5826: inst = 32'h10408000;
      5827: inst = 32'hc404d90;
      5828: inst = 32'h8220000;
      5829: inst = 32'h10408000;
      5830: inst = 32'hc404d91;
      5831: inst = 32'h8220000;
      5832: inst = 32'h10408000;
      5833: inst = 32'hc404d92;
      5834: inst = 32'h8220000;
      5835: inst = 32'h10408000;
      5836: inst = 32'hc404d93;
      5837: inst = 32'h8220000;
      5838: inst = 32'h10408000;
      5839: inst = 32'hc404d94;
      5840: inst = 32'h8220000;
      5841: inst = 32'h10408000;
      5842: inst = 32'hc404d95;
      5843: inst = 32'h8220000;
      5844: inst = 32'h10408000;
      5845: inst = 32'hc404d96;
      5846: inst = 32'h8220000;
      5847: inst = 32'h10408000;
      5848: inst = 32'hc404d97;
      5849: inst = 32'h8220000;
      5850: inst = 32'h10408000;
      5851: inst = 32'hc404d98;
      5852: inst = 32'h8220000;
      5853: inst = 32'h10408000;
      5854: inst = 32'hc404d99;
      5855: inst = 32'h8220000;
      5856: inst = 32'h10408000;
      5857: inst = 32'hc404d9a;
      5858: inst = 32'h8220000;
      5859: inst = 32'h10408000;
      5860: inst = 32'hc404d9b;
      5861: inst = 32'h8220000;
      5862: inst = 32'h10408000;
      5863: inst = 32'hc404d9c;
      5864: inst = 32'h8220000;
      5865: inst = 32'h10408000;
      5866: inst = 32'hc404d9d;
      5867: inst = 32'h8220000;
      5868: inst = 32'h10408000;
      5869: inst = 32'hc404d9e;
      5870: inst = 32'h8220000;
      5871: inst = 32'h10408000;
      5872: inst = 32'hc404d9f;
      5873: inst = 32'h8220000;
      5874: inst = 32'h10408000;
      5875: inst = 32'hc404da0;
      5876: inst = 32'h8220000;
      5877: inst = 32'h10408000;
      5878: inst = 32'hc404da1;
      5879: inst = 32'h8220000;
      5880: inst = 32'h10408000;
      5881: inst = 32'hc404da2;
      5882: inst = 32'h8220000;
      5883: inst = 32'h10408000;
      5884: inst = 32'hc404da3;
      5885: inst = 32'h8220000;
      5886: inst = 32'h10408000;
      5887: inst = 32'hc404da4;
      5888: inst = 32'h8220000;
      5889: inst = 32'h10408000;
      5890: inst = 32'hc404da5;
      5891: inst = 32'h8220000;
      5892: inst = 32'h10408000;
      5893: inst = 32'hc404da6;
      5894: inst = 32'h8220000;
      5895: inst = 32'h10408000;
      5896: inst = 32'hc404da7;
      5897: inst = 32'h8220000;
      5898: inst = 32'h10408000;
      5899: inst = 32'hc404da8;
      5900: inst = 32'h8220000;
      5901: inst = 32'h10408000;
      5902: inst = 32'hc404da9;
      5903: inst = 32'h8220000;
      5904: inst = 32'h10408000;
      5905: inst = 32'hc404daa;
      5906: inst = 32'h8220000;
      5907: inst = 32'h10408000;
      5908: inst = 32'hc404dab;
      5909: inst = 32'h8220000;
      5910: inst = 32'h10408000;
      5911: inst = 32'hc404dac;
      5912: inst = 32'h8220000;
      5913: inst = 32'h10408000;
      5914: inst = 32'hc404dad;
      5915: inst = 32'h8220000;
      5916: inst = 32'h10408000;
      5917: inst = 32'hc404dae;
      5918: inst = 32'h8220000;
      5919: inst = 32'h10408000;
      5920: inst = 32'hc404dd7;
      5921: inst = 32'h8220000;
      5922: inst = 32'h10408000;
      5923: inst = 32'hc404dd8;
      5924: inst = 32'h8220000;
      5925: inst = 32'h10408000;
      5926: inst = 32'hc404dd9;
      5927: inst = 32'h8220000;
      5928: inst = 32'h10408000;
      5929: inst = 32'hc404dda;
      5930: inst = 32'h8220000;
      5931: inst = 32'h10408000;
      5932: inst = 32'hc404ddb;
      5933: inst = 32'h8220000;
      5934: inst = 32'h10408000;
      5935: inst = 32'hc404ddc;
      5936: inst = 32'h8220000;
      5937: inst = 32'h10408000;
      5938: inst = 32'hc404ddd;
      5939: inst = 32'h8220000;
      5940: inst = 32'h10408000;
      5941: inst = 32'hc404dde;
      5942: inst = 32'h8220000;
      5943: inst = 32'h10408000;
      5944: inst = 32'hc404ddf;
      5945: inst = 32'h8220000;
      5946: inst = 32'h10408000;
      5947: inst = 32'hc404de0;
      5948: inst = 32'h8220000;
      5949: inst = 32'h10408000;
      5950: inst = 32'hc404de1;
      5951: inst = 32'h8220000;
      5952: inst = 32'h10408000;
      5953: inst = 32'hc404de2;
      5954: inst = 32'h8220000;
      5955: inst = 32'h10408000;
      5956: inst = 32'hc404de3;
      5957: inst = 32'h8220000;
      5958: inst = 32'h10408000;
      5959: inst = 32'hc404de4;
      5960: inst = 32'h8220000;
      5961: inst = 32'h10408000;
      5962: inst = 32'hc404de5;
      5963: inst = 32'h8220000;
      5964: inst = 32'h10408000;
      5965: inst = 32'hc404de6;
      5966: inst = 32'h8220000;
      5967: inst = 32'h10408000;
      5968: inst = 32'hc404de7;
      5969: inst = 32'h8220000;
      5970: inst = 32'h10408000;
      5971: inst = 32'hc404de8;
      5972: inst = 32'h8220000;
      5973: inst = 32'h10408000;
      5974: inst = 32'hc404de9;
      5975: inst = 32'h8220000;
      5976: inst = 32'h10408000;
      5977: inst = 32'hc404dea;
      5978: inst = 32'h8220000;
      5979: inst = 32'h10408000;
      5980: inst = 32'hc404deb;
      5981: inst = 32'h8220000;
      5982: inst = 32'h10408000;
      5983: inst = 32'hc404dec;
      5984: inst = 32'h8220000;
      5985: inst = 32'h10408000;
      5986: inst = 32'hc404ded;
      5987: inst = 32'h8220000;
      5988: inst = 32'h10408000;
      5989: inst = 32'hc404dee;
      5990: inst = 32'h8220000;
      5991: inst = 32'h10408000;
      5992: inst = 32'hc404def;
      5993: inst = 32'h8220000;
      5994: inst = 32'h10408000;
      5995: inst = 32'hc404df0;
      5996: inst = 32'h8220000;
      5997: inst = 32'h10408000;
      5998: inst = 32'hc404df1;
      5999: inst = 32'h8220000;
      6000: inst = 32'h10408000;
      6001: inst = 32'hc404df2;
      6002: inst = 32'h8220000;
      6003: inst = 32'h10408000;
      6004: inst = 32'hc404df3;
      6005: inst = 32'h8220000;
      6006: inst = 32'h10408000;
      6007: inst = 32'hc404df4;
      6008: inst = 32'h8220000;
      6009: inst = 32'h10408000;
      6010: inst = 32'hc404df5;
      6011: inst = 32'h8220000;
      6012: inst = 32'h10408000;
      6013: inst = 32'hc404df6;
      6014: inst = 32'h8220000;
      6015: inst = 32'h10408000;
      6016: inst = 32'hc404df7;
      6017: inst = 32'h8220000;
      6018: inst = 32'h10408000;
      6019: inst = 32'hc404df8;
      6020: inst = 32'h8220000;
      6021: inst = 32'h10408000;
      6022: inst = 32'hc404df9;
      6023: inst = 32'h8220000;
      6024: inst = 32'h10408000;
      6025: inst = 32'hc404dfa;
      6026: inst = 32'h8220000;
      6027: inst = 32'h10408000;
      6028: inst = 32'hc404dfb;
      6029: inst = 32'h8220000;
      6030: inst = 32'h10408000;
      6031: inst = 32'hc404dfc;
      6032: inst = 32'h8220000;
      6033: inst = 32'h10408000;
      6034: inst = 32'hc404dfd;
      6035: inst = 32'h8220000;
      6036: inst = 32'h10408000;
      6037: inst = 32'hc404dfe;
      6038: inst = 32'h8220000;
      6039: inst = 32'h10408000;
      6040: inst = 32'hc404dff;
      6041: inst = 32'h8220000;
      6042: inst = 32'h10408000;
      6043: inst = 32'hc404e00;
      6044: inst = 32'h8220000;
      6045: inst = 32'h10408000;
      6046: inst = 32'hc404e01;
      6047: inst = 32'h8220000;
      6048: inst = 32'h10408000;
      6049: inst = 32'hc404e02;
      6050: inst = 32'h8220000;
      6051: inst = 32'h10408000;
      6052: inst = 32'hc404e03;
      6053: inst = 32'h8220000;
      6054: inst = 32'h10408000;
      6055: inst = 32'hc404e04;
      6056: inst = 32'h8220000;
      6057: inst = 32'h10408000;
      6058: inst = 32'hc404e05;
      6059: inst = 32'h8220000;
      6060: inst = 32'h10408000;
      6061: inst = 32'hc404e06;
      6062: inst = 32'h8220000;
      6063: inst = 32'h10408000;
      6064: inst = 32'hc404e07;
      6065: inst = 32'h8220000;
      6066: inst = 32'h10408000;
      6067: inst = 32'hc404e08;
      6068: inst = 32'h8220000;
      6069: inst = 32'h10408000;
      6070: inst = 32'hc404e09;
      6071: inst = 32'h8220000;
      6072: inst = 32'h10408000;
      6073: inst = 32'hc404e0a;
      6074: inst = 32'h8220000;
      6075: inst = 32'h10408000;
      6076: inst = 32'hc404e0b;
      6077: inst = 32'h8220000;
      6078: inst = 32'h10408000;
      6079: inst = 32'hc404e0c;
      6080: inst = 32'h8220000;
      6081: inst = 32'h10408000;
      6082: inst = 32'hc404e0d;
      6083: inst = 32'h8220000;
      6084: inst = 32'h10408000;
      6085: inst = 32'hc404e0e;
      6086: inst = 32'h8220000;
      6087: inst = 32'h10408000;
      6088: inst = 32'hc404e37;
      6089: inst = 32'h8220000;
      6090: inst = 32'h10408000;
      6091: inst = 32'hc404e38;
      6092: inst = 32'h8220000;
      6093: inst = 32'h10408000;
      6094: inst = 32'hc404e39;
      6095: inst = 32'h8220000;
      6096: inst = 32'h10408000;
      6097: inst = 32'hc404e3a;
      6098: inst = 32'h8220000;
      6099: inst = 32'h10408000;
      6100: inst = 32'hc404e3b;
      6101: inst = 32'h8220000;
      6102: inst = 32'h10408000;
      6103: inst = 32'hc404e3c;
      6104: inst = 32'h8220000;
      6105: inst = 32'h10408000;
      6106: inst = 32'hc404e3d;
      6107: inst = 32'h8220000;
      6108: inst = 32'h10408000;
      6109: inst = 32'hc404e3e;
      6110: inst = 32'h8220000;
      6111: inst = 32'h10408000;
      6112: inst = 32'hc404e3f;
      6113: inst = 32'h8220000;
      6114: inst = 32'h10408000;
      6115: inst = 32'hc404e40;
      6116: inst = 32'h8220000;
      6117: inst = 32'h10408000;
      6118: inst = 32'hc404e41;
      6119: inst = 32'h8220000;
      6120: inst = 32'h10408000;
      6121: inst = 32'hc404e42;
      6122: inst = 32'h8220000;
      6123: inst = 32'h10408000;
      6124: inst = 32'hc404e43;
      6125: inst = 32'h8220000;
      6126: inst = 32'h10408000;
      6127: inst = 32'hc404e44;
      6128: inst = 32'h8220000;
      6129: inst = 32'h10408000;
      6130: inst = 32'hc404e45;
      6131: inst = 32'h8220000;
      6132: inst = 32'h10408000;
      6133: inst = 32'hc404e46;
      6134: inst = 32'h8220000;
      6135: inst = 32'h10408000;
      6136: inst = 32'hc404e47;
      6137: inst = 32'h8220000;
      6138: inst = 32'h10408000;
      6139: inst = 32'hc404e48;
      6140: inst = 32'h8220000;
      6141: inst = 32'h10408000;
      6142: inst = 32'hc404e49;
      6143: inst = 32'h8220000;
      6144: inst = 32'h10408000;
      6145: inst = 32'hc404e4a;
      6146: inst = 32'h8220000;
      6147: inst = 32'h10408000;
      6148: inst = 32'hc404e4b;
      6149: inst = 32'h8220000;
      6150: inst = 32'h10408000;
      6151: inst = 32'hc404e4c;
      6152: inst = 32'h8220000;
      6153: inst = 32'h10408000;
      6154: inst = 32'hc404e4d;
      6155: inst = 32'h8220000;
      6156: inst = 32'h10408000;
      6157: inst = 32'hc404e4e;
      6158: inst = 32'h8220000;
      6159: inst = 32'h10408000;
      6160: inst = 32'hc404e4f;
      6161: inst = 32'h8220000;
      6162: inst = 32'h10408000;
      6163: inst = 32'hc404e50;
      6164: inst = 32'h8220000;
      6165: inst = 32'h10408000;
      6166: inst = 32'hc404e51;
      6167: inst = 32'h8220000;
      6168: inst = 32'h10408000;
      6169: inst = 32'hc404e52;
      6170: inst = 32'h8220000;
      6171: inst = 32'h10408000;
      6172: inst = 32'hc404e53;
      6173: inst = 32'h8220000;
      6174: inst = 32'h10408000;
      6175: inst = 32'hc404e54;
      6176: inst = 32'h8220000;
      6177: inst = 32'h10408000;
      6178: inst = 32'hc404e55;
      6179: inst = 32'h8220000;
      6180: inst = 32'h10408000;
      6181: inst = 32'hc404e56;
      6182: inst = 32'h8220000;
      6183: inst = 32'h10408000;
      6184: inst = 32'hc404e57;
      6185: inst = 32'h8220000;
      6186: inst = 32'h10408000;
      6187: inst = 32'hc404e58;
      6188: inst = 32'h8220000;
      6189: inst = 32'h10408000;
      6190: inst = 32'hc404e59;
      6191: inst = 32'h8220000;
      6192: inst = 32'h10408000;
      6193: inst = 32'hc404e5a;
      6194: inst = 32'h8220000;
      6195: inst = 32'h10408000;
      6196: inst = 32'hc404e5b;
      6197: inst = 32'h8220000;
      6198: inst = 32'h10408000;
      6199: inst = 32'hc404e5c;
      6200: inst = 32'h8220000;
      6201: inst = 32'h10408000;
      6202: inst = 32'hc404e5d;
      6203: inst = 32'h8220000;
      6204: inst = 32'h10408000;
      6205: inst = 32'hc404e5e;
      6206: inst = 32'h8220000;
      6207: inst = 32'h10408000;
      6208: inst = 32'hc404e5f;
      6209: inst = 32'h8220000;
      6210: inst = 32'h10408000;
      6211: inst = 32'hc404e60;
      6212: inst = 32'h8220000;
      6213: inst = 32'h10408000;
      6214: inst = 32'hc404e61;
      6215: inst = 32'h8220000;
      6216: inst = 32'h10408000;
      6217: inst = 32'hc404e62;
      6218: inst = 32'h8220000;
      6219: inst = 32'h10408000;
      6220: inst = 32'hc404e63;
      6221: inst = 32'h8220000;
      6222: inst = 32'h10408000;
      6223: inst = 32'hc404e64;
      6224: inst = 32'h8220000;
      6225: inst = 32'h10408000;
      6226: inst = 32'hc404e65;
      6227: inst = 32'h8220000;
      6228: inst = 32'h10408000;
      6229: inst = 32'hc404e66;
      6230: inst = 32'h8220000;
      6231: inst = 32'h10408000;
      6232: inst = 32'hc404e67;
      6233: inst = 32'h8220000;
      6234: inst = 32'h10408000;
      6235: inst = 32'hc404e68;
      6236: inst = 32'h8220000;
      6237: inst = 32'h10408000;
      6238: inst = 32'hc404e69;
      6239: inst = 32'h8220000;
      6240: inst = 32'h10408000;
      6241: inst = 32'hc404e6a;
      6242: inst = 32'h8220000;
      6243: inst = 32'h10408000;
      6244: inst = 32'hc404e6b;
      6245: inst = 32'h8220000;
      6246: inst = 32'h10408000;
      6247: inst = 32'hc404e6c;
      6248: inst = 32'h8220000;
      6249: inst = 32'h10408000;
      6250: inst = 32'hc404e6d;
      6251: inst = 32'h8220000;
      6252: inst = 32'h10408000;
      6253: inst = 32'hc404e6e;
      6254: inst = 32'h8220000;
      6255: inst = 32'h10408000;
      6256: inst = 32'hc404e97;
      6257: inst = 32'h8220000;
      6258: inst = 32'h10408000;
      6259: inst = 32'hc404e98;
      6260: inst = 32'h8220000;
      6261: inst = 32'h10408000;
      6262: inst = 32'hc404e99;
      6263: inst = 32'h8220000;
      6264: inst = 32'h10408000;
      6265: inst = 32'hc404e9a;
      6266: inst = 32'h8220000;
      6267: inst = 32'h10408000;
      6268: inst = 32'hc404e9b;
      6269: inst = 32'h8220000;
      6270: inst = 32'h10408000;
      6271: inst = 32'hc404e9c;
      6272: inst = 32'h8220000;
      6273: inst = 32'h10408000;
      6274: inst = 32'hc404e9d;
      6275: inst = 32'h8220000;
      6276: inst = 32'h10408000;
      6277: inst = 32'hc404e9e;
      6278: inst = 32'h8220000;
      6279: inst = 32'h10408000;
      6280: inst = 32'hc404ea8;
      6281: inst = 32'h8220000;
      6282: inst = 32'h10408000;
      6283: inst = 32'hc404ea9;
      6284: inst = 32'h8220000;
      6285: inst = 32'h10408000;
      6286: inst = 32'hc404eaa;
      6287: inst = 32'h8220000;
      6288: inst = 32'h10408000;
      6289: inst = 32'hc404eab;
      6290: inst = 32'h8220000;
      6291: inst = 32'h10408000;
      6292: inst = 32'hc404eac;
      6293: inst = 32'h8220000;
      6294: inst = 32'h10408000;
      6295: inst = 32'hc404ead;
      6296: inst = 32'h8220000;
      6297: inst = 32'h10408000;
      6298: inst = 32'hc404eae;
      6299: inst = 32'h8220000;
      6300: inst = 32'h10408000;
      6301: inst = 32'hc404eaf;
      6302: inst = 32'h8220000;
      6303: inst = 32'h10408000;
      6304: inst = 32'hc404eb0;
      6305: inst = 32'h8220000;
      6306: inst = 32'h10408000;
      6307: inst = 32'hc404eb1;
      6308: inst = 32'h8220000;
      6309: inst = 32'h10408000;
      6310: inst = 32'hc404eb2;
      6311: inst = 32'h8220000;
      6312: inst = 32'h10408000;
      6313: inst = 32'hc404eb3;
      6314: inst = 32'h8220000;
      6315: inst = 32'h10408000;
      6316: inst = 32'hc404eb4;
      6317: inst = 32'h8220000;
      6318: inst = 32'h10408000;
      6319: inst = 32'hc404eb5;
      6320: inst = 32'h8220000;
      6321: inst = 32'h10408000;
      6322: inst = 32'hc404eb6;
      6323: inst = 32'h8220000;
      6324: inst = 32'h10408000;
      6325: inst = 32'hc404eb7;
      6326: inst = 32'h8220000;
      6327: inst = 32'h10408000;
      6328: inst = 32'hc404ec1;
      6329: inst = 32'h8220000;
      6330: inst = 32'h10408000;
      6331: inst = 32'hc404ec2;
      6332: inst = 32'h8220000;
      6333: inst = 32'h10408000;
      6334: inst = 32'hc404ec3;
      6335: inst = 32'h8220000;
      6336: inst = 32'h10408000;
      6337: inst = 32'hc404ec4;
      6338: inst = 32'h8220000;
      6339: inst = 32'h10408000;
      6340: inst = 32'hc404ec5;
      6341: inst = 32'h8220000;
      6342: inst = 32'h10408000;
      6343: inst = 32'hc404ec6;
      6344: inst = 32'h8220000;
      6345: inst = 32'h10408000;
      6346: inst = 32'hc404ec7;
      6347: inst = 32'h8220000;
      6348: inst = 32'h10408000;
      6349: inst = 32'hc404ec8;
      6350: inst = 32'h8220000;
      6351: inst = 32'h10408000;
      6352: inst = 32'hc404ec9;
      6353: inst = 32'h8220000;
      6354: inst = 32'h10408000;
      6355: inst = 32'hc404eca;
      6356: inst = 32'h8220000;
      6357: inst = 32'h10408000;
      6358: inst = 32'hc404ecb;
      6359: inst = 32'h8220000;
      6360: inst = 32'h10408000;
      6361: inst = 32'hc404ecc;
      6362: inst = 32'h8220000;
      6363: inst = 32'h10408000;
      6364: inst = 32'hc404ecd;
      6365: inst = 32'h8220000;
      6366: inst = 32'h10408000;
      6367: inst = 32'hc404ece;
      6368: inst = 32'h8220000;
      6369: inst = 32'h10408000;
      6370: inst = 32'hc404ef7;
      6371: inst = 32'h8220000;
      6372: inst = 32'h10408000;
      6373: inst = 32'hc404ef8;
      6374: inst = 32'h8220000;
      6375: inst = 32'h10408000;
      6376: inst = 32'hc404ef9;
      6377: inst = 32'h8220000;
      6378: inst = 32'h10408000;
      6379: inst = 32'hc404efa;
      6380: inst = 32'h8220000;
      6381: inst = 32'h10408000;
      6382: inst = 32'hc404efb;
      6383: inst = 32'h8220000;
      6384: inst = 32'h10408000;
      6385: inst = 32'hc404efc;
      6386: inst = 32'h8220000;
      6387: inst = 32'h10408000;
      6388: inst = 32'hc404efd;
      6389: inst = 32'h8220000;
      6390: inst = 32'h10408000;
      6391: inst = 32'hc404efe;
      6392: inst = 32'h8220000;
      6393: inst = 32'h10408000;
      6394: inst = 32'hc404f08;
      6395: inst = 32'h8220000;
      6396: inst = 32'h10408000;
      6397: inst = 32'hc404f09;
      6398: inst = 32'h8220000;
      6399: inst = 32'h10408000;
      6400: inst = 32'hc404f0a;
      6401: inst = 32'h8220000;
      6402: inst = 32'h10408000;
      6403: inst = 32'hc404f0b;
      6404: inst = 32'h8220000;
      6405: inst = 32'h10408000;
      6406: inst = 32'hc404f0c;
      6407: inst = 32'h8220000;
      6408: inst = 32'h10408000;
      6409: inst = 32'hc404f0d;
      6410: inst = 32'h8220000;
      6411: inst = 32'h10408000;
      6412: inst = 32'hc404f0e;
      6413: inst = 32'h8220000;
      6414: inst = 32'h10408000;
      6415: inst = 32'hc404f0f;
      6416: inst = 32'h8220000;
      6417: inst = 32'h10408000;
      6418: inst = 32'hc404f10;
      6419: inst = 32'h8220000;
      6420: inst = 32'h10408000;
      6421: inst = 32'hc404f11;
      6422: inst = 32'h8220000;
      6423: inst = 32'h10408000;
      6424: inst = 32'hc404f12;
      6425: inst = 32'h8220000;
      6426: inst = 32'h10408000;
      6427: inst = 32'hc404f13;
      6428: inst = 32'h8220000;
      6429: inst = 32'h10408000;
      6430: inst = 32'hc404f14;
      6431: inst = 32'h8220000;
      6432: inst = 32'h10408000;
      6433: inst = 32'hc404f15;
      6434: inst = 32'h8220000;
      6435: inst = 32'h10408000;
      6436: inst = 32'hc404f16;
      6437: inst = 32'h8220000;
      6438: inst = 32'h10408000;
      6439: inst = 32'hc404f17;
      6440: inst = 32'h8220000;
      6441: inst = 32'h10408000;
      6442: inst = 32'hc404f21;
      6443: inst = 32'h8220000;
      6444: inst = 32'h10408000;
      6445: inst = 32'hc404f22;
      6446: inst = 32'h8220000;
      6447: inst = 32'h10408000;
      6448: inst = 32'hc404f23;
      6449: inst = 32'h8220000;
      6450: inst = 32'h10408000;
      6451: inst = 32'hc404f24;
      6452: inst = 32'h8220000;
      6453: inst = 32'h10408000;
      6454: inst = 32'hc404f25;
      6455: inst = 32'h8220000;
      6456: inst = 32'h10408000;
      6457: inst = 32'hc404f26;
      6458: inst = 32'h8220000;
      6459: inst = 32'h10408000;
      6460: inst = 32'hc404f27;
      6461: inst = 32'h8220000;
      6462: inst = 32'h10408000;
      6463: inst = 32'hc404f28;
      6464: inst = 32'h8220000;
      6465: inst = 32'h10408000;
      6466: inst = 32'hc404f29;
      6467: inst = 32'h8220000;
      6468: inst = 32'h10408000;
      6469: inst = 32'hc404f2a;
      6470: inst = 32'h8220000;
      6471: inst = 32'h10408000;
      6472: inst = 32'hc404f2b;
      6473: inst = 32'h8220000;
      6474: inst = 32'h10408000;
      6475: inst = 32'hc404f2c;
      6476: inst = 32'h8220000;
      6477: inst = 32'h10408000;
      6478: inst = 32'hc404f2d;
      6479: inst = 32'h8220000;
      6480: inst = 32'h10408000;
      6481: inst = 32'hc404f2e;
      6482: inst = 32'h8220000;
      6483: inst = 32'h10408000;
      6484: inst = 32'hc404f57;
      6485: inst = 32'h8220000;
      6486: inst = 32'h10408000;
      6487: inst = 32'hc404f58;
      6488: inst = 32'h8220000;
      6489: inst = 32'h10408000;
      6490: inst = 32'hc404f59;
      6491: inst = 32'h8220000;
      6492: inst = 32'h10408000;
      6493: inst = 32'hc404f5a;
      6494: inst = 32'h8220000;
      6495: inst = 32'h10408000;
      6496: inst = 32'hc404f5b;
      6497: inst = 32'h8220000;
      6498: inst = 32'h10408000;
      6499: inst = 32'hc404f5c;
      6500: inst = 32'h8220000;
      6501: inst = 32'h10408000;
      6502: inst = 32'hc404f5d;
      6503: inst = 32'h8220000;
      6504: inst = 32'h10408000;
      6505: inst = 32'hc404f5e;
      6506: inst = 32'h8220000;
      6507: inst = 32'h10408000;
      6508: inst = 32'hc404f68;
      6509: inst = 32'h8220000;
      6510: inst = 32'h10408000;
      6511: inst = 32'hc404f69;
      6512: inst = 32'h8220000;
      6513: inst = 32'h10408000;
      6514: inst = 32'hc404f6a;
      6515: inst = 32'h8220000;
      6516: inst = 32'h10408000;
      6517: inst = 32'hc404f6b;
      6518: inst = 32'h8220000;
      6519: inst = 32'h10408000;
      6520: inst = 32'hc404f6c;
      6521: inst = 32'h8220000;
      6522: inst = 32'h10408000;
      6523: inst = 32'hc404f6d;
      6524: inst = 32'h8220000;
      6525: inst = 32'h10408000;
      6526: inst = 32'hc404f6e;
      6527: inst = 32'h8220000;
      6528: inst = 32'h10408000;
      6529: inst = 32'hc404f6f;
      6530: inst = 32'h8220000;
      6531: inst = 32'h10408000;
      6532: inst = 32'hc404f70;
      6533: inst = 32'h8220000;
      6534: inst = 32'h10408000;
      6535: inst = 32'hc404f71;
      6536: inst = 32'h8220000;
      6537: inst = 32'h10408000;
      6538: inst = 32'hc404f72;
      6539: inst = 32'h8220000;
      6540: inst = 32'h10408000;
      6541: inst = 32'hc404f73;
      6542: inst = 32'h8220000;
      6543: inst = 32'h10408000;
      6544: inst = 32'hc404f74;
      6545: inst = 32'h8220000;
      6546: inst = 32'h10408000;
      6547: inst = 32'hc404f75;
      6548: inst = 32'h8220000;
      6549: inst = 32'h10408000;
      6550: inst = 32'hc404f76;
      6551: inst = 32'h8220000;
      6552: inst = 32'h10408000;
      6553: inst = 32'hc404f77;
      6554: inst = 32'h8220000;
      6555: inst = 32'h10408000;
      6556: inst = 32'hc404f81;
      6557: inst = 32'h8220000;
      6558: inst = 32'h10408000;
      6559: inst = 32'hc404f82;
      6560: inst = 32'h8220000;
      6561: inst = 32'h10408000;
      6562: inst = 32'hc404f83;
      6563: inst = 32'h8220000;
      6564: inst = 32'h10408000;
      6565: inst = 32'hc404f84;
      6566: inst = 32'h8220000;
      6567: inst = 32'h10408000;
      6568: inst = 32'hc404f85;
      6569: inst = 32'h8220000;
      6570: inst = 32'h10408000;
      6571: inst = 32'hc404f86;
      6572: inst = 32'h8220000;
      6573: inst = 32'h10408000;
      6574: inst = 32'hc404f87;
      6575: inst = 32'h8220000;
      6576: inst = 32'h10408000;
      6577: inst = 32'hc404f88;
      6578: inst = 32'h8220000;
      6579: inst = 32'h10408000;
      6580: inst = 32'hc404f89;
      6581: inst = 32'h8220000;
      6582: inst = 32'h10408000;
      6583: inst = 32'hc404f8a;
      6584: inst = 32'h8220000;
      6585: inst = 32'h10408000;
      6586: inst = 32'hc404f8b;
      6587: inst = 32'h8220000;
      6588: inst = 32'h10408000;
      6589: inst = 32'hc404f8c;
      6590: inst = 32'h8220000;
      6591: inst = 32'h10408000;
      6592: inst = 32'hc404f8d;
      6593: inst = 32'h8220000;
      6594: inst = 32'h10408000;
      6595: inst = 32'hc404f8e;
      6596: inst = 32'h8220000;
      6597: inst = 32'h10408000;
      6598: inst = 32'hc404fb7;
      6599: inst = 32'h8220000;
      6600: inst = 32'h10408000;
      6601: inst = 32'hc404fb8;
      6602: inst = 32'h8220000;
      6603: inst = 32'h10408000;
      6604: inst = 32'hc404fb9;
      6605: inst = 32'h8220000;
      6606: inst = 32'h10408000;
      6607: inst = 32'hc404fba;
      6608: inst = 32'h8220000;
      6609: inst = 32'h10408000;
      6610: inst = 32'hc404fbb;
      6611: inst = 32'h8220000;
      6612: inst = 32'h10408000;
      6613: inst = 32'hc404fbc;
      6614: inst = 32'h8220000;
      6615: inst = 32'h10408000;
      6616: inst = 32'hc404fbd;
      6617: inst = 32'h8220000;
      6618: inst = 32'h10408000;
      6619: inst = 32'hc404fbe;
      6620: inst = 32'h8220000;
      6621: inst = 32'h10408000;
      6622: inst = 32'hc404fc8;
      6623: inst = 32'h8220000;
      6624: inst = 32'h10408000;
      6625: inst = 32'hc404fc9;
      6626: inst = 32'h8220000;
      6627: inst = 32'h10408000;
      6628: inst = 32'hc404fca;
      6629: inst = 32'h8220000;
      6630: inst = 32'h10408000;
      6631: inst = 32'hc404fcb;
      6632: inst = 32'h8220000;
      6633: inst = 32'h10408000;
      6634: inst = 32'hc404fcc;
      6635: inst = 32'h8220000;
      6636: inst = 32'h10408000;
      6637: inst = 32'hc404fcd;
      6638: inst = 32'h8220000;
      6639: inst = 32'h10408000;
      6640: inst = 32'hc404fce;
      6641: inst = 32'h8220000;
      6642: inst = 32'h10408000;
      6643: inst = 32'hc404fcf;
      6644: inst = 32'h8220000;
      6645: inst = 32'h10408000;
      6646: inst = 32'hc404fd0;
      6647: inst = 32'h8220000;
      6648: inst = 32'h10408000;
      6649: inst = 32'hc404fd1;
      6650: inst = 32'h8220000;
      6651: inst = 32'h10408000;
      6652: inst = 32'hc404fd2;
      6653: inst = 32'h8220000;
      6654: inst = 32'h10408000;
      6655: inst = 32'hc404fd3;
      6656: inst = 32'h8220000;
      6657: inst = 32'h10408000;
      6658: inst = 32'hc404fd4;
      6659: inst = 32'h8220000;
      6660: inst = 32'h10408000;
      6661: inst = 32'hc404fd5;
      6662: inst = 32'h8220000;
      6663: inst = 32'h10408000;
      6664: inst = 32'hc404fd6;
      6665: inst = 32'h8220000;
      6666: inst = 32'h10408000;
      6667: inst = 32'hc404fd7;
      6668: inst = 32'h8220000;
      6669: inst = 32'h10408000;
      6670: inst = 32'hc404fe1;
      6671: inst = 32'h8220000;
      6672: inst = 32'h10408000;
      6673: inst = 32'hc404fe2;
      6674: inst = 32'h8220000;
      6675: inst = 32'h10408000;
      6676: inst = 32'hc404fe3;
      6677: inst = 32'h8220000;
      6678: inst = 32'h10408000;
      6679: inst = 32'hc404fe4;
      6680: inst = 32'h8220000;
      6681: inst = 32'h10408000;
      6682: inst = 32'hc404fe5;
      6683: inst = 32'h8220000;
      6684: inst = 32'h10408000;
      6685: inst = 32'hc404fe6;
      6686: inst = 32'h8220000;
      6687: inst = 32'h10408000;
      6688: inst = 32'hc404fe7;
      6689: inst = 32'h8220000;
      6690: inst = 32'h10408000;
      6691: inst = 32'hc404fe8;
      6692: inst = 32'h8220000;
      6693: inst = 32'h10408000;
      6694: inst = 32'hc404fe9;
      6695: inst = 32'h8220000;
      6696: inst = 32'h10408000;
      6697: inst = 32'hc404fea;
      6698: inst = 32'h8220000;
      6699: inst = 32'h10408000;
      6700: inst = 32'hc404feb;
      6701: inst = 32'h8220000;
      6702: inst = 32'h10408000;
      6703: inst = 32'hc404fec;
      6704: inst = 32'h8220000;
      6705: inst = 32'h10408000;
      6706: inst = 32'hc404fed;
      6707: inst = 32'h8220000;
      6708: inst = 32'h10408000;
      6709: inst = 32'hc404fee;
      6710: inst = 32'h8220000;
      6711: inst = 32'h10408000;
      6712: inst = 32'hc405017;
      6713: inst = 32'h8220000;
      6714: inst = 32'h10408000;
      6715: inst = 32'hc405018;
      6716: inst = 32'h8220000;
      6717: inst = 32'h10408000;
      6718: inst = 32'hc405019;
      6719: inst = 32'h8220000;
      6720: inst = 32'h10408000;
      6721: inst = 32'hc40501a;
      6722: inst = 32'h8220000;
      6723: inst = 32'h10408000;
      6724: inst = 32'hc40501b;
      6725: inst = 32'h8220000;
      6726: inst = 32'h10408000;
      6727: inst = 32'hc40501c;
      6728: inst = 32'h8220000;
      6729: inst = 32'h10408000;
      6730: inst = 32'hc40501d;
      6731: inst = 32'h8220000;
      6732: inst = 32'h10408000;
      6733: inst = 32'hc40501e;
      6734: inst = 32'h8220000;
      6735: inst = 32'h10408000;
      6736: inst = 32'hc405028;
      6737: inst = 32'h8220000;
      6738: inst = 32'h10408000;
      6739: inst = 32'hc405029;
      6740: inst = 32'h8220000;
      6741: inst = 32'h10408000;
      6742: inst = 32'hc40502a;
      6743: inst = 32'h8220000;
      6744: inst = 32'h10408000;
      6745: inst = 32'hc40502b;
      6746: inst = 32'h8220000;
      6747: inst = 32'h10408000;
      6748: inst = 32'hc40502c;
      6749: inst = 32'h8220000;
      6750: inst = 32'h10408000;
      6751: inst = 32'hc40502d;
      6752: inst = 32'h8220000;
      6753: inst = 32'h10408000;
      6754: inst = 32'hc40502e;
      6755: inst = 32'h8220000;
      6756: inst = 32'h10408000;
      6757: inst = 32'hc40502f;
      6758: inst = 32'h8220000;
      6759: inst = 32'h10408000;
      6760: inst = 32'hc405030;
      6761: inst = 32'h8220000;
      6762: inst = 32'h10408000;
      6763: inst = 32'hc405031;
      6764: inst = 32'h8220000;
      6765: inst = 32'h10408000;
      6766: inst = 32'hc405032;
      6767: inst = 32'h8220000;
      6768: inst = 32'h10408000;
      6769: inst = 32'hc405033;
      6770: inst = 32'h8220000;
      6771: inst = 32'h10408000;
      6772: inst = 32'hc405034;
      6773: inst = 32'h8220000;
      6774: inst = 32'h10408000;
      6775: inst = 32'hc405035;
      6776: inst = 32'h8220000;
      6777: inst = 32'h10408000;
      6778: inst = 32'hc405036;
      6779: inst = 32'h8220000;
      6780: inst = 32'h10408000;
      6781: inst = 32'hc405037;
      6782: inst = 32'h8220000;
      6783: inst = 32'h10408000;
      6784: inst = 32'hc405041;
      6785: inst = 32'h8220000;
      6786: inst = 32'h10408000;
      6787: inst = 32'hc405042;
      6788: inst = 32'h8220000;
      6789: inst = 32'h10408000;
      6790: inst = 32'hc405043;
      6791: inst = 32'h8220000;
      6792: inst = 32'h10408000;
      6793: inst = 32'hc405044;
      6794: inst = 32'h8220000;
      6795: inst = 32'h10408000;
      6796: inst = 32'hc405045;
      6797: inst = 32'h8220000;
      6798: inst = 32'h10408000;
      6799: inst = 32'hc405046;
      6800: inst = 32'h8220000;
      6801: inst = 32'h10408000;
      6802: inst = 32'hc405047;
      6803: inst = 32'h8220000;
      6804: inst = 32'h10408000;
      6805: inst = 32'hc405048;
      6806: inst = 32'h8220000;
      6807: inst = 32'h10408000;
      6808: inst = 32'hc405049;
      6809: inst = 32'h8220000;
      6810: inst = 32'h10408000;
      6811: inst = 32'hc40504a;
      6812: inst = 32'h8220000;
      6813: inst = 32'h10408000;
      6814: inst = 32'hc40504b;
      6815: inst = 32'h8220000;
      6816: inst = 32'h10408000;
      6817: inst = 32'hc40504c;
      6818: inst = 32'h8220000;
      6819: inst = 32'h10408000;
      6820: inst = 32'hc40504d;
      6821: inst = 32'h8220000;
      6822: inst = 32'h10408000;
      6823: inst = 32'hc40504e;
      6824: inst = 32'h8220000;
      6825: inst = 32'h10408000;
      6826: inst = 32'hc405077;
      6827: inst = 32'h8220000;
      6828: inst = 32'h10408000;
      6829: inst = 32'hc405078;
      6830: inst = 32'h8220000;
      6831: inst = 32'h10408000;
      6832: inst = 32'hc405079;
      6833: inst = 32'h8220000;
      6834: inst = 32'h10408000;
      6835: inst = 32'hc40507a;
      6836: inst = 32'h8220000;
      6837: inst = 32'h10408000;
      6838: inst = 32'hc40507b;
      6839: inst = 32'h8220000;
      6840: inst = 32'h10408000;
      6841: inst = 32'hc40507c;
      6842: inst = 32'h8220000;
      6843: inst = 32'h10408000;
      6844: inst = 32'hc40507d;
      6845: inst = 32'h8220000;
      6846: inst = 32'h10408000;
      6847: inst = 32'hc40507e;
      6848: inst = 32'h8220000;
      6849: inst = 32'h10408000;
      6850: inst = 32'hc405088;
      6851: inst = 32'h8220000;
      6852: inst = 32'h10408000;
      6853: inst = 32'hc405089;
      6854: inst = 32'h8220000;
      6855: inst = 32'h10408000;
      6856: inst = 32'hc40508a;
      6857: inst = 32'h8220000;
      6858: inst = 32'h10408000;
      6859: inst = 32'hc40508b;
      6860: inst = 32'h8220000;
      6861: inst = 32'h10408000;
      6862: inst = 32'hc40508c;
      6863: inst = 32'h8220000;
      6864: inst = 32'h10408000;
      6865: inst = 32'hc40508d;
      6866: inst = 32'h8220000;
      6867: inst = 32'h10408000;
      6868: inst = 32'hc40508e;
      6869: inst = 32'h8220000;
      6870: inst = 32'h10408000;
      6871: inst = 32'hc40508f;
      6872: inst = 32'h8220000;
      6873: inst = 32'h10408000;
      6874: inst = 32'hc405090;
      6875: inst = 32'h8220000;
      6876: inst = 32'h10408000;
      6877: inst = 32'hc405091;
      6878: inst = 32'h8220000;
      6879: inst = 32'h10408000;
      6880: inst = 32'hc405092;
      6881: inst = 32'h8220000;
      6882: inst = 32'h10408000;
      6883: inst = 32'hc405093;
      6884: inst = 32'h8220000;
      6885: inst = 32'h10408000;
      6886: inst = 32'hc405094;
      6887: inst = 32'h8220000;
      6888: inst = 32'h10408000;
      6889: inst = 32'hc405095;
      6890: inst = 32'h8220000;
      6891: inst = 32'h10408000;
      6892: inst = 32'hc405096;
      6893: inst = 32'h8220000;
      6894: inst = 32'h10408000;
      6895: inst = 32'hc405097;
      6896: inst = 32'h8220000;
      6897: inst = 32'h10408000;
      6898: inst = 32'hc4050a1;
      6899: inst = 32'h8220000;
      6900: inst = 32'h10408000;
      6901: inst = 32'hc4050a2;
      6902: inst = 32'h8220000;
      6903: inst = 32'h10408000;
      6904: inst = 32'hc4050a3;
      6905: inst = 32'h8220000;
      6906: inst = 32'h10408000;
      6907: inst = 32'hc4050a4;
      6908: inst = 32'h8220000;
      6909: inst = 32'h10408000;
      6910: inst = 32'hc4050a5;
      6911: inst = 32'h8220000;
      6912: inst = 32'h10408000;
      6913: inst = 32'hc4050a6;
      6914: inst = 32'h8220000;
      6915: inst = 32'h10408000;
      6916: inst = 32'hc4050a7;
      6917: inst = 32'h8220000;
      6918: inst = 32'h10408000;
      6919: inst = 32'hc4050a8;
      6920: inst = 32'h8220000;
      6921: inst = 32'h10408000;
      6922: inst = 32'hc4050a9;
      6923: inst = 32'h8220000;
      6924: inst = 32'h10408000;
      6925: inst = 32'hc4050aa;
      6926: inst = 32'h8220000;
      6927: inst = 32'h10408000;
      6928: inst = 32'hc4050ab;
      6929: inst = 32'h8220000;
      6930: inst = 32'h10408000;
      6931: inst = 32'hc4050ac;
      6932: inst = 32'h8220000;
      6933: inst = 32'h10408000;
      6934: inst = 32'hc4050ad;
      6935: inst = 32'h8220000;
      6936: inst = 32'h10408000;
      6937: inst = 32'hc4050ae;
      6938: inst = 32'h8220000;
      6939: inst = 32'h10408000;
      6940: inst = 32'hc4050d7;
      6941: inst = 32'h8220000;
      6942: inst = 32'h10408000;
      6943: inst = 32'hc4050d8;
      6944: inst = 32'h8220000;
      6945: inst = 32'h10408000;
      6946: inst = 32'hc4050d9;
      6947: inst = 32'h8220000;
      6948: inst = 32'h10408000;
      6949: inst = 32'hc4050da;
      6950: inst = 32'h8220000;
      6951: inst = 32'h10408000;
      6952: inst = 32'hc4050db;
      6953: inst = 32'h8220000;
      6954: inst = 32'h10408000;
      6955: inst = 32'hc4050dc;
      6956: inst = 32'h8220000;
      6957: inst = 32'h10408000;
      6958: inst = 32'hc4050dd;
      6959: inst = 32'h8220000;
      6960: inst = 32'h10408000;
      6961: inst = 32'hc4050de;
      6962: inst = 32'h8220000;
      6963: inst = 32'h10408000;
      6964: inst = 32'hc4050e8;
      6965: inst = 32'h8220000;
      6966: inst = 32'h10408000;
      6967: inst = 32'hc4050e9;
      6968: inst = 32'h8220000;
      6969: inst = 32'h10408000;
      6970: inst = 32'hc4050ea;
      6971: inst = 32'h8220000;
      6972: inst = 32'h10408000;
      6973: inst = 32'hc4050eb;
      6974: inst = 32'h8220000;
      6975: inst = 32'h10408000;
      6976: inst = 32'hc4050ec;
      6977: inst = 32'h8220000;
      6978: inst = 32'h10408000;
      6979: inst = 32'hc4050ed;
      6980: inst = 32'h8220000;
      6981: inst = 32'h10408000;
      6982: inst = 32'hc4050ee;
      6983: inst = 32'h8220000;
      6984: inst = 32'h10408000;
      6985: inst = 32'hc4050ef;
      6986: inst = 32'h8220000;
      6987: inst = 32'h10408000;
      6988: inst = 32'hc4050f0;
      6989: inst = 32'h8220000;
      6990: inst = 32'h10408000;
      6991: inst = 32'hc4050f1;
      6992: inst = 32'h8220000;
      6993: inst = 32'h10408000;
      6994: inst = 32'hc4050f2;
      6995: inst = 32'h8220000;
      6996: inst = 32'h10408000;
      6997: inst = 32'hc4050f3;
      6998: inst = 32'h8220000;
      6999: inst = 32'h10408000;
      7000: inst = 32'hc4050f4;
      7001: inst = 32'h8220000;
      7002: inst = 32'h10408000;
      7003: inst = 32'hc4050f5;
      7004: inst = 32'h8220000;
      7005: inst = 32'h10408000;
      7006: inst = 32'hc4050f6;
      7007: inst = 32'h8220000;
      7008: inst = 32'h10408000;
      7009: inst = 32'hc4050f7;
      7010: inst = 32'h8220000;
      7011: inst = 32'h10408000;
      7012: inst = 32'hc405101;
      7013: inst = 32'h8220000;
      7014: inst = 32'h10408000;
      7015: inst = 32'hc405102;
      7016: inst = 32'h8220000;
      7017: inst = 32'h10408000;
      7018: inst = 32'hc405103;
      7019: inst = 32'h8220000;
      7020: inst = 32'h10408000;
      7021: inst = 32'hc405104;
      7022: inst = 32'h8220000;
      7023: inst = 32'h10408000;
      7024: inst = 32'hc405105;
      7025: inst = 32'h8220000;
      7026: inst = 32'h10408000;
      7027: inst = 32'hc405106;
      7028: inst = 32'h8220000;
      7029: inst = 32'h10408000;
      7030: inst = 32'hc405107;
      7031: inst = 32'h8220000;
      7032: inst = 32'h10408000;
      7033: inst = 32'hc405108;
      7034: inst = 32'h8220000;
      7035: inst = 32'h10408000;
      7036: inst = 32'hc405109;
      7037: inst = 32'h8220000;
      7038: inst = 32'h10408000;
      7039: inst = 32'hc40510a;
      7040: inst = 32'h8220000;
      7041: inst = 32'h10408000;
      7042: inst = 32'hc40510b;
      7043: inst = 32'h8220000;
      7044: inst = 32'h10408000;
      7045: inst = 32'hc40510c;
      7046: inst = 32'h8220000;
      7047: inst = 32'h10408000;
      7048: inst = 32'hc40510d;
      7049: inst = 32'h8220000;
      7050: inst = 32'h10408000;
      7051: inst = 32'hc40510e;
      7052: inst = 32'h8220000;
      7053: inst = 32'h10408000;
      7054: inst = 32'hc405137;
      7055: inst = 32'h8220000;
      7056: inst = 32'h10408000;
      7057: inst = 32'hc405138;
      7058: inst = 32'h8220000;
      7059: inst = 32'h10408000;
      7060: inst = 32'hc405139;
      7061: inst = 32'h8220000;
      7062: inst = 32'h10408000;
      7063: inst = 32'hc40513a;
      7064: inst = 32'h8220000;
      7065: inst = 32'h10408000;
      7066: inst = 32'hc40513b;
      7067: inst = 32'h8220000;
      7068: inst = 32'h10408000;
      7069: inst = 32'hc40513c;
      7070: inst = 32'h8220000;
      7071: inst = 32'h10408000;
      7072: inst = 32'hc40513d;
      7073: inst = 32'h8220000;
      7074: inst = 32'h10408000;
      7075: inst = 32'hc40513e;
      7076: inst = 32'h8220000;
      7077: inst = 32'h10408000;
      7078: inst = 32'hc405148;
      7079: inst = 32'h8220000;
      7080: inst = 32'h10408000;
      7081: inst = 32'hc405149;
      7082: inst = 32'h8220000;
      7083: inst = 32'h10408000;
      7084: inst = 32'hc40514a;
      7085: inst = 32'h8220000;
      7086: inst = 32'h10408000;
      7087: inst = 32'hc40514b;
      7088: inst = 32'h8220000;
      7089: inst = 32'h10408000;
      7090: inst = 32'hc40514c;
      7091: inst = 32'h8220000;
      7092: inst = 32'h10408000;
      7093: inst = 32'hc40514d;
      7094: inst = 32'h8220000;
      7095: inst = 32'h10408000;
      7096: inst = 32'hc40514e;
      7097: inst = 32'h8220000;
      7098: inst = 32'h10408000;
      7099: inst = 32'hc40514f;
      7100: inst = 32'h8220000;
      7101: inst = 32'h10408000;
      7102: inst = 32'hc405150;
      7103: inst = 32'h8220000;
      7104: inst = 32'h10408000;
      7105: inst = 32'hc405151;
      7106: inst = 32'h8220000;
      7107: inst = 32'h10408000;
      7108: inst = 32'hc405152;
      7109: inst = 32'h8220000;
      7110: inst = 32'h10408000;
      7111: inst = 32'hc405153;
      7112: inst = 32'h8220000;
      7113: inst = 32'h10408000;
      7114: inst = 32'hc405154;
      7115: inst = 32'h8220000;
      7116: inst = 32'h10408000;
      7117: inst = 32'hc405155;
      7118: inst = 32'h8220000;
      7119: inst = 32'h10408000;
      7120: inst = 32'hc405156;
      7121: inst = 32'h8220000;
      7122: inst = 32'h10408000;
      7123: inst = 32'hc405157;
      7124: inst = 32'h8220000;
      7125: inst = 32'h10408000;
      7126: inst = 32'hc405161;
      7127: inst = 32'h8220000;
      7128: inst = 32'h10408000;
      7129: inst = 32'hc405162;
      7130: inst = 32'h8220000;
      7131: inst = 32'h10408000;
      7132: inst = 32'hc405163;
      7133: inst = 32'h8220000;
      7134: inst = 32'h10408000;
      7135: inst = 32'hc405164;
      7136: inst = 32'h8220000;
      7137: inst = 32'h10408000;
      7138: inst = 32'hc405165;
      7139: inst = 32'h8220000;
      7140: inst = 32'h10408000;
      7141: inst = 32'hc405166;
      7142: inst = 32'h8220000;
      7143: inst = 32'h10408000;
      7144: inst = 32'hc405167;
      7145: inst = 32'h8220000;
      7146: inst = 32'h10408000;
      7147: inst = 32'hc405168;
      7148: inst = 32'h8220000;
      7149: inst = 32'h10408000;
      7150: inst = 32'hc405169;
      7151: inst = 32'h8220000;
      7152: inst = 32'h10408000;
      7153: inst = 32'hc40516a;
      7154: inst = 32'h8220000;
      7155: inst = 32'h10408000;
      7156: inst = 32'hc40516b;
      7157: inst = 32'h8220000;
      7158: inst = 32'h10408000;
      7159: inst = 32'hc40516c;
      7160: inst = 32'h8220000;
      7161: inst = 32'h10408000;
      7162: inst = 32'hc40516d;
      7163: inst = 32'h8220000;
      7164: inst = 32'h10408000;
      7165: inst = 32'hc40516e;
      7166: inst = 32'h8220000;
      7167: inst = 32'h10408000;
      7168: inst = 32'hc405197;
      7169: inst = 32'h8220000;
      7170: inst = 32'h10408000;
      7171: inst = 32'hc405198;
      7172: inst = 32'h8220000;
      7173: inst = 32'h10408000;
      7174: inst = 32'hc405199;
      7175: inst = 32'h8220000;
      7176: inst = 32'h10408000;
      7177: inst = 32'hc40519a;
      7178: inst = 32'h8220000;
      7179: inst = 32'h10408000;
      7180: inst = 32'hc40519b;
      7181: inst = 32'h8220000;
      7182: inst = 32'h10408000;
      7183: inst = 32'hc40519c;
      7184: inst = 32'h8220000;
      7185: inst = 32'h10408000;
      7186: inst = 32'hc40519d;
      7187: inst = 32'h8220000;
      7188: inst = 32'h10408000;
      7189: inst = 32'hc4051aa;
      7190: inst = 32'h8220000;
      7191: inst = 32'h10408000;
      7192: inst = 32'hc4051ab;
      7193: inst = 32'h8220000;
      7194: inst = 32'h10408000;
      7195: inst = 32'hc4051ac;
      7196: inst = 32'h8220000;
      7197: inst = 32'h10408000;
      7198: inst = 32'hc4051ad;
      7199: inst = 32'h8220000;
      7200: inst = 32'h10408000;
      7201: inst = 32'hc4051ae;
      7202: inst = 32'h8220000;
      7203: inst = 32'h10408000;
      7204: inst = 32'hc4051af;
      7205: inst = 32'h8220000;
      7206: inst = 32'h10408000;
      7207: inst = 32'hc4051b0;
      7208: inst = 32'h8220000;
      7209: inst = 32'h10408000;
      7210: inst = 32'hc4051b1;
      7211: inst = 32'h8220000;
      7212: inst = 32'h10408000;
      7213: inst = 32'hc4051b2;
      7214: inst = 32'h8220000;
      7215: inst = 32'h10408000;
      7216: inst = 32'hc4051b3;
      7217: inst = 32'h8220000;
      7218: inst = 32'h10408000;
      7219: inst = 32'hc4051b4;
      7220: inst = 32'h8220000;
      7221: inst = 32'h10408000;
      7222: inst = 32'hc4051b5;
      7223: inst = 32'h8220000;
      7224: inst = 32'h10408000;
      7225: inst = 32'hc4051c2;
      7226: inst = 32'h8220000;
      7227: inst = 32'h10408000;
      7228: inst = 32'hc4051c3;
      7229: inst = 32'h8220000;
      7230: inst = 32'h10408000;
      7231: inst = 32'hc4051c4;
      7232: inst = 32'h8220000;
      7233: inst = 32'h10408000;
      7234: inst = 32'hc4051c5;
      7235: inst = 32'h8220000;
      7236: inst = 32'h10408000;
      7237: inst = 32'hc4051c6;
      7238: inst = 32'h8220000;
      7239: inst = 32'h10408000;
      7240: inst = 32'hc4051c7;
      7241: inst = 32'h8220000;
      7242: inst = 32'h10408000;
      7243: inst = 32'hc4051c8;
      7244: inst = 32'h8220000;
      7245: inst = 32'h10408000;
      7246: inst = 32'hc4051c9;
      7247: inst = 32'h8220000;
      7248: inst = 32'h10408000;
      7249: inst = 32'hc4051ca;
      7250: inst = 32'h8220000;
      7251: inst = 32'h10408000;
      7252: inst = 32'hc4051cb;
      7253: inst = 32'h8220000;
      7254: inst = 32'h10408000;
      7255: inst = 32'hc4051cc;
      7256: inst = 32'h8220000;
      7257: inst = 32'h10408000;
      7258: inst = 32'hc4051cd;
      7259: inst = 32'h8220000;
      7260: inst = 32'h10408000;
      7261: inst = 32'hc4051ce;
      7262: inst = 32'h8220000;
      7263: inst = 32'h10408000;
      7264: inst = 32'hc4051f7;
      7265: inst = 32'h8220000;
      7266: inst = 32'h10408000;
      7267: inst = 32'hc4051f8;
      7268: inst = 32'h8220000;
      7269: inst = 32'h10408000;
      7270: inst = 32'hc4051f9;
      7271: inst = 32'h8220000;
      7272: inst = 32'h10408000;
      7273: inst = 32'hc4051fa;
      7274: inst = 32'h8220000;
      7275: inst = 32'h10408000;
      7276: inst = 32'hc4051fb;
      7277: inst = 32'h8220000;
      7278: inst = 32'h10408000;
      7279: inst = 32'hc4051fc;
      7280: inst = 32'h8220000;
      7281: inst = 32'h10408000;
      7282: inst = 32'hc40520a;
      7283: inst = 32'h8220000;
      7284: inst = 32'h10408000;
      7285: inst = 32'hc40520b;
      7286: inst = 32'h8220000;
      7287: inst = 32'h10408000;
      7288: inst = 32'hc40520c;
      7289: inst = 32'h8220000;
      7290: inst = 32'h10408000;
      7291: inst = 32'hc40520d;
      7292: inst = 32'h8220000;
      7293: inst = 32'h10408000;
      7294: inst = 32'hc40520e;
      7295: inst = 32'h8220000;
      7296: inst = 32'h10408000;
      7297: inst = 32'hc40520f;
      7298: inst = 32'h8220000;
      7299: inst = 32'h10408000;
      7300: inst = 32'hc405210;
      7301: inst = 32'h8220000;
      7302: inst = 32'h10408000;
      7303: inst = 32'hc405211;
      7304: inst = 32'h8220000;
      7305: inst = 32'h10408000;
      7306: inst = 32'hc405212;
      7307: inst = 32'h8220000;
      7308: inst = 32'h10408000;
      7309: inst = 32'hc405213;
      7310: inst = 32'h8220000;
      7311: inst = 32'h10408000;
      7312: inst = 32'hc405214;
      7313: inst = 32'h8220000;
      7314: inst = 32'h10408000;
      7315: inst = 32'hc405215;
      7316: inst = 32'h8220000;
      7317: inst = 32'h10408000;
      7318: inst = 32'hc405223;
      7319: inst = 32'h8220000;
      7320: inst = 32'h10408000;
      7321: inst = 32'hc405224;
      7322: inst = 32'h8220000;
      7323: inst = 32'h10408000;
      7324: inst = 32'hc405225;
      7325: inst = 32'h8220000;
      7326: inst = 32'h10408000;
      7327: inst = 32'hc405226;
      7328: inst = 32'h8220000;
      7329: inst = 32'h10408000;
      7330: inst = 32'hc405227;
      7331: inst = 32'h8220000;
      7332: inst = 32'h10408000;
      7333: inst = 32'hc405228;
      7334: inst = 32'h8220000;
      7335: inst = 32'h10408000;
      7336: inst = 32'hc405229;
      7337: inst = 32'h8220000;
      7338: inst = 32'h10408000;
      7339: inst = 32'hc40522a;
      7340: inst = 32'h8220000;
      7341: inst = 32'h10408000;
      7342: inst = 32'hc40522b;
      7343: inst = 32'h8220000;
      7344: inst = 32'h10408000;
      7345: inst = 32'hc40522c;
      7346: inst = 32'h8220000;
      7347: inst = 32'h10408000;
      7348: inst = 32'hc40522d;
      7349: inst = 32'h8220000;
      7350: inst = 32'h10408000;
      7351: inst = 32'hc40522e;
      7352: inst = 32'h8220000;
      7353: inst = 32'h10408000;
      7354: inst = 32'hc405257;
      7355: inst = 32'h8220000;
      7356: inst = 32'h10408000;
      7357: inst = 32'hc405258;
      7358: inst = 32'h8220000;
      7359: inst = 32'h10408000;
      7360: inst = 32'hc405259;
      7361: inst = 32'h8220000;
      7362: inst = 32'h10408000;
      7363: inst = 32'hc40525a;
      7364: inst = 32'h8220000;
      7365: inst = 32'h10408000;
      7366: inst = 32'hc40525b;
      7367: inst = 32'h8220000;
      7368: inst = 32'h10408000;
      7369: inst = 32'hc40526a;
      7370: inst = 32'h8220000;
      7371: inst = 32'h10408000;
      7372: inst = 32'hc40526b;
      7373: inst = 32'h8220000;
      7374: inst = 32'h10408000;
      7375: inst = 32'hc40526c;
      7376: inst = 32'h8220000;
      7377: inst = 32'h10408000;
      7378: inst = 32'hc40526d;
      7379: inst = 32'h8220000;
      7380: inst = 32'h10408000;
      7381: inst = 32'hc40526e;
      7382: inst = 32'h8220000;
      7383: inst = 32'h10408000;
      7384: inst = 32'hc40526f;
      7385: inst = 32'h8220000;
      7386: inst = 32'h10408000;
      7387: inst = 32'hc405270;
      7388: inst = 32'h8220000;
      7389: inst = 32'h10408000;
      7390: inst = 32'hc405271;
      7391: inst = 32'h8220000;
      7392: inst = 32'h10408000;
      7393: inst = 32'hc405272;
      7394: inst = 32'h8220000;
      7395: inst = 32'h10408000;
      7396: inst = 32'hc405273;
      7397: inst = 32'h8220000;
      7398: inst = 32'h10408000;
      7399: inst = 32'hc405274;
      7400: inst = 32'h8220000;
      7401: inst = 32'h10408000;
      7402: inst = 32'hc405275;
      7403: inst = 32'h8220000;
      7404: inst = 32'h10408000;
      7405: inst = 32'hc405284;
      7406: inst = 32'h8220000;
      7407: inst = 32'h10408000;
      7408: inst = 32'hc405285;
      7409: inst = 32'h8220000;
      7410: inst = 32'h10408000;
      7411: inst = 32'hc405286;
      7412: inst = 32'h8220000;
      7413: inst = 32'h10408000;
      7414: inst = 32'hc405287;
      7415: inst = 32'h8220000;
      7416: inst = 32'h10408000;
      7417: inst = 32'hc405288;
      7418: inst = 32'h8220000;
      7419: inst = 32'h10408000;
      7420: inst = 32'hc405289;
      7421: inst = 32'h8220000;
      7422: inst = 32'h10408000;
      7423: inst = 32'hc40528a;
      7424: inst = 32'h8220000;
      7425: inst = 32'h10408000;
      7426: inst = 32'hc40528b;
      7427: inst = 32'h8220000;
      7428: inst = 32'h10408000;
      7429: inst = 32'hc40528c;
      7430: inst = 32'h8220000;
      7431: inst = 32'h10408000;
      7432: inst = 32'hc40528d;
      7433: inst = 32'h8220000;
      7434: inst = 32'h10408000;
      7435: inst = 32'hc40528e;
      7436: inst = 32'h8220000;
      7437: inst = 32'h10408000;
      7438: inst = 32'hc4052b7;
      7439: inst = 32'h8220000;
      7440: inst = 32'h10408000;
      7441: inst = 32'hc4052b8;
      7442: inst = 32'h8220000;
      7443: inst = 32'h10408000;
      7444: inst = 32'hc4052b9;
      7445: inst = 32'h8220000;
      7446: inst = 32'h10408000;
      7447: inst = 32'hc4052ba;
      7448: inst = 32'h8220000;
      7449: inst = 32'h10408000;
      7450: inst = 32'hc4052bb;
      7451: inst = 32'h8220000;
      7452: inst = 32'h10408000;
      7453: inst = 32'hc4052ca;
      7454: inst = 32'h8220000;
      7455: inst = 32'h10408000;
      7456: inst = 32'hc4052cb;
      7457: inst = 32'h8220000;
      7458: inst = 32'h10408000;
      7459: inst = 32'hc4052cc;
      7460: inst = 32'h8220000;
      7461: inst = 32'h10408000;
      7462: inst = 32'hc4052cd;
      7463: inst = 32'h8220000;
      7464: inst = 32'h10408000;
      7465: inst = 32'hc4052ce;
      7466: inst = 32'h8220000;
      7467: inst = 32'h10408000;
      7468: inst = 32'hc4052cf;
      7469: inst = 32'h8220000;
      7470: inst = 32'h10408000;
      7471: inst = 32'hc4052d0;
      7472: inst = 32'h8220000;
      7473: inst = 32'h10408000;
      7474: inst = 32'hc4052d1;
      7475: inst = 32'h8220000;
      7476: inst = 32'h10408000;
      7477: inst = 32'hc4052d2;
      7478: inst = 32'h8220000;
      7479: inst = 32'h10408000;
      7480: inst = 32'hc4052d3;
      7481: inst = 32'h8220000;
      7482: inst = 32'h10408000;
      7483: inst = 32'hc4052d4;
      7484: inst = 32'h8220000;
      7485: inst = 32'h10408000;
      7486: inst = 32'hc4052d5;
      7487: inst = 32'h8220000;
      7488: inst = 32'h10408000;
      7489: inst = 32'hc4052e4;
      7490: inst = 32'h8220000;
      7491: inst = 32'h10408000;
      7492: inst = 32'hc4052e5;
      7493: inst = 32'h8220000;
      7494: inst = 32'h10408000;
      7495: inst = 32'hc4052e6;
      7496: inst = 32'h8220000;
      7497: inst = 32'h10408000;
      7498: inst = 32'hc4052e7;
      7499: inst = 32'h8220000;
      7500: inst = 32'h10408000;
      7501: inst = 32'hc4052e8;
      7502: inst = 32'h8220000;
      7503: inst = 32'h10408000;
      7504: inst = 32'hc4052e9;
      7505: inst = 32'h8220000;
      7506: inst = 32'h10408000;
      7507: inst = 32'hc4052ea;
      7508: inst = 32'h8220000;
      7509: inst = 32'h10408000;
      7510: inst = 32'hc4052eb;
      7511: inst = 32'h8220000;
      7512: inst = 32'h10408000;
      7513: inst = 32'hc4052ec;
      7514: inst = 32'h8220000;
      7515: inst = 32'h10408000;
      7516: inst = 32'hc4052ed;
      7517: inst = 32'h8220000;
      7518: inst = 32'h10408000;
      7519: inst = 32'hc4052ee;
      7520: inst = 32'h8220000;
      7521: inst = 32'hc2094b2;
      7522: inst = 32'h10408000;
      7523: inst = 32'hc403feb;
      7524: inst = 32'h8220000;
      7525: inst = 32'h10408000;
      7526: inst = 32'hc40404b;
      7527: inst = 32'h8220000;
      7528: inst = 32'h10408000;
      7529: inst = 32'hc4040ab;
      7530: inst = 32'h8220000;
      7531: inst = 32'h10408000;
      7532: inst = 32'hc40410b;
      7533: inst = 32'h8220000;
      7534: inst = 32'h10408000;
      7535: inst = 32'hc40416b;
      7536: inst = 32'h8220000;
      7537: inst = 32'h10408000;
      7538: inst = 32'hc4041cb;
      7539: inst = 32'h8220000;
      7540: inst = 32'h10408000;
      7541: inst = 32'hc40422b;
      7542: inst = 32'h8220000;
      7543: inst = 32'h10408000;
      7544: inst = 32'hc40428b;
      7545: inst = 32'h8220000;
      7546: inst = 32'hc20b596;
      7547: inst = 32'h10408000;
      7548: inst = 32'hc4041da;
      7549: inst = 32'h8220000;
      7550: inst = 32'h10408000;
      7551: inst = 32'hc4041db;
      7552: inst = 32'h8220000;
      7553: inst = 32'h10408000;
      7554: inst = 32'hc4041dc;
      7555: inst = 32'h8220000;
      7556: inst = 32'h10408000;
      7557: inst = 32'hc4041dd;
      7558: inst = 32'h8220000;
      7559: inst = 32'h10408000;
      7560: inst = 32'hc4041de;
      7561: inst = 32'h8220000;
      7562: inst = 32'h10408000;
      7563: inst = 32'hc4041df;
      7564: inst = 32'h8220000;
      7565: inst = 32'h10408000;
      7566: inst = 32'hc4041e0;
      7567: inst = 32'h8220000;
      7568: inst = 32'h10408000;
      7569: inst = 32'hc4041e1;
      7570: inst = 32'h8220000;
      7571: inst = 32'h10408000;
      7572: inst = 32'hc4041e2;
      7573: inst = 32'h8220000;
      7574: inst = 32'h10408000;
      7575: inst = 32'hc4041e3;
      7576: inst = 32'h8220000;
      7577: inst = 32'h10408000;
      7578: inst = 32'hc4041e4;
      7579: inst = 32'h8220000;
      7580: inst = 32'h10408000;
      7581: inst = 32'hc4041e5;
      7582: inst = 32'h8220000;
      7583: inst = 32'h10408000;
      7584: inst = 32'hc4041e6;
      7585: inst = 32'h8220000;
      7586: inst = 32'h10408000;
      7587: inst = 32'hc4041e7;
      7588: inst = 32'h8220000;
      7589: inst = 32'h10408000;
      7590: inst = 32'hc4041e8;
      7591: inst = 32'h8220000;
      7592: inst = 32'h10408000;
      7593: inst = 32'hc4041e9;
      7594: inst = 32'h8220000;
      7595: inst = 32'h10408000;
      7596: inst = 32'hc4041ea;
      7597: inst = 32'h8220000;
      7598: inst = 32'h10408000;
      7599: inst = 32'hc4041eb;
      7600: inst = 32'h8220000;
      7601: inst = 32'h10408000;
      7602: inst = 32'hc4041ec;
      7603: inst = 32'h8220000;
      7604: inst = 32'h10408000;
      7605: inst = 32'hc4041ed;
      7606: inst = 32'h8220000;
      7607: inst = 32'h10408000;
      7608: inst = 32'hc4041ee;
      7609: inst = 32'h8220000;
      7610: inst = 32'h10408000;
      7611: inst = 32'hc4041ef;
      7612: inst = 32'h8220000;
      7613: inst = 32'h10408000;
      7614: inst = 32'hc4041f0;
      7615: inst = 32'h8220000;
      7616: inst = 32'h10408000;
      7617: inst = 32'hc4041f1;
      7618: inst = 32'h8220000;
      7619: inst = 32'h10408000;
      7620: inst = 32'hc4041f2;
      7621: inst = 32'h8220000;
      7622: inst = 32'h10408000;
      7623: inst = 32'hc4041f3;
      7624: inst = 32'h8220000;
      7625: inst = 32'h10408000;
      7626: inst = 32'hc4041f4;
      7627: inst = 32'h8220000;
      7628: inst = 32'h10408000;
      7629: inst = 32'hc4041f5;
      7630: inst = 32'h8220000;
      7631: inst = 32'h10408000;
      7632: inst = 32'hc4041f6;
      7633: inst = 32'h8220000;
      7634: inst = 32'h10408000;
      7635: inst = 32'hc4041f7;
      7636: inst = 32'h8220000;
      7637: inst = 32'h10408000;
      7638: inst = 32'hc4041f8;
      7639: inst = 32'h8220000;
      7640: inst = 32'h10408000;
      7641: inst = 32'hc4041f9;
      7642: inst = 32'h8220000;
      7643: inst = 32'h10408000;
      7644: inst = 32'hc4041fa;
      7645: inst = 32'h8220000;
      7646: inst = 32'h10408000;
      7647: inst = 32'hc4041fb;
      7648: inst = 32'h8220000;
      7649: inst = 32'h10408000;
      7650: inst = 32'hc4041fc;
      7651: inst = 32'h8220000;
      7652: inst = 32'h10408000;
      7653: inst = 32'hc4041fd;
      7654: inst = 32'h8220000;
      7655: inst = 32'h10408000;
      7656: inst = 32'hc4041fe;
      7657: inst = 32'h8220000;
      7658: inst = 32'h10408000;
      7659: inst = 32'hc4041ff;
      7660: inst = 32'h8220000;
      7661: inst = 32'h10408000;
      7662: inst = 32'hc404200;
      7663: inst = 32'h8220000;
      7664: inst = 32'h10408000;
      7665: inst = 32'hc404201;
      7666: inst = 32'h8220000;
      7667: inst = 32'h10408000;
      7668: inst = 32'hc404202;
      7669: inst = 32'h8220000;
      7670: inst = 32'h10408000;
      7671: inst = 32'hc404203;
      7672: inst = 32'h8220000;
      7673: inst = 32'h10408000;
      7674: inst = 32'hc404204;
      7675: inst = 32'h8220000;
      7676: inst = 32'h10408000;
      7677: inst = 32'hc404205;
      7678: inst = 32'h8220000;
      7679: inst = 32'h10408000;
      7680: inst = 32'hc404bfa;
      7681: inst = 32'h8220000;
      7682: inst = 32'h10408000;
      7683: inst = 32'hc404bfb;
      7684: inst = 32'h8220000;
      7685: inst = 32'h10408000;
      7686: inst = 32'hc404bfc;
      7687: inst = 32'h8220000;
      7688: inst = 32'h10408000;
      7689: inst = 32'hc404bfd;
      7690: inst = 32'h8220000;
      7691: inst = 32'h10408000;
      7692: inst = 32'hc404bfe;
      7693: inst = 32'h8220000;
      7694: inst = 32'h10408000;
      7695: inst = 32'hc404bff;
      7696: inst = 32'h8220000;
      7697: inst = 32'h10408000;
      7698: inst = 32'hc404c00;
      7699: inst = 32'h8220000;
      7700: inst = 32'h10408000;
      7701: inst = 32'hc404c01;
      7702: inst = 32'h8220000;
      7703: inst = 32'h10408000;
      7704: inst = 32'hc404c02;
      7705: inst = 32'h8220000;
      7706: inst = 32'h10408000;
      7707: inst = 32'hc404c03;
      7708: inst = 32'h8220000;
      7709: inst = 32'h10408000;
      7710: inst = 32'hc404c04;
      7711: inst = 32'h8220000;
      7712: inst = 32'h10408000;
      7713: inst = 32'hc404c05;
      7714: inst = 32'h8220000;
      7715: inst = 32'h10408000;
      7716: inst = 32'hc404c06;
      7717: inst = 32'h8220000;
      7718: inst = 32'h10408000;
      7719: inst = 32'hc404c07;
      7720: inst = 32'h8220000;
      7721: inst = 32'h10408000;
      7722: inst = 32'hc404c08;
      7723: inst = 32'h8220000;
      7724: inst = 32'h10408000;
      7725: inst = 32'hc404c09;
      7726: inst = 32'h8220000;
      7727: inst = 32'h10408000;
      7728: inst = 32'hc404c0a;
      7729: inst = 32'h8220000;
      7730: inst = 32'h10408000;
      7731: inst = 32'hc404c0b;
      7732: inst = 32'h8220000;
      7733: inst = 32'h10408000;
      7734: inst = 32'hc404c0c;
      7735: inst = 32'h8220000;
      7736: inst = 32'h10408000;
      7737: inst = 32'hc404c0d;
      7738: inst = 32'h8220000;
      7739: inst = 32'h10408000;
      7740: inst = 32'hc404c0e;
      7741: inst = 32'h8220000;
      7742: inst = 32'h10408000;
      7743: inst = 32'hc404c0f;
      7744: inst = 32'h8220000;
      7745: inst = 32'h10408000;
      7746: inst = 32'hc404c10;
      7747: inst = 32'h8220000;
      7748: inst = 32'h10408000;
      7749: inst = 32'hc404c11;
      7750: inst = 32'h8220000;
      7751: inst = 32'h10408000;
      7752: inst = 32'hc404c12;
      7753: inst = 32'h8220000;
      7754: inst = 32'h10408000;
      7755: inst = 32'hc404c13;
      7756: inst = 32'h8220000;
      7757: inst = 32'h10408000;
      7758: inst = 32'hc404c14;
      7759: inst = 32'h8220000;
      7760: inst = 32'h10408000;
      7761: inst = 32'hc404c15;
      7762: inst = 32'h8220000;
      7763: inst = 32'h10408000;
      7764: inst = 32'hc404c16;
      7765: inst = 32'h8220000;
      7766: inst = 32'h10408000;
      7767: inst = 32'hc404c17;
      7768: inst = 32'h8220000;
      7769: inst = 32'h10408000;
      7770: inst = 32'hc404c18;
      7771: inst = 32'h8220000;
      7772: inst = 32'h10408000;
      7773: inst = 32'hc404c19;
      7774: inst = 32'h8220000;
      7775: inst = 32'h10408000;
      7776: inst = 32'hc404c1a;
      7777: inst = 32'h8220000;
      7778: inst = 32'h10408000;
      7779: inst = 32'hc404c1b;
      7780: inst = 32'h8220000;
      7781: inst = 32'h10408000;
      7782: inst = 32'hc404c1c;
      7783: inst = 32'h8220000;
      7784: inst = 32'h10408000;
      7785: inst = 32'hc404c1d;
      7786: inst = 32'h8220000;
      7787: inst = 32'h10408000;
      7788: inst = 32'hc404c1e;
      7789: inst = 32'h8220000;
      7790: inst = 32'h10408000;
      7791: inst = 32'hc404c1f;
      7792: inst = 32'h8220000;
      7793: inst = 32'h10408000;
      7794: inst = 32'hc404c20;
      7795: inst = 32'h8220000;
      7796: inst = 32'h10408000;
      7797: inst = 32'hc404c21;
      7798: inst = 32'h8220000;
      7799: inst = 32'h10408000;
      7800: inst = 32'hc404c22;
      7801: inst = 32'h8220000;
      7802: inst = 32'h10408000;
      7803: inst = 32'hc404c23;
      7804: inst = 32'h8220000;
      7805: inst = 32'h10408000;
      7806: inst = 32'hc404c24;
      7807: inst = 32'h8220000;
      7808: inst = 32'h10408000;
      7809: inst = 32'hc404c25;
      7810: inst = 32'h8220000;
      7811: inst = 32'hc20ffff;
      7812: inst = 32'h10408000;
      7813: inst = 32'hc40423c;
      7814: inst = 32'h8220000;
      7815: inst = 32'h10408000;
      7816: inst = 32'hc40423d;
      7817: inst = 32'h8220000;
      7818: inst = 32'h10408000;
      7819: inst = 32'hc40423e;
      7820: inst = 32'h8220000;
      7821: inst = 32'h10408000;
      7822: inst = 32'hc40423f;
      7823: inst = 32'h8220000;
      7824: inst = 32'h10408000;
      7825: inst = 32'hc404240;
      7826: inst = 32'h8220000;
      7827: inst = 32'h10408000;
      7828: inst = 32'hc404241;
      7829: inst = 32'h8220000;
      7830: inst = 32'h10408000;
      7831: inst = 32'hc404242;
      7832: inst = 32'h8220000;
      7833: inst = 32'h10408000;
      7834: inst = 32'hc404243;
      7835: inst = 32'h8220000;
      7836: inst = 32'h10408000;
      7837: inst = 32'hc404244;
      7838: inst = 32'h8220000;
      7839: inst = 32'h10408000;
      7840: inst = 32'hc404245;
      7841: inst = 32'h8220000;
      7842: inst = 32'h10408000;
      7843: inst = 32'hc404246;
      7844: inst = 32'h8220000;
      7845: inst = 32'h10408000;
      7846: inst = 32'hc404247;
      7847: inst = 32'h8220000;
      7848: inst = 32'h10408000;
      7849: inst = 32'hc404248;
      7850: inst = 32'h8220000;
      7851: inst = 32'h10408000;
      7852: inst = 32'hc404249;
      7853: inst = 32'h8220000;
      7854: inst = 32'h10408000;
      7855: inst = 32'hc40424a;
      7856: inst = 32'h8220000;
      7857: inst = 32'h10408000;
      7858: inst = 32'hc40424b;
      7859: inst = 32'h8220000;
      7860: inst = 32'h10408000;
      7861: inst = 32'hc40424c;
      7862: inst = 32'h8220000;
      7863: inst = 32'h10408000;
      7864: inst = 32'hc40424d;
      7865: inst = 32'h8220000;
      7866: inst = 32'h10408000;
      7867: inst = 32'hc40424e;
      7868: inst = 32'h8220000;
      7869: inst = 32'h10408000;
      7870: inst = 32'hc40424f;
      7871: inst = 32'h8220000;
      7872: inst = 32'h10408000;
      7873: inst = 32'hc404250;
      7874: inst = 32'h8220000;
      7875: inst = 32'h10408000;
      7876: inst = 32'hc404251;
      7877: inst = 32'h8220000;
      7878: inst = 32'h10408000;
      7879: inst = 32'hc404252;
      7880: inst = 32'h8220000;
      7881: inst = 32'h10408000;
      7882: inst = 32'hc404253;
      7883: inst = 32'h8220000;
      7884: inst = 32'h10408000;
      7885: inst = 32'hc404254;
      7886: inst = 32'h8220000;
      7887: inst = 32'h10408000;
      7888: inst = 32'hc404255;
      7889: inst = 32'h8220000;
      7890: inst = 32'h10408000;
      7891: inst = 32'hc404256;
      7892: inst = 32'h8220000;
      7893: inst = 32'h10408000;
      7894: inst = 32'hc404257;
      7895: inst = 32'h8220000;
      7896: inst = 32'h10408000;
      7897: inst = 32'hc404258;
      7898: inst = 32'h8220000;
      7899: inst = 32'h10408000;
      7900: inst = 32'hc404259;
      7901: inst = 32'h8220000;
      7902: inst = 32'h10408000;
      7903: inst = 32'hc40425a;
      7904: inst = 32'h8220000;
      7905: inst = 32'h10408000;
      7906: inst = 32'hc40425b;
      7907: inst = 32'h8220000;
      7908: inst = 32'h10408000;
      7909: inst = 32'hc40425c;
      7910: inst = 32'h8220000;
      7911: inst = 32'h10408000;
      7912: inst = 32'hc40425d;
      7913: inst = 32'h8220000;
      7914: inst = 32'h10408000;
      7915: inst = 32'hc40425e;
      7916: inst = 32'h8220000;
      7917: inst = 32'h10408000;
      7918: inst = 32'hc40425f;
      7919: inst = 32'h8220000;
      7920: inst = 32'h10408000;
      7921: inst = 32'hc404260;
      7922: inst = 32'h8220000;
      7923: inst = 32'h10408000;
      7924: inst = 32'hc404261;
      7925: inst = 32'h8220000;
      7926: inst = 32'h10408000;
      7927: inst = 32'hc404262;
      7928: inst = 32'h8220000;
      7929: inst = 32'h10408000;
      7930: inst = 32'hc404263;
      7931: inst = 32'h8220000;
      7932: inst = 32'h10408000;
      7933: inst = 32'hc40429c;
      7934: inst = 32'h8220000;
      7935: inst = 32'h10408000;
      7936: inst = 32'hc40429d;
      7937: inst = 32'h8220000;
      7938: inst = 32'h10408000;
      7939: inst = 32'hc40429e;
      7940: inst = 32'h8220000;
      7941: inst = 32'h10408000;
      7942: inst = 32'hc40429f;
      7943: inst = 32'h8220000;
      7944: inst = 32'h10408000;
      7945: inst = 32'hc4042a0;
      7946: inst = 32'h8220000;
      7947: inst = 32'h10408000;
      7948: inst = 32'hc4042a1;
      7949: inst = 32'h8220000;
      7950: inst = 32'h10408000;
      7951: inst = 32'hc4042a2;
      7952: inst = 32'h8220000;
      7953: inst = 32'h10408000;
      7954: inst = 32'hc4042a3;
      7955: inst = 32'h8220000;
      7956: inst = 32'h10408000;
      7957: inst = 32'hc4042a4;
      7958: inst = 32'h8220000;
      7959: inst = 32'h10408000;
      7960: inst = 32'hc4042a5;
      7961: inst = 32'h8220000;
      7962: inst = 32'h10408000;
      7963: inst = 32'hc4042a6;
      7964: inst = 32'h8220000;
      7965: inst = 32'h10408000;
      7966: inst = 32'hc4042a7;
      7967: inst = 32'h8220000;
      7968: inst = 32'h10408000;
      7969: inst = 32'hc4042a8;
      7970: inst = 32'h8220000;
      7971: inst = 32'h10408000;
      7972: inst = 32'hc4042a9;
      7973: inst = 32'h8220000;
      7974: inst = 32'h10408000;
      7975: inst = 32'hc4042aa;
      7976: inst = 32'h8220000;
      7977: inst = 32'h10408000;
      7978: inst = 32'hc4042ab;
      7979: inst = 32'h8220000;
      7980: inst = 32'h10408000;
      7981: inst = 32'hc4042ac;
      7982: inst = 32'h8220000;
      7983: inst = 32'h10408000;
      7984: inst = 32'hc4042ad;
      7985: inst = 32'h8220000;
      7986: inst = 32'h10408000;
      7987: inst = 32'hc4042ae;
      7988: inst = 32'h8220000;
      7989: inst = 32'h10408000;
      7990: inst = 32'hc4042af;
      7991: inst = 32'h8220000;
      7992: inst = 32'h10408000;
      7993: inst = 32'hc4042b0;
      7994: inst = 32'h8220000;
      7995: inst = 32'h10408000;
      7996: inst = 32'hc4042b1;
      7997: inst = 32'h8220000;
      7998: inst = 32'h10408000;
      7999: inst = 32'hc4042b2;
      8000: inst = 32'h8220000;
      8001: inst = 32'h10408000;
      8002: inst = 32'hc4042b3;
      8003: inst = 32'h8220000;
      8004: inst = 32'h10408000;
      8005: inst = 32'hc4042b4;
      8006: inst = 32'h8220000;
      8007: inst = 32'h10408000;
      8008: inst = 32'hc4042b5;
      8009: inst = 32'h8220000;
      8010: inst = 32'h10408000;
      8011: inst = 32'hc4042b6;
      8012: inst = 32'h8220000;
      8013: inst = 32'h10408000;
      8014: inst = 32'hc4042b7;
      8015: inst = 32'h8220000;
      8016: inst = 32'h10408000;
      8017: inst = 32'hc4042b8;
      8018: inst = 32'h8220000;
      8019: inst = 32'h10408000;
      8020: inst = 32'hc4042b9;
      8021: inst = 32'h8220000;
      8022: inst = 32'h10408000;
      8023: inst = 32'hc4042ba;
      8024: inst = 32'h8220000;
      8025: inst = 32'h10408000;
      8026: inst = 32'hc4042bb;
      8027: inst = 32'h8220000;
      8028: inst = 32'h10408000;
      8029: inst = 32'hc4042bc;
      8030: inst = 32'h8220000;
      8031: inst = 32'h10408000;
      8032: inst = 32'hc4042bd;
      8033: inst = 32'h8220000;
      8034: inst = 32'h10408000;
      8035: inst = 32'hc4042be;
      8036: inst = 32'h8220000;
      8037: inst = 32'h10408000;
      8038: inst = 32'hc4042bf;
      8039: inst = 32'h8220000;
      8040: inst = 32'h10408000;
      8041: inst = 32'hc4042c0;
      8042: inst = 32'h8220000;
      8043: inst = 32'h10408000;
      8044: inst = 32'hc4042c1;
      8045: inst = 32'h8220000;
      8046: inst = 32'h10408000;
      8047: inst = 32'hc4042c2;
      8048: inst = 32'h8220000;
      8049: inst = 32'h10408000;
      8050: inst = 32'hc4042c3;
      8051: inst = 32'h8220000;
      8052: inst = 32'h10408000;
      8053: inst = 32'hc4042fc;
      8054: inst = 32'h8220000;
      8055: inst = 32'h10408000;
      8056: inst = 32'hc4042fd;
      8057: inst = 32'h8220000;
      8058: inst = 32'h10408000;
      8059: inst = 32'hc4042fe;
      8060: inst = 32'h8220000;
      8061: inst = 32'h10408000;
      8062: inst = 32'hc4042ff;
      8063: inst = 32'h8220000;
      8064: inst = 32'h10408000;
      8065: inst = 32'hc404300;
      8066: inst = 32'h8220000;
      8067: inst = 32'h10408000;
      8068: inst = 32'hc404301;
      8069: inst = 32'h8220000;
      8070: inst = 32'h10408000;
      8071: inst = 32'hc404302;
      8072: inst = 32'h8220000;
      8073: inst = 32'h10408000;
      8074: inst = 32'hc404303;
      8075: inst = 32'h8220000;
      8076: inst = 32'h10408000;
      8077: inst = 32'hc404304;
      8078: inst = 32'h8220000;
      8079: inst = 32'h10408000;
      8080: inst = 32'hc404305;
      8081: inst = 32'h8220000;
      8082: inst = 32'h10408000;
      8083: inst = 32'hc404306;
      8084: inst = 32'h8220000;
      8085: inst = 32'h10408000;
      8086: inst = 32'hc404307;
      8087: inst = 32'h8220000;
      8088: inst = 32'h10408000;
      8089: inst = 32'hc404308;
      8090: inst = 32'h8220000;
      8091: inst = 32'h10408000;
      8092: inst = 32'hc404309;
      8093: inst = 32'h8220000;
      8094: inst = 32'h10408000;
      8095: inst = 32'hc40430a;
      8096: inst = 32'h8220000;
      8097: inst = 32'h10408000;
      8098: inst = 32'hc40430b;
      8099: inst = 32'h8220000;
      8100: inst = 32'h10408000;
      8101: inst = 32'hc40430c;
      8102: inst = 32'h8220000;
      8103: inst = 32'h10408000;
      8104: inst = 32'hc40430d;
      8105: inst = 32'h8220000;
      8106: inst = 32'h10408000;
      8107: inst = 32'hc40430e;
      8108: inst = 32'h8220000;
      8109: inst = 32'h10408000;
      8110: inst = 32'hc40430f;
      8111: inst = 32'h8220000;
      8112: inst = 32'h10408000;
      8113: inst = 32'hc404310;
      8114: inst = 32'h8220000;
      8115: inst = 32'h10408000;
      8116: inst = 32'hc404311;
      8117: inst = 32'h8220000;
      8118: inst = 32'h10408000;
      8119: inst = 32'hc404312;
      8120: inst = 32'h8220000;
      8121: inst = 32'h10408000;
      8122: inst = 32'hc404313;
      8123: inst = 32'h8220000;
      8124: inst = 32'h10408000;
      8125: inst = 32'hc404314;
      8126: inst = 32'h8220000;
      8127: inst = 32'h10408000;
      8128: inst = 32'hc404315;
      8129: inst = 32'h8220000;
      8130: inst = 32'h10408000;
      8131: inst = 32'hc404316;
      8132: inst = 32'h8220000;
      8133: inst = 32'h10408000;
      8134: inst = 32'hc404317;
      8135: inst = 32'h8220000;
      8136: inst = 32'h10408000;
      8137: inst = 32'hc404318;
      8138: inst = 32'h8220000;
      8139: inst = 32'h10408000;
      8140: inst = 32'hc404319;
      8141: inst = 32'h8220000;
      8142: inst = 32'h10408000;
      8143: inst = 32'hc40431a;
      8144: inst = 32'h8220000;
      8145: inst = 32'h10408000;
      8146: inst = 32'hc40431b;
      8147: inst = 32'h8220000;
      8148: inst = 32'h10408000;
      8149: inst = 32'hc40431c;
      8150: inst = 32'h8220000;
      8151: inst = 32'h10408000;
      8152: inst = 32'hc40431d;
      8153: inst = 32'h8220000;
      8154: inst = 32'h10408000;
      8155: inst = 32'hc40431e;
      8156: inst = 32'h8220000;
      8157: inst = 32'h10408000;
      8158: inst = 32'hc40431f;
      8159: inst = 32'h8220000;
      8160: inst = 32'h10408000;
      8161: inst = 32'hc404320;
      8162: inst = 32'h8220000;
      8163: inst = 32'h10408000;
      8164: inst = 32'hc404321;
      8165: inst = 32'h8220000;
      8166: inst = 32'h10408000;
      8167: inst = 32'hc404322;
      8168: inst = 32'h8220000;
      8169: inst = 32'h10408000;
      8170: inst = 32'hc404323;
      8171: inst = 32'h8220000;
      8172: inst = 32'h10408000;
      8173: inst = 32'hc40435c;
      8174: inst = 32'h8220000;
      8175: inst = 32'h10408000;
      8176: inst = 32'hc40435d;
      8177: inst = 32'h8220000;
      8178: inst = 32'h10408000;
      8179: inst = 32'hc40435e;
      8180: inst = 32'h8220000;
      8181: inst = 32'h10408000;
      8182: inst = 32'hc40435f;
      8183: inst = 32'h8220000;
      8184: inst = 32'h10408000;
      8185: inst = 32'hc404360;
      8186: inst = 32'h8220000;
      8187: inst = 32'h10408000;
      8188: inst = 32'hc404361;
      8189: inst = 32'h8220000;
      8190: inst = 32'h10408000;
      8191: inst = 32'hc404362;
      8192: inst = 32'h8220000;
      8193: inst = 32'h10408000;
      8194: inst = 32'hc404363;
      8195: inst = 32'h8220000;
      8196: inst = 32'h10408000;
      8197: inst = 32'hc404364;
      8198: inst = 32'h8220000;
      8199: inst = 32'h10408000;
      8200: inst = 32'hc404365;
      8201: inst = 32'h8220000;
      8202: inst = 32'h10408000;
      8203: inst = 32'hc404366;
      8204: inst = 32'h8220000;
      8205: inst = 32'h10408000;
      8206: inst = 32'hc404367;
      8207: inst = 32'h8220000;
      8208: inst = 32'h10408000;
      8209: inst = 32'hc404368;
      8210: inst = 32'h8220000;
      8211: inst = 32'h10408000;
      8212: inst = 32'hc404369;
      8213: inst = 32'h8220000;
      8214: inst = 32'h10408000;
      8215: inst = 32'hc40436a;
      8216: inst = 32'h8220000;
      8217: inst = 32'h10408000;
      8218: inst = 32'hc40436b;
      8219: inst = 32'h8220000;
      8220: inst = 32'h10408000;
      8221: inst = 32'hc40436c;
      8222: inst = 32'h8220000;
      8223: inst = 32'h10408000;
      8224: inst = 32'hc40436d;
      8225: inst = 32'h8220000;
      8226: inst = 32'h10408000;
      8227: inst = 32'hc40436e;
      8228: inst = 32'h8220000;
      8229: inst = 32'h10408000;
      8230: inst = 32'hc40436f;
      8231: inst = 32'h8220000;
      8232: inst = 32'h10408000;
      8233: inst = 32'hc404370;
      8234: inst = 32'h8220000;
      8235: inst = 32'h10408000;
      8236: inst = 32'hc404371;
      8237: inst = 32'h8220000;
      8238: inst = 32'h10408000;
      8239: inst = 32'hc404372;
      8240: inst = 32'h8220000;
      8241: inst = 32'h10408000;
      8242: inst = 32'hc404373;
      8243: inst = 32'h8220000;
      8244: inst = 32'h10408000;
      8245: inst = 32'hc404374;
      8246: inst = 32'h8220000;
      8247: inst = 32'h10408000;
      8248: inst = 32'hc404375;
      8249: inst = 32'h8220000;
      8250: inst = 32'h10408000;
      8251: inst = 32'hc404376;
      8252: inst = 32'h8220000;
      8253: inst = 32'h10408000;
      8254: inst = 32'hc404377;
      8255: inst = 32'h8220000;
      8256: inst = 32'h10408000;
      8257: inst = 32'hc404378;
      8258: inst = 32'h8220000;
      8259: inst = 32'h10408000;
      8260: inst = 32'hc404379;
      8261: inst = 32'h8220000;
      8262: inst = 32'h10408000;
      8263: inst = 32'hc40437a;
      8264: inst = 32'h8220000;
      8265: inst = 32'h10408000;
      8266: inst = 32'hc40437b;
      8267: inst = 32'h8220000;
      8268: inst = 32'h10408000;
      8269: inst = 32'hc40437c;
      8270: inst = 32'h8220000;
      8271: inst = 32'h10408000;
      8272: inst = 32'hc40437d;
      8273: inst = 32'h8220000;
      8274: inst = 32'h10408000;
      8275: inst = 32'hc40437e;
      8276: inst = 32'h8220000;
      8277: inst = 32'h10408000;
      8278: inst = 32'hc40437f;
      8279: inst = 32'h8220000;
      8280: inst = 32'h10408000;
      8281: inst = 32'hc404380;
      8282: inst = 32'h8220000;
      8283: inst = 32'h10408000;
      8284: inst = 32'hc404381;
      8285: inst = 32'h8220000;
      8286: inst = 32'h10408000;
      8287: inst = 32'hc404382;
      8288: inst = 32'h8220000;
      8289: inst = 32'h10408000;
      8290: inst = 32'hc404383;
      8291: inst = 32'h8220000;
      8292: inst = 32'h10408000;
      8293: inst = 32'hc4043bc;
      8294: inst = 32'h8220000;
      8295: inst = 32'h10408000;
      8296: inst = 32'hc4043bd;
      8297: inst = 32'h8220000;
      8298: inst = 32'h10408000;
      8299: inst = 32'hc4043be;
      8300: inst = 32'h8220000;
      8301: inst = 32'h10408000;
      8302: inst = 32'hc4043bf;
      8303: inst = 32'h8220000;
      8304: inst = 32'h10408000;
      8305: inst = 32'hc4043c0;
      8306: inst = 32'h8220000;
      8307: inst = 32'h10408000;
      8308: inst = 32'hc4043c1;
      8309: inst = 32'h8220000;
      8310: inst = 32'h10408000;
      8311: inst = 32'hc4043c2;
      8312: inst = 32'h8220000;
      8313: inst = 32'h10408000;
      8314: inst = 32'hc4043c3;
      8315: inst = 32'h8220000;
      8316: inst = 32'h10408000;
      8317: inst = 32'hc4043c4;
      8318: inst = 32'h8220000;
      8319: inst = 32'h10408000;
      8320: inst = 32'hc4043c5;
      8321: inst = 32'h8220000;
      8322: inst = 32'h10408000;
      8323: inst = 32'hc4043c6;
      8324: inst = 32'h8220000;
      8325: inst = 32'h10408000;
      8326: inst = 32'hc4043c7;
      8327: inst = 32'h8220000;
      8328: inst = 32'h10408000;
      8329: inst = 32'hc4043c8;
      8330: inst = 32'h8220000;
      8331: inst = 32'h10408000;
      8332: inst = 32'hc4043c9;
      8333: inst = 32'h8220000;
      8334: inst = 32'h10408000;
      8335: inst = 32'hc4043ca;
      8336: inst = 32'h8220000;
      8337: inst = 32'h10408000;
      8338: inst = 32'hc4043cb;
      8339: inst = 32'h8220000;
      8340: inst = 32'h10408000;
      8341: inst = 32'hc4043cc;
      8342: inst = 32'h8220000;
      8343: inst = 32'h10408000;
      8344: inst = 32'hc4043cd;
      8345: inst = 32'h8220000;
      8346: inst = 32'h10408000;
      8347: inst = 32'hc4043ce;
      8348: inst = 32'h8220000;
      8349: inst = 32'h10408000;
      8350: inst = 32'hc4043cf;
      8351: inst = 32'h8220000;
      8352: inst = 32'h10408000;
      8353: inst = 32'hc4043d0;
      8354: inst = 32'h8220000;
      8355: inst = 32'h10408000;
      8356: inst = 32'hc4043d1;
      8357: inst = 32'h8220000;
      8358: inst = 32'h10408000;
      8359: inst = 32'hc4043d2;
      8360: inst = 32'h8220000;
      8361: inst = 32'h10408000;
      8362: inst = 32'hc4043d3;
      8363: inst = 32'h8220000;
      8364: inst = 32'h10408000;
      8365: inst = 32'hc4043d4;
      8366: inst = 32'h8220000;
      8367: inst = 32'h10408000;
      8368: inst = 32'hc4043d5;
      8369: inst = 32'h8220000;
      8370: inst = 32'h10408000;
      8371: inst = 32'hc4043d6;
      8372: inst = 32'h8220000;
      8373: inst = 32'h10408000;
      8374: inst = 32'hc4043d7;
      8375: inst = 32'h8220000;
      8376: inst = 32'h10408000;
      8377: inst = 32'hc4043d8;
      8378: inst = 32'h8220000;
      8379: inst = 32'h10408000;
      8380: inst = 32'hc4043d9;
      8381: inst = 32'h8220000;
      8382: inst = 32'h10408000;
      8383: inst = 32'hc4043da;
      8384: inst = 32'h8220000;
      8385: inst = 32'h10408000;
      8386: inst = 32'hc4043db;
      8387: inst = 32'h8220000;
      8388: inst = 32'h10408000;
      8389: inst = 32'hc4043dc;
      8390: inst = 32'h8220000;
      8391: inst = 32'h10408000;
      8392: inst = 32'hc4043dd;
      8393: inst = 32'h8220000;
      8394: inst = 32'h10408000;
      8395: inst = 32'hc4043de;
      8396: inst = 32'h8220000;
      8397: inst = 32'h10408000;
      8398: inst = 32'hc4043df;
      8399: inst = 32'h8220000;
      8400: inst = 32'h10408000;
      8401: inst = 32'hc4043e0;
      8402: inst = 32'h8220000;
      8403: inst = 32'h10408000;
      8404: inst = 32'hc4043e1;
      8405: inst = 32'h8220000;
      8406: inst = 32'h10408000;
      8407: inst = 32'hc4043e2;
      8408: inst = 32'h8220000;
      8409: inst = 32'h10408000;
      8410: inst = 32'hc4043e3;
      8411: inst = 32'h8220000;
      8412: inst = 32'h10408000;
      8413: inst = 32'hc40441c;
      8414: inst = 32'h8220000;
      8415: inst = 32'h10408000;
      8416: inst = 32'hc40441d;
      8417: inst = 32'h8220000;
      8418: inst = 32'h10408000;
      8419: inst = 32'hc40441e;
      8420: inst = 32'h8220000;
      8421: inst = 32'h10408000;
      8422: inst = 32'hc40441f;
      8423: inst = 32'h8220000;
      8424: inst = 32'h10408000;
      8425: inst = 32'hc404420;
      8426: inst = 32'h8220000;
      8427: inst = 32'h10408000;
      8428: inst = 32'hc404421;
      8429: inst = 32'h8220000;
      8430: inst = 32'h10408000;
      8431: inst = 32'hc404422;
      8432: inst = 32'h8220000;
      8433: inst = 32'h10408000;
      8434: inst = 32'hc404423;
      8435: inst = 32'h8220000;
      8436: inst = 32'h10408000;
      8437: inst = 32'hc404424;
      8438: inst = 32'h8220000;
      8439: inst = 32'h10408000;
      8440: inst = 32'hc404425;
      8441: inst = 32'h8220000;
      8442: inst = 32'h10408000;
      8443: inst = 32'hc404426;
      8444: inst = 32'h8220000;
      8445: inst = 32'h10408000;
      8446: inst = 32'hc404427;
      8447: inst = 32'h8220000;
      8448: inst = 32'h10408000;
      8449: inst = 32'hc404428;
      8450: inst = 32'h8220000;
      8451: inst = 32'h10408000;
      8452: inst = 32'hc404429;
      8453: inst = 32'h8220000;
      8454: inst = 32'h10408000;
      8455: inst = 32'hc40442a;
      8456: inst = 32'h8220000;
      8457: inst = 32'h10408000;
      8458: inst = 32'hc40442b;
      8459: inst = 32'h8220000;
      8460: inst = 32'h10408000;
      8461: inst = 32'hc40442c;
      8462: inst = 32'h8220000;
      8463: inst = 32'h10408000;
      8464: inst = 32'hc40442d;
      8465: inst = 32'h8220000;
      8466: inst = 32'h10408000;
      8467: inst = 32'hc40442e;
      8468: inst = 32'h8220000;
      8469: inst = 32'h10408000;
      8470: inst = 32'hc40442f;
      8471: inst = 32'h8220000;
      8472: inst = 32'h10408000;
      8473: inst = 32'hc404430;
      8474: inst = 32'h8220000;
      8475: inst = 32'h10408000;
      8476: inst = 32'hc404431;
      8477: inst = 32'h8220000;
      8478: inst = 32'h10408000;
      8479: inst = 32'hc404432;
      8480: inst = 32'h8220000;
      8481: inst = 32'h10408000;
      8482: inst = 32'hc404433;
      8483: inst = 32'h8220000;
      8484: inst = 32'h10408000;
      8485: inst = 32'hc404434;
      8486: inst = 32'h8220000;
      8487: inst = 32'h10408000;
      8488: inst = 32'hc404435;
      8489: inst = 32'h8220000;
      8490: inst = 32'h10408000;
      8491: inst = 32'hc404436;
      8492: inst = 32'h8220000;
      8493: inst = 32'h10408000;
      8494: inst = 32'hc404437;
      8495: inst = 32'h8220000;
      8496: inst = 32'h10408000;
      8497: inst = 32'hc404438;
      8498: inst = 32'h8220000;
      8499: inst = 32'h10408000;
      8500: inst = 32'hc404439;
      8501: inst = 32'h8220000;
      8502: inst = 32'h10408000;
      8503: inst = 32'hc40443a;
      8504: inst = 32'h8220000;
      8505: inst = 32'h10408000;
      8506: inst = 32'hc40443b;
      8507: inst = 32'h8220000;
      8508: inst = 32'h10408000;
      8509: inst = 32'hc40443c;
      8510: inst = 32'h8220000;
      8511: inst = 32'h10408000;
      8512: inst = 32'hc40443d;
      8513: inst = 32'h8220000;
      8514: inst = 32'h10408000;
      8515: inst = 32'hc40443e;
      8516: inst = 32'h8220000;
      8517: inst = 32'h10408000;
      8518: inst = 32'hc40443f;
      8519: inst = 32'h8220000;
      8520: inst = 32'h10408000;
      8521: inst = 32'hc404440;
      8522: inst = 32'h8220000;
      8523: inst = 32'h10408000;
      8524: inst = 32'hc404441;
      8525: inst = 32'h8220000;
      8526: inst = 32'h10408000;
      8527: inst = 32'hc404442;
      8528: inst = 32'h8220000;
      8529: inst = 32'h10408000;
      8530: inst = 32'hc404443;
      8531: inst = 32'h8220000;
      8532: inst = 32'h10408000;
      8533: inst = 32'hc40447c;
      8534: inst = 32'h8220000;
      8535: inst = 32'h10408000;
      8536: inst = 32'hc40447d;
      8537: inst = 32'h8220000;
      8538: inst = 32'h10408000;
      8539: inst = 32'hc40447e;
      8540: inst = 32'h8220000;
      8541: inst = 32'h10408000;
      8542: inst = 32'hc40447f;
      8543: inst = 32'h8220000;
      8544: inst = 32'h10408000;
      8545: inst = 32'hc404480;
      8546: inst = 32'h8220000;
      8547: inst = 32'h10408000;
      8548: inst = 32'hc404481;
      8549: inst = 32'h8220000;
      8550: inst = 32'h10408000;
      8551: inst = 32'hc404482;
      8552: inst = 32'h8220000;
      8553: inst = 32'h10408000;
      8554: inst = 32'hc404483;
      8555: inst = 32'h8220000;
      8556: inst = 32'h10408000;
      8557: inst = 32'hc404484;
      8558: inst = 32'h8220000;
      8559: inst = 32'h10408000;
      8560: inst = 32'hc404485;
      8561: inst = 32'h8220000;
      8562: inst = 32'h10408000;
      8563: inst = 32'hc404486;
      8564: inst = 32'h8220000;
      8565: inst = 32'h10408000;
      8566: inst = 32'hc404487;
      8567: inst = 32'h8220000;
      8568: inst = 32'h10408000;
      8569: inst = 32'hc404488;
      8570: inst = 32'h8220000;
      8571: inst = 32'h10408000;
      8572: inst = 32'hc404489;
      8573: inst = 32'h8220000;
      8574: inst = 32'h10408000;
      8575: inst = 32'hc40448a;
      8576: inst = 32'h8220000;
      8577: inst = 32'h10408000;
      8578: inst = 32'hc40448b;
      8579: inst = 32'h8220000;
      8580: inst = 32'h10408000;
      8581: inst = 32'hc40448c;
      8582: inst = 32'h8220000;
      8583: inst = 32'h10408000;
      8584: inst = 32'hc40448d;
      8585: inst = 32'h8220000;
      8586: inst = 32'h10408000;
      8587: inst = 32'hc40448e;
      8588: inst = 32'h8220000;
      8589: inst = 32'h10408000;
      8590: inst = 32'hc40448f;
      8591: inst = 32'h8220000;
      8592: inst = 32'h10408000;
      8593: inst = 32'hc404490;
      8594: inst = 32'h8220000;
      8595: inst = 32'h10408000;
      8596: inst = 32'hc404491;
      8597: inst = 32'h8220000;
      8598: inst = 32'h10408000;
      8599: inst = 32'hc404492;
      8600: inst = 32'h8220000;
      8601: inst = 32'h10408000;
      8602: inst = 32'hc404493;
      8603: inst = 32'h8220000;
      8604: inst = 32'h10408000;
      8605: inst = 32'hc404494;
      8606: inst = 32'h8220000;
      8607: inst = 32'h10408000;
      8608: inst = 32'hc404495;
      8609: inst = 32'h8220000;
      8610: inst = 32'h10408000;
      8611: inst = 32'hc404496;
      8612: inst = 32'h8220000;
      8613: inst = 32'h10408000;
      8614: inst = 32'hc404497;
      8615: inst = 32'h8220000;
      8616: inst = 32'h10408000;
      8617: inst = 32'hc404498;
      8618: inst = 32'h8220000;
      8619: inst = 32'h10408000;
      8620: inst = 32'hc404499;
      8621: inst = 32'h8220000;
      8622: inst = 32'h10408000;
      8623: inst = 32'hc40449a;
      8624: inst = 32'h8220000;
      8625: inst = 32'h10408000;
      8626: inst = 32'hc40449b;
      8627: inst = 32'h8220000;
      8628: inst = 32'h10408000;
      8629: inst = 32'hc40449c;
      8630: inst = 32'h8220000;
      8631: inst = 32'h10408000;
      8632: inst = 32'hc40449d;
      8633: inst = 32'h8220000;
      8634: inst = 32'h10408000;
      8635: inst = 32'hc40449e;
      8636: inst = 32'h8220000;
      8637: inst = 32'h10408000;
      8638: inst = 32'hc40449f;
      8639: inst = 32'h8220000;
      8640: inst = 32'h10408000;
      8641: inst = 32'hc4044a0;
      8642: inst = 32'h8220000;
      8643: inst = 32'h10408000;
      8644: inst = 32'hc4044a1;
      8645: inst = 32'h8220000;
      8646: inst = 32'h10408000;
      8647: inst = 32'hc4044a2;
      8648: inst = 32'h8220000;
      8649: inst = 32'h10408000;
      8650: inst = 32'hc4044a3;
      8651: inst = 32'h8220000;
      8652: inst = 32'h10408000;
      8653: inst = 32'hc4044dc;
      8654: inst = 32'h8220000;
      8655: inst = 32'h10408000;
      8656: inst = 32'hc4044dd;
      8657: inst = 32'h8220000;
      8658: inst = 32'h10408000;
      8659: inst = 32'hc4044de;
      8660: inst = 32'h8220000;
      8661: inst = 32'h10408000;
      8662: inst = 32'hc4044df;
      8663: inst = 32'h8220000;
      8664: inst = 32'h10408000;
      8665: inst = 32'hc4044e0;
      8666: inst = 32'h8220000;
      8667: inst = 32'h10408000;
      8668: inst = 32'hc4044e1;
      8669: inst = 32'h8220000;
      8670: inst = 32'h10408000;
      8671: inst = 32'hc4044e2;
      8672: inst = 32'h8220000;
      8673: inst = 32'h10408000;
      8674: inst = 32'hc4044e3;
      8675: inst = 32'h8220000;
      8676: inst = 32'h10408000;
      8677: inst = 32'hc4044e4;
      8678: inst = 32'h8220000;
      8679: inst = 32'h10408000;
      8680: inst = 32'hc4044e5;
      8681: inst = 32'h8220000;
      8682: inst = 32'h10408000;
      8683: inst = 32'hc4044e6;
      8684: inst = 32'h8220000;
      8685: inst = 32'h10408000;
      8686: inst = 32'hc4044e7;
      8687: inst = 32'h8220000;
      8688: inst = 32'h10408000;
      8689: inst = 32'hc4044e8;
      8690: inst = 32'h8220000;
      8691: inst = 32'h10408000;
      8692: inst = 32'hc4044e9;
      8693: inst = 32'h8220000;
      8694: inst = 32'h10408000;
      8695: inst = 32'hc4044ea;
      8696: inst = 32'h8220000;
      8697: inst = 32'h10408000;
      8698: inst = 32'hc4044eb;
      8699: inst = 32'h8220000;
      8700: inst = 32'h10408000;
      8701: inst = 32'hc4044ec;
      8702: inst = 32'h8220000;
      8703: inst = 32'h10408000;
      8704: inst = 32'hc4044ed;
      8705: inst = 32'h8220000;
      8706: inst = 32'h10408000;
      8707: inst = 32'hc4044ee;
      8708: inst = 32'h8220000;
      8709: inst = 32'h10408000;
      8710: inst = 32'hc4044ef;
      8711: inst = 32'h8220000;
      8712: inst = 32'h10408000;
      8713: inst = 32'hc4044f0;
      8714: inst = 32'h8220000;
      8715: inst = 32'h10408000;
      8716: inst = 32'hc4044f1;
      8717: inst = 32'h8220000;
      8718: inst = 32'h10408000;
      8719: inst = 32'hc4044f2;
      8720: inst = 32'h8220000;
      8721: inst = 32'h10408000;
      8722: inst = 32'hc4044f3;
      8723: inst = 32'h8220000;
      8724: inst = 32'h10408000;
      8725: inst = 32'hc4044f4;
      8726: inst = 32'h8220000;
      8727: inst = 32'h10408000;
      8728: inst = 32'hc4044f5;
      8729: inst = 32'h8220000;
      8730: inst = 32'h10408000;
      8731: inst = 32'hc4044f6;
      8732: inst = 32'h8220000;
      8733: inst = 32'h10408000;
      8734: inst = 32'hc4044f7;
      8735: inst = 32'h8220000;
      8736: inst = 32'h10408000;
      8737: inst = 32'hc4044f8;
      8738: inst = 32'h8220000;
      8739: inst = 32'h10408000;
      8740: inst = 32'hc4044f9;
      8741: inst = 32'h8220000;
      8742: inst = 32'h10408000;
      8743: inst = 32'hc4044fa;
      8744: inst = 32'h8220000;
      8745: inst = 32'h10408000;
      8746: inst = 32'hc4044fb;
      8747: inst = 32'h8220000;
      8748: inst = 32'h10408000;
      8749: inst = 32'hc4044fc;
      8750: inst = 32'h8220000;
      8751: inst = 32'h10408000;
      8752: inst = 32'hc4044fd;
      8753: inst = 32'h8220000;
      8754: inst = 32'h10408000;
      8755: inst = 32'hc4044fe;
      8756: inst = 32'h8220000;
      8757: inst = 32'h10408000;
      8758: inst = 32'hc4044ff;
      8759: inst = 32'h8220000;
      8760: inst = 32'h10408000;
      8761: inst = 32'hc404500;
      8762: inst = 32'h8220000;
      8763: inst = 32'h10408000;
      8764: inst = 32'hc404501;
      8765: inst = 32'h8220000;
      8766: inst = 32'h10408000;
      8767: inst = 32'hc404502;
      8768: inst = 32'h8220000;
      8769: inst = 32'h10408000;
      8770: inst = 32'hc404503;
      8771: inst = 32'h8220000;
      8772: inst = 32'h10408000;
      8773: inst = 32'hc40453c;
      8774: inst = 32'h8220000;
      8775: inst = 32'h10408000;
      8776: inst = 32'hc40453d;
      8777: inst = 32'h8220000;
      8778: inst = 32'h10408000;
      8779: inst = 32'hc40453e;
      8780: inst = 32'h8220000;
      8781: inst = 32'h10408000;
      8782: inst = 32'hc40453f;
      8783: inst = 32'h8220000;
      8784: inst = 32'h10408000;
      8785: inst = 32'hc404540;
      8786: inst = 32'h8220000;
      8787: inst = 32'h10408000;
      8788: inst = 32'hc404541;
      8789: inst = 32'h8220000;
      8790: inst = 32'h10408000;
      8791: inst = 32'hc404542;
      8792: inst = 32'h8220000;
      8793: inst = 32'h10408000;
      8794: inst = 32'hc404543;
      8795: inst = 32'h8220000;
      8796: inst = 32'h10408000;
      8797: inst = 32'hc404544;
      8798: inst = 32'h8220000;
      8799: inst = 32'h10408000;
      8800: inst = 32'hc404545;
      8801: inst = 32'h8220000;
      8802: inst = 32'h10408000;
      8803: inst = 32'hc404546;
      8804: inst = 32'h8220000;
      8805: inst = 32'h10408000;
      8806: inst = 32'hc404547;
      8807: inst = 32'h8220000;
      8808: inst = 32'h10408000;
      8809: inst = 32'hc404548;
      8810: inst = 32'h8220000;
      8811: inst = 32'h10408000;
      8812: inst = 32'hc404549;
      8813: inst = 32'h8220000;
      8814: inst = 32'h10408000;
      8815: inst = 32'hc40454a;
      8816: inst = 32'h8220000;
      8817: inst = 32'h10408000;
      8818: inst = 32'hc40454b;
      8819: inst = 32'h8220000;
      8820: inst = 32'h10408000;
      8821: inst = 32'hc40454c;
      8822: inst = 32'h8220000;
      8823: inst = 32'h10408000;
      8824: inst = 32'hc40454d;
      8825: inst = 32'h8220000;
      8826: inst = 32'h10408000;
      8827: inst = 32'hc40454e;
      8828: inst = 32'h8220000;
      8829: inst = 32'h10408000;
      8830: inst = 32'hc40454f;
      8831: inst = 32'h8220000;
      8832: inst = 32'h10408000;
      8833: inst = 32'hc404550;
      8834: inst = 32'h8220000;
      8835: inst = 32'h10408000;
      8836: inst = 32'hc404551;
      8837: inst = 32'h8220000;
      8838: inst = 32'h10408000;
      8839: inst = 32'hc404552;
      8840: inst = 32'h8220000;
      8841: inst = 32'h10408000;
      8842: inst = 32'hc404553;
      8843: inst = 32'h8220000;
      8844: inst = 32'h10408000;
      8845: inst = 32'hc404554;
      8846: inst = 32'h8220000;
      8847: inst = 32'h10408000;
      8848: inst = 32'hc404555;
      8849: inst = 32'h8220000;
      8850: inst = 32'h10408000;
      8851: inst = 32'hc404556;
      8852: inst = 32'h8220000;
      8853: inst = 32'h10408000;
      8854: inst = 32'hc404557;
      8855: inst = 32'h8220000;
      8856: inst = 32'h10408000;
      8857: inst = 32'hc404558;
      8858: inst = 32'h8220000;
      8859: inst = 32'h10408000;
      8860: inst = 32'hc404559;
      8861: inst = 32'h8220000;
      8862: inst = 32'h10408000;
      8863: inst = 32'hc40455a;
      8864: inst = 32'h8220000;
      8865: inst = 32'h10408000;
      8866: inst = 32'hc40455b;
      8867: inst = 32'h8220000;
      8868: inst = 32'h10408000;
      8869: inst = 32'hc40455c;
      8870: inst = 32'h8220000;
      8871: inst = 32'h10408000;
      8872: inst = 32'hc40455d;
      8873: inst = 32'h8220000;
      8874: inst = 32'h10408000;
      8875: inst = 32'hc40455e;
      8876: inst = 32'h8220000;
      8877: inst = 32'h10408000;
      8878: inst = 32'hc40455f;
      8879: inst = 32'h8220000;
      8880: inst = 32'h10408000;
      8881: inst = 32'hc404560;
      8882: inst = 32'h8220000;
      8883: inst = 32'h10408000;
      8884: inst = 32'hc404561;
      8885: inst = 32'h8220000;
      8886: inst = 32'h10408000;
      8887: inst = 32'hc404562;
      8888: inst = 32'h8220000;
      8889: inst = 32'h10408000;
      8890: inst = 32'hc404563;
      8891: inst = 32'h8220000;
      8892: inst = 32'h10408000;
      8893: inst = 32'hc40459c;
      8894: inst = 32'h8220000;
      8895: inst = 32'h10408000;
      8896: inst = 32'hc40459d;
      8897: inst = 32'h8220000;
      8898: inst = 32'h10408000;
      8899: inst = 32'hc40459e;
      8900: inst = 32'h8220000;
      8901: inst = 32'h10408000;
      8902: inst = 32'hc40459f;
      8903: inst = 32'h8220000;
      8904: inst = 32'h10408000;
      8905: inst = 32'hc4045a0;
      8906: inst = 32'h8220000;
      8907: inst = 32'h10408000;
      8908: inst = 32'hc4045a1;
      8909: inst = 32'h8220000;
      8910: inst = 32'h10408000;
      8911: inst = 32'hc4045a2;
      8912: inst = 32'h8220000;
      8913: inst = 32'h10408000;
      8914: inst = 32'hc4045a3;
      8915: inst = 32'h8220000;
      8916: inst = 32'h10408000;
      8917: inst = 32'hc4045a4;
      8918: inst = 32'h8220000;
      8919: inst = 32'h10408000;
      8920: inst = 32'hc4045a5;
      8921: inst = 32'h8220000;
      8922: inst = 32'h10408000;
      8923: inst = 32'hc4045a6;
      8924: inst = 32'h8220000;
      8925: inst = 32'h10408000;
      8926: inst = 32'hc4045a7;
      8927: inst = 32'h8220000;
      8928: inst = 32'h10408000;
      8929: inst = 32'hc4045a8;
      8930: inst = 32'h8220000;
      8931: inst = 32'h10408000;
      8932: inst = 32'hc4045a9;
      8933: inst = 32'h8220000;
      8934: inst = 32'h10408000;
      8935: inst = 32'hc4045aa;
      8936: inst = 32'h8220000;
      8937: inst = 32'h10408000;
      8938: inst = 32'hc4045ab;
      8939: inst = 32'h8220000;
      8940: inst = 32'h10408000;
      8941: inst = 32'hc4045ac;
      8942: inst = 32'h8220000;
      8943: inst = 32'h10408000;
      8944: inst = 32'hc4045ad;
      8945: inst = 32'h8220000;
      8946: inst = 32'h10408000;
      8947: inst = 32'hc4045ae;
      8948: inst = 32'h8220000;
      8949: inst = 32'h10408000;
      8950: inst = 32'hc4045af;
      8951: inst = 32'h8220000;
      8952: inst = 32'h10408000;
      8953: inst = 32'hc4045b0;
      8954: inst = 32'h8220000;
      8955: inst = 32'h10408000;
      8956: inst = 32'hc4045b1;
      8957: inst = 32'h8220000;
      8958: inst = 32'h10408000;
      8959: inst = 32'hc4045b2;
      8960: inst = 32'h8220000;
      8961: inst = 32'h10408000;
      8962: inst = 32'hc4045b3;
      8963: inst = 32'h8220000;
      8964: inst = 32'h10408000;
      8965: inst = 32'hc4045b4;
      8966: inst = 32'h8220000;
      8967: inst = 32'h10408000;
      8968: inst = 32'hc4045b5;
      8969: inst = 32'h8220000;
      8970: inst = 32'h10408000;
      8971: inst = 32'hc4045b6;
      8972: inst = 32'h8220000;
      8973: inst = 32'h10408000;
      8974: inst = 32'hc4045b7;
      8975: inst = 32'h8220000;
      8976: inst = 32'h10408000;
      8977: inst = 32'hc4045b8;
      8978: inst = 32'h8220000;
      8979: inst = 32'h10408000;
      8980: inst = 32'hc4045b9;
      8981: inst = 32'h8220000;
      8982: inst = 32'h10408000;
      8983: inst = 32'hc4045ba;
      8984: inst = 32'h8220000;
      8985: inst = 32'h10408000;
      8986: inst = 32'hc4045bb;
      8987: inst = 32'h8220000;
      8988: inst = 32'h10408000;
      8989: inst = 32'hc4045bc;
      8990: inst = 32'h8220000;
      8991: inst = 32'h10408000;
      8992: inst = 32'hc4045bd;
      8993: inst = 32'h8220000;
      8994: inst = 32'h10408000;
      8995: inst = 32'hc4045be;
      8996: inst = 32'h8220000;
      8997: inst = 32'h10408000;
      8998: inst = 32'hc4045bf;
      8999: inst = 32'h8220000;
      9000: inst = 32'h10408000;
      9001: inst = 32'hc4045c0;
      9002: inst = 32'h8220000;
      9003: inst = 32'h10408000;
      9004: inst = 32'hc4045c1;
      9005: inst = 32'h8220000;
      9006: inst = 32'h10408000;
      9007: inst = 32'hc4045c2;
      9008: inst = 32'h8220000;
      9009: inst = 32'h10408000;
      9010: inst = 32'hc4045c3;
      9011: inst = 32'h8220000;
      9012: inst = 32'h10408000;
      9013: inst = 32'hc4045fc;
      9014: inst = 32'h8220000;
      9015: inst = 32'h10408000;
      9016: inst = 32'hc4045fd;
      9017: inst = 32'h8220000;
      9018: inst = 32'h10408000;
      9019: inst = 32'hc4045fe;
      9020: inst = 32'h8220000;
      9021: inst = 32'h10408000;
      9022: inst = 32'hc4045ff;
      9023: inst = 32'h8220000;
      9024: inst = 32'h10408000;
      9025: inst = 32'hc404600;
      9026: inst = 32'h8220000;
      9027: inst = 32'h10408000;
      9028: inst = 32'hc404601;
      9029: inst = 32'h8220000;
      9030: inst = 32'h10408000;
      9031: inst = 32'hc404602;
      9032: inst = 32'h8220000;
      9033: inst = 32'h10408000;
      9034: inst = 32'hc404603;
      9035: inst = 32'h8220000;
      9036: inst = 32'h10408000;
      9037: inst = 32'hc404604;
      9038: inst = 32'h8220000;
      9039: inst = 32'h10408000;
      9040: inst = 32'hc404605;
      9041: inst = 32'h8220000;
      9042: inst = 32'h10408000;
      9043: inst = 32'hc404606;
      9044: inst = 32'h8220000;
      9045: inst = 32'h10408000;
      9046: inst = 32'hc404607;
      9047: inst = 32'h8220000;
      9048: inst = 32'h10408000;
      9049: inst = 32'hc404608;
      9050: inst = 32'h8220000;
      9051: inst = 32'h10408000;
      9052: inst = 32'hc404609;
      9053: inst = 32'h8220000;
      9054: inst = 32'h10408000;
      9055: inst = 32'hc40460a;
      9056: inst = 32'h8220000;
      9057: inst = 32'h10408000;
      9058: inst = 32'hc40460b;
      9059: inst = 32'h8220000;
      9060: inst = 32'h10408000;
      9061: inst = 32'hc40460c;
      9062: inst = 32'h8220000;
      9063: inst = 32'h10408000;
      9064: inst = 32'hc40460d;
      9065: inst = 32'h8220000;
      9066: inst = 32'h10408000;
      9067: inst = 32'hc40460e;
      9068: inst = 32'h8220000;
      9069: inst = 32'h10408000;
      9070: inst = 32'hc40460f;
      9071: inst = 32'h8220000;
      9072: inst = 32'h10408000;
      9073: inst = 32'hc404610;
      9074: inst = 32'h8220000;
      9075: inst = 32'h10408000;
      9076: inst = 32'hc404611;
      9077: inst = 32'h8220000;
      9078: inst = 32'h10408000;
      9079: inst = 32'hc404612;
      9080: inst = 32'h8220000;
      9081: inst = 32'h10408000;
      9082: inst = 32'hc404613;
      9083: inst = 32'h8220000;
      9084: inst = 32'h10408000;
      9085: inst = 32'hc404614;
      9086: inst = 32'h8220000;
      9087: inst = 32'h10408000;
      9088: inst = 32'hc404615;
      9089: inst = 32'h8220000;
      9090: inst = 32'h10408000;
      9091: inst = 32'hc404616;
      9092: inst = 32'h8220000;
      9093: inst = 32'h10408000;
      9094: inst = 32'hc404617;
      9095: inst = 32'h8220000;
      9096: inst = 32'h10408000;
      9097: inst = 32'hc404618;
      9098: inst = 32'h8220000;
      9099: inst = 32'h10408000;
      9100: inst = 32'hc404619;
      9101: inst = 32'h8220000;
      9102: inst = 32'h10408000;
      9103: inst = 32'hc40461a;
      9104: inst = 32'h8220000;
      9105: inst = 32'h10408000;
      9106: inst = 32'hc40461b;
      9107: inst = 32'h8220000;
      9108: inst = 32'h10408000;
      9109: inst = 32'hc40461c;
      9110: inst = 32'h8220000;
      9111: inst = 32'h10408000;
      9112: inst = 32'hc40461d;
      9113: inst = 32'h8220000;
      9114: inst = 32'h10408000;
      9115: inst = 32'hc40461e;
      9116: inst = 32'h8220000;
      9117: inst = 32'h10408000;
      9118: inst = 32'hc40461f;
      9119: inst = 32'h8220000;
      9120: inst = 32'h10408000;
      9121: inst = 32'hc404620;
      9122: inst = 32'h8220000;
      9123: inst = 32'h10408000;
      9124: inst = 32'hc404621;
      9125: inst = 32'h8220000;
      9126: inst = 32'h10408000;
      9127: inst = 32'hc404622;
      9128: inst = 32'h8220000;
      9129: inst = 32'h10408000;
      9130: inst = 32'hc404623;
      9131: inst = 32'h8220000;
      9132: inst = 32'h10408000;
      9133: inst = 32'hc40465c;
      9134: inst = 32'h8220000;
      9135: inst = 32'h10408000;
      9136: inst = 32'hc40465d;
      9137: inst = 32'h8220000;
      9138: inst = 32'h10408000;
      9139: inst = 32'hc40465e;
      9140: inst = 32'h8220000;
      9141: inst = 32'h10408000;
      9142: inst = 32'hc40465f;
      9143: inst = 32'h8220000;
      9144: inst = 32'h10408000;
      9145: inst = 32'hc404660;
      9146: inst = 32'h8220000;
      9147: inst = 32'h10408000;
      9148: inst = 32'hc404661;
      9149: inst = 32'h8220000;
      9150: inst = 32'h10408000;
      9151: inst = 32'hc404662;
      9152: inst = 32'h8220000;
      9153: inst = 32'h10408000;
      9154: inst = 32'hc404663;
      9155: inst = 32'h8220000;
      9156: inst = 32'h10408000;
      9157: inst = 32'hc404664;
      9158: inst = 32'h8220000;
      9159: inst = 32'h10408000;
      9160: inst = 32'hc404665;
      9161: inst = 32'h8220000;
      9162: inst = 32'h10408000;
      9163: inst = 32'hc404666;
      9164: inst = 32'h8220000;
      9165: inst = 32'h10408000;
      9166: inst = 32'hc404667;
      9167: inst = 32'h8220000;
      9168: inst = 32'h10408000;
      9169: inst = 32'hc404668;
      9170: inst = 32'h8220000;
      9171: inst = 32'h10408000;
      9172: inst = 32'hc404669;
      9173: inst = 32'h8220000;
      9174: inst = 32'h10408000;
      9175: inst = 32'hc40466a;
      9176: inst = 32'h8220000;
      9177: inst = 32'h10408000;
      9178: inst = 32'hc40466b;
      9179: inst = 32'h8220000;
      9180: inst = 32'h10408000;
      9181: inst = 32'hc40466c;
      9182: inst = 32'h8220000;
      9183: inst = 32'h10408000;
      9184: inst = 32'hc40466d;
      9185: inst = 32'h8220000;
      9186: inst = 32'h10408000;
      9187: inst = 32'hc40466e;
      9188: inst = 32'h8220000;
      9189: inst = 32'h10408000;
      9190: inst = 32'hc40466f;
      9191: inst = 32'h8220000;
      9192: inst = 32'h10408000;
      9193: inst = 32'hc404670;
      9194: inst = 32'h8220000;
      9195: inst = 32'h10408000;
      9196: inst = 32'hc404671;
      9197: inst = 32'h8220000;
      9198: inst = 32'h10408000;
      9199: inst = 32'hc404672;
      9200: inst = 32'h8220000;
      9201: inst = 32'h10408000;
      9202: inst = 32'hc404673;
      9203: inst = 32'h8220000;
      9204: inst = 32'h10408000;
      9205: inst = 32'hc404674;
      9206: inst = 32'h8220000;
      9207: inst = 32'h10408000;
      9208: inst = 32'hc404675;
      9209: inst = 32'h8220000;
      9210: inst = 32'h10408000;
      9211: inst = 32'hc404676;
      9212: inst = 32'h8220000;
      9213: inst = 32'h10408000;
      9214: inst = 32'hc404677;
      9215: inst = 32'h8220000;
      9216: inst = 32'h10408000;
      9217: inst = 32'hc404678;
      9218: inst = 32'h8220000;
      9219: inst = 32'h10408000;
      9220: inst = 32'hc404679;
      9221: inst = 32'h8220000;
      9222: inst = 32'h10408000;
      9223: inst = 32'hc40467a;
      9224: inst = 32'h8220000;
      9225: inst = 32'h10408000;
      9226: inst = 32'hc40467b;
      9227: inst = 32'h8220000;
      9228: inst = 32'h10408000;
      9229: inst = 32'hc40467c;
      9230: inst = 32'h8220000;
      9231: inst = 32'h10408000;
      9232: inst = 32'hc40467d;
      9233: inst = 32'h8220000;
      9234: inst = 32'h10408000;
      9235: inst = 32'hc40467e;
      9236: inst = 32'h8220000;
      9237: inst = 32'h10408000;
      9238: inst = 32'hc40467f;
      9239: inst = 32'h8220000;
      9240: inst = 32'h10408000;
      9241: inst = 32'hc404680;
      9242: inst = 32'h8220000;
      9243: inst = 32'h10408000;
      9244: inst = 32'hc404681;
      9245: inst = 32'h8220000;
      9246: inst = 32'h10408000;
      9247: inst = 32'hc404682;
      9248: inst = 32'h8220000;
      9249: inst = 32'h10408000;
      9250: inst = 32'hc404683;
      9251: inst = 32'h8220000;
      9252: inst = 32'h10408000;
      9253: inst = 32'hc4046bc;
      9254: inst = 32'h8220000;
      9255: inst = 32'h10408000;
      9256: inst = 32'hc4046bd;
      9257: inst = 32'h8220000;
      9258: inst = 32'h10408000;
      9259: inst = 32'hc4046be;
      9260: inst = 32'h8220000;
      9261: inst = 32'h10408000;
      9262: inst = 32'hc4046bf;
      9263: inst = 32'h8220000;
      9264: inst = 32'h10408000;
      9265: inst = 32'hc4046c0;
      9266: inst = 32'h8220000;
      9267: inst = 32'h10408000;
      9268: inst = 32'hc4046c1;
      9269: inst = 32'h8220000;
      9270: inst = 32'h10408000;
      9271: inst = 32'hc4046c2;
      9272: inst = 32'h8220000;
      9273: inst = 32'h10408000;
      9274: inst = 32'hc4046c3;
      9275: inst = 32'h8220000;
      9276: inst = 32'h10408000;
      9277: inst = 32'hc4046c4;
      9278: inst = 32'h8220000;
      9279: inst = 32'h10408000;
      9280: inst = 32'hc4046c5;
      9281: inst = 32'h8220000;
      9282: inst = 32'h10408000;
      9283: inst = 32'hc4046c6;
      9284: inst = 32'h8220000;
      9285: inst = 32'h10408000;
      9286: inst = 32'hc4046c7;
      9287: inst = 32'h8220000;
      9288: inst = 32'h10408000;
      9289: inst = 32'hc4046c8;
      9290: inst = 32'h8220000;
      9291: inst = 32'h10408000;
      9292: inst = 32'hc4046c9;
      9293: inst = 32'h8220000;
      9294: inst = 32'h10408000;
      9295: inst = 32'hc4046ca;
      9296: inst = 32'h8220000;
      9297: inst = 32'h10408000;
      9298: inst = 32'hc4046cb;
      9299: inst = 32'h8220000;
      9300: inst = 32'h10408000;
      9301: inst = 32'hc4046cc;
      9302: inst = 32'h8220000;
      9303: inst = 32'h10408000;
      9304: inst = 32'hc4046cd;
      9305: inst = 32'h8220000;
      9306: inst = 32'h10408000;
      9307: inst = 32'hc4046ce;
      9308: inst = 32'h8220000;
      9309: inst = 32'h10408000;
      9310: inst = 32'hc4046cf;
      9311: inst = 32'h8220000;
      9312: inst = 32'h10408000;
      9313: inst = 32'hc4046d0;
      9314: inst = 32'h8220000;
      9315: inst = 32'h10408000;
      9316: inst = 32'hc4046d1;
      9317: inst = 32'h8220000;
      9318: inst = 32'h10408000;
      9319: inst = 32'hc4046d2;
      9320: inst = 32'h8220000;
      9321: inst = 32'h10408000;
      9322: inst = 32'hc4046d3;
      9323: inst = 32'h8220000;
      9324: inst = 32'h10408000;
      9325: inst = 32'hc4046d4;
      9326: inst = 32'h8220000;
      9327: inst = 32'h10408000;
      9328: inst = 32'hc4046d5;
      9329: inst = 32'h8220000;
      9330: inst = 32'h10408000;
      9331: inst = 32'hc4046d6;
      9332: inst = 32'h8220000;
      9333: inst = 32'h10408000;
      9334: inst = 32'hc4046d7;
      9335: inst = 32'h8220000;
      9336: inst = 32'h10408000;
      9337: inst = 32'hc4046d8;
      9338: inst = 32'h8220000;
      9339: inst = 32'h10408000;
      9340: inst = 32'hc4046d9;
      9341: inst = 32'h8220000;
      9342: inst = 32'h10408000;
      9343: inst = 32'hc4046da;
      9344: inst = 32'h8220000;
      9345: inst = 32'h10408000;
      9346: inst = 32'hc4046db;
      9347: inst = 32'h8220000;
      9348: inst = 32'h10408000;
      9349: inst = 32'hc4046dc;
      9350: inst = 32'h8220000;
      9351: inst = 32'h10408000;
      9352: inst = 32'hc4046dd;
      9353: inst = 32'h8220000;
      9354: inst = 32'h10408000;
      9355: inst = 32'hc4046de;
      9356: inst = 32'h8220000;
      9357: inst = 32'h10408000;
      9358: inst = 32'hc4046df;
      9359: inst = 32'h8220000;
      9360: inst = 32'h10408000;
      9361: inst = 32'hc4046e0;
      9362: inst = 32'h8220000;
      9363: inst = 32'h10408000;
      9364: inst = 32'hc4046e1;
      9365: inst = 32'h8220000;
      9366: inst = 32'h10408000;
      9367: inst = 32'hc4046e2;
      9368: inst = 32'h8220000;
      9369: inst = 32'h10408000;
      9370: inst = 32'hc4046e3;
      9371: inst = 32'h8220000;
      9372: inst = 32'h10408000;
      9373: inst = 32'hc40471c;
      9374: inst = 32'h8220000;
      9375: inst = 32'h10408000;
      9376: inst = 32'hc40471d;
      9377: inst = 32'h8220000;
      9378: inst = 32'h10408000;
      9379: inst = 32'hc40471e;
      9380: inst = 32'h8220000;
      9381: inst = 32'h10408000;
      9382: inst = 32'hc40471f;
      9383: inst = 32'h8220000;
      9384: inst = 32'h10408000;
      9385: inst = 32'hc404720;
      9386: inst = 32'h8220000;
      9387: inst = 32'h10408000;
      9388: inst = 32'hc404721;
      9389: inst = 32'h8220000;
      9390: inst = 32'h10408000;
      9391: inst = 32'hc404722;
      9392: inst = 32'h8220000;
      9393: inst = 32'h10408000;
      9394: inst = 32'hc404723;
      9395: inst = 32'h8220000;
      9396: inst = 32'h10408000;
      9397: inst = 32'hc404724;
      9398: inst = 32'h8220000;
      9399: inst = 32'h10408000;
      9400: inst = 32'hc404725;
      9401: inst = 32'h8220000;
      9402: inst = 32'h10408000;
      9403: inst = 32'hc404726;
      9404: inst = 32'h8220000;
      9405: inst = 32'h10408000;
      9406: inst = 32'hc404727;
      9407: inst = 32'h8220000;
      9408: inst = 32'h10408000;
      9409: inst = 32'hc404728;
      9410: inst = 32'h8220000;
      9411: inst = 32'h10408000;
      9412: inst = 32'hc404729;
      9413: inst = 32'h8220000;
      9414: inst = 32'h10408000;
      9415: inst = 32'hc40472a;
      9416: inst = 32'h8220000;
      9417: inst = 32'h10408000;
      9418: inst = 32'hc40472b;
      9419: inst = 32'h8220000;
      9420: inst = 32'h10408000;
      9421: inst = 32'hc40472c;
      9422: inst = 32'h8220000;
      9423: inst = 32'h10408000;
      9424: inst = 32'hc40472d;
      9425: inst = 32'h8220000;
      9426: inst = 32'h10408000;
      9427: inst = 32'hc40472e;
      9428: inst = 32'h8220000;
      9429: inst = 32'h10408000;
      9430: inst = 32'hc40472f;
      9431: inst = 32'h8220000;
      9432: inst = 32'h10408000;
      9433: inst = 32'hc404730;
      9434: inst = 32'h8220000;
      9435: inst = 32'h10408000;
      9436: inst = 32'hc404731;
      9437: inst = 32'h8220000;
      9438: inst = 32'h10408000;
      9439: inst = 32'hc404732;
      9440: inst = 32'h8220000;
      9441: inst = 32'h10408000;
      9442: inst = 32'hc404733;
      9443: inst = 32'h8220000;
      9444: inst = 32'h10408000;
      9445: inst = 32'hc404734;
      9446: inst = 32'h8220000;
      9447: inst = 32'h10408000;
      9448: inst = 32'hc404735;
      9449: inst = 32'h8220000;
      9450: inst = 32'h10408000;
      9451: inst = 32'hc404736;
      9452: inst = 32'h8220000;
      9453: inst = 32'h10408000;
      9454: inst = 32'hc404737;
      9455: inst = 32'h8220000;
      9456: inst = 32'h10408000;
      9457: inst = 32'hc404738;
      9458: inst = 32'h8220000;
      9459: inst = 32'h10408000;
      9460: inst = 32'hc404739;
      9461: inst = 32'h8220000;
      9462: inst = 32'h10408000;
      9463: inst = 32'hc40473a;
      9464: inst = 32'h8220000;
      9465: inst = 32'h10408000;
      9466: inst = 32'hc40473b;
      9467: inst = 32'h8220000;
      9468: inst = 32'h10408000;
      9469: inst = 32'hc40473c;
      9470: inst = 32'h8220000;
      9471: inst = 32'h10408000;
      9472: inst = 32'hc40473d;
      9473: inst = 32'h8220000;
      9474: inst = 32'h10408000;
      9475: inst = 32'hc40473e;
      9476: inst = 32'h8220000;
      9477: inst = 32'h10408000;
      9478: inst = 32'hc40473f;
      9479: inst = 32'h8220000;
      9480: inst = 32'h10408000;
      9481: inst = 32'hc404740;
      9482: inst = 32'h8220000;
      9483: inst = 32'h10408000;
      9484: inst = 32'hc404741;
      9485: inst = 32'h8220000;
      9486: inst = 32'h10408000;
      9487: inst = 32'hc404742;
      9488: inst = 32'h8220000;
      9489: inst = 32'h10408000;
      9490: inst = 32'hc404743;
      9491: inst = 32'h8220000;
      9492: inst = 32'h10408000;
      9493: inst = 32'hc40477c;
      9494: inst = 32'h8220000;
      9495: inst = 32'h10408000;
      9496: inst = 32'hc40477d;
      9497: inst = 32'h8220000;
      9498: inst = 32'h10408000;
      9499: inst = 32'hc40477e;
      9500: inst = 32'h8220000;
      9501: inst = 32'h10408000;
      9502: inst = 32'hc40477f;
      9503: inst = 32'h8220000;
      9504: inst = 32'h10408000;
      9505: inst = 32'hc404780;
      9506: inst = 32'h8220000;
      9507: inst = 32'h10408000;
      9508: inst = 32'hc404781;
      9509: inst = 32'h8220000;
      9510: inst = 32'h10408000;
      9511: inst = 32'hc404782;
      9512: inst = 32'h8220000;
      9513: inst = 32'h10408000;
      9514: inst = 32'hc404783;
      9515: inst = 32'h8220000;
      9516: inst = 32'h10408000;
      9517: inst = 32'hc404784;
      9518: inst = 32'h8220000;
      9519: inst = 32'h10408000;
      9520: inst = 32'hc404785;
      9521: inst = 32'h8220000;
      9522: inst = 32'h10408000;
      9523: inst = 32'hc404786;
      9524: inst = 32'h8220000;
      9525: inst = 32'h10408000;
      9526: inst = 32'hc404787;
      9527: inst = 32'h8220000;
      9528: inst = 32'h10408000;
      9529: inst = 32'hc404788;
      9530: inst = 32'h8220000;
      9531: inst = 32'h10408000;
      9532: inst = 32'hc404789;
      9533: inst = 32'h8220000;
      9534: inst = 32'h10408000;
      9535: inst = 32'hc40478a;
      9536: inst = 32'h8220000;
      9537: inst = 32'h10408000;
      9538: inst = 32'hc40478b;
      9539: inst = 32'h8220000;
      9540: inst = 32'h10408000;
      9541: inst = 32'hc40478c;
      9542: inst = 32'h8220000;
      9543: inst = 32'h10408000;
      9544: inst = 32'hc40478d;
      9545: inst = 32'h8220000;
      9546: inst = 32'h10408000;
      9547: inst = 32'hc40478e;
      9548: inst = 32'h8220000;
      9549: inst = 32'h10408000;
      9550: inst = 32'hc40478f;
      9551: inst = 32'h8220000;
      9552: inst = 32'h10408000;
      9553: inst = 32'hc404790;
      9554: inst = 32'h8220000;
      9555: inst = 32'h10408000;
      9556: inst = 32'hc404791;
      9557: inst = 32'h8220000;
      9558: inst = 32'h10408000;
      9559: inst = 32'hc404792;
      9560: inst = 32'h8220000;
      9561: inst = 32'h10408000;
      9562: inst = 32'hc404793;
      9563: inst = 32'h8220000;
      9564: inst = 32'h10408000;
      9565: inst = 32'hc404794;
      9566: inst = 32'h8220000;
      9567: inst = 32'h10408000;
      9568: inst = 32'hc404795;
      9569: inst = 32'h8220000;
      9570: inst = 32'h10408000;
      9571: inst = 32'hc404796;
      9572: inst = 32'h8220000;
      9573: inst = 32'h10408000;
      9574: inst = 32'hc404797;
      9575: inst = 32'h8220000;
      9576: inst = 32'h10408000;
      9577: inst = 32'hc404798;
      9578: inst = 32'h8220000;
      9579: inst = 32'h10408000;
      9580: inst = 32'hc404799;
      9581: inst = 32'h8220000;
      9582: inst = 32'h10408000;
      9583: inst = 32'hc40479a;
      9584: inst = 32'h8220000;
      9585: inst = 32'h10408000;
      9586: inst = 32'hc40479b;
      9587: inst = 32'h8220000;
      9588: inst = 32'h10408000;
      9589: inst = 32'hc40479c;
      9590: inst = 32'h8220000;
      9591: inst = 32'h10408000;
      9592: inst = 32'hc40479d;
      9593: inst = 32'h8220000;
      9594: inst = 32'h10408000;
      9595: inst = 32'hc40479e;
      9596: inst = 32'h8220000;
      9597: inst = 32'h10408000;
      9598: inst = 32'hc40479f;
      9599: inst = 32'h8220000;
      9600: inst = 32'h10408000;
      9601: inst = 32'hc4047a0;
      9602: inst = 32'h8220000;
      9603: inst = 32'h10408000;
      9604: inst = 32'hc4047a1;
      9605: inst = 32'h8220000;
      9606: inst = 32'h10408000;
      9607: inst = 32'hc4047a2;
      9608: inst = 32'h8220000;
      9609: inst = 32'h10408000;
      9610: inst = 32'hc4047a3;
      9611: inst = 32'h8220000;
      9612: inst = 32'h10408000;
      9613: inst = 32'hc4047dc;
      9614: inst = 32'h8220000;
      9615: inst = 32'h10408000;
      9616: inst = 32'hc4047dd;
      9617: inst = 32'h8220000;
      9618: inst = 32'h10408000;
      9619: inst = 32'hc4047de;
      9620: inst = 32'h8220000;
      9621: inst = 32'h10408000;
      9622: inst = 32'hc4047df;
      9623: inst = 32'h8220000;
      9624: inst = 32'h10408000;
      9625: inst = 32'hc4047e0;
      9626: inst = 32'h8220000;
      9627: inst = 32'h10408000;
      9628: inst = 32'hc4047e1;
      9629: inst = 32'h8220000;
      9630: inst = 32'h10408000;
      9631: inst = 32'hc4047e2;
      9632: inst = 32'h8220000;
      9633: inst = 32'h10408000;
      9634: inst = 32'hc4047e3;
      9635: inst = 32'h8220000;
      9636: inst = 32'h10408000;
      9637: inst = 32'hc4047e4;
      9638: inst = 32'h8220000;
      9639: inst = 32'h10408000;
      9640: inst = 32'hc4047e5;
      9641: inst = 32'h8220000;
      9642: inst = 32'h10408000;
      9643: inst = 32'hc4047e6;
      9644: inst = 32'h8220000;
      9645: inst = 32'h10408000;
      9646: inst = 32'hc4047e7;
      9647: inst = 32'h8220000;
      9648: inst = 32'h10408000;
      9649: inst = 32'hc4047e8;
      9650: inst = 32'h8220000;
      9651: inst = 32'h10408000;
      9652: inst = 32'hc4047e9;
      9653: inst = 32'h8220000;
      9654: inst = 32'h10408000;
      9655: inst = 32'hc4047ea;
      9656: inst = 32'h8220000;
      9657: inst = 32'h10408000;
      9658: inst = 32'hc4047eb;
      9659: inst = 32'h8220000;
      9660: inst = 32'h10408000;
      9661: inst = 32'hc4047ec;
      9662: inst = 32'h8220000;
      9663: inst = 32'h10408000;
      9664: inst = 32'hc4047ed;
      9665: inst = 32'h8220000;
      9666: inst = 32'h10408000;
      9667: inst = 32'hc4047ee;
      9668: inst = 32'h8220000;
      9669: inst = 32'h10408000;
      9670: inst = 32'hc4047ef;
      9671: inst = 32'h8220000;
      9672: inst = 32'h10408000;
      9673: inst = 32'hc4047f0;
      9674: inst = 32'h8220000;
      9675: inst = 32'h10408000;
      9676: inst = 32'hc4047f1;
      9677: inst = 32'h8220000;
      9678: inst = 32'h10408000;
      9679: inst = 32'hc4047f2;
      9680: inst = 32'h8220000;
      9681: inst = 32'h10408000;
      9682: inst = 32'hc4047f3;
      9683: inst = 32'h8220000;
      9684: inst = 32'h10408000;
      9685: inst = 32'hc4047f4;
      9686: inst = 32'h8220000;
      9687: inst = 32'h10408000;
      9688: inst = 32'hc4047f5;
      9689: inst = 32'h8220000;
      9690: inst = 32'h10408000;
      9691: inst = 32'hc4047f6;
      9692: inst = 32'h8220000;
      9693: inst = 32'h10408000;
      9694: inst = 32'hc4047f7;
      9695: inst = 32'h8220000;
      9696: inst = 32'h10408000;
      9697: inst = 32'hc4047f8;
      9698: inst = 32'h8220000;
      9699: inst = 32'h10408000;
      9700: inst = 32'hc4047f9;
      9701: inst = 32'h8220000;
      9702: inst = 32'h10408000;
      9703: inst = 32'hc4047fa;
      9704: inst = 32'h8220000;
      9705: inst = 32'h10408000;
      9706: inst = 32'hc4047fb;
      9707: inst = 32'h8220000;
      9708: inst = 32'h10408000;
      9709: inst = 32'hc4047fc;
      9710: inst = 32'h8220000;
      9711: inst = 32'h10408000;
      9712: inst = 32'hc4047fd;
      9713: inst = 32'h8220000;
      9714: inst = 32'h10408000;
      9715: inst = 32'hc4047fe;
      9716: inst = 32'h8220000;
      9717: inst = 32'h10408000;
      9718: inst = 32'hc4047ff;
      9719: inst = 32'h8220000;
      9720: inst = 32'h10408000;
      9721: inst = 32'hc404800;
      9722: inst = 32'h8220000;
      9723: inst = 32'h10408000;
      9724: inst = 32'hc404801;
      9725: inst = 32'h8220000;
      9726: inst = 32'h10408000;
      9727: inst = 32'hc404802;
      9728: inst = 32'h8220000;
      9729: inst = 32'h10408000;
      9730: inst = 32'hc404803;
      9731: inst = 32'h8220000;
      9732: inst = 32'h10408000;
      9733: inst = 32'hc40483c;
      9734: inst = 32'h8220000;
      9735: inst = 32'h10408000;
      9736: inst = 32'hc40483d;
      9737: inst = 32'h8220000;
      9738: inst = 32'h10408000;
      9739: inst = 32'hc40483e;
      9740: inst = 32'h8220000;
      9741: inst = 32'h10408000;
      9742: inst = 32'hc40483f;
      9743: inst = 32'h8220000;
      9744: inst = 32'h10408000;
      9745: inst = 32'hc404840;
      9746: inst = 32'h8220000;
      9747: inst = 32'h10408000;
      9748: inst = 32'hc404841;
      9749: inst = 32'h8220000;
      9750: inst = 32'h10408000;
      9751: inst = 32'hc404842;
      9752: inst = 32'h8220000;
      9753: inst = 32'h10408000;
      9754: inst = 32'hc404843;
      9755: inst = 32'h8220000;
      9756: inst = 32'h10408000;
      9757: inst = 32'hc404844;
      9758: inst = 32'h8220000;
      9759: inst = 32'h10408000;
      9760: inst = 32'hc404845;
      9761: inst = 32'h8220000;
      9762: inst = 32'h10408000;
      9763: inst = 32'hc404846;
      9764: inst = 32'h8220000;
      9765: inst = 32'h10408000;
      9766: inst = 32'hc404847;
      9767: inst = 32'h8220000;
      9768: inst = 32'h10408000;
      9769: inst = 32'hc404848;
      9770: inst = 32'h8220000;
      9771: inst = 32'h10408000;
      9772: inst = 32'hc404849;
      9773: inst = 32'h8220000;
      9774: inst = 32'h10408000;
      9775: inst = 32'hc40484a;
      9776: inst = 32'h8220000;
      9777: inst = 32'h10408000;
      9778: inst = 32'hc40484b;
      9779: inst = 32'h8220000;
      9780: inst = 32'h10408000;
      9781: inst = 32'hc40484c;
      9782: inst = 32'h8220000;
      9783: inst = 32'h10408000;
      9784: inst = 32'hc40484d;
      9785: inst = 32'h8220000;
      9786: inst = 32'h10408000;
      9787: inst = 32'hc40484e;
      9788: inst = 32'h8220000;
      9789: inst = 32'h10408000;
      9790: inst = 32'hc40484f;
      9791: inst = 32'h8220000;
      9792: inst = 32'h10408000;
      9793: inst = 32'hc404850;
      9794: inst = 32'h8220000;
      9795: inst = 32'h10408000;
      9796: inst = 32'hc404851;
      9797: inst = 32'h8220000;
      9798: inst = 32'h10408000;
      9799: inst = 32'hc404852;
      9800: inst = 32'h8220000;
      9801: inst = 32'h10408000;
      9802: inst = 32'hc404853;
      9803: inst = 32'h8220000;
      9804: inst = 32'h10408000;
      9805: inst = 32'hc404854;
      9806: inst = 32'h8220000;
      9807: inst = 32'h10408000;
      9808: inst = 32'hc404855;
      9809: inst = 32'h8220000;
      9810: inst = 32'h10408000;
      9811: inst = 32'hc404856;
      9812: inst = 32'h8220000;
      9813: inst = 32'h10408000;
      9814: inst = 32'hc404857;
      9815: inst = 32'h8220000;
      9816: inst = 32'h10408000;
      9817: inst = 32'hc404858;
      9818: inst = 32'h8220000;
      9819: inst = 32'h10408000;
      9820: inst = 32'hc404859;
      9821: inst = 32'h8220000;
      9822: inst = 32'h10408000;
      9823: inst = 32'hc40485a;
      9824: inst = 32'h8220000;
      9825: inst = 32'h10408000;
      9826: inst = 32'hc40485b;
      9827: inst = 32'h8220000;
      9828: inst = 32'h10408000;
      9829: inst = 32'hc40485c;
      9830: inst = 32'h8220000;
      9831: inst = 32'h10408000;
      9832: inst = 32'hc40485d;
      9833: inst = 32'h8220000;
      9834: inst = 32'h10408000;
      9835: inst = 32'hc40485e;
      9836: inst = 32'h8220000;
      9837: inst = 32'h10408000;
      9838: inst = 32'hc40485f;
      9839: inst = 32'h8220000;
      9840: inst = 32'h10408000;
      9841: inst = 32'hc404860;
      9842: inst = 32'h8220000;
      9843: inst = 32'h10408000;
      9844: inst = 32'hc404861;
      9845: inst = 32'h8220000;
      9846: inst = 32'h10408000;
      9847: inst = 32'hc404862;
      9848: inst = 32'h8220000;
      9849: inst = 32'h10408000;
      9850: inst = 32'hc404863;
      9851: inst = 32'h8220000;
      9852: inst = 32'h10408000;
      9853: inst = 32'hc40489c;
      9854: inst = 32'h8220000;
      9855: inst = 32'h10408000;
      9856: inst = 32'hc40489d;
      9857: inst = 32'h8220000;
      9858: inst = 32'h10408000;
      9859: inst = 32'hc40489e;
      9860: inst = 32'h8220000;
      9861: inst = 32'h10408000;
      9862: inst = 32'hc40489f;
      9863: inst = 32'h8220000;
      9864: inst = 32'h10408000;
      9865: inst = 32'hc4048a0;
      9866: inst = 32'h8220000;
      9867: inst = 32'h10408000;
      9868: inst = 32'hc4048a1;
      9869: inst = 32'h8220000;
      9870: inst = 32'h10408000;
      9871: inst = 32'hc4048a2;
      9872: inst = 32'h8220000;
      9873: inst = 32'h10408000;
      9874: inst = 32'hc4048a3;
      9875: inst = 32'h8220000;
      9876: inst = 32'h10408000;
      9877: inst = 32'hc4048a4;
      9878: inst = 32'h8220000;
      9879: inst = 32'h10408000;
      9880: inst = 32'hc4048a5;
      9881: inst = 32'h8220000;
      9882: inst = 32'h10408000;
      9883: inst = 32'hc4048a6;
      9884: inst = 32'h8220000;
      9885: inst = 32'h10408000;
      9886: inst = 32'hc4048a7;
      9887: inst = 32'h8220000;
      9888: inst = 32'h10408000;
      9889: inst = 32'hc4048a8;
      9890: inst = 32'h8220000;
      9891: inst = 32'h10408000;
      9892: inst = 32'hc4048a9;
      9893: inst = 32'h8220000;
      9894: inst = 32'h10408000;
      9895: inst = 32'hc4048aa;
      9896: inst = 32'h8220000;
      9897: inst = 32'h10408000;
      9898: inst = 32'hc4048ab;
      9899: inst = 32'h8220000;
      9900: inst = 32'h10408000;
      9901: inst = 32'hc4048ac;
      9902: inst = 32'h8220000;
      9903: inst = 32'h10408000;
      9904: inst = 32'hc4048ad;
      9905: inst = 32'h8220000;
      9906: inst = 32'h10408000;
      9907: inst = 32'hc4048ae;
      9908: inst = 32'h8220000;
      9909: inst = 32'h10408000;
      9910: inst = 32'hc4048af;
      9911: inst = 32'h8220000;
      9912: inst = 32'h10408000;
      9913: inst = 32'hc4048b0;
      9914: inst = 32'h8220000;
      9915: inst = 32'h10408000;
      9916: inst = 32'hc4048b1;
      9917: inst = 32'h8220000;
      9918: inst = 32'h10408000;
      9919: inst = 32'hc4048b2;
      9920: inst = 32'h8220000;
      9921: inst = 32'h10408000;
      9922: inst = 32'hc4048b3;
      9923: inst = 32'h8220000;
      9924: inst = 32'h10408000;
      9925: inst = 32'hc4048b4;
      9926: inst = 32'h8220000;
      9927: inst = 32'h10408000;
      9928: inst = 32'hc4048b5;
      9929: inst = 32'h8220000;
      9930: inst = 32'h10408000;
      9931: inst = 32'hc4048b6;
      9932: inst = 32'h8220000;
      9933: inst = 32'h10408000;
      9934: inst = 32'hc4048b7;
      9935: inst = 32'h8220000;
      9936: inst = 32'h10408000;
      9937: inst = 32'hc4048b8;
      9938: inst = 32'h8220000;
      9939: inst = 32'h10408000;
      9940: inst = 32'hc4048b9;
      9941: inst = 32'h8220000;
      9942: inst = 32'h10408000;
      9943: inst = 32'hc4048ba;
      9944: inst = 32'h8220000;
      9945: inst = 32'h10408000;
      9946: inst = 32'hc4048bb;
      9947: inst = 32'h8220000;
      9948: inst = 32'h10408000;
      9949: inst = 32'hc4048bc;
      9950: inst = 32'h8220000;
      9951: inst = 32'h10408000;
      9952: inst = 32'hc4048bd;
      9953: inst = 32'h8220000;
      9954: inst = 32'h10408000;
      9955: inst = 32'hc4048be;
      9956: inst = 32'h8220000;
      9957: inst = 32'h10408000;
      9958: inst = 32'hc4048bf;
      9959: inst = 32'h8220000;
      9960: inst = 32'h10408000;
      9961: inst = 32'hc4048c0;
      9962: inst = 32'h8220000;
      9963: inst = 32'h10408000;
      9964: inst = 32'hc4048c1;
      9965: inst = 32'h8220000;
      9966: inst = 32'h10408000;
      9967: inst = 32'hc4048c2;
      9968: inst = 32'h8220000;
      9969: inst = 32'h10408000;
      9970: inst = 32'hc4048c3;
      9971: inst = 32'h8220000;
      9972: inst = 32'h10408000;
      9973: inst = 32'hc4048fc;
      9974: inst = 32'h8220000;
      9975: inst = 32'h10408000;
      9976: inst = 32'hc4048fd;
      9977: inst = 32'h8220000;
      9978: inst = 32'h10408000;
      9979: inst = 32'hc4048fe;
      9980: inst = 32'h8220000;
      9981: inst = 32'h10408000;
      9982: inst = 32'hc4048ff;
      9983: inst = 32'h8220000;
      9984: inst = 32'h10408000;
      9985: inst = 32'hc404900;
      9986: inst = 32'h8220000;
      9987: inst = 32'h10408000;
      9988: inst = 32'hc404901;
      9989: inst = 32'h8220000;
      9990: inst = 32'h10408000;
      9991: inst = 32'hc404902;
      9992: inst = 32'h8220000;
      9993: inst = 32'h10408000;
      9994: inst = 32'hc404903;
      9995: inst = 32'h8220000;
      9996: inst = 32'h10408000;
      9997: inst = 32'hc404904;
      9998: inst = 32'h8220000;
      9999: inst = 32'h10408000;
      10000: inst = 32'hc404905;
      10001: inst = 32'h8220000;
      10002: inst = 32'h10408000;
      10003: inst = 32'hc404906;
      10004: inst = 32'h8220000;
      10005: inst = 32'h10408000;
      10006: inst = 32'hc404907;
      10007: inst = 32'h8220000;
      10008: inst = 32'h10408000;
      10009: inst = 32'hc404908;
      10010: inst = 32'h8220000;
      10011: inst = 32'h10408000;
      10012: inst = 32'hc404909;
      10013: inst = 32'h8220000;
      10014: inst = 32'h10408000;
      10015: inst = 32'hc40490a;
      10016: inst = 32'h8220000;
      10017: inst = 32'h10408000;
      10018: inst = 32'hc40490b;
      10019: inst = 32'h8220000;
      10020: inst = 32'h10408000;
      10021: inst = 32'hc40490c;
      10022: inst = 32'h8220000;
      10023: inst = 32'h10408000;
      10024: inst = 32'hc40490d;
      10025: inst = 32'h8220000;
      10026: inst = 32'h10408000;
      10027: inst = 32'hc40490e;
      10028: inst = 32'h8220000;
      10029: inst = 32'h10408000;
      10030: inst = 32'hc40490f;
      10031: inst = 32'h8220000;
      10032: inst = 32'h10408000;
      10033: inst = 32'hc404910;
      10034: inst = 32'h8220000;
      10035: inst = 32'h10408000;
      10036: inst = 32'hc404911;
      10037: inst = 32'h8220000;
      10038: inst = 32'h10408000;
      10039: inst = 32'hc404912;
      10040: inst = 32'h8220000;
      10041: inst = 32'h10408000;
      10042: inst = 32'hc404913;
      10043: inst = 32'h8220000;
      10044: inst = 32'h10408000;
      10045: inst = 32'hc404914;
      10046: inst = 32'h8220000;
      10047: inst = 32'h10408000;
      10048: inst = 32'hc404915;
      10049: inst = 32'h8220000;
      10050: inst = 32'h10408000;
      10051: inst = 32'hc404916;
      10052: inst = 32'h8220000;
      10053: inst = 32'h10408000;
      10054: inst = 32'hc404917;
      10055: inst = 32'h8220000;
      10056: inst = 32'h10408000;
      10057: inst = 32'hc404918;
      10058: inst = 32'h8220000;
      10059: inst = 32'h10408000;
      10060: inst = 32'hc404919;
      10061: inst = 32'h8220000;
      10062: inst = 32'h10408000;
      10063: inst = 32'hc40491a;
      10064: inst = 32'h8220000;
      10065: inst = 32'h10408000;
      10066: inst = 32'hc40491b;
      10067: inst = 32'h8220000;
      10068: inst = 32'h10408000;
      10069: inst = 32'hc40491c;
      10070: inst = 32'h8220000;
      10071: inst = 32'h10408000;
      10072: inst = 32'hc40491d;
      10073: inst = 32'h8220000;
      10074: inst = 32'h10408000;
      10075: inst = 32'hc40491e;
      10076: inst = 32'h8220000;
      10077: inst = 32'h10408000;
      10078: inst = 32'hc40491f;
      10079: inst = 32'h8220000;
      10080: inst = 32'h10408000;
      10081: inst = 32'hc404920;
      10082: inst = 32'h8220000;
      10083: inst = 32'h10408000;
      10084: inst = 32'hc404921;
      10085: inst = 32'h8220000;
      10086: inst = 32'h10408000;
      10087: inst = 32'hc404922;
      10088: inst = 32'h8220000;
      10089: inst = 32'h10408000;
      10090: inst = 32'hc404923;
      10091: inst = 32'h8220000;
      10092: inst = 32'h10408000;
      10093: inst = 32'hc40495c;
      10094: inst = 32'h8220000;
      10095: inst = 32'h10408000;
      10096: inst = 32'hc40495d;
      10097: inst = 32'h8220000;
      10098: inst = 32'h10408000;
      10099: inst = 32'hc40495e;
      10100: inst = 32'h8220000;
      10101: inst = 32'h10408000;
      10102: inst = 32'hc40495f;
      10103: inst = 32'h8220000;
      10104: inst = 32'h10408000;
      10105: inst = 32'hc404960;
      10106: inst = 32'h8220000;
      10107: inst = 32'h10408000;
      10108: inst = 32'hc404961;
      10109: inst = 32'h8220000;
      10110: inst = 32'h10408000;
      10111: inst = 32'hc404962;
      10112: inst = 32'h8220000;
      10113: inst = 32'h10408000;
      10114: inst = 32'hc404963;
      10115: inst = 32'h8220000;
      10116: inst = 32'h10408000;
      10117: inst = 32'hc404964;
      10118: inst = 32'h8220000;
      10119: inst = 32'h10408000;
      10120: inst = 32'hc404965;
      10121: inst = 32'h8220000;
      10122: inst = 32'h10408000;
      10123: inst = 32'hc404966;
      10124: inst = 32'h8220000;
      10125: inst = 32'h10408000;
      10126: inst = 32'hc404967;
      10127: inst = 32'h8220000;
      10128: inst = 32'h10408000;
      10129: inst = 32'hc404968;
      10130: inst = 32'h8220000;
      10131: inst = 32'h10408000;
      10132: inst = 32'hc404969;
      10133: inst = 32'h8220000;
      10134: inst = 32'h10408000;
      10135: inst = 32'hc40496a;
      10136: inst = 32'h8220000;
      10137: inst = 32'h10408000;
      10138: inst = 32'hc40496b;
      10139: inst = 32'h8220000;
      10140: inst = 32'h10408000;
      10141: inst = 32'hc40496c;
      10142: inst = 32'h8220000;
      10143: inst = 32'h10408000;
      10144: inst = 32'hc40496d;
      10145: inst = 32'h8220000;
      10146: inst = 32'h10408000;
      10147: inst = 32'hc40496e;
      10148: inst = 32'h8220000;
      10149: inst = 32'h10408000;
      10150: inst = 32'hc40496f;
      10151: inst = 32'h8220000;
      10152: inst = 32'h10408000;
      10153: inst = 32'hc404970;
      10154: inst = 32'h8220000;
      10155: inst = 32'h10408000;
      10156: inst = 32'hc404971;
      10157: inst = 32'h8220000;
      10158: inst = 32'h10408000;
      10159: inst = 32'hc404972;
      10160: inst = 32'h8220000;
      10161: inst = 32'h10408000;
      10162: inst = 32'hc404973;
      10163: inst = 32'h8220000;
      10164: inst = 32'h10408000;
      10165: inst = 32'hc404974;
      10166: inst = 32'h8220000;
      10167: inst = 32'h10408000;
      10168: inst = 32'hc404975;
      10169: inst = 32'h8220000;
      10170: inst = 32'h10408000;
      10171: inst = 32'hc404976;
      10172: inst = 32'h8220000;
      10173: inst = 32'h10408000;
      10174: inst = 32'hc404977;
      10175: inst = 32'h8220000;
      10176: inst = 32'h10408000;
      10177: inst = 32'hc404978;
      10178: inst = 32'h8220000;
      10179: inst = 32'h10408000;
      10180: inst = 32'hc404979;
      10181: inst = 32'h8220000;
      10182: inst = 32'h10408000;
      10183: inst = 32'hc40497a;
      10184: inst = 32'h8220000;
      10185: inst = 32'h10408000;
      10186: inst = 32'hc40497b;
      10187: inst = 32'h8220000;
      10188: inst = 32'h10408000;
      10189: inst = 32'hc40497c;
      10190: inst = 32'h8220000;
      10191: inst = 32'h10408000;
      10192: inst = 32'hc40497d;
      10193: inst = 32'h8220000;
      10194: inst = 32'h10408000;
      10195: inst = 32'hc40497e;
      10196: inst = 32'h8220000;
      10197: inst = 32'h10408000;
      10198: inst = 32'hc40497f;
      10199: inst = 32'h8220000;
      10200: inst = 32'h10408000;
      10201: inst = 32'hc404980;
      10202: inst = 32'h8220000;
      10203: inst = 32'h10408000;
      10204: inst = 32'hc404981;
      10205: inst = 32'h8220000;
      10206: inst = 32'h10408000;
      10207: inst = 32'hc404982;
      10208: inst = 32'h8220000;
      10209: inst = 32'h10408000;
      10210: inst = 32'hc404983;
      10211: inst = 32'h8220000;
      10212: inst = 32'h10408000;
      10213: inst = 32'hc404992;
      10214: inst = 32'h8220000;
      10215: inst = 32'h10408000;
      10216: inst = 32'hc4049bc;
      10217: inst = 32'h8220000;
      10218: inst = 32'h10408000;
      10219: inst = 32'hc4049bd;
      10220: inst = 32'h8220000;
      10221: inst = 32'h10408000;
      10222: inst = 32'hc4049be;
      10223: inst = 32'h8220000;
      10224: inst = 32'h10408000;
      10225: inst = 32'hc4049bf;
      10226: inst = 32'h8220000;
      10227: inst = 32'h10408000;
      10228: inst = 32'hc4049c0;
      10229: inst = 32'h8220000;
      10230: inst = 32'h10408000;
      10231: inst = 32'hc4049c1;
      10232: inst = 32'h8220000;
      10233: inst = 32'h10408000;
      10234: inst = 32'hc4049c2;
      10235: inst = 32'h8220000;
      10236: inst = 32'h10408000;
      10237: inst = 32'hc4049c3;
      10238: inst = 32'h8220000;
      10239: inst = 32'h10408000;
      10240: inst = 32'hc4049c4;
      10241: inst = 32'h8220000;
      10242: inst = 32'h10408000;
      10243: inst = 32'hc4049c5;
      10244: inst = 32'h8220000;
      10245: inst = 32'h10408000;
      10246: inst = 32'hc4049c6;
      10247: inst = 32'h8220000;
      10248: inst = 32'h10408000;
      10249: inst = 32'hc4049c7;
      10250: inst = 32'h8220000;
      10251: inst = 32'h10408000;
      10252: inst = 32'hc4049c8;
      10253: inst = 32'h8220000;
      10254: inst = 32'h10408000;
      10255: inst = 32'hc4049c9;
      10256: inst = 32'h8220000;
      10257: inst = 32'h10408000;
      10258: inst = 32'hc4049ca;
      10259: inst = 32'h8220000;
      10260: inst = 32'h10408000;
      10261: inst = 32'hc4049cb;
      10262: inst = 32'h8220000;
      10263: inst = 32'h10408000;
      10264: inst = 32'hc4049cc;
      10265: inst = 32'h8220000;
      10266: inst = 32'h10408000;
      10267: inst = 32'hc4049cd;
      10268: inst = 32'h8220000;
      10269: inst = 32'h10408000;
      10270: inst = 32'hc4049ce;
      10271: inst = 32'h8220000;
      10272: inst = 32'h10408000;
      10273: inst = 32'hc4049cf;
      10274: inst = 32'h8220000;
      10275: inst = 32'h10408000;
      10276: inst = 32'hc4049d0;
      10277: inst = 32'h8220000;
      10278: inst = 32'h10408000;
      10279: inst = 32'hc4049d1;
      10280: inst = 32'h8220000;
      10281: inst = 32'h10408000;
      10282: inst = 32'hc4049d2;
      10283: inst = 32'h8220000;
      10284: inst = 32'h10408000;
      10285: inst = 32'hc4049d3;
      10286: inst = 32'h8220000;
      10287: inst = 32'h10408000;
      10288: inst = 32'hc4049d4;
      10289: inst = 32'h8220000;
      10290: inst = 32'h10408000;
      10291: inst = 32'hc4049d5;
      10292: inst = 32'h8220000;
      10293: inst = 32'h10408000;
      10294: inst = 32'hc4049d6;
      10295: inst = 32'h8220000;
      10296: inst = 32'h10408000;
      10297: inst = 32'hc4049d7;
      10298: inst = 32'h8220000;
      10299: inst = 32'h10408000;
      10300: inst = 32'hc4049d8;
      10301: inst = 32'h8220000;
      10302: inst = 32'h10408000;
      10303: inst = 32'hc4049d9;
      10304: inst = 32'h8220000;
      10305: inst = 32'h10408000;
      10306: inst = 32'hc4049da;
      10307: inst = 32'h8220000;
      10308: inst = 32'h10408000;
      10309: inst = 32'hc4049db;
      10310: inst = 32'h8220000;
      10311: inst = 32'h10408000;
      10312: inst = 32'hc4049dc;
      10313: inst = 32'h8220000;
      10314: inst = 32'h10408000;
      10315: inst = 32'hc4049dd;
      10316: inst = 32'h8220000;
      10317: inst = 32'h10408000;
      10318: inst = 32'hc4049de;
      10319: inst = 32'h8220000;
      10320: inst = 32'h10408000;
      10321: inst = 32'hc4049df;
      10322: inst = 32'h8220000;
      10323: inst = 32'h10408000;
      10324: inst = 32'hc4049e0;
      10325: inst = 32'h8220000;
      10326: inst = 32'h10408000;
      10327: inst = 32'hc4049e1;
      10328: inst = 32'h8220000;
      10329: inst = 32'h10408000;
      10330: inst = 32'hc4049e2;
      10331: inst = 32'h8220000;
      10332: inst = 32'h10408000;
      10333: inst = 32'hc4049e3;
      10334: inst = 32'h8220000;
      10335: inst = 32'h10408000;
      10336: inst = 32'hc4049f2;
      10337: inst = 32'h8220000;
      10338: inst = 32'h10408000;
      10339: inst = 32'hc404a1c;
      10340: inst = 32'h8220000;
      10341: inst = 32'h10408000;
      10342: inst = 32'hc404a1d;
      10343: inst = 32'h8220000;
      10344: inst = 32'h10408000;
      10345: inst = 32'hc404a1e;
      10346: inst = 32'h8220000;
      10347: inst = 32'h10408000;
      10348: inst = 32'hc404a1f;
      10349: inst = 32'h8220000;
      10350: inst = 32'h10408000;
      10351: inst = 32'hc404a20;
      10352: inst = 32'h8220000;
      10353: inst = 32'h10408000;
      10354: inst = 32'hc404a21;
      10355: inst = 32'h8220000;
      10356: inst = 32'h10408000;
      10357: inst = 32'hc404a22;
      10358: inst = 32'h8220000;
      10359: inst = 32'h10408000;
      10360: inst = 32'hc404a23;
      10361: inst = 32'h8220000;
      10362: inst = 32'h10408000;
      10363: inst = 32'hc404a24;
      10364: inst = 32'h8220000;
      10365: inst = 32'h10408000;
      10366: inst = 32'hc404a25;
      10367: inst = 32'h8220000;
      10368: inst = 32'h10408000;
      10369: inst = 32'hc404a26;
      10370: inst = 32'h8220000;
      10371: inst = 32'h10408000;
      10372: inst = 32'hc404a27;
      10373: inst = 32'h8220000;
      10374: inst = 32'h10408000;
      10375: inst = 32'hc404a28;
      10376: inst = 32'h8220000;
      10377: inst = 32'h10408000;
      10378: inst = 32'hc404a29;
      10379: inst = 32'h8220000;
      10380: inst = 32'h10408000;
      10381: inst = 32'hc404a2a;
      10382: inst = 32'h8220000;
      10383: inst = 32'h10408000;
      10384: inst = 32'hc404a2b;
      10385: inst = 32'h8220000;
      10386: inst = 32'h10408000;
      10387: inst = 32'hc404a2c;
      10388: inst = 32'h8220000;
      10389: inst = 32'h10408000;
      10390: inst = 32'hc404a2d;
      10391: inst = 32'h8220000;
      10392: inst = 32'h10408000;
      10393: inst = 32'hc404a2e;
      10394: inst = 32'h8220000;
      10395: inst = 32'h10408000;
      10396: inst = 32'hc404a2f;
      10397: inst = 32'h8220000;
      10398: inst = 32'h10408000;
      10399: inst = 32'hc404a30;
      10400: inst = 32'h8220000;
      10401: inst = 32'h10408000;
      10402: inst = 32'hc404a31;
      10403: inst = 32'h8220000;
      10404: inst = 32'h10408000;
      10405: inst = 32'hc404a32;
      10406: inst = 32'h8220000;
      10407: inst = 32'h10408000;
      10408: inst = 32'hc404a33;
      10409: inst = 32'h8220000;
      10410: inst = 32'h10408000;
      10411: inst = 32'hc404a34;
      10412: inst = 32'h8220000;
      10413: inst = 32'h10408000;
      10414: inst = 32'hc404a35;
      10415: inst = 32'h8220000;
      10416: inst = 32'h10408000;
      10417: inst = 32'hc404a36;
      10418: inst = 32'h8220000;
      10419: inst = 32'h10408000;
      10420: inst = 32'hc404a37;
      10421: inst = 32'h8220000;
      10422: inst = 32'h10408000;
      10423: inst = 32'hc404a38;
      10424: inst = 32'h8220000;
      10425: inst = 32'h10408000;
      10426: inst = 32'hc404a39;
      10427: inst = 32'h8220000;
      10428: inst = 32'h10408000;
      10429: inst = 32'hc404a3a;
      10430: inst = 32'h8220000;
      10431: inst = 32'h10408000;
      10432: inst = 32'hc404a3b;
      10433: inst = 32'h8220000;
      10434: inst = 32'h10408000;
      10435: inst = 32'hc404a3c;
      10436: inst = 32'h8220000;
      10437: inst = 32'h10408000;
      10438: inst = 32'hc404a3d;
      10439: inst = 32'h8220000;
      10440: inst = 32'h10408000;
      10441: inst = 32'hc404a3e;
      10442: inst = 32'h8220000;
      10443: inst = 32'h10408000;
      10444: inst = 32'hc404a3f;
      10445: inst = 32'h8220000;
      10446: inst = 32'h10408000;
      10447: inst = 32'hc404a40;
      10448: inst = 32'h8220000;
      10449: inst = 32'h10408000;
      10450: inst = 32'hc404a41;
      10451: inst = 32'h8220000;
      10452: inst = 32'h10408000;
      10453: inst = 32'hc404a42;
      10454: inst = 32'h8220000;
      10455: inst = 32'h10408000;
      10456: inst = 32'hc404a43;
      10457: inst = 32'h8220000;
      10458: inst = 32'h10408000;
      10459: inst = 32'hc404a52;
      10460: inst = 32'h8220000;
      10461: inst = 32'h10408000;
      10462: inst = 32'hc404a7c;
      10463: inst = 32'h8220000;
      10464: inst = 32'h10408000;
      10465: inst = 32'hc404a7d;
      10466: inst = 32'h8220000;
      10467: inst = 32'h10408000;
      10468: inst = 32'hc404a7e;
      10469: inst = 32'h8220000;
      10470: inst = 32'h10408000;
      10471: inst = 32'hc404a7f;
      10472: inst = 32'h8220000;
      10473: inst = 32'h10408000;
      10474: inst = 32'hc404a80;
      10475: inst = 32'h8220000;
      10476: inst = 32'h10408000;
      10477: inst = 32'hc404a81;
      10478: inst = 32'h8220000;
      10479: inst = 32'h10408000;
      10480: inst = 32'hc404a82;
      10481: inst = 32'h8220000;
      10482: inst = 32'h10408000;
      10483: inst = 32'hc404a83;
      10484: inst = 32'h8220000;
      10485: inst = 32'h10408000;
      10486: inst = 32'hc404a84;
      10487: inst = 32'h8220000;
      10488: inst = 32'h10408000;
      10489: inst = 32'hc404a85;
      10490: inst = 32'h8220000;
      10491: inst = 32'h10408000;
      10492: inst = 32'hc404a86;
      10493: inst = 32'h8220000;
      10494: inst = 32'h10408000;
      10495: inst = 32'hc404a87;
      10496: inst = 32'h8220000;
      10497: inst = 32'h10408000;
      10498: inst = 32'hc404a88;
      10499: inst = 32'h8220000;
      10500: inst = 32'h10408000;
      10501: inst = 32'hc404a89;
      10502: inst = 32'h8220000;
      10503: inst = 32'h10408000;
      10504: inst = 32'hc404a8a;
      10505: inst = 32'h8220000;
      10506: inst = 32'h10408000;
      10507: inst = 32'hc404a8b;
      10508: inst = 32'h8220000;
      10509: inst = 32'h10408000;
      10510: inst = 32'hc404a8c;
      10511: inst = 32'h8220000;
      10512: inst = 32'h10408000;
      10513: inst = 32'hc404a8d;
      10514: inst = 32'h8220000;
      10515: inst = 32'h10408000;
      10516: inst = 32'hc404a8e;
      10517: inst = 32'h8220000;
      10518: inst = 32'h10408000;
      10519: inst = 32'hc404a8f;
      10520: inst = 32'h8220000;
      10521: inst = 32'h10408000;
      10522: inst = 32'hc404a90;
      10523: inst = 32'h8220000;
      10524: inst = 32'h10408000;
      10525: inst = 32'hc404a91;
      10526: inst = 32'h8220000;
      10527: inst = 32'h10408000;
      10528: inst = 32'hc404a92;
      10529: inst = 32'h8220000;
      10530: inst = 32'h10408000;
      10531: inst = 32'hc404a93;
      10532: inst = 32'h8220000;
      10533: inst = 32'h10408000;
      10534: inst = 32'hc404a94;
      10535: inst = 32'h8220000;
      10536: inst = 32'h10408000;
      10537: inst = 32'hc404a95;
      10538: inst = 32'h8220000;
      10539: inst = 32'h10408000;
      10540: inst = 32'hc404a96;
      10541: inst = 32'h8220000;
      10542: inst = 32'h10408000;
      10543: inst = 32'hc404a97;
      10544: inst = 32'h8220000;
      10545: inst = 32'h10408000;
      10546: inst = 32'hc404a98;
      10547: inst = 32'h8220000;
      10548: inst = 32'h10408000;
      10549: inst = 32'hc404a99;
      10550: inst = 32'h8220000;
      10551: inst = 32'h10408000;
      10552: inst = 32'hc404a9a;
      10553: inst = 32'h8220000;
      10554: inst = 32'h10408000;
      10555: inst = 32'hc404a9b;
      10556: inst = 32'h8220000;
      10557: inst = 32'h10408000;
      10558: inst = 32'hc404a9c;
      10559: inst = 32'h8220000;
      10560: inst = 32'h10408000;
      10561: inst = 32'hc404a9d;
      10562: inst = 32'h8220000;
      10563: inst = 32'h10408000;
      10564: inst = 32'hc404a9e;
      10565: inst = 32'h8220000;
      10566: inst = 32'h10408000;
      10567: inst = 32'hc404a9f;
      10568: inst = 32'h8220000;
      10569: inst = 32'h10408000;
      10570: inst = 32'hc404aa0;
      10571: inst = 32'h8220000;
      10572: inst = 32'h10408000;
      10573: inst = 32'hc404aa1;
      10574: inst = 32'h8220000;
      10575: inst = 32'h10408000;
      10576: inst = 32'hc404aa2;
      10577: inst = 32'h8220000;
      10578: inst = 32'h10408000;
      10579: inst = 32'hc404aa3;
      10580: inst = 32'h8220000;
      10581: inst = 32'h10408000;
      10582: inst = 32'hc404ab4;
      10583: inst = 32'h8220000;
      10584: inst = 32'h10408000;
      10585: inst = 32'hc404adc;
      10586: inst = 32'h8220000;
      10587: inst = 32'h10408000;
      10588: inst = 32'hc404add;
      10589: inst = 32'h8220000;
      10590: inst = 32'h10408000;
      10591: inst = 32'hc404ade;
      10592: inst = 32'h8220000;
      10593: inst = 32'h10408000;
      10594: inst = 32'hc404adf;
      10595: inst = 32'h8220000;
      10596: inst = 32'h10408000;
      10597: inst = 32'hc404ae0;
      10598: inst = 32'h8220000;
      10599: inst = 32'h10408000;
      10600: inst = 32'hc404ae1;
      10601: inst = 32'h8220000;
      10602: inst = 32'h10408000;
      10603: inst = 32'hc404ae2;
      10604: inst = 32'h8220000;
      10605: inst = 32'h10408000;
      10606: inst = 32'hc404ae3;
      10607: inst = 32'h8220000;
      10608: inst = 32'h10408000;
      10609: inst = 32'hc404ae4;
      10610: inst = 32'h8220000;
      10611: inst = 32'h10408000;
      10612: inst = 32'hc404ae5;
      10613: inst = 32'h8220000;
      10614: inst = 32'h10408000;
      10615: inst = 32'hc404ae6;
      10616: inst = 32'h8220000;
      10617: inst = 32'h10408000;
      10618: inst = 32'hc404ae7;
      10619: inst = 32'h8220000;
      10620: inst = 32'h10408000;
      10621: inst = 32'hc404ae8;
      10622: inst = 32'h8220000;
      10623: inst = 32'h10408000;
      10624: inst = 32'hc404ae9;
      10625: inst = 32'h8220000;
      10626: inst = 32'h10408000;
      10627: inst = 32'hc404aea;
      10628: inst = 32'h8220000;
      10629: inst = 32'h10408000;
      10630: inst = 32'hc404aeb;
      10631: inst = 32'h8220000;
      10632: inst = 32'h10408000;
      10633: inst = 32'hc404aec;
      10634: inst = 32'h8220000;
      10635: inst = 32'h10408000;
      10636: inst = 32'hc404aed;
      10637: inst = 32'h8220000;
      10638: inst = 32'h10408000;
      10639: inst = 32'hc404aee;
      10640: inst = 32'h8220000;
      10641: inst = 32'h10408000;
      10642: inst = 32'hc404aef;
      10643: inst = 32'h8220000;
      10644: inst = 32'h10408000;
      10645: inst = 32'hc404af0;
      10646: inst = 32'h8220000;
      10647: inst = 32'h10408000;
      10648: inst = 32'hc404af1;
      10649: inst = 32'h8220000;
      10650: inst = 32'h10408000;
      10651: inst = 32'hc404af2;
      10652: inst = 32'h8220000;
      10653: inst = 32'h10408000;
      10654: inst = 32'hc404af3;
      10655: inst = 32'h8220000;
      10656: inst = 32'h10408000;
      10657: inst = 32'hc404af4;
      10658: inst = 32'h8220000;
      10659: inst = 32'h10408000;
      10660: inst = 32'hc404af5;
      10661: inst = 32'h8220000;
      10662: inst = 32'h10408000;
      10663: inst = 32'hc404af6;
      10664: inst = 32'h8220000;
      10665: inst = 32'h10408000;
      10666: inst = 32'hc404af7;
      10667: inst = 32'h8220000;
      10668: inst = 32'h10408000;
      10669: inst = 32'hc404af8;
      10670: inst = 32'h8220000;
      10671: inst = 32'h10408000;
      10672: inst = 32'hc404af9;
      10673: inst = 32'h8220000;
      10674: inst = 32'h10408000;
      10675: inst = 32'hc404afa;
      10676: inst = 32'h8220000;
      10677: inst = 32'h10408000;
      10678: inst = 32'hc404afb;
      10679: inst = 32'h8220000;
      10680: inst = 32'h10408000;
      10681: inst = 32'hc404afc;
      10682: inst = 32'h8220000;
      10683: inst = 32'h10408000;
      10684: inst = 32'hc404afd;
      10685: inst = 32'h8220000;
      10686: inst = 32'h10408000;
      10687: inst = 32'hc404afe;
      10688: inst = 32'h8220000;
      10689: inst = 32'h10408000;
      10690: inst = 32'hc404aff;
      10691: inst = 32'h8220000;
      10692: inst = 32'h10408000;
      10693: inst = 32'hc404b00;
      10694: inst = 32'h8220000;
      10695: inst = 32'h10408000;
      10696: inst = 32'hc404b01;
      10697: inst = 32'h8220000;
      10698: inst = 32'h10408000;
      10699: inst = 32'hc404b02;
      10700: inst = 32'h8220000;
      10701: inst = 32'h10408000;
      10702: inst = 32'hc404b03;
      10703: inst = 32'h8220000;
      10704: inst = 32'h10408000;
      10705: inst = 32'hc404b14;
      10706: inst = 32'h8220000;
      10707: inst = 32'h10408000;
      10708: inst = 32'hc404b3c;
      10709: inst = 32'h8220000;
      10710: inst = 32'h10408000;
      10711: inst = 32'hc404b3d;
      10712: inst = 32'h8220000;
      10713: inst = 32'h10408000;
      10714: inst = 32'hc404b3e;
      10715: inst = 32'h8220000;
      10716: inst = 32'h10408000;
      10717: inst = 32'hc404b3f;
      10718: inst = 32'h8220000;
      10719: inst = 32'h10408000;
      10720: inst = 32'hc404b40;
      10721: inst = 32'h8220000;
      10722: inst = 32'h10408000;
      10723: inst = 32'hc404b41;
      10724: inst = 32'h8220000;
      10725: inst = 32'h10408000;
      10726: inst = 32'hc404b42;
      10727: inst = 32'h8220000;
      10728: inst = 32'h10408000;
      10729: inst = 32'hc404b43;
      10730: inst = 32'h8220000;
      10731: inst = 32'h10408000;
      10732: inst = 32'hc404b44;
      10733: inst = 32'h8220000;
      10734: inst = 32'h10408000;
      10735: inst = 32'hc404b45;
      10736: inst = 32'h8220000;
      10737: inst = 32'h10408000;
      10738: inst = 32'hc404b46;
      10739: inst = 32'h8220000;
      10740: inst = 32'h10408000;
      10741: inst = 32'hc404b47;
      10742: inst = 32'h8220000;
      10743: inst = 32'h10408000;
      10744: inst = 32'hc404b48;
      10745: inst = 32'h8220000;
      10746: inst = 32'h10408000;
      10747: inst = 32'hc404b49;
      10748: inst = 32'h8220000;
      10749: inst = 32'h10408000;
      10750: inst = 32'hc404b4a;
      10751: inst = 32'h8220000;
      10752: inst = 32'h10408000;
      10753: inst = 32'hc404b4b;
      10754: inst = 32'h8220000;
      10755: inst = 32'h10408000;
      10756: inst = 32'hc404b4c;
      10757: inst = 32'h8220000;
      10758: inst = 32'h10408000;
      10759: inst = 32'hc404b4d;
      10760: inst = 32'h8220000;
      10761: inst = 32'h10408000;
      10762: inst = 32'hc404b4e;
      10763: inst = 32'h8220000;
      10764: inst = 32'h10408000;
      10765: inst = 32'hc404b4f;
      10766: inst = 32'h8220000;
      10767: inst = 32'h10408000;
      10768: inst = 32'hc404b50;
      10769: inst = 32'h8220000;
      10770: inst = 32'h10408000;
      10771: inst = 32'hc404b51;
      10772: inst = 32'h8220000;
      10773: inst = 32'h10408000;
      10774: inst = 32'hc404b52;
      10775: inst = 32'h8220000;
      10776: inst = 32'h10408000;
      10777: inst = 32'hc404b53;
      10778: inst = 32'h8220000;
      10779: inst = 32'h10408000;
      10780: inst = 32'hc404b54;
      10781: inst = 32'h8220000;
      10782: inst = 32'h10408000;
      10783: inst = 32'hc404b55;
      10784: inst = 32'h8220000;
      10785: inst = 32'h10408000;
      10786: inst = 32'hc404b56;
      10787: inst = 32'h8220000;
      10788: inst = 32'h10408000;
      10789: inst = 32'hc404b57;
      10790: inst = 32'h8220000;
      10791: inst = 32'h10408000;
      10792: inst = 32'hc404b58;
      10793: inst = 32'h8220000;
      10794: inst = 32'h10408000;
      10795: inst = 32'hc404b59;
      10796: inst = 32'h8220000;
      10797: inst = 32'h10408000;
      10798: inst = 32'hc404b5a;
      10799: inst = 32'h8220000;
      10800: inst = 32'h10408000;
      10801: inst = 32'hc404b5b;
      10802: inst = 32'h8220000;
      10803: inst = 32'h10408000;
      10804: inst = 32'hc404b5c;
      10805: inst = 32'h8220000;
      10806: inst = 32'h10408000;
      10807: inst = 32'hc404b5d;
      10808: inst = 32'h8220000;
      10809: inst = 32'h10408000;
      10810: inst = 32'hc404b5e;
      10811: inst = 32'h8220000;
      10812: inst = 32'h10408000;
      10813: inst = 32'hc404b5f;
      10814: inst = 32'h8220000;
      10815: inst = 32'h10408000;
      10816: inst = 32'hc404b60;
      10817: inst = 32'h8220000;
      10818: inst = 32'h10408000;
      10819: inst = 32'hc404b61;
      10820: inst = 32'h8220000;
      10821: inst = 32'h10408000;
      10822: inst = 32'hc404b62;
      10823: inst = 32'h8220000;
      10824: inst = 32'h10408000;
      10825: inst = 32'hc404b63;
      10826: inst = 32'h8220000;
      10827: inst = 32'h10408000;
      10828: inst = 32'hc404b9c;
      10829: inst = 32'h8220000;
      10830: inst = 32'h10408000;
      10831: inst = 32'hc404b9d;
      10832: inst = 32'h8220000;
      10833: inst = 32'h10408000;
      10834: inst = 32'hc404b9e;
      10835: inst = 32'h8220000;
      10836: inst = 32'h10408000;
      10837: inst = 32'hc404b9f;
      10838: inst = 32'h8220000;
      10839: inst = 32'h10408000;
      10840: inst = 32'hc404ba0;
      10841: inst = 32'h8220000;
      10842: inst = 32'h10408000;
      10843: inst = 32'hc404ba1;
      10844: inst = 32'h8220000;
      10845: inst = 32'h10408000;
      10846: inst = 32'hc404ba2;
      10847: inst = 32'h8220000;
      10848: inst = 32'h10408000;
      10849: inst = 32'hc404ba3;
      10850: inst = 32'h8220000;
      10851: inst = 32'h10408000;
      10852: inst = 32'hc404ba4;
      10853: inst = 32'h8220000;
      10854: inst = 32'h10408000;
      10855: inst = 32'hc404ba5;
      10856: inst = 32'h8220000;
      10857: inst = 32'h10408000;
      10858: inst = 32'hc404ba6;
      10859: inst = 32'h8220000;
      10860: inst = 32'h10408000;
      10861: inst = 32'hc404ba7;
      10862: inst = 32'h8220000;
      10863: inst = 32'h10408000;
      10864: inst = 32'hc404ba8;
      10865: inst = 32'h8220000;
      10866: inst = 32'h10408000;
      10867: inst = 32'hc404ba9;
      10868: inst = 32'h8220000;
      10869: inst = 32'h10408000;
      10870: inst = 32'hc404baa;
      10871: inst = 32'h8220000;
      10872: inst = 32'h10408000;
      10873: inst = 32'hc404bab;
      10874: inst = 32'h8220000;
      10875: inst = 32'h10408000;
      10876: inst = 32'hc404bac;
      10877: inst = 32'h8220000;
      10878: inst = 32'h10408000;
      10879: inst = 32'hc404bad;
      10880: inst = 32'h8220000;
      10881: inst = 32'h10408000;
      10882: inst = 32'hc404bae;
      10883: inst = 32'h8220000;
      10884: inst = 32'h10408000;
      10885: inst = 32'hc404baf;
      10886: inst = 32'h8220000;
      10887: inst = 32'h10408000;
      10888: inst = 32'hc404bb0;
      10889: inst = 32'h8220000;
      10890: inst = 32'h10408000;
      10891: inst = 32'hc404bb1;
      10892: inst = 32'h8220000;
      10893: inst = 32'h10408000;
      10894: inst = 32'hc404bb2;
      10895: inst = 32'h8220000;
      10896: inst = 32'h10408000;
      10897: inst = 32'hc404bb3;
      10898: inst = 32'h8220000;
      10899: inst = 32'h10408000;
      10900: inst = 32'hc404bb4;
      10901: inst = 32'h8220000;
      10902: inst = 32'h10408000;
      10903: inst = 32'hc404bb5;
      10904: inst = 32'h8220000;
      10905: inst = 32'h10408000;
      10906: inst = 32'hc404bb6;
      10907: inst = 32'h8220000;
      10908: inst = 32'h10408000;
      10909: inst = 32'hc404bb7;
      10910: inst = 32'h8220000;
      10911: inst = 32'h10408000;
      10912: inst = 32'hc404bb8;
      10913: inst = 32'h8220000;
      10914: inst = 32'h10408000;
      10915: inst = 32'hc404bb9;
      10916: inst = 32'h8220000;
      10917: inst = 32'h10408000;
      10918: inst = 32'hc404bba;
      10919: inst = 32'h8220000;
      10920: inst = 32'h10408000;
      10921: inst = 32'hc404bbb;
      10922: inst = 32'h8220000;
      10923: inst = 32'h10408000;
      10924: inst = 32'hc404bbc;
      10925: inst = 32'h8220000;
      10926: inst = 32'h10408000;
      10927: inst = 32'hc404bbd;
      10928: inst = 32'h8220000;
      10929: inst = 32'h10408000;
      10930: inst = 32'hc404bbe;
      10931: inst = 32'h8220000;
      10932: inst = 32'h10408000;
      10933: inst = 32'hc404bbf;
      10934: inst = 32'h8220000;
      10935: inst = 32'h10408000;
      10936: inst = 32'hc404bc0;
      10937: inst = 32'h8220000;
      10938: inst = 32'h10408000;
      10939: inst = 32'hc404bc1;
      10940: inst = 32'h8220000;
      10941: inst = 32'h10408000;
      10942: inst = 32'hc404bc2;
      10943: inst = 32'h8220000;
      10944: inst = 32'h10408000;
      10945: inst = 32'hc404bc3;
      10946: inst = 32'h8220000;
      10947: inst = 32'hc20ee75;
      10948: inst = 32'h10408000;
      10949: inst = 32'hc4042ea;
      10950: inst = 32'h8220000;
      10951: inst = 32'h10408000;
      10952: inst = 32'hc4043a7;
      10953: inst = 32'h8220000;
      10954: inst = 32'hc20d42c;
      10955: inst = 32'h10408000;
      10956: inst = 32'hc4042eb;
      10957: inst = 32'h8220000;
      10958: inst = 32'h10408000;
      10959: inst = 32'hc4042ec;
      10960: inst = 32'h8220000;
      10961: inst = 32'h10408000;
      10962: inst = 32'hc4043a8;
      10963: inst = 32'h8220000;
      10964: inst = 32'hc20ee55;
      10965: inst = 32'h10408000;
      10966: inst = 32'hc4042ed;
      10967: inst = 32'h8220000;
      10968: inst = 32'h10408000;
      10969: inst = 32'hc4043b0;
      10970: inst = 32'h8220000;
      10971: inst = 32'hc20e571;
      10972: inst = 32'h10408000;
      10973: inst = 32'hc404349;
      10974: inst = 32'h8220000;
      10975: inst = 32'h10408000;
      10976: inst = 32'hc40434e;
      10977: inst = 32'h8220000;
      10978: inst = 32'h10408000;
      10979: inst = 32'hc404406;
      10980: inst = 32'h8220000;
      10981: inst = 32'h10408000;
      10982: inst = 32'hc404411;
      10983: inst = 32'h8220000;
      10984: inst = 32'hc20cb28;
      10985: inst = 32'h10408000;
      10986: inst = 32'hc40434a;
      10987: inst = 32'h8220000;
      10988: inst = 32'h10408000;
      10989: inst = 32'hc40434d;
      10990: inst = 32'h8220000;
      10991: inst = 32'h10408000;
      10992: inst = 32'hc404407;
      10993: inst = 32'h8220000;
      10994: inst = 32'h10408000;
      10995: inst = 32'hc404410;
      10996: inst = 32'h8220000;
      10997: inst = 32'hc20cac7;
      10998: inst = 32'h10408000;
      10999: inst = 32'hc40434b;
      11000: inst = 32'h8220000;
      11001: inst = 32'h10408000;
      11002: inst = 32'hc40434c;
      11003: inst = 32'h8220000;
      11004: inst = 32'h10408000;
      11005: inst = 32'hc4043a9;
      11006: inst = 32'h8220000;
      11007: inst = 32'h10408000;
      11008: inst = 32'hc4043aa;
      11009: inst = 32'h8220000;
      11010: inst = 32'h10408000;
      11011: inst = 32'hc4043ab;
      11012: inst = 32'h8220000;
      11013: inst = 32'h10408000;
      11014: inst = 32'hc4043ac;
      11015: inst = 32'h8220000;
      11016: inst = 32'h10408000;
      11017: inst = 32'hc4043ad;
      11018: inst = 32'h8220000;
      11019: inst = 32'h10408000;
      11020: inst = 32'hc4043ae;
      11021: inst = 32'h8220000;
      11022: inst = 32'h10408000;
      11023: inst = 32'hc404408;
      11024: inst = 32'h8220000;
      11025: inst = 32'h10408000;
      11026: inst = 32'hc404409;
      11027: inst = 32'h8220000;
      11028: inst = 32'h10408000;
      11029: inst = 32'hc40440a;
      11030: inst = 32'h8220000;
      11031: inst = 32'h10408000;
      11032: inst = 32'hc40440b;
      11033: inst = 32'h8220000;
      11034: inst = 32'h10408000;
      11035: inst = 32'hc40440c;
      11036: inst = 32'h8220000;
      11037: inst = 32'h10408000;
      11038: inst = 32'hc40440d;
      11039: inst = 32'h8220000;
      11040: inst = 32'h10408000;
      11041: inst = 32'hc40440e;
      11042: inst = 32'h8220000;
      11043: inst = 32'h10408000;
      11044: inst = 32'hc40440f;
      11045: inst = 32'h8220000;
      11046: inst = 32'hc20d40c;
      11047: inst = 32'h10408000;
      11048: inst = 32'hc4043af;
      11049: inst = 32'h8220000;
      11050: inst = 32'hc20ee8e;
      11051: inst = 32'h10408000;
      11052: inst = 32'hc40446a;
      11053: inst = 32'h8220000;
      11054: inst = 32'h10408000;
      11055: inst = 32'hc4044b5;
      11056: inst = 32'h8220000;
      11057: inst = 32'hc20ee48;
      11058: inst = 32'h10408000;
      11059: inst = 32'hc40446b;
      11060: inst = 32'h8220000;
      11061: inst = 32'h10408000;
      11062: inst = 32'hc40446c;
      11063: inst = 32'h8220000;
      11064: inst = 32'h10408000;
      11065: inst = 32'hc4044b3;
      11066: inst = 32'h8220000;
      11067: inst = 32'h10408000;
      11068: inst = 32'hc4044b4;
      11069: inst = 32'h8220000;
      11070: inst = 32'hc20ee90;
      11071: inst = 32'h10408000;
      11072: inst = 32'hc40446d;
      11073: inst = 32'h8220000;
      11074: inst = 32'h10408000;
      11075: inst = 32'hc4044b2;
      11076: inst = 32'h8220000;
      11077: inst = 32'hc20eeb5;
      11078: inst = 32'h10408000;
      11079: inst = 32'hc4044cb;
      11080: inst = 32'h8220000;
      11081: inst = 32'h10408000;
      11082: inst = 32'hc4044cc;
      11083: inst = 32'h8220000;
      11084: inst = 32'h10408000;
      11085: inst = 32'hc404513;
      11086: inst = 32'h8220000;
      11087: inst = 32'h10408000;
      11088: inst = 32'hc404514;
      11089: inst = 32'h8220000;
      11090: inst = 32'hc20c2e2;
      11091: inst = 32'h10408000;
      11092: inst = 32'hc4046ef;
      11093: inst = 32'h8220000;
      11094: inst = 32'h10408000;
      11095: inst = 32'hc4046f0;
      11096: inst = 32'h8220000;
      11097: inst = 32'h10408000;
      11098: inst = 32'hc4046f1;
      11099: inst = 32'h8220000;
      11100: inst = 32'h10408000;
      11101: inst = 32'hc4046f2;
      11102: inst = 32'h8220000;
      11103: inst = 32'h10408000;
      11104: inst = 32'hc4046f3;
      11105: inst = 32'h8220000;
      11106: inst = 32'h10408000;
      11107: inst = 32'hc4046f4;
      11108: inst = 32'h8220000;
      11109: inst = 32'h10408000;
      11110: inst = 32'hc4046f5;
      11111: inst = 32'h8220000;
      11112: inst = 32'h10408000;
      11113: inst = 32'hc4046f6;
      11114: inst = 32'h8220000;
      11115: inst = 32'h10408000;
      11116: inst = 32'hc4046f7;
      11117: inst = 32'h8220000;
      11118: inst = 32'h10408000;
      11119: inst = 32'hc4046f8;
      11120: inst = 32'h8220000;
      11121: inst = 32'h10408000;
      11122: inst = 32'hc4046f9;
      11123: inst = 32'h8220000;
      11124: inst = 32'h10408000;
      11125: inst = 32'hc4046fa;
      11126: inst = 32'h8220000;
      11127: inst = 32'h10408000;
      11128: inst = 32'hc4046fb;
      11129: inst = 32'h8220000;
      11130: inst = 32'h10408000;
      11131: inst = 32'hc4046fc;
      11132: inst = 32'h8220000;
      11133: inst = 32'h10408000;
      11134: inst = 32'hc4046fd;
      11135: inst = 32'h8220000;
      11136: inst = 32'h10408000;
      11137: inst = 32'hc4046fe;
      11138: inst = 32'h8220000;
      11139: inst = 32'h10408000;
      11140: inst = 32'hc4046ff;
      11141: inst = 32'h8220000;
      11142: inst = 32'h10408000;
      11143: inst = 32'hc40474f;
      11144: inst = 32'h8220000;
      11145: inst = 32'h10408000;
      11146: inst = 32'hc40475f;
      11147: inst = 32'h8220000;
      11148: inst = 32'h10408000;
      11149: inst = 32'hc4047af;
      11150: inst = 32'h8220000;
      11151: inst = 32'h10408000;
      11152: inst = 32'hc4047bf;
      11153: inst = 32'h8220000;
      11154: inst = 32'h10408000;
      11155: inst = 32'hc40480f;
      11156: inst = 32'h8220000;
      11157: inst = 32'h10408000;
      11158: inst = 32'hc40481f;
      11159: inst = 32'h8220000;
      11160: inst = 32'h10408000;
      11161: inst = 32'hc40486f;
      11162: inst = 32'h8220000;
      11163: inst = 32'h10408000;
      11164: inst = 32'hc40487f;
      11165: inst = 32'h8220000;
      11166: inst = 32'h10408000;
      11167: inst = 32'hc4048cf;
      11168: inst = 32'h8220000;
      11169: inst = 32'h10408000;
      11170: inst = 32'hc4048df;
      11171: inst = 32'h8220000;
      11172: inst = 32'h10408000;
      11173: inst = 32'hc40492f;
      11174: inst = 32'h8220000;
      11175: inst = 32'h10408000;
      11176: inst = 32'hc40493f;
      11177: inst = 32'h8220000;
      11178: inst = 32'h10408000;
      11179: inst = 32'hc40498f;
      11180: inst = 32'h8220000;
      11181: inst = 32'h10408000;
      11182: inst = 32'hc40499f;
      11183: inst = 32'h8220000;
      11184: inst = 32'h10408000;
      11185: inst = 32'hc4049ef;
      11186: inst = 32'h8220000;
      11187: inst = 32'h10408000;
      11188: inst = 32'hc4049ff;
      11189: inst = 32'h8220000;
      11190: inst = 32'h10408000;
      11191: inst = 32'hc404a4f;
      11192: inst = 32'h8220000;
      11193: inst = 32'h10408000;
      11194: inst = 32'hc404a5f;
      11195: inst = 32'h8220000;
      11196: inst = 32'h10408000;
      11197: inst = 32'hc404aaf;
      11198: inst = 32'h8220000;
      11199: inst = 32'h10408000;
      11200: inst = 32'hc404abf;
      11201: inst = 32'h8220000;
      11202: inst = 32'h10408000;
      11203: inst = 32'hc404b0f;
      11204: inst = 32'h8220000;
      11205: inst = 32'h10408000;
      11206: inst = 32'hc404b1f;
      11207: inst = 32'h8220000;
      11208: inst = 32'h10408000;
      11209: inst = 32'hc404b6f;
      11210: inst = 32'h8220000;
      11211: inst = 32'h10408000;
      11212: inst = 32'hc404b7f;
      11213: inst = 32'h8220000;
      11214: inst = 32'h10408000;
      11215: inst = 32'hc404bcf;
      11216: inst = 32'h8220000;
      11217: inst = 32'h10408000;
      11218: inst = 32'hc404bdf;
      11219: inst = 32'h8220000;
      11220: inst = 32'h10408000;
      11221: inst = 32'hc404c2f;
      11222: inst = 32'h8220000;
      11223: inst = 32'h10408000;
      11224: inst = 32'hc404c3f;
      11225: inst = 32'h8220000;
      11226: inst = 32'h10408000;
      11227: inst = 32'hc404c8f;
      11228: inst = 32'h8220000;
      11229: inst = 32'h10408000;
      11230: inst = 32'hc404c9f;
      11231: inst = 32'h8220000;
      11232: inst = 32'h10408000;
      11233: inst = 32'hc404cef;
      11234: inst = 32'h8220000;
      11235: inst = 32'h10408000;
      11236: inst = 32'hc404cff;
      11237: inst = 32'h8220000;
      11238: inst = 32'h10408000;
      11239: inst = 32'hc404d4f;
      11240: inst = 32'h8220000;
      11241: inst = 32'h10408000;
      11242: inst = 32'hc404d5f;
      11243: inst = 32'h8220000;
      11244: inst = 32'h10408000;
      11245: inst = 32'hc404daf;
      11246: inst = 32'h8220000;
      11247: inst = 32'h10408000;
      11248: inst = 32'hc404dbf;
      11249: inst = 32'h8220000;
      11250: inst = 32'h10408000;
      11251: inst = 32'hc404e0f;
      11252: inst = 32'h8220000;
      11253: inst = 32'h10408000;
      11254: inst = 32'hc404e1f;
      11255: inst = 32'h8220000;
      11256: inst = 32'h10408000;
      11257: inst = 32'hc404e6f;
      11258: inst = 32'h8220000;
      11259: inst = 32'h10408000;
      11260: inst = 32'hc404e7f;
      11261: inst = 32'h8220000;
      11262: inst = 32'h10408000;
      11263: inst = 32'hc404ecf;
      11264: inst = 32'h8220000;
      11265: inst = 32'h10408000;
      11266: inst = 32'hc404edf;
      11267: inst = 32'h8220000;
      11268: inst = 32'h10408000;
      11269: inst = 32'hc404f2f;
      11270: inst = 32'h8220000;
      11271: inst = 32'h10408000;
      11272: inst = 32'hc404f3f;
      11273: inst = 32'h8220000;
      11274: inst = 32'h10408000;
      11275: inst = 32'hc404f8f;
      11276: inst = 32'h8220000;
      11277: inst = 32'h10408000;
      11278: inst = 32'hc404f9f;
      11279: inst = 32'h8220000;
      11280: inst = 32'h10408000;
      11281: inst = 32'hc404fef;
      11282: inst = 32'h8220000;
      11283: inst = 32'h10408000;
      11284: inst = 32'hc404fff;
      11285: inst = 32'h8220000;
      11286: inst = 32'h10408000;
      11287: inst = 32'hc40504f;
      11288: inst = 32'h8220000;
      11289: inst = 32'h10408000;
      11290: inst = 32'hc40505f;
      11291: inst = 32'h8220000;
      11292: inst = 32'h10408000;
      11293: inst = 32'hc4050af;
      11294: inst = 32'h8220000;
      11295: inst = 32'h10408000;
      11296: inst = 32'hc4050bf;
      11297: inst = 32'h8220000;
      11298: inst = 32'h10408000;
      11299: inst = 32'hc40510f;
      11300: inst = 32'h8220000;
      11301: inst = 32'h10408000;
      11302: inst = 32'hc40511f;
      11303: inst = 32'h8220000;
      11304: inst = 32'h10408000;
      11305: inst = 32'hc40516f;
      11306: inst = 32'h8220000;
      11307: inst = 32'h10408000;
      11308: inst = 32'hc40517f;
      11309: inst = 32'h8220000;
      11310: inst = 32'h10408000;
      11311: inst = 32'hc4051cf;
      11312: inst = 32'h8220000;
      11313: inst = 32'h10408000;
      11314: inst = 32'hc4051df;
      11315: inst = 32'h8220000;
      11316: inst = 32'h10408000;
      11317: inst = 32'hc40522f;
      11318: inst = 32'h8220000;
      11319: inst = 32'h10408000;
      11320: inst = 32'hc40523f;
      11321: inst = 32'h8220000;
      11322: inst = 32'h10408000;
      11323: inst = 32'hc40528f;
      11324: inst = 32'h8220000;
      11325: inst = 32'h10408000;
      11326: inst = 32'hc40529f;
      11327: inst = 32'h8220000;
      11328: inst = 32'h10408000;
      11329: inst = 32'hc4052ef;
      11330: inst = 32'h8220000;
      11331: inst = 32'h10408000;
      11332: inst = 32'hc4052f0;
      11333: inst = 32'h8220000;
      11334: inst = 32'h10408000;
      11335: inst = 32'hc4052f1;
      11336: inst = 32'h8220000;
      11337: inst = 32'h10408000;
      11338: inst = 32'hc4052f2;
      11339: inst = 32'h8220000;
      11340: inst = 32'h10408000;
      11341: inst = 32'hc4052f3;
      11342: inst = 32'h8220000;
      11343: inst = 32'h10408000;
      11344: inst = 32'hc4052f4;
      11345: inst = 32'h8220000;
      11346: inst = 32'h10408000;
      11347: inst = 32'hc4052f5;
      11348: inst = 32'h8220000;
      11349: inst = 32'h10408000;
      11350: inst = 32'hc4052f6;
      11351: inst = 32'h8220000;
      11352: inst = 32'h10408000;
      11353: inst = 32'hc4052f7;
      11354: inst = 32'h8220000;
      11355: inst = 32'h10408000;
      11356: inst = 32'hc4052f8;
      11357: inst = 32'h8220000;
      11358: inst = 32'h10408000;
      11359: inst = 32'hc4052f9;
      11360: inst = 32'h8220000;
      11361: inst = 32'h10408000;
      11362: inst = 32'hc4052fa;
      11363: inst = 32'h8220000;
      11364: inst = 32'h10408000;
      11365: inst = 32'hc4052fb;
      11366: inst = 32'h8220000;
      11367: inst = 32'h10408000;
      11368: inst = 32'hc4052fc;
      11369: inst = 32'h8220000;
      11370: inst = 32'h10408000;
      11371: inst = 32'hc4052fd;
      11372: inst = 32'h8220000;
      11373: inst = 32'h10408000;
      11374: inst = 32'hc4052fe;
      11375: inst = 32'h8220000;
      11376: inst = 32'h10408000;
      11377: inst = 32'hc4052ff;
      11378: inst = 32'h8220000;
      11379: inst = 32'hc20dbc5;
      11380: inst = 32'h10408000;
      11381: inst = 32'hc404750;
      11382: inst = 32'h8220000;
      11383: inst = 32'h10408000;
      11384: inst = 32'hc404751;
      11385: inst = 32'h8220000;
      11386: inst = 32'h10408000;
      11387: inst = 32'hc404752;
      11388: inst = 32'h8220000;
      11389: inst = 32'h10408000;
      11390: inst = 32'hc404753;
      11391: inst = 32'h8220000;
      11392: inst = 32'h10408000;
      11393: inst = 32'hc404754;
      11394: inst = 32'h8220000;
      11395: inst = 32'h10408000;
      11396: inst = 32'hc404755;
      11397: inst = 32'h8220000;
      11398: inst = 32'h10408000;
      11399: inst = 32'hc404756;
      11400: inst = 32'h8220000;
      11401: inst = 32'h10408000;
      11402: inst = 32'hc404757;
      11403: inst = 32'h8220000;
      11404: inst = 32'h10408000;
      11405: inst = 32'hc404758;
      11406: inst = 32'h8220000;
      11407: inst = 32'h10408000;
      11408: inst = 32'hc404759;
      11409: inst = 32'h8220000;
      11410: inst = 32'h10408000;
      11411: inst = 32'hc40475a;
      11412: inst = 32'h8220000;
      11413: inst = 32'h10408000;
      11414: inst = 32'hc40475b;
      11415: inst = 32'h8220000;
      11416: inst = 32'h10408000;
      11417: inst = 32'hc40475c;
      11418: inst = 32'h8220000;
      11419: inst = 32'h10408000;
      11420: inst = 32'hc40475d;
      11421: inst = 32'h8220000;
      11422: inst = 32'h10408000;
      11423: inst = 32'hc40475e;
      11424: inst = 32'h8220000;
      11425: inst = 32'h10408000;
      11426: inst = 32'hc4047b0;
      11427: inst = 32'h8220000;
      11428: inst = 32'h10408000;
      11429: inst = 32'hc4047b1;
      11430: inst = 32'h8220000;
      11431: inst = 32'h10408000;
      11432: inst = 32'hc4047b2;
      11433: inst = 32'h8220000;
      11434: inst = 32'h10408000;
      11435: inst = 32'hc4047b3;
      11436: inst = 32'h8220000;
      11437: inst = 32'h10408000;
      11438: inst = 32'hc4047b4;
      11439: inst = 32'h8220000;
      11440: inst = 32'h10408000;
      11441: inst = 32'hc4047b5;
      11442: inst = 32'h8220000;
      11443: inst = 32'h10408000;
      11444: inst = 32'hc4047b6;
      11445: inst = 32'h8220000;
      11446: inst = 32'h10408000;
      11447: inst = 32'hc4047b7;
      11448: inst = 32'h8220000;
      11449: inst = 32'h10408000;
      11450: inst = 32'hc4047b8;
      11451: inst = 32'h8220000;
      11452: inst = 32'h10408000;
      11453: inst = 32'hc4047b9;
      11454: inst = 32'h8220000;
      11455: inst = 32'h10408000;
      11456: inst = 32'hc4047ba;
      11457: inst = 32'h8220000;
      11458: inst = 32'h10408000;
      11459: inst = 32'hc4047bb;
      11460: inst = 32'h8220000;
      11461: inst = 32'h10408000;
      11462: inst = 32'hc4047bc;
      11463: inst = 32'h8220000;
      11464: inst = 32'h10408000;
      11465: inst = 32'hc4047bd;
      11466: inst = 32'h8220000;
      11467: inst = 32'h10408000;
      11468: inst = 32'hc4047be;
      11469: inst = 32'h8220000;
      11470: inst = 32'h10408000;
      11471: inst = 32'hc404810;
      11472: inst = 32'h8220000;
      11473: inst = 32'h10408000;
      11474: inst = 32'hc404811;
      11475: inst = 32'h8220000;
      11476: inst = 32'h10408000;
      11477: inst = 32'hc404812;
      11478: inst = 32'h8220000;
      11479: inst = 32'h10408000;
      11480: inst = 32'hc404813;
      11481: inst = 32'h8220000;
      11482: inst = 32'h10408000;
      11483: inst = 32'hc404814;
      11484: inst = 32'h8220000;
      11485: inst = 32'h10408000;
      11486: inst = 32'hc404815;
      11487: inst = 32'h8220000;
      11488: inst = 32'h10408000;
      11489: inst = 32'hc404816;
      11490: inst = 32'h8220000;
      11491: inst = 32'h10408000;
      11492: inst = 32'hc404817;
      11493: inst = 32'h8220000;
      11494: inst = 32'h10408000;
      11495: inst = 32'hc404818;
      11496: inst = 32'h8220000;
      11497: inst = 32'h10408000;
      11498: inst = 32'hc404819;
      11499: inst = 32'h8220000;
      11500: inst = 32'h10408000;
      11501: inst = 32'hc40481a;
      11502: inst = 32'h8220000;
      11503: inst = 32'h10408000;
      11504: inst = 32'hc40481b;
      11505: inst = 32'h8220000;
      11506: inst = 32'h10408000;
      11507: inst = 32'hc40481c;
      11508: inst = 32'h8220000;
      11509: inst = 32'h10408000;
      11510: inst = 32'hc40481d;
      11511: inst = 32'h8220000;
      11512: inst = 32'h10408000;
      11513: inst = 32'hc40481e;
      11514: inst = 32'h8220000;
      11515: inst = 32'h10408000;
      11516: inst = 32'hc404870;
      11517: inst = 32'h8220000;
      11518: inst = 32'h10408000;
      11519: inst = 32'hc404871;
      11520: inst = 32'h8220000;
      11521: inst = 32'h10408000;
      11522: inst = 32'hc404872;
      11523: inst = 32'h8220000;
      11524: inst = 32'h10408000;
      11525: inst = 32'hc404873;
      11526: inst = 32'h8220000;
      11527: inst = 32'h10408000;
      11528: inst = 32'hc404874;
      11529: inst = 32'h8220000;
      11530: inst = 32'h10408000;
      11531: inst = 32'hc404875;
      11532: inst = 32'h8220000;
      11533: inst = 32'h10408000;
      11534: inst = 32'hc404876;
      11535: inst = 32'h8220000;
      11536: inst = 32'h10408000;
      11537: inst = 32'hc404877;
      11538: inst = 32'h8220000;
      11539: inst = 32'h10408000;
      11540: inst = 32'hc404878;
      11541: inst = 32'h8220000;
      11542: inst = 32'h10408000;
      11543: inst = 32'hc404879;
      11544: inst = 32'h8220000;
      11545: inst = 32'h10408000;
      11546: inst = 32'hc40487a;
      11547: inst = 32'h8220000;
      11548: inst = 32'h10408000;
      11549: inst = 32'hc40487b;
      11550: inst = 32'h8220000;
      11551: inst = 32'h10408000;
      11552: inst = 32'hc40487c;
      11553: inst = 32'h8220000;
      11554: inst = 32'h10408000;
      11555: inst = 32'hc40487d;
      11556: inst = 32'h8220000;
      11557: inst = 32'h10408000;
      11558: inst = 32'hc40487e;
      11559: inst = 32'h8220000;
      11560: inst = 32'h10408000;
      11561: inst = 32'hc4048d0;
      11562: inst = 32'h8220000;
      11563: inst = 32'h10408000;
      11564: inst = 32'hc4048d1;
      11565: inst = 32'h8220000;
      11566: inst = 32'h10408000;
      11567: inst = 32'hc4048d2;
      11568: inst = 32'h8220000;
      11569: inst = 32'h10408000;
      11570: inst = 32'hc4048d3;
      11571: inst = 32'h8220000;
      11572: inst = 32'h10408000;
      11573: inst = 32'hc4048d4;
      11574: inst = 32'h8220000;
      11575: inst = 32'h10408000;
      11576: inst = 32'hc4048d5;
      11577: inst = 32'h8220000;
      11578: inst = 32'h10408000;
      11579: inst = 32'hc4048d6;
      11580: inst = 32'h8220000;
      11581: inst = 32'h10408000;
      11582: inst = 32'hc4048d7;
      11583: inst = 32'h8220000;
      11584: inst = 32'h10408000;
      11585: inst = 32'hc4048d8;
      11586: inst = 32'h8220000;
      11587: inst = 32'h10408000;
      11588: inst = 32'hc4048d9;
      11589: inst = 32'h8220000;
      11590: inst = 32'h10408000;
      11591: inst = 32'hc4048da;
      11592: inst = 32'h8220000;
      11593: inst = 32'h10408000;
      11594: inst = 32'hc4048db;
      11595: inst = 32'h8220000;
      11596: inst = 32'h10408000;
      11597: inst = 32'hc4048dc;
      11598: inst = 32'h8220000;
      11599: inst = 32'h10408000;
      11600: inst = 32'hc4048dd;
      11601: inst = 32'h8220000;
      11602: inst = 32'h10408000;
      11603: inst = 32'hc4048de;
      11604: inst = 32'h8220000;
      11605: inst = 32'h10408000;
      11606: inst = 32'hc404930;
      11607: inst = 32'h8220000;
      11608: inst = 32'h10408000;
      11609: inst = 32'hc404931;
      11610: inst = 32'h8220000;
      11611: inst = 32'h10408000;
      11612: inst = 32'hc404936;
      11613: inst = 32'h8220000;
      11614: inst = 32'h10408000;
      11615: inst = 32'hc404937;
      11616: inst = 32'h8220000;
      11617: inst = 32'h10408000;
      11618: inst = 32'hc404938;
      11619: inst = 32'h8220000;
      11620: inst = 32'h10408000;
      11621: inst = 32'hc404939;
      11622: inst = 32'h8220000;
      11623: inst = 32'h10408000;
      11624: inst = 32'hc40493a;
      11625: inst = 32'h8220000;
      11626: inst = 32'h10408000;
      11627: inst = 32'hc40493b;
      11628: inst = 32'h8220000;
      11629: inst = 32'h10408000;
      11630: inst = 32'hc40493c;
      11631: inst = 32'h8220000;
      11632: inst = 32'h10408000;
      11633: inst = 32'hc40493d;
      11634: inst = 32'h8220000;
      11635: inst = 32'h10408000;
      11636: inst = 32'hc40493e;
      11637: inst = 32'h8220000;
      11638: inst = 32'h10408000;
      11639: inst = 32'hc404990;
      11640: inst = 32'h8220000;
      11641: inst = 32'h10408000;
      11642: inst = 32'hc404991;
      11643: inst = 32'h8220000;
      11644: inst = 32'h10408000;
      11645: inst = 32'hc404996;
      11646: inst = 32'h8220000;
      11647: inst = 32'h10408000;
      11648: inst = 32'hc404997;
      11649: inst = 32'h8220000;
      11650: inst = 32'h10408000;
      11651: inst = 32'hc404998;
      11652: inst = 32'h8220000;
      11653: inst = 32'h10408000;
      11654: inst = 32'hc404999;
      11655: inst = 32'h8220000;
      11656: inst = 32'h10408000;
      11657: inst = 32'hc40499a;
      11658: inst = 32'h8220000;
      11659: inst = 32'h10408000;
      11660: inst = 32'hc40499b;
      11661: inst = 32'h8220000;
      11662: inst = 32'h10408000;
      11663: inst = 32'hc40499c;
      11664: inst = 32'h8220000;
      11665: inst = 32'h10408000;
      11666: inst = 32'hc40499d;
      11667: inst = 32'h8220000;
      11668: inst = 32'h10408000;
      11669: inst = 32'hc40499e;
      11670: inst = 32'h8220000;
      11671: inst = 32'h10408000;
      11672: inst = 32'hc4049f0;
      11673: inst = 32'h8220000;
      11674: inst = 32'h10408000;
      11675: inst = 32'hc4049f1;
      11676: inst = 32'h8220000;
      11677: inst = 32'h10408000;
      11678: inst = 32'hc4049f6;
      11679: inst = 32'h8220000;
      11680: inst = 32'h10408000;
      11681: inst = 32'hc4049f7;
      11682: inst = 32'h8220000;
      11683: inst = 32'h10408000;
      11684: inst = 32'hc4049f8;
      11685: inst = 32'h8220000;
      11686: inst = 32'h10408000;
      11687: inst = 32'hc4049f9;
      11688: inst = 32'h8220000;
      11689: inst = 32'h10408000;
      11690: inst = 32'hc4049fa;
      11691: inst = 32'h8220000;
      11692: inst = 32'h10408000;
      11693: inst = 32'hc4049fb;
      11694: inst = 32'h8220000;
      11695: inst = 32'h10408000;
      11696: inst = 32'hc4049fc;
      11697: inst = 32'h8220000;
      11698: inst = 32'h10408000;
      11699: inst = 32'hc4049fd;
      11700: inst = 32'h8220000;
      11701: inst = 32'h10408000;
      11702: inst = 32'hc4049fe;
      11703: inst = 32'h8220000;
      11704: inst = 32'h10408000;
      11705: inst = 32'hc404a50;
      11706: inst = 32'h8220000;
      11707: inst = 32'h10408000;
      11708: inst = 32'hc404a51;
      11709: inst = 32'h8220000;
      11710: inst = 32'h10408000;
      11711: inst = 32'hc404a56;
      11712: inst = 32'h8220000;
      11713: inst = 32'h10408000;
      11714: inst = 32'hc404a57;
      11715: inst = 32'h8220000;
      11716: inst = 32'h10408000;
      11717: inst = 32'hc404a58;
      11718: inst = 32'h8220000;
      11719: inst = 32'h10408000;
      11720: inst = 32'hc404a59;
      11721: inst = 32'h8220000;
      11722: inst = 32'h10408000;
      11723: inst = 32'hc404a5a;
      11724: inst = 32'h8220000;
      11725: inst = 32'h10408000;
      11726: inst = 32'hc404a5b;
      11727: inst = 32'h8220000;
      11728: inst = 32'h10408000;
      11729: inst = 32'hc404a5c;
      11730: inst = 32'h8220000;
      11731: inst = 32'h10408000;
      11732: inst = 32'hc404a5d;
      11733: inst = 32'h8220000;
      11734: inst = 32'h10408000;
      11735: inst = 32'hc404a5e;
      11736: inst = 32'h8220000;
      11737: inst = 32'h10408000;
      11738: inst = 32'hc404ab0;
      11739: inst = 32'h8220000;
      11740: inst = 32'h10408000;
      11741: inst = 32'hc404ab1;
      11742: inst = 32'h8220000;
      11743: inst = 32'h10408000;
      11744: inst = 32'hc404ab6;
      11745: inst = 32'h8220000;
      11746: inst = 32'h10408000;
      11747: inst = 32'hc404ab7;
      11748: inst = 32'h8220000;
      11749: inst = 32'h10408000;
      11750: inst = 32'hc404ab8;
      11751: inst = 32'h8220000;
      11752: inst = 32'h10408000;
      11753: inst = 32'hc404ab9;
      11754: inst = 32'h8220000;
      11755: inst = 32'h10408000;
      11756: inst = 32'hc404aba;
      11757: inst = 32'h8220000;
      11758: inst = 32'h10408000;
      11759: inst = 32'hc404abb;
      11760: inst = 32'h8220000;
      11761: inst = 32'h10408000;
      11762: inst = 32'hc404abc;
      11763: inst = 32'h8220000;
      11764: inst = 32'h10408000;
      11765: inst = 32'hc404abd;
      11766: inst = 32'h8220000;
      11767: inst = 32'h10408000;
      11768: inst = 32'hc404abe;
      11769: inst = 32'h8220000;
      11770: inst = 32'h10408000;
      11771: inst = 32'hc404b10;
      11772: inst = 32'h8220000;
      11773: inst = 32'h10408000;
      11774: inst = 32'hc404b11;
      11775: inst = 32'h8220000;
      11776: inst = 32'h10408000;
      11777: inst = 32'hc404b16;
      11778: inst = 32'h8220000;
      11779: inst = 32'h10408000;
      11780: inst = 32'hc404b17;
      11781: inst = 32'h8220000;
      11782: inst = 32'h10408000;
      11783: inst = 32'hc404b18;
      11784: inst = 32'h8220000;
      11785: inst = 32'h10408000;
      11786: inst = 32'hc404b19;
      11787: inst = 32'h8220000;
      11788: inst = 32'h10408000;
      11789: inst = 32'hc404b1a;
      11790: inst = 32'h8220000;
      11791: inst = 32'h10408000;
      11792: inst = 32'hc404b1b;
      11793: inst = 32'h8220000;
      11794: inst = 32'h10408000;
      11795: inst = 32'hc404b1c;
      11796: inst = 32'h8220000;
      11797: inst = 32'h10408000;
      11798: inst = 32'hc404b1d;
      11799: inst = 32'h8220000;
      11800: inst = 32'h10408000;
      11801: inst = 32'hc404b1e;
      11802: inst = 32'h8220000;
      11803: inst = 32'h10408000;
      11804: inst = 32'hc404b70;
      11805: inst = 32'h8220000;
      11806: inst = 32'h10408000;
      11807: inst = 32'hc404b71;
      11808: inst = 32'h8220000;
      11809: inst = 32'h10408000;
      11810: inst = 32'hc404b76;
      11811: inst = 32'h8220000;
      11812: inst = 32'h10408000;
      11813: inst = 32'hc404b77;
      11814: inst = 32'h8220000;
      11815: inst = 32'h10408000;
      11816: inst = 32'hc404b78;
      11817: inst = 32'h8220000;
      11818: inst = 32'h10408000;
      11819: inst = 32'hc404b79;
      11820: inst = 32'h8220000;
      11821: inst = 32'h10408000;
      11822: inst = 32'hc404b7a;
      11823: inst = 32'h8220000;
      11824: inst = 32'h10408000;
      11825: inst = 32'hc404b7b;
      11826: inst = 32'h8220000;
      11827: inst = 32'h10408000;
      11828: inst = 32'hc404b7c;
      11829: inst = 32'h8220000;
      11830: inst = 32'h10408000;
      11831: inst = 32'hc404b7d;
      11832: inst = 32'h8220000;
      11833: inst = 32'h10408000;
      11834: inst = 32'hc404b7e;
      11835: inst = 32'h8220000;
      11836: inst = 32'h10408000;
      11837: inst = 32'hc404bd0;
      11838: inst = 32'h8220000;
      11839: inst = 32'h10408000;
      11840: inst = 32'hc404bd1;
      11841: inst = 32'h8220000;
      11842: inst = 32'h10408000;
      11843: inst = 32'hc404bd2;
      11844: inst = 32'h8220000;
      11845: inst = 32'h10408000;
      11846: inst = 32'hc404bd3;
      11847: inst = 32'h8220000;
      11848: inst = 32'h10408000;
      11849: inst = 32'hc404bd4;
      11850: inst = 32'h8220000;
      11851: inst = 32'h10408000;
      11852: inst = 32'hc404bd5;
      11853: inst = 32'h8220000;
      11854: inst = 32'h10408000;
      11855: inst = 32'hc404bd6;
      11856: inst = 32'h8220000;
      11857: inst = 32'h10408000;
      11858: inst = 32'hc404bd7;
      11859: inst = 32'h8220000;
      11860: inst = 32'h10408000;
      11861: inst = 32'hc404bd8;
      11862: inst = 32'h8220000;
      11863: inst = 32'h10408000;
      11864: inst = 32'hc404bd9;
      11865: inst = 32'h8220000;
      11866: inst = 32'h10408000;
      11867: inst = 32'hc404bda;
      11868: inst = 32'h8220000;
      11869: inst = 32'h10408000;
      11870: inst = 32'hc404bdb;
      11871: inst = 32'h8220000;
      11872: inst = 32'h10408000;
      11873: inst = 32'hc404bdc;
      11874: inst = 32'h8220000;
      11875: inst = 32'h10408000;
      11876: inst = 32'hc404bdd;
      11877: inst = 32'h8220000;
      11878: inst = 32'h10408000;
      11879: inst = 32'hc404bde;
      11880: inst = 32'h8220000;
      11881: inst = 32'h10408000;
      11882: inst = 32'hc404c30;
      11883: inst = 32'h8220000;
      11884: inst = 32'h10408000;
      11885: inst = 32'hc404c31;
      11886: inst = 32'h8220000;
      11887: inst = 32'h10408000;
      11888: inst = 32'hc404c32;
      11889: inst = 32'h8220000;
      11890: inst = 32'h10408000;
      11891: inst = 32'hc404c33;
      11892: inst = 32'h8220000;
      11893: inst = 32'h10408000;
      11894: inst = 32'hc404c34;
      11895: inst = 32'h8220000;
      11896: inst = 32'h10408000;
      11897: inst = 32'hc404c35;
      11898: inst = 32'h8220000;
      11899: inst = 32'h10408000;
      11900: inst = 32'hc404c36;
      11901: inst = 32'h8220000;
      11902: inst = 32'h10408000;
      11903: inst = 32'hc404c37;
      11904: inst = 32'h8220000;
      11905: inst = 32'h10408000;
      11906: inst = 32'hc404c38;
      11907: inst = 32'h8220000;
      11908: inst = 32'h10408000;
      11909: inst = 32'hc404c39;
      11910: inst = 32'h8220000;
      11911: inst = 32'h10408000;
      11912: inst = 32'hc404c3a;
      11913: inst = 32'h8220000;
      11914: inst = 32'h10408000;
      11915: inst = 32'hc404c3b;
      11916: inst = 32'h8220000;
      11917: inst = 32'h10408000;
      11918: inst = 32'hc404c3c;
      11919: inst = 32'h8220000;
      11920: inst = 32'h10408000;
      11921: inst = 32'hc404c3d;
      11922: inst = 32'h8220000;
      11923: inst = 32'h10408000;
      11924: inst = 32'hc404c3e;
      11925: inst = 32'h8220000;
      11926: inst = 32'h10408000;
      11927: inst = 32'hc404c90;
      11928: inst = 32'h8220000;
      11929: inst = 32'h10408000;
      11930: inst = 32'hc404c91;
      11931: inst = 32'h8220000;
      11932: inst = 32'h10408000;
      11933: inst = 32'hc404c92;
      11934: inst = 32'h8220000;
      11935: inst = 32'h10408000;
      11936: inst = 32'hc404c93;
      11937: inst = 32'h8220000;
      11938: inst = 32'h10408000;
      11939: inst = 32'hc404c94;
      11940: inst = 32'h8220000;
      11941: inst = 32'h10408000;
      11942: inst = 32'hc404c95;
      11943: inst = 32'h8220000;
      11944: inst = 32'h10408000;
      11945: inst = 32'hc404c96;
      11946: inst = 32'h8220000;
      11947: inst = 32'h10408000;
      11948: inst = 32'hc404c97;
      11949: inst = 32'h8220000;
      11950: inst = 32'h10408000;
      11951: inst = 32'hc404c98;
      11952: inst = 32'h8220000;
      11953: inst = 32'h10408000;
      11954: inst = 32'hc404c99;
      11955: inst = 32'h8220000;
      11956: inst = 32'h10408000;
      11957: inst = 32'hc404c9a;
      11958: inst = 32'h8220000;
      11959: inst = 32'h10408000;
      11960: inst = 32'hc404c9b;
      11961: inst = 32'h8220000;
      11962: inst = 32'h10408000;
      11963: inst = 32'hc404c9c;
      11964: inst = 32'h8220000;
      11965: inst = 32'h10408000;
      11966: inst = 32'hc404c9d;
      11967: inst = 32'h8220000;
      11968: inst = 32'h10408000;
      11969: inst = 32'hc404c9e;
      11970: inst = 32'h8220000;
      11971: inst = 32'h10408000;
      11972: inst = 32'hc404cf0;
      11973: inst = 32'h8220000;
      11974: inst = 32'h10408000;
      11975: inst = 32'hc404cf1;
      11976: inst = 32'h8220000;
      11977: inst = 32'h10408000;
      11978: inst = 32'hc404cf2;
      11979: inst = 32'h8220000;
      11980: inst = 32'h10408000;
      11981: inst = 32'hc404cf3;
      11982: inst = 32'h8220000;
      11983: inst = 32'h10408000;
      11984: inst = 32'hc404cf4;
      11985: inst = 32'h8220000;
      11986: inst = 32'h10408000;
      11987: inst = 32'hc404cf5;
      11988: inst = 32'h8220000;
      11989: inst = 32'h10408000;
      11990: inst = 32'hc404cf6;
      11991: inst = 32'h8220000;
      11992: inst = 32'h10408000;
      11993: inst = 32'hc404cf7;
      11994: inst = 32'h8220000;
      11995: inst = 32'h10408000;
      11996: inst = 32'hc404cf8;
      11997: inst = 32'h8220000;
      11998: inst = 32'h10408000;
      11999: inst = 32'hc404cf9;
      12000: inst = 32'h8220000;
      12001: inst = 32'h10408000;
      12002: inst = 32'hc404cfa;
      12003: inst = 32'h8220000;
      12004: inst = 32'h10408000;
      12005: inst = 32'hc404cfe;
      12006: inst = 32'h8220000;
      12007: inst = 32'h10408000;
      12008: inst = 32'hc404d50;
      12009: inst = 32'h8220000;
      12010: inst = 32'h10408000;
      12011: inst = 32'hc404d51;
      12012: inst = 32'h8220000;
      12013: inst = 32'h10408000;
      12014: inst = 32'hc404d52;
      12015: inst = 32'h8220000;
      12016: inst = 32'h10408000;
      12017: inst = 32'hc404d53;
      12018: inst = 32'h8220000;
      12019: inst = 32'h10408000;
      12020: inst = 32'hc404d54;
      12021: inst = 32'h8220000;
      12022: inst = 32'h10408000;
      12023: inst = 32'hc404d55;
      12024: inst = 32'h8220000;
      12025: inst = 32'h10408000;
      12026: inst = 32'hc404d56;
      12027: inst = 32'h8220000;
      12028: inst = 32'h10408000;
      12029: inst = 32'hc404d57;
      12030: inst = 32'h8220000;
      12031: inst = 32'h10408000;
      12032: inst = 32'hc404d58;
      12033: inst = 32'h8220000;
      12034: inst = 32'h10408000;
      12035: inst = 32'hc404d59;
      12036: inst = 32'h8220000;
      12037: inst = 32'h10408000;
      12038: inst = 32'hc404d5a;
      12039: inst = 32'h8220000;
      12040: inst = 32'h10408000;
      12041: inst = 32'hc404d5c;
      12042: inst = 32'h8220000;
      12043: inst = 32'h10408000;
      12044: inst = 32'hc404d5d;
      12045: inst = 32'h8220000;
      12046: inst = 32'h10408000;
      12047: inst = 32'hc404d5e;
      12048: inst = 32'h8220000;
      12049: inst = 32'h10408000;
      12050: inst = 32'hc404db0;
      12051: inst = 32'h8220000;
      12052: inst = 32'h10408000;
      12053: inst = 32'hc404db1;
      12054: inst = 32'h8220000;
      12055: inst = 32'h10408000;
      12056: inst = 32'hc404db2;
      12057: inst = 32'h8220000;
      12058: inst = 32'h10408000;
      12059: inst = 32'hc404db3;
      12060: inst = 32'h8220000;
      12061: inst = 32'h10408000;
      12062: inst = 32'hc404db4;
      12063: inst = 32'h8220000;
      12064: inst = 32'h10408000;
      12065: inst = 32'hc404db5;
      12066: inst = 32'h8220000;
      12067: inst = 32'h10408000;
      12068: inst = 32'hc404db6;
      12069: inst = 32'h8220000;
      12070: inst = 32'h10408000;
      12071: inst = 32'hc404db7;
      12072: inst = 32'h8220000;
      12073: inst = 32'h10408000;
      12074: inst = 32'hc404db8;
      12075: inst = 32'h8220000;
      12076: inst = 32'h10408000;
      12077: inst = 32'hc404db9;
      12078: inst = 32'h8220000;
      12079: inst = 32'h10408000;
      12080: inst = 32'hc404dba;
      12081: inst = 32'h8220000;
      12082: inst = 32'h10408000;
      12083: inst = 32'hc404dbb;
      12084: inst = 32'h8220000;
      12085: inst = 32'h10408000;
      12086: inst = 32'hc404dbc;
      12087: inst = 32'h8220000;
      12088: inst = 32'h10408000;
      12089: inst = 32'hc404dbd;
      12090: inst = 32'h8220000;
      12091: inst = 32'h10408000;
      12092: inst = 32'hc404dbe;
      12093: inst = 32'h8220000;
      12094: inst = 32'h10408000;
      12095: inst = 32'hc404e10;
      12096: inst = 32'h8220000;
      12097: inst = 32'h10408000;
      12098: inst = 32'hc404e11;
      12099: inst = 32'h8220000;
      12100: inst = 32'h10408000;
      12101: inst = 32'hc404e12;
      12102: inst = 32'h8220000;
      12103: inst = 32'h10408000;
      12104: inst = 32'hc404e13;
      12105: inst = 32'h8220000;
      12106: inst = 32'h10408000;
      12107: inst = 32'hc404e14;
      12108: inst = 32'h8220000;
      12109: inst = 32'h10408000;
      12110: inst = 32'hc404e15;
      12111: inst = 32'h8220000;
      12112: inst = 32'h10408000;
      12113: inst = 32'hc404e16;
      12114: inst = 32'h8220000;
      12115: inst = 32'h10408000;
      12116: inst = 32'hc404e17;
      12117: inst = 32'h8220000;
      12118: inst = 32'h10408000;
      12119: inst = 32'hc404e18;
      12120: inst = 32'h8220000;
      12121: inst = 32'h10408000;
      12122: inst = 32'hc404e19;
      12123: inst = 32'h8220000;
      12124: inst = 32'h10408000;
      12125: inst = 32'hc404e1a;
      12126: inst = 32'h8220000;
      12127: inst = 32'h10408000;
      12128: inst = 32'hc404e1b;
      12129: inst = 32'h8220000;
      12130: inst = 32'h10408000;
      12131: inst = 32'hc404e1c;
      12132: inst = 32'h8220000;
      12133: inst = 32'h10408000;
      12134: inst = 32'hc404e1d;
      12135: inst = 32'h8220000;
      12136: inst = 32'h10408000;
      12137: inst = 32'hc404e1e;
      12138: inst = 32'h8220000;
      12139: inst = 32'h10408000;
      12140: inst = 32'hc404e70;
      12141: inst = 32'h8220000;
      12142: inst = 32'h10408000;
      12143: inst = 32'hc404e71;
      12144: inst = 32'h8220000;
      12145: inst = 32'h10408000;
      12146: inst = 32'hc404e72;
      12147: inst = 32'h8220000;
      12148: inst = 32'h10408000;
      12149: inst = 32'hc404e73;
      12150: inst = 32'h8220000;
      12151: inst = 32'h10408000;
      12152: inst = 32'hc404e74;
      12153: inst = 32'h8220000;
      12154: inst = 32'h10408000;
      12155: inst = 32'hc404e75;
      12156: inst = 32'h8220000;
      12157: inst = 32'h10408000;
      12158: inst = 32'hc404e76;
      12159: inst = 32'h8220000;
      12160: inst = 32'h10408000;
      12161: inst = 32'hc404e77;
      12162: inst = 32'h8220000;
      12163: inst = 32'h10408000;
      12164: inst = 32'hc404e78;
      12165: inst = 32'h8220000;
      12166: inst = 32'h10408000;
      12167: inst = 32'hc404e79;
      12168: inst = 32'h8220000;
      12169: inst = 32'h10408000;
      12170: inst = 32'hc404e7a;
      12171: inst = 32'h8220000;
      12172: inst = 32'h10408000;
      12173: inst = 32'hc404e7b;
      12174: inst = 32'h8220000;
      12175: inst = 32'h10408000;
      12176: inst = 32'hc404e7c;
      12177: inst = 32'h8220000;
      12178: inst = 32'h10408000;
      12179: inst = 32'hc404e7d;
      12180: inst = 32'h8220000;
      12181: inst = 32'h10408000;
      12182: inst = 32'hc404e7e;
      12183: inst = 32'h8220000;
      12184: inst = 32'h10408000;
      12185: inst = 32'hc404ed0;
      12186: inst = 32'h8220000;
      12187: inst = 32'h10408000;
      12188: inst = 32'hc404ed1;
      12189: inst = 32'h8220000;
      12190: inst = 32'h10408000;
      12191: inst = 32'hc404ed2;
      12192: inst = 32'h8220000;
      12193: inst = 32'h10408000;
      12194: inst = 32'hc404ed3;
      12195: inst = 32'h8220000;
      12196: inst = 32'h10408000;
      12197: inst = 32'hc404ed4;
      12198: inst = 32'h8220000;
      12199: inst = 32'h10408000;
      12200: inst = 32'hc404ed5;
      12201: inst = 32'h8220000;
      12202: inst = 32'h10408000;
      12203: inst = 32'hc404ed6;
      12204: inst = 32'h8220000;
      12205: inst = 32'h10408000;
      12206: inst = 32'hc404ed7;
      12207: inst = 32'h8220000;
      12208: inst = 32'h10408000;
      12209: inst = 32'hc404ed8;
      12210: inst = 32'h8220000;
      12211: inst = 32'h10408000;
      12212: inst = 32'hc404ed9;
      12213: inst = 32'h8220000;
      12214: inst = 32'h10408000;
      12215: inst = 32'hc404eda;
      12216: inst = 32'h8220000;
      12217: inst = 32'h10408000;
      12218: inst = 32'hc404edb;
      12219: inst = 32'h8220000;
      12220: inst = 32'h10408000;
      12221: inst = 32'hc404edc;
      12222: inst = 32'h8220000;
      12223: inst = 32'h10408000;
      12224: inst = 32'hc404edd;
      12225: inst = 32'h8220000;
      12226: inst = 32'h10408000;
      12227: inst = 32'hc404ede;
      12228: inst = 32'h8220000;
      12229: inst = 32'h10408000;
      12230: inst = 32'hc404f30;
      12231: inst = 32'h8220000;
      12232: inst = 32'h10408000;
      12233: inst = 32'hc404f31;
      12234: inst = 32'h8220000;
      12235: inst = 32'h10408000;
      12236: inst = 32'hc404f32;
      12237: inst = 32'h8220000;
      12238: inst = 32'h10408000;
      12239: inst = 32'hc404f33;
      12240: inst = 32'h8220000;
      12241: inst = 32'h10408000;
      12242: inst = 32'hc404f34;
      12243: inst = 32'h8220000;
      12244: inst = 32'h10408000;
      12245: inst = 32'hc404f35;
      12246: inst = 32'h8220000;
      12247: inst = 32'h10408000;
      12248: inst = 32'hc404f36;
      12249: inst = 32'h8220000;
      12250: inst = 32'h10408000;
      12251: inst = 32'hc404f37;
      12252: inst = 32'h8220000;
      12253: inst = 32'h10408000;
      12254: inst = 32'hc404f38;
      12255: inst = 32'h8220000;
      12256: inst = 32'h10408000;
      12257: inst = 32'hc404f39;
      12258: inst = 32'h8220000;
      12259: inst = 32'h10408000;
      12260: inst = 32'hc404f3a;
      12261: inst = 32'h8220000;
      12262: inst = 32'h10408000;
      12263: inst = 32'hc404f3b;
      12264: inst = 32'h8220000;
      12265: inst = 32'h10408000;
      12266: inst = 32'hc404f3c;
      12267: inst = 32'h8220000;
      12268: inst = 32'h10408000;
      12269: inst = 32'hc404f3d;
      12270: inst = 32'h8220000;
      12271: inst = 32'h10408000;
      12272: inst = 32'hc404f3e;
      12273: inst = 32'h8220000;
      12274: inst = 32'h10408000;
      12275: inst = 32'hc404f90;
      12276: inst = 32'h8220000;
      12277: inst = 32'h10408000;
      12278: inst = 32'hc404f91;
      12279: inst = 32'h8220000;
      12280: inst = 32'h10408000;
      12281: inst = 32'hc404f92;
      12282: inst = 32'h8220000;
      12283: inst = 32'h10408000;
      12284: inst = 32'hc404f93;
      12285: inst = 32'h8220000;
      12286: inst = 32'h10408000;
      12287: inst = 32'hc404f94;
      12288: inst = 32'h8220000;
      12289: inst = 32'h10408000;
      12290: inst = 32'hc404f95;
      12291: inst = 32'h8220000;
      12292: inst = 32'h10408000;
      12293: inst = 32'hc404f96;
      12294: inst = 32'h8220000;
      12295: inst = 32'h10408000;
      12296: inst = 32'hc404f97;
      12297: inst = 32'h8220000;
      12298: inst = 32'h10408000;
      12299: inst = 32'hc404f98;
      12300: inst = 32'h8220000;
      12301: inst = 32'h10408000;
      12302: inst = 32'hc404f99;
      12303: inst = 32'h8220000;
      12304: inst = 32'h10408000;
      12305: inst = 32'hc404f9a;
      12306: inst = 32'h8220000;
      12307: inst = 32'h10408000;
      12308: inst = 32'hc404f9b;
      12309: inst = 32'h8220000;
      12310: inst = 32'h10408000;
      12311: inst = 32'hc404f9c;
      12312: inst = 32'h8220000;
      12313: inst = 32'h10408000;
      12314: inst = 32'hc404f9d;
      12315: inst = 32'h8220000;
      12316: inst = 32'h10408000;
      12317: inst = 32'hc404f9e;
      12318: inst = 32'h8220000;
      12319: inst = 32'h10408000;
      12320: inst = 32'hc404ff0;
      12321: inst = 32'h8220000;
      12322: inst = 32'h10408000;
      12323: inst = 32'hc404ff1;
      12324: inst = 32'h8220000;
      12325: inst = 32'h10408000;
      12326: inst = 32'hc404ff2;
      12327: inst = 32'h8220000;
      12328: inst = 32'h10408000;
      12329: inst = 32'hc404ff3;
      12330: inst = 32'h8220000;
      12331: inst = 32'h10408000;
      12332: inst = 32'hc404ff4;
      12333: inst = 32'h8220000;
      12334: inst = 32'h10408000;
      12335: inst = 32'hc404ff5;
      12336: inst = 32'h8220000;
      12337: inst = 32'h10408000;
      12338: inst = 32'hc404ff6;
      12339: inst = 32'h8220000;
      12340: inst = 32'h10408000;
      12341: inst = 32'hc404ff7;
      12342: inst = 32'h8220000;
      12343: inst = 32'h10408000;
      12344: inst = 32'hc404ff8;
      12345: inst = 32'h8220000;
      12346: inst = 32'h10408000;
      12347: inst = 32'hc404ff9;
      12348: inst = 32'h8220000;
      12349: inst = 32'h10408000;
      12350: inst = 32'hc404ffa;
      12351: inst = 32'h8220000;
      12352: inst = 32'h10408000;
      12353: inst = 32'hc404ffb;
      12354: inst = 32'h8220000;
      12355: inst = 32'h10408000;
      12356: inst = 32'hc404ffc;
      12357: inst = 32'h8220000;
      12358: inst = 32'h10408000;
      12359: inst = 32'hc404ffd;
      12360: inst = 32'h8220000;
      12361: inst = 32'h10408000;
      12362: inst = 32'hc404ffe;
      12363: inst = 32'h8220000;
      12364: inst = 32'h10408000;
      12365: inst = 32'hc405050;
      12366: inst = 32'h8220000;
      12367: inst = 32'h10408000;
      12368: inst = 32'hc405051;
      12369: inst = 32'h8220000;
      12370: inst = 32'h10408000;
      12371: inst = 32'hc405052;
      12372: inst = 32'h8220000;
      12373: inst = 32'h10408000;
      12374: inst = 32'hc405053;
      12375: inst = 32'h8220000;
      12376: inst = 32'h10408000;
      12377: inst = 32'hc405054;
      12378: inst = 32'h8220000;
      12379: inst = 32'h10408000;
      12380: inst = 32'hc405055;
      12381: inst = 32'h8220000;
      12382: inst = 32'h10408000;
      12383: inst = 32'hc405056;
      12384: inst = 32'h8220000;
      12385: inst = 32'h10408000;
      12386: inst = 32'hc405057;
      12387: inst = 32'h8220000;
      12388: inst = 32'h10408000;
      12389: inst = 32'hc405058;
      12390: inst = 32'h8220000;
      12391: inst = 32'h10408000;
      12392: inst = 32'hc405059;
      12393: inst = 32'h8220000;
      12394: inst = 32'h10408000;
      12395: inst = 32'hc40505a;
      12396: inst = 32'h8220000;
      12397: inst = 32'h10408000;
      12398: inst = 32'hc40505b;
      12399: inst = 32'h8220000;
      12400: inst = 32'h10408000;
      12401: inst = 32'hc40505c;
      12402: inst = 32'h8220000;
      12403: inst = 32'h10408000;
      12404: inst = 32'hc40505d;
      12405: inst = 32'h8220000;
      12406: inst = 32'h10408000;
      12407: inst = 32'hc40505e;
      12408: inst = 32'h8220000;
      12409: inst = 32'h10408000;
      12410: inst = 32'hc4050b0;
      12411: inst = 32'h8220000;
      12412: inst = 32'h10408000;
      12413: inst = 32'hc4050b1;
      12414: inst = 32'h8220000;
      12415: inst = 32'h10408000;
      12416: inst = 32'hc4050b2;
      12417: inst = 32'h8220000;
      12418: inst = 32'h10408000;
      12419: inst = 32'hc4050b3;
      12420: inst = 32'h8220000;
      12421: inst = 32'h10408000;
      12422: inst = 32'hc4050b4;
      12423: inst = 32'h8220000;
      12424: inst = 32'h10408000;
      12425: inst = 32'hc4050b5;
      12426: inst = 32'h8220000;
      12427: inst = 32'h10408000;
      12428: inst = 32'hc4050b6;
      12429: inst = 32'h8220000;
      12430: inst = 32'h10408000;
      12431: inst = 32'hc4050b7;
      12432: inst = 32'h8220000;
      12433: inst = 32'h10408000;
      12434: inst = 32'hc4050b8;
      12435: inst = 32'h8220000;
      12436: inst = 32'h10408000;
      12437: inst = 32'hc4050b9;
      12438: inst = 32'h8220000;
      12439: inst = 32'h10408000;
      12440: inst = 32'hc4050ba;
      12441: inst = 32'h8220000;
      12442: inst = 32'h10408000;
      12443: inst = 32'hc4050bb;
      12444: inst = 32'h8220000;
      12445: inst = 32'h10408000;
      12446: inst = 32'hc4050bc;
      12447: inst = 32'h8220000;
      12448: inst = 32'h10408000;
      12449: inst = 32'hc4050bd;
      12450: inst = 32'h8220000;
      12451: inst = 32'h10408000;
      12452: inst = 32'hc4050be;
      12453: inst = 32'h8220000;
      12454: inst = 32'h10408000;
      12455: inst = 32'hc405110;
      12456: inst = 32'h8220000;
      12457: inst = 32'h10408000;
      12458: inst = 32'hc405111;
      12459: inst = 32'h8220000;
      12460: inst = 32'h10408000;
      12461: inst = 32'hc405112;
      12462: inst = 32'h8220000;
      12463: inst = 32'h10408000;
      12464: inst = 32'hc405113;
      12465: inst = 32'h8220000;
      12466: inst = 32'h10408000;
      12467: inst = 32'hc405114;
      12468: inst = 32'h8220000;
      12469: inst = 32'h10408000;
      12470: inst = 32'hc405115;
      12471: inst = 32'h8220000;
      12472: inst = 32'h10408000;
      12473: inst = 32'hc405116;
      12474: inst = 32'h8220000;
      12475: inst = 32'h10408000;
      12476: inst = 32'hc405117;
      12477: inst = 32'h8220000;
      12478: inst = 32'h10408000;
      12479: inst = 32'hc405118;
      12480: inst = 32'h8220000;
      12481: inst = 32'h10408000;
      12482: inst = 32'hc405119;
      12483: inst = 32'h8220000;
      12484: inst = 32'h10408000;
      12485: inst = 32'hc40511a;
      12486: inst = 32'h8220000;
      12487: inst = 32'h10408000;
      12488: inst = 32'hc40511b;
      12489: inst = 32'h8220000;
      12490: inst = 32'h10408000;
      12491: inst = 32'hc40511c;
      12492: inst = 32'h8220000;
      12493: inst = 32'h10408000;
      12494: inst = 32'hc40511d;
      12495: inst = 32'h8220000;
      12496: inst = 32'h10408000;
      12497: inst = 32'hc40511e;
      12498: inst = 32'h8220000;
      12499: inst = 32'h10408000;
      12500: inst = 32'hc405170;
      12501: inst = 32'h8220000;
      12502: inst = 32'h10408000;
      12503: inst = 32'hc405171;
      12504: inst = 32'h8220000;
      12505: inst = 32'h10408000;
      12506: inst = 32'hc405172;
      12507: inst = 32'h8220000;
      12508: inst = 32'h10408000;
      12509: inst = 32'hc405173;
      12510: inst = 32'h8220000;
      12511: inst = 32'h10408000;
      12512: inst = 32'hc405174;
      12513: inst = 32'h8220000;
      12514: inst = 32'h10408000;
      12515: inst = 32'hc405175;
      12516: inst = 32'h8220000;
      12517: inst = 32'h10408000;
      12518: inst = 32'hc405176;
      12519: inst = 32'h8220000;
      12520: inst = 32'h10408000;
      12521: inst = 32'hc405177;
      12522: inst = 32'h8220000;
      12523: inst = 32'h10408000;
      12524: inst = 32'hc405178;
      12525: inst = 32'h8220000;
      12526: inst = 32'h10408000;
      12527: inst = 32'hc405179;
      12528: inst = 32'h8220000;
      12529: inst = 32'h10408000;
      12530: inst = 32'hc40517a;
      12531: inst = 32'h8220000;
      12532: inst = 32'h10408000;
      12533: inst = 32'hc40517b;
      12534: inst = 32'h8220000;
      12535: inst = 32'h10408000;
      12536: inst = 32'hc40517c;
      12537: inst = 32'h8220000;
      12538: inst = 32'h10408000;
      12539: inst = 32'hc40517d;
      12540: inst = 32'h8220000;
      12541: inst = 32'h10408000;
      12542: inst = 32'hc40517e;
      12543: inst = 32'h8220000;
      12544: inst = 32'h10408000;
      12545: inst = 32'hc4051d0;
      12546: inst = 32'h8220000;
      12547: inst = 32'h10408000;
      12548: inst = 32'hc4051d1;
      12549: inst = 32'h8220000;
      12550: inst = 32'h10408000;
      12551: inst = 32'hc4051d2;
      12552: inst = 32'h8220000;
      12553: inst = 32'h10408000;
      12554: inst = 32'hc4051d3;
      12555: inst = 32'h8220000;
      12556: inst = 32'h10408000;
      12557: inst = 32'hc4051d4;
      12558: inst = 32'h8220000;
      12559: inst = 32'h10408000;
      12560: inst = 32'hc4051d5;
      12561: inst = 32'h8220000;
      12562: inst = 32'h10408000;
      12563: inst = 32'hc4051d6;
      12564: inst = 32'h8220000;
      12565: inst = 32'h10408000;
      12566: inst = 32'hc4051d7;
      12567: inst = 32'h8220000;
      12568: inst = 32'h10408000;
      12569: inst = 32'hc4051d8;
      12570: inst = 32'h8220000;
      12571: inst = 32'h10408000;
      12572: inst = 32'hc4051d9;
      12573: inst = 32'h8220000;
      12574: inst = 32'h10408000;
      12575: inst = 32'hc4051da;
      12576: inst = 32'h8220000;
      12577: inst = 32'h10408000;
      12578: inst = 32'hc4051db;
      12579: inst = 32'h8220000;
      12580: inst = 32'h10408000;
      12581: inst = 32'hc4051dc;
      12582: inst = 32'h8220000;
      12583: inst = 32'h10408000;
      12584: inst = 32'hc4051dd;
      12585: inst = 32'h8220000;
      12586: inst = 32'h10408000;
      12587: inst = 32'hc4051de;
      12588: inst = 32'h8220000;
      12589: inst = 32'h10408000;
      12590: inst = 32'hc405230;
      12591: inst = 32'h8220000;
      12592: inst = 32'h10408000;
      12593: inst = 32'hc405231;
      12594: inst = 32'h8220000;
      12595: inst = 32'h10408000;
      12596: inst = 32'hc405232;
      12597: inst = 32'h8220000;
      12598: inst = 32'h10408000;
      12599: inst = 32'hc405233;
      12600: inst = 32'h8220000;
      12601: inst = 32'h10408000;
      12602: inst = 32'hc405234;
      12603: inst = 32'h8220000;
      12604: inst = 32'h10408000;
      12605: inst = 32'hc405235;
      12606: inst = 32'h8220000;
      12607: inst = 32'h10408000;
      12608: inst = 32'hc405236;
      12609: inst = 32'h8220000;
      12610: inst = 32'h10408000;
      12611: inst = 32'hc405237;
      12612: inst = 32'h8220000;
      12613: inst = 32'h10408000;
      12614: inst = 32'hc405238;
      12615: inst = 32'h8220000;
      12616: inst = 32'h10408000;
      12617: inst = 32'hc405239;
      12618: inst = 32'h8220000;
      12619: inst = 32'h10408000;
      12620: inst = 32'hc40523a;
      12621: inst = 32'h8220000;
      12622: inst = 32'h10408000;
      12623: inst = 32'hc40523b;
      12624: inst = 32'h8220000;
      12625: inst = 32'h10408000;
      12626: inst = 32'hc40523c;
      12627: inst = 32'h8220000;
      12628: inst = 32'h10408000;
      12629: inst = 32'hc40523d;
      12630: inst = 32'h8220000;
      12631: inst = 32'h10408000;
      12632: inst = 32'hc40523e;
      12633: inst = 32'h8220000;
      12634: inst = 32'h10408000;
      12635: inst = 32'hc405290;
      12636: inst = 32'h8220000;
      12637: inst = 32'h10408000;
      12638: inst = 32'hc405291;
      12639: inst = 32'h8220000;
      12640: inst = 32'h10408000;
      12641: inst = 32'hc405292;
      12642: inst = 32'h8220000;
      12643: inst = 32'h10408000;
      12644: inst = 32'hc405293;
      12645: inst = 32'h8220000;
      12646: inst = 32'h10408000;
      12647: inst = 32'hc405294;
      12648: inst = 32'h8220000;
      12649: inst = 32'h10408000;
      12650: inst = 32'hc405295;
      12651: inst = 32'h8220000;
      12652: inst = 32'h10408000;
      12653: inst = 32'hc405296;
      12654: inst = 32'h8220000;
      12655: inst = 32'h10408000;
      12656: inst = 32'hc405297;
      12657: inst = 32'h8220000;
      12658: inst = 32'h10408000;
      12659: inst = 32'hc405298;
      12660: inst = 32'h8220000;
      12661: inst = 32'h10408000;
      12662: inst = 32'hc405299;
      12663: inst = 32'h8220000;
      12664: inst = 32'h10408000;
      12665: inst = 32'hc40529a;
      12666: inst = 32'h8220000;
      12667: inst = 32'h10408000;
      12668: inst = 32'hc40529b;
      12669: inst = 32'h8220000;
      12670: inst = 32'h10408000;
      12671: inst = 32'hc40529c;
      12672: inst = 32'h8220000;
      12673: inst = 32'h10408000;
      12674: inst = 32'hc40529d;
      12675: inst = 32'h8220000;
      12676: inst = 32'h10408000;
      12677: inst = 32'hc40529e;
      12678: inst = 32'h8220000;
      12679: inst = 32'hc20ef7c;
      12680: inst = 32'h10408000;
      12681: inst = 32'hc404932;
      12682: inst = 32'h8220000;
      12683: inst = 32'h10408000;
      12684: inst = 32'hc404933;
      12685: inst = 32'h8220000;
      12686: inst = 32'h10408000;
      12687: inst = 32'hc404934;
      12688: inst = 32'h8220000;
      12689: inst = 32'h10408000;
      12690: inst = 32'hc404935;
      12691: inst = 32'h8220000;
      12692: inst = 32'h10408000;
      12693: inst = 32'hc404993;
      12694: inst = 32'h8220000;
      12695: inst = 32'h10408000;
      12696: inst = 32'hc404994;
      12697: inst = 32'h8220000;
      12698: inst = 32'h10408000;
      12699: inst = 32'hc404995;
      12700: inst = 32'h8220000;
      12701: inst = 32'h10408000;
      12702: inst = 32'hc4049f3;
      12703: inst = 32'h8220000;
      12704: inst = 32'h10408000;
      12705: inst = 32'hc4049f4;
      12706: inst = 32'h8220000;
      12707: inst = 32'h10408000;
      12708: inst = 32'hc4049f5;
      12709: inst = 32'h8220000;
      12710: inst = 32'h10408000;
      12711: inst = 32'hc404a53;
      12712: inst = 32'h8220000;
      12713: inst = 32'h10408000;
      12714: inst = 32'hc404a54;
      12715: inst = 32'h8220000;
      12716: inst = 32'h10408000;
      12717: inst = 32'hc404a55;
      12718: inst = 32'h8220000;
      12719: inst = 32'h10408000;
      12720: inst = 32'hc404ab2;
      12721: inst = 32'h8220000;
      12722: inst = 32'h10408000;
      12723: inst = 32'hc404ab3;
      12724: inst = 32'h8220000;
      12725: inst = 32'h10408000;
      12726: inst = 32'hc404ab5;
      12727: inst = 32'h8220000;
      12728: inst = 32'h10408000;
      12729: inst = 32'hc404b12;
      12730: inst = 32'h8220000;
      12731: inst = 32'h10408000;
      12732: inst = 32'hc404b13;
      12733: inst = 32'h8220000;
      12734: inst = 32'h10408000;
      12735: inst = 32'hc404b15;
      12736: inst = 32'h8220000;
      12737: inst = 32'h10408000;
      12738: inst = 32'hc404b72;
      12739: inst = 32'h8220000;
      12740: inst = 32'h10408000;
      12741: inst = 32'hc404b73;
      12742: inst = 32'h8220000;
      12743: inst = 32'h10408000;
      12744: inst = 32'hc404b74;
      12745: inst = 32'h8220000;
      12746: inst = 32'h10408000;
      12747: inst = 32'hc404b75;
      12748: inst = 32'h8220000;
      12749: inst = 32'hc20eed7;
      12750: inst = 32'h10408000;
      12751: inst = 32'hc404a08;
      12752: inst = 32'h8220000;
      12753: inst = 32'h10408000;
      12754: inst = 32'hc404a0e;
      12755: inst = 32'h8220000;
      12756: inst = 32'hc20e6fa;
      12757: inst = 32'h10408000;
      12758: inst = 32'hc404a09;
      12759: inst = 32'h8220000;
      12760: inst = 32'h10408000;
      12761: inst = 32'hc404a0d;
      12762: inst = 32'h8220000;
      12763: inst = 32'h10408000;
      12764: inst = 32'hc404be7;
      12765: inst = 32'h8220000;
      12766: inst = 32'hc20e6fb;
      12767: inst = 32'h10408000;
      12768: inst = 32'hc404a0a;
      12769: inst = 32'h8220000;
      12770: inst = 32'h10408000;
      12771: inst = 32'hc404a0c;
      12772: inst = 32'h8220000;
      12773: inst = 32'h10408000;
      12774: inst = 32'hc404ac7;
      12775: inst = 32'h8220000;
      12776: inst = 32'h10408000;
      12777: inst = 32'hc404acf;
      12778: inst = 32'h8220000;
      12779: inst = 32'h10408000;
      12780: inst = 32'hc404b87;
      12781: inst = 32'h8220000;
      12782: inst = 32'h10408000;
      12783: inst = 32'hc404b8f;
      12784: inst = 32'h8220000;
      12785: inst = 32'h10408000;
      12786: inst = 32'hc404c4d;
      12787: inst = 32'h8220000;
      12788: inst = 32'hc20defb;
      12789: inst = 32'h10408000;
      12790: inst = 32'hc404a0b;
      12791: inst = 32'h8220000;
      12792: inst = 32'h10408000;
      12793: inst = 32'hc404a68;
      12794: inst = 32'h8220000;
      12795: inst = 32'h10408000;
      12796: inst = 32'hc404a69;
      12797: inst = 32'h8220000;
      12798: inst = 32'h10408000;
      12799: inst = 32'hc404a6a;
      12800: inst = 32'h8220000;
      12801: inst = 32'h10408000;
      12802: inst = 32'hc404a6b;
      12803: inst = 32'h8220000;
      12804: inst = 32'h10408000;
      12805: inst = 32'hc404a6c;
      12806: inst = 32'h8220000;
      12807: inst = 32'h10408000;
      12808: inst = 32'hc404a6d;
      12809: inst = 32'h8220000;
      12810: inst = 32'h10408000;
      12811: inst = 32'hc404a6e;
      12812: inst = 32'h8220000;
      12813: inst = 32'h10408000;
      12814: inst = 32'hc404ac8;
      12815: inst = 32'h8220000;
      12816: inst = 32'h10408000;
      12817: inst = 32'hc404ac9;
      12818: inst = 32'h8220000;
      12819: inst = 32'h10408000;
      12820: inst = 32'hc404aca;
      12821: inst = 32'h8220000;
      12822: inst = 32'h10408000;
      12823: inst = 32'hc404acb;
      12824: inst = 32'h8220000;
      12825: inst = 32'h10408000;
      12826: inst = 32'hc404acc;
      12827: inst = 32'h8220000;
      12828: inst = 32'h10408000;
      12829: inst = 32'hc404acd;
      12830: inst = 32'h8220000;
      12831: inst = 32'h10408000;
      12832: inst = 32'hc404ace;
      12833: inst = 32'h8220000;
      12834: inst = 32'h10408000;
      12835: inst = 32'hc404b27;
      12836: inst = 32'h8220000;
      12837: inst = 32'h10408000;
      12838: inst = 32'hc404b2a;
      12839: inst = 32'h8220000;
      12840: inst = 32'h10408000;
      12841: inst = 32'hc404b2d;
      12842: inst = 32'h8220000;
      12843: inst = 32'h10408000;
      12844: inst = 32'hc404b2e;
      12845: inst = 32'h8220000;
      12846: inst = 32'h10408000;
      12847: inst = 32'hc404b2f;
      12848: inst = 32'h8220000;
      12849: inst = 32'h10408000;
      12850: inst = 32'hc404b8a;
      12851: inst = 32'h8220000;
      12852: inst = 32'h10408000;
      12853: inst = 32'hc404b8d;
      12854: inst = 32'h8220000;
      12855: inst = 32'h10408000;
      12856: inst = 32'hc404b8e;
      12857: inst = 32'h8220000;
      12858: inst = 32'h10408000;
      12859: inst = 32'hc404be8;
      12860: inst = 32'h8220000;
      12861: inst = 32'h10408000;
      12862: inst = 32'hc404be9;
      12863: inst = 32'h8220000;
      12864: inst = 32'h10408000;
      12865: inst = 32'hc404bea;
      12866: inst = 32'h8220000;
      12867: inst = 32'h10408000;
      12868: inst = 32'hc404beb;
      12869: inst = 32'h8220000;
      12870: inst = 32'h10408000;
      12871: inst = 32'hc404bec;
      12872: inst = 32'h8220000;
      12873: inst = 32'h10408000;
      12874: inst = 32'hc404bed;
      12875: inst = 32'h8220000;
      12876: inst = 32'h10408000;
      12877: inst = 32'hc404bee;
      12878: inst = 32'h8220000;
      12879: inst = 32'h10408000;
      12880: inst = 32'hc404c49;
      12881: inst = 32'h8220000;
      12882: inst = 32'h10408000;
      12883: inst = 32'hc404c4b;
      12884: inst = 32'h8220000;
      12885: inst = 32'h10408000;
      12886: inst = 32'hc404ca9;
      12887: inst = 32'h8220000;
      12888: inst = 32'h10408000;
      12889: inst = 32'hc404cab;
      12890: inst = 32'h8220000;
      12891: inst = 32'hc20eed8;
      12892: inst = 32'h10408000;
      12893: inst = 32'hc404a67;
      12894: inst = 32'h8220000;
      12895: inst = 32'h10408000;
      12896: inst = 32'hc404a6f;
      12897: inst = 32'h8220000;
      12898: inst = 32'hc204a69;
      12899: inst = 32'h10408000;
      12900: inst = 32'hc404b28;
      12901: inst = 32'h8220000;
      12902: inst = 32'h10408000;
      12903: inst = 32'hc404b29;
      12904: inst = 32'h8220000;
      12905: inst = 32'h10408000;
      12906: inst = 32'hc404b2b;
      12907: inst = 32'h8220000;
      12908: inst = 32'h10408000;
      12909: inst = 32'hc404b2c;
      12910: inst = 32'h8220000;
      12911: inst = 32'h10408000;
      12912: inst = 32'hc404b88;
      12913: inst = 32'h8220000;
      12914: inst = 32'h10408000;
      12915: inst = 32'hc404b89;
      12916: inst = 32'h8220000;
      12917: inst = 32'h10408000;
      12918: inst = 32'hc404b8b;
      12919: inst = 32'h8220000;
      12920: inst = 32'h10408000;
      12921: inst = 32'hc404b8c;
      12922: inst = 32'h8220000;
      12923: inst = 32'h10408000;
      12924: inst = 32'hc404c48;
      12925: inst = 32'h8220000;
      12926: inst = 32'h10408000;
      12927: inst = 32'hc404c4a;
      12928: inst = 32'h8220000;
      12929: inst = 32'h10408000;
      12930: inst = 32'hc404c4c;
      12931: inst = 32'h8220000;
      12932: inst = 32'h10408000;
      12933: inst = 32'hc404ca8;
      12934: inst = 32'h8220000;
      12935: inst = 32'h10408000;
      12936: inst = 32'hc404caa;
      12937: inst = 32'h8220000;
      12938: inst = 32'h10408000;
      12939: inst = 32'hc404cac;
      12940: inst = 32'h8220000;
      12941: inst = 32'h10408000;
      12942: inst = 32'hc405085;
      12943: inst = 32'h8220000;
      12944: inst = 32'h10408000;
      12945: inst = 32'hc40509a;
      12946: inst = 32'h8220000;
      12947: inst = 32'h10408000;
      12948: inst = 32'hc4050e4;
      12949: inst = 32'h8220000;
      12950: inst = 32'h10408000;
      12951: inst = 32'hc4050e5;
      12952: inst = 32'h8220000;
      12953: inst = 32'h10408000;
      12954: inst = 32'hc4050fa;
      12955: inst = 32'h8220000;
      12956: inst = 32'h10408000;
      12957: inst = 32'hc4050fb;
      12958: inst = 32'h8220000;
      12959: inst = 32'h10408000;
      12960: inst = 32'hc405143;
      12961: inst = 32'h8220000;
      12962: inst = 32'h10408000;
      12963: inst = 32'hc405144;
      12964: inst = 32'h8220000;
      12965: inst = 32'h10408000;
      12966: inst = 32'hc405145;
      12967: inst = 32'h8220000;
      12968: inst = 32'h10408000;
      12969: inst = 32'hc40515a;
      12970: inst = 32'h8220000;
      12971: inst = 32'h10408000;
      12972: inst = 32'hc40515b;
      12973: inst = 32'h8220000;
      12974: inst = 32'h10408000;
      12975: inst = 32'hc40515c;
      12976: inst = 32'h8220000;
      12977: inst = 32'h10408000;
      12978: inst = 32'hc4051a2;
      12979: inst = 32'h8220000;
      12980: inst = 32'h10408000;
      12981: inst = 32'hc4051a3;
      12982: inst = 32'h8220000;
      12983: inst = 32'h10408000;
      12984: inst = 32'hc4051a4;
      12985: inst = 32'h8220000;
      12986: inst = 32'h10408000;
      12987: inst = 32'hc4051a5;
      12988: inst = 32'h8220000;
      12989: inst = 32'h10408000;
      12990: inst = 32'hc4051ba;
      12991: inst = 32'h8220000;
      12992: inst = 32'h10408000;
      12993: inst = 32'hc4051bb;
      12994: inst = 32'h8220000;
      12995: inst = 32'h10408000;
      12996: inst = 32'hc4051bc;
      12997: inst = 32'h8220000;
      12998: inst = 32'h10408000;
      12999: inst = 32'hc4051bd;
      13000: inst = 32'h8220000;
      13001: inst = 32'h10408000;
      13002: inst = 32'hc405202;
      13003: inst = 32'h8220000;
      13004: inst = 32'h10408000;
      13005: inst = 32'hc405203;
      13006: inst = 32'h8220000;
      13007: inst = 32'h10408000;
      13008: inst = 32'hc405204;
      13009: inst = 32'h8220000;
      13010: inst = 32'h10408000;
      13011: inst = 32'hc405205;
      13012: inst = 32'h8220000;
      13013: inst = 32'h10408000;
      13014: inst = 32'hc40521a;
      13015: inst = 32'h8220000;
      13016: inst = 32'h10408000;
      13017: inst = 32'hc40521b;
      13018: inst = 32'h8220000;
      13019: inst = 32'h10408000;
      13020: inst = 32'hc40521c;
      13021: inst = 32'h8220000;
      13022: inst = 32'h10408000;
      13023: inst = 32'hc40521d;
      13024: inst = 32'h8220000;
      13025: inst = 32'h10408000;
      13026: inst = 32'hc405262;
      13027: inst = 32'h8220000;
      13028: inst = 32'h10408000;
      13029: inst = 32'hc405263;
      13030: inst = 32'h8220000;
      13031: inst = 32'h10408000;
      13032: inst = 32'hc405264;
      13033: inst = 32'h8220000;
      13034: inst = 32'h10408000;
      13035: inst = 32'hc405265;
      13036: inst = 32'h8220000;
      13037: inst = 32'h10408000;
      13038: inst = 32'hc40527a;
      13039: inst = 32'h8220000;
      13040: inst = 32'h10408000;
      13041: inst = 32'hc40527b;
      13042: inst = 32'h8220000;
      13043: inst = 32'h10408000;
      13044: inst = 32'hc40527c;
      13045: inst = 32'h8220000;
      13046: inst = 32'h10408000;
      13047: inst = 32'hc40527d;
      13048: inst = 32'h8220000;
      13049: inst = 32'h10408000;
      13050: inst = 32'hc4052c2;
      13051: inst = 32'h8220000;
      13052: inst = 32'h10408000;
      13053: inst = 32'hc4052c3;
      13054: inst = 32'h8220000;
      13055: inst = 32'h10408000;
      13056: inst = 32'hc4052c4;
      13057: inst = 32'h8220000;
      13058: inst = 32'h10408000;
      13059: inst = 32'hc4052db;
      13060: inst = 32'h8220000;
      13061: inst = 32'h10408000;
      13062: inst = 32'hc4052dc;
      13063: inst = 32'h8220000;
      13064: inst = 32'h10408000;
      13065: inst = 32'hc4052dd;
      13066: inst = 32'h8220000;
      13067: inst = 32'h10408000;
      13068: inst = 32'hc405322;
      13069: inst = 32'h8220000;
      13070: inst = 32'h10408000;
      13071: inst = 32'hc405323;
      13072: inst = 32'h8220000;
      13073: inst = 32'h10408000;
      13074: inst = 32'hc405324;
      13075: inst = 32'h8220000;
      13076: inst = 32'h10408000;
      13077: inst = 32'hc40533b;
      13078: inst = 32'h8220000;
      13079: inst = 32'h10408000;
      13080: inst = 32'hc40533c;
      13081: inst = 32'h8220000;
      13082: inst = 32'h10408000;
      13083: inst = 32'hc40533d;
      13084: inst = 32'h8220000;
      13085: inst = 32'h10408000;
      13086: inst = 32'hc40537f;
      13087: inst = 32'h8220000;
      13088: inst = 32'h10408000;
      13089: inst = 32'hc405382;
      13090: inst = 32'h8220000;
      13091: inst = 32'h10408000;
      13092: inst = 32'hc405383;
      13093: inst = 32'h8220000;
      13094: inst = 32'h10408000;
      13095: inst = 32'hc405384;
      13096: inst = 32'h8220000;
      13097: inst = 32'h10408000;
      13098: inst = 32'hc40539b;
      13099: inst = 32'h8220000;
      13100: inst = 32'h10408000;
      13101: inst = 32'hc40539c;
      13102: inst = 32'h8220000;
      13103: inst = 32'h10408000;
      13104: inst = 32'hc40539d;
      13105: inst = 32'h8220000;
      13106: inst = 32'h10408000;
      13107: inst = 32'hc4053a0;
      13108: inst = 32'h8220000;
      13109: inst = 32'h10408000;
      13110: inst = 32'hc4053de;
      13111: inst = 32'h8220000;
      13112: inst = 32'h10408000;
      13113: inst = 32'hc4053df;
      13114: inst = 32'h8220000;
      13115: inst = 32'h10408000;
      13116: inst = 32'hc4053e2;
      13117: inst = 32'h8220000;
      13118: inst = 32'h10408000;
      13119: inst = 32'hc4053e3;
      13120: inst = 32'h8220000;
      13121: inst = 32'h10408000;
      13122: inst = 32'hc4053fc;
      13123: inst = 32'h8220000;
      13124: inst = 32'h10408000;
      13125: inst = 32'hc4053fd;
      13126: inst = 32'h8220000;
      13127: inst = 32'h10408000;
      13128: inst = 32'hc405400;
      13129: inst = 32'h8220000;
      13130: inst = 32'h10408000;
      13131: inst = 32'hc405401;
      13132: inst = 32'h8220000;
      13133: inst = 32'h10408000;
      13134: inst = 32'hc40543d;
      13135: inst = 32'h8220000;
      13136: inst = 32'h10408000;
      13137: inst = 32'hc40543e;
      13138: inst = 32'h8220000;
      13139: inst = 32'h10408000;
      13140: inst = 32'hc40543f;
      13141: inst = 32'h8220000;
      13142: inst = 32'h10408000;
      13143: inst = 32'hc405442;
      13144: inst = 32'h8220000;
      13145: inst = 32'h10408000;
      13146: inst = 32'hc405443;
      13147: inst = 32'h8220000;
      13148: inst = 32'h10408000;
      13149: inst = 32'hc40545c;
      13150: inst = 32'h8220000;
      13151: inst = 32'h10408000;
      13152: inst = 32'hc40545d;
      13153: inst = 32'h8220000;
      13154: inst = 32'h10408000;
      13155: inst = 32'hc405460;
      13156: inst = 32'h8220000;
      13157: inst = 32'h10408000;
      13158: inst = 32'hc405461;
      13159: inst = 32'h8220000;
      13160: inst = 32'h10408000;
      13161: inst = 32'hc405462;
      13162: inst = 32'h8220000;
      13163: inst = 32'h10408000;
      13164: inst = 32'hc40549d;
      13165: inst = 32'h8220000;
      13166: inst = 32'h10408000;
      13167: inst = 32'hc40549e;
      13168: inst = 32'h8220000;
      13169: inst = 32'h10408000;
      13170: inst = 32'hc4054a0;
      13171: inst = 32'h8220000;
      13172: inst = 32'h10408000;
      13173: inst = 32'hc4054a1;
      13174: inst = 32'h8220000;
      13175: inst = 32'h10408000;
      13176: inst = 32'hc4054a2;
      13177: inst = 32'h8220000;
      13178: inst = 32'h10408000;
      13179: inst = 32'hc4054a3;
      13180: inst = 32'h8220000;
      13181: inst = 32'h10408000;
      13182: inst = 32'hc4054bc;
      13183: inst = 32'h8220000;
      13184: inst = 32'h10408000;
      13185: inst = 32'hc4054bd;
      13186: inst = 32'h8220000;
      13187: inst = 32'h10408000;
      13188: inst = 32'hc4054be;
      13189: inst = 32'h8220000;
      13190: inst = 32'h10408000;
      13191: inst = 32'hc4054bf;
      13192: inst = 32'h8220000;
      13193: inst = 32'h10408000;
      13194: inst = 32'hc4054c1;
      13195: inst = 32'h8220000;
      13196: inst = 32'h10408000;
      13197: inst = 32'hc4054c2;
      13198: inst = 32'h8220000;
      13199: inst = 32'h10408000;
      13200: inst = 32'hc4054fc;
      13201: inst = 32'h8220000;
      13202: inst = 32'h10408000;
      13203: inst = 32'hc4054fd;
      13204: inst = 32'h8220000;
      13205: inst = 32'h10408000;
      13206: inst = 32'hc4054fe;
      13207: inst = 32'h8220000;
      13208: inst = 32'h10408000;
      13209: inst = 32'hc405502;
      13210: inst = 32'h8220000;
      13211: inst = 32'h10408000;
      13212: inst = 32'hc40551d;
      13213: inst = 32'h8220000;
      13214: inst = 32'h10408000;
      13215: inst = 32'hc405521;
      13216: inst = 32'h8220000;
      13217: inst = 32'h10408000;
      13218: inst = 32'hc405522;
      13219: inst = 32'h8220000;
      13220: inst = 32'h10408000;
      13221: inst = 32'hc405523;
      13222: inst = 32'h8220000;
      13223: inst = 32'h10408000;
      13224: inst = 32'hc40555b;
      13225: inst = 32'h8220000;
      13226: inst = 32'h10408000;
      13227: inst = 32'hc40555c;
      13228: inst = 32'h8220000;
      13229: inst = 32'h10408000;
      13230: inst = 32'hc40555d;
      13231: inst = 32'h8220000;
      13232: inst = 32'h10408000;
      13233: inst = 32'hc405562;
      13234: inst = 32'h8220000;
      13235: inst = 32'h10408000;
      13236: inst = 32'hc40557d;
      13237: inst = 32'h8220000;
      13238: inst = 32'h10408000;
      13239: inst = 32'hc405582;
      13240: inst = 32'h8220000;
      13241: inst = 32'h10408000;
      13242: inst = 32'hc405583;
      13243: inst = 32'h8220000;
      13244: inst = 32'h10408000;
      13245: inst = 32'hc405584;
      13246: inst = 32'h8220000;
      13247: inst = 32'h10408000;
      13248: inst = 32'hc4055ba;
      13249: inst = 32'h8220000;
      13250: inst = 32'h10408000;
      13251: inst = 32'hc4055bb;
      13252: inst = 32'h8220000;
      13253: inst = 32'h10408000;
      13254: inst = 32'hc4055bc;
      13255: inst = 32'h8220000;
      13256: inst = 32'h10408000;
      13257: inst = 32'hc4055bd;
      13258: inst = 32'h8220000;
      13259: inst = 32'h10408000;
      13260: inst = 32'hc4055c2;
      13261: inst = 32'h8220000;
      13262: inst = 32'h10408000;
      13263: inst = 32'hc4055dd;
      13264: inst = 32'h8220000;
      13265: inst = 32'h10408000;
      13266: inst = 32'hc4055e2;
      13267: inst = 32'h8220000;
      13268: inst = 32'h10408000;
      13269: inst = 32'hc4055e3;
      13270: inst = 32'h8220000;
      13271: inst = 32'h10408000;
      13272: inst = 32'hc4055e4;
      13273: inst = 32'h8220000;
      13274: inst = 32'h10408000;
      13275: inst = 32'hc4055e5;
      13276: inst = 32'h8220000;
      13277: inst = 32'h10408000;
      13278: inst = 32'hc40561a;
      13279: inst = 32'h8220000;
      13280: inst = 32'h10408000;
      13281: inst = 32'hc40561b;
      13282: inst = 32'h8220000;
      13283: inst = 32'h10408000;
      13284: inst = 32'hc40561c;
      13285: inst = 32'h8220000;
      13286: inst = 32'h10408000;
      13287: inst = 32'hc40561d;
      13288: inst = 32'h8220000;
      13289: inst = 32'h10408000;
      13290: inst = 32'hc405642;
      13291: inst = 32'h8220000;
      13292: inst = 32'h10408000;
      13293: inst = 32'hc405643;
      13294: inst = 32'h8220000;
      13295: inst = 32'h10408000;
      13296: inst = 32'hc405644;
      13297: inst = 32'h8220000;
      13298: inst = 32'h10408000;
      13299: inst = 32'hc405645;
      13300: inst = 32'h8220000;
      13301: inst = 32'h10408000;
      13302: inst = 32'hc405679;
      13303: inst = 32'h8220000;
      13304: inst = 32'h10408000;
      13305: inst = 32'hc40567a;
      13306: inst = 32'h8220000;
      13307: inst = 32'h10408000;
      13308: inst = 32'hc40567b;
      13309: inst = 32'h8220000;
      13310: inst = 32'h10408000;
      13311: inst = 32'hc40567c;
      13312: inst = 32'h8220000;
      13313: inst = 32'h10408000;
      13314: inst = 32'hc4056a3;
      13315: inst = 32'h8220000;
      13316: inst = 32'h10408000;
      13317: inst = 32'hc4056a4;
      13318: inst = 32'h8220000;
      13319: inst = 32'h10408000;
      13320: inst = 32'hc4056a5;
      13321: inst = 32'h8220000;
      13322: inst = 32'h10408000;
      13323: inst = 32'hc4056a6;
      13324: inst = 32'h8220000;
      13325: inst = 32'hc20e6d9;
      13326: inst = 32'h10408000;
      13327: inst = 32'hc404bef;
      13328: inst = 32'h8220000;
      13329: inst = 32'h10408000;
      13330: inst = 32'hc404c4e;
      13331: inst = 32'h8220000;
      13332: inst = 32'hc20eeb7;
      13333: inst = 32'h10408000;
      13334: inst = 32'hc404c47;
      13335: inst = 32'h8220000;
      13336: inst = 32'hc20d615;
      13337: inst = 32'h10408000;
      13338: inst = 32'hc404ca2;
      13339: inst = 32'h8220000;
      13340: inst = 32'h10408000;
      13341: inst = 32'hc404d00;
      13342: inst = 32'h8220000;
      13343: inst = 32'hc209c91;
      13344: inst = 32'h10408000;
      13345: inst = 32'hc404ca3;
      13346: inst = 32'h8220000;
      13347: inst = 32'h10408000;
      13348: inst = 32'hc404d01;
      13349: inst = 32'h8220000;
      13350: inst = 32'hc207bf0;
      13351: inst = 32'h10408000;
      13352: inst = 32'hc404ca4;
      13353: inst = 32'h8220000;
      13354: inst = 32'h10408000;
      13355: inst = 32'hc404ca5;
      13356: inst = 32'h8220000;
      13357: inst = 32'h10408000;
      13358: inst = 32'hc404ca6;
      13359: inst = 32'h8220000;
      13360: inst = 32'h10408000;
      13361: inst = 32'hc404ca7;
      13362: inst = 32'h8220000;
      13363: inst = 32'h10408000;
      13364: inst = 32'hc404d02;
      13365: inst = 32'h8220000;
      13366: inst = 32'h10408000;
      13367: inst = 32'hc404d03;
      13368: inst = 32'h8220000;
      13369: inst = 32'h10408000;
      13370: inst = 32'hc404d04;
      13371: inst = 32'h8220000;
      13372: inst = 32'h10408000;
      13373: inst = 32'hc404d05;
      13374: inst = 32'h8220000;
      13375: inst = 32'h10408000;
      13376: inst = 32'hc404d06;
      13377: inst = 32'h8220000;
      13378: inst = 32'h10408000;
      13379: inst = 32'hc404d07;
      13380: inst = 32'h8220000;
      13381: inst = 32'h10408000;
      13382: inst = 32'hc404d08;
      13383: inst = 32'h8220000;
      13384: inst = 32'h10408000;
      13385: inst = 32'hc404d09;
      13386: inst = 32'h8220000;
      13387: inst = 32'h10408000;
      13388: inst = 32'hc404d0a;
      13389: inst = 32'h8220000;
      13390: inst = 32'h10408000;
      13391: inst = 32'hc404d0b;
      13392: inst = 32'h8220000;
      13393: inst = 32'h10408000;
      13394: inst = 32'hc404d0c;
      13395: inst = 32'h8220000;
      13396: inst = 32'h10408000;
      13397: inst = 32'hc404d0d;
      13398: inst = 32'h8220000;
      13399: inst = 32'h10408000;
      13400: inst = 32'hc404d0e;
      13401: inst = 32'h8220000;
      13402: inst = 32'h10408000;
      13403: inst = 32'hc404d0f;
      13404: inst = 32'h8220000;
      13405: inst = 32'h10408000;
      13406: inst = 32'hc404d10;
      13407: inst = 32'h8220000;
      13408: inst = 32'h10408000;
      13409: inst = 32'hc404d11;
      13410: inst = 32'h8220000;
      13411: inst = 32'h10408000;
      13412: inst = 32'hc404d12;
      13413: inst = 32'h8220000;
      13414: inst = 32'h10408000;
      13415: inst = 32'hc404d13;
      13416: inst = 32'h8220000;
      13417: inst = 32'h10408000;
      13418: inst = 32'hc404d14;
      13419: inst = 32'h8220000;
      13420: inst = 32'h10408000;
      13421: inst = 32'hc4055c3;
      13422: inst = 32'h8220000;
      13423: inst = 32'h10408000;
      13424: inst = 32'hc4055dc;
      13425: inst = 32'h8220000;
      13426: inst = 32'hc20ad55;
      13427: inst = 32'h10408000;
      13428: inst = 32'hc404cad;
      13429: inst = 32'h8220000;
      13430: inst = 32'hc208410;
      13431: inst = 32'h10408000;
      13432: inst = 32'hc404cae;
      13433: inst = 32'h8220000;
      13434: inst = 32'h10408000;
      13435: inst = 32'hc404caf;
      13436: inst = 32'h8220000;
      13437: inst = 32'h10408000;
      13438: inst = 32'hc404cb0;
      13439: inst = 32'h8220000;
      13440: inst = 32'h10408000;
      13441: inst = 32'hc404cb1;
      13442: inst = 32'h8220000;
      13443: inst = 32'h10408000;
      13444: inst = 32'hc404cb2;
      13445: inst = 32'h8220000;
      13446: inst = 32'h10408000;
      13447: inst = 32'hc404cb3;
      13448: inst = 32'h8220000;
      13449: inst = 32'h10408000;
      13450: inst = 32'hc404cb4;
      13451: inst = 32'h8220000;
      13452: inst = 32'h10408000;
      13453: inst = 32'hc404cb5;
      13454: inst = 32'h8220000;
      13455: inst = 32'h10408000;
      13456: inst = 32'hc40537d;
      13457: inst = 32'h8220000;
      13458: inst = 32'h10408000;
      13459: inst = 32'hc405385;
      13460: inst = 32'h8220000;
      13461: inst = 32'h10408000;
      13462: inst = 32'hc40539a;
      13463: inst = 32'h8220000;
      13464: inst = 32'h10408000;
      13465: inst = 32'hc4053a2;
      13466: inst = 32'h8220000;
      13467: inst = 32'h10408000;
      13468: inst = 32'hc4054a4;
      13469: inst = 32'h8220000;
      13470: inst = 32'h10408000;
      13471: inst = 32'hc4054bb;
      13472: inst = 32'h8220000;
      13473: inst = 32'h10408000;
      13474: inst = 32'hc405741;
      13475: inst = 32'h8220000;
      13476: inst = 32'h10408000;
      13477: inst = 32'hc40575e;
      13478: inst = 32'h8220000;
      13479: inst = 32'hc209470;
      13480: inst = 32'h10408000;
      13481: inst = 32'hc404cb6;
      13482: inst = 32'h8220000;
      13483: inst = 32'h10408000;
      13484: inst = 32'hc404d15;
      13485: inst = 32'h8220000;
      13486: inst = 32'hc20a534;
      13487: inst = 32'h10408000;
      13488: inst = 32'hc404cfb;
      13489: inst = 32'h8220000;
      13490: inst = 32'hc208c51;
      13491: inst = 32'h10408000;
      13492: inst = 32'hc404cfc;
      13493: inst = 32'h8220000;
      13494: inst = 32'h10408000;
      13495: inst = 32'hc404cfd;
      13496: inst = 32'h8220000;
      13497: inst = 32'h10408000;
      13498: inst = 32'hc4053da;
      13499: inst = 32'h8220000;
      13500: inst = 32'h10408000;
      13501: inst = 32'hc4053dc;
      13502: inst = 32'h8220000;
      13503: inst = 32'h10408000;
      13504: inst = 32'hc405403;
      13505: inst = 32'h8220000;
      13506: inst = 32'h10408000;
      13507: inst = 32'hc405405;
      13508: inst = 32'h8220000;
      13509: inst = 32'h10408000;
      13510: inst = 32'hc4054fa;
      13511: inst = 32'h8220000;
      13512: inst = 32'h10408000;
      13513: inst = 32'hc405525;
      13514: inst = 32'h8220000;
      13515: inst = 32'h10408000;
      13516: inst = 32'hc405557;
      13517: inst = 32'h8220000;
      13518: inst = 32'h10408000;
      13519: inst = 32'hc40555f;
      13520: inst = 32'h8220000;
      13521: inst = 32'h10408000;
      13522: inst = 32'hc405580;
      13523: inst = 32'h8220000;
      13524: inst = 32'h10408000;
      13525: inst = 32'hc405588;
      13526: inst = 32'h8220000;
      13527: inst = 32'h10408000;
      13528: inst = 32'hc405618;
      13529: inst = 32'h8220000;
      13530: inst = 32'h10408000;
      13531: inst = 32'hc405627;
      13532: inst = 32'h8220000;
      13533: inst = 32'h10408000;
      13534: inst = 32'hc405638;
      13535: inst = 32'h8220000;
      13536: inst = 32'h10408000;
      13537: inst = 32'hc405647;
      13538: inst = 32'h8220000;
      13539: inst = 32'h10408000;
      13540: inst = 32'hc40570b;
      13541: inst = 32'h8220000;
      13542: inst = 32'hc206b6d;
      13543: inst = 32'h10408000;
      13544: inst = 32'hc404d16;
      13545: inst = 32'h8220000;
      13546: inst = 32'h10408000;
      13547: inst = 32'hc404d75;
      13548: inst = 32'h8220000;
      13549: inst = 32'h10408000;
      13550: inst = 32'hc404d76;
      13551: inst = 32'h8220000;
      13552: inst = 32'h10408000;
      13553: inst = 32'hc404dd5;
      13554: inst = 32'h8220000;
      13555: inst = 32'h10408000;
      13556: inst = 32'hc404dd6;
      13557: inst = 32'h8220000;
      13558: inst = 32'h10408000;
      13559: inst = 32'hc404e35;
      13560: inst = 32'h8220000;
      13561: inst = 32'h10408000;
      13562: inst = 32'hc404e36;
      13563: inst = 32'h8220000;
      13564: inst = 32'h10408000;
      13565: inst = 32'hc404e95;
      13566: inst = 32'h8220000;
      13567: inst = 32'h10408000;
      13568: inst = 32'hc404e96;
      13569: inst = 32'h8220000;
      13570: inst = 32'h10408000;
      13571: inst = 32'hc404ef5;
      13572: inst = 32'h8220000;
      13573: inst = 32'h10408000;
      13574: inst = 32'hc404ef6;
      13575: inst = 32'h8220000;
      13576: inst = 32'h10408000;
      13577: inst = 32'hc404f55;
      13578: inst = 32'h8220000;
      13579: inst = 32'h10408000;
      13580: inst = 32'hc404f56;
      13581: inst = 32'h8220000;
      13582: inst = 32'h10408000;
      13583: inst = 32'hc404fb5;
      13584: inst = 32'h8220000;
      13585: inst = 32'h10408000;
      13586: inst = 32'hc404fb6;
      13587: inst = 32'h8220000;
      13588: inst = 32'h10408000;
      13589: inst = 32'hc405015;
      13590: inst = 32'h8220000;
      13591: inst = 32'h10408000;
      13592: inst = 32'hc405016;
      13593: inst = 32'h8220000;
      13594: inst = 32'h10408000;
      13595: inst = 32'hc405075;
      13596: inst = 32'h8220000;
      13597: inst = 32'h10408000;
      13598: inst = 32'hc405076;
      13599: inst = 32'h8220000;
      13600: inst = 32'h10408000;
      13601: inst = 32'hc4050d5;
      13602: inst = 32'h8220000;
      13603: inst = 32'h10408000;
      13604: inst = 32'hc4050d6;
      13605: inst = 32'h8220000;
      13606: inst = 32'h10408000;
      13607: inst = 32'hc405135;
      13608: inst = 32'h8220000;
      13609: inst = 32'h10408000;
      13610: inst = 32'hc405136;
      13611: inst = 32'h8220000;
      13612: inst = 32'h10408000;
      13613: inst = 32'hc405195;
      13614: inst = 32'h8220000;
      13615: inst = 32'h10408000;
      13616: inst = 32'hc405196;
      13617: inst = 32'h8220000;
      13618: inst = 32'h10408000;
      13619: inst = 32'hc4051f5;
      13620: inst = 32'h8220000;
      13621: inst = 32'h10408000;
      13622: inst = 32'hc4051f6;
      13623: inst = 32'h8220000;
      13624: inst = 32'h10408000;
      13625: inst = 32'hc405255;
      13626: inst = 32'h8220000;
      13627: inst = 32'h10408000;
      13628: inst = 32'hc405256;
      13629: inst = 32'h8220000;
      13630: inst = 32'h10408000;
      13631: inst = 32'hc4052b5;
      13632: inst = 32'h8220000;
      13633: inst = 32'h10408000;
      13634: inst = 32'hc4052b6;
      13635: inst = 32'h8220000;
      13636: inst = 32'h10408000;
      13637: inst = 32'hc405325;
      13638: inst = 32'h8220000;
      13639: inst = 32'h10408000;
      13640: inst = 32'hc40533a;
      13641: inst = 32'h8220000;
      13642: inst = 32'hc20c638;
      13643: inst = 32'h10408000;
      13644: inst = 32'hc404d5b;
      13645: inst = 32'h8220000;
      13646: inst = 32'hc208c71;
      13647: inst = 32'h10408000;
      13648: inst = 32'hc404d60;
      13649: inst = 32'h8220000;
      13650: inst = 32'h10408000;
      13651: inst = 32'hc404d61;
      13652: inst = 32'h8220000;
      13653: inst = 32'h10408000;
      13654: inst = 32'hc404d62;
      13655: inst = 32'h8220000;
      13656: inst = 32'h10408000;
      13657: inst = 32'hc404d63;
      13658: inst = 32'h8220000;
      13659: inst = 32'h10408000;
      13660: inst = 32'hc404d64;
      13661: inst = 32'h8220000;
      13662: inst = 32'h10408000;
      13663: inst = 32'hc404d65;
      13664: inst = 32'h8220000;
      13665: inst = 32'h10408000;
      13666: inst = 32'hc404d66;
      13667: inst = 32'h8220000;
      13668: inst = 32'h10408000;
      13669: inst = 32'hc404d67;
      13670: inst = 32'h8220000;
      13671: inst = 32'h10408000;
      13672: inst = 32'hc404d68;
      13673: inst = 32'h8220000;
      13674: inst = 32'h10408000;
      13675: inst = 32'hc404d69;
      13676: inst = 32'h8220000;
      13677: inst = 32'h10408000;
      13678: inst = 32'hc404d6a;
      13679: inst = 32'h8220000;
      13680: inst = 32'h10408000;
      13681: inst = 32'hc404d6b;
      13682: inst = 32'h8220000;
      13683: inst = 32'h10408000;
      13684: inst = 32'hc404d6c;
      13685: inst = 32'h8220000;
      13686: inst = 32'h10408000;
      13687: inst = 32'hc404d6d;
      13688: inst = 32'h8220000;
      13689: inst = 32'h10408000;
      13690: inst = 32'hc404d6e;
      13691: inst = 32'h8220000;
      13692: inst = 32'h10408000;
      13693: inst = 32'hc404d6f;
      13694: inst = 32'h8220000;
      13695: inst = 32'h10408000;
      13696: inst = 32'hc404d70;
      13697: inst = 32'h8220000;
      13698: inst = 32'h10408000;
      13699: inst = 32'hc404d71;
      13700: inst = 32'h8220000;
      13701: inst = 32'h10408000;
      13702: inst = 32'hc404d72;
      13703: inst = 32'h8220000;
      13704: inst = 32'h10408000;
      13705: inst = 32'hc404d73;
      13706: inst = 32'h8220000;
      13707: inst = 32'h10408000;
      13708: inst = 32'hc404d74;
      13709: inst = 32'h8220000;
      13710: inst = 32'h10408000;
      13711: inst = 32'hc404dc0;
      13712: inst = 32'h8220000;
      13713: inst = 32'h10408000;
      13714: inst = 32'hc404dca;
      13715: inst = 32'h8220000;
      13716: inst = 32'h10408000;
      13717: inst = 32'hc404dd4;
      13718: inst = 32'h8220000;
      13719: inst = 32'h10408000;
      13720: inst = 32'hc404e20;
      13721: inst = 32'h8220000;
      13722: inst = 32'h10408000;
      13723: inst = 32'hc404e2a;
      13724: inst = 32'h8220000;
      13725: inst = 32'h10408000;
      13726: inst = 32'hc404e34;
      13727: inst = 32'h8220000;
      13728: inst = 32'h10408000;
      13729: inst = 32'hc404e80;
      13730: inst = 32'h8220000;
      13731: inst = 32'h10408000;
      13732: inst = 32'hc404e8a;
      13733: inst = 32'h8220000;
      13734: inst = 32'h10408000;
      13735: inst = 32'hc404e94;
      13736: inst = 32'h8220000;
      13737: inst = 32'h10408000;
      13738: inst = 32'hc404ee0;
      13739: inst = 32'h8220000;
      13740: inst = 32'h10408000;
      13741: inst = 32'hc404eea;
      13742: inst = 32'h8220000;
      13743: inst = 32'h10408000;
      13744: inst = 32'hc404ef4;
      13745: inst = 32'h8220000;
      13746: inst = 32'h10408000;
      13747: inst = 32'hc404f40;
      13748: inst = 32'h8220000;
      13749: inst = 32'h10408000;
      13750: inst = 32'hc404f4a;
      13751: inst = 32'h8220000;
      13752: inst = 32'h10408000;
      13753: inst = 32'hc404f54;
      13754: inst = 32'h8220000;
      13755: inst = 32'h10408000;
      13756: inst = 32'hc404fa0;
      13757: inst = 32'h8220000;
      13758: inst = 32'h10408000;
      13759: inst = 32'hc404faa;
      13760: inst = 32'h8220000;
      13761: inst = 32'h10408000;
      13762: inst = 32'hc404fb4;
      13763: inst = 32'h8220000;
      13764: inst = 32'h10408000;
      13765: inst = 32'hc405000;
      13766: inst = 32'h8220000;
      13767: inst = 32'h10408000;
      13768: inst = 32'hc40500a;
      13769: inst = 32'h8220000;
      13770: inst = 32'h10408000;
      13771: inst = 32'hc405014;
      13772: inst = 32'h8220000;
      13773: inst = 32'h10408000;
      13774: inst = 32'hc405060;
      13775: inst = 32'h8220000;
      13776: inst = 32'h10408000;
      13777: inst = 32'hc40506a;
      13778: inst = 32'h8220000;
      13779: inst = 32'h10408000;
      13780: inst = 32'hc405074;
      13781: inst = 32'h8220000;
      13782: inst = 32'h10408000;
      13783: inst = 32'hc4050c0;
      13784: inst = 32'h8220000;
      13785: inst = 32'h10408000;
      13786: inst = 32'hc4050ca;
      13787: inst = 32'h8220000;
      13788: inst = 32'h10408000;
      13789: inst = 32'hc4050d4;
      13790: inst = 32'h8220000;
      13791: inst = 32'h10408000;
      13792: inst = 32'hc405120;
      13793: inst = 32'h8220000;
      13794: inst = 32'h10408000;
      13795: inst = 32'hc40512a;
      13796: inst = 32'h8220000;
      13797: inst = 32'h10408000;
      13798: inst = 32'hc405134;
      13799: inst = 32'h8220000;
      13800: inst = 32'h10408000;
      13801: inst = 32'hc405180;
      13802: inst = 32'h8220000;
      13803: inst = 32'h10408000;
      13804: inst = 32'hc40518a;
      13805: inst = 32'h8220000;
      13806: inst = 32'h10408000;
      13807: inst = 32'hc405194;
      13808: inst = 32'h8220000;
      13809: inst = 32'h10408000;
      13810: inst = 32'hc4051a8;
      13811: inst = 32'h8220000;
      13812: inst = 32'h10408000;
      13813: inst = 32'hc4051a9;
      13814: inst = 32'h8220000;
      13815: inst = 32'h10408000;
      13816: inst = 32'hc4051b7;
      13817: inst = 32'h8220000;
      13818: inst = 32'h10408000;
      13819: inst = 32'hc4051e0;
      13820: inst = 32'h8220000;
      13821: inst = 32'h10408000;
      13822: inst = 32'hc4051ea;
      13823: inst = 32'h8220000;
      13824: inst = 32'h10408000;
      13825: inst = 32'hc4051f4;
      13826: inst = 32'h8220000;
      13827: inst = 32'h10408000;
      13828: inst = 32'hc405208;
      13829: inst = 32'h8220000;
      13830: inst = 32'h10408000;
      13831: inst = 32'hc405217;
      13832: inst = 32'h8220000;
      13833: inst = 32'h10408000;
      13834: inst = 32'hc405240;
      13835: inst = 32'h8220000;
      13836: inst = 32'h10408000;
      13837: inst = 32'hc40524a;
      13838: inst = 32'h8220000;
      13839: inst = 32'h10408000;
      13840: inst = 32'hc405254;
      13841: inst = 32'h8220000;
      13842: inst = 32'h10408000;
      13843: inst = 32'hc40525e;
      13844: inst = 32'h8220000;
      13845: inst = 32'h10408000;
      13846: inst = 32'hc405268;
      13847: inst = 32'h8220000;
      13848: inst = 32'h10408000;
      13849: inst = 32'hc405277;
      13850: inst = 32'h8220000;
      13851: inst = 32'h10408000;
      13852: inst = 32'hc405281;
      13853: inst = 32'h8220000;
      13854: inst = 32'h10408000;
      13855: inst = 32'hc4052a0;
      13856: inst = 32'h8220000;
      13857: inst = 32'h10408000;
      13858: inst = 32'hc4052a1;
      13859: inst = 32'h8220000;
      13860: inst = 32'h10408000;
      13861: inst = 32'hc4052a2;
      13862: inst = 32'h8220000;
      13863: inst = 32'h10408000;
      13864: inst = 32'hc4052a3;
      13865: inst = 32'h8220000;
      13866: inst = 32'h10408000;
      13867: inst = 32'hc4052a4;
      13868: inst = 32'h8220000;
      13869: inst = 32'h10408000;
      13870: inst = 32'hc4052a5;
      13871: inst = 32'h8220000;
      13872: inst = 32'h10408000;
      13873: inst = 32'hc4052a6;
      13874: inst = 32'h8220000;
      13875: inst = 32'h10408000;
      13876: inst = 32'hc4052a7;
      13877: inst = 32'h8220000;
      13878: inst = 32'h10408000;
      13879: inst = 32'hc4052a8;
      13880: inst = 32'h8220000;
      13881: inst = 32'h10408000;
      13882: inst = 32'hc4052a9;
      13883: inst = 32'h8220000;
      13884: inst = 32'h10408000;
      13885: inst = 32'hc4052aa;
      13886: inst = 32'h8220000;
      13887: inst = 32'h10408000;
      13888: inst = 32'hc4052ab;
      13889: inst = 32'h8220000;
      13890: inst = 32'h10408000;
      13891: inst = 32'hc4052ac;
      13892: inst = 32'h8220000;
      13893: inst = 32'h10408000;
      13894: inst = 32'hc4052ad;
      13895: inst = 32'h8220000;
      13896: inst = 32'h10408000;
      13897: inst = 32'hc4052ae;
      13898: inst = 32'h8220000;
      13899: inst = 32'h10408000;
      13900: inst = 32'hc4052af;
      13901: inst = 32'h8220000;
      13902: inst = 32'h10408000;
      13903: inst = 32'hc4052b0;
      13904: inst = 32'h8220000;
      13905: inst = 32'h10408000;
      13906: inst = 32'hc4052b1;
      13907: inst = 32'h8220000;
      13908: inst = 32'h10408000;
      13909: inst = 32'hc4052b2;
      13910: inst = 32'h8220000;
      13911: inst = 32'h10408000;
      13912: inst = 32'hc4052b3;
      13913: inst = 32'h8220000;
      13914: inst = 32'h10408000;
      13915: inst = 32'hc4052b4;
      13916: inst = 32'h8220000;
      13917: inst = 32'h10408000;
      13918: inst = 32'hc4052bd;
      13919: inst = 32'h8220000;
      13920: inst = 32'h10408000;
      13921: inst = 32'hc4052be;
      13922: inst = 32'h8220000;
      13923: inst = 32'h10408000;
      13924: inst = 32'hc4052c8;
      13925: inst = 32'h8220000;
      13926: inst = 32'h10408000;
      13927: inst = 32'hc4052d7;
      13928: inst = 32'h8220000;
      13929: inst = 32'h10408000;
      13930: inst = 32'hc4052e1;
      13931: inst = 32'h8220000;
      13932: inst = 32'h10408000;
      13933: inst = 32'hc4052e2;
      13934: inst = 32'h8220000;
      13935: inst = 32'h10408000;
      13936: inst = 32'hc40531c;
      13937: inst = 32'h8220000;
      13938: inst = 32'h10408000;
      13939: inst = 32'hc40531d;
      13940: inst = 32'h8220000;
      13941: inst = 32'h10408000;
      13942: inst = 32'hc40531e;
      13943: inst = 32'h8220000;
      13944: inst = 32'h10408000;
      13945: inst = 32'hc40531f;
      13946: inst = 32'h8220000;
      13947: inst = 32'h10408000;
      13948: inst = 32'hc405320;
      13949: inst = 32'h8220000;
      13950: inst = 32'h10408000;
      13951: inst = 32'hc405326;
      13952: inst = 32'h8220000;
      13953: inst = 32'h10408000;
      13954: inst = 32'hc405327;
      13955: inst = 32'h8220000;
      13956: inst = 32'h10408000;
      13957: inst = 32'hc405328;
      13958: inst = 32'h8220000;
      13959: inst = 32'h10408000;
      13960: inst = 32'hc405337;
      13961: inst = 32'h8220000;
      13962: inst = 32'h10408000;
      13963: inst = 32'hc405338;
      13964: inst = 32'h8220000;
      13965: inst = 32'h10408000;
      13966: inst = 32'hc405339;
      13967: inst = 32'h8220000;
      13968: inst = 32'h10408000;
      13969: inst = 32'hc40533f;
      13970: inst = 32'h8220000;
      13971: inst = 32'h10408000;
      13972: inst = 32'hc405340;
      13973: inst = 32'h8220000;
      13974: inst = 32'h10408000;
      13975: inst = 32'hc405341;
      13976: inst = 32'h8220000;
      13977: inst = 32'h10408000;
      13978: inst = 32'hc405342;
      13979: inst = 32'h8220000;
      13980: inst = 32'h10408000;
      13981: inst = 32'hc405343;
      13982: inst = 32'h8220000;
      13983: inst = 32'h10408000;
      13984: inst = 32'hc40537b;
      13985: inst = 32'h8220000;
      13986: inst = 32'h10408000;
      13987: inst = 32'hc40537c;
      13988: inst = 32'h8220000;
      13989: inst = 32'h10408000;
      13990: inst = 32'hc405386;
      13991: inst = 32'h8220000;
      13992: inst = 32'h10408000;
      13993: inst = 32'hc405387;
      13994: inst = 32'h8220000;
      13995: inst = 32'h10408000;
      13996: inst = 32'hc405388;
      13997: inst = 32'h8220000;
      13998: inst = 32'h10408000;
      13999: inst = 32'hc405397;
      14000: inst = 32'h8220000;
      14001: inst = 32'h10408000;
      14002: inst = 32'hc405398;
      14003: inst = 32'h8220000;
      14004: inst = 32'h10408000;
      14005: inst = 32'hc405399;
      14006: inst = 32'h8220000;
      14007: inst = 32'h10408000;
      14008: inst = 32'hc4053a3;
      14009: inst = 32'h8220000;
      14010: inst = 32'h10408000;
      14011: inst = 32'hc4053a4;
      14012: inst = 32'h8220000;
      14013: inst = 32'h10408000;
      14014: inst = 32'hc4053db;
      14015: inst = 32'h8220000;
      14016: inst = 32'h10408000;
      14017: inst = 32'hc4053e5;
      14018: inst = 32'h8220000;
      14019: inst = 32'h10408000;
      14020: inst = 32'hc4053e6;
      14021: inst = 32'h8220000;
      14022: inst = 32'h10408000;
      14023: inst = 32'hc4053e7;
      14024: inst = 32'h8220000;
      14025: inst = 32'h10408000;
      14026: inst = 32'hc4053f8;
      14027: inst = 32'h8220000;
      14028: inst = 32'h10408000;
      14029: inst = 32'hc4053f9;
      14030: inst = 32'h8220000;
      14031: inst = 32'h10408000;
      14032: inst = 32'hc4053fa;
      14033: inst = 32'h8220000;
      14034: inst = 32'h10408000;
      14035: inst = 32'hc405404;
      14036: inst = 32'h8220000;
      14037: inst = 32'h10408000;
      14038: inst = 32'hc40543a;
      14039: inst = 32'h8220000;
      14040: inst = 32'h10408000;
      14041: inst = 32'hc40543b;
      14042: inst = 32'h8220000;
      14043: inst = 32'h10408000;
      14044: inst = 32'hc405445;
      14045: inst = 32'h8220000;
      14046: inst = 32'h10408000;
      14047: inst = 32'hc405446;
      14048: inst = 32'h8220000;
      14049: inst = 32'h10408000;
      14050: inst = 32'hc405447;
      14051: inst = 32'h8220000;
      14052: inst = 32'h10408000;
      14053: inst = 32'hc405458;
      14054: inst = 32'h8220000;
      14055: inst = 32'h10408000;
      14056: inst = 32'hc405459;
      14057: inst = 32'h8220000;
      14058: inst = 32'h10408000;
      14059: inst = 32'hc40545a;
      14060: inst = 32'h8220000;
      14061: inst = 32'h10408000;
      14062: inst = 32'hc405464;
      14063: inst = 32'h8220000;
      14064: inst = 32'h10408000;
      14065: inst = 32'hc405465;
      14066: inst = 32'h8220000;
      14067: inst = 32'h10408000;
      14068: inst = 32'hc405499;
      14069: inst = 32'h8220000;
      14070: inst = 32'h10408000;
      14071: inst = 32'hc40549a;
      14072: inst = 32'h8220000;
      14073: inst = 32'h10408000;
      14074: inst = 32'hc4054a5;
      14075: inst = 32'h8220000;
      14076: inst = 32'h10408000;
      14077: inst = 32'hc4054a6;
      14078: inst = 32'h8220000;
      14079: inst = 32'h10408000;
      14080: inst = 32'hc4054a7;
      14081: inst = 32'h8220000;
      14082: inst = 32'h10408000;
      14083: inst = 32'hc4054b8;
      14084: inst = 32'h8220000;
      14085: inst = 32'h10408000;
      14086: inst = 32'hc4054b9;
      14087: inst = 32'h8220000;
      14088: inst = 32'h10408000;
      14089: inst = 32'hc4054ba;
      14090: inst = 32'h8220000;
      14091: inst = 32'h10408000;
      14092: inst = 32'hc4054c5;
      14093: inst = 32'h8220000;
      14094: inst = 32'h10408000;
      14095: inst = 32'hc4054c6;
      14096: inst = 32'h8220000;
      14097: inst = 32'h10408000;
      14098: inst = 32'hc4054f8;
      14099: inst = 32'h8220000;
      14100: inst = 32'h10408000;
      14101: inst = 32'hc4054f9;
      14102: inst = 32'h8220000;
      14103: inst = 32'h10408000;
      14104: inst = 32'hc405500;
      14105: inst = 32'h8220000;
      14106: inst = 32'h10408000;
      14107: inst = 32'hc405504;
      14108: inst = 32'h8220000;
      14109: inst = 32'h10408000;
      14110: inst = 32'hc405505;
      14111: inst = 32'h8220000;
      14112: inst = 32'h10408000;
      14113: inst = 32'hc405506;
      14114: inst = 32'h8220000;
      14115: inst = 32'h10408000;
      14116: inst = 32'hc405507;
      14117: inst = 32'h8220000;
      14118: inst = 32'h10408000;
      14119: inst = 32'hc405518;
      14120: inst = 32'h8220000;
      14121: inst = 32'h10408000;
      14122: inst = 32'hc405519;
      14123: inst = 32'h8220000;
      14124: inst = 32'h10408000;
      14125: inst = 32'hc40551a;
      14126: inst = 32'h8220000;
      14127: inst = 32'h10408000;
      14128: inst = 32'hc40551b;
      14129: inst = 32'h8220000;
      14130: inst = 32'h10408000;
      14131: inst = 32'hc40551f;
      14132: inst = 32'h8220000;
      14133: inst = 32'h10408000;
      14134: inst = 32'hc405526;
      14135: inst = 32'h8220000;
      14136: inst = 32'h10408000;
      14137: inst = 32'hc405527;
      14138: inst = 32'h8220000;
      14139: inst = 32'h10408000;
      14140: inst = 32'hc405558;
      14141: inst = 32'h8220000;
      14142: inst = 32'h10408000;
      14143: inst = 32'hc405559;
      14144: inst = 32'h8220000;
      14145: inst = 32'h10408000;
      14146: inst = 32'hc405560;
      14147: inst = 32'h8220000;
      14148: inst = 32'h10408000;
      14149: inst = 32'hc405564;
      14150: inst = 32'h8220000;
      14151: inst = 32'h10408000;
      14152: inst = 32'hc405565;
      14153: inst = 32'h8220000;
      14154: inst = 32'h10408000;
      14155: inst = 32'hc405566;
      14156: inst = 32'h8220000;
      14157: inst = 32'h10408000;
      14158: inst = 32'hc405567;
      14159: inst = 32'h8220000;
      14160: inst = 32'h10408000;
      14161: inst = 32'hc405578;
      14162: inst = 32'h8220000;
      14163: inst = 32'h10408000;
      14164: inst = 32'hc405579;
      14165: inst = 32'h8220000;
      14166: inst = 32'h10408000;
      14167: inst = 32'hc40557a;
      14168: inst = 32'h8220000;
      14169: inst = 32'h10408000;
      14170: inst = 32'hc40557b;
      14171: inst = 32'h8220000;
      14172: inst = 32'h10408000;
      14173: inst = 32'hc40557f;
      14174: inst = 32'h8220000;
      14175: inst = 32'h10408000;
      14176: inst = 32'hc405586;
      14177: inst = 32'h8220000;
      14178: inst = 32'h10408000;
      14179: inst = 32'hc405587;
      14180: inst = 32'h8220000;
      14181: inst = 32'h10408000;
      14182: inst = 32'hc4055b7;
      14183: inst = 32'h8220000;
      14184: inst = 32'h10408000;
      14185: inst = 32'hc4055b8;
      14186: inst = 32'h8220000;
      14187: inst = 32'h10408000;
      14188: inst = 32'hc4055bf;
      14189: inst = 32'h8220000;
      14190: inst = 32'h10408000;
      14191: inst = 32'hc4055c0;
      14192: inst = 32'h8220000;
      14193: inst = 32'h10408000;
      14194: inst = 32'hc4055c4;
      14195: inst = 32'h8220000;
      14196: inst = 32'h10408000;
      14197: inst = 32'hc4055c5;
      14198: inst = 32'h8220000;
      14199: inst = 32'h10408000;
      14200: inst = 32'hc4055c6;
      14201: inst = 32'h8220000;
      14202: inst = 32'h10408000;
      14203: inst = 32'hc4055c7;
      14204: inst = 32'h8220000;
      14205: inst = 32'h10408000;
      14206: inst = 32'hc4055d8;
      14207: inst = 32'h8220000;
      14208: inst = 32'h10408000;
      14209: inst = 32'hc4055d9;
      14210: inst = 32'h8220000;
      14211: inst = 32'h10408000;
      14212: inst = 32'hc4055da;
      14213: inst = 32'h8220000;
      14214: inst = 32'h10408000;
      14215: inst = 32'hc4055db;
      14216: inst = 32'h8220000;
      14217: inst = 32'h10408000;
      14218: inst = 32'hc4055df;
      14219: inst = 32'h8220000;
      14220: inst = 32'h10408000;
      14221: inst = 32'hc4055e0;
      14222: inst = 32'h8220000;
      14223: inst = 32'h10408000;
      14224: inst = 32'hc4055e7;
      14225: inst = 32'h8220000;
      14226: inst = 32'h10408000;
      14227: inst = 32'hc4055e8;
      14228: inst = 32'h8220000;
      14229: inst = 32'h10408000;
      14230: inst = 32'hc405616;
      14231: inst = 32'h8220000;
      14232: inst = 32'h10408000;
      14233: inst = 32'hc405617;
      14234: inst = 32'h8220000;
      14235: inst = 32'h10408000;
      14236: inst = 32'hc40561f;
      14237: inst = 32'h8220000;
      14238: inst = 32'h10408000;
      14239: inst = 32'hc405620;
      14240: inst = 32'h8220000;
      14241: inst = 32'h10408000;
      14242: inst = 32'hc405623;
      14243: inst = 32'h8220000;
      14244: inst = 32'h10408000;
      14245: inst = 32'hc405624;
      14246: inst = 32'h8220000;
      14247: inst = 32'h10408000;
      14248: inst = 32'hc405625;
      14249: inst = 32'h8220000;
      14250: inst = 32'h10408000;
      14251: inst = 32'hc405626;
      14252: inst = 32'h8220000;
      14253: inst = 32'h10408000;
      14254: inst = 32'hc405639;
      14255: inst = 32'h8220000;
      14256: inst = 32'h10408000;
      14257: inst = 32'hc40563a;
      14258: inst = 32'h8220000;
      14259: inst = 32'h10408000;
      14260: inst = 32'hc40563b;
      14261: inst = 32'h8220000;
      14262: inst = 32'h10408000;
      14263: inst = 32'hc40563c;
      14264: inst = 32'h8220000;
      14265: inst = 32'h10408000;
      14266: inst = 32'hc40563f;
      14267: inst = 32'h8220000;
      14268: inst = 32'h10408000;
      14269: inst = 32'hc405640;
      14270: inst = 32'h8220000;
      14271: inst = 32'h10408000;
      14272: inst = 32'hc405648;
      14273: inst = 32'h8220000;
      14274: inst = 32'h10408000;
      14275: inst = 32'hc405649;
      14276: inst = 32'h8220000;
      14277: inst = 32'h10408000;
      14278: inst = 32'hc405675;
      14279: inst = 32'h8220000;
      14280: inst = 32'h10408000;
      14281: inst = 32'hc405676;
      14282: inst = 32'h8220000;
      14283: inst = 32'h10408000;
      14284: inst = 32'hc405677;
      14285: inst = 32'h8220000;
      14286: inst = 32'h10408000;
      14287: inst = 32'hc40567e;
      14288: inst = 32'h8220000;
      14289: inst = 32'h10408000;
      14290: inst = 32'hc40567f;
      14291: inst = 32'h8220000;
      14292: inst = 32'h10408000;
      14293: inst = 32'hc405680;
      14294: inst = 32'h8220000;
      14295: inst = 32'h10408000;
      14296: inst = 32'hc405683;
      14297: inst = 32'h8220000;
      14298: inst = 32'h10408000;
      14299: inst = 32'hc405684;
      14300: inst = 32'h8220000;
      14301: inst = 32'h10408000;
      14302: inst = 32'hc405685;
      14303: inst = 32'h8220000;
      14304: inst = 32'h10408000;
      14305: inst = 32'hc405686;
      14306: inst = 32'h8220000;
      14307: inst = 32'h10408000;
      14308: inst = 32'hc405699;
      14309: inst = 32'h8220000;
      14310: inst = 32'h10408000;
      14311: inst = 32'hc40569a;
      14312: inst = 32'h8220000;
      14313: inst = 32'h10408000;
      14314: inst = 32'hc40569b;
      14315: inst = 32'h8220000;
      14316: inst = 32'h10408000;
      14317: inst = 32'hc40569c;
      14318: inst = 32'h8220000;
      14319: inst = 32'h10408000;
      14320: inst = 32'hc40569f;
      14321: inst = 32'h8220000;
      14322: inst = 32'h10408000;
      14323: inst = 32'hc4056a0;
      14324: inst = 32'h8220000;
      14325: inst = 32'h10408000;
      14326: inst = 32'hc4056a1;
      14327: inst = 32'h8220000;
      14328: inst = 32'h10408000;
      14329: inst = 32'hc4056a8;
      14330: inst = 32'h8220000;
      14331: inst = 32'h10408000;
      14332: inst = 32'hc4056a9;
      14333: inst = 32'h8220000;
      14334: inst = 32'h10408000;
      14335: inst = 32'hc4056aa;
      14336: inst = 32'h8220000;
      14337: inst = 32'h10408000;
      14338: inst = 32'hc4056d4;
      14339: inst = 32'h8220000;
      14340: inst = 32'h10408000;
      14341: inst = 32'hc4056d5;
      14342: inst = 32'h8220000;
      14343: inst = 32'h10408000;
      14344: inst = 32'hc4056d6;
      14345: inst = 32'h8220000;
      14346: inst = 32'h10408000;
      14347: inst = 32'hc4056d7;
      14348: inst = 32'h8220000;
      14349: inst = 32'h10408000;
      14350: inst = 32'hc4056d8;
      14351: inst = 32'h8220000;
      14352: inst = 32'h10408000;
      14353: inst = 32'hc4056d9;
      14354: inst = 32'h8220000;
      14355: inst = 32'h10408000;
      14356: inst = 32'hc4056da;
      14357: inst = 32'h8220000;
      14358: inst = 32'h10408000;
      14359: inst = 32'hc4056db;
      14360: inst = 32'h8220000;
      14361: inst = 32'h10408000;
      14362: inst = 32'hc4056dc;
      14363: inst = 32'h8220000;
      14364: inst = 32'h10408000;
      14365: inst = 32'hc4056dd;
      14366: inst = 32'h8220000;
      14367: inst = 32'h10408000;
      14368: inst = 32'hc4056de;
      14369: inst = 32'h8220000;
      14370: inst = 32'h10408000;
      14371: inst = 32'hc4056df;
      14372: inst = 32'h8220000;
      14373: inst = 32'h10408000;
      14374: inst = 32'hc4056e0;
      14375: inst = 32'h8220000;
      14376: inst = 32'h10408000;
      14377: inst = 32'hc4056e3;
      14378: inst = 32'h8220000;
      14379: inst = 32'h10408000;
      14380: inst = 32'hc4056e4;
      14381: inst = 32'h8220000;
      14382: inst = 32'h10408000;
      14383: inst = 32'hc4056e5;
      14384: inst = 32'h8220000;
      14385: inst = 32'h10408000;
      14386: inst = 32'hc4056e6;
      14387: inst = 32'h8220000;
      14388: inst = 32'h10408000;
      14389: inst = 32'hc4056f9;
      14390: inst = 32'h8220000;
      14391: inst = 32'h10408000;
      14392: inst = 32'hc4056fa;
      14393: inst = 32'h8220000;
      14394: inst = 32'h10408000;
      14395: inst = 32'hc4056fb;
      14396: inst = 32'h8220000;
      14397: inst = 32'h10408000;
      14398: inst = 32'hc4056fc;
      14399: inst = 32'h8220000;
      14400: inst = 32'h10408000;
      14401: inst = 32'hc4056ff;
      14402: inst = 32'h8220000;
      14403: inst = 32'h10408000;
      14404: inst = 32'hc405700;
      14405: inst = 32'h8220000;
      14406: inst = 32'h10408000;
      14407: inst = 32'hc405701;
      14408: inst = 32'h8220000;
      14409: inst = 32'h10408000;
      14410: inst = 32'hc405702;
      14411: inst = 32'h8220000;
      14412: inst = 32'h10408000;
      14413: inst = 32'hc405703;
      14414: inst = 32'h8220000;
      14415: inst = 32'h10408000;
      14416: inst = 32'hc405704;
      14417: inst = 32'h8220000;
      14418: inst = 32'h10408000;
      14419: inst = 32'hc405705;
      14420: inst = 32'h8220000;
      14421: inst = 32'h10408000;
      14422: inst = 32'hc405706;
      14423: inst = 32'h8220000;
      14424: inst = 32'h10408000;
      14425: inst = 32'hc405707;
      14426: inst = 32'h8220000;
      14427: inst = 32'h10408000;
      14428: inst = 32'hc405708;
      14429: inst = 32'h8220000;
      14430: inst = 32'h10408000;
      14431: inst = 32'hc405709;
      14432: inst = 32'h8220000;
      14433: inst = 32'h10408000;
      14434: inst = 32'hc40570a;
      14435: inst = 32'h8220000;
      14436: inst = 32'h10408000;
      14437: inst = 32'hc405734;
      14438: inst = 32'h8220000;
      14439: inst = 32'h10408000;
      14440: inst = 32'hc405735;
      14441: inst = 32'h8220000;
      14442: inst = 32'h10408000;
      14443: inst = 32'hc405736;
      14444: inst = 32'h8220000;
      14445: inst = 32'h10408000;
      14446: inst = 32'hc405737;
      14447: inst = 32'h8220000;
      14448: inst = 32'h10408000;
      14449: inst = 32'hc405738;
      14450: inst = 32'h8220000;
      14451: inst = 32'h10408000;
      14452: inst = 32'hc405739;
      14453: inst = 32'h8220000;
      14454: inst = 32'h10408000;
      14455: inst = 32'hc40573a;
      14456: inst = 32'h8220000;
      14457: inst = 32'h10408000;
      14458: inst = 32'hc40573b;
      14459: inst = 32'h8220000;
      14460: inst = 32'h10408000;
      14461: inst = 32'hc40573c;
      14462: inst = 32'h8220000;
      14463: inst = 32'h10408000;
      14464: inst = 32'hc40573d;
      14465: inst = 32'h8220000;
      14466: inst = 32'h10408000;
      14467: inst = 32'hc40573e;
      14468: inst = 32'h8220000;
      14469: inst = 32'h10408000;
      14470: inst = 32'hc40573f;
      14471: inst = 32'h8220000;
      14472: inst = 32'h10408000;
      14473: inst = 32'hc405740;
      14474: inst = 32'h8220000;
      14475: inst = 32'h10408000;
      14476: inst = 32'hc405742;
      14477: inst = 32'h8220000;
      14478: inst = 32'h10408000;
      14479: inst = 32'hc405743;
      14480: inst = 32'h8220000;
      14481: inst = 32'h10408000;
      14482: inst = 32'hc405744;
      14483: inst = 32'h8220000;
      14484: inst = 32'h10408000;
      14485: inst = 32'hc405745;
      14486: inst = 32'h8220000;
      14487: inst = 32'h10408000;
      14488: inst = 32'hc405746;
      14489: inst = 32'h8220000;
      14490: inst = 32'h10408000;
      14491: inst = 32'hc405759;
      14492: inst = 32'h8220000;
      14493: inst = 32'h10408000;
      14494: inst = 32'hc40575a;
      14495: inst = 32'h8220000;
      14496: inst = 32'h10408000;
      14497: inst = 32'hc40575b;
      14498: inst = 32'h8220000;
      14499: inst = 32'h10408000;
      14500: inst = 32'hc40575c;
      14501: inst = 32'h8220000;
      14502: inst = 32'h10408000;
      14503: inst = 32'hc40575d;
      14504: inst = 32'h8220000;
      14505: inst = 32'h10408000;
      14506: inst = 32'hc40575f;
      14507: inst = 32'h8220000;
      14508: inst = 32'h10408000;
      14509: inst = 32'hc405760;
      14510: inst = 32'h8220000;
      14511: inst = 32'h10408000;
      14512: inst = 32'hc405761;
      14513: inst = 32'h8220000;
      14514: inst = 32'h10408000;
      14515: inst = 32'hc405762;
      14516: inst = 32'h8220000;
      14517: inst = 32'h10408000;
      14518: inst = 32'hc405763;
      14519: inst = 32'h8220000;
      14520: inst = 32'h10408000;
      14521: inst = 32'hc405764;
      14522: inst = 32'h8220000;
      14523: inst = 32'h10408000;
      14524: inst = 32'hc405765;
      14525: inst = 32'h8220000;
      14526: inst = 32'h10408000;
      14527: inst = 32'hc405766;
      14528: inst = 32'h8220000;
      14529: inst = 32'h10408000;
      14530: inst = 32'hc405767;
      14531: inst = 32'h8220000;
      14532: inst = 32'h10408000;
      14533: inst = 32'hc405768;
      14534: inst = 32'h8220000;
      14535: inst = 32'h10408000;
      14536: inst = 32'hc405769;
      14537: inst = 32'h8220000;
      14538: inst = 32'h10408000;
      14539: inst = 32'hc40576a;
      14540: inst = 32'h8220000;
      14541: inst = 32'h10408000;
      14542: inst = 32'hc40576b;
      14543: inst = 32'h8220000;
      14544: inst = 32'h10408000;
      14545: inst = 32'hc405793;
      14546: inst = 32'h8220000;
      14547: inst = 32'h10408000;
      14548: inst = 32'hc405794;
      14549: inst = 32'h8220000;
      14550: inst = 32'h10408000;
      14551: inst = 32'hc405795;
      14552: inst = 32'h8220000;
      14553: inst = 32'h10408000;
      14554: inst = 32'hc405796;
      14555: inst = 32'h8220000;
      14556: inst = 32'h10408000;
      14557: inst = 32'hc405797;
      14558: inst = 32'h8220000;
      14559: inst = 32'h10408000;
      14560: inst = 32'hc405798;
      14561: inst = 32'h8220000;
      14562: inst = 32'h10408000;
      14563: inst = 32'hc405799;
      14564: inst = 32'h8220000;
      14565: inst = 32'h10408000;
      14566: inst = 32'hc40579a;
      14567: inst = 32'h8220000;
      14568: inst = 32'h10408000;
      14569: inst = 32'hc40579b;
      14570: inst = 32'h8220000;
      14571: inst = 32'h10408000;
      14572: inst = 32'hc40579c;
      14573: inst = 32'h8220000;
      14574: inst = 32'h10408000;
      14575: inst = 32'hc40579d;
      14576: inst = 32'h8220000;
      14577: inst = 32'h10408000;
      14578: inst = 32'hc40579e;
      14579: inst = 32'h8220000;
      14580: inst = 32'h10408000;
      14581: inst = 32'hc40579f;
      14582: inst = 32'h8220000;
      14583: inst = 32'h10408000;
      14584: inst = 32'hc4057a0;
      14585: inst = 32'h8220000;
      14586: inst = 32'h10408000;
      14587: inst = 32'hc4057a1;
      14588: inst = 32'h8220000;
      14589: inst = 32'h10408000;
      14590: inst = 32'hc4057a2;
      14591: inst = 32'h8220000;
      14592: inst = 32'h10408000;
      14593: inst = 32'hc4057a3;
      14594: inst = 32'h8220000;
      14595: inst = 32'h10408000;
      14596: inst = 32'hc4057a4;
      14597: inst = 32'h8220000;
      14598: inst = 32'h10408000;
      14599: inst = 32'hc4057a5;
      14600: inst = 32'h8220000;
      14601: inst = 32'h10408000;
      14602: inst = 32'hc4057a6;
      14603: inst = 32'h8220000;
      14604: inst = 32'h10408000;
      14605: inst = 32'hc4057b9;
      14606: inst = 32'h8220000;
      14607: inst = 32'h10408000;
      14608: inst = 32'hc4057ba;
      14609: inst = 32'h8220000;
      14610: inst = 32'h10408000;
      14611: inst = 32'hc4057bb;
      14612: inst = 32'h8220000;
      14613: inst = 32'h10408000;
      14614: inst = 32'hc4057bc;
      14615: inst = 32'h8220000;
      14616: inst = 32'h10408000;
      14617: inst = 32'hc4057bd;
      14618: inst = 32'h8220000;
      14619: inst = 32'h10408000;
      14620: inst = 32'hc4057be;
      14621: inst = 32'h8220000;
      14622: inst = 32'h10408000;
      14623: inst = 32'hc4057bf;
      14624: inst = 32'h8220000;
      14625: inst = 32'h10408000;
      14626: inst = 32'hc4057c0;
      14627: inst = 32'h8220000;
      14628: inst = 32'h10408000;
      14629: inst = 32'hc4057c1;
      14630: inst = 32'h8220000;
      14631: inst = 32'h10408000;
      14632: inst = 32'hc4057c2;
      14633: inst = 32'h8220000;
      14634: inst = 32'h10408000;
      14635: inst = 32'hc4057c3;
      14636: inst = 32'h8220000;
      14637: inst = 32'h10408000;
      14638: inst = 32'hc4057c4;
      14639: inst = 32'h8220000;
      14640: inst = 32'h10408000;
      14641: inst = 32'hc4057c5;
      14642: inst = 32'h8220000;
      14643: inst = 32'h10408000;
      14644: inst = 32'hc4057c6;
      14645: inst = 32'h8220000;
      14646: inst = 32'h10408000;
      14647: inst = 32'hc4057c7;
      14648: inst = 32'h8220000;
      14649: inst = 32'h10408000;
      14650: inst = 32'hc4057c8;
      14651: inst = 32'h8220000;
      14652: inst = 32'h10408000;
      14653: inst = 32'hc4057c9;
      14654: inst = 32'h8220000;
      14655: inst = 32'h10408000;
      14656: inst = 32'hc4057ca;
      14657: inst = 32'h8220000;
      14658: inst = 32'h10408000;
      14659: inst = 32'hc4057cb;
      14660: inst = 32'h8220000;
      14661: inst = 32'h10408000;
      14662: inst = 32'hc4057cc;
      14663: inst = 32'h8220000;
      14664: inst = 32'hc20bdd7;
      14665: inst = 32'h10408000;
      14666: inst = 32'hc404dc1;
      14667: inst = 32'h8220000;
      14668: inst = 32'h10408000;
      14669: inst = 32'hc404dc2;
      14670: inst = 32'h8220000;
      14671: inst = 32'h10408000;
      14672: inst = 32'hc404dc3;
      14673: inst = 32'h8220000;
      14674: inst = 32'h10408000;
      14675: inst = 32'hc404dc4;
      14676: inst = 32'h8220000;
      14677: inst = 32'h10408000;
      14678: inst = 32'hc404dc5;
      14679: inst = 32'h8220000;
      14680: inst = 32'h10408000;
      14681: inst = 32'hc404dc6;
      14682: inst = 32'h8220000;
      14683: inst = 32'h10408000;
      14684: inst = 32'hc404dc7;
      14685: inst = 32'h8220000;
      14686: inst = 32'h10408000;
      14687: inst = 32'hc404dc8;
      14688: inst = 32'h8220000;
      14689: inst = 32'h10408000;
      14690: inst = 32'hc404dc9;
      14691: inst = 32'h8220000;
      14692: inst = 32'h10408000;
      14693: inst = 32'hc404dcb;
      14694: inst = 32'h8220000;
      14695: inst = 32'h10408000;
      14696: inst = 32'hc404dcc;
      14697: inst = 32'h8220000;
      14698: inst = 32'h10408000;
      14699: inst = 32'hc404dcd;
      14700: inst = 32'h8220000;
      14701: inst = 32'h10408000;
      14702: inst = 32'hc404dce;
      14703: inst = 32'h8220000;
      14704: inst = 32'h10408000;
      14705: inst = 32'hc404dcf;
      14706: inst = 32'h8220000;
      14707: inst = 32'h10408000;
      14708: inst = 32'hc404dd0;
      14709: inst = 32'h8220000;
      14710: inst = 32'h10408000;
      14711: inst = 32'hc404dd1;
      14712: inst = 32'h8220000;
      14713: inst = 32'h10408000;
      14714: inst = 32'hc404dd2;
      14715: inst = 32'h8220000;
      14716: inst = 32'h10408000;
      14717: inst = 32'hc404dd3;
      14718: inst = 32'h8220000;
      14719: inst = 32'h10408000;
      14720: inst = 32'hc404e21;
      14721: inst = 32'h8220000;
      14722: inst = 32'h10408000;
      14723: inst = 32'hc404e22;
      14724: inst = 32'h8220000;
      14725: inst = 32'h10408000;
      14726: inst = 32'hc404e23;
      14727: inst = 32'h8220000;
      14728: inst = 32'h10408000;
      14729: inst = 32'hc404e24;
      14730: inst = 32'h8220000;
      14731: inst = 32'h10408000;
      14732: inst = 32'hc404e25;
      14733: inst = 32'h8220000;
      14734: inst = 32'h10408000;
      14735: inst = 32'hc404e26;
      14736: inst = 32'h8220000;
      14737: inst = 32'h10408000;
      14738: inst = 32'hc404e27;
      14739: inst = 32'h8220000;
      14740: inst = 32'h10408000;
      14741: inst = 32'hc404e28;
      14742: inst = 32'h8220000;
      14743: inst = 32'h10408000;
      14744: inst = 32'hc404e29;
      14745: inst = 32'h8220000;
      14746: inst = 32'h10408000;
      14747: inst = 32'hc404e2b;
      14748: inst = 32'h8220000;
      14749: inst = 32'h10408000;
      14750: inst = 32'hc404e2c;
      14751: inst = 32'h8220000;
      14752: inst = 32'h10408000;
      14753: inst = 32'hc404e2d;
      14754: inst = 32'h8220000;
      14755: inst = 32'h10408000;
      14756: inst = 32'hc404e2e;
      14757: inst = 32'h8220000;
      14758: inst = 32'h10408000;
      14759: inst = 32'hc404e2f;
      14760: inst = 32'h8220000;
      14761: inst = 32'h10408000;
      14762: inst = 32'hc404e30;
      14763: inst = 32'h8220000;
      14764: inst = 32'h10408000;
      14765: inst = 32'hc404e31;
      14766: inst = 32'h8220000;
      14767: inst = 32'h10408000;
      14768: inst = 32'hc404e32;
      14769: inst = 32'h8220000;
      14770: inst = 32'h10408000;
      14771: inst = 32'hc404e33;
      14772: inst = 32'h8220000;
      14773: inst = 32'h10408000;
      14774: inst = 32'hc404e81;
      14775: inst = 32'h8220000;
      14776: inst = 32'h10408000;
      14777: inst = 32'hc404e82;
      14778: inst = 32'h8220000;
      14779: inst = 32'h10408000;
      14780: inst = 32'hc404e83;
      14781: inst = 32'h8220000;
      14782: inst = 32'h10408000;
      14783: inst = 32'hc404e84;
      14784: inst = 32'h8220000;
      14785: inst = 32'h10408000;
      14786: inst = 32'hc404e85;
      14787: inst = 32'h8220000;
      14788: inst = 32'h10408000;
      14789: inst = 32'hc404e86;
      14790: inst = 32'h8220000;
      14791: inst = 32'h10408000;
      14792: inst = 32'hc404e87;
      14793: inst = 32'h8220000;
      14794: inst = 32'h10408000;
      14795: inst = 32'hc404e88;
      14796: inst = 32'h8220000;
      14797: inst = 32'h10408000;
      14798: inst = 32'hc404e89;
      14799: inst = 32'h8220000;
      14800: inst = 32'h10408000;
      14801: inst = 32'hc404e8b;
      14802: inst = 32'h8220000;
      14803: inst = 32'h10408000;
      14804: inst = 32'hc404e8c;
      14805: inst = 32'h8220000;
      14806: inst = 32'h10408000;
      14807: inst = 32'hc404e8d;
      14808: inst = 32'h8220000;
      14809: inst = 32'h10408000;
      14810: inst = 32'hc404e8e;
      14811: inst = 32'h8220000;
      14812: inst = 32'h10408000;
      14813: inst = 32'hc404e8f;
      14814: inst = 32'h8220000;
      14815: inst = 32'h10408000;
      14816: inst = 32'hc404e90;
      14817: inst = 32'h8220000;
      14818: inst = 32'h10408000;
      14819: inst = 32'hc404e91;
      14820: inst = 32'h8220000;
      14821: inst = 32'h10408000;
      14822: inst = 32'hc404e92;
      14823: inst = 32'h8220000;
      14824: inst = 32'h10408000;
      14825: inst = 32'hc404e93;
      14826: inst = 32'h8220000;
      14827: inst = 32'h10408000;
      14828: inst = 32'hc404ee1;
      14829: inst = 32'h8220000;
      14830: inst = 32'h10408000;
      14831: inst = 32'hc404ee2;
      14832: inst = 32'h8220000;
      14833: inst = 32'h10408000;
      14834: inst = 32'hc404ee3;
      14835: inst = 32'h8220000;
      14836: inst = 32'h10408000;
      14837: inst = 32'hc404ee4;
      14838: inst = 32'h8220000;
      14839: inst = 32'h10408000;
      14840: inst = 32'hc404ee5;
      14841: inst = 32'h8220000;
      14842: inst = 32'h10408000;
      14843: inst = 32'hc404ee6;
      14844: inst = 32'h8220000;
      14845: inst = 32'h10408000;
      14846: inst = 32'hc404ee7;
      14847: inst = 32'h8220000;
      14848: inst = 32'h10408000;
      14849: inst = 32'hc404ee8;
      14850: inst = 32'h8220000;
      14851: inst = 32'h10408000;
      14852: inst = 32'hc404ee9;
      14853: inst = 32'h8220000;
      14854: inst = 32'h10408000;
      14855: inst = 32'hc404eeb;
      14856: inst = 32'h8220000;
      14857: inst = 32'h10408000;
      14858: inst = 32'hc404eec;
      14859: inst = 32'h8220000;
      14860: inst = 32'h10408000;
      14861: inst = 32'hc404eed;
      14862: inst = 32'h8220000;
      14863: inst = 32'h10408000;
      14864: inst = 32'hc404eee;
      14865: inst = 32'h8220000;
      14866: inst = 32'h10408000;
      14867: inst = 32'hc404eef;
      14868: inst = 32'h8220000;
      14869: inst = 32'h10408000;
      14870: inst = 32'hc404ef0;
      14871: inst = 32'h8220000;
      14872: inst = 32'h10408000;
      14873: inst = 32'hc404ef1;
      14874: inst = 32'h8220000;
      14875: inst = 32'h10408000;
      14876: inst = 32'hc404ef2;
      14877: inst = 32'h8220000;
      14878: inst = 32'h10408000;
      14879: inst = 32'hc404ef3;
      14880: inst = 32'h8220000;
      14881: inst = 32'h10408000;
      14882: inst = 32'hc404f41;
      14883: inst = 32'h8220000;
      14884: inst = 32'h10408000;
      14885: inst = 32'hc404f42;
      14886: inst = 32'h8220000;
      14887: inst = 32'h10408000;
      14888: inst = 32'hc404f43;
      14889: inst = 32'h8220000;
      14890: inst = 32'h10408000;
      14891: inst = 32'hc404f44;
      14892: inst = 32'h8220000;
      14893: inst = 32'h10408000;
      14894: inst = 32'hc404f45;
      14895: inst = 32'h8220000;
      14896: inst = 32'h10408000;
      14897: inst = 32'hc404f46;
      14898: inst = 32'h8220000;
      14899: inst = 32'h10408000;
      14900: inst = 32'hc404f47;
      14901: inst = 32'h8220000;
      14902: inst = 32'h10408000;
      14903: inst = 32'hc404f48;
      14904: inst = 32'h8220000;
      14905: inst = 32'h10408000;
      14906: inst = 32'hc404f49;
      14907: inst = 32'h8220000;
      14908: inst = 32'h10408000;
      14909: inst = 32'hc404f4b;
      14910: inst = 32'h8220000;
      14911: inst = 32'h10408000;
      14912: inst = 32'hc404f4c;
      14913: inst = 32'h8220000;
      14914: inst = 32'h10408000;
      14915: inst = 32'hc404f4d;
      14916: inst = 32'h8220000;
      14917: inst = 32'h10408000;
      14918: inst = 32'hc404f4e;
      14919: inst = 32'h8220000;
      14920: inst = 32'h10408000;
      14921: inst = 32'hc404f4f;
      14922: inst = 32'h8220000;
      14923: inst = 32'h10408000;
      14924: inst = 32'hc404f50;
      14925: inst = 32'h8220000;
      14926: inst = 32'h10408000;
      14927: inst = 32'hc404f51;
      14928: inst = 32'h8220000;
      14929: inst = 32'h10408000;
      14930: inst = 32'hc404f52;
      14931: inst = 32'h8220000;
      14932: inst = 32'h10408000;
      14933: inst = 32'hc404f53;
      14934: inst = 32'h8220000;
      14935: inst = 32'h10408000;
      14936: inst = 32'hc404fa1;
      14937: inst = 32'h8220000;
      14938: inst = 32'h10408000;
      14939: inst = 32'hc404fa2;
      14940: inst = 32'h8220000;
      14941: inst = 32'h10408000;
      14942: inst = 32'hc404fa3;
      14943: inst = 32'h8220000;
      14944: inst = 32'h10408000;
      14945: inst = 32'hc404fa4;
      14946: inst = 32'h8220000;
      14947: inst = 32'h10408000;
      14948: inst = 32'hc404fa5;
      14949: inst = 32'h8220000;
      14950: inst = 32'h10408000;
      14951: inst = 32'hc404fa6;
      14952: inst = 32'h8220000;
      14953: inst = 32'h10408000;
      14954: inst = 32'hc404fa7;
      14955: inst = 32'h8220000;
      14956: inst = 32'h10408000;
      14957: inst = 32'hc404fa9;
      14958: inst = 32'h8220000;
      14959: inst = 32'h10408000;
      14960: inst = 32'hc404fab;
      14961: inst = 32'h8220000;
      14962: inst = 32'h10408000;
      14963: inst = 32'hc404fad;
      14964: inst = 32'h8220000;
      14965: inst = 32'h10408000;
      14966: inst = 32'hc404fae;
      14967: inst = 32'h8220000;
      14968: inst = 32'h10408000;
      14969: inst = 32'hc404faf;
      14970: inst = 32'h8220000;
      14971: inst = 32'h10408000;
      14972: inst = 32'hc404fb0;
      14973: inst = 32'h8220000;
      14974: inst = 32'h10408000;
      14975: inst = 32'hc404fb1;
      14976: inst = 32'h8220000;
      14977: inst = 32'h10408000;
      14978: inst = 32'hc404fb2;
      14979: inst = 32'h8220000;
      14980: inst = 32'h10408000;
      14981: inst = 32'hc404fb3;
      14982: inst = 32'h8220000;
      14983: inst = 32'h10408000;
      14984: inst = 32'hc405001;
      14985: inst = 32'h8220000;
      14986: inst = 32'h10408000;
      14987: inst = 32'hc405002;
      14988: inst = 32'h8220000;
      14989: inst = 32'h10408000;
      14990: inst = 32'hc405003;
      14991: inst = 32'h8220000;
      14992: inst = 32'h10408000;
      14993: inst = 32'hc405004;
      14994: inst = 32'h8220000;
      14995: inst = 32'h10408000;
      14996: inst = 32'hc405005;
      14997: inst = 32'h8220000;
      14998: inst = 32'h10408000;
      14999: inst = 32'hc405006;
      15000: inst = 32'h8220000;
      15001: inst = 32'h10408000;
      15002: inst = 32'hc405007;
      15003: inst = 32'h8220000;
      15004: inst = 32'h10408000;
      15005: inst = 32'hc405009;
      15006: inst = 32'h8220000;
      15007: inst = 32'h10408000;
      15008: inst = 32'hc40500b;
      15009: inst = 32'h8220000;
      15010: inst = 32'h10408000;
      15011: inst = 32'hc40500d;
      15012: inst = 32'h8220000;
      15013: inst = 32'h10408000;
      15014: inst = 32'hc40500e;
      15015: inst = 32'h8220000;
      15016: inst = 32'h10408000;
      15017: inst = 32'hc40500f;
      15018: inst = 32'h8220000;
      15019: inst = 32'h10408000;
      15020: inst = 32'hc405010;
      15021: inst = 32'h8220000;
      15022: inst = 32'h10408000;
      15023: inst = 32'hc405011;
      15024: inst = 32'h8220000;
      15025: inst = 32'h10408000;
      15026: inst = 32'hc405012;
      15027: inst = 32'h8220000;
      15028: inst = 32'h10408000;
      15029: inst = 32'hc405013;
      15030: inst = 32'h8220000;
      15031: inst = 32'h10408000;
      15032: inst = 32'hc405061;
      15033: inst = 32'h8220000;
      15034: inst = 32'h10408000;
      15035: inst = 32'hc405062;
      15036: inst = 32'h8220000;
      15037: inst = 32'h10408000;
      15038: inst = 32'hc405063;
      15039: inst = 32'h8220000;
      15040: inst = 32'h10408000;
      15041: inst = 32'hc405064;
      15042: inst = 32'h8220000;
      15043: inst = 32'h10408000;
      15044: inst = 32'hc405065;
      15045: inst = 32'h8220000;
      15046: inst = 32'h10408000;
      15047: inst = 32'hc405066;
      15048: inst = 32'h8220000;
      15049: inst = 32'h10408000;
      15050: inst = 32'hc405067;
      15051: inst = 32'h8220000;
      15052: inst = 32'h10408000;
      15053: inst = 32'hc405068;
      15054: inst = 32'h8220000;
      15055: inst = 32'h10408000;
      15056: inst = 32'hc405069;
      15057: inst = 32'h8220000;
      15058: inst = 32'h10408000;
      15059: inst = 32'hc40506b;
      15060: inst = 32'h8220000;
      15061: inst = 32'h10408000;
      15062: inst = 32'hc40506c;
      15063: inst = 32'h8220000;
      15064: inst = 32'h10408000;
      15065: inst = 32'hc40506d;
      15066: inst = 32'h8220000;
      15067: inst = 32'h10408000;
      15068: inst = 32'hc40506e;
      15069: inst = 32'h8220000;
      15070: inst = 32'h10408000;
      15071: inst = 32'hc40506f;
      15072: inst = 32'h8220000;
      15073: inst = 32'h10408000;
      15074: inst = 32'hc405070;
      15075: inst = 32'h8220000;
      15076: inst = 32'h10408000;
      15077: inst = 32'hc405071;
      15078: inst = 32'h8220000;
      15079: inst = 32'h10408000;
      15080: inst = 32'hc405072;
      15081: inst = 32'h8220000;
      15082: inst = 32'h10408000;
      15083: inst = 32'hc405073;
      15084: inst = 32'h8220000;
      15085: inst = 32'h10408000;
      15086: inst = 32'hc4050c1;
      15087: inst = 32'h8220000;
      15088: inst = 32'h10408000;
      15089: inst = 32'hc4050c2;
      15090: inst = 32'h8220000;
      15091: inst = 32'h10408000;
      15092: inst = 32'hc4050c3;
      15093: inst = 32'h8220000;
      15094: inst = 32'h10408000;
      15095: inst = 32'hc4050c4;
      15096: inst = 32'h8220000;
      15097: inst = 32'h10408000;
      15098: inst = 32'hc4050c5;
      15099: inst = 32'h8220000;
      15100: inst = 32'h10408000;
      15101: inst = 32'hc4050c6;
      15102: inst = 32'h8220000;
      15103: inst = 32'h10408000;
      15104: inst = 32'hc4050c7;
      15105: inst = 32'h8220000;
      15106: inst = 32'h10408000;
      15107: inst = 32'hc4050c8;
      15108: inst = 32'h8220000;
      15109: inst = 32'h10408000;
      15110: inst = 32'hc4050c9;
      15111: inst = 32'h8220000;
      15112: inst = 32'h10408000;
      15113: inst = 32'hc4050cb;
      15114: inst = 32'h8220000;
      15115: inst = 32'h10408000;
      15116: inst = 32'hc4050cc;
      15117: inst = 32'h8220000;
      15118: inst = 32'h10408000;
      15119: inst = 32'hc4050cd;
      15120: inst = 32'h8220000;
      15121: inst = 32'h10408000;
      15122: inst = 32'hc4050ce;
      15123: inst = 32'h8220000;
      15124: inst = 32'h10408000;
      15125: inst = 32'hc4050cf;
      15126: inst = 32'h8220000;
      15127: inst = 32'h10408000;
      15128: inst = 32'hc4050d0;
      15129: inst = 32'h8220000;
      15130: inst = 32'h10408000;
      15131: inst = 32'hc4050d1;
      15132: inst = 32'h8220000;
      15133: inst = 32'h10408000;
      15134: inst = 32'hc4050d2;
      15135: inst = 32'h8220000;
      15136: inst = 32'h10408000;
      15137: inst = 32'hc4050d3;
      15138: inst = 32'h8220000;
      15139: inst = 32'h10408000;
      15140: inst = 32'hc405121;
      15141: inst = 32'h8220000;
      15142: inst = 32'h10408000;
      15143: inst = 32'hc405122;
      15144: inst = 32'h8220000;
      15145: inst = 32'h10408000;
      15146: inst = 32'hc405123;
      15147: inst = 32'h8220000;
      15148: inst = 32'h10408000;
      15149: inst = 32'hc405124;
      15150: inst = 32'h8220000;
      15151: inst = 32'h10408000;
      15152: inst = 32'hc405125;
      15153: inst = 32'h8220000;
      15154: inst = 32'h10408000;
      15155: inst = 32'hc405126;
      15156: inst = 32'h8220000;
      15157: inst = 32'h10408000;
      15158: inst = 32'hc405127;
      15159: inst = 32'h8220000;
      15160: inst = 32'h10408000;
      15161: inst = 32'hc405128;
      15162: inst = 32'h8220000;
      15163: inst = 32'h10408000;
      15164: inst = 32'hc405129;
      15165: inst = 32'h8220000;
      15166: inst = 32'h10408000;
      15167: inst = 32'hc40512b;
      15168: inst = 32'h8220000;
      15169: inst = 32'h10408000;
      15170: inst = 32'hc40512c;
      15171: inst = 32'h8220000;
      15172: inst = 32'h10408000;
      15173: inst = 32'hc40512d;
      15174: inst = 32'h8220000;
      15175: inst = 32'h10408000;
      15176: inst = 32'hc40512e;
      15177: inst = 32'h8220000;
      15178: inst = 32'h10408000;
      15179: inst = 32'hc40512f;
      15180: inst = 32'h8220000;
      15181: inst = 32'h10408000;
      15182: inst = 32'hc405130;
      15183: inst = 32'h8220000;
      15184: inst = 32'h10408000;
      15185: inst = 32'hc405131;
      15186: inst = 32'h8220000;
      15187: inst = 32'h10408000;
      15188: inst = 32'hc405132;
      15189: inst = 32'h8220000;
      15190: inst = 32'h10408000;
      15191: inst = 32'hc405133;
      15192: inst = 32'h8220000;
      15193: inst = 32'h10408000;
      15194: inst = 32'hc405181;
      15195: inst = 32'h8220000;
      15196: inst = 32'h10408000;
      15197: inst = 32'hc405182;
      15198: inst = 32'h8220000;
      15199: inst = 32'h10408000;
      15200: inst = 32'hc405183;
      15201: inst = 32'h8220000;
      15202: inst = 32'h10408000;
      15203: inst = 32'hc405184;
      15204: inst = 32'h8220000;
      15205: inst = 32'h10408000;
      15206: inst = 32'hc405185;
      15207: inst = 32'h8220000;
      15208: inst = 32'h10408000;
      15209: inst = 32'hc405186;
      15210: inst = 32'h8220000;
      15211: inst = 32'h10408000;
      15212: inst = 32'hc405187;
      15213: inst = 32'h8220000;
      15214: inst = 32'h10408000;
      15215: inst = 32'hc405188;
      15216: inst = 32'h8220000;
      15217: inst = 32'h10408000;
      15218: inst = 32'hc405189;
      15219: inst = 32'h8220000;
      15220: inst = 32'h10408000;
      15221: inst = 32'hc40518b;
      15222: inst = 32'h8220000;
      15223: inst = 32'h10408000;
      15224: inst = 32'hc40518c;
      15225: inst = 32'h8220000;
      15226: inst = 32'h10408000;
      15227: inst = 32'hc40518d;
      15228: inst = 32'h8220000;
      15229: inst = 32'h10408000;
      15230: inst = 32'hc40518e;
      15231: inst = 32'h8220000;
      15232: inst = 32'h10408000;
      15233: inst = 32'hc40518f;
      15234: inst = 32'h8220000;
      15235: inst = 32'h10408000;
      15236: inst = 32'hc405190;
      15237: inst = 32'h8220000;
      15238: inst = 32'h10408000;
      15239: inst = 32'hc405191;
      15240: inst = 32'h8220000;
      15241: inst = 32'h10408000;
      15242: inst = 32'hc405192;
      15243: inst = 32'h8220000;
      15244: inst = 32'h10408000;
      15245: inst = 32'hc405193;
      15246: inst = 32'h8220000;
      15247: inst = 32'h10408000;
      15248: inst = 32'hc4051e1;
      15249: inst = 32'h8220000;
      15250: inst = 32'h10408000;
      15251: inst = 32'hc4051e2;
      15252: inst = 32'h8220000;
      15253: inst = 32'h10408000;
      15254: inst = 32'hc4051e3;
      15255: inst = 32'h8220000;
      15256: inst = 32'h10408000;
      15257: inst = 32'hc4051e4;
      15258: inst = 32'h8220000;
      15259: inst = 32'h10408000;
      15260: inst = 32'hc4051e5;
      15261: inst = 32'h8220000;
      15262: inst = 32'h10408000;
      15263: inst = 32'hc4051e6;
      15264: inst = 32'h8220000;
      15265: inst = 32'h10408000;
      15266: inst = 32'hc4051e7;
      15267: inst = 32'h8220000;
      15268: inst = 32'h10408000;
      15269: inst = 32'hc4051e8;
      15270: inst = 32'h8220000;
      15271: inst = 32'h10408000;
      15272: inst = 32'hc4051e9;
      15273: inst = 32'h8220000;
      15274: inst = 32'h10408000;
      15275: inst = 32'hc4051eb;
      15276: inst = 32'h8220000;
      15277: inst = 32'h10408000;
      15278: inst = 32'hc4051ec;
      15279: inst = 32'h8220000;
      15280: inst = 32'h10408000;
      15281: inst = 32'hc4051ed;
      15282: inst = 32'h8220000;
      15283: inst = 32'h10408000;
      15284: inst = 32'hc4051ee;
      15285: inst = 32'h8220000;
      15286: inst = 32'h10408000;
      15287: inst = 32'hc4051ef;
      15288: inst = 32'h8220000;
      15289: inst = 32'h10408000;
      15290: inst = 32'hc4051f0;
      15291: inst = 32'h8220000;
      15292: inst = 32'h10408000;
      15293: inst = 32'hc4051f1;
      15294: inst = 32'h8220000;
      15295: inst = 32'h10408000;
      15296: inst = 32'hc4051f2;
      15297: inst = 32'h8220000;
      15298: inst = 32'h10408000;
      15299: inst = 32'hc4051f3;
      15300: inst = 32'h8220000;
      15301: inst = 32'h10408000;
      15302: inst = 32'hc405241;
      15303: inst = 32'h8220000;
      15304: inst = 32'h10408000;
      15305: inst = 32'hc405242;
      15306: inst = 32'h8220000;
      15307: inst = 32'h10408000;
      15308: inst = 32'hc405243;
      15309: inst = 32'h8220000;
      15310: inst = 32'h10408000;
      15311: inst = 32'hc405244;
      15312: inst = 32'h8220000;
      15313: inst = 32'h10408000;
      15314: inst = 32'hc405245;
      15315: inst = 32'h8220000;
      15316: inst = 32'h10408000;
      15317: inst = 32'hc405246;
      15318: inst = 32'h8220000;
      15319: inst = 32'h10408000;
      15320: inst = 32'hc405247;
      15321: inst = 32'h8220000;
      15322: inst = 32'h10408000;
      15323: inst = 32'hc405248;
      15324: inst = 32'h8220000;
      15325: inst = 32'h10408000;
      15326: inst = 32'hc405249;
      15327: inst = 32'h8220000;
      15328: inst = 32'h10408000;
      15329: inst = 32'hc40524b;
      15330: inst = 32'h8220000;
      15331: inst = 32'h10408000;
      15332: inst = 32'hc40524c;
      15333: inst = 32'h8220000;
      15334: inst = 32'h10408000;
      15335: inst = 32'hc40524d;
      15336: inst = 32'h8220000;
      15337: inst = 32'h10408000;
      15338: inst = 32'hc40524e;
      15339: inst = 32'h8220000;
      15340: inst = 32'h10408000;
      15341: inst = 32'hc40524f;
      15342: inst = 32'h8220000;
      15343: inst = 32'h10408000;
      15344: inst = 32'hc405250;
      15345: inst = 32'h8220000;
      15346: inst = 32'h10408000;
      15347: inst = 32'hc405251;
      15348: inst = 32'h8220000;
      15349: inst = 32'h10408000;
      15350: inst = 32'hc405252;
      15351: inst = 32'h8220000;
      15352: inst = 32'h10408000;
      15353: inst = 32'hc405253;
      15354: inst = 32'h8220000;
      15355: inst = 32'hc20bd73;
      15356: inst = 32'h10408000;
      15357: inst = 32'hc404e9f;
      15358: inst = 32'h8220000;
      15359: inst = 32'h10408000;
      15360: inst = 32'hc404ec0;
      15361: inst = 32'h8220000;
      15362: inst = 32'hc205aed;
      15363: inst = 32'h10408000;
      15364: inst = 32'hc404ea0;
      15365: inst = 32'h8220000;
      15366: inst = 32'h10408000;
      15367: inst = 32'hc404ea1;
      15368: inst = 32'h8220000;
      15369: inst = 32'h10408000;
      15370: inst = 32'hc404ea2;
      15371: inst = 32'h8220000;
      15372: inst = 32'h10408000;
      15373: inst = 32'hc404ea3;
      15374: inst = 32'h8220000;
      15375: inst = 32'h10408000;
      15376: inst = 32'hc404ea4;
      15377: inst = 32'h8220000;
      15378: inst = 32'h10408000;
      15379: inst = 32'hc404ebb;
      15380: inst = 32'h8220000;
      15381: inst = 32'h10408000;
      15382: inst = 32'hc404ebc;
      15383: inst = 32'h8220000;
      15384: inst = 32'h10408000;
      15385: inst = 32'hc404ebd;
      15386: inst = 32'h8220000;
      15387: inst = 32'h10408000;
      15388: inst = 32'hc404ebe;
      15389: inst = 32'h8220000;
      15390: inst = 32'h10408000;
      15391: inst = 32'hc404ebf;
      15392: inst = 32'h8220000;
      15393: inst = 32'h10408000;
      15394: inst = 32'hc404f00;
      15395: inst = 32'h8220000;
      15396: inst = 32'h10408000;
      15397: inst = 32'hc404f01;
      15398: inst = 32'h8220000;
      15399: inst = 32'h10408000;
      15400: inst = 32'hc404f02;
      15401: inst = 32'h8220000;
      15402: inst = 32'h10408000;
      15403: inst = 32'hc404f03;
      15404: inst = 32'h8220000;
      15405: inst = 32'h10408000;
      15406: inst = 32'hc404f04;
      15407: inst = 32'h8220000;
      15408: inst = 32'h10408000;
      15409: inst = 32'hc404f05;
      15410: inst = 32'h8220000;
      15411: inst = 32'h10408000;
      15412: inst = 32'hc404f1a;
      15413: inst = 32'h8220000;
      15414: inst = 32'h10408000;
      15415: inst = 32'hc404f1b;
      15416: inst = 32'h8220000;
      15417: inst = 32'h10408000;
      15418: inst = 32'hc404f1c;
      15419: inst = 32'h8220000;
      15420: inst = 32'h10408000;
      15421: inst = 32'hc404f1d;
      15422: inst = 32'h8220000;
      15423: inst = 32'h10408000;
      15424: inst = 32'hc404f1e;
      15425: inst = 32'h8220000;
      15426: inst = 32'h10408000;
      15427: inst = 32'hc404f1f;
      15428: inst = 32'h8220000;
      15429: inst = 32'h10408000;
      15430: inst = 32'hc404f60;
      15431: inst = 32'h8220000;
      15432: inst = 32'h10408000;
      15433: inst = 32'hc404f61;
      15434: inst = 32'h8220000;
      15435: inst = 32'h10408000;
      15436: inst = 32'hc404f62;
      15437: inst = 32'h8220000;
      15438: inst = 32'h10408000;
      15439: inst = 32'hc404f63;
      15440: inst = 32'h8220000;
      15441: inst = 32'h10408000;
      15442: inst = 32'hc404f64;
      15443: inst = 32'h8220000;
      15444: inst = 32'h10408000;
      15445: inst = 32'hc404f65;
      15446: inst = 32'h8220000;
      15447: inst = 32'h10408000;
      15448: inst = 32'hc404f66;
      15449: inst = 32'h8220000;
      15450: inst = 32'h10408000;
      15451: inst = 32'hc404f67;
      15452: inst = 32'h8220000;
      15453: inst = 32'h10408000;
      15454: inst = 32'hc404f78;
      15455: inst = 32'h8220000;
      15456: inst = 32'h10408000;
      15457: inst = 32'hc404f79;
      15458: inst = 32'h8220000;
      15459: inst = 32'h10408000;
      15460: inst = 32'hc404f7a;
      15461: inst = 32'h8220000;
      15462: inst = 32'h10408000;
      15463: inst = 32'hc404f7b;
      15464: inst = 32'h8220000;
      15465: inst = 32'h10408000;
      15466: inst = 32'hc404f7c;
      15467: inst = 32'h8220000;
      15468: inst = 32'h10408000;
      15469: inst = 32'hc404f7d;
      15470: inst = 32'h8220000;
      15471: inst = 32'h10408000;
      15472: inst = 32'hc404f7e;
      15473: inst = 32'h8220000;
      15474: inst = 32'h10408000;
      15475: inst = 32'hc404f7f;
      15476: inst = 32'h8220000;
      15477: inst = 32'h10408000;
      15478: inst = 32'hc404fc0;
      15479: inst = 32'h8220000;
      15480: inst = 32'h10408000;
      15481: inst = 32'hc404fc1;
      15482: inst = 32'h8220000;
      15483: inst = 32'h10408000;
      15484: inst = 32'hc404fc2;
      15485: inst = 32'h8220000;
      15486: inst = 32'h10408000;
      15487: inst = 32'hc404fc3;
      15488: inst = 32'h8220000;
      15489: inst = 32'h10408000;
      15490: inst = 32'hc404fc4;
      15491: inst = 32'h8220000;
      15492: inst = 32'h10408000;
      15493: inst = 32'hc404fc6;
      15494: inst = 32'h8220000;
      15495: inst = 32'h10408000;
      15496: inst = 32'hc404fc7;
      15497: inst = 32'h8220000;
      15498: inst = 32'h10408000;
      15499: inst = 32'hc404fd8;
      15500: inst = 32'h8220000;
      15501: inst = 32'h10408000;
      15502: inst = 32'hc404fd9;
      15503: inst = 32'h8220000;
      15504: inst = 32'h10408000;
      15505: inst = 32'hc404fdb;
      15506: inst = 32'h8220000;
      15507: inst = 32'h10408000;
      15508: inst = 32'hc404fdc;
      15509: inst = 32'h8220000;
      15510: inst = 32'h10408000;
      15511: inst = 32'hc404fdd;
      15512: inst = 32'h8220000;
      15513: inst = 32'h10408000;
      15514: inst = 32'hc404fde;
      15515: inst = 32'h8220000;
      15516: inst = 32'h10408000;
      15517: inst = 32'hc404fdf;
      15518: inst = 32'h8220000;
      15519: inst = 32'h10408000;
      15520: inst = 32'hc405020;
      15521: inst = 32'h8220000;
      15522: inst = 32'h10408000;
      15523: inst = 32'hc405021;
      15524: inst = 32'h8220000;
      15525: inst = 32'h10408000;
      15526: inst = 32'hc405022;
      15527: inst = 32'h8220000;
      15528: inst = 32'h10408000;
      15529: inst = 32'hc405023;
      15530: inst = 32'h8220000;
      15531: inst = 32'h10408000;
      15532: inst = 32'hc405026;
      15533: inst = 32'h8220000;
      15534: inst = 32'h10408000;
      15535: inst = 32'hc405027;
      15536: inst = 32'h8220000;
      15537: inst = 32'h10408000;
      15538: inst = 32'hc405038;
      15539: inst = 32'h8220000;
      15540: inst = 32'h10408000;
      15541: inst = 32'hc405039;
      15542: inst = 32'h8220000;
      15543: inst = 32'h10408000;
      15544: inst = 32'hc40503c;
      15545: inst = 32'h8220000;
      15546: inst = 32'h10408000;
      15547: inst = 32'hc40503d;
      15548: inst = 32'h8220000;
      15549: inst = 32'h10408000;
      15550: inst = 32'hc40503e;
      15551: inst = 32'h8220000;
      15552: inst = 32'h10408000;
      15553: inst = 32'hc40503f;
      15554: inst = 32'h8220000;
      15555: inst = 32'h10408000;
      15556: inst = 32'hc40507f;
      15557: inst = 32'h8220000;
      15558: inst = 32'h10408000;
      15559: inst = 32'hc405080;
      15560: inst = 32'h8220000;
      15561: inst = 32'h10408000;
      15562: inst = 32'hc405081;
      15563: inst = 32'h8220000;
      15564: inst = 32'h10408000;
      15565: inst = 32'hc405082;
      15566: inst = 32'h8220000;
      15567: inst = 32'h10408000;
      15568: inst = 32'hc405086;
      15569: inst = 32'h8220000;
      15570: inst = 32'h10408000;
      15571: inst = 32'hc405087;
      15572: inst = 32'h8220000;
      15573: inst = 32'h10408000;
      15574: inst = 32'hc405098;
      15575: inst = 32'h8220000;
      15576: inst = 32'h10408000;
      15577: inst = 32'hc405099;
      15578: inst = 32'h8220000;
      15579: inst = 32'h10408000;
      15580: inst = 32'hc40509d;
      15581: inst = 32'h8220000;
      15582: inst = 32'h10408000;
      15583: inst = 32'hc40509e;
      15584: inst = 32'h8220000;
      15585: inst = 32'h10408000;
      15586: inst = 32'hc40509f;
      15587: inst = 32'h8220000;
      15588: inst = 32'h10408000;
      15589: inst = 32'hc4050a0;
      15590: inst = 32'h8220000;
      15591: inst = 32'h10408000;
      15592: inst = 32'hc4050df;
      15593: inst = 32'h8220000;
      15594: inst = 32'h10408000;
      15595: inst = 32'hc4050e0;
      15596: inst = 32'h8220000;
      15597: inst = 32'h10408000;
      15598: inst = 32'hc4050e1;
      15599: inst = 32'h8220000;
      15600: inst = 32'h10408000;
      15601: inst = 32'hc4050e2;
      15602: inst = 32'h8220000;
      15603: inst = 32'h10408000;
      15604: inst = 32'hc4050e6;
      15605: inst = 32'h8220000;
      15606: inst = 32'h10408000;
      15607: inst = 32'hc4050e7;
      15608: inst = 32'h8220000;
      15609: inst = 32'h10408000;
      15610: inst = 32'hc4050f8;
      15611: inst = 32'h8220000;
      15612: inst = 32'h10408000;
      15613: inst = 32'hc4050f9;
      15614: inst = 32'h8220000;
      15615: inst = 32'h10408000;
      15616: inst = 32'hc4050fd;
      15617: inst = 32'h8220000;
      15618: inst = 32'h10408000;
      15619: inst = 32'hc4050fe;
      15620: inst = 32'h8220000;
      15621: inst = 32'h10408000;
      15622: inst = 32'hc4050ff;
      15623: inst = 32'h8220000;
      15624: inst = 32'h10408000;
      15625: inst = 32'hc405100;
      15626: inst = 32'h8220000;
      15627: inst = 32'h10408000;
      15628: inst = 32'hc40513f;
      15629: inst = 32'h8220000;
      15630: inst = 32'h10408000;
      15631: inst = 32'hc405140;
      15632: inst = 32'h8220000;
      15633: inst = 32'h10408000;
      15634: inst = 32'hc405141;
      15635: inst = 32'h8220000;
      15636: inst = 32'h10408000;
      15637: inst = 32'hc405146;
      15638: inst = 32'h8220000;
      15639: inst = 32'h10408000;
      15640: inst = 32'hc405147;
      15641: inst = 32'h8220000;
      15642: inst = 32'h10408000;
      15643: inst = 32'hc405158;
      15644: inst = 32'h8220000;
      15645: inst = 32'h10408000;
      15646: inst = 32'hc405159;
      15647: inst = 32'h8220000;
      15648: inst = 32'h10408000;
      15649: inst = 32'hc40515e;
      15650: inst = 32'h8220000;
      15651: inst = 32'h10408000;
      15652: inst = 32'hc40515f;
      15653: inst = 32'h8220000;
      15654: inst = 32'h10408000;
      15655: inst = 32'hc405160;
      15656: inst = 32'h8220000;
      15657: inst = 32'h10408000;
      15658: inst = 32'hc40519f;
      15659: inst = 32'h8220000;
      15660: inst = 32'h10408000;
      15661: inst = 32'hc4051a0;
      15662: inst = 32'h8220000;
      15663: inst = 32'h10408000;
      15664: inst = 32'hc4051a6;
      15665: inst = 32'h8220000;
      15666: inst = 32'h10408000;
      15667: inst = 32'hc4051a7;
      15668: inst = 32'h8220000;
      15669: inst = 32'h10408000;
      15670: inst = 32'hc4051b8;
      15671: inst = 32'h8220000;
      15672: inst = 32'h10408000;
      15673: inst = 32'hc4051b9;
      15674: inst = 32'h8220000;
      15675: inst = 32'h10408000;
      15676: inst = 32'hc4051bf;
      15677: inst = 32'h8220000;
      15678: inst = 32'h10408000;
      15679: inst = 32'hc4051c0;
      15680: inst = 32'h8220000;
      15681: inst = 32'h10408000;
      15682: inst = 32'hc4051ff;
      15683: inst = 32'h8220000;
      15684: inst = 32'h10408000;
      15685: inst = 32'hc405200;
      15686: inst = 32'h8220000;
      15687: inst = 32'h10408000;
      15688: inst = 32'hc405206;
      15689: inst = 32'h8220000;
      15690: inst = 32'h10408000;
      15691: inst = 32'hc405207;
      15692: inst = 32'h8220000;
      15693: inst = 32'h10408000;
      15694: inst = 32'hc405218;
      15695: inst = 32'h8220000;
      15696: inst = 32'h10408000;
      15697: inst = 32'hc405219;
      15698: inst = 32'h8220000;
      15699: inst = 32'h10408000;
      15700: inst = 32'hc40521f;
      15701: inst = 32'h8220000;
      15702: inst = 32'h10408000;
      15703: inst = 32'hc405220;
      15704: inst = 32'h8220000;
      15705: inst = 32'h10408000;
      15706: inst = 32'hc40525f;
      15707: inst = 32'h8220000;
      15708: inst = 32'h10408000;
      15709: inst = 32'hc405260;
      15710: inst = 32'h8220000;
      15711: inst = 32'h10408000;
      15712: inst = 32'hc405266;
      15713: inst = 32'h8220000;
      15714: inst = 32'h10408000;
      15715: inst = 32'hc405267;
      15716: inst = 32'h8220000;
      15717: inst = 32'h10408000;
      15718: inst = 32'hc405278;
      15719: inst = 32'h8220000;
      15720: inst = 32'h10408000;
      15721: inst = 32'hc405279;
      15722: inst = 32'h8220000;
      15723: inst = 32'h10408000;
      15724: inst = 32'hc40527f;
      15725: inst = 32'h8220000;
      15726: inst = 32'h10408000;
      15727: inst = 32'hc405280;
      15728: inst = 32'h8220000;
      15729: inst = 32'h10408000;
      15730: inst = 32'hc4052bf;
      15731: inst = 32'h8220000;
      15732: inst = 32'h10408000;
      15733: inst = 32'hc4052c0;
      15734: inst = 32'h8220000;
      15735: inst = 32'h10408000;
      15736: inst = 32'hc4052c6;
      15737: inst = 32'h8220000;
      15738: inst = 32'h10408000;
      15739: inst = 32'hc4052c7;
      15740: inst = 32'h8220000;
      15741: inst = 32'h10408000;
      15742: inst = 32'hc4052d8;
      15743: inst = 32'h8220000;
      15744: inst = 32'h10408000;
      15745: inst = 32'hc4052d9;
      15746: inst = 32'h8220000;
      15747: inst = 32'h10408000;
      15748: inst = 32'hc4052df;
      15749: inst = 32'h8220000;
      15750: inst = 32'h10408000;
      15751: inst = 32'hc4052e0;
      15752: inst = 32'h8220000;
      15753: inst = 32'hc207bae;
      15754: inst = 32'h10408000;
      15755: inst = 32'hc404ea5;
      15756: inst = 32'h8220000;
      15757: inst = 32'h10408000;
      15758: inst = 32'hc404eba;
      15759: inst = 32'h8220000;
      15760: inst = 32'hc20c5b4;
      15761: inst = 32'h10408000;
      15762: inst = 32'hc404ea6;
      15763: inst = 32'h8220000;
      15764: inst = 32'h10408000;
      15765: inst = 32'hc404eb9;
      15766: inst = 32'h8220000;
      15767: inst = 32'hc20d5f4;
      15768: inst = 32'h10408000;
      15769: inst = 32'hc404ea7;
      15770: inst = 32'h8220000;
      15771: inst = 32'h10408000;
      15772: inst = 32'hc404eb8;
      15773: inst = 32'h8220000;
      15774: inst = 32'hc20a4b1;
      15775: inst = 32'h10408000;
      15776: inst = 32'hc404eff;
      15777: inst = 32'h8220000;
      15778: inst = 32'h10408000;
      15779: inst = 32'hc404f20;
      15780: inst = 32'h8220000;
      15781: inst = 32'h10408000;
      15782: inst = 32'hc404fbf;
      15783: inst = 32'h8220000;
      15784: inst = 32'h10408000;
      15785: inst = 32'hc404fe0;
      15786: inst = 32'h8220000;
      15787: inst = 32'hc2062ed;
      15788: inst = 32'h10408000;
      15789: inst = 32'hc404f06;
      15790: inst = 32'h8220000;
      15791: inst = 32'h10408000;
      15792: inst = 32'hc404f19;
      15793: inst = 32'h8220000;
      15794: inst = 32'hc209450;
      15795: inst = 32'h10408000;
      15796: inst = 32'hc404f07;
      15797: inst = 32'h8220000;
      15798: inst = 32'h10408000;
      15799: inst = 32'hc404f18;
      15800: inst = 32'h8220000;
      15801: inst = 32'h10408000;
      15802: inst = 32'hc405209;
      15803: inst = 32'h8220000;
      15804: inst = 32'h10408000;
      15805: inst = 32'hc405216;
      15806: inst = 32'h8220000;
      15807: inst = 32'hc20a4d1;
      15808: inst = 32'h10408000;
      15809: inst = 32'hc404f5f;
      15810: inst = 32'h8220000;
      15811: inst = 32'h10408000;
      15812: inst = 32'hc404f80;
      15813: inst = 32'h8220000;
      15814: inst = 32'hc204a49;
      15815: inst = 32'h10408000;
      15816: inst = 32'hc404fa8;
      15817: inst = 32'h8220000;
      15818: inst = 32'h10408000;
      15819: inst = 32'hc404fac;
      15820: inst = 32'h8220000;
      15821: inst = 32'h10408000;
      15822: inst = 32'hc405008;
      15823: inst = 32'h8220000;
      15824: inst = 32'h10408000;
      15825: inst = 32'hc40500c;
      15826: inst = 32'h8220000;
      15827: inst = 32'hc205acb;
      15828: inst = 32'h10408000;
      15829: inst = 32'hc404fc5;
      15830: inst = 32'h8220000;
      15831: inst = 32'h10408000;
      15832: inst = 32'hc404fda;
      15833: inst = 32'h8220000;
      15834: inst = 32'h10408000;
      15835: inst = 32'hc405336;
      15836: inst = 32'h8220000;
      15837: inst = 32'h10408000;
      15838: inst = 32'hc405380;
      15839: inst = 32'h8220000;
      15840: inst = 32'h10408000;
      15841: inst = 32'hc40539f;
      15842: inst = 32'h8220000;
      15843: inst = 32'h10408000;
      15844: inst = 32'hc4053dd;
      15845: inst = 32'h8220000;
      15846: inst = 32'h10408000;
      15847: inst = 32'hc405402;
      15848: inst = 32'h8220000;
      15849: inst = 32'hc20630d;
      15850: inst = 32'h10408000;
      15851: inst = 32'hc40501f;
      15852: inst = 32'h8220000;
      15853: inst = 32'h10408000;
      15854: inst = 32'hc405040;
      15855: inst = 32'h8220000;
      15856: inst = 32'hc205aec;
      15857: inst = 32'h10408000;
      15858: inst = 32'hc405024;
      15859: inst = 32'h8220000;
      15860: inst = 32'h10408000;
      15861: inst = 32'hc40503b;
      15862: inst = 32'h8220000;
      15863: inst = 32'h10408000;
      15864: inst = 32'hc405083;
      15865: inst = 32'h8220000;
      15866: inst = 32'h10408000;
      15867: inst = 32'hc40509c;
      15868: inst = 32'h8220000;
      15869: inst = 32'h10408000;
      15870: inst = 32'hc4051a1;
      15871: inst = 32'h8220000;
      15872: inst = 32'h10408000;
      15873: inst = 32'hc4051be;
      15874: inst = 32'h8220000;
      15875: inst = 32'h10408000;
      15876: inst = 32'hc405329;
      15877: inst = 32'h8220000;
      15878: inst = 32'h10408000;
      15879: inst = 32'hc405568;
      15880: inst = 32'h8220000;
      15881: inst = 32'h10408000;
      15882: inst = 32'hc405577;
      15883: inst = 32'h8220000;
      15884: inst = 32'h10408000;
      15885: inst = 32'hc4057a7;
      15886: inst = 32'h8220000;
      15887: inst = 32'h10408000;
      15888: inst = 32'hc4057b8;
      15889: inst = 32'h8220000;
      15890: inst = 32'hc205269;
      15891: inst = 32'h10408000;
      15892: inst = 32'hc405025;
      15893: inst = 32'h8220000;
      15894: inst = 32'h10408000;
      15895: inst = 32'hc40503a;
      15896: inst = 32'h8220000;
      15897: inst = 32'h10408000;
      15898: inst = 32'hc40537e;
      15899: inst = 32'h8220000;
      15900: inst = 32'h10408000;
      15901: inst = 32'hc4053a1;
      15902: inst = 32'h8220000;
      15903: inst = 32'h10408000;
      15904: inst = 32'hc40549c;
      15905: inst = 32'h8220000;
      15906: inst = 32'h10408000;
      15907: inst = 32'hc4054c3;
      15908: inst = 32'h8220000;
      15909: inst = 32'hc20528a;
      15910: inst = 32'h10408000;
      15911: inst = 32'hc405084;
      15912: inst = 32'h8220000;
      15913: inst = 32'h10408000;
      15914: inst = 32'hc40509b;
      15915: inst = 32'h8220000;
      15916: inst = 32'h10408000;
      15917: inst = 32'hc4050e3;
      15918: inst = 32'h8220000;
      15919: inst = 32'h10408000;
      15920: inst = 32'hc4050fc;
      15921: inst = 32'h8220000;
      15922: inst = 32'h10408000;
      15923: inst = 32'hc4052c5;
      15924: inst = 32'h8220000;
      15925: inst = 32'h10408000;
      15926: inst = 32'hc4052da;
      15927: inst = 32'h8220000;
      15928: inst = 32'h10408000;
      15929: inst = 32'hc4053e9;
      15930: inst = 32'h8220000;
      15931: inst = 32'h10408000;
      15932: inst = 32'hc4053f6;
      15933: inst = 32'h8220000;
      15934: inst = 32'h10408000;
      15935: inst = 32'hc405449;
      15936: inst = 32'h8220000;
      15937: inst = 32'h10408000;
      15938: inst = 32'hc405456;
      15939: inst = 32'h8220000;
      15940: inst = 32'h10408000;
      15941: inst = 32'hc4054a9;
      15942: inst = 32'h8220000;
      15943: inst = 32'h10408000;
      15944: inst = 32'hc4054b6;
      15945: inst = 32'h8220000;
      15946: inst = 32'h10408000;
      15947: inst = 32'hc405509;
      15948: inst = 32'h8220000;
      15949: inst = 32'h10408000;
      15950: inst = 32'hc405516;
      15951: inst = 32'h8220000;
      15952: inst = 32'h10408000;
      15953: inst = 32'hc40555e;
      15954: inst = 32'h8220000;
      15955: inst = 32'h10408000;
      15956: inst = 32'hc405569;
      15957: inst = 32'h8220000;
      15958: inst = 32'h10408000;
      15959: inst = 32'hc405576;
      15960: inst = 32'h8220000;
      15961: inst = 32'h10408000;
      15962: inst = 32'hc405581;
      15963: inst = 32'h8220000;
      15964: inst = 32'h10408000;
      15965: inst = 32'hc4055c9;
      15966: inst = 32'h8220000;
      15967: inst = 32'h10408000;
      15968: inst = 32'hc4055d6;
      15969: inst = 32'h8220000;
      15970: inst = 32'h10408000;
      15971: inst = 32'hc405628;
      15972: inst = 32'h8220000;
      15973: inst = 32'h10408000;
      15974: inst = 32'hc405629;
      15975: inst = 32'h8220000;
      15976: inst = 32'h10408000;
      15977: inst = 32'hc405636;
      15978: inst = 32'h8220000;
      15979: inst = 32'h10408000;
      15980: inst = 32'hc405637;
      15981: inst = 32'h8220000;
      15982: inst = 32'h10408000;
      15983: inst = 32'hc40567d;
      15984: inst = 32'h8220000;
      15985: inst = 32'h10408000;
      15986: inst = 32'hc405688;
      15987: inst = 32'h8220000;
      15988: inst = 32'h10408000;
      15989: inst = 32'hc405689;
      15990: inst = 32'h8220000;
      15991: inst = 32'h10408000;
      15992: inst = 32'hc405696;
      15993: inst = 32'h8220000;
      15994: inst = 32'h10408000;
      15995: inst = 32'hc405697;
      15996: inst = 32'h8220000;
      15997: inst = 32'h10408000;
      15998: inst = 32'hc4056a2;
      15999: inst = 32'h8220000;
      16000: inst = 32'h10408000;
      16001: inst = 32'hc4056e8;
      16002: inst = 32'h8220000;
      16003: inst = 32'h10408000;
      16004: inst = 32'hc4056e9;
      16005: inst = 32'h8220000;
      16006: inst = 32'h10408000;
      16007: inst = 32'hc4056f6;
      16008: inst = 32'h8220000;
      16009: inst = 32'h10408000;
      16010: inst = 32'hc4056f7;
      16011: inst = 32'h8220000;
      16012: inst = 32'h10408000;
      16013: inst = 32'hc405748;
      16014: inst = 32'h8220000;
      16015: inst = 32'h10408000;
      16016: inst = 32'hc405749;
      16017: inst = 32'h8220000;
      16018: inst = 32'h10408000;
      16019: inst = 32'hc405756;
      16020: inst = 32'h8220000;
      16021: inst = 32'h10408000;
      16022: inst = 32'hc405757;
      16023: inst = 32'h8220000;
      16024: inst = 32'h10408000;
      16025: inst = 32'hc4057a8;
      16026: inst = 32'h8220000;
      16027: inst = 32'h10408000;
      16028: inst = 32'hc4057a9;
      16029: inst = 32'h8220000;
      16030: inst = 32'h10408000;
      16031: inst = 32'hc4057b6;
      16032: inst = 32'h8220000;
      16033: inst = 32'h10408000;
      16034: inst = 32'hc4057b7;
      16035: inst = 32'h8220000;
      16036: inst = 32'hc205aab;
      16037: inst = 32'h10408000;
      16038: inst = 32'hc405142;
      16039: inst = 32'h8220000;
      16040: inst = 32'h10408000;
      16041: inst = 32'hc40515d;
      16042: inst = 32'h8220000;
      16043: inst = 32'hc20cdd4;
      16044: inst = 32'h10408000;
      16045: inst = 32'hc40519e;
      16046: inst = 32'h8220000;
      16047: inst = 32'h10408000;
      16048: inst = 32'hc4051c1;
      16049: inst = 32'h8220000;
      16050: inst = 32'hc209471;
      16051: inst = 32'h10408000;
      16052: inst = 32'hc4051b6;
      16053: inst = 32'h8220000;
      16054: inst = 32'hc20de55;
      16055: inst = 32'h10408000;
      16056: inst = 32'hc4051fd;
      16057: inst = 32'h8220000;
      16058: inst = 32'h10408000;
      16059: inst = 32'hc405222;
      16060: inst = 32'h8220000;
      16061: inst = 32'hc209492;
      16062: inst = 32'h10408000;
      16063: inst = 32'hc4051fe;
      16064: inst = 32'h8220000;
      16065: inst = 32'h10408000;
      16066: inst = 32'hc405221;
      16067: inst = 32'h8220000;
      16068: inst = 32'hc205acc;
      16069: inst = 32'h10408000;
      16070: inst = 32'hc405201;
      16071: inst = 32'h8220000;
      16072: inst = 32'h10408000;
      16073: inst = 32'hc40521e;
      16074: inst = 32'h8220000;
      16075: inst = 32'h10408000;
      16076: inst = 32'hc405261;
      16077: inst = 32'h8220000;
      16078: inst = 32'h10408000;
      16079: inst = 32'hc40527e;
      16080: inst = 32'h8220000;
      16081: inst = 32'h10408000;
      16082: inst = 32'hc4052c1;
      16083: inst = 32'h8220000;
      16084: inst = 32'h10408000;
      16085: inst = 32'hc4052de;
      16086: inst = 32'h8220000;
      16087: inst = 32'hc20e696;
      16088: inst = 32'h10408000;
      16089: inst = 32'hc40525c;
      16090: inst = 32'h8220000;
      16091: inst = 32'h10408000;
      16092: inst = 32'hc405283;
      16093: inst = 32'h8220000;
      16094: inst = 32'hc209cb2;
      16095: inst = 32'h10408000;
      16096: inst = 32'hc40525d;
      16097: inst = 32'h8220000;
      16098: inst = 32'h10408000;
      16099: inst = 32'hc405282;
      16100: inst = 32'h8220000;
      16101: inst = 32'hc208c2f;
      16102: inst = 32'h10408000;
      16103: inst = 32'hc405269;
      16104: inst = 32'h8220000;
      16105: inst = 32'h10408000;
      16106: inst = 32'hc405276;
      16107: inst = 32'h8220000;
      16108: inst = 32'hc20ad33;
      16109: inst = 32'h10408000;
      16110: inst = 32'hc4052bc;
      16111: inst = 32'h8220000;
      16112: inst = 32'h10408000;
      16113: inst = 32'hc4052e3;
      16114: inst = 32'h8220000;
      16115: inst = 32'hc2083ee;
      16116: inst = 32'h10408000;
      16117: inst = 32'hc4052c9;
      16118: inst = 32'h8220000;
      16119: inst = 32'h10408000;
      16120: inst = 32'hc4052d6;
      16121: inst = 32'h8220000;
      16122: inst = 32'hc206b50;
      16123: inst = 32'h10408000;
      16124: inst = 32'hc405300;
      16125: inst = 32'h8220000;
      16126: inst = 32'h10408000;
      16127: inst = 32'hc405301;
      16128: inst = 32'h8220000;
      16129: inst = 32'h10408000;
      16130: inst = 32'hc405302;
      16131: inst = 32'h8220000;
      16132: inst = 32'h10408000;
      16133: inst = 32'hc405303;
      16134: inst = 32'h8220000;
      16135: inst = 32'h10408000;
      16136: inst = 32'hc405304;
      16137: inst = 32'h8220000;
      16138: inst = 32'h10408000;
      16139: inst = 32'hc405305;
      16140: inst = 32'h8220000;
      16141: inst = 32'h10408000;
      16142: inst = 32'hc405306;
      16143: inst = 32'h8220000;
      16144: inst = 32'h10408000;
      16145: inst = 32'hc405307;
      16146: inst = 32'h8220000;
      16147: inst = 32'h10408000;
      16148: inst = 32'hc405308;
      16149: inst = 32'h8220000;
      16150: inst = 32'h10408000;
      16151: inst = 32'hc405309;
      16152: inst = 32'h8220000;
      16153: inst = 32'h10408000;
      16154: inst = 32'hc40530a;
      16155: inst = 32'h8220000;
      16156: inst = 32'h10408000;
      16157: inst = 32'hc40530b;
      16158: inst = 32'h8220000;
      16159: inst = 32'h10408000;
      16160: inst = 32'hc40530c;
      16161: inst = 32'h8220000;
      16162: inst = 32'h10408000;
      16163: inst = 32'hc40530d;
      16164: inst = 32'h8220000;
      16165: inst = 32'h10408000;
      16166: inst = 32'hc40530e;
      16167: inst = 32'h8220000;
      16168: inst = 32'h10408000;
      16169: inst = 32'hc40530f;
      16170: inst = 32'h8220000;
      16171: inst = 32'h10408000;
      16172: inst = 32'hc405310;
      16173: inst = 32'h8220000;
      16174: inst = 32'h10408000;
      16175: inst = 32'hc405311;
      16176: inst = 32'h8220000;
      16177: inst = 32'h10408000;
      16178: inst = 32'hc405312;
      16179: inst = 32'h8220000;
      16180: inst = 32'h10408000;
      16181: inst = 32'hc405313;
      16182: inst = 32'h8220000;
      16183: inst = 32'h10408000;
      16184: inst = 32'hc405314;
      16185: inst = 32'h8220000;
      16186: inst = 32'h10408000;
      16187: inst = 32'hc405315;
      16188: inst = 32'h8220000;
      16189: inst = 32'h10408000;
      16190: inst = 32'hc405316;
      16191: inst = 32'h8220000;
      16192: inst = 32'h10408000;
      16193: inst = 32'hc405317;
      16194: inst = 32'h8220000;
      16195: inst = 32'h10408000;
      16196: inst = 32'hc405318;
      16197: inst = 32'h8220000;
      16198: inst = 32'h10408000;
      16199: inst = 32'hc405319;
      16200: inst = 32'h8220000;
      16201: inst = 32'h10408000;
      16202: inst = 32'hc40531a;
      16203: inst = 32'h8220000;
      16204: inst = 32'h10408000;
      16205: inst = 32'hc40532a;
      16206: inst = 32'h8220000;
      16207: inst = 32'h10408000;
      16208: inst = 32'hc40532b;
      16209: inst = 32'h8220000;
      16210: inst = 32'h10408000;
      16211: inst = 32'hc40532c;
      16212: inst = 32'h8220000;
      16213: inst = 32'h10408000;
      16214: inst = 32'hc40532d;
      16215: inst = 32'h8220000;
      16216: inst = 32'h10408000;
      16217: inst = 32'hc40532e;
      16218: inst = 32'h8220000;
      16219: inst = 32'h10408000;
      16220: inst = 32'hc40532f;
      16221: inst = 32'h8220000;
      16222: inst = 32'h10408000;
      16223: inst = 32'hc405330;
      16224: inst = 32'h8220000;
      16225: inst = 32'h10408000;
      16226: inst = 32'hc405331;
      16227: inst = 32'h8220000;
      16228: inst = 32'h10408000;
      16229: inst = 32'hc405332;
      16230: inst = 32'h8220000;
      16231: inst = 32'h10408000;
      16232: inst = 32'hc405333;
      16233: inst = 32'h8220000;
      16234: inst = 32'h10408000;
      16235: inst = 32'hc405334;
      16236: inst = 32'h8220000;
      16237: inst = 32'h10408000;
      16238: inst = 32'hc405335;
      16239: inst = 32'h8220000;
      16240: inst = 32'h10408000;
      16241: inst = 32'hc405345;
      16242: inst = 32'h8220000;
      16243: inst = 32'h10408000;
      16244: inst = 32'hc405346;
      16245: inst = 32'h8220000;
      16246: inst = 32'h10408000;
      16247: inst = 32'hc405347;
      16248: inst = 32'h8220000;
      16249: inst = 32'h10408000;
      16250: inst = 32'hc405348;
      16251: inst = 32'h8220000;
      16252: inst = 32'h10408000;
      16253: inst = 32'hc405349;
      16254: inst = 32'h8220000;
      16255: inst = 32'h10408000;
      16256: inst = 32'hc40534a;
      16257: inst = 32'h8220000;
      16258: inst = 32'h10408000;
      16259: inst = 32'hc40534b;
      16260: inst = 32'h8220000;
      16261: inst = 32'h10408000;
      16262: inst = 32'hc40534c;
      16263: inst = 32'h8220000;
      16264: inst = 32'h10408000;
      16265: inst = 32'hc40534d;
      16266: inst = 32'h8220000;
      16267: inst = 32'h10408000;
      16268: inst = 32'hc40534e;
      16269: inst = 32'h8220000;
      16270: inst = 32'h10408000;
      16271: inst = 32'hc40534f;
      16272: inst = 32'h8220000;
      16273: inst = 32'h10408000;
      16274: inst = 32'hc405350;
      16275: inst = 32'h8220000;
      16276: inst = 32'h10408000;
      16277: inst = 32'hc405351;
      16278: inst = 32'h8220000;
      16279: inst = 32'h10408000;
      16280: inst = 32'hc405352;
      16281: inst = 32'h8220000;
      16282: inst = 32'h10408000;
      16283: inst = 32'hc405353;
      16284: inst = 32'h8220000;
      16285: inst = 32'h10408000;
      16286: inst = 32'hc405354;
      16287: inst = 32'h8220000;
      16288: inst = 32'h10408000;
      16289: inst = 32'hc405355;
      16290: inst = 32'h8220000;
      16291: inst = 32'h10408000;
      16292: inst = 32'hc405356;
      16293: inst = 32'h8220000;
      16294: inst = 32'h10408000;
      16295: inst = 32'hc405357;
      16296: inst = 32'h8220000;
      16297: inst = 32'h10408000;
      16298: inst = 32'hc405358;
      16299: inst = 32'h8220000;
      16300: inst = 32'h10408000;
      16301: inst = 32'hc405359;
      16302: inst = 32'h8220000;
      16303: inst = 32'h10408000;
      16304: inst = 32'hc40535a;
      16305: inst = 32'h8220000;
      16306: inst = 32'h10408000;
      16307: inst = 32'hc40535b;
      16308: inst = 32'h8220000;
      16309: inst = 32'h10408000;
      16310: inst = 32'hc40535c;
      16311: inst = 32'h8220000;
      16312: inst = 32'h10408000;
      16313: inst = 32'hc40535d;
      16314: inst = 32'h8220000;
      16315: inst = 32'h10408000;
      16316: inst = 32'hc40535e;
      16317: inst = 32'h8220000;
      16318: inst = 32'h10408000;
      16319: inst = 32'hc40535f;
      16320: inst = 32'h8220000;
      16321: inst = 32'h10408000;
      16322: inst = 32'hc405360;
      16323: inst = 32'h8220000;
      16324: inst = 32'h10408000;
      16325: inst = 32'hc405361;
      16326: inst = 32'h8220000;
      16327: inst = 32'h10408000;
      16328: inst = 32'hc405362;
      16329: inst = 32'h8220000;
      16330: inst = 32'h10408000;
      16331: inst = 32'hc405363;
      16332: inst = 32'h8220000;
      16333: inst = 32'h10408000;
      16334: inst = 32'hc405364;
      16335: inst = 32'h8220000;
      16336: inst = 32'h10408000;
      16337: inst = 32'hc405365;
      16338: inst = 32'h8220000;
      16339: inst = 32'h10408000;
      16340: inst = 32'hc405366;
      16341: inst = 32'h8220000;
      16342: inst = 32'h10408000;
      16343: inst = 32'hc405367;
      16344: inst = 32'h8220000;
      16345: inst = 32'h10408000;
      16346: inst = 32'hc405368;
      16347: inst = 32'h8220000;
      16348: inst = 32'h10408000;
      16349: inst = 32'hc405369;
      16350: inst = 32'h8220000;
      16351: inst = 32'h10408000;
      16352: inst = 32'hc40536a;
      16353: inst = 32'h8220000;
      16354: inst = 32'h10408000;
      16355: inst = 32'hc40536b;
      16356: inst = 32'h8220000;
      16357: inst = 32'h10408000;
      16358: inst = 32'hc40536c;
      16359: inst = 32'h8220000;
      16360: inst = 32'h10408000;
      16361: inst = 32'hc40536d;
      16362: inst = 32'h8220000;
      16363: inst = 32'h10408000;
      16364: inst = 32'hc40536e;
      16365: inst = 32'h8220000;
      16366: inst = 32'h10408000;
      16367: inst = 32'hc40536f;
      16368: inst = 32'h8220000;
      16369: inst = 32'h10408000;
      16370: inst = 32'hc405370;
      16371: inst = 32'h8220000;
      16372: inst = 32'h10408000;
      16373: inst = 32'hc405371;
      16374: inst = 32'h8220000;
      16375: inst = 32'h10408000;
      16376: inst = 32'hc405372;
      16377: inst = 32'h8220000;
      16378: inst = 32'h10408000;
      16379: inst = 32'hc405373;
      16380: inst = 32'h8220000;
      16381: inst = 32'h10408000;
      16382: inst = 32'hc405374;
      16383: inst = 32'h8220000;
      16384: inst = 32'h10408000;
      16385: inst = 32'hc405375;
      16386: inst = 32'h8220000;
      16387: inst = 32'h10408000;
      16388: inst = 32'hc405376;
      16389: inst = 32'h8220000;
      16390: inst = 32'h10408000;
      16391: inst = 32'hc405377;
      16392: inst = 32'h8220000;
      16393: inst = 32'h10408000;
      16394: inst = 32'hc405378;
      16395: inst = 32'h8220000;
      16396: inst = 32'h10408000;
      16397: inst = 32'hc405379;
      16398: inst = 32'h8220000;
      16399: inst = 32'h10408000;
      16400: inst = 32'hc40538a;
      16401: inst = 32'h8220000;
      16402: inst = 32'h10408000;
      16403: inst = 32'hc40538b;
      16404: inst = 32'h8220000;
      16405: inst = 32'h10408000;
      16406: inst = 32'hc40538c;
      16407: inst = 32'h8220000;
      16408: inst = 32'h10408000;
      16409: inst = 32'hc40538d;
      16410: inst = 32'h8220000;
      16411: inst = 32'h10408000;
      16412: inst = 32'hc40538e;
      16413: inst = 32'h8220000;
      16414: inst = 32'h10408000;
      16415: inst = 32'hc40538f;
      16416: inst = 32'h8220000;
      16417: inst = 32'h10408000;
      16418: inst = 32'hc405390;
      16419: inst = 32'h8220000;
      16420: inst = 32'h10408000;
      16421: inst = 32'hc405391;
      16422: inst = 32'h8220000;
      16423: inst = 32'h10408000;
      16424: inst = 32'hc405392;
      16425: inst = 32'h8220000;
      16426: inst = 32'h10408000;
      16427: inst = 32'hc405393;
      16428: inst = 32'h8220000;
      16429: inst = 32'h10408000;
      16430: inst = 32'hc405394;
      16431: inst = 32'h8220000;
      16432: inst = 32'h10408000;
      16433: inst = 32'hc405395;
      16434: inst = 32'h8220000;
      16435: inst = 32'h10408000;
      16436: inst = 32'hc4053a6;
      16437: inst = 32'h8220000;
      16438: inst = 32'h10408000;
      16439: inst = 32'hc4053a7;
      16440: inst = 32'h8220000;
      16441: inst = 32'h10408000;
      16442: inst = 32'hc4053a8;
      16443: inst = 32'h8220000;
      16444: inst = 32'h10408000;
      16445: inst = 32'hc4053a9;
      16446: inst = 32'h8220000;
      16447: inst = 32'h10408000;
      16448: inst = 32'hc4053aa;
      16449: inst = 32'h8220000;
      16450: inst = 32'h10408000;
      16451: inst = 32'hc4053ab;
      16452: inst = 32'h8220000;
      16453: inst = 32'h10408000;
      16454: inst = 32'hc4053ac;
      16455: inst = 32'h8220000;
      16456: inst = 32'h10408000;
      16457: inst = 32'hc4053ad;
      16458: inst = 32'h8220000;
      16459: inst = 32'h10408000;
      16460: inst = 32'hc4053ae;
      16461: inst = 32'h8220000;
      16462: inst = 32'h10408000;
      16463: inst = 32'hc4053af;
      16464: inst = 32'h8220000;
      16465: inst = 32'h10408000;
      16466: inst = 32'hc4053b0;
      16467: inst = 32'h8220000;
      16468: inst = 32'h10408000;
      16469: inst = 32'hc4053b1;
      16470: inst = 32'h8220000;
      16471: inst = 32'h10408000;
      16472: inst = 32'hc4053b2;
      16473: inst = 32'h8220000;
      16474: inst = 32'h10408000;
      16475: inst = 32'hc4053b3;
      16476: inst = 32'h8220000;
      16477: inst = 32'h10408000;
      16478: inst = 32'hc4053b4;
      16479: inst = 32'h8220000;
      16480: inst = 32'h10408000;
      16481: inst = 32'hc4053b5;
      16482: inst = 32'h8220000;
      16483: inst = 32'h10408000;
      16484: inst = 32'hc4053b6;
      16485: inst = 32'h8220000;
      16486: inst = 32'h10408000;
      16487: inst = 32'hc4053b7;
      16488: inst = 32'h8220000;
      16489: inst = 32'h10408000;
      16490: inst = 32'hc4053b8;
      16491: inst = 32'h8220000;
      16492: inst = 32'h10408000;
      16493: inst = 32'hc4053b9;
      16494: inst = 32'h8220000;
      16495: inst = 32'h10408000;
      16496: inst = 32'hc4053ba;
      16497: inst = 32'h8220000;
      16498: inst = 32'h10408000;
      16499: inst = 32'hc4053bb;
      16500: inst = 32'h8220000;
      16501: inst = 32'h10408000;
      16502: inst = 32'hc4053bc;
      16503: inst = 32'h8220000;
      16504: inst = 32'h10408000;
      16505: inst = 32'hc4053bd;
      16506: inst = 32'h8220000;
      16507: inst = 32'h10408000;
      16508: inst = 32'hc4053be;
      16509: inst = 32'h8220000;
      16510: inst = 32'h10408000;
      16511: inst = 32'hc4053bf;
      16512: inst = 32'h8220000;
      16513: inst = 32'h10408000;
      16514: inst = 32'hc4053c0;
      16515: inst = 32'h8220000;
      16516: inst = 32'h10408000;
      16517: inst = 32'hc4053c1;
      16518: inst = 32'h8220000;
      16519: inst = 32'h10408000;
      16520: inst = 32'hc4053c2;
      16521: inst = 32'h8220000;
      16522: inst = 32'h10408000;
      16523: inst = 32'hc4053c3;
      16524: inst = 32'h8220000;
      16525: inst = 32'h10408000;
      16526: inst = 32'hc4053c4;
      16527: inst = 32'h8220000;
      16528: inst = 32'h10408000;
      16529: inst = 32'hc4053c5;
      16530: inst = 32'h8220000;
      16531: inst = 32'h10408000;
      16532: inst = 32'hc4053c6;
      16533: inst = 32'h8220000;
      16534: inst = 32'h10408000;
      16535: inst = 32'hc4053c7;
      16536: inst = 32'h8220000;
      16537: inst = 32'h10408000;
      16538: inst = 32'hc4053c8;
      16539: inst = 32'h8220000;
      16540: inst = 32'h10408000;
      16541: inst = 32'hc4053c9;
      16542: inst = 32'h8220000;
      16543: inst = 32'h10408000;
      16544: inst = 32'hc4053ca;
      16545: inst = 32'h8220000;
      16546: inst = 32'h10408000;
      16547: inst = 32'hc4053cb;
      16548: inst = 32'h8220000;
      16549: inst = 32'h10408000;
      16550: inst = 32'hc4053cc;
      16551: inst = 32'h8220000;
      16552: inst = 32'h10408000;
      16553: inst = 32'hc4053cd;
      16554: inst = 32'h8220000;
      16555: inst = 32'h10408000;
      16556: inst = 32'hc4053ce;
      16557: inst = 32'h8220000;
      16558: inst = 32'h10408000;
      16559: inst = 32'hc4053cf;
      16560: inst = 32'h8220000;
      16561: inst = 32'h10408000;
      16562: inst = 32'hc4053d0;
      16563: inst = 32'h8220000;
      16564: inst = 32'h10408000;
      16565: inst = 32'hc4053d1;
      16566: inst = 32'h8220000;
      16567: inst = 32'h10408000;
      16568: inst = 32'hc4053d2;
      16569: inst = 32'h8220000;
      16570: inst = 32'h10408000;
      16571: inst = 32'hc4053d3;
      16572: inst = 32'h8220000;
      16573: inst = 32'h10408000;
      16574: inst = 32'hc4053d4;
      16575: inst = 32'h8220000;
      16576: inst = 32'h10408000;
      16577: inst = 32'hc4053d5;
      16578: inst = 32'h8220000;
      16579: inst = 32'h10408000;
      16580: inst = 32'hc4053d6;
      16581: inst = 32'h8220000;
      16582: inst = 32'h10408000;
      16583: inst = 32'hc4053d7;
      16584: inst = 32'h8220000;
      16585: inst = 32'h10408000;
      16586: inst = 32'hc4053d8;
      16587: inst = 32'h8220000;
      16588: inst = 32'h10408000;
      16589: inst = 32'hc4053ea;
      16590: inst = 32'h8220000;
      16591: inst = 32'h10408000;
      16592: inst = 32'hc4053eb;
      16593: inst = 32'h8220000;
      16594: inst = 32'h10408000;
      16595: inst = 32'hc4053ec;
      16596: inst = 32'h8220000;
      16597: inst = 32'h10408000;
      16598: inst = 32'hc4053ed;
      16599: inst = 32'h8220000;
      16600: inst = 32'h10408000;
      16601: inst = 32'hc4053ee;
      16602: inst = 32'h8220000;
      16603: inst = 32'h10408000;
      16604: inst = 32'hc4053ef;
      16605: inst = 32'h8220000;
      16606: inst = 32'h10408000;
      16607: inst = 32'hc4053f0;
      16608: inst = 32'h8220000;
      16609: inst = 32'h10408000;
      16610: inst = 32'hc4053f1;
      16611: inst = 32'h8220000;
      16612: inst = 32'h10408000;
      16613: inst = 32'hc4053f2;
      16614: inst = 32'h8220000;
      16615: inst = 32'h10408000;
      16616: inst = 32'hc4053f3;
      16617: inst = 32'h8220000;
      16618: inst = 32'h10408000;
      16619: inst = 32'hc4053f4;
      16620: inst = 32'h8220000;
      16621: inst = 32'h10408000;
      16622: inst = 32'hc4053f5;
      16623: inst = 32'h8220000;
      16624: inst = 32'h10408000;
      16625: inst = 32'hc405407;
      16626: inst = 32'h8220000;
      16627: inst = 32'h10408000;
      16628: inst = 32'hc405408;
      16629: inst = 32'h8220000;
      16630: inst = 32'h10408000;
      16631: inst = 32'hc405409;
      16632: inst = 32'h8220000;
      16633: inst = 32'h10408000;
      16634: inst = 32'hc40540a;
      16635: inst = 32'h8220000;
      16636: inst = 32'h10408000;
      16637: inst = 32'hc40540b;
      16638: inst = 32'h8220000;
      16639: inst = 32'h10408000;
      16640: inst = 32'hc40540c;
      16641: inst = 32'h8220000;
      16642: inst = 32'h10408000;
      16643: inst = 32'hc40540d;
      16644: inst = 32'h8220000;
      16645: inst = 32'h10408000;
      16646: inst = 32'hc40540e;
      16647: inst = 32'h8220000;
      16648: inst = 32'h10408000;
      16649: inst = 32'hc40540f;
      16650: inst = 32'h8220000;
      16651: inst = 32'h10408000;
      16652: inst = 32'hc405410;
      16653: inst = 32'h8220000;
      16654: inst = 32'h10408000;
      16655: inst = 32'hc405411;
      16656: inst = 32'h8220000;
      16657: inst = 32'h10408000;
      16658: inst = 32'hc405412;
      16659: inst = 32'h8220000;
      16660: inst = 32'h10408000;
      16661: inst = 32'hc405413;
      16662: inst = 32'h8220000;
      16663: inst = 32'h10408000;
      16664: inst = 32'hc405414;
      16665: inst = 32'h8220000;
      16666: inst = 32'h10408000;
      16667: inst = 32'hc405415;
      16668: inst = 32'h8220000;
      16669: inst = 32'h10408000;
      16670: inst = 32'hc405416;
      16671: inst = 32'h8220000;
      16672: inst = 32'h10408000;
      16673: inst = 32'hc405417;
      16674: inst = 32'h8220000;
      16675: inst = 32'h10408000;
      16676: inst = 32'hc405418;
      16677: inst = 32'h8220000;
      16678: inst = 32'h10408000;
      16679: inst = 32'hc405419;
      16680: inst = 32'h8220000;
      16681: inst = 32'h10408000;
      16682: inst = 32'hc40541a;
      16683: inst = 32'h8220000;
      16684: inst = 32'h10408000;
      16685: inst = 32'hc40541b;
      16686: inst = 32'h8220000;
      16687: inst = 32'h10408000;
      16688: inst = 32'hc40541c;
      16689: inst = 32'h8220000;
      16690: inst = 32'h10408000;
      16691: inst = 32'hc40541d;
      16692: inst = 32'h8220000;
      16693: inst = 32'h10408000;
      16694: inst = 32'hc40541e;
      16695: inst = 32'h8220000;
      16696: inst = 32'h10408000;
      16697: inst = 32'hc40541f;
      16698: inst = 32'h8220000;
      16699: inst = 32'h10408000;
      16700: inst = 32'hc405420;
      16701: inst = 32'h8220000;
      16702: inst = 32'h10408000;
      16703: inst = 32'hc405421;
      16704: inst = 32'h8220000;
      16705: inst = 32'h10408000;
      16706: inst = 32'hc405422;
      16707: inst = 32'h8220000;
      16708: inst = 32'h10408000;
      16709: inst = 32'hc405423;
      16710: inst = 32'h8220000;
      16711: inst = 32'h10408000;
      16712: inst = 32'hc405424;
      16713: inst = 32'h8220000;
      16714: inst = 32'h10408000;
      16715: inst = 32'hc405425;
      16716: inst = 32'h8220000;
      16717: inst = 32'h10408000;
      16718: inst = 32'hc405426;
      16719: inst = 32'h8220000;
      16720: inst = 32'h10408000;
      16721: inst = 32'hc405427;
      16722: inst = 32'h8220000;
      16723: inst = 32'h10408000;
      16724: inst = 32'hc405428;
      16725: inst = 32'h8220000;
      16726: inst = 32'h10408000;
      16727: inst = 32'hc405429;
      16728: inst = 32'h8220000;
      16729: inst = 32'h10408000;
      16730: inst = 32'hc40542a;
      16731: inst = 32'h8220000;
      16732: inst = 32'h10408000;
      16733: inst = 32'hc40542b;
      16734: inst = 32'h8220000;
      16735: inst = 32'h10408000;
      16736: inst = 32'hc40542c;
      16737: inst = 32'h8220000;
      16738: inst = 32'h10408000;
      16739: inst = 32'hc40542d;
      16740: inst = 32'h8220000;
      16741: inst = 32'h10408000;
      16742: inst = 32'hc40542e;
      16743: inst = 32'h8220000;
      16744: inst = 32'h10408000;
      16745: inst = 32'hc40542f;
      16746: inst = 32'h8220000;
      16747: inst = 32'h10408000;
      16748: inst = 32'hc405430;
      16749: inst = 32'h8220000;
      16750: inst = 32'h10408000;
      16751: inst = 32'hc405431;
      16752: inst = 32'h8220000;
      16753: inst = 32'h10408000;
      16754: inst = 32'hc405432;
      16755: inst = 32'h8220000;
      16756: inst = 32'h10408000;
      16757: inst = 32'hc405433;
      16758: inst = 32'h8220000;
      16759: inst = 32'h10408000;
      16760: inst = 32'hc405434;
      16761: inst = 32'h8220000;
      16762: inst = 32'h10408000;
      16763: inst = 32'hc405435;
      16764: inst = 32'h8220000;
      16765: inst = 32'h10408000;
      16766: inst = 32'hc405436;
      16767: inst = 32'h8220000;
      16768: inst = 32'h10408000;
      16769: inst = 32'hc405437;
      16770: inst = 32'h8220000;
      16771: inst = 32'h10408000;
      16772: inst = 32'hc405438;
      16773: inst = 32'h8220000;
      16774: inst = 32'h10408000;
      16775: inst = 32'hc40544a;
      16776: inst = 32'h8220000;
      16777: inst = 32'h10408000;
      16778: inst = 32'hc40544b;
      16779: inst = 32'h8220000;
      16780: inst = 32'h10408000;
      16781: inst = 32'hc40544c;
      16782: inst = 32'h8220000;
      16783: inst = 32'h10408000;
      16784: inst = 32'hc40544d;
      16785: inst = 32'h8220000;
      16786: inst = 32'h10408000;
      16787: inst = 32'hc40544e;
      16788: inst = 32'h8220000;
      16789: inst = 32'h10408000;
      16790: inst = 32'hc40544f;
      16791: inst = 32'h8220000;
      16792: inst = 32'h10408000;
      16793: inst = 32'hc405450;
      16794: inst = 32'h8220000;
      16795: inst = 32'h10408000;
      16796: inst = 32'hc405451;
      16797: inst = 32'h8220000;
      16798: inst = 32'h10408000;
      16799: inst = 32'hc405452;
      16800: inst = 32'h8220000;
      16801: inst = 32'h10408000;
      16802: inst = 32'hc405453;
      16803: inst = 32'h8220000;
      16804: inst = 32'h10408000;
      16805: inst = 32'hc405454;
      16806: inst = 32'h8220000;
      16807: inst = 32'h10408000;
      16808: inst = 32'hc405455;
      16809: inst = 32'h8220000;
      16810: inst = 32'h10408000;
      16811: inst = 32'hc405467;
      16812: inst = 32'h8220000;
      16813: inst = 32'h10408000;
      16814: inst = 32'hc405468;
      16815: inst = 32'h8220000;
      16816: inst = 32'h10408000;
      16817: inst = 32'hc405469;
      16818: inst = 32'h8220000;
      16819: inst = 32'h10408000;
      16820: inst = 32'hc40546a;
      16821: inst = 32'h8220000;
      16822: inst = 32'h10408000;
      16823: inst = 32'hc40546b;
      16824: inst = 32'h8220000;
      16825: inst = 32'h10408000;
      16826: inst = 32'hc40546c;
      16827: inst = 32'h8220000;
      16828: inst = 32'h10408000;
      16829: inst = 32'hc40546d;
      16830: inst = 32'h8220000;
      16831: inst = 32'h10408000;
      16832: inst = 32'hc40546e;
      16833: inst = 32'h8220000;
      16834: inst = 32'h10408000;
      16835: inst = 32'hc40546f;
      16836: inst = 32'h8220000;
      16837: inst = 32'h10408000;
      16838: inst = 32'hc405470;
      16839: inst = 32'h8220000;
      16840: inst = 32'h10408000;
      16841: inst = 32'hc405471;
      16842: inst = 32'h8220000;
      16843: inst = 32'h10408000;
      16844: inst = 32'hc405472;
      16845: inst = 32'h8220000;
      16846: inst = 32'h10408000;
      16847: inst = 32'hc405473;
      16848: inst = 32'h8220000;
      16849: inst = 32'h10408000;
      16850: inst = 32'hc405474;
      16851: inst = 32'h8220000;
      16852: inst = 32'h10408000;
      16853: inst = 32'hc405475;
      16854: inst = 32'h8220000;
      16855: inst = 32'h10408000;
      16856: inst = 32'hc405476;
      16857: inst = 32'h8220000;
      16858: inst = 32'h10408000;
      16859: inst = 32'hc405477;
      16860: inst = 32'h8220000;
      16861: inst = 32'h10408000;
      16862: inst = 32'hc405478;
      16863: inst = 32'h8220000;
      16864: inst = 32'h10408000;
      16865: inst = 32'hc405479;
      16866: inst = 32'h8220000;
      16867: inst = 32'h10408000;
      16868: inst = 32'hc40547a;
      16869: inst = 32'h8220000;
      16870: inst = 32'h10408000;
      16871: inst = 32'hc40547b;
      16872: inst = 32'h8220000;
      16873: inst = 32'h10408000;
      16874: inst = 32'hc40547c;
      16875: inst = 32'h8220000;
      16876: inst = 32'h10408000;
      16877: inst = 32'hc40547d;
      16878: inst = 32'h8220000;
      16879: inst = 32'h10408000;
      16880: inst = 32'hc40547e;
      16881: inst = 32'h8220000;
      16882: inst = 32'h10408000;
      16883: inst = 32'hc40547f;
      16884: inst = 32'h8220000;
      16885: inst = 32'h10408000;
      16886: inst = 32'hc405480;
      16887: inst = 32'h8220000;
      16888: inst = 32'h10408000;
      16889: inst = 32'hc405481;
      16890: inst = 32'h8220000;
      16891: inst = 32'h10408000;
      16892: inst = 32'hc405482;
      16893: inst = 32'h8220000;
      16894: inst = 32'h10408000;
      16895: inst = 32'hc405483;
      16896: inst = 32'h8220000;
      16897: inst = 32'h10408000;
      16898: inst = 32'hc405484;
      16899: inst = 32'h8220000;
      16900: inst = 32'h10408000;
      16901: inst = 32'hc405485;
      16902: inst = 32'h8220000;
      16903: inst = 32'h10408000;
      16904: inst = 32'hc405486;
      16905: inst = 32'h8220000;
      16906: inst = 32'h10408000;
      16907: inst = 32'hc405487;
      16908: inst = 32'h8220000;
      16909: inst = 32'h10408000;
      16910: inst = 32'hc405488;
      16911: inst = 32'h8220000;
      16912: inst = 32'h10408000;
      16913: inst = 32'hc405489;
      16914: inst = 32'h8220000;
      16915: inst = 32'h10408000;
      16916: inst = 32'hc40548a;
      16917: inst = 32'h8220000;
      16918: inst = 32'h10408000;
      16919: inst = 32'hc40548b;
      16920: inst = 32'h8220000;
      16921: inst = 32'h10408000;
      16922: inst = 32'hc40548c;
      16923: inst = 32'h8220000;
      16924: inst = 32'h10408000;
      16925: inst = 32'hc40548d;
      16926: inst = 32'h8220000;
      16927: inst = 32'h10408000;
      16928: inst = 32'hc40548e;
      16929: inst = 32'h8220000;
      16930: inst = 32'h10408000;
      16931: inst = 32'hc40548f;
      16932: inst = 32'h8220000;
      16933: inst = 32'h10408000;
      16934: inst = 32'hc405490;
      16935: inst = 32'h8220000;
      16936: inst = 32'h10408000;
      16937: inst = 32'hc405491;
      16938: inst = 32'h8220000;
      16939: inst = 32'h10408000;
      16940: inst = 32'hc405492;
      16941: inst = 32'h8220000;
      16942: inst = 32'h10408000;
      16943: inst = 32'hc405493;
      16944: inst = 32'h8220000;
      16945: inst = 32'h10408000;
      16946: inst = 32'hc405494;
      16947: inst = 32'h8220000;
      16948: inst = 32'h10408000;
      16949: inst = 32'hc405495;
      16950: inst = 32'h8220000;
      16951: inst = 32'h10408000;
      16952: inst = 32'hc405496;
      16953: inst = 32'h8220000;
      16954: inst = 32'h10408000;
      16955: inst = 32'hc405497;
      16956: inst = 32'h8220000;
      16957: inst = 32'h10408000;
      16958: inst = 32'hc4054aa;
      16959: inst = 32'h8220000;
      16960: inst = 32'h10408000;
      16961: inst = 32'hc4054ab;
      16962: inst = 32'h8220000;
      16963: inst = 32'h10408000;
      16964: inst = 32'hc4054ac;
      16965: inst = 32'h8220000;
      16966: inst = 32'h10408000;
      16967: inst = 32'hc4054ad;
      16968: inst = 32'h8220000;
      16969: inst = 32'h10408000;
      16970: inst = 32'hc4054ae;
      16971: inst = 32'h8220000;
      16972: inst = 32'h10408000;
      16973: inst = 32'hc4054af;
      16974: inst = 32'h8220000;
      16975: inst = 32'h10408000;
      16976: inst = 32'hc4054b0;
      16977: inst = 32'h8220000;
      16978: inst = 32'h10408000;
      16979: inst = 32'hc4054b1;
      16980: inst = 32'h8220000;
      16981: inst = 32'h10408000;
      16982: inst = 32'hc4054b2;
      16983: inst = 32'h8220000;
      16984: inst = 32'h10408000;
      16985: inst = 32'hc4054b3;
      16986: inst = 32'h8220000;
      16987: inst = 32'h10408000;
      16988: inst = 32'hc4054b4;
      16989: inst = 32'h8220000;
      16990: inst = 32'h10408000;
      16991: inst = 32'hc4054b5;
      16992: inst = 32'h8220000;
      16993: inst = 32'h10408000;
      16994: inst = 32'hc4054c8;
      16995: inst = 32'h8220000;
      16996: inst = 32'h10408000;
      16997: inst = 32'hc4054c9;
      16998: inst = 32'h8220000;
      16999: inst = 32'h10408000;
      17000: inst = 32'hc4054ca;
      17001: inst = 32'h8220000;
      17002: inst = 32'h10408000;
      17003: inst = 32'hc4054cb;
      17004: inst = 32'h8220000;
      17005: inst = 32'h10408000;
      17006: inst = 32'hc4054cc;
      17007: inst = 32'h8220000;
      17008: inst = 32'h10408000;
      17009: inst = 32'hc4054cd;
      17010: inst = 32'h8220000;
      17011: inst = 32'h10408000;
      17012: inst = 32'hc4054ce;
      17013: inst = 32'h8220000;
      17014: inst = 32'h10408000;
      17015: inst = 32'hc4054cf;
      17016: inst = 32'h8220000;
      17017: inst = 32'h10408000;
      17018: inst = 32'hc4054d0;
      17019: inst = 32'h8220000;
      17020: inst = 32'h10408000;
      17021: inst = 32'hc4054d1;
      17022: inst = 32'h8220000;
      17023: inst = 32'h10408000;
      17024: inst = 32'hc4054d2;
      17025: inst = 32'h8220000;
      17026: inst = 32'h10408000;
      17027: inst = 32'hc4054d3;
      17028: inst = 32'h8220000;
      17029: inst = 32'h10408000;
      17030: inst = 32'hc4054d4;
      17031: inst = 32'h8220000;
      17032: inst = 32'h10408000;
      17033: inst = 32'hc4054d5;
      17034: inst = 32'h8220000;
      17035: inst = 32'h10408000;
      17036: inst = 32'hc4054d6;
      17037: inst = 32'h8220000;
      17038: inst = 32'h10408000;
      17039: inst = 32'hc4054d7;
      17040: inst = 32'h8220000;
      17041: inst = 32'h10408000;
      17042: inst = 32'hc4054d8;
      17043: inst = 32'h8220000;
      17044: inst = 32'h10408000;
      17045: inst = 32'hc4054d9;
      17046: inst = 32'h8220000;
      17047: inst = 32'h10408000;
      17048: inst = 32'hc4054da;
      17049: inst = 32'h8220000;
      17050: inst = 32'h10408000;
      17051: inst = 32'hc4054db;
      17052: inst = 32'h8220000;
      17053: inst = 32'h10408000;
      17054: inst = 32'hc4054dc;
      17055: inst = 32'h8220000;
      17056: inst = 32'h10408000;
      17057: inst = 32'hc4054dd;
      17058: inst = 32'h8220000;
      17059: inst = 32'h10408000;
      17060: inst = 32'hc4054de;
      17061: inst = 32'h8220000;
      17062: inst = 32'h10408000;
      17063: inst = 32'hc4054df;
      17064: inst = 32'h8220000;
      17065: inst = 32'h10408000;
      17066: inst = 32'hc4054e0;
      17067: inst = 32'h8220000;
      17068: inst = 32'h10408000;
      17069: inst = 32'hc4054e1;
      17070: inst = 32'h8220000;
      17071: inst = 32'h10408000;
      17072: inst = 32'hc4054e2;
      17073: inst = 32'h8220000;
      17074: inst = 32'h10408000;
      17075: inst = 32'hc4054e3;
      17076: inst = 32'h8220000;
      17077: inst = 32'h10408000;
      17078: inst = 32'hc4054e4;
      17079: inst = 32'h8220000;
      17080: inst = 32'h10408000;
      17081: inst = 32'hc4054e5;
      17082: inst = 32'h8220000;
      17083: inst = 32'h10408000;
      17084: inst = 32'hc4054e6;
      17085: inst = 32'h8220000;
      17086: inst = 32'h10408000;
      17087: inst = 32'hc4054e7;
      17088: inst = 32'h8220000;
      17089: inst = 32'h10408000;
      17090: inst = 32'hc4054e8;
      17091: inst = 32'h8220000;
      17092: inst = 32'h10408000;
      17093: inst = 32'hc4054e9;
      17094: inst = 32'h8220000;
      17095: inst = 32'h10408000;
      17096: inst = 32'hc4054ea;
      17097: inst = 32'h8220000;
      17098: inst = 32'h10408000;
      17099: inst = 32'hc4054eb;
      17100: inst = 32'h8220000;
      17101: inst = 32'h10408000;
      17102: inst = 32'hc4054ec;
      17103: inst = 32'h8220000;
      17104: inst = 32'h10408000;
      17105: inst = 32'hc4054ed;
      17106: inst = 32'h8220000;
      17107: inst = 32'h10408000;
      17108: inst = 32'hc4054ee;
      17109: inst = 32'h8220000;
      17110: inst = 32'h10408000;
      17111: inst = 32'hc4054ef;
      17112: inst = 32'h8220000;
      17113: inst = 32'h10408000;
      17114: inst = 32'hc4054f0;
      17115: inst = 32'h8220000;
      17116: inst = 32'h10408000;
      17117: inst = 32'hc4054f1;
      17118: inst = 32'h8220000;
      17119: inst = 32'h10408000;
      17120: inst = 32'hc4054f2;
      17121: inst = 32'h8220000;
      17122: inst = 32'h10408000;
      17123: inst = 32'hc4054f3;
      17124: inst = 32'h8220000;
      17125: inst = 32'h10408000;
      17126: inst = 32'hc4054f4;
      17127: inst = 32'h8220000;
      17128: inst = 32'h10408000;
      17129: inst = 32'hc4054f5;
      17130: inst = 32'h8220000;
      17131: inst = 32'h10408000;
      17132: inst = 32'hc4054f6;
      17133: inst = 32'h8220000;
      17134: inst = 32'h10408000;
      17135: inst = 32'hc40550a;
      17136: inst = 32'h8220000;
      17137: inst = 32'h10408000;
      17138: inst = 32'hc40550b;
      17139: inst = 32'h8220000;
      17140: inst = 32'h10408000;
      17141: inst = 32'hc40550c;
      17142: inst = 32'h8220000;
      17143: inst = 32'h10408000;
      17144: inst = 32'hc40550d;
      17145: inst = 32'h8220000;
      17146: inst = 32'h10408000;
      17147: inst = 32'hc40550e;
      17148: inst = 32'h8220000;
      17149: inst = 32'h10408000;
      17150: inst = 32'hc40550f;
      17151: inst = 32'h8220000;
      17152: inst = 32'h10408000;
      17153: inst = 32'hc405510;
      17154: inst = 32'h8220000;
      17155: inst = 32'h10408000;
      17156: inst = 32'hc405511;
      17157: inst = 32'h8220000;
      17158: inst = 32'h10408000;
      17159: inst = 32'hc405512;
      17160: inst = 32'h8220000;
      17161: inst = 32'h10408000;
      17162: inst = 32'hc405513;
      17163: inst = 32'h8220000;
      17164: inst = 32'h10408000;
      17165: inst = 32'hc405514;
      17166: inst = 32'h8220000;
      17167: inst = 32'h10408000;
      17168: inst = 32'hc405515;
      17169: inst = 32'h8220000;
      17170: inst = 32'h10408000;
      17171: inst = 32'hc405529;
      17172: inst = 32'h8220000;
      17173: inst = 32'h10408000;
      17174: inst = 32'hc40552a;
      17175: inst = 32'h8220000;
      17176: inst = 32'h10408000;
      17177: inst = 32'hc40552b;
      17178: inst = 32'h8220000;
      17179: inst = 32'h10408000;
      17180: inst = 32'hc40552c;
      17181: inst = 32'h8220000;
      17182: inst = 32'h10408000;
      17183: inst = 32'hc40552d;
      17184: inst = 32'h8220000;
      17185: inst = 32'h10408000;
      17186: inst = 32'hc40552e;
      17187: inst = 32'h8220000;
      17188: inst = 32'h10408000;
      17189: inst = 32'hc40552f;
      17190: inst = 32'h8220000;
      17191: inst = 32'h10408000;
      17192: inst = 32'hc405530;
      17193: inst = 32'h8220000;
      17194: inst = 32'h10408000;
      17195: inst = 32'hc405531;
      17196: inst = 32'h8220000;
      17197: inst = 32'h10408000;
      17198: inst = 32'hc405532;
      17199: inst = 32'h8220000;
      17200: inst = 32'h10408000;
      17201: inst = 32'hc405533;
      17202: inst = 32'h8220000;
      17203: inst = 32'h10408000;
      17204: inst = 32'hc405534;
      17205: inst = 32'h8220000;
      17206: inst = 32'h10408000;
      17207: inst = 32'hc405535;
      17208: inst = 32'h8220000;
      17209: inst = 32'h10408000;
      17210: inst = 32'hc405536;
      17211: inst = 32'h8220000;
      17212: inst = 32'h10408000;
      17213: inst = 32'hc405537;
      17214: inst = 32'h8220000;
      17215: inst = 32'h10408000;
      17216: inst = 32'hc405538;
      17217: inst = 32'h8220000;
      17218: inst = 32'h10408000;
      17219: inst = 32'hc405539;
      17220: inst = 32'h8220000;
      17221: inst = 32'h10408000;
      17222: inst = 32'hc40553a;
      17223: inst = 32'h8220000;
      17224: inst = 32'h10408000;
      17225: inst = 32'hc40553b;
      17226: inst = 32'h8220000;
      17227: inst = 32'h10408000;
      17228: inst = 32'hc40553c;
      17229: inst = 32'h8220000;
      17230: inst = 32'h10408000;
      17231: inst = 32'hc40553d;
      17232: inst = 32'h8220000;
      17233: inst = 32'h10408000;
      17234: inst = 32'hc40553e;
      17235: inst = 32'h8220000;
      17236: inst = 32'h10408000;
      17237: inst = 32'hc40553f;
      17238: inst = 32'h8220000;
      17239: inst = 32'h10408000;
      17240: inst = 32'hc405540;
      17241: inst = 32'h8220000;
      17242: inst = 32'h10408000;
      17243: inst = 32'hc405541;
      17244: inst = 32'h8220000;
      17245: inst = 32'h10408000;
      17246: inst = 32'hc405542;
      17247: inst = 32'h8220000;
      17248: inst = 32'h10408000;
      17249: inst = 32'hc405543;
      17250: inst = 32'h8220000;
      17251: inst = 32'h10408000;
      17252: inst = 32'hc405544;
      17253: inst = 32'h8220000;
      17254: inst = 32'h10408000;
      17255: inst = 32'hc405545;
      17256: inst = 32'h8220000;
      17257: inst = 32'h10408000;
      17258: inst = 32'hc405546;
      17259: inst = 32'h8220000;
      17260: inst = 32'h10408000;
      17261: inst = 32'hc405547;
      17262: inst = 32'h8220000;
      17263: inst = 32'h10408000;
      17264: inst = 32'hc405548;
      17265: inst = 32'h8220000;
      17266: inst = 32'h10408000;
      17267: inst = 32'hc405549;
      17268: inst = 32'h8220000;
      17269: inst = 32'h10408000;
      17270: inst = 32'hc40554a;
      17271: inst = 32'h8220000;
      17272: inst = 32'h10408000;
      17273: inst = 32'hc40554b;
      17274: inst = 32'h8220000;
      17275: inst = 32'h10408000;
      17276: inst = 32'hc40554c;
      17277: inst = 32'h8220000;
      17278: inst = 32'h10408000;
      17279: inst = 32'hc40554d;
      17280: inst = 32'h8220000;
      17281: inst = 32'h10408000;
      17282: inst = 32'hc40554e;
      17283: inst = 32'h8220000;
      17284: inst = 32'h10408000;
      17285: inst = 32'hc40554f;
      17286: inst = 32'h8220000;
      17287: inst = 32'h10408000;
      17288: inst = 32'hc405550;
      17289: inst = 32'h8220000;
      17290: inst = 32'h10408000;
      17291: inst = 32'hc405551;
      17292: inst = 32'h8220000;
      17293: inst = 32'h10408000;
      17294: inst = 32'hc405552;
      17295: inst = 32'h8220000;
      17296: inst = 32'h10408000;
      17297: inst = 32'hc405553;
      17298: inst = 32'h8220000;
      17299: inst = 32'h10408000;
      17300: inst = 32'hc405554;
      17301: inst = 32'h8220000;
      17302: inst = 32'h10408000;
      17303: inst = 32'hc405555;
      17304: inst = 32'h8220000;
      17305: inst = 32'h10408000;
      17306: inst = 32'hc40556a;
      17307: inst = 32'h8220000;
      17308: inst = 32'h10408000;
      17309: inst = 32'hc40556b;
      17310: inst = 32'h8220000;
      17311: inst = 32'h10408000;
      17312: inst = 32'hc40556c;
      17313: inst = 32'h8220000;
      17314: inst = 32'h10408000;
      17315: inst = 32'hc40556d;
      17316: inst = 32'h8220000;
      17317: inst = 32'h10408000;
      17318: inst = 32'hc40556e;
      17319: inst = 32'h8220000;
      17320: inst = 32'h10408000;
      17321: inst = 32'hc40556f;
      17322: inst = 32'h8220000;
      17323: inst = 32'h10408000;
      17324: inst = 32'hc405570;
      17325: inst = 32'h8220000;
      17326: inst = 32'h10408000;
      17327: inst = 32'hc405571;
      17328: inst = 32'h8220000;
      17329: inst = 32'h10408000;
      17330: inst = 32'hc405572;
      17331: inst = 32'h8220000;
      17332: inst = 32'h10408000;
      17333: inst = 32'hc405573;
      17334: inst = 32'h8220000;
      17335: inst = 32'h10408000;
      17336: inst = 32'hc405574;
      17337: inst = 32'h8220000;
      17338: inst = 32'h10408000;
      17339: inst = 32'hc405575;
      17340: inst = 32'h8220000;
      17341: inst = 32'h10408000;
      17342: inst = 32'hc40558a;
      17343: inst = 32'h8220000;
      17344: inst = 32'h10408000;
      17345: inst = 32'hc40558b;
      17346: inst = 32'h8220000;
      17347: inst = 32'h10408000;
      17348: inst = 32'hc40558c;
      17349: inst = 32'h8220000;
      17350: inst = 32'h10408000;
      17351: inst = 32'hc40558d;
      17352: inst = 32'h8220000;
      17353: inst = 32'h10408000;
      17354: inst = 32'hc40558e;
      17355: inst = 32'h8220000;
      17356: inst = 32'h10408000;
      17357: inst = 32'hc40558f;
      17358: inst = 32'h8220000;
      17359: inst = 32'h10408000;
      17360: inst = 32'hc405590;
      17361: inst = 32'h8220000;
      17362: inst = 32'h10408000;
      17363: inst = 32'hc405591;
      17364: inst = 32'h8220000;
      17365: inst = 32'h10408000;
      17366: inst = 32'hc405592;
      17367: inst = 32'h8220000;
      17368: inst = 32'h10408000;
      17369: inst = 32'hc405593;
      17370: inst = 32'h8220000;
      17371: inst = 32'h10408000;
      17372: inst = 32'hc405594;
      17373: inst = 32'h8220000;
      17374: inst = 32'h10408000;
      17375: inst = 32'hc405595;
      17376: inst = 32'h8220000;
      17377: inst = 32'h10408000;
      17378: inst = 32'hc405596;
      17379: inst = 32'h8220000;
      17380: inst = 32'h10408000;
      17381: inst = 32'hc405597;
      17382: inst = 32'h8220000;
      17383: inst = 32'h10408000;
      17384: inst = 32'hc405598;
      17385: inst = 32'h8220000;
      17386: inst = 32'h10408000;
      17387: inst = 32'hc405599;
      17388: inst = 32'h8220000;
      17389: inst = 32'h10408000;
      17390: inst = 32'hc40559a;
      17391: inst = 32'h8220000;
      17392: inst = 32'h10408000;
      17393: inst = 32'hc40559b;
      17394: inst = 32'h8220000;
      17395: inst = 32'h10408000;
      17396: inst = 32'hc40559c;
      17397: inst = 32'h8220000;
      17398: inst = 32'h10408000;
      17399: inst = 32'hc40559d;
      17400: inst = 32'h8220000;
      17401: inst = 32'h10408000;
      17402: inst = 32'hc40559e;
      17403: inst = 32'h8220000;
      17404: inst = 32'h10408000;
      17405: inst = 32'hc40559f;
      17406: inst = 32'h8220000;
      17407: inst = 32'h10408000;
      17408: inst = 32'hc4055a0;
      17409: inst = 32'h8220000;
      17410: inst = 32'h10408000;
      17411: inst = 32'hc4055a1;
      17412: inst = 32'h8220000;
      17413: inst = 32'h10408000;
      17414: inst = 32'hc4055a2;
      17415: inst = 32'h8220000;
      17416: inst = 32'h10408000;
      17417: inst = 32'hc4055a3;
      17418: inst = 32'h8220000;
      17419: inst = 32'h10408000;
      17420: inst = 32'hc4055a4;
      17421: inst = 32'h8220000;
      17422: inst = 32'h10408000;
      17423: inst = 32'hc4055a5;
      17424: inst = 32'h8220000;
      17425: inst = 32'h10408000;
      17426: inst = 32'hc4055a6;
      17427: inst = 32'h8220000;
      17428: inst = 32'h10408000;
      17429: inst = 32'hc4055a7;
      17430: inst = 32'h8220000;
      17431: inst = 32'h10408000;
      17432: inst = 32'hc4055a8;
      17433: inst = 32'h8220000;
      17434: inst = 32'h10408000;
      17435: inst = 32'hc4055a9;
      17436: inst = 32'h8220000;
      17437: inst = 32'h10408000;
      17438: inst = 32'hc4055aa;
      17439: inst = 32'h8220000;
      17440: inst = 32'h10408000;
      17441: inst = 32'hc4055ab;
      17442: inst = 32'h8220000;
      17443: inst = 32'h10408000;
      17444: inst = 32'hc4055ac;
      17445: inst = 32'h8220000;
      17446: inst = 32'h10408000;
      17447: inst = 32'hc4055ad;
      17448: inst = 32'h8220000;
      17449: inst = 32'h10408000;
      17450: inst = 32'hc4055ae;
      17451: inst = 32'h8220000;
      17452: inst = 32'h10408000;
      17453: inst = 32'hc4055af;
      17454: inst = 32'h8220000;
      17455: inst = 32'h10408000;
      17456: inst = 32'hc4055b0;
      17457: inst = 32'h8220000;
      17458: inst = 32'h10408000;
      17459: inst = 32'hc4055b1;
      17460: inst = 32'h8220000;
      17461: inst = 32'h10408000;
      17462: inst = 32'hc4055b2;
      17463: inst = 32'h8220000;
      17464: inst = 32'h10408000;
      17465: inst = 32'hc4055b3;
      17466: inst = 32'h8220000;
      17467: inst = 32'h10408000;
      17468: inst = 32'hc4055b4;
      17469: inst = 32'h8220000;
      17470: inst = 32'h10408000;
      17471: inst = 32'hc4055ca;
      17472: inst = 32'h8220000;
      17473: inst = 32'h10408000;
      17474: inst = 32'hc4055cb;
      17475: inst = 32'h8220000;
      17476: inst = 32'h10408000;
      17477: inst = 32'hc4055cc;
      17478: inst = 32'h8220000;
      17479: inst = 32'h10408000;
      17480: inst = 32'hc4055cd;
      17481: inst = 32'h8220000;
      17482: inst = 32'h10408000;
      17483: inst = 32'hc4055ce;
      17484: inst = 32'h8220000;
      17485: inst = 32'h10408000;
      17486: inst = 32'hc4055cf;
      17487: inst = 32'h8220000;
      17488: inst = 32'h10408000;
      17489: inst = 32'hc4055d0;
      17490: inst = 32'h8220000;
      17491: inst = 32'h10408000;
      17492: inst = 32'hc4055d1;
      17493: inst = 32'h8220000;
      17494: inst = 32'h10408000;
      17495: inst = 32'hc4055d2;
      17496: inst = 32'h8220000;
      17497: inst = 32'h10408000;
      17498: inst = 32'hc4055d3;
      17499: inst = 32'h8220000;
      17500: inst = 32'h10408000;
      17501: inst = 32'hc4055d4;
      17502: inst = 32'h8220000;
      17503: inst = 32'h10408000;
      17504: inst = 32'hc4055d5;
      17505: inst = 32'h8220000;
      17506: inst = 32'h10408000;
      17507: inst = 32'hc4055eb;
      17508: inst = 32'h8220000;
      17509: inst = 32'h10408000;
      17510: inst = 32'hc4055ec;
      17511: inst = 32'h8220000;
      17512: inst = 32'h10408000;
      17513: inst = 32'hc4055ed;
      17514: inst = 32'h8220000;
      17515: inst = 32'h10408000;
      17516: inst = 32'hc4055ee;
      17517: inst = 32'h8220000;
      17518: inst = 32'h10408000;
      17519: inst = 32'hc4055ef;
      17520: inst = 32'h8220000;
      17521: inst = 32'h10408000;
      17522: inst = 32'hc4055f0;
      17523: inst = 32'h8220000;
      17524: inst = 32'h10408000;
      17525: inst = 32'hc4055f1;
      17526: inst = 32'h8220000;
      17527: inst = 32'h10408000;
      17528: inst = 32'hc4055f2;
      17529: inst = 32'h8220000;
      17530: inst = 32'h10408000;
      17531: inst = 32'hc4055f3;
      17532: inst = 32'h8220000;
      17533: inst = 32'h10408000;
      17534: inst = 32'hc4055f4;
      17535: inst = 32'h8220000;
      17536: inst = 32'h10408000;
      17537: inst = 32'hc4055f5;
      17538: inst = 32'h8220000;
      17539: inst = 32'h10408000;
      17540: inst = 32'hc4055f6;
      17541: inst = 32'h8220000;
      17542: inst = 32'h10408000;
      17543: inst = 32'hc4055f7;
      17544: inst = 32'h8220000;
      17545: inst = 32'h10408000;
      17546: inst = 32'hc4055f8;
      17547: inst = 32'h8220000;
      17548: inst = 32'h10408000;
      17549: inst = 32'hc4055f9;
      17550: inst = 32'h8220000;
      17551: inst = 32'h10408000;
      17552: inst = 32'hc4055fa;
      17553: inst = 32'h8220000;
      17554: inst = 32'h10408000;
      17555: inst = 32'hc4055fb;
      17556: inst = 32'h8220000;
      17557: inst = 32'h10408000;
      17558: inst = 32'hc4055fc;
      17559: inst = 32'h8220000;
      17560: inst = 32'h10408000;
      17561: inst = 32'hc4055fd;
      17562: inst = 32'h8220000;
      17563: inst = 32'h10408000;
      17564: inst = 32'hc4055fe;
      17565: inst = 32'h8220000;
      17566: inst = 32'h10408000;
      17567: inst = 32'hc4055ff;
      17568: inst = 32'h8220000;
      17569: inst = 32'h10408000;
      17570: inst = 32'hc405600;
      17571: inst = 32'h8220000;
      17572: inst = 32'h10408000;
      17573: inst = 32'hc405601;
      17574: inst = 32'h8220000;
      17575: inst = 32'h10408000;
      17576: inst = 32'hc405602;
      17577: inst = 32'h8220000;
      17578: inst = 32'h10408000;
      17579: inst = 32'hc405603;
      17580: inst = 32'h8220000;
      17581: inst = 32'h10408000;
      17582: inst = 32'hc405604;
      17583: inst = 32'h8220000;
      17584: inst = 32'h10408000;
      17585: inst = 32'hc405605;
      17586: inst = 32'h8220000;
      17587: inst = 32'h10408000;
      17588: inst = 32'hc405606;
      17589: inst = 32'h8220000;
      17590: inst = 32'h10408000;
      17591: inst = 32'hc405607;
      17592: inst = 32'h8220000;
      17593: inst = 32'h10408000;
      17594: inst = 32'hc405608;
      17595: inst = 32'h8220000;
      17596: inst = 32'h10408000;
      17597: inst = 32'hc405609;
      17598: inst = 32'h8220000;
      17599: inst = 32'h10408000;
      17600: inst = 32'hc40560a;
      17601: inst = 32'h8220000;
      17602: inst = 32'h10408000;
      17603: inst = 32'hc40560b;
      17604: inst = 32'h8220000;
      17605: inst = 32'h10408000;
      17606: inst = 32'hc40560c;
      17607: inst = 32'h8220000;
      17608: inst = 32'h10408000;
      17609: inst = 32'hc40560d;
      17610: inst = 32'h8220000;
      17611: inst = 32'h10408000;
      17612: inst = 32'hc40560e;
      17613: inst = 32'h8220000;
      17614: inst = 32'h10408000;
      17615: inst = 32'hc40560f;
      17616: inst = 32'h8220000;
      17617: inst = 32'h10408000;
      17618: inst = 32'hc405610;
      17619: inst = 32'h8220000;
      17620: inst = 32'h10408000;
      17621: inst = 32'hc405611;
      17622: inst = 32'h8220000;
      17623: inst = 32'h10408000;
      17624: inst = 32'hc405612;
      17625: inst = 32'h8220000;
      17626: inst = 32'h10408000;
      17627: inst = 32'hc405613;
      17628: inst = 32'h8220000;
      17629: inst = 32'h10408000;
      17630: inst = 32'hc405614;
      17631: inst = 32'h8220000;
      17632: inst = 32'h10408000;
      17633: inst = 32'hc40562a;
      17634: inst = 32'h8220000;
      17635: inst = 32'h10408000;
      17636: inst = 32'hc40562b;
      17637: inst = 32'h8220000;
      17638: inst = 32'h10408000;
      17639: inst = 32'hc40562c;
      17640: inst = 32'h8220000;
      17641: inst = 32'h10408000;
      17642: inst = 32'hc40562d;
      17643: inst = 32'h8220000;
      17644: inst = 32'h10408000;
      17645: inst = 32'hc40562e;
      17646: inst = 32'h8220000;
      17647: inst = 32'h10408000;
      17648: inst = 32'hc40562f;
      17649: inst = 32'h8220000;
      17650: inst = 32'h10408000;
      17651: inst = 32'hc405630;
      17652: inst = 32'h8220000;
      17653: inst = 32'h10408000;
      17654: inst = 32'hc405631;
      17655: inst = 32'h8220000;
      17656: inst = 32'h10408000;
      17657: inst = 32'hc405632;
      17658: inst = 32'h8220000;
      17659: inst = 32'h10408000;
      17660: inst = 32'hc405633;
      17661: inst = 32'h8220000;
      17662: inst = 32'h10408000;
      17663: inst = 32'hc405634;
      17664: inst = 32'h8220000;
      17665: inst = 32'h10408000;
      17666: inst = 32'hc405635;
      17667: inst = 32'h8220000;
      17668: inst = 32'h10408000;
      17669: inst = 32'hc40564b;
      17670: inst = 32'h8220000;
      17671: inst = 32'h10408000;
      17672: inst = 32'hc40564c;
      17673: inst = 32'h8220000;
      17674: inst = 32'h10408000;
      17675: inst = 32'hc40564d;
      17676: inst = 32'h8220000;
      17677: inst = 32'h10408000;
      17678: inst = 32'hc40564e;
      17679: inst = 32'h8220000;
      17680: inst = 32'h10408000;
      17681: inst = 32'hc40564f;
      17682: inst = 32'h8220000;
      17683: inst = 32'h10408000;
      17684: inst = 32'hc405650;
      17685: inst = 32'h8220000;
      17686: inst = 32'h10408000;
      17687: inst = 32'hc405651;
      17688: inst = 32'h8220000;
      17689: inst = 32'h10408000;
      17690: inst = 32'hc405652;
      17691: inst = 32'h8220000;
      17692: inst = 32'h10408000;
      17693: inst = 32'hc405653;
      17694: inst = 32'h8220000;
      17695: inst = 32'h10408000;
      17696: inst = 32'hc405654;
      17697: inst = 32'h8220000;
      17698: inst = 32'h10408000;
      17699: inst = 32'hc405655;
      17700: inst = 32'h8220000;
      17701: inst = 32'h10408000;
      17702: inst = 32'hc405656;
      17703: inst = 32'h8220000;
      17704: inst = 32'h10408000;
      17705: inst = 32'hc405657;
      17706: inst = 32'h8220000;
      17707: inst = 32'h10408000;
      17708: inst = 32'hc405658;
      17709: inst = 32'h8220000;
      17710: inst = 32'h10408000;
      17711: inst = 32'hc405659;
      17712: inst = 32'h8220000;
      17713: inst = 32'h10408000;
      17714: inst = 32'hc40565a;
      17715: inst = 32'h8220000;
      17716: inst = 32'h10408000;
      17717: inst = 32'hc40565b;
      17718: inst = 32'h8220000;
      17719: inst = 32'h10408000;
      17720: inst = 32'hc40565c;
      17721: inst = 32'h8220000;
      17722: inst = 32'h10408000;
      17723: inst = 32'hc40565d;
      17724: inst = 32'h8220000;
      17725: inst = 32'h10408000;
      17726: inst = 32'hc40565e;
      17727: inst = 32'h8220000;
      17728: inst = 32'h10408000;
      17729: inst = 32'hc40565f;
      17730: inst = 32'h8220000;
      17731: inst = 32'h10408000;
      17732: inst = 32'hc405660;
      17733: inst = 32'h8220000;
      17734: inst = 32'h10408000;
      17735: inst = 32'hc405661;
      17736: inst = 32'h8220000;
      17737: inst = 32'h10408000;
      17738: inst = 32'hc405662;
      17739: inst = 32'h8220000;
      17740: inst = 32'h10408000;
      17741: inst = 32'hc405663;
      17742: inst = 32'h8220000;
      17743: inst = 32'h10408000;
      17744: inst = 32'hc405664;
      17745: inst = 32'h8220000;
      17746: inst = 32'h10408000;
      17747: inst = 32'hc405665;
      17748: inst = 32'h8220000;
      17749: inst = 32'h10408000;
      17750: inst = 32'hc405666;
      17751: inst = 32'h8220000;
      17752: inst = 32'h10408000;
      17753: inst = 32'hc405667;
      17754: inst = 32'h8220000;
      17755: inst = 32'h10408000;
      17756: inst = 32'hc405668;
      17757: inst = 32'h8220000;
      17758: inst = 32'h10408000;
      17759: inst = 32'hc405669;
      17760: inst = 32'h8220000;
      17761: inst = 32'h10408000;
      17762: inst = 32'hc40566a;
      17763: inst = 32'h8220000;
      17764: inst = 32'h10408000;
      17765: inst = 32'hc40566b;
      17766: inst = 32'h8220000;
      17767: inst = 32'h10408000;
      17768: inst = 32'hc40566c;
      17769: inst = 32'h8220000;
      17770: inst = 32'h10408000;
      17771: inst = 32'hc40566d;
      17772: inst = 32'h8220000;
      17773: inst = 32'h10408000;
      17774: inst = 32'hc40566e;
      17775: inst = 32'h8220000;
      17776: inst = 32'h10408000;
      17777: inst = 32'hc40566f;
      17778: inst = 32'h8220000;
      17779: inst = 32'h10408000;
      17780: inst = 32'hc405670;
      17781: inst = 32'h8220000;
      17782: inst = 32'h10408000;
      17783: inst = 32'hc405671;
      17784: inst = 32'h8220000;
      17785: inst = 32'h10408000;
      17786: inst = 32'hc405672;
      17787: inst = 32'h8220000;
      17788: inst = 32'h10408000;
      17789: inst = 32'hc405673;
      17790: inst = 32'h8220000;
      17791: inst = 32'h10408000;
      17792: inst = 32'hc40568a;
      17793: inst = 32'h8220000;
      17794: inst = 32'h10408000;
      17795: inst = 32'hc40568b;
      17796: inst = 32'h8220000;
      17797: inst = 32'h10408000;
      17798: inst = 32'hc40568c;
      17799: inst = 32'h8220000;
      17800: inst = 32'h10408000;
      17801: inst = 32'hc40568d;
      17802: inst = 32'h8220000;
      17803: inst = 32'h10408000;
      17804: inst = 32'hc40568e;
      17805: inst = 32'h8220000;
      17806: inst = 32'h10408000;
      17807: inst = 32'hc40568f;
      17808: inst = 32'h8220000;
      17809: inst = 32'h10408000;
      17810: inst = 32'hc405690;
      17811: inst = 32'h8220000;
      17812: inst = 32'h10408000;
      17813: inst = 32'hc405691;
      17814: inst = 32'h8220000;
      17815: inst = 32'h10408000;
      17816: inst = 32'hc405692;
      17817: inst = 32'h8220000;
      17818: inst = 32'h10408000;
      17819: inst = 32'hc405693;
      17820: inst = 32'h8220000;
      17821: inst = 32'h10408000;
      17822: inst = 32'hc405694;
      17823: inst = 32'h8220000;
      17824: inst = 32'h10408000;
      17825: inst = 32'hc405695;
      17826: inst = 32'h8220000;
      17827: inst = 32'h10408000;
      17828: inst = 32'hc4056ac;
      17829: inst = 32'h8220000;
      17830: inst = 32'h10408000;
      17831: inst = 32'hc4056ad;
      17832: inst = 32'h8220000;
      17833: inst = 32'h10408000;
      17834: inst = 32'hc4056ae;
      17835: inst = 32'h8220000;
      17836: inst = 32'h10408000;
      17837: inst = 32'hc4056af;
      17838: inst = 32'h8220000;
      17839: inst = 32'h10408000;
      17840: inst = 32'hc4056b0;
      17841: inst = 32'h8220000;
      17842: inst = 32'h10408000;
      17843: inst = 32'hc4056b1;
      17844: inst = 32'h8220000;
      17845: inst = 32'h10408000;
      17846: inst = 32'hc4056b2;
      17847: inst = 32'h8220000;
      17848: inst = 32'h10408000;
      17849: inst = 32'hc4056b3;
      17850: inst = 32'h8220000;
      17851: inst = 32'h10408000;
      17852: inst = 32'hc4056b4;
      17853: inst = 32'h8220000;
      17854: inst = 32'h10408000;
      17855: inst = 32'hc4056b5;
      17856: inst = 32'h8220000;
      17857: inst = 32'h10408000;
      17858: inst = 32'hc4056b6;
      17859: inst = 32'h8220000;
      17860: inst = 32'h10408000;
      17861: inst = 32'hc4056b7;
      17862: inst = 32'h8220000;
      17863: inst = 32'h10408000;
      17864: inst = 32'hc4056b8;
      17865: inst = 32'h8220000;
      17866: inst = 32'h10408000;
      17867: inst = 32'hc4056b9;
      17868: inst = 32'h8220000;
      17869: inst = 32'h10408000;
      17870: inst = 32'hc4056ba;
      17871: inst = 32'h8220000;
      17872: inst = 32'h10408000;
      17873: inst = 32'hc4056bb;
      17874: inst = 32'h8220000;
      17875: inst = 32'h10408000;
      17876: inst = 32'hc4056bc;
      17877: inst = 32'h8220000;
      17878: inst = 32'h10408000;
      17879: inst = 32'hc4056bd;
      17880: inst = 32'h8220000;
      17881: inst = 32'h10408000;
      17882: inst = 32'hc4056be;
      17883: inst = 32'h8220000;
      17884: inst = 32'h10408000;
      17885: inst = 32'hc4056bf;
      17886: inst = 32'h8220000;
      17887: inst = 32'h10408000;
      17888: inst = 32'hc4056c0;
      17889: inst = 32'h8220000;
      17890: inst = 32'h10408000;
      17891: inst = 32'hc4056c1;
      17892: inst = 32'h8220000;
      17893: inst = 32'h10408000;
      17894: inst = 32'hc4056c2;
      17895: inst = 32'h8220000;
      17896: inst = 32'h10408000;
      17897: inst = 32'hc4056c3;
      17898: inst = 32'h8220000;
      17899: inst = 32'h10408000;
      17900: inst = 32'hc4056c4;
      17901: inst = 32'h8220000;
      17902: inst = 32'h10408000;
      17903: inst = 32'hc4056c5;
      17904: inst = 32'h8220000;
      17905: inst = 32'h10408000;
      17906: inst = 32'hc4056c6;
      17907: inst = 32'h8220000;
      17908: inst = 32'h10408000;
      17909: inst = 32'hc4056c7;
      17910: inst = 32'h8220000;
      17911: inst = 32'h10408000;
      17912: inst = 32'hc4056c8;
      17913: inst = 32'h8220000;
      17914: inst = 32'h10408000;
      17915: inst = 32'hc4056c9;
      17916: inst = 32'h8220000;
      17917: inst = 32'h10408000;
      17918: inst = 32'hc4056ca;
      17919: inst = 32'h8220000;
      17920: inst = 32'h10408000;
      17921: inst = 32'hc4056cb;
      17922: inst = 32'h8220000;
      17923: inst = 32'h10408000;
      17924: inst = 32'hc4056cc;
      17925: inst = 32'h8220000;
      17926: inst = 32'h10408000;
      17927: inst = 32'hc4056cd;
      17928: inst = 32'h8220000;
      17929: inst = 32'h10408000;
      17930: inst = 32'hc4056ce;
      17931: inst = 32'h8220000;
      17932: inst = 32'h10408000;
      17933: inst = 32'hc4056cf;
      17934: inst = 32'h8220000;
      17935: inst = 32'h10408000;
      17936: inst = 32'hc4056d0;
      17937: inst = 32'h8220000;
      17938: inst = 32'h10408000;
      17939: inst = 32'hc4056d1;
      17940: inst = 32'h8220000;
      17941: inst = 32'h10408000;
      17942: inst = 32'hc4056d2;
      17943: inst = 32'h8220000;
      17944: inst = 32'h10408000;
      17945: inst = 32'hc4056ea;
      17946: inst = 32'h8220000;
      17947: inst = 32'h10408000;
      17948: inst = 32'hc4056eb;
      17949: inst = 32'h8220000;
      17950: inst = 32'h10408000;
      17951: inst = 32'hc4056ec;
      17952: inst = 32'h8220000;
      17953: inst = 32'h10408000;
      17954: inst = 32'hc4056ed;
      17955: inst = 32'h8220000;
      17956: inst = 32'h10408000;
      17957: inst = 32'hc4056ee;
      17958: inst = 32'h8220000;
      17959: inst = 32'h10408000;
      17960: inst = 32'hc4056ef;
      17961: inst = 32'h8220000;
      17962: inst = 32'h10408000;
      17963: inst = 32'hc4056f0;
      17964: inst = 32'h8220000;
      17965: inst = 32'h10408000;
      17966: inst = 32'hc4056f1;
      17967: inst = 32'h8220000;
      17968: inst = 32'h10408000;
      17969: inst = 32'hc4056f2;
      17970: inst = 32'h8220000;
      17971: inst = 32'h10408000;
      17972: inst = 32'hc4056f3;
      17973: inst = 32'h8220000;
      17974: inst = 32'h10408000;
      17975: inst = 32'hc4056f4;
      17976: inst = 32'h8220000;
      17977: inst = 32'h10408000;
      17978: inst = 32'hc4056f5;
      17979: inst = 32'h8220000;
      17980: inst = 32'h10408000;
      17981: inst = 32'hc40570d;
      17982: inst = 32'h8220000;
      17983: inst = 32'h10408000;
      17984: inst = 32'hc40570e;
      17985: inst = 32'h8220000;
      17986: inst = 32'h10408000;
      17987: inst = 32'hc40570f;
      17988: inst = 32'h8220000;
      17989: inst = 32'h10408000;
      17990: inst = 32'hc405710;
      17991: inst = 32'h8220000;
      17992: inst = 32'h10408000;
      17993: inst = 32'hc405711;
      17994: inst = 32'h8220000;
      17995: inst = 32'h10408000;
      17996: inst = 32'hc405712;
      17997: inst = 32'h8220000;
      17998: inst = 32'h10408000;
      17999: inst = 32'hc405713;
      18000: inst = 32'h8220000;
      18001: inst = 32'h10408000;
      18002: inst = 32'hc405714;
      18003: inst = 32'h8220000;
      18004: inst = 32'h10408000;
      18005: inst = 32'hc405715;
      18006: inst = 32'h8220000;
      18007: inst = 32'h10408000;
      18008: inst = 32'hc405716;
      18009: inst = 32'h8220000;
      18010: inst = 32'h10408000;
      18011: inst = 32'hc405717;
      18012: inst = 32'h8220000;
      18013: inst = 32'h10408000;
      18014: inst = 32'hc405718;
      18015: inst = 32'h8220000;
      18016: inst = 32'h10408000;
      18017: inst = 32'hc405719;
      18018: inst = 32'h8220000;
      18019: inst = 32'h10408000;
      18020: inst = 32'hc40571a;
      18021: inst = 32'h8220000;
      18022: inst = 32'h10408000;
      18023: inst = 32'hc40571b;
      18024: inst = 32'h8220000;
      18025: inst = 32'h10408000;
      18026: inst = 32'hc40571c;
      18027: inst = 32'h8220000;
      18028: inst = 32'h10408000;
      18029: inst = 32'hc40571d;
      18030: inst = 32'h8220000;
      18031: inst = 32'h10408000;
      18032: inst = 32'hc40571e;
      18033: inst = 32'h8220000;
      18034: inst = 32'h10408000;
      18035: inst = 32'hc40571f;
      18036: inst = 32'h8220000;
      18037: inst = 32'h10408000;
      18038: inst = 32'hc405720;
      18039: inst = 32'h8220000;
      18040: inst = 32'h10408000;
      18041: inst = 32'hc405721;
      18042: inst = 32'h8220000;
      18043: inst = 32'h10408000;
      18044: inst = 32'hc405722;
      18045: inst = 32'h8220000;
      18046: inst = 32'h10408000;
      18047: inst = 32'hc405723;
      18048: inst = 32'h8220000;
      18049: inst = 32'h10408000;
      18050: inst = 32'hc405724;
      18051: inst = 32'h8220000;
      18052: inst = 32'h10408000;
      18053: inst = 32'hc405725;
      18054: inst = 32'h8220000;
      18055: inst = 32'h10408000;
      18056: inst = 32'hc405726;
      18057: inst = 32'h8220000;
      18058: inst = 32'h10408000;
      18059: inst = 32'hc405727;
      18060: inst = 32'h8220000;
      18061: inst = 32'h10408000;
      18062: inst = 32'hc405728;
      18063: inst = 32'h8220000;
      18064: inst = 32'h10408000;
      18065: inst = 32'hc405729;
      18066: inst = 32'h8220000;
      18067: inst = 32'h10408000;
      18068: inst = 32'hc40572a;
      18069: inst = 32'h8220000;
      18070: inst = 32'h10408000;
      18071: inst = 32'hc40572b;
      18072: inst = 32'h8220000;
      18073: inst = 32'h10408000;
      18074: inst = 32'hc40572c;
      18075: inst = 32'h8220000;
      18076: inst = 32'h10408000;
      18077: inst = 32'hc40572d;
      18078: inst = 32'h8220000;
      18079: inst = 32'h10408000;
      18080: inst = 32'hc40572e;
      18081: inst = 32'h8220000;
      18082: inst = 32'h10408000;
      18083: inst = 32'hc40572f;
      18084: inst = 32'h8220000;
      18085: inst = 32'h10408000;
      18086: inst = 32'hc405730;
      18087: inst = 32'h8220000;
      18088: inst = 32'h10408000;
      18089: inst = 32'hc405731;
      18090: inst = 32'h8220000;
      18091: inst = 32'h10408000;
      18092: inst = 32'hc40574a;
      18093: inst = 32'h8220000;
      18094: inst = 32'h10408000;
      18095: inst = 32'hc40574b;
      18096: inst = 32'h8220000;
      18097: inst = 32'h10408000;
      18098: inst = 32'hc40574c;
      18099: inst = 32'h8220000;
      18100: inst = 32'h10408000;
      18101: inst = 32'hc40574d;
      18102: inst = 32'h8220000;
      18103: inst = 32'h10408000;
      18104: inst = 32'hc40574e;
      18105: inst = 32'h8220000;
      18106: inst = 32'h10408000;
      18107: inst = 32'hc40574f;
      18108: inst = 32'h8220000;
      18109: inst = 32'h10408000;
      18110: inst = 32'hc405750;
      18111: inst = 32'h8220000;
      18112: inst = 32'h10408000;
      18113: inst = 32'hc405751;
      18114: inst = 32'h8220000;
      18115: inst = 32'h10408000;
      18116: inst = 32'hc405752;
      18117: inst = 32'h8220000;
      18118: inst = 32'h10408000;
      18119: inst = 32'hc405753;
      18120: inst = 32'h8220000;
      18121: inst = 32'h10408000;
      18122: inst = 32'hc405754;
      18123: inst = 32'h8220000;
      18124: inst = 32'h10408000;
      18125: inst = 32'hc405755;
      18126: inst = 32'h8220000;
      18127: inst = 32'h10408000;
      18128: inst = 32'hc40576e;
      18129: inst = 32'h8220000;
      18130: inst = 32'h10408000;
      18131: inst = 32'hc40576f;
      18132: inst = 32'h8220000;
      18133: inst = 32'h10408000;
      18134: inst = 32'hc405770;
      18135: inst = 32'h8220000;
      18136: inst = 32'h10408000;
      18137: inst = 32'hc405771;
      18138: inst = 32'h8220000;
      18139: inst = 32'h10408000;
      18140: inst = 32'hc405772;
      18141: inst = 32'h8220000;
      18142: inst = 32'h10408000;
      18143: inst = 32'hc405773;
      18144: inst = 32'h8220000;
      18145: inst = 32'h10408000;
      18146: inst = 32'hc405774;
      18147: inst = 32'h8220000;
      18148: inst = 32'h10408000;
      18149: inst = 32'hc405775;
      18150: inst = 32'h8220000;
      18151: inst = 32'h10408000;
      18152: inst = 32'hc405776;
      18153: inst = 32'h8220000;
      18154: inst = 32'h10408000;
      18155: inst = 32'hc405777;
      18156: inst = 32'h8220000;
      18157: inst = 32'h10408000;
      18158: inst = 32'hc405778;
      18159: inst = 32'h8220000;
      18160: inst = 32'h10408000;
      18161: inst = 32'hc405779;
      18162: inst = 32'h8220000;
      18163: inst = 32'h10408000;
      18164: inst = 32'hc40577a;
      18165: inst = 32'h8220000;
      18166: inst = 32'h10408000;
      18167: inst = 32'hc40577b;
      18168: inst = 32'h8220000;
      18169: inst = 32'h10408000;
      18170: inst = 32'hc40577c;
      18171: inst = 32'h8220000;
      18172: inst = 32'h10408000;
      18173: inst = 32'hc40577d;
      18174: inst = 32'h8220000;
      18175: inst = 32'h10408000;
      18176: inst = 32'hc40577e;
      18177: inst = 32'h8220000;
      18178: inst = 32'h10408000;
      18179: inst = 32'hc40577f;
      18180: inst = 32'h8220000;
      18181: inst = 32'h10408000;
      18182: inst = 32'hc405780;
      18183: inst = 32'h8220000;
      18184: inst = 32'h10408000;
      18185: inst = 32'hc405781;
      18186: inst = 32'h8220000;
      18187: inst = 32'h10408000;
      18188: inst = 32'hc405782;
      18189: inst = 32'h8220000;
      18190: inst = 32'h10408000;
      18191: inst = 32'hc405783;
      18192: inst = 32'h8220000;
      18193: inst = 32'h10408000;
      18194: inst = 32'hc405784;
      18195: inst = 32'h8220000;
      18196: inst = 32'h10408000;
      18197: inst = 32'hc405785;
      18198: inst = 32'h8220000;
      18199: inst = 32'h10408000;
      18200: inst = 32'hc405786;
      18201: inst = 32'h8220000;
      18202: inst = 32'h10408000;
      18203: inst = 32'hc405787;
      18204: inst = 32'h8220000;
      18205: inst = 32'h10408000;
      18206: inst = 32'hc405788;
      18207: inst = 32'h8220000;
      18208: inst = 32'h10408000;
      18209: inst = 32'hc405789;
      18210: inst = 32'h8220000;
      18211: inst = 32'h10408000;
      18212: inst = 32'hc40578a;
      18213: inst = 32'h8220000;
      18214: inst = 32'h10408000;
      18215: inst = 32'hc40578b;
      18216: inst = 32'h8220000;
      18217: inst = 32'h10408000;
      18218: inst = 32'hc40578c;
      18219: inst = 32'h8220000;
      18220: inst = 32'h10408000;
      18221: inst = 32'hc40578d;
      18222: inst = 32'h8220000;
      18223: inst = 32'h10408000;
      18224: inst = 32'hc40578e;
      18225: inst = 32'h8220000;
      18226: inst = 32'h10408000;
      18227: inst = 32'hc40578f;
      18228: inst = 32'h8220000;
      18229: inst = 32'h10408000;
      18230: inst = 32'hc405790;
      18231: inst = 32'h8220000;
      18232: inst = 32'h10408000;
      18233: inst = 32'hc405791;
      18234: inst = 32'h8220000;
      18235: inst = 32'h10408000;
      18236: inst = 32'hc4057aa;
      18237: inst = 32'h8220000;
      18238: inst = 32'h10408000;
      18239: inst = 32'hc4057ab;
      18240: inst = 32'h8220000;
      18241: inst = 32'h10408000;
      18242: inst = 32'hc4057ac;
      18243: inst = 32'h8220000;
      18244: inst = 32'h10408000;
      18245: inst = 32'hc4057ad;
      18246: inst = 32'h8220000;
      18247: inst = 32'h10408000;
      18248: inst = 32'hc4057ae;
      18249: inst = 32'h8220000;
      18250: inst = 32'h10408000;
      18251: inst = 32'hc4057af;
      18252: inst = 32'h8220000;
      18253: inst = 32'h10408000;
      18254: inst = 32'hc4057b0;
      18255: inst = 32'h8220000;
      18256: inst = 32'h10408000;
      18257: inst = 32'hc4057b1;
      18258: inst = 32'h8220000;
      18259: inst = 32'h10408000;
      18260: inst = 32'hc4057b2;
      18261: inst = 32'h8220000;
      18262: inst = 32'h10408000;
      18263: inst = 32'hc4057b3;
      18264: inst = 32'h8220000;
      18265: inst = 32'h10408000;
      18266: inst = 32'hc4057b4;
      18267: inst = 32'h8220000;
      18268: inst = 32'h10408000;
      18269: inst = 32'hc4057b5;
      18270: inst = 32'h8220000;
      18271: inst = 32'h10408000;
      18272: inst = 32'hc4057ce;
      18273: inst = 32'h8220000;
      18274: inst = 32'h10408000;
      18275: inst = 32'hc4057cf;
      18276: inst = 32'h8220000;
      18277: inst = 32'h10408000;
      18278: inst = 32'hc4057d0;
      18279: inst = 32'h8220000;
      18280: inst = 32'h10408000;
      18281: inst = 32'hc4057d1;
      18282: inst = 32'h8220000;
      18283: inst = 32'h10408000;
      18284: inst = 32'hc4057d2;
      18285: inst = 32'h8220000;
      18286: inst = 32'h10408000;
      18287: inst = 32'hc4057d3;
      18288: inst = 32'h8220000;
      18289: inst = 32'h10408000;
      18290: inst = 32'hc4057d4;
      18291: inst = 32'h8220000;
      18292: inst = 32'h10408000;
      18293: inst = 32'hc4057d5;
      18294: inst = 32'h8220000;
      18295: inst = 32'h10408000;
      18296: inst = 32'hc4057d6;
      18297: inst = 32'h8220000;
      18298: inst = 32'h10408000;
      18299: inst = 32'hc4057d7;
      18300: inst = 32'h8220000;
      18301: inst = 32'h10408000;
      18302: inst = 32'hc4057d8;
      18303: inst = 32'h8220000;
      18304: inst = 32'h10408000;
      18305: inst = 32'hc4057d9;
      18306: inst = 32'h8220000;
      18307: inst = 32'h10408000;
      18308: inst = 32'hc4057da;
      18309: inst = 32'h8220000;
      18310: inst = 32'h10408000;
      18311: inst = 32'hc4057db;
      18312: inst = 32'h8220000;
      18313: inst = 32'h10408000;
      18314: inst = 32'hc4057dc;
      18315: inst = 32'h8220000;
      18316: inst = 32'h10408000;
      18317: inst = 32'hc4057dd;
      18318: inst = 32'h8220000;
      18319: inst = 32'h10408000;
      18320: inst = 32'hc4057de;
      18321: inst = 32'h8220000;
      18322: inst = 32'h10408000;
      18323: inst = 32'hc4057df;
      18324: inst = 32'h8220000;
      18325: inst = 32'hc207bd0;
      18326: inst = 32'h10408000;
      18327: inst = 32'hc40531b;
      18328: inst = 32'h8220000;
      18329: inst = 32'h10408000;
      18330: inst = 32'hc405344;
      18331: inst = 32'h8220000;
      18332: inst = 32'hc207bcf;
      18333: inst = 32'h10408000;
      18334: inst = 32'hc405321;
      18335: inst = 32'h8220000;
      18336: inst = 32'h10408000;
      18337: inst = 32'hc40533e;
      18338: inst = 32'h8220000;
      18339: inst = 32'h10408000;
      18340: inst = 32'hc405381;
      18341: inst = 32'h8220000;
      18342: inst = 32'h10408000;
      18343: inst = 32'hc40539e;
      18344: inst = 32'h8220000;
      18345: inst = 32'h10408000;
      18346: inst = 32'hc4053e1;
      18347: inst = 32'h8220000;
      18348: inst = 32'h10408000;
      18349: inst = 32'hc4053fe;
      18350: inst = 32'h8220000;
      18351: inst = 32'h10408000;
      18352: inst = 32'hc405441;
      18353: inst = 32'h8220000;
      18354: inst = 32'h10408000;
      18355: inst = 32'hc405448;
      18356: inst = 32'h8220000;
      18357: inst = 32'h10408000;
      18358: inst = 32'hc405457;
      18359: inst = 32'h8220000;
      18360: inst = 32'h10408000;
      18361: inst = 32'hc40545e;
      18362: inst = 32'h8220000;
      18363: inst = 32'h10408000;
      18364: inst = 32'hc405501;
      18365: inst = 32'h8220000;
      18366: inst = 32'h10408000;
      18367: inst = 32'hc40551e;
      18368: inst = 32'h8220000;
      18369: inst = 32'h10408000;
      18370: inst = 32'hc405561;
      18371: inst = 32'h8220000;
      18372: inst = 32'h10408000;
      18373: inst = 32'hc40557e;
      18374: inst = 32'h8220000;
      18375: inst = 32'h10408000;
      18376: inst = 32'hc4055b9;
      18377: inst = 32'h8220000;
      18378: inst = 32'h10408000;
      18379: inst = 32'hc4055c1;
      18380: inst = 32'h8220000;
      18381: inst = 32'h10408000;
      18382: inst = 32'hc4055de;
      18383: inst = 32'h8220000;
      18384: inst = 32'h10408000;
      18385: inst = 32'hc4055e6;
      18386: inst = 32'h8220000;
      18387: inst = 32'h10408000;
      18388: inst = 32'hc40561e;
      18389: inst = 32'h8220000;
      18390: inst = 32'h10408000;
      18391: inst = 32'hc405621;
      18392: inst = 32'h8220000;
      18393: inst = 32'h10408000;
      18394: inst = 32'hc40563e;
      18395: inst = 32'h8220000;
      18396: inst = 32'h10408000;
      18397: inst = 32'hc405641;
      18398: inst = 32'h8220000;
      18399: inst = 32'h10408000;
      18400: inst = 32'hc405681;
      18401: inst = 32'h8220000;
      18402: inst = 32'h10408000;
      18403: inst = 32'hc405698;
      18404: inst = 32'h8220000;
      18405: inst = 32'h10408000;
      18406: inst = 32'hc40569e;
      18407: inst = 32'h8220000;
      18408: inst = 32'h10408000;
      18409: inst = 32'hc4056e1;
      18410: inst = 32'h8220000;
      18411: inst = 32'h10408000;
      18412: inst = 32'hc4056fe;
      18413: inst = 32'h8220000;
      18414: inst = 32'hc207390;
      18415: inst = 32'h10408000;
      18416: inst = 32'hc40537a;
      18417: inst = 32'h8220000;
      18418: inst = 32'h10408000;
      18419: inst = 32'hc4053a5;
      18420: inst = 32'h8220000;
      18421: inst = 32'hc2052aa;
      18422: inst = 32'h10408000;
      18423: inst = 32'hc405389;
      18424: inst = 32'h8220000;
      18425: inst = 32'h10408000;
      18426: inst = 32'hc405396;
      18427: inst = 32'h8220000;
      18428: inst = 32'h10408000;
      18429: inst = 32'hc4054fb;
      18430: inst = 32'h8220000;
      18431: inst = 32'h10408000;
      18432: inst = 32'hc405503;
      18433: inst = 32'h8220000;
      18434: inst = 32'h10408000;
      18435: inst = 32'hc40551c;
      18436: inst = 32'h8220000;
      18437: inst = 32'h10408000;
      18438: inst = 32'hc405524;
      18439: inst = 32'h8220000;
      18440: inst = 32'h10408000;
      18441: inst = 32'hc4055c8;
      18442: inst = 32'h8220000;
      18443: inst = 32'h10408000;
      18444: inst = 32'hc4055d7;
      18445: inst = 32'h8220000;
      18446: inst = 32'h10408000;
      18447: inst = 32'hc405619;
      18448: inst = 32'h8220000;
      18449: inst = 32'h10408000;
      18450: inst = 32'hc405622;
      18451: inst = 32'h8220000;
      18452: inst = 32'h10408000;
      18453: inst = 32'hc40563d;
      18454: inst = 32'h8220000;
      18455: inst = 32'h10408000;
      18456: inst = 32'hc405646;
      18457: inst = 32'h8220000;
      18458: inst = 32'hc206b70;
      18459: inst = 32'h10408000;
      18460: inst = 32'hc4053d9;
      18461: inst = 32'h8220000;
      18462: inst = 32'h10408000;
      18463: inst = 32'hc405406;
      18464: inst = 32'h8220000;
      18465: inst = 32'h10408000;
      18466: inst = 32'hc405556;
      18467: inst = 32'h8220000;
      18468: inst = 32'h10408000;
      18469: inst = 32'hc405589;
      18470: inst = 32'h8220000;
      18471: inst = 32'h10408000;
      18472: inst = 32'hc4055b5;
      18473: inst = 32'h8220000;
      18474: inst = 32'h10408000;
      18475: inst = 32'hc4055ea;
      18476: inst = 32'h8220000;
      18477: inst = 32'h10408000;
      18478: inst = 32'hc405732;
      18479: inst = 32'h8220000;
      18480: inst = 32'h10408000;
      18481: inst = 32'hc40576d;
      18482: inst = 32'h8220000;
      18483: inst = 32'hc20736e;
      18484: inst = 32'h10408000;
      18485: inst = 32'hc4053e0;
      18486: inst = 32'h8220000;
      18487: inst = 32'h10408000;
      18488: inst = 32'hc4053ff;
      18489: inst = 32'h8220000;
      18490: inst = 32'hc205aaa;
      18491: inst = 32'h10408000;
      18492: inst = 32'hc4053e4;
      18493: inst = 32'h8220000;
      18494: inst = 32'h10408000;
      18495: inst = 32'hc4053fb;
      18496: inst = 32'h8220000;
      18497: inst = 32'hc208431;
      18498: inst = 32'h10408000;
      18499: inst = 32'hc4053e8;
      18500: inst = 32'h8220000;
      18501: inst = 32'h10408000;
      18502: inst = 32'hc4053f7;
      18503: inst = 32'h8220000;
      18504: inst = 32'h10408000;
      18505: inst = 32'hc405439;
      18506: inst = 32'h8220000;
      18507: inst = 32'h10408000;
      18508: inst = 32'hc405466;
      18509: inst = 32'h8220000;
      18510: inst = 32'h10408000;
      18511: inst = 32'hc4055b6;
      18512: inst = 32'h8220000;
      18513: inst = 32'h10408000;
      18514: inst = 32'hc4055e9;
      18515: inst = 32'h8220000;
      18516: inst = 32'h10408000;
      18517: inst = 32'hc405733;
      18518: inst = 32'h8220000;
      18519: inst = 32'h10408000;
      18520: inst = 32'hc40576c;
      18521: inst = 32'h8220000;
      18522: inst = 32'hc206b4d;
      18523: inst = 32'h10408000;
      18524: inst = 32'hc40543c;
      18525: inst = 32'h8220000;
      18526: inst = 32'h10408000;
      18527: inst = 32'hc405444;
      18528: inst = 32'h8220000;
      18529: inst = 32'h10408000;
      18530: inst = 32'hc40545b;
      18531: inst = 32'h8220000;
      18532: inst = 32'h10408000;
      18533: inst = 32'hc405463;
      18534: inst = 32'h8220000;
      18535: inst = 32'h10408000;
      18536: inst = 32'hc405563;
      18537: inst = 32'h8220000;
      18538: inst = 32'h10408000;
      18539: inst = 32'hc40557c;
      18540: inst = 32'h8220000;
      18541: inst = 32'h10408000;
      18542: inst = 32'hc405682;
      18543: inst = 32'h8220000;
      18544: inst = 32'h10408000;
      18545: inst = 32'hc40569d;
      18546: inst = 32'h8220000;
      18547: inst = 32'hc208430;
      18548: inst = 32'h10408000;
      18549: inst = 32'hc405440;
      18550: inst = 32'h8220000;
      18551: inst = 32'h10408000;
      18552: inst = 32'hc40545f;
      18553: inst = 32'h8220000;
      18554: inst = 32'hc207bf1;
      18555: inst = 32'h10408000;
      18556: inst = 32'hc405498;
      18557: inst = 32'h8220000;
      18558: inst = 32'h10408000;
      18559: inst = 32'hc4054c7;
      18560: inst = 32'h8220000;
      18561: inst = 32'h10408000;
      18562: inst = 32'hc405615;
      18563: inst = 32'h8220000;
      18564: inst = 32'h10408000;
      18565: inst = 32'hc40564a;
      18566: inst = 32'h8220000;
      18567: inst = 32'hc207bef;
      18568: inst = 32'h10408000;
      18569: inst = 32'hc40549b;
      18570: inst = 32'h8220000;
      18571: inst = 32'h10408000;
      18572: inst = 32'hc4054c4;
      18573: inst = 32'h8220000;
      18574: inst = 32'h10408000;
      18575: inst = 32'hc405687;
      18576: inst = 32'h8220000;
      18577: inst = 32'h10408000;
      18578: inst = 32'hc4056e2;
      18579: inst = 32'h8220000;
      18580: inst = 32'h10408000;
      18581: inst = 32'hc4056fd;
      18582: inst = 32'h8220000;
      18583: inst = 32'hc205aeb;
      18584: inst = 32'h10408000;
      18585: inst = 32'hc40549f;
      18586: inst = 32'h8220000;
      18587: inst = 32'h10408000;
      18588: inst = 32'hc4054c0;
      18589: inst = 32'h8220000;
      18590: inst = 32'hc206b6e;
      18591: inst = 32'h10408000;
      18592: inst = 32'hc4054a8;
      18593: inst = 32'h8220000;
      18594: inst = 32'h10408000;
      18595: inst = 32'hc4054b7;
      18596: inst = 32'h8220000;
      18597: inst = 32'h10408000;
      18598: inst = 32'hc4056e7;
      18599: inst = 32'h8220000;
      18600: inst = 32'h10408000;
      18601: inst = 32'hc4056f8;
      18602: inst = 32'h8220000;
      18603: inst = 32'hc2073b0;
      18604: inst = 32'h10408000;
      18605: inst = 32'hc4054f7;
      18606: inst = 32'h8220000;
      18607: inst = 32'h10408000;
      18608: inst = 32'hc405528;
      18609: inst = 32'h8220000;
      18610: inst = 32'h10408000;
      18611: inst = 32'hc405674;
      18612: inst = 32'h8220000;
      18613: inst = 32'h10408000;
      18614: inst = 32'hc4056ab;
      18615: inst = 32'h8220000;
      18616: inst = 32'hc2073ae;
      18617: inst = 32'h10408000;
      18618: inst = 32'hc4054ff;
      18619: inst = 32'h8220000;
      18620: inst = 32'h10408000;
      18621: inst = 32'hc405520;
      18622: inst = 32'h8220000;
      18623: inst = 32'hc20632d;
      18624: inst = 32'h10408000;
      18625: inst = 32'hc405508;
      18626: inst = 32'h8220000;
      18627: inst = 32'h10408000;
      18628: inst = 32'hc405517;
      18629: inst = 32'h8220000;
      18630: inst = 32'h10408000;
      18631: inst = 32'hc405747;
      18632: inst = 32'h8220000;
      18633: inst = 32'h10408000;
      18634: inst = 32'hc405758;
      18635: inst = 32'h8220000;
      18636: inst = 32'hc206b2d;
      18637: inst = 32'h10408000;
      18638: inst = 32'hc40555a;
      18639: inst = 32'h8220000;
      18640: inst = 32'h10408000;
      18641: inst = 32'hc405585;
      18642: inst = 32'h8220000;
      18643: inst = 32'hc20630c;
      18644: inst = 32'h10408000;
      18645: inst = 32'hc4055be;
      18646: inst = 32'h8220000;
      18647: inst = 32'h10408000;
      18648: inst = 32'hc4055e1;
      18649: inst = 32'h8220000;
      18650: inst = 32'h10408000;
      18651: inst = 32'hc405678;
      18652: inst = 32'h8220000;
      18653: inst = 32'hc20632c;
      18654: inst = 32'h10408000;
      18655: inst = 32'hc4056a7;
      18656: inst = 32'h8220000;
      18657: inst = 32'hc206b90;
      18658: inst = 32'h10408000;
      18659: inst = 32'hc4056d3;
      18660: inst = 32'h8220000;
      18661: inst = 32'h10408000;
      18662: inst = 32'hc40570c;
      18663: inst = 32'h8220000;
      18664: inst = 32'hc207c11;
      18665: inst = 32'h10408000;
      18666: inst = 32'hc405792;
      18667: inst = 32'h8220000;
      18668: inst = 32'h10408000;
      18669: inst = 32'hc4057cd;
      18670: inst = 32'h8220000;
      18671: inst = 32'h58000000;
      18672: inst = 32'hc20ea25;
      18673: inst = 32'h10408000;
      18674: inst = 32'hc40464d;
      18675: inst = 32'h8220000;
      18676: inst = 32'h10408000;
      18677: inst = 32'hc40464e;
      18678: inst = 32'h8220000;
      18679: inst = 32'h10408000;
      18680: inst = 32'hc40464f;
      18681: inst = 32'h8220000;
      18682: inst = 32'h10408000;
      18683: inst = 32'hc404650;
      18684: inst = 32'h8220000;
      18685: inst = 32'h10408000;
      18686: inst = 32'hc404651;
      18687: inst = 32'h8220000;
      18688: inst = 32'h10408000;
      18689: inst = 32'hc404652;
      18690: inst = 32'h8220000;
      18691: inst = 32'h10408000;
      18692: inst = 32'hc404653;
      18693: inst = 32'h8220000;
      18694: inst = 32'h10408000;
      18695: inst = 32'hc404654;
      18696: inst = 32'h8220000;
      18697: inst = 32'h10408000;
      18698: inst = 32'hc404655;
      18699: inst = 32'h8220000;
      18700: inst = 32'h10408000;
      18701: inst = 32'hc404659;
      18702: inst = 32'h8220000;
      18703: inst = 32'h10408000;
      18704: inst = 32'hc40465a;
      18705: inst = 32'h8220000;
      18706: inst = 32'h10408000;
      18707: inst = 32'hc40465b;
      18708: inst = 32'h8220000;
      18709: inst = 32'h10408000;
      18710: inst = 32'hc40465c;
      18711: inst = 32'h8220000;
      18712: inst = 32'h10408000;
      18713: inst = 32'hc40465d;
      18714: inst = 32'h8220000;
      18715: inst = 32'h10408000;
      18716: inst = 32'hc40465e;
      18717: inst = 32'h8220000;
      18718: inst = 32'h10408000;
      18719: inst = 32'hc40465f;
      18720: inst = 32'h8220000;
      18721: inst = 32'h10408000;
      18722: inst = 32'hc404660;
      18723: inst = 32'h8220000;
      18724: inst = 32'h10408000;
      18725: inst = 32'hc404661;
      18726: inst = 32'h8220000;
      18727: inst = 32'h10408000;
      18728: inst = 32'hc404663;
      18729: inst = 32'h8220000;
      18730: inst = 32'h10408000;
      18731: inst = 32'hc404664;
      18732: inst = 32'h8220000;
      18733: inst = 32'h10408000;
      18734: inst = 32'hc404665;
      18735: inst = 32'h8220000;
      18736: inst = 32'h10408000;
      18737: inst = 32'hc404666;
      18738: inst = 32'h8220000;
      18739: inst = 32'h10408000;
      18740: inst = 32'hc404667;
      18741: inst = 32'h8220000;
      18742: inst = 32'h10408000;
      18743: inst = 32'hc404668;
      18744: inst = 32'h8220000;
      18745: inst = 32'h10408000;
      18746: inst = 32'hc404669;
      18747: inst = 32'h8220000;
      18748: inst = 32'h10408000;
      18749: inst = 32'hc40466a;
      18750: inst = 32'h8220000;
      18751: inst = 32'h10408000;
      18752: inst = 32'hc40466b;
      18753: inst = 32'h8220000;
      18754: inst = 32'h10408000;
      18755: inst = 32'hc404671;
      18756: inst = 32'h8220000;
      18757: inst = 32'h10408000;
      18758: inst = 32'hc404672;
      18759: inst = 32'h8220000;
      18760: inst = 32'h10408000;
      18761: inst = 32'hc404673;
      18762: inst = 32'h8220000;
      18763: inst = 32'h10408000;
      18764: inst = 32'hc404674;
      18765: inst = 32'h8220000;
      18766: inst = 32'h10408000;
      18767: inst = 32'hc404675;
      18768: inst = 32'h8220000;
      18769: inst = 32'h10408000;
      18770: inst = 32'hc404676;
      18771: inst = 32'h8220000;
      18772: inst = 32'h10408000;
      18773: inst = 32'hc404677;
      18774: inst = 32'h8220000;
      18775: inst = 32'h10408000;
      18776: inst = 32'hc404678;
      18777: inst = 32'h8220000;
      18778: inst = 32'h10408000;
      18779: inst = 32'hc404679;
      18780: inst = 32'h8220000;
      18781: inst = 32'h10408000;
      18782: inst = 32'hc40467c;
      18783: inst = 32'h8220000;
      18784: inst = 32'h10408000;
      18785: inst = 32'hc40467d;
      18786: inst = 32'h8220000;
      18787: inst = 32'h10408000;
      18788: inst = 32'hc40467e;
      18789: inst = 32'h8220000;
      18790: inst = 32'h10408000;
      18791: inst = 32'hc40467f;
      18792: inst = 32'h8220000;
      18793: inst = 32'h10408000;
      18794: inst = 32'hc404680;
      18795: inst = 32'h8220000;
      18796: inst = 32'h10408000;
      18797: inst = 32'hc404681;
      18798: inst = 32'h8220000;
      18799: inst = 32'h10408000;
      18800: inst = 32'hc404682;
      18801: inst = 32'h8220000;
      18802: inst = 32'h10408000;
      18803: inst = 32'hc404683;
      18804: inst = 32'h8220000;
      18805: inst = 32'h10408000;
      18806: inst = 32'hc404684;
      18807: inst = 32'h8220000;
      18808: inst = 32'h10408000;
      18809: inst = 32'hc404685;
      18810: inst = 32'h8220000;
      18811: inst = 32'h10408000;
      18812: inst = 32'hc40468b;
      18813: inst = 32'h8220000;
      18814: inst = 32'h10408000;
      18815: inst = 32'hc40468c;
      18816: inst = 32'h8220000;
      18817: inst = 32'h10408000;
      18818: inst = 32'hc40468d;
      18819: inst = 32'h8220000;
      18820: inst = 32'h10408000;
      18821: inst = 32'hc40468e;
      18822: inst = 32'h8220000;
      18823: inst = 32'h10408000;
      18824: inst = 32'hc40468f;
      18825: inst = 32'h8220000;
      18826: inst = 32'h10408000;
      18827: inst = 32'hc404690;
      18828: inst = 32'h8220000;
      18829: inst = 32'h10408000;
      18830: inst = 32'hc404691;
      18831: inst = 32'h8220000;
      18832: inst = 32'h10408000;
      18833: inst = 32'hc404692;
      18834: inst = 32'h8220000;
      18835: inst = 32'h10408000;
      18836: inst = 32'hc404693;
      18837: inst = 32'h8220000;
      18838: inst = 32'h10408000;
      18839: inst = 32'hc4046ac;
      18840: inst = 32'h8220000;
      18841: inst = 32'h10408000;
      18842: inst = 32'hc4046ad;
      18843: inst = 32'h8220000;
      18844: inst = 32'h10408000;
      18845: inst = 32'hc4046ae;
      18846: inst = 32'h8220000;
      18847: inst = 32'h10408000;
      18848: inst = 32'hc4046af;
      18849: inst = 32'h8220000;
      18850: inst = 32'h10408000;
      18851: inst = 32'hc4046b0;
      18852: inst = 32'h8220000;
      18853: inst = 32'h10408000;
      18854: inst = 32'hc4046b1;
      18855: inst = 32'h8220000;
      18856: inst = 32'h10408000;
      18857: inst = 32'hc4046b2;
      18858: inst = 32'h8220000;
      18859: inst = 32'h10408000;
      18860: inst = 32'hc4046b3;
      18861: inst = 32'h8220000;
      18862: inst = 32'h10408000;
      18863: inst = 32'hc4046b4;
      18864: inst = 32'h8220000;
      18865: inst = 32'h10408000;
      18866: inst = 32'hc4046b5;
      18867: inst = 32'h8220000;
      18868: inst = 32'h10408000;
      18869: inst = 32'hc4046b8;
      18870: inst = 32'h8220000;
      18871: inst = 32'h10408000;
      18872: inst = 32'hc4046b9;
      18873: inst = 32'h8220000;
      18874: inst = 32'h10408000;
      18875: inst = 32'hc4046ba;
      18876: inst = 32'h8220000;
      18877: inst = 32'h10408000;
      18878: inst = 32'hc4046bb;
      18879: inst = 32'h8220000;
      18880: inst = 32'h10408000;
      18881: inst = 32'hc4046bc;
      18882: inst = 32'h8220000;
      18883: inst = 32'h10408000;
      18884: inst = 32'hc4046bd;
      18885: inst = 32'h8220000;
      18886: inst = 32'h10408000;
      18887: inst = 32'hc4046be;
      18888: inst = 32'h8220000;
      18889: inst = 32'h10408000;
      18890: inst = 32'hc4046bf;
      18891: inst = 32'h8220000;
      18892: inst = 32'h10408000;
      18893: inst = 32'hc4046c0;
      18894: inst = 32'h8220000;
      18895: inst = 32'h10408000;
      18896: inst = 32'hc4046c1;
      18897: inst = 32'h8220000;
      18898: inst = 32'h10408000;
      18899: inst = 32'hc4046c3;
      18900: inst = 32'h8220000;
      18901: inst = 32'h10408000;
      18902: inst = 32'hc4046c4;
      18903: inst = 32'h8220000;
      18904: inst = 32'h10408000;
      18905: inst = 32'hc4046c5;
      18906: inst = 32'h8220000;
      18907: inst = 32'h10408000;
      18908: inst = 32'hc4046c6;
      18909: inst = 32'h8220000;
      18910: inst = 32'h10408000;
      18911: inst = 32'hc4046c7;
      18912: inst = 32'h8220000;
      18913: inst = 32'h10408000;
      18914: inst = 32'hc4046c8;
      18915: inst = 32'h8220000;
      18916: inst = 32'h10408000;
      18917: inst = 32'hc4046c9;
      18918: inst = 32'h8220000;
      18919: inst = 32'h10408000;
      18920: inst = 32'hc4046ca;
      18921: inst = 32'h8220000;
      18922: inst = 32'h10408000;
      18923: inst = 32'hc4046cb;
      18924: inst = 32'h8220000;
      18925: inst = 32'h10408000;
      18926: inst = 32'hc4046d0;
      18927: inst = 32'h8220000;
      18928: inst = 32'h10408000;
      18929: inst = 32'hc4046d1;
      18930: inst = 32'h8220000;
      18931: inst = 32'h10408000;
      18932: inst = 32'hc4046d2;
      18933: inst = 32'h8220000;
      18934: inst = 32'h10408000;
      18935: inst = 32'hc4046d3;
      18936: inst = 32'h8220000;
      18937: inst = 32'h10408000;
      18938: inst = 32'hc4046d4;
      18939: inst = 32'h8220000;
      18940: inst = 32'h10408000;
      18941: inst = 32'hc4046d5;
      18942: inst = 32'h8220000;
      18943: inst = 32'h10408000;
      18944: inst = 32'hc4046d6;
      18945: inst = 32'h8220000;
      18946: inst = 32'h10408000;
      18947: inst = 32'hc4046d7;
      18948: inst = 32'h8220000;
      18949: inst = 32'h10408000;
      18950: inst = 32'hc4046d8;
      18951: inst = 32'h8220000;
      18952: inst = 32'h10408000;
      18953: inst = 32'hc4046da;
      18954: inst = 32'h8220000;
      18955: inst = 32'h10408000;
      18956: inst = 32'hc4046dc;
      18957: inst = 32'h8220000;
      18958: inst = 32'h10408000;
      18959: inst = 32'hc4046dd;
      18960: inst = 32'h8220000;
      18961: inst = 32'h10408000;
      18962: inst = 32'hc4046de;
      18963: inst = 32'h8220000;
      18964: inst = 32'h10408000;
      18965: inst = 32'hc4046df;
      18966: inst = 32'h8220000;
      18967: inst = 32'h10408000;
      18968: inst = 32'hc4046e0;
      18969: inst = 32'h8220000;
      18970: inst = 32'h10408000;
      18971: inst = 32'hc4046e1;
      18972: inst = 32'h8220000;
      18973: inst = 32'h10408000;
      18974: inst = 32'hc4046e2;
      18975: inst = 32'h8220000;
      18976: inst = 32'h10408000;
      18977: inst = 32'hc4046e3;
      18978: inst = 32'h8220000;
      18979: inst = 32'h10408000;
      18980: inst = 32'hc4046e4;
      18981: inst = 32'h8220000;
      18982: inst = 32'h10408000;
      18983: inst = 32'hc4046e5;
      18984: inst = 32'h8220000;
      18985: inst = 32'h10408000;
      18986: inst = 32'hc4046ea;
      18987: inst = 32'h8220000;
      18988: inst = 32'h10408000;
      18989: inst = 32'hc4046eb;
      18990: inst = 32'h8220000;
      18991: inst = 32'h10408000;
      18992: inst = 32'hc4046ec;
      18993: inst = 32'h8220000;
      18994: inst = 32'h10408000;
      18995: inst = 32'hc4046ed;
      18996: inst = 32'h8220000;
      18997: inst = 32'h10408000;
      18998: inst = 32'hc4046ee;
      18999: inst = 32'h8220000;
      19000: inst = 32'h10408000;
      19001: inst = 32'hc4046ef;
      19002: inst = 32'h8220000;
      19003: inst = 32'h10408000;
      19004: inst = 32'hc4046f0;
      19005: inst = 32'h8220000;
      19006: inst = 32'h10408000;
      19007: inst = 32'hc4046f1;
      19008: inst = 32'h8220000;
      19009: inst = 32'h10408000;
      19010: inst = 32'hc4046f2;
      19011: inst = 32'h8220000;
      19012: inst = 32'h10408000;
      19013: inst = 32'hc4046f3;
      19014: inst = 32'h8220000;
      19015: inst = 32'h10408000;
      19016: inst = 32'hc40470b;
      19017: inst = 32'h8220000;
      19018: inst = 32'h10408000;
      19019: inst = 32'hc40470c;
      19020: inst = 32'h8220000;
      19021: inst = 32'h10408000;
      19022: inst = 32'hc40470d;
      19023: inst = 32'h8220000;
      19024: inst = 32'h10408000;
      19025: inst = 32'hc404717;
      19026: inst = 32'h8220000;
      19027: inst = 32'h10408000;
      19028: inst = 32'hc404718;
      19029: inst = 32'h8220000;
      19030: inst = 32'h10408000;
      19031: inst = 32'hc404719;
      19032: inst = 32'h8220000;
      19033: inst = 32'h10408000;
      19034: inst = 32'hc404728;
      19035: inst = 32'h8220000;
      19036: inst = 32'h10408000;
      19037: inst = 32'hc404729;
      19038: inst = 32'h8220000;
      19039: inst = 32'h10408000;
      19040: inst = 32'hc40472a;
      19041: inst = 32'h8220000;
      19042: inst = 32'h10408000;
      19043: inst = 32'hc40472b;
      19044: inst = 32'h8220000;
      19045: inst = 32'h10408000;
      19046: inst = 32'hc404730;
      19047: inst = 32'h8220000;
      19048: inst = 32'h10408000;
      19049: inst = 32'hc404731;
      19050: inst = 32'h8220000;
      19051: inst = 32'h10408000;
      19052: inst = 32'hc404735;
      19053: inst = 32'h8220000;
      19054: inst = 32'h10408000;
      19055: inst = 32'hc404736;
      19056: inst = 32'h8220000;
      19057: inst = 32'h10408000;
      19058: inst = 32'hc404737;
      19059: inst = 32'h8220000;
      19060: inst = 32'h10408000;
      19061: inst = 32'hc404739;
      19062: inst = 32'h8220000;
      19063: inst = 32'h10408000;
      19064: inst = 32'hc40473a;
      19065: inst = 32'h8220000;
      19066: inst = 32'h10408000;
      19067: inst = 32'hc404742;
      19068: inst = 32'h8220000;
      19069: inst = 32'h10408000;
      19070: inst = 32'hc404743;
      19071: inst = 32'h8220000;
      19072: inst = 32'h10408000;
      19073: inst = 32'hc404744;
      19074: inst = 32'h8220000;
      19075: inst = 32'h10408000;
      19076: inst = 32'hc404745;
      19077: inst = 32'h8220000;
      19078: inst = 32'h10408000;
      19079: inst = 32'hc404749;
      19080: inst = 32'h8220000;
      19081: inst = 32'h10408000;
      19082: inst = 32'hc40474a;
      19083: inst = 32'h8220000;
      19084: inst = 32'h10408000;
      19085: inst = 32'hc40474b;
      19086: inst = 32'h8220000;
      19087: inst = 32'h10408000;
      19088: inst = 32'hc40476b;
      19089: inst = 32'h8220000;
      19090: inst = 32'h10408000;
      19091: inst = 32'hc40476c;
      19092: inst = 32'h8220000;
      19093: inst = 32'h10408000;
      19094: inst = 32'hc404777;
      19095: inst = 32'h8220000;
      19096: inst = 32'h10408000;
      19097: inst = 32'hc404778;
      19098: inst = 32'h8220000;
      19099: inst = 32'h10408000;
      19100: inst = 32'hc404788;
      19101: inst = 32'h8220000;
      19102: inst = 32'h10408000;
      19103: inst = 32'hc404789;
      19104: inst = 32'h8220000;
      19105: inst = 32'h10408000;
      19106: inst = 32'hc40478a;
      19107: inst = 32'h8220000;
      19108: inst = 32'h10408000;
      19109: inst = 32'hc404790;
      19110: inst = 32'h8220000;
      19111: inst = 32'h10408000;
      19112: inst = 32'hc404791;
      19113: inst = 32'h8220000;
      19114: inst = 32'h10408000;
      19115: inst = 32'hc404795;
      19116: inst = 32'h8220000;
      19117: inst = 32'h10408000;
      19118: inst = 32'hc404799;
      19119: inst = 32'h8220000;
      19120: inst = 32'h10408000;
      19121: inst = 32'hc40479a;
      19122: inst = 32'h8220000;
      19123: inst = 32'h10408000;
      19124: inst = 32'hc4047a2;
      19125: inst = 32'h8220000;
      19126: inst = 32'h10408000;
      19127: inst = 32'hc4047a3;
      19128: inst = 32'h8220000;
      19129: inst = 32'h10408000;
      19130: inst = 32'hc4047a4;
      19131: inst = 32'h8220000;
      19132: inst = 32'h10408000;
      19133: inst = 32'hc4047a9;
      19134: inst = 32'h8220000;
      19135: inst = 32'h10408000;
      19136: inst = 32'hc4047aa;
      19137: inst = 32'h8220000;
      19138: inst = 32'h10408000;
      19139: inst = 32'hc4047cb;
      19140: inst = 32'h8220000;
      19141: inst = 32'h10408000;
      19142: inst = 32'hc4047cc;
      19143: inst = 32'h8220000;
      19144: inst = 32'h10408000;
      19145: inst = 32'hc4047ce;
      19146: inst = 32'h8220000;
      19147: inst = 32'h10408000;
      19148: inst = 32'hc4047cf;
      19149: inst = 32'h8220000;
      19150: inst = 32'h10408000;
      19151: inst = 32'hc4047d0;
      19152: inst = 32'h8220000;
      19153: inst = 32'h10408000;
      19154: inst = 32'hc4047d1;
      19155: inst = 32'h8220000;
      19156: inst = 32'h10408000;
      19157: inst = 32'hc4047d2;
      19158: inst = 32'h8220000;
      19159: inst = 32'h10408000;
      19160: inst = 32'hc4047d7;
      19161: inst = 32'h8220000;
      19162: inst = 32'h10408000;
      19163: inst = 32'hc4047d8;
      19164: inst = 32'h8220000;
      19165: inst = 32'h10408000;
      19166: inst = 32'hc4047da;
      19167: inst = 32'h8220000;
      19168: inst = 32'h10408000;
      19169: inst = 32'hc4047db;
      19170: inst = 32'h8220000;
      19171: inst = 32'h10408000;
      19172: inst = 32'hc4047dc;
      19173: inst = 32'h8220000;
      19174: inst = 32'h10408000;
      19175: inst = 32'hc4047dd;
      19176: inst = 32'h8220000;
      19177: inst = 32'h10408000;
      19178: inst = 32'hc4047de;
      19179: inst = 32'h8220000;
      19180: inst = 32'h10408000;
      19181: inst = 32'hc4047e7;
      19182: inst = 32'h8220000;
      19183: inst = 32'h10408000;
      19184: inst = 32'hc4047e8;
      19185: inst = 32'h8220000;
      19186: inst = 32'h10408000;
      19187: inst = 32'hc4047e9;
      19188: inst = 32'h8220000;
      19189: inst = 32'h10408000;
      19190: inst = 32'hc4047f0;
      19191: inst = 32'h8220000;
      19192: inst = 32'h10408000;
      19193: inst = 32'hc4047f1;
      19194: inst = 32'h8220000;
      19195: inst = 32'h10408000;
      19196: inst = 32'hc4047f9;
      19197: inst = 32'h8220000;
      19198: inst = 32'h10408000;
      19199: inst = 32'hc4047fa;
      19200: inst = 32'h8220000;
      19201: inst = 32'h10408000;
      19202: inst = 32'hc404800;
      19203: inst = 32'h8220000;
      19204: inst = 32'h10408000;
      19205: inst = 32'hc404801;
      19206: inst = 32'h8220000;
      19207: inst = 32'h10408000;
      19208: inst = 32'hc404802;
      19209: inst = 32'h8220000;
      19210: inst = 32'h10408000;
      19211: inst = 32'hc404803;
      19212: inst = 32'h8220000;
      19213: inst = 32'h10408000;
      19214: inst = 32'hc404809;
      19215: inst = 32'h8220000;
      19216: inst = 32'h10408000;
      19217: inst = 32'hc40480a;
      19218: inst = 32'h8220000;
      19219: inst = 32'h10408000;
      19220: inst = 32'hc40480c;
      19221: inst = 32'h8220000;
      19222: inst = 32'h10408000;
      19223: inst = 32'hc40480d;
      19224: inst = 32'h8220000;
      19225: inst = 32'h10408000;
      19226: inst = 32'hc40480e;
      19227: inst = 32'h8220000;
      19228: inst = 32'h10408000;
      19229: inst = 32'hc40480f;
      19230: inst = 32'h8220000;
      19231: inst = 32'h10408000;
      19232: inst = 32'hc404810;
      19233: inst = 32'h8220000;
      19234: inst = 32'h10408000;
      19235: inst = 32'hc404811;
      19236: inst = 32'h8220000;
      19237: inst = 32'h10408000;
      19238: inst = 32'hc40482b;
      19239: inst = 32'h8220000;
      19240: inst = 32'h10408000;
      19241: inst = 32'hc40482c;
      19242: inst = 32'h8220000;
      19243: inst = 32'h10408000;
      19244: inst = 32'hc40482e;
      19245: inst = 32'h8220000;
      19246: inst = 32'h10408000;
      19247: inst = 32'hc40482f;
      19248: inst = 32'h8220000;
      19249: inst = 32'h10408000;
      19250: inst = 32'hc404830;
      19251: inst = 32'h8220000;
      19252: inst = 32'h10408000;
      19253: inst = 32'hc404831;
      19254: inst = 32'h8220000;
      19255: inst = 32'h10408000;
      19256: inst = 32'hc404832;
      19257: inst = 32'h8220000;
      19258: inst = 32'h10408000;
      19259: inst = 32'hc404837;
      19260: inst = 32'h8220000;
      19261: inst = 32'h10408000;
      19262: inst = 32'hc404838;
      19263: inst = 32'h8220000;
      19264: inst = 32'h10408000;
      19265: inst = 32'hc40483a;
      19266: inst = 32'h8220000;
      19267: inst = 32'h10408000;
      19268: inst = 32'hc40483b;
      19269: inst = 32'h8220000;
      19270: inst = 32'h10408000;
      19271: inst = 32'hc40483c;
      19272: inst = 32'h8220000;
      19273: inst = 32'h10408000;
      19274: inst = 32'hc40483d;
      19275: inst = 32'h8220000;
      19276: inst = 32'h10408000;
      19277: inst = 32'hc40483e;
      19278: inst = 32'h8220000;
      19279: inst = 32'h10408000;
      19280: inst = 32'hc404846;
      19281: inst = 32'h8220000;
      19282: inst = 32'h10408000;
      19283: inst = 32'hc404847;
      19284: inst = 32'h8220000;
      19285: inst = 32'h10408000;
      19286: inst = 32'hc404848;
      19287: inst = 32'h8220000;
      19288: inst = 32'h10408000;
      19289: inst = 32'hc404850;
      19290: inst = 32'h8220000;
      19291: inst = 32'h10408000;
      19292: inst = 32'hc404851;
      19293: inst = 32'h8220000;
      19294: inst = 32'h10408000;
      19295: inst = 32'hc404859;
      19296: inst = 32'h8220000;
      19297: inst = 32'h10408000;
      19298: inst = 32'hc40485a;
      19299: inst = 32'h8220000;
      19300: inst = 32'h10408000;
      19301: inst = 32'hc40485f;
      19302: inst = 32'h8220000;
      19303: inst = 32'h10408000;
      19304: inst = 32'hc404860;
      19305: inst = 32'h8220000;
      19306: inst = 32'h10408000;
      19307: inst = 32'hc404861;
      19308: inst = 32'h8220000;
      19309: inst = 32'h10408000;
      19310: inst = 32'hc404862;
      19311: inst = 32'h8220000;
      19312: inst = 32'h10408000;
      19313: inst = 32'hc404869;
      19314: inst = 32'h8220000;
      19315: inst = 32'h10408000;
      19316: inst = 32'hc40486a;
      19317: inst = 32'h8220000;
      19318: inst = 32'h10408000;
      19319: inst = 32'hc40486c;
      19320: inst = 32'h8220000;
      19321: inst = 32'h10408000;
      19322: inst = 32'hc40486d;
      19323: inst = 32'h8220000;
      19324: inst = 32'h10408000;
      19325: inst = 32'hc40486e;
      19326: inst = 32'h8220000;
      19327: inst = 32'h10408000;
      19328: inst = 32'hc40486f;
      19329: inst = 32'h8220000;
      19330: inst = 32'h10408000;
      19331: inst = 32'hc404870;
      19332: inst = 32'h8220000;
      19333: inst = 32'h10408000;
      19334: inst = 32'hc404871;
      19335: inst = 32'h8220000;
      19336: inst = 32'h10408000;
      19337: inst = 32'hc404872;
      19338: inst = 32'h8220000;
      19339: inst = 32'h10408000;
      19340: inst = 32'hc40488b;
      19341: inst = 32'h8220000;
      19342: inst = 32'h10408000;
      19343: inst = 32'hc40488c;
      19344: inst = 32'h8220000;
      19345: inst = 32'h10408000;
      19346: inst = 32'hc404897;
      19347: inst = 32'h8220000;
      19348: inst = 32'h10408000;
      19349: inst = 32'hc404898;
      19350: inst = 32'h8220000;
      19351: inst = 32'h10408000;
      19352: inst = 32'hc4048a6;
      19353: inst = 32'h8220000;
      19354: inst = 32'h10408000;
      19355: inst = 32'hc4048b0;
      19356: inst = 32'h8220000;
      19357: inst = 32'h10408000;
      19358: inst = 32'hc4048b1;
      19359: inst = 32'h8220000;
      19360: inst = 32'h10408000;
      19361: inst = 32'hc4048b4;
      19362: inst = 32'h8220000;
      19363: inst = 32'h10408000;
      19364: inst = 32'hc4048b5;
      19365: inst = 32'h8220000;
      19366: inst = 32'h10408000;
      19367: inst = 32'hc4048b9;
      19368: inst = 32'h8220000;
      19369: inst = 32'h10408000;
      19370: inst = 32'hc4048ba;
      19371: inst = 32'h8220000;
      19372: inst = 32'h10408000;
      19373: inst = 32'hc4048bf;
      19374: inst = 32'h8220000;
      19375: inst = 32'h10408000;
      19376: inst = 32'hc4048c9;
      19377: inst = 32'h8220000;
      19378: inst = 32'h10408000;
      19379: inst = 32'hc4048ca;
      19380: inst = 32'h8220000;
      19381: inst = 32'h10408000;
      19382: inst = 32'hc4048d1;
      19383: inst = 32'h8220000;
      19384: inst = 32'h10408000;
      19385: inst = 32'hc4048d2;
      19386: inst = 32'h8220000;
      19387: inst = 32'h10408000;
      19388: inst = 32'hc4048d3;
      19389: inst = 32'h8220000;
      19390: inst = 32'h10408000;
      19391: inst = 32'hc4048eb;
      19392: inst = 32'h8220000;
      19393: inst = 32'h10408000;
      19394: inst = 32'hc4048ec;
      19395: inst = 32'h8220000;
      19396: inst = 32'h10408000;
      19397: inst = 32'hc4048ed;
      19398: inst = 32'h8220000;
      19399: inst = 32'h10408000;
      19400: inst = 32'hc4048ee;
      19401: inst = 32'h8220000;
      19402: inst = 32'h10408000;
      19403: inst = 32'hc4048ef;
      19404: inst = 32'h8220000;
      19405: inst = 32'h10408000;
      19406: inst = 32'hc4048f0;
      19407: inst = 32'h8220000;
      19408: inst = 32'h10408000;
      19409: inst = 32'hc4048f1;
      19410: inst = 32'h8220000;
      19411: inst = 32'h10408000;
      19412: inst = 32'hc4048f2;
      19413: inst = 32'h8220000;
      19414: inst = 32'h10408000;
      19415: inst = 32'hc4048f3;
      19416: inst = 32'h8220000;
      19417: inst = 32'h10408000;
      19418: inst = 32'hc4048f4;
      19419: inst = 32'h8220000;
      19420: inst = 32'h10408000;
      19421: inst = 32'hc4048f5;
      19422: inst = 32'h8220000;
      19423: inst = 32'h10408000;
      19424: inst = 32'hc4048f7;
      19425: inst = 32'h8220000;
      19426: inst = 32'h10408000;
      19427: inst = 32'hc4048f8;
      19428: inst = 32'h8220000;
      19429: inst = 32'h10408000;
      19430: inst = 32'hc4048f9;
      19431: inst = 32'h8220000;
      19432: inst = 32'h10408000;
      19433: inst = 32'hc4048fa;
      19434: inst = 32'h8220000;
      19435: inst = 32'h10408000;
      19436: inst = 32'hc4048fb;
      19437: inst = 32'h8220000;
      19438: inst = 32'h10408000;
      19439: inst = 32'hc4048fc;
      19440: inst = 32'h8220000;
      19441: inst = 32'h10408000;
      19442: inst = 32'hc4048fd;
      19443: inst = 32'h8220000;
      19444: inst = 32'h10408000;
      19445: inst = 32'hc4048fe;
      19446: inst = 32'h8220000;
      19447: inst = 32'h10408000;
      19448: inst = 32'hc4048ff;
      19449: inst = 32'h8220000;
      19450: inst = 32'h10408000;
      19451: inst = 32'hc404900;
      19452: inst = 32'h8220000;
      19453: inst = 32'h10408000;
      19454: inst = 32'hc404901;
      19455: inst = 32'h8220000;
      19456: inst = 32'h10408000;
      19457: inst = 32'hc404904;
      19458: inst = 32'h8220000;
      19459: inst = 32'h10408000;
      19460: inst = 32'hc404905;
      19461: inst = 32'h8220000;
      19462: inst = 32'h10408000;
      19463: inst = 32'hc404906;
      19464: inst = 32'h8220000;
      19465: inst = 32'h10408000;
      19466: inst = 32'hc404907;
      19467: inst = 32'h8220000;
      19468: inst = 32'h10408000;
      19469: inst = 32'hc404908;
      19470: inst = 32'h8220000;
      19471: inst = 32'h10408000;
      19472: inst = 32'hc404909;
      19473: inst = 32'h8220000;
      19474: inst = 32'h10408000;
      19475: inst = 32'hc40490a;
      19476: inst = 32'h8220000;
      19477: inst = 32'h10408000;
      19478: inst = 32'hc40490b;
      19479: inst = 32'h8220000;
      19480: inst = 32'h10408000;
      19481: inst = 32'hc40490c;
      19482: inst = 32'h8220000;
      19483: inst = 32'h10408000;
      19484: inst = 32'hc40490d;
      19485: inst = 32'h8220000;
      19486: inst = 32'h10408000;
      19487: inst = 32'hc404910;
      19488: inst = 32'h8220000;
      19489: inst = 32'h10408000;
      19490: inst = 32'hc404911;
      19491: inst = 32'h8220000;
      19492: inst = 32'h10408000;
      19493: inst = 32'hc404912;
      19494: inst = 32'h8220000;
      19495: inst = 32'h10408000;
      19496: inst = 32'hc404913;
      19497: inst = 32'h8220000;
      19498: inst = 32'h10408000;
      19499: inst = 32'hc404914;
      19500: inst = 32'h8220000;
      19501: inst = 32'h10408000;
      19502: inst = 32'hc404915;
      19503: inst = 32'h8220000;
      19504: inst = 32'h10408000;
      19505: inst = 32'hc404916;
      19506: inst = 32'h8220000;
      19507: inst = 32'h10408000;
      19508: inst = 32'hc404917;
      19509: inst = 32'h8220000;
      19510: inst = 32'h10408000;
      19511: inst = 32'hc404918;
      19512: inst = 32'h8220000;
      19513: inst = 32'h10408000;
      19514: inst = 32'hc404919;
      19515: inst = 32'h8220000;
      19516: inst = 32'h10408000;
      19517: inst = 32'hc40491a;
      19518: inst = 32'h8220000;
      19519: inst = 32'h10408000;
      19520: inst = 32'hc40491e;
      19521: inst = 32'h8220000;
      19522: inst = 32'h10408000;
      19523: inst = 32'hc40491f;
      19524: inst = 32'h8220000;
      19525: inst = 32'h10408000;
      19526: inst = 32'hc404920;
      19527: inst = 32'h8220000;
      19528: inst = 32'h10408000;
      19529: inst = 32'hc404921;
      19530: inst = 32'h8220000;
      19531: inst = 32'h10408000;
      19532: inst = 32'hc404922;
      19533: inst = 32'h8220000;
      19534: inst = 32'h10408000;
      19535: inst = 32'hc404923;
      19536: inst = 32'h8220000;
      19537: inst = 32'h10408000;
      19538: inst = 32'hc404924;
      19539: inst = 32'h8220000;
      19540: inst = 32'h10408000;
      19541: inst = 32'hc404925;
      19542: inst = 32'h8220000;
      19543: inst = 32'h10408000;
      19544: inst = 32'hc404926;
      19545: inst = 32'h8220000;
      19546: inst = 32'h10408000;
      19547: inst = 32'hc404927;
      19548: inst = 32'h8220000;
      19549: inst = 32'h10408000;
      19550: inst = 32'hc404929;
      19551: inst = 32'h8220000;
      19552: inst = 32'h10408000;
      19553: inst = 32'hc40492a;
      19554: inst = 32'h8220000;
      19555: inst = 32'h10408000;
      19556: inst = 32'hc40492b;
      19557: inst = 32'h8220000;
      19558: inst = 32'h10408000;
      19559: inst = 32'hc40492c;
      19560: inst = 32'h8220000;
      19561: inst = 32'h10408000;
      19562: inst = 32'hc40492d;
      19563: inst = 32'h8220000;
      19564: inst = 32'h10408000;
      19565: inst = 32'hc40492e;
      19566: inst = 32'h8220000;
      19567: inst = 32'h10408000;
      19568: inst = 32'hc40492f;
      19569: inst = 32'h8220000;
      19570: inst = 32'h10408000;
      19571: inst = 32'hc404930;
      19572: inst = 32'h8220000;
      19573: inst = 32'h10408000;
      19574: inst = 32'hc404931;
      19575: inst = 32'h8220000;
      19576: inst = 32'h10408000;
      19577: inst = 32'hc404932;
      19578: inst = 32'h8220000;
      19579: inst = 32'h10408000;
      19580: inst = 32'hc404933;
      19581: inst = 32'h8220000;
      19582: inst = 32'h10408000;
      19583: inst = 32'hc40494b;
      19584: inst = 32'h8220000;
      19585: inst = 32'h10408000;
      19586: inst = 32'hc40494c;
      19587: inst = 32'h8220000;
      19588: inst = 32'h10408000;
      19589: inst = 32'hc40494d;
      19590: inst = 32'h8220000;
      19591: inst = 32'h10408000;
      19592: inst = 32'hc40494e;
      19593: inst = 32'h8220000;
      19594: inst = 32'h10408000;
      19595: inst = 32'hc40494f;
      19596: inst = 32'h8220000;
      19597: inst = 32'h10408000;
      19598: inst = 32'hc404950;
      19599: inst = 32'h8220000;
      19600: inst = 32'h10408000;
      19601: inst = 32'hc404951;
      19602: inst = 32'h8220000;
      19603: inst = 32'h10408000;
      19604: inst = 32'hc404952;
      19605: inst = 32'h8220000;
      19606: inst = 32'h10408000;
      19607: inst = 32'hc404953;
      19608: inst = 32'h8220000;
      19609: inst = 32'h10408000;
      19610: inst = 32'hc404954;
      19611: inst = 32'h8220000;
      19612: inst = 32'h10408000;
      19613: inst = 32'hc404957;
      19614: inst = 32'h8220000;
      19615: inst = 32'h10408000;
      19616: inst = 32'hc404958;
      19617: inst = 32'h8220000;
      19618: inst = 32'h10408000;
      19619: inst = 32'hc404959;
      19620: inst = 32'h8220000;
      19621: inst = 32'h10408000;
      19622: inst = 32'hc40495a;
      19623: inst = 32'h8220000;
      19624: inst = 32'h10408000;
      19625: inst = 32'hc40495b;
      19626: inst = 32'h8220000;
      19627: inst = 32'h10408000;
      19628: inst = 32'hc40495c;
      19629: inst = 32'h8220000;
      19630: inst = 32'h10408000;
      19631: inst = 32'hc40495d;
      19632: inst = 32'h8220000;
      19633: inst = 32'h10408000;
      19634: inst = 32'hc40495e;
      19635: inst = 32'h8220000;
      19636: inst = 32'h10408000;
      19637: inst = 32'hc40495f;
      19638: inst = 32'h8220000;
      19639: inst = 32'h10408000;
      19640: inst = 32'hc404960;
      19641: inst = 32'h8220000;
      19642: inst = 32'h10408000;
      19643: inst = 32'hc404961;
      19644: inst = 32'h8220000;
      19645: inst = 32'h10408000;
      19646: inst = 32'hc404963;
      19647: inst = 32'h8220000;
      19648: inst = 32'h10408000;
      19649: inst = 32'hc404964;
      19650: inst = 32'h8220000;
      19651: inst = 32'h10408000;
      19652: inst = 32'hc404965;
      19653: inst = 32'h8220000;
      19654: inst = 32'h10408000;
      19655: inst = 32'hc404966;
      19656: inst = 32'h8220000;
      19657: inst = 32'h10408000;
      19658: inst = 32'hc404967;
      19659: inst = 32'h8220000;
      19660: inst = 32'h10408000;
      19661: inst = 32'hc404968;
      19662: inst = 32'h8220000;
      19663: inst = 32'h10408000;
      19664: inst = 32'hc404969;
      19665: inst = 32'h8220000;
      19666: inst = 32'h10408000;
      19667: inst = 32'hc40496a;
      19668: inst = 32'h8220000;
      19669: inst = 32'h10408000;
      19670: inst = 32'hc40496b;
      19671: inst = 32'h8220000;
      19672: inst = 32'h10408000;
      19673: inst = 32'hc40496c;
      19674: inst = 32'h8220000;
      19675: inst = 32'h10408000;
      19676: inst = 32'hc40496d;
      19677: inst = 32'h8220000;
      19678: inst = 32'h10408000;
      19679: inst = 32'hc404970;
      19680: inst = 32'h8220000;
      19681: inst = 32'h10408000;
      19682: inst = 32'hc404971;
      19683: inst = 32'h8220000;
      19684: inst = 32'h10408000;
      19685: inst = 32'hc404972;
      19686: inst = 32'h8220000;
      19687: inst = 32'h10408000;
      19688: inst = 32'hc404973;
      19689: inst = 32'h8220000;
      19690: inst = 32'h10408000;
      19691: inst = 32'hc404974;
      19692: inst = 32'h8220000;
      19693: inst = 32'h10408000;
      19694: inst = 32'hc404975;
      19695: inst = 32'h8220000;
      19696: inst = 32'h10408000;
      19697: inst = 32'hc404976;
      19698: inst = 32'h8220000;
      19699: inst = 32'h10408000;
      19700: inst = 32'hc404977;
      19701: inst = 32'h8220000;
      19702: inst = 32'h10408000;
      19703: inst = 32'hc404978;
      19704: inst = 32'h8220000;
      19705: inst = 32'h10408000;
      19706: inst = 32'hc404979;
      19707: inst = 32'h8220000;
      19708: inst = 32'h10408000;
      19709: inst = 32'hc40497d;
      19710: inst = 32'h8220000;
      19711: inst = 32'h10408000;
      19712: inst = 32'hc40497e;
      19713: inst = 32'h8220000;
      19714: inst = 32'h10408000;
      19715: inst = 32'hc40497f;
      19716: inst = 32'h8220000;
      19717: inst = 32'h10408000;
      19718: inst = 32'hc404980;
      19719: inst = 32'h8220000;
      19720: inst = 32'h10408000;
      19721: inst = 32'hc404981;
      19722: inst = 32'h8220000;
      19723: inst = 32'h10408000;
      19724: inst = 32'hc404982;
      19725: inst = 32'h8220000;
      19726: inst = 32'h10408000;
      19727: inst = 32'hc404983;
      19728: inst = 32'h8220000;
      19729: inst = 32'h10408000;
      19730: inst = 32'hc404984;
      19731: inst = 32'h8220000;
      19732: inst = 32'h10408000;
      19733: inst = 32'hc404985;
      19734: inst = 32'h8220000;
      19735: inst = 32'h10408000;
      19736: inst = 32'hc404986;
      19737: inst = 32'h8220000;
      19738: inst = 32'h10408000;
      19739: inst = 32'hc404987;
      19740: inst = 32'h8220000;
      19741: inst = 32'h10408000;
      19742: inst = 32'hc404989;
      19743: inst = 32'h8220000;
      19744: inst = 32'h10408000;
      19745: inst = 32'hc40498a;
      19746: inst = 32'h8220000;
      19747: inst = 32'h10408000;
      19748: inst = 32'hc40498b;
      19749: inst = 32'h8220000;
      19750: inst = 32'h10408000;
      19751: inst = 32'hc40498c;
      19752: inst = 32'h8220000;
      19753: inst = 32'h10408000;
      19754: inst = 32'hc40498d;
      19755: inst = 32'h8220000;
      19756: inst = 32'h10408000;
      19757: inst = 32'hc40498e;
      19758: inst = 32'h8220000;
      19759: inst = 32'h10408000;
      19760: inst = 32'hc40498f;
      19761: inst = 32'h8220000;
      19762: inst = 32'h10408000;
      19763: inst = 32'hc404990;
      19764: inst = 32'h8220000;
      19765: inst = 32'h10408000;
      19766: inst = 32'hc404991;
      19767: inst = 32'h8220000;
      19768: inst = 32'h10408000;
      19769: inst = 32'hc404992;
      19770: inst = 32'h8220000;
      19771: inst = 32'h10408000;
      19772: inst = 32'hc404993;
      19773: inst = 32'h8220000;
      19774: inst = 32'h10408000;
      19775: inst = 32'hc404dcd;
      19776: inst = 32'h8220000;
      19777: inst = 32'h10408000;
      19778: inst = 32'hc404dce;
      19779: inst = 32'h8220000;
      19780: inst = 32'h10408000;
      19781: inst = 32'hc404dcf;
      19782: inst = 32'h8220000;
      19783: inst = 32'h10408000;
      19784: inst = 32'hc404dd0;
      19785: inst = 32'h8220000;
      19786: inst = 32'h10408000;
      19787: inst = 32'hc404dd1;
      19788: inst = 32'h8220000;
      19789: inst = 32'h10408000;
      19790: inst = 32'hc404dd2;
      19791: inst = 32'h8220000;
      19792: inst = 32'h10408000;
      19793: inst = 32'hc404dd3;
      19794: inst = 32'h8220000;
      19795: inst = 32'h10408000;
      19796: inst = 32'hc404dd4;
      19797: inst = 32'h8220000;
      19798: inst = 32'h10408000;
      19799: inst = 32'hc404dd5;
      19800: inst = 32'h8220000;
      19801: inst = 32'h10408000;
      19802: inst = 32'hc404dd7;
      19803: inst = 32'h8220000;
      19804: inst = 32'h10408000;
      19805: inst = 32'hc404dd8;
      19806: inst = 32'h8220000;
      19807: inst = 32'h10408000;
      19808: inst = 32'hc404dd9;
      19809: inst = 32'h8220000;
      19810: inst = 32'h10408000;
      19811: inst = 32'hc404dda;
      19812: inst = 32'h8220000;
      19813: inst = 32'h10408000;
      19814: inst = 32'hc404ddb;
      19815: inst = 32'h8220000;
      19816: inst = 32'h10408000;
      19817: inst = 32'hc404ddc;
      19818: inst = 32'h8220000;
      19819: inst = 32'h10408000;
      19820: inst = 32'hc404ddd;
      19821: inst = 32'h8220000;
      19822: inst = 32'h10408000;
      19823: inst = 32'hc404dde;
      19824: inst = 32'h8220000;
      19825: inst = 32'h10408000;
      19826: inst = 32'hc404ddf;
      19827: inst = 32'h8220000;
      19828: inst = 32'h10408000;
      19829: inst = 32'hc404de0;
      19830: inst = 32'h8220000;
      19831: inst = 32'h10408000;
      19832: inst = 32'hc404de1;
      19833: inst = 32'h8220000;
      19834: inst = 32'h10408000;
      19835: inst = 32'hc404de2;
      19836: inst = 32'h8220000;
      19837: inst = 32'h10408000;
      19838: inst = 32'hc404de4;
      19839: inst = 32'h8220000;
      19840: inst = 32'h10408000;
      19841: inst = 32'hc404de5;
      19842: inst = 32'h8220000;
      19843: inst = 32'h10408000;
      19844: inst = 32'hc404de6;
      19845: inst = 32'h8220000;
      19846: inst = 32'h10408000;
      19847: inst = 32'hc404de7;
      19848: inst = 32'h8220000;
      19849: inst = 32'h10408000;
      19850: inst = 32'hc404de8;
      19851: inst = 32'h8220000;
      19852: inst = 32'h10408000;
      19853: inst = 32'hc404de9;
      19854: inst = 32'h8220000;
      19855: inst = 32'h10408000;
      19856: inst = 32'hc404dea;
      19857: inst = 32'h8220000;
      19858: inst = 32'h10408000;
      19859: inst = 32'hc404deb;
      19860: inst = 32'h8220000;
      19861: inst = 32'h10408000;
      19862: inst = 32'hc404dec;
      19863: inst = 32'h8220000;
      19864: inst = 32'h10408000;
      19865: inst = 32'hc404ded;
      19866: inst = 32'h8220000;
      19867: inst = 32'h10408000;
      19868: inst = 32'hc404df0;
      19869: inst = 32'h8220000;
      19870: inst = 32'h10408000;
      19871: inst = 32'hc404df1;
      19872: inst = 32'h8220000;
      19873: inst = 32'h10408000;
      19874: inst = 32'hc404df2;
      19875: inst = 32'h8220000;
      19876: inst = 32'h10408000;
      19877: inst = 32'hc404dfc;
      19878: inst = 32'h8220000;
      19879: inst = 32'h10408000;
      19880: inst = 32'hc404dfd;
      19881: inst = 32'h8220000;
      19882: inst = 32'h10408000;
      19883: inst = 32'hc404dfe;
      19884: inst = 32'h8220000;
      19885: inst = 32'h10408000;
      19886: inst = 32'hc404dff;
      19887: inst = 32'h8220000;
      19888: inst = 32'h10408000;
      19889: inst = 32'hc404e00;
      19890: inst = 32'h8220000;
      19891: inst = 32'h10408000;
      19892: inst = 32'hc404e01;
      19893: inst = 32'h8220000;
      19894: inst = 32'h10408000;
      19895: inst = 32'hc404e02;
      19896: inst = 32'h8220000;
      19897: inst = 32'h10408000;
      19898: inst = 32'hc404e03;
      19899: inst = 32'h8220000;
      19900: inst = 32'h10408000;
      19901: inst = 32'hc404e04;
      19902: inst = 32'h8220000;
      19903: inst = 32'h10408000;
      19904: inst = 32'hc404e05;
      19905: inst = 32'h8220000;
      19906: inst = 32'h10408000;
      19907: inst = 32'hc404e06;
      19908: inst = 32'h8220000;
      19909: inst = 32'h10408000;
      19910: inst = 32'hc404e07;
      19911: inst = 32'h8220000;
      19912: inst = 32'h10408000;
      19913: inst = 32'hc404e0b;
      19914: inst = 32'h8220000;
      19915: inst = 32'h10408000;
      19916: inst = 32'hc404e0c;
      19917: inst = 32'h8220000;
      19918: inst = 32'h10408000;
      19919: inst = 32'hc404e0d;
      19920: inst = 32'h8220000;
      19921: inst = 32'h10408000;
      19922: inst = 32'hc404e0e;
      19923: inst = 32'h8220000;
      19924: inst = 32'h10408000;
      19925: inst = 32'hc404e0f;
      19926: inst = 32'h8220000;
      19927: inst = 32'h10408000;
      19928: inst = 32'hc404e10;
      19929: inst = 32'h8220000;
      19930: inst = 32'h10408000;
      19931: inst = 32'hc404e11;
      19932: inst = 32'h8220000;
      19933: inst = 32'h10408000;
      19934: inst = 32'hc404e12;
      19935: inst = 32'h8220000;
      19936: inst = 32'h10408000;
      19937: inst = 32'hc404e13;
      19938: inst = 32'h8220000;
      19939: inst = 32'h10408000;
      19940: inst = 32'hc404e2c;
      19941: inst = 32'h8220000;
      19942: inst = 32'h10408000;
      19943: inst = 32'hc404e2d;
      19944: inst = 32'h8220000;
      19945: inst = 32'h10408000;
      19946: inst = 32'hc404e2e;
      19947: inst = 32'h8220000;
      19948: inst = 32'h10408000;
      19949: inst = 32'hc404e2f;
      19950: inst = 32'h8220000;
      19951: inst = 32'h10408000;
      19952: inst = 32'hc404e30;
      19953: inst = 32'h8220000;
      19954: inst = 32'h10408000;
      19955: inst = 32'hc404e31;
      19956: inst = 32'h8220000;
      19957: inst = 32'h10408000;
      19958: inst = 32'hc404e32;
      19959: inst = 32'h8220000;
      19960: inst = 32'h10408000;
      19961: inst = 32'hc404e33;
      19962: inst = 32'h8220000;
      19963: inst = 32'h10408000;
      19964: inst = 32'hc404e34;
      19965: inst = 32'h8220000;
      19966: inst = 32'h10408000;
      19967: inst = 32'hc404e35;
      19968: inst = 32'h8220000;
      19969: inst = 32'h10408000;
      19970: inst = 32'hc404e38;
      19971: inst = 32'h8220000;
      19972: inst = 32'h10408000;
      19973: inst = 32'hc404e39;
      19974: inst = 32'h8220000;
      19975: inst = 32'h10408000;
      19976: inst = 32'hc404e3a;
      19977: inst = 32'h8220000;
      19978: inst = 32'h10408000;
      19979: inst = 32'hc404e3b;
      19980: inst = 32'h8220000;
      19981: inst = 32'h10408000;
      19982: inst = 32'hc404e3c;
      19983: inst = 32'h8220000;
      19984: inst = 32'h10408000;
      19985: inst = 32'hc404e3d;
      19986: inst = 32'h8220000;
      19987: inst = 32'h10408000;
      19988: inst = 32'hc404e3e;
      19989: inst = 32'h8220000;
      19990: inst = 32'h10408000;
      19991: inst = 32'hc404e3f;
      19992: inst = 32'h8220000;
      19993: inst = 32'h10408000;
      19994: inst = 32'hc404e40;
      19995: inst = 32'h8220000;
      19996: inst = 32'h10408000;
      19997: inst = 32'hc404e41;
      19998: inst = 32'h8220000;
      19999: inst = 32'h10408000;
      20000: inst = 32'hc404e42;
      20001: inst = 32'h8220000;
      20002: inst = 32'h10408000;
      20003: inst = 32'hc404e44;
      20004: inst = 32'h8220000;
      20005: inst = 32'h10408000;
      20006: inst = 32'hc404e45;
      20007: inst = 32'h8220000;
      20008: inst = 32'h10408000;
      20009: inst = 32'hc404e46;
      20010: inst = 32'h8220000;
      20011: inst = 32'h10408000;
      20012: inst = 32'hc404e47;
      20013: inst = 32'h8220000;
      20014: inst = 32'h10408000;
      20015: inst = 32'hc404e48;
      20016: inst = 32'h8220000;
      20017: inst = 32'h10408000;
      20018: inst = 32'hc404e49;
      20019: inst = 32'h8220000;
      20020: inst = 32'h10408000;
      20021: inst = 32'hc404e4a;
      20022: inst = 32'h8220000;
      20023: inst = 32'h10408000;
      20024: inst = 32'hc404e4b;
      20025: inst = 32'h8220000;
      20026: inst = 32'h10408000;
      20027: inst = 32'hc404e4c;
      20028: inst = 32'h8220000;
      20029: inst = 32'h10408000;
      20030: inst = 32'hc404e4d;
      20031: inst = 32'h8220000;
      20032: inst = 32'h10408000;
      20033: inst = 32'hc404e50;
      20034: inst = 32'h8220000;
      20035: inst = 32'h10408000;
      20036: inst = 32'hc404e51;
      20037: inst = 32'h8220000;
      20038: inst = 32'h10408000;
      20039: inst = 32'hc404e52;
      20040: inst = 32'h8220000;
      20041: inst = 32'h10408000;
      20042: inst = 32'hc404e53;
      20043: inst = 32'h8220000;
      20044: inst = 32'h10408000;
      20045: inst = 32'hc404e5c;
      20046: inst = 32'h8220000;
      20047: inst = 32'h10408000;
      20048: inst = 32'hc404e5d;
      20049: inst = 32'h8220000;
      20050: inst = 32'h10408000;
      20051: inst = 32'hc404e5e;
      20052: inst = 32'h8220000;
      20053: inst = 32'h10408000;
      20054: inst = 32'hc404e5f;
      20055: inst = 32'h8220000;
      20056: inst = 32'h10408000;
      20057: inst = 32'hc404e60;
      20058: inst = 32'h8220000;
      20059: inst = 32'h10408000;
      20060: inst = 32'hc404e61;
      20061: inst = 32'h8220000;
      20062: inst = 32'h10408000;
      20063: inst = 32'hc404e62;
      20064: inst = 32'h8220000;
      20065: inst = 32'h10408000;
      20066: inst = 32'hc404e63;
      20067: inst = 32'h8220000;
      20068: inst = 32'h10408000;
      20069: inst = 32'hc404e64;
      20070: inst = 32'h8220000;
      20071: inst = 32'h10408000;
      20072: inst = 32'hc404e65;
      20073: inst = 32'h8220000;
      20074: inst = 32'h10408000;
      20075: inst = 32'hc404e66;
      20076: inst = 32'h8220000;
      20077: inst = 32'h10408000;
      20078: inst = 32'hc404e6a;
      20079: inst = 32'h8220000;
      20080: inst = 32'h10408000;
      20081: inst = 32'hc404e6b;
      20082: inst = 32'h8220000;
      20083: inst = 32'h10408000;
      20084: inst = 32'hc404e6c;
      20085: inst = 32'h8220000;
      20086: inst = 32'h10408000;
      20087: inst = 32'hc404e6d;
      20088: inst = 32'h8220000;
      20089: inst = 32'h10408000;
      20090: inst = 32'hc404e6e;
      20091: inst = 32'h8220000;
      20092: inst = 32'h10408000;
      20093: inst = 32'hc404e6f;
      20094: inst = 32'h8220000;
      20095: inst = 32'h10408000;
      20096: inst = 32'hc404e70;
      20097: inst = 32'h8220000;
      20098: inst = 32'h10408000;
      20099: inst = 32'hc404e71;
      20100: inst = 32'h8220000;
      20101: inst = 32'h10408000;
      20102: inst = 32'hc404e72;
      20103: inst = 32'h8220000;
      20104: inst = 32'h10408000;
      20105: inst = 32'hc404e73;
      20106: inst = 32'h8220000;
      20107: inst = 32'h10408000;
      20108: inst = 32'hc404e8b;
      20109: inst = 32'h8220000;
      20110: inst = 32'h10408000;
      20111: inst = 32'hc404e8c;
      20112: inst = 32'h8220000;
      20113: inst = 32'h10408000;
      20114: inst = 32'hc404e8d;
      20115: inst = 32'h8220000;
      20116: inst = 32'h10408000;
      20117: inst = 32'hc404e99;
      20118: inst = 32'h8220000;
      20119: inst = 32'h10408000;
      20120: inst = 32'hc404e9a;
      20121: inst = 32'h8220000;
      20122: inst = 32'h10408000;
      20123: inst = 32'hc404e9b;
      20124: inst = 32'h8220000;
      20125: inst = 32'h10408000;
      20126: inst = 32'hc404e9c;
      20127: inst = 32'h8220000;
      20128: inst = 32'h10408000;
      20129: inst = 32'hc404ea4;
      20130: inst = 32'h8220000;
      20131: inst = 32'h10408000;
      20132: inst = 32'hc404ea5;
      20133: inst = 32'h8220000;
      20134: inst = 32'h10408000;
      20135: inst = 32'hc404eac;
      20136: inst = 32'h8220000;
      20137: inst = 32'h10408000;
      20138: inst = 32'hc404ead;
      20139: inst = 32'h8220000;
      20140: inst = 32'h10408000;
      20141: inst = 32'hc404eb0;
      20142: inst = 32'h8220000;
      20143: inst = 32'h10408000;
      20144: inst = 32'hc404eb1;
      20145: inst = 32'h8220000;
      20146: inst = 32'h10408000;
      20147: inst = 32'hc404eb2;
      20148: inst = 32'h8220000;
      20149: inst = 32'h10408000;
      20150: inst = 32'hc404eb3;
      20151: inst = 32'h8220000;
      20152: inst = 32'h10408000;
      20153: inst = 32'hc404eb4;
      20154: inst = 32'h8220000;
      20155: inst = 32'h10408000;
      20156: inst = 32'hc404ebc;
      20157: inst = 32'h8220000;
      20158: inst = 32'h10408000;
      20159: inst = 32'hc404ebd;
      20160: inst = 32'h8220000;
      20161: inst = 32'h10408000;
      20162: inst = 32'hc404ec2;
      20163: inst = 32'h8220000;
      20164: inst = 32'h10408000;
      20165: inst = 32'hc404ec3;
      20166: inst = 32'h8220000;
      20167: inst = 32'h10408000;
      20168: inst = 32'hc404ec4;
      20169: inst = 32'h8220000;
      20170: inst = 32'h10408000;
      20171: inst = 32'hc404ec5;
      20172: inst = 32'h8220000;
      20173: inst = 32'h10408000;
      20174: inst = 32'hc404ec9;
      20175: inst = 32'h8220000;
      20176: inst = 32'h10408000;
      20177: inst = 32'hc404eca;
      20178: inst = 32'h8220000;
      20179: inst = 32'h10408000;
      20180: inst = 32'hc404eeb;
      20181: inst = 32'h8220000;
      20182: inst = 32'h10408000;
      20183: inst = 32'hc404eec;
      20184: inst = 32'h8220000;
      20185: inst = 32'h10408000;
      20186: inst = 32'hc404efa;
      20187: inst = 32'h8220000;
      20188: inst = 32'h10408000;
      20189: inst = 32'hc404efb;
      20190: inst = 32'h8220000;
      20191: inst = 32'h10408000;
      20192: inst = 32'hc404efc;
      20193: inst = 32'h8220000;
      20194: inst = 32'h10408000;
      20195: inst = 32'hc404f04;
      20196: inst = 32'h8220000;
      20197: inst = 32'h10408000;
      20198: inst = 32'hc404f05;
      20199: inst = 32'h8220000;
      20200: inst = 32'h10408000;
      20201: inst = 32'hc404f0c;
      20202: inst = 32'h8220000;
      20203: inst = 32'h10408000;
      20204: inst = 32'hc404f0d;
      20205: inst = 32'h8220000;
      20206: inst = 32'h10408000;
      20207: inst = 32'hc404f10;
      20208: inst = 32'h8220000;
      20209: inst = 32'h10408000;
      20210: inst = 32'hc404f12;
      20211: inst = 32'h8220000;
      20212: inst = 32'h10408000;
      20213: inst = 32'hc404f13;
      20214: inst = 32'h8220000;
      20215: inst = 32'h10408000;
      20216: inst = 32'hc404f14;
      20217: inst = 32'h8220000;
      20218: inst = 32'h10408000;
      20219: inst = 32'hc404f15;
      20220: inst = 32'h8220000;
      20221: inst = 32'h10408000;
      20222: inst = 32'hc404f1c;
      20223: inst = 32'h8220000;
      20224: inst = 32'h10408000;
      20225: inst = 32'hc404f1d;
      20226: inst = 32'h8220000;
      20227: inst = 32'h10408000;
      20228: inst = 32'hc404f22;
      20229: inst = 32'h8220000;
      20230: inst = 32'h10408000;
      20231: inst = 32'hc404f23;
      20232: inst = 32'h8220000;
      20233: inst = 32'h10408000;
      20234: inst = 32'hc404f24;
      20235: inst = 32'h8220000;
      20236: inst = 32'h10408000;
      20237: inst = 32'hc404f29;
      20238: inst = 32'h8220000;
      20239: inst = 32'h10408000;
      20240: inst = 32'hc404f2a;
      20241: inst = 32'h8220000;
      20242: inst = 32'h10408000;
      20243: inst = 32'hc404f4b;
      20244: inst = 32'h8220000;
      20245: inst = 32'h10408000;
      20246: inst = 32'hc404f4c;
      20247: inst = 32'h8220000;
      20248: inst = 32'h10408000;
      20249: inst = 32'hc404f4e;
      20250: inst = 32'h8220000;
      20251: inst = 32'h10408000;
      20252: inst = 32'hc404f4f;
      20253: inst = 32'h8220000;
      20254: inst = 32'h10408000;
      20255: inst = 32'hc404f50;
      20256: inst = 32'h8220000;
      20257: inst = 32'h10408000;
      20258: inst = 32'hc404f51;
      20259: inst = 32'h8220000;
      20260: inst = 32'h10408000;
      20261: inst = 32'hc404f52;
      20262: inst = 32'h8220000;
      20263: inst = 32'h10408000;
      20264: inst = 32'hc404f5b;
      20265: inst = 32'h8220000;
      20266: inst = 32'h10408000;
      20267: inst = 32'hc404f5c;
      20268: inst = 32'h8220000;
      20269: inst = 32'h10408000;
      20270: inst = 32'hc404f5d;
      20271: inst = 32'h8220000;
      20272: inst = 32'h10408000;
      20273: inst = 32'hc404f64;
      20274: inst = 32'h8220000;
      20275: inst = 32'h10408000;
      20276: inst = 32'hc404f65;
      20277: inst = 32'h8220000;
      20278: inst = 32'h10408000;
      20279: inst = 32'hc404f6c;
      20280: inst = 32'h8220000;
      20281: inst = 32'h10408000;
      20282: inst = 32'hc404f70;
      20283: inst = 32'h8220000;
      20284: inst = 32'h10408000;
      20285: inst = 32'hc404f71;
      20286: inst = 32'h8220000;
      20287: inst = 32'h10408000;
      20288: inst = 32'hc404f72;
      20289: inst = 32'h8220000;
      20290: inst = 32'h10408000;
      20291: inst = 32'hc404f73;
      20292: inst = 32'h8220000;
      20293: inst = 32'h10408000;
      20294: inst = 32'hc404f74;
      20295: inst = 32'h8220000;
      20296: inst = 32'h10408000;
      20297: inst = 32'hc404f75;
      20298: inst = 32'h8220000;
      20299: inst = 32'h10408000;
      20300: inst = 32'hc404f76;
      20301: inst = 32'h8220000;
      20302: inst = 32'h10408000;
      20303: inst = 32'hc404f7c;
      20304: inst = 32'h8220000;
      20305: inst = 32'h10408000;
      20306: inst = 32'hc404f7d;
      20307: inst = 32'h8220000;
      20308: inst = 32'h10408000;
      20309: inst = 32'hc404f7f;
      20310: inst = 32'h8220000;
      20311: inst = 32'h10408000;
      20312: inst = 32'hc404f80;
      20313: inst = 32'h8220000;
      20314: inst = 32'h10408000;
      20315: inst = 32'hc404f81;
      20316: inst = 32'h8220000;
      20317: inst = 32'h10408000;
      20318: inst = 32'hc404f82;
      20319: inst = 32'h8220000;
      20320: inst = 32'h10408000;
      20321: inst = 32'hc404f83;
      20322: inst = 32'h8220000;
      20323: inst = 32'h10408000;
      20324: inst = 32'hc404f89;
      20325: inst = 32'h8220000;
      20326: inst = 32'h10408000;
      20327: inst = 32'hc404f8a;
      20328: inst = 32'h8220000;
      20329: inst = 32'h10408000;
      20330: inst = 32'hc404f8c;
      20331: inst = 32'h8220000;
      20332: inst = 32'h10408000;
      20333: inst = 32'hc404f8d;
      20334: inst = 32'h8220000;
      20335: inst = 32'h10408000;
      20336: inst = 32'hc404f8e;
      20337: inst = 32'h8220000;
      20338: inst = 32'h10408000;
      20339: inst = 32'hc404f8f;
      20340: inst = 32'h8220000;
      20341: inst = 32'h10408000;
      20342: inst = 32'hc404f90;
      20343: inst = 32'h8220000;
      20344: inst = 32'h10408000;
      20345: inst = 32'hc404fab;
      20346: inst = 32'h8220000;
      20347: inst = 32'h10408000;
      20348: inst = 32'hc404fac;
      20349: inst = 32'h8220000;
      20350: inst = 32'h10408000;
      20351: inst = 32'hc404fae;
      20352: inst = 32'h8220000;
      20353: inst = 32'h10408000;
      20354: inst = 32'hc404faf;
      20355: inst = 32'h8220000;
      20356: inst = 32'h10408000;
      20357: inst = 32'hc404fb0;
      20358: inst = 32'h8220000;
      20359: inst = 32'h10408000;
      20360: inst = 32'hc404fb1;
      20361: inst = 32'h8220000;
      20362: inst = 32'h10408000;
      20363: inst = 32'hc404fb2;
      20364: inst = 32'h8220000;
      20365: inst = 32'h10408000;
      20366: inst = 32'hc404fbc;
      20367: inst = 32'h8220000;
      20368: inst = 32'h10408000;
      20369: inst = 32'hc404fbd;
      20370: inst = 32'h8220000;
      20371: inst = 32'h10408000;
      20372: inst = 32'hc404fbe;
      20373: inst = 32'h8220000;
      20374: inst = 32'h10408000;
      20375: inst = 32'hc404fc4;
      20376: inst = 32'h8220000;
      20377: inst = 32'h10408000;
      20378: inst = 32'hc404fc5;
      20379: inst = 32'h8220000;
      20380: inst = 32'h10408000;
      20381: inst = 32'hc404fd0;
      20382: inst = 32'h8220000;
      20383: inst = 32'h10408000;
      20384: inst = 32'hc404fd1;
      20385: inst = 32'h8220000;
      20386: inst = 32'h10408000;
      20387: inst = 32'hc404fd2;
      20388: inst = 32'h8220000;
      20389: inst = 32'h10408000;
      20390: inst = 32'hc404fd4;
      20391: inst = 32'h8220000;
      20392: inst = 32'h10408000;
      20393: inst = 32'hc404fd5;
      20394: inst = 32'h8220000;
      20395: inst = 32'h10408000;
      20396: inst = 32'hc404fd6;
      20397: inst = 32'h8220000;
      20398: inst = 32'h10408000;
      20399: inst = 32'hc404fd7;
      20400: inst = 32'h8220000;
      20401: inst = 32'h10408000;
      20402: inst = 32'hc404fdc;
      20403: inst = 32'h8220000;
      20404: inst = 32'h10408000;
      20405: inst = 32'hc404fdd;
      20406: inst = 32'h8220000;
      20407: inst = 32'h10408000;
      20408: inst = 32'hc404fdf;
      20409: inst = 32'h8220000;
      20410: inst = 32'h10408000;
      20411: inst = 32'hc404fe0;
      20412: inst = 32'h8220000;
      20413: inst = 32'h10408000;
      20414: inst = 32'hc404fe1;
      20415: inst = 32'h8220000;
      20416: inst = 32'h10408000;
      20417: inst = 32'hc404fe2;
      20418: inst = 32'h8220000;
      20419: inst = 32'h10408000;
      20420: inst = 32'hc404fe9;
      20421: inst = 32'h8220000;
      20422: inst = 32'h10408000;
      20423: inst = 32'hc404fea;
      20424: inst = 32'h8220000;
      20425: inst = 32'h10408000;
      20426: inst = 32'hc404fec;
      20427: inst = 32'h8220000;
      20428: inst = 32'h10408000;
      20429: inst = 32'hc404fed;
      20430: inst = 32'h8220000;
      20431: inst = 32'h10408000;
      20432: inst = 32'hc404fee;
      20433: inst = 32'h8220000;
      20434: inst = 32'h10408000;
      20435: inst = 32'hc404fef;
      20436: inst = 32'h8220000;
      20437: inst = 32'h10408000;
      20438: inst = 32'hc404ff0;
      20439: inst = 32'h8220000;
      20440: inst = 32'h10408000;
      20441: inst = 32'hc40500b;
      20442: inst = 32'h8220000;
      20443: inst = 32'h10408000;
      20444: inst = 32'hc40500c;
      20445: inst = 32'h8220000;
      20446: inst = 32'h10408000;
      20447: inst = 32'hc40501d;
      20448: inst = 32'h8220000;
      20449: inst = 32'h10408000;
      20450: inst = 32'hc40501e;
      20451: inst = 32'h8220000;
      20452: inst = 32'h10408000;
      20453: inst = 32'hc40501f;
      20454: inst = 32'h8220000;
      20455: inst = 32'h10408000;
      20456: inst = 32'hc405024;
      20457: inst = 32'h8220000;
      20458: inst = 32'h10408000;
      20459: inst = 32'hc405025;
      20460: inst = 32'h8220000;
      20461: inst = 32'h10408000;
      20462: inst = 32'hc405030;
      20463: inst = 32'h8220000;
      20464: inst = 32'h10408000;
      20465: inst = 32'hc405031;
      20466: inst = 32'h8220000;
      20467: inst = 32'h10408000;
      20468: inst = 32'hc405032;
      20469: inst = 32'h8220000;
      20470: inst = 32'h10408000;
      20471: inst = 32'hc405033;
      20472: inst = 32'h8220000;
      20473: inst = 32'h10408000;
      20474: inst = 32'hc405034;
      20475: inst = 32'h8220000;
      20476: inst = 32'h10408000;
      20477: inst = 32'hc405035;
      20478: inst = 32'h8220000;
      20479: inst = 32'h10408000;
      20480: inst = 32'hc405036;
      20481: inst = 32'h8220000;
      20482: inst = 32'h10408000;
      20483: inst = 32'hc405037;
      20484: inst = 32'h8220000;
      20485: inst = 32'h10408000;
      20486: inst = 32'hc405038;
      20487: inst = 32'h8220000;
      20488: inst = 32'h10408000;
      20489: inst = 32'hc40503c;
      20490: inst = 32'h8220000;
      20491: inst = 32'h10408000;
      20492: inst = 32'hc40503d;
      20493: inst = 32'h8220000;
      20494: inst = 32'h10408000;
      20495: inst = 32'hc405049;
      20496: inst = 32'h8220000;
      20497: inst = 32'h10408000;
      20498: inst = 32'hc40504a;
      20499: inst = 32'h8220000;
      20500: inst = 32'h10408000;
      20501: inst = 32'hc40506b;
      20502: inst = 32'h8220000;
      20503: inst = 32'h10408000;
      20504: inst = 32'hc40506c;
      20505: inst = 32'h8220000;
      20506: inst = 32'h10408000;
      20507: inst = 32'hc40506d;
      20508: inst = 32'h8220000;
      20509: inst = 32'h10408000;
      20510: inst = 32'hc40506e;
      20511: inst = 32'h8220000;
      20512: inst = 32'h10408000;
      20513: inst = 32'hc40506f;
      20514: inst = 32'h8220000;
      20515: inst = 32'h10408000;
      20516: inst = 32'hc405070;
      20517: inst = 32'h8220000;
      20518: inst = 32'h10408000;
      20519: inst = 32'hc405071;
      20520: inst = 32'h8220000;
      20521: inst = 32'h10408000;
      20522: inst = 32'hc405072;
      20523: inst = 32'h8220000;
      20524: inst = 32'h10408000;
      20525: inst = 32'hc405073;
      20526: inst = 32'h8220000;
      20527: inst = 32'h10408000;
      20528: inst = 32'hc405074;
      20529: inst = 32'h8220000;
      20530: inst = 32'h10408000;
      20531: inst = 32'hc405075;
      20532: inst = 32'h8220000;
      20533: inst = 32'h10408000;
      20534: inst = 32'hc405077;
      20535: inst = 32'h8220000;
      20536: inst = 32'h10408000;
      20537: inst = 32'hc405078;
      20538: inst = 32'h8220000;
      20539: inst = 32'h10408000;
      20540: inst = 32'hc405079;
      20541: inst = 32'h8220000;
      20542: inst = 32'h10408000;
      20543: inst = 32'hc40507a;
      20544: inst = 32'h8220000;
      20545: inst = 32'h10408000;
      20546: inst = 32'hc40507b;
      20547: inst = 32'h8220000;
      20548: inst = 32'h10408000;
      20549: inst = 32'hc40507c;
      20550: inst = 32'h8220000;
      20551: inst = 32'h10408000;
      20552: inst = 32'hc40507d;
      20553: inst = 32'h8220000;
      20554: inst = 32'h10408000;
      20555: inst = 32'hc40507e;
      20556: inst = 32'h8220000;
      20557: inst = 32'h10408000;
      20558: inst = 32'hc40507f;
      20559: inst = 32'h8220000;
      20560: inst = 32'h10408000;
      20561: inst = 32'hc405080;
      20562: inst = 32'h8220000;
      20563: inst = 32'h10408000;
      20564: inst = 32'hc405084;
      20565: inst = 32'h8220000;
      20566: inst = 32'h10408000;
      20567: inst = 32'hc405085;
      20568: inst = 32'h8220000;
      20569: inst = 32'h10408000;
      20570: inst = 32'hc405086;
      20571: inst = 32'h8220000;
      20572: inst = 32'h10408000;
      20573: inst = 32'hc405087;
      20574: inst = 32'h8220000;
      20575: inst = 32'h10408000;
      20576: inst = 32'hc405088;
      20577: inst = 32'h8220000;
      20578: inst = 32'h10408000;
      20579: inst = 32'hc405089;
      20580: inst = 32'h8220000;
      20581: inst = 32'h10408000;
      20582: inst = 32'hc40508a;
      20583: inst = 32'h8220000;
      20584: inst = 32'h10408000;
      20585: inst = 32'hc40508b;
      20586: inst = 32'h8220000;
      20587: inst = 32'h10408000;
      20588: inst = 32'hc40508c;
      20589: inst = 32'h8220000;
      20590: inst = 32'h10408000;
      20591: inst = 32'hc40508d;
      20592: inst = 32'h8220000;
      20593: inst = 32'h10408000;
      20594: inst = 32'hc405090;
      20595: inst = 32'h8220000;
      20596: inst = 32'h10408000;
      20597: inst = 32'hc405091;
      20598: inst = 32'h8220000;
      20599: inst = 32'h10408000;
      20600: inst = 32'hc405096;
      20601: inst = 32'h8220000;
      20602: inst = 32'h10408000;
      20603: inst = 32'hc405097;
      20604: inst = 32'h8220000;
      20605: inst = 32'h10408000;
      20606: inst = 32'hc405098;
      20607: inst = 32'h8220000;
      20608: inst = 32'h10408000;
      20609: inst = 32'hc405099;
      20610: inst = 32'h8220000;
      20611: inst = 32'h10408000;
      20612: inst = 32'hc40509c;
      20613: inst = 32'h8220000;
      20614: inst = 32'h10408000;
      20615: inst = 32'hc40509d;
      20616: inst = 32'h8220000;
      20617: inst = 32'h10408000;
      20618: inst = 32'hc4050a9;
      20619: inst = 32'h8220000;
      20620: inst = 32'h10408000;
      20621: inst = 32'hc4050aa;
      20622: inst = 32'h8220000;
      20623: inst = 32'h10408000;
      20624: inst = 32'hc4050ab;
      20625: inst = 32'h8220000;
      20626: inst = 32'h10408000;
      20627: inst = 32'hc4050ac;
      20628: inst = 32'h8220000;
      20629: inst = 32'h10408000;
      20630: inst = 32'hc4050ad;
      20631: inst = 32'h8220000;
      20632: inst = 32'h10408000;
      20633: inst = 32'hc4050ae;
      20634: inst = 32'h8220000;
      20635: inst = 32'h10408000;
      20636: inst = 32'hc4050af;
      20637: inst = 32'h8220000;
      20638: inst = 32'h10408000;
      20639: inst = 32'hc4050b0;
      20640: inst = 32'h8220000;
      20641: inst = 32'h10408000;
      20642: inst = 32'hc4050b1;
      20643: inst = 32'h8220000;
      20644: inst = 32'h10408000;
      20645: inst = 32'hc4050b2;
      20646: inst = 32'h8220000;
      20647: inst = 32'h10408000;
      20648: inst = 32'hc4050b3;
      20649: inst = 32'h8220000;
      20650: inst = 32'h10408000;
      20651: inst = 32'hc4050cb;
      20652: inst = 32'h8220000;
      20653: inst = 32'h10408000;
      20654: inst = 32'hc4050cc;
      20655: inst = 32'h8220000;
      20656: inst = 32'h10408000;
      20657: inst = 32'hc4050cd;
      20658: inst = 32'h8220000;
      20659: inst = 32'h10408000;
      20660: inst = 32'hc4050ce;
      20661: inst = 32'h8220000;
      20662: inst = 32'h10408000;
      20663: inst = 32'hc4050cf;
      20664: inst = 32'h8220000;
      20665: inst = 32'h10408000;
      20666: inst = 32'hc4050d0;
      20667: inst = 32'h8220000;
      20668: inst = 32'h10408000;
      20669: inst = 32'hc4050d1;
      20670: inst = 32'h8220000;
      20671: inst = 32'h10408000;
      20672: inst = 32'hc4050d2;
      20673: inst = 32'h8220000;
      20674: inst = 32'h10408000;
      20675: inst = 32'hc4050d3;
      20676: inst = 32'h8220000;
      20677: inst = 32'h10408000;
      20678: inst = 32'hc4050d4;
      20679: inst = 32'h8220000;
      20680: inst = 32'h10408000;
      20681: inst = 32'hc4050d7;
      20682: inst = 32'h8220000;
      20683: inst = 32'h10408000;
      20684: inst = 32'hc4050d8;
      20685: inst = 32'h8220000;
      20686: inst = 32'h10408000;
      20687: inst = 32'hc4050d9;
      20688: inst = 32'h8220000;
      20689: inst = 32'h10408000;
      20690: inst = 32'hc4050da;
      20691: inst = 32'h8220000;
      20692: inst = 32'h10408000;
      20693: inst = 32'hc4050db;
      20694: inst = 32'h8220000;
      20695: inst = 32'h10408000;
      20696: inst = 32'hc4050dc;
      20697: inst = 32'h8220000;
      20698: inst = 32'h10408000;
      20699: inst = 32'hc4050dd;
      20700: inst = 32'h8220000;
      20701: inst = 32'h10408000;
      20702: inst = 32'hc4050de;
      20703: inst = 32'h8220000;
      20704: inst = 32'h10408000;
      20705: inst = 32'hc4050df;
      20706: inst = 32'h8220000;
      20707: inst = 32'h10408000;
      20708: inst = 32'hc4050e0;
      20709: inst = 32'h8220000;
      20710: inst = 32'h10408000;
      20711: inst = 32'hc4050e1;
      20712: inst = 32'h8220000;
      20713: inst = 32'h10408000;
      20714: inst = 32'hc4050e5;
      20715: inst = 32'h8220000;
      20716: inst = 32'h10408000;
      20717: inst = 32'hc4050e6;
      20718: inst = 32'h8220000;
      20719: inst = 32'h10408000;
      20720: inst = 32'hc4050e7;
      20721: inst = 32'h8220000;
      20722: inst = 32'h10408000;
      20723: inst = 32'hc4050e8;
      20724: inst = 32'h8220000;
      20725: inst = 32'h10408000;
      20726: inst = 32'hc4050e9;
      20727: inst = 32'h8220000;
      20728: inst = 32'h10408000;
      20729: inst = 32'hc4050ea;
      20730: inst = 32'h8220000;
      20731: inst = 32'h10408000;
      20732: inst = 32'hc4050eb;
      20733: inst = 32'h8220000;
      20734: inst = 32'h10408000;
      20735: inst = 32'hc4050ec;
      20736: inst = 32'h8220000;
      20737: inst = 32'h10408000;
      20738: inst = 32'hc4050ed;
      20739: inst = 32'h8220000;
      20740: inst = 32'h10408000;
      20741: inst = 32'hc4050f0;
      20742: inst = 32'h8220000;
      20743: inst = 32'h10408000;
      20744: inst = 32'hc4050f1;
      20745: inst = 32'h8220000;
      20746: inst = 32'h10408000;
      20747: inst = 32'hc4050f6;
      20748: inst = 32'h8220000;
      20749: inst = 32'h10408000;
      20750: inst = 32'hc4050f7;
      20751: inst = 32'h8220000;
      20752: inst = 32'h10408000;
      20753: inst = 32'hc4050f8;
      20754: inst = 32'h8220000;
      20755: inst = 32'h10408000;
      20756: inst = 32'hc4050f9;
      20757: inst = 32'h8220000;
      20758: inst = 32'h10408000;
      20759: inst = 32'hc4050fa;
      20760: inst = 32'h8220000;
      20761: inst = 32'h10408000;
      20762: inst = 32'hc4050fc;
      20763: inst = 32'h8220000;
      20764: inst = 32'h10408000;
      20765: inst = 32'hc4050fd;
      20766: inst = 32'h8220000;
      20767: inst = 32'h10408000;
      20768: inst = 32'hc405109;
      20769: inst = 32'h8220000;
      20770: inst = 32'h10408000;
      20771: inst = 32'hc40510a;
      20772: inst = 32'h8220000;
      20773: inst = 32'h10408000;
      20774: inst = 32'hc40510b;
      20775: inst = 32'h8220000;
      20776: inst = 32'h10408000;
      20777: inst = 32'hc40510c;
      20778: inst = 32'h8220000;
      20779: inst = 32'h10408000;
      20780: inst = 32'hc40510d;
      20781: inst = 32'h8220000;
      20782: inst = 32'h10408000;
      20783: inst = 32'hc40510e;
      20784: inst = 32'h8220000;
      20785: inst = 32'h10408000;
      20786: inst = 32'hc40510f;
      20787: inst = 32'h8220000;
      20788: inst = 32'h10408000;
      20789: inst = 32'hc405110;
      20790: inst = 32'h8220000;
      20791: inst = 32'h10408000;
      20792: inst = 32'hc405111;
      20793: inst = 32'h8220000;
      20794: inst = 32'h10408000;
      20795: inst = 32'hc405112;
      20796: inst = 32'h8220000;
      20797: inst = 32'h10408000;
      20798: inst = 32'hc405113;
      20799: inst = 32'h8220000;
      20800: inst = 32'h58000000;
      20801: inst = 32'h29c20000;
      20802: inst = 32'h29e30000;
      20803: inst = 32'h11600000;
      20804: inst = 32'hd600060;
      20805: inst = 32'h12208000;
      20806: inst = 32'he203fe0;
      20807: inst = 32'h13e00000;
      20808: inst = 32'hfe0515f;
      20809: inst = 32'h20200000;
      20810: inst = 32'h5be00000;
      20811: inst = 32'h13e00000;
      20812: inst = 32'hfe05d2e;
      20813: inst = 32'h20200001;
      20814: inst = 32'h5be00000;
      20815: inst = 32'h13e00000;
      20816: inst = 32'hfe05d2e;
      20817: inst = 32'h20200002;
      20818: inst = 32'h5be00000;
      20819: inst = 32'h13e00000;
      20820: inst = 32'hfe05954;
      20821: inst = 32'h20200003;
      20822: inst = 32'h5be00000;
      20823: inst = 32'h13e00000;
      20824: inst = 32'hfe05954;
      20825: inst = 32'h20200004;
      20826: inst = 32'h5be00000;
      20827: inst = 32'h13e00000;
      20828: inst = 32'hfe05564;
      20829: inst = 32'h20200005;
      20830: inst = 32'h5be00000;
      20831: inst = 32'hc6018c3;
      20832: inst = 32'h2a0e0000;
      20833: inst = 32'h294f0000;
      20834: inst = 32'h11200000;
      20835: inst = 32'hd205167;
      20836: inst = 32'h13e00000;
      20837: inst = 32'hfe0a9fb;
      20838: inst = 32'h5be00000;
      20839: inst = 32'h244c8000;
      20840: inst = 32'h24428800;
      20841: inst = 32'h8620000;
      20842: inst = 32'h2a0e0001;
      20843: inst = 32'h294f0000;
      20844: inst = 32'h11200000;
      20845: inst = 32'hd205171;
      20846: inst = 32'h13e00000;
      20847: inst = 32'hfe0a9fb;
      20848: inst = 32'h5be00000;
      20849: inst = 32'h244c8000;
      20850: inst = 32'h24428800;
      20851: inst = 32'h8620000;
      20852: inst = 32'h2a0e0002;
      20853: inst = 32'h294f0000;
      20854: inst = 32'h11200000;
      20855: inst = 32'hd20517b;
      20856: inst = 32'h13e00000;
      20857: inst = 32'hfe0a9fb;
      20858: inst = 32'h5be00000;
      20859: inst = 32'h244c8000;
      20860: inst = 32'h24428800;
      20861: inst = 32'h8620000;
      20862: inst = 32'h2a0e0003;
      20863: inst = 32'h294f0000;
      20864: inst = 32'h11200000;
      20865: inst = 32'hd205185;
      20866: inst = 32'h13e00000;
      20867: inst = 32'hfe0a9fb;
      20868: inst = 32'h5be00000;
      20869: inst = 32'h244c8000;
      20870: inst = 32'h24428800;
      20871: inst = 32'h8620000;
      20872: inst = 32'h2a0e0004;
      20873: inst = 32'h294f0000;
      20874: inst = 32'h11200000;
      20875: inst = 32'hd20518f;
      20876: inst = 32'h13e00000;
      20877: inst = 32'hfe0a9fb;
      20878: inst = 32'h5be00000;
      20879: inst = 32'h244c8000;
      20880: inst = 32'h24428800;
      20881: inst = 32'h8620000;
      20882: inst = 32'h2a0e0005;
      20883: inst = 32'h294f0000;
      20884: inst = 32'h11200000;
      20885: inst = 32'hd205199;
      20886: inst = 32'h13e00000;
      20887: inst = 32'hfe0a9fb;
      20888: inst = 32'h5be00000;
      20889: inst = 32'h244c8000;
      20890: inst = 32'h24428800;
      20891: inst = 32'h8620000;
      20892: inst = 32'h2a0e0006;
      20893: inst = 32'h294f0000;
      20894: inst = 32'h11200000;
      20895: inst = 32'hd2051a3;
      20896: inst = 32'h13e00000;
      20897: inst = 32'hfe0a9fb;
      20898: inst = 32'h5be00000;
      20899: inst = 32'h244c8000;
      20900: inst = 32'h24428800;
      20901: inst = 32'h8620000;
      20902: inst = 32'h2a0e0007;
      20903: inst = 32'h294f0000;
      20904: inst = 32'h11200000;
      20905: inst = 32'hd2051ad;
      20906: inst = 32'h13e00000;
      20907: inst = 32'hfe0a9fb;
      20908: inst = 32'h5be00000;
      20909: inst = 32'h244c8000;
      20910: inst = 32'h24428800;
      20911: inst = 32'h8620000;
      20912: inst = 32'h2a0e0008;
      20913: inst = 32'h294f0000;
      20914: inst = 32'h11200000;
      20915: inst = 32'hd2051b7;
      20916: inst = 32'h13e00000;
      20917: inst = 32'hfe0a9fb;
      20918: inst = 32'h5be00000;
      20919: inst = 32'h244c8000;
      20920: inst = 32'h24428800;
      20921: inst = 32'h8620000;
      20922: inst = 32'h2a0e0009;
      20923: inst = 32'h294f0000;
      20924: inst = 32'h11200000;
      20925: inst = 32'hd2051c1;
      20926: inst = 32'h13e00000;
      20927: inst = 32'hfe0a9fb;
      20928: inst = 32'h5be00000;
      20929: inst = 32'h244c8000;
      20930: inst = 32'h24428800;
      20931: inst = 32'h8620000;
      20932: inst = 32'h2a0e0000;
      20933: inst = 32'h294f0001;
      20934: inst = 32'h11200000;
      20935: inst = 32'hd2051cb;
      20936: inst = 32'h13e00000;
      20937: inst = 32'hfe0a9fb;
      20938: inst = 32'h5be00000;
      20939: inst = 32'h244c8000;
      20940: inst = 32'h24428800;
      20941: inst = 32'h8620000;
      20942: inst = 32'h2a0e0001;
      20943: inst = 32'h294f0001;
      20944: inst = 32'h11200000;
      20945: inst = 32'hd2051d5;
      20946: inst = 32'h13e00000;
      20947: inst = 32'hfe0a9fb;
      20948: inst = 32'h5be00000;
      20949: inst = 32'h244c8000;
      20950: inst = 32'h24428800;
      20951: inst = 32'h8620000;
      20952: inst = 32'h2a0e0002;
      20953: inst = 32'h294f0001;
      20954: inst = 32'h11200000;
      20955: inst = 32'hd2051df;
      20956: inst = 32'h13e00000;
      20957: inst = 32'hfe0a9fb;
      20958: inst = 32'h5be00000;
      20959: inst = 32'h244c8000;
      20960: inst = 32'h24428800;
      20961: inst = 32'h8620000;
      20962: inst = 32'h2a0e0003;
      20963: inst = 32'h294f0001;
      20964: inst = 32'h11200000;
      20965: inst = 32'hd2051e9;
      20966: inst = 32'h13e00000;
      20967: inst = 32'hfe0a9fb;
      20968: inst = 32'h5be00000;
      20969: inst = 32'h244c8000;
      20970: inst = 32'h24428800;
      20971: inst = 32'h8620000;
      20972: inst = 32'h2a0e0004;
      20973: inst = 32'h294f0001;
      20974: inst = 32'h11200000;
      20975: inst = 32'hd2051f3;
      20976: inst = 32'h13e00000;
      20977: inst = 32'hfe0a9fb;
      20978: inst = 32'h5be00000;
      20979: inst = 32'h244c8000;
      20980: inst = 32'h24428800;
      20981: inst = 32'h8620000;
      20982: inst = 32'h2a0e0005;
      20983: inst = 32'h294f0001;
      20984: inst = 32'h11200000;
      20985: inst = 32'hd2051fd;
      20986: inst = 32'h13e00000;
      20987: inst = 32'hfe0a9fb;
      20988: inst = 32'h5be00000;
      20989: inst = 32'h244c8000;
      20990: inst = 32'h24428800;
      20991: inst = 32'h8620000;
      20992: inst = 32'h2a0e0006;
      20993: inst = 32'h294f0001;
      20994: inst = 32'h11200000;
      20995: inst = 32'hd205207;
      20996: inst = 32'h13e00000;
      20997: inst = 32'hfe0a9fb;
      20998: inst = 32'h5be00000;
      20999: inst = 32'h244c8000;
      21000: inst = 32'h24428800;
      21001: inst = 32'h8620000;
      21002: inst = 32'h2a0e0007;
      21003: inst = 32'h294f0001;
      21004: inst = 32'h11200000;
      21005: inst = 32'hd205211;
      21006: inst = 32'h13e00000;
      21007: inst = 32'hfe0a9fb;
      21008: inst = 32'h5be00000;
      21009: inst = 32'h244c8000;
      21010: inst = 32'h24428800;
      21011: inst = 32'h8620000;
      21012: inst = 32'h2a0e0008;
      21013: inst = 32'h294f0001;
      21014: inst = 32'h11200000;
      21015: inst = 32'hd20521b;
      21016: inst = 32'h13e00000;
      21017: inst = 32'hfe0a9fb;
      21018: inst = 32'h5be00000;
      21019: inst = 32'h244c8000;
      21020: inst = 32'h24428800;
      21021: inst = 32'h8620000;
      21022: inst = 32'h2a0e0009;
      21023: inst = 32'h294f0001;
      21024: inst = 32'h11200000;
      21025: inst = 32'hd205225;
      21026: inst = 32'h13e00000;
      21027: inst = 32'hfe0a9fb;
      21028: inst = 32'h5be00000;
      21029: inst = 32'h244c8000;
      21030: inst = 32'h24428800;
      21031: inst = 32'h8620000;
      21032: inst = 32'h2a0e0000;
      21033: inst = 32'h294f0002;
      21034: inst = 32'h11200000;
      21035: inst = 32'hd20522f;
      21036: inst = 32'h13e00000;
      21037: inst = 32'hfe0a9fb;
      21038: inst = 32'h5be00000;
      21039: inst = 32'h244c8000;
      21040: inst = 32'h24428800;
      21041: inst = 32'h8620000;
      21042: inst = 32'h2a0e0009;
      21043: inst = 32'h294f0002;
      21044: inst = 32'h11200000;
      21045: inst = 32'hd205239;
      21046: inst = 32'h13e00000;
      21047: inst = 32'hfe0a9fb;
      21048: inst = 32'h5be00000;
      21049: inst = 32'h244c8000;
      21050: inst = 32'h24428800;
      21051: inst = 32'h8620000;
      21052: inst = 32'h2a0e0000;
      21053: inst = 32'h294f0003;
      21054: inst = 32'h11200000;
      21055: inst = 32'hd205243;
      21056: inst = 32'h13e00000;
      21057: inst = 32'hfe0a9fb;
      21058: inst = 32'h5be00000;
      21059: inst = 32'h244c8000;
      21060: inst = 32'h24428800;
      21061: inst = 32'h8620000;
      21062: inst = 32'h2a0e0002;
      21063: inst = 32'h294f0003;
      21064: inst = 32'h11200000;
      21065: inst = 32'hd20524d;
      21066: inst = 32'h13e00000;
      21067: inst = 32'hfe0a9fb;
      21068: inst = 32'h5be00000;
      21069: inst = 32'h244c8000;
      21070: inst = 32'h24428800;
      21071: inst = 32'h8620000;
      21072: inst = 32'h2a0e0007;
      21073: inst = 32'h294f0003;
      21074: inst = 32'h11200000;
      21075: inst = 32'hd205257;
      21076: inst = 32'h13e00000;
      21077: inst = 32'hfe0a9fb;
      21078: inst = 32'h5be00000;
      21079: inst = 32'h244c8000;
      21080: inst = 32'h24428800;
      21081: inst = 32'h8620000;
      21082: inst = 32'h2a0e0009;
      21083: inst = 32'h294f0003;
      21084: inst = 32'h11200000;
      21085: inst = 32'hd205261;
      21086: inst = 32'h13e00000;
      21087: inst = 32'hfe0a9fb;
      21088: inst = 32'h5be00000;
      21089: inst = 32'h244c8000;
      21090: inst = 32'h24428800;
      21091: inst = 32'h8620000;
      21092: inst = 32'h2a0e0000;
      21093: inst = 32'h294f0004;
      21094: inst = 32'h11200000;
      21095: inst = 32'hd20526b;
      21096: inst = 32'h13e00000;
      21097: inst = 32'hfe0a9fb;
      21098: inst = 32'h5be00000;
      21099: inst = 32'h244c8000;
      21100: inst = 32'h24428800;
      21101: inst = 32'h8620000;
      21102: inst = 32'h2a0e0002;
      21103: inst = 32'h294f0004;
      21104: inst = 32'h11200000;
      21105: inst = 32'hd205275;
      21106: inst = 32'h13e00000;
      21107: inst = 32'hfe0a9fb;
      21108: inst = 32'h5be00000;
      21109: inst = 32'h244c8000;
      21110: inst = 32'h24428800;
      21111: inst = 32'h8620000;
      21112: inst = 32'h2a0e0007;
      21113: inst = 32'h294f0004;
      21114: inst = 32'h11200000;
      21115: inst = 32'hd20527f;
      21116: inst = 32'h13e00000;
      21117: inst = 32'hfe0a9fb;
      21118: inst = 32'h5be00000;
      21119: inst = 32'h244c8000;
      21120: inst = 32'h24428800;
      21121: inst = 32'h8620000;
      21122: inst = 32'h2a0e0009;
      21123: inst = 32'h294f0004;
      21124: inst = 32'h11200000;
      21125: inst = 32'hd205289;
      21126: inst = 32'h13e00000;
      21127: inst = 32'hfe0a9fb;
      21128: inst = 32'h5be00000;
      21129: inst = 32'h244c8000;
      21130: inst = 32'h24428800;
      21131: inst = 32'h8620000;
      21132: inst = 32'h2a0e0000;
      21133: inst = 32'h294f0005;
      21134: inst = 32'h11200000;
      21135: inst = 32'hd205293;
      21136: inst = 32'h13e00000;
      21137: inst = 32'hfe0a9fb;
      21138: inst = 32'h5be00000;
      21139: inst = 32'h244c8000;
      21140: inst = 32'h24428800;
      21141: inst = 32'h8620000;
      21142: inst = 32'h2a0e0009;
      21143: inst = 32'h294f0005;
      21144: inst = 32'h11200000;
      21145: inst = 32'hd20529d;
      21146: inst = 32'h13e00000;
      21147: inst = 32'hfe0a9fb;
      21148: inst = 32'h5be00000;
      21149: inst = 32'h244c8000;
      21150: inst = 32'h24428800;
      21151: inst = 32'h8620000;
      21152: inst = 32'h2a0e0000;
      21153: inst = 32'h294f0006;
      21154: inst = 32'h11200000;
      21155: inst = 32'hd2052a7;
      21156: inst = 32'h13e00000;
      21157: inst = 32'hfe0a9fb;
      21158: inst = 32'h5be00000;
      21159: inst = 32'h244c8000;
      21160: inst = 32'h24428800;
      21161: inst = 32'h8620000;
      21162: inst = 32'h2a0e0009;
      21163: inst = 32'h294f0006;
      21164: inst = 32'h11200000;
      21165: inst = 32'hd2052b1;
      21166: inst = 32'h13e00000;
      21167: inst = 32'hfe0a9fb;
      21168: inst = 32'h5be00000;
      21169: inst = 32'h244c8000;
      21170: inst = 32'h24428800;
      21171: inst = 32'h8620000;
      21172: inst = 32'hc60f4ce;
      21173: inst = 32'h2a0e0001;
      21174: inst = 32'h294f0002;
      21175: inst = 32'h11200000;
      21176: inst = 32'hd2052bc;
      21177: inst = 32'h13e00000;
      21178: inst = 32'hfe0a9fb;
      21179: inst = 32'h5be00000;
      21180: inst = 32'h244c8000;
      21181: inst = 32'h24428800;
      21182: inst = 32'h8620000;
      21183: inst = 32'h2a0e0002;
      21184: inst = 32'h294f0002;
      21185: inst = 32'h11200000;
      21186: inst = 32'hd2052c6;
      21187: inst = 32'h13e00000;
      21188: inst = 32'hfe0a9fb;
      21189: inst = 32'h5be00000;
      21190: inst = 32'h244c8000;
      21191: inst = 32'h24428800;
      21192: inst = 32'h8620000;
      21193: inst = 32'h2a0e0003;
      21194: inst = 32'h294f0002;
      21195: inst = 32'h11200000;
      21196: inst = 32'hd2052d0;
      21197: inst = 32'h13e00000;
      21198: inst = 32'hfe0a9fb;
      21199: inst = 32'h5be00000;
      21200: inst = 32'h244c8000;
      21201: inst = 32'h24428800;
      21202: inst = 32'h8620000;
      21203: inst = 32'h2a0e0004;
      21204: inst = 32'h294f0002;
      21205: inst = 32'h11200000;
      21206: inst = 32'hd2052da;
      21207: inst = 32'h13e00000;
      21208: inst = 32'hfe0a9fb;
      21209: inst = 32'h5be00000;
      21210: inst = 32'h244c8000;
      21211: inst = 32'h24428800;
      21212: inst = 32'h8620000;
      21213: inst = 32'h2a0e0005;
      21214: inst = 32'h294f0002;
      21215: inst = 32'h11200000;
      21216: inst = 32'hd2052e4;
      21217: inst = 32'h13e00000;
      21218: inst = 32'hfe0a9fb;
      21219: inst = 32'h5be00000;
      21220: inst = 32'h244c8000;
      21221: inst = 32'h24428800;
      21222: inst = 32'h8620000;
      21223: inst = 32'h2a0e0006;
      21224: inst = 32'h294f0002;
      21225: inst = 32'h11200000;
      21226: inst = 32'hd2052ee;
      21227: inst = 32'h13e00000;
      21228: inst = 32'hfe0a9fb;
      21229: inst = 32'h5be00000;
      21230: inst = 32'h244c8000;
      21231: inst = 32'h24428800;
      21232: inst = 32'h8620000;
      21233: inst = 32'h2a0e0007;
      21234: inst = 32'h294f0002;
      21235: inst = 32'h11200000;
      21236: inst = 32'hd2052f8;
      21237: inst = 32'h13e00000;
      21238: inst = 32'hfe0a9fb;
      21239: inst = 32'h5be00000;
      21240: inst = 32'h244c8000;
      21241: inst = 32'h24428800;
      21242: inst = 32'h8620000;
      21243: inst = 32'h2a0e0008;
      21244: inst = 32'h294f0002;
      21245: inst = 32'h11200000;
      21246: inst = 32'hd205302;
      21247: inst = 32'h13e00000;
      21248: inst = 32'hfe0a9fb;
      21249: inst = 32'h5be00000;
      21250: inst = 32'h244c8000;
      21251: inst = 32'h24428800;
      21252: inst = 32'h8620000;
      21253: inst = 32'h2a0e0001;
      21254: inst = 32'h294f0003;
      21255: inst = 32'h11200000;
      21256: inst = 32'hd20530c;
      21257: inst = 32'h13e00000;
      21258: inst = 32'hfe0a9fb;
      21259: inst = 32'h5be00000;
      21260: inst = 32'h244c8000;
      21261: inst = 32'h24428800;
      21262: inst = 32'h8620000;
      21263: inst = 32'h2a0e0003;
      21264: inst = 32'h294f0003;
      21265: inst = 32'h11200000;
      21266: inst = 32'hd205316;
      21267: inst = 32'h13e00000;
      21268: inst = 32'hfe0a9fb;
      21269: inst = 32'h5be00000;
      21270: inst = 32'h244c8000;
      21271: inst = 32'h24428800;
      21272: inst = 32'h8620000;
      21273: inst = 32'h2a0e0004;
      21274: inst = 32'h294f0003;
      21275: inst = 32'h11200000;
      21276: inst = 32'hd205320;
      21277: inst = 32'h13e00000;
      21278: inst = 32'hfe0a9fb;
      21279: inst = 32'h5be00000;
      21280: inst = 32'h244c8000;
      21281: inst = 32'h24428800;
      21282: inst = 32'h8620000;
      21283: inst = 32'h2a0e0005;
      21284: inst = 32'h294f0003;
      21285: inst = 32'h11200000;
      21286: inst = 32'hd20532a;
      21287: inst = 32'h13e00000;
      21288: inst = 32'hfe0a9fb;
      21289: inst = 32'h5be00000;
      21290: inst = 32'h244c8000;
      21291: inst = 32'h24428800;
      21292: inst = 32'h8620000;
      21293: inst = 32'h2a0e0006;
      21294: inst = 32'h294f0003;
      21295: inst = 32'h11200000;
      21296: inst = 32'hd205334;
      21297: inst = 32'h13e00000;
      21298: inst = 32'hfe0a9fb;
      21299: inst = 32'h5be00000;
      21300: inst = 32'h244c8000;
      21301: inst = 32'h24428800;
      21302: inst = 32'h8620000;
      21303: inst = 32'h2a0e0008;
      21304: inst = 32'h294f0003;
      21305: inst = 32'h11200000;
      21306: inst = 32'hd20533e;
      21307: inst = 32'h13e00000;
      21308: inst = 32'hfe0a9fb;
      21309: inst = 32'h5be00000;
      21310: inst = 32'h244c8000;
      21311: inst = 32'h24428800;
      21312: inst = 32'h8620000;
      21313: inst = 32'h2a0e0001;
      21314: inst = 32'h294f0004;
      21315: inst = 32'h11200000;
      21316: inst = 32'hd205348;
      21317: inst = 32'h13e00000;
      21318: inst = 32'hfe0a9fb;
      21319: inst = 32'h5be00000;
      21320: inst = 32'h244c8000;
      21321: inst = 32'h24428800;
      21322: inst = 32'h8620000;
      21323: inst = 32'h2a0e0003;
      21324: inst = 32'h294f0004;
      21325: inst = 32'h11200000;
      21326: inst = 32'hd205352;
      21327: inst = 32'h13e00000;
      21328: inst = 32'hfe0a9fb;
      21329: inst = 32'h5be00000;
      21330: inst = 32'h244c8000;
      21331: inst = 32'h24428800;
      21332: inst = 32'h8620000;
      21333: inst = 32'h2a0e0004;
      21334: inst = 32'h294f0004;
      21335: inst = 32'h11200000;
      21336: inst = 32'hd20535c;
      21337: inst = 32'h13e00000;
      21338: inst = 32'hfe0a9fb;
      21339: inst = 32'h5be00000;
      21340: inst = 32'h244c8000;
      21341: inst = 32'h24428800;
      21342: inst = 32'h8620000;
      21343: inst = 32'h2a0e0005;
      21344: inst = 32'h294f0004;
      21345: inst = 32'h11200000;
      21346: inst = 32'hd205366;
      21347: inst = 32'h13e00000;
      21348: inst = 32'hfe0a9fb;
      21349: inst = 32'h5be00000;
      21350: inst = 32'h244c8000;
      21351: inst = 32'h24428800;
      21352: inst = 32'h8620000;
      21353: inst = 32'h2a0e0006;
      21354: inst = 32'h294f0004;
      21355: inst = 32'h11200000;
      21356: inst = 32'hd205370;
      21357: inst = 32'h13e00000;
      21358: inst = 32'hfe0a9fb;
      21359: inst = 32'h5be00000;
      21360: inst = 32'h244c8000;
      21361: inst = 32'h24428800;
      21362: inst = 32'h8620000;
      21363: inst = 32'h2a0e0008;
      21364: inst = 32'h294f0004;
      21365: inst = 32'h11200000;
      21366: inst = 32'hd20537a;
      21367: inst = 32'h13e00000;
      21368: inst = 32'hfe0a9fb;
      21369: inst = 32'h5be00000;
      21370: inst = 32'h244c8000;
      21371: inst = 32'h24428800;
      21372: inst = 32'h8620000;
      21373: inst = 32'h2a0e0001;
      21374: inst = 32'h294f0005;
      21375: inst = 32'h11200000;
      21376: inst = 32'hd205384;
      21377: inst = 32'h13e00000;
      21378: inst = 32'hfe0a9fb;
      21379: inst = 32'h5be00000;
      21380: inst = 32'h244c8000;
      21381: inst = 32'h24428800;
      21382: inst = 32'h8620000;
      21383: inst = 32'h2a0e0002;
      21384: inst = 32'h294f0005;
      21385: inst = 32'h11200000;
      21386: inst = 32'hd20538e;
      21387: inst = 32'h13e00000;
      21388: inst = 32'hfe0a9fb;
      21389: inst = 32'h5be00000;
      21390: inst = 32'h244c8000;
      21391: inst = 32'h24428800;
      21392: inst = 32'h8620000;
      21393: inst = 32'h2a0e0003;
      21394: inst = 32'h294f0005;
      21395: inst = 32'h11200000;
      21396: inst = 32'hd205398;
      21397: inst = 32'h13e00000;
      21398: inst = 32'hfe0a9fb;
      21399: inst = 32'h5be00000;
      21400: inst = 32'h244c8000;
      21401: inst = 32'h24428800;
      21402: inst = 32'h8620000;
      21403: inst = 32'h2a0e0004;
      21404: inst = 32'h294f0005;
      21405: inst = 32'h11200000;
      21406: inst = 32'hd2053a2;
      21407: inst = 32'h13e00000;
      21408: inst = 32'hfe0a9fb;
      21409: inst = 32'h5be00000;
      21410: inst = 32'h244c8000;
      21411: inst = 32'h24428800;
      21412: inst = 32'h8620000;
      21413: inst = 32'h2a0e0005;
      21414: inst = 32'h294f0005;
      21415: inst = 32'h11200000;
      21416: inst = 32'hd2053ac;
      21417: inst = 32'h13e00000;
      21418: inst = 32'hfe0a9fb;
      21419: inst = 32'h5be00000;
      21420: inst = 32'h244c8000;
      21421: inst = 32'h24428800;
      21422: inst = 32'h8620000;
      21423: inst = 32'h2a0e0006;
      21424: inst = 32'h294f0005;
      21425: inst = 32'h11200000;
      21426: inst = 32'hd2053b6;
      21427: inst = 32'h13e00000;
      21428: inst = 32'hfe0a9fb;
      21429: inst = 32'h5be00000;
      21430: inst = 32'h244c8000;
      21431: inst = 32'h24428800;
      21432: inst = 32'h8620000;
      21433: inst = 32'h2a0e0007;
      21434: inst = 32'h294f0005;
      21435: inst = 32'h11200000;
      21436: inst = 32'hd2053c0;
      21437: inst = 32'h13e00000;
      21438: inst = 32'hfe0a9fb;
      21439: inst = 32'h5be00000;
      21440: inst = 32'h244c8000;
      21441: inst = 32'h24428800;
      21442: inst = 32'h8620000;
      21443: inst = 32'h2a0e0008;
      21444: inst = 32'h294f0005;
      21445: inst = 32'h11200000;
      21446: inst = 32'hd2053ca;
      21447: inst = 32'h13e00000;
      21448: inst = 32'hfe0a9fb;
      21449: inst = 32'h5be00000;
      21450: inst = 32'h244c8000;
      21451: inst = 32'h24428800;
      21452: inst = 32'h8620000;
      21453: inst = 32'h2a0e0001;
      21454: inst = 32'h294f0006;
      21455: inst = 32'h11200000;
      21456: inst = 32'hd2053d4;
      21457: inst = 32'h13e00000;
      21458: inst = 32'hfe0a9fb;
      21459: inst = 32'h5be00000;
      21460: inst = 32'h244c8000;
      21461: inst = 32'h24428800;
      21462: inst = 32'h8620000;
      21463: inst = 32'h2a0e0002;
      21464: inst = 32'h294f0006;
      21465: inst = 32'h11200000;
      21466: inst = 32'hd2053de;
      21467: inst = 32'h13e00000;
      21468: inst = 32'hfe0a9fb;
      21469: inst = 32'h5be00000;
      21470: inst = 32'h244c8000;
      21471: inst = 32'h24428800;
      21472: inst = 32'h8620000;
      21473: inst = 32'h2a0e0003;
      21474: inst = 32'h294f0006;
      21475: inst = 32'h11200000;
      21476: inst = 32'hd2053e8;
      21477: inst = 32'h13e00000;
      21478: inst = 32'hfe0a9fb;
      21479: inst = 32'h5be00000;
      21480: inst = 32'h244c8000;
      21481: inst = 32'h24428800;
      21482: inst = 32'h8620000;
      21483: inst = 32'h2a0e0004;
      21484: inst = 32'h294f0006;
      21485: inst = 32'h11200000;
      21486: inst = 32'hd2053f2;
      21487: inst = 32'h13e00000;
      21488: inst = 32'hfe0a9fb;
      21489: inst = 32'h5be00000;
      21490: inst = 32'h244c8000;
      21491: inst = 32'h24428800;
      21492: inst = 32'h8620000;
      21493: inst = 32'h2a0e0005;
      21494: inst = 32'h294f0006;
      21495: inst = 32'h11200000;
      21496: inst = 32'hd2053fc;
      21497: inst = 32'h13e00000;
      21498: inst = 32'hfe0a9fb;
      21499: inst = 32'h5be00000;
      21500: inst = 32'h244c8000;
      21501: inst = 32'h24428800;
      21502: inst = 32'h8620000;
      21503: inst = 32'h2a0e0006;
      21504: inst = 32'h294f0006;
      21505: inst = 32'h11200000;
      21506: inst = 32'hd205406;
      21507: inst = 32'h13e00000;
      21508: inst = 32'hfe0a9fb;
      21509: inst = 32'h5be00000;
      21510: inst = 32'h244c8000;
      21511: inst = 32'h24428800;
      21512: inst = 32'h8620000;
      21513: inst = 32'h2a0e0007;
      21514: inst = 32'h294f0006;
      21515: inst = 32'h11200000;
      21516: inst = 32'hd205410;
      21517: inst = 32'h13e00000;
      21518: inst = 32'hfe0a9fb;
      21519: inst = 32'h5be00000;
      21520: inst = 32'h244c8000;
      21521: inst = 32'h24428800;
      21522: inst = 32'h8620000;
      21523: inst = 32'h2a0e0008;
      21524: inst = 32'h294f0006;
      21525: inst = 32'h11200000;
      21526: inst = 32'hd20541a;
      21527: inst = 32'h13e00000;
      21528: inst = 32'hfe0a9fb;
      21529: inst = 32'h5be00000;
      21530: inst = 32'h244c8000;
      21531: inst = 32'h24428800;
      21532: inst = 32'h8620000;
      21533: inst = 32'h2a0e0000;
      21534: inst = 32'h294f0008;
      21535: inst = 32'h11200000;
      21536: inst = 32'hd205424;
      21537: inst = 32'h13e00000;
      21538: inst = 32'hfe0a9fb;
      21539: inst = 32'h5be00000;
      21540: inst = 32'h244c8000;
      21541: inst = 32'h24428800;
      21542: inst = 32'h8620000;
      21543: inst = 32'h2a0e0001;
      21544: inst = 32'h294f0008;
      21545: inst = 32'h11200000;
      21546: inst = 32'hd20542e;
      21547: inst = 32'h13e00000;
      21548: inst = 32'hfe0a9fb;
      21549: inst = 32'h5be00000;
      21550: inst = 32'h244c8000;
      21551: inst = 32'h24428800;
      21552: inst = 32'h8620000;
      21553: inst = 32'h2a0e0008;
      21554: inst = 32'h294f0008;
      21555: inst = 32'h11200000;
      21556: inst = 32'hd205438;
      21557: inst = 32'h13e00000;
      21558: inst = 32'hfe0a9fb;
      21559: inst = 32'h5be00000;
      21560: inst = 32'h244c8000;
      21561: inst = 32'h24428800;
      21562: inst = 32'h8620000;
      21563: inst = 32'h2a0e0009;
      21564: inst = 32'h294f0008;
      21565: inst = 32'h11200000;
      21566: inst = 32'hd205442;
      21567: inst = 32'h13e00000;
      21568: inst = 32'hfe0a9fb;
      21569: inst = 32'h5be00000;
      21570: inst = 32'h244c8000;
      21571: inst = 32'h24428800;
      21572: inst = 32'h8620000;
      21573: inst = 32'h2a0e0003;
      21574: inst = 32'h294f000c;
      21575: inst = 32'h11200000;
      21576: inst = 32'hd20544c;
      21577: inst = 32'h13e00000;
      21578: inst = 32'hfe0a9fb;
      21579: inst = 32'h5be00000;
      21580: inst = 32'h244c8000;
      21581: inst = 32'h24428800;
      21582: inst = 32'h8620000;
      21583: inst = 32'h2a0e0006;
      21584: inst = 32'h294f000c;
      21585: inst = 32'h11200000;
      21586: inst = 32'hd205456;
      21587: inst = 32'h13e00000;
      21588: inst = 32'hfe0a9fb;
      21589: inst = 32'h5be00000;
      21590: inst = 32'h244c8000;
      21591: inst = 32'h24428800;
      21592: inst = 32'h8620000;
      21593: inst = 32'hc607800;
      21594: inst = 32'h2a0e0002;
      21595: inst = 32'h294f0007;
      21596: inst = 32'h11200000;
      21597: inst = 32'hd205461;
      21598: inst = 32'h13e00000;
      21599: inst = 32'hfe0a9fb;
      21600: inst = 32'h5be00000;
      21601: inst = 32'h244c8000;
      21602: inst = 32'h24428800;
      21603: inst = 32'h8620000;
      21604: inst = 32'h2a0e0003;
      21605: inst = 32'h294f0007;
      21606: inst = 32'h11200000;
      21607: inst = 32'hd20546b;
      21608: inst = 32'h13e00000;
      21609: inst = 32'hfe0a9fb;
      21610: inst = 32'h5be00000;
      21611: inst = 32'h244c8000;
      21612: inst = 32'h24428800;
      21613: inst = 32'h8620000;
      21614: inst = 32'h2a0e0006;
      21615: inst = 32'h294f0007;
      21616: inst = 32'h11200000;
      21617: inst = 32'hd205475;
      21618: inst = 32'h13e00000;
      21619: inst = 32'hfe0a9fb;
      21620: inst = 32'h5be00000;
      21621: inst = 32'h244c8000;
      21622: inst = 32'h24428800;
      21623: inst = 32'h8620000;
      21624: inst = 32'h2a0e0007;
      21625: inst = 32'h294f0007;
      21626: inst = 32'h11200000;
      21627: inst = 32'hd20547f;
      21628: inst = 32'h13e00000;
      21629: inst = 32'hfe0a9fb;
      21630: inst = 32'h5be00000;
      21631: inst = 32'h244c8000;
      21632: inst = 32'h24428800;
      21633: inst = 32'h8620000;
      21634: inst = 32'hc60a000;
      21635: inst = 32'h2a0e0004;
      21636: inst = 32'h294f0007;
      21637: inst = 32'h11200000;
      21638: inst = 32'hd20548a;
      21639: inst = 32'h13e00000;
      21640: inst = 32'hfe0a9fb;
      21641: inst = 32'h5be00000;
      21642: inst = 32'h244c8000;
      21643: inst = 32'h24428800;
      21644: inst = 32'h8620000;
      21645: inst = 32'h2a0e0005;
      21646: inst = 32'h294f0007;
      21647: inst = 32'h11200000;
      21648: inst = 32'hd205494;
      21649: inst = 32'h13e00000;
      21650: inst = 32'hfe0a9fb;
      21651: inst = 32'h5be00000;
      21652: inst = 32'h244c8000;
      21653: inst = 32'h24428800;
      21654: inst = 32'h8620000;
      21655: inst = 32'h2a0e0002;
      21656: inst = 32'h294f0008;
      21657: inst = 32'h11200000;
      21658: inst = 32'hd20549e;
      21659: inst = 32'h13e00000;
      21660: inst = 32'hfe0a9fb;
      21661: inst = 32'h5be00000;
      21662: inst = 32'h244c8000;
      21663: inst = 32'h24428800;
      21664: inst = 32'h8620000;
      21665: inst = 32'h2a0e0003;
      21666: inst = 32'h294f0008;
      21667: inst = 32'h11200000;
      21668: inst = 32'hd2054a8;
      21669: inst = 32'h13e00000;
      21670: inst = 32'hfe0a9fb;
      21671: inst = 32'h5be00000;
      21672: inst = 32'h244c8000;
      21673: inst = 32'h24428800;
      21674: inst = 32'h8620000;
      21675: inst = 32'h2a0e0004;
      21676: inst = 32'h294f0008;
      21677: inst = 32'h11200000;
      21678: inst = 32'hd2054b2;
      21679: inst = 32'h13e00000;
      21680: inst = 32'hfe0a9fb;
      21681: inst = 32'h5be00000;
      21682: inst = 32'h244c8000;
      21683: inst = 32'h24428800;
      21684: inst = 32'h8620000;
      21685: inst = 32'h2a0e0005;
      21686: inst = 32'h294f0008;
      21687: inst = 32'h11200000;
      21688: inst = 32'hd2054bc;
      21689: inst = 32'h13e00000;
      21690: inst = 32'hfe0a9fb;
      21691: inst = 32'h5be00000;
      21692: inst = 32'h244c8000;
      21693: inst = 32'h24428800;
      21694: inst = 32'h8620000;
      21695: inst = 32'h2a0e0006;
      21696: inst = 32'h294f0008;
      21697: inst = 32'h11200000;
      21698: inst = 32'hd2054c6;
      21699: inst = 32'h13e00000;
      21700: inst = 32'hfe0a9fb;
      21701: inst = 32'h5be00000;
      21702: inst = 32'h244c8000;
      21703: inst = 32'h24428800;
      21704: inst = 32'h8620000;
      21705: inst = 32'h2a0e0007;
      21706: inst = 32'h294f0008;
      21707: inst = 32'h11200000;
      21708: inst = 32'hd2054d0;
      21709: inst = 32'h13e00000;
      21710: inst = 32'hfe0a9fb;
      21711: inst = 32'h5be00000;
      21712: inst = 32'h244c8000;
      21713: inst = 32'h24428800;
      21714: inst = 32'h8620000;
      21715: inst = 32'h2a0e0002;
      21716: inst = 32'h294f0009;
      21717: inst = 32'h11200000;
      21718: inst = 32'hd2054da;
      21719: inst = 32'h13e00000;
      21720: inst = 32'hfe0a9fb;
      21721: inst = 32'h5be00000;
      21722: inst = 32'h244c8000;
      21723: inst = 32'h24428800;
      21724: inst = 32'h8620000;
      21725: inst = 32'h2a0e0003;
      21726: inst = 32'h294f0009;
      21727: inst = 32'h11200000;
      21728: inst = 32'hd2054e4;
      21729: inst = 32'h13e00000;
      21730: inst = 32'hfe0a9fb;
      21731: inst = 32'h5be00000;
      21732: inst = 32'h244c8000;
      21733: inst = 32'h24428800;
      21734: inst = 32'h8620000;
      21735: inst = 32'h2a0e0004;
      21736: inst = 32'h294f0009;
      21737: inst = 32'h11200000;
      21738: inst = 32'hd2054ee;
      21739: inst = 32'h13e00000;
      21740: inst = 32'hfe0a9fb;
      21741: inst = 32'h5be00000;
      21742: inst = 32'h244c8000;
      21743: inst = 32'h24428800;
      21744: inst = 32'h8620000;
      21745: inst = 32'h2a0e0005;
      21746: inst = 32'h294f0009;
      21747: inst = 32'h11200000;
      21748: inst = 32'hd2054f8;
      21749: inst = 32'h13e00000;
      21750: inst = 32'hfe0a9fb;
      21751: inst = 32'h5be00000;
      21752: inst = 32'h244c8000;
      21753: inst = 32'h24428800;
      21754: inst = 32'h8620000;
      21755: inst = 32'h2a0e0006;
      21756: inst = 32'h294f0009;
      21757: inst = 32'h11200000;
      21758: inst = 32'hd205502;
      21759: inst = 32'h13e00000;
      21760: inst = 32'hfe0a9fb;
      21761: inst = 32'h5be00000;
      21762: inst = 32'h244c8000;
      21763: inst = 32'h24428800;
      21764: inst = 32'h8620000;
      21765: inst = 32'h2a0e0007;
      21766: inst = 32'h294f0009;
      21767: inst = 32'h11200000;
      21768: inst = 32'hd20550c;
      21769: inst = 32'h13e00000;
      21770: inst = 32'hfe0a9fb;
      21771: inst = 32'h5be00000;
      21772: inst = 32'h244c8000;
      21773: inst = 32'h24428800;
      21774: inst = 32'h8620000;
      21775: inst = 32'hc6010ac;
      21776: inst = 32'h2a0e0002;
      21777: inst = 32'h294f000a;
      21778: inst = 32'h11200000;
      21779: inst = 32'hd205517;
      21780: inst = 32'h13e00000;
      21781: inst = 32'hfe0a9fb;
      21782: inst = 32'h5be00000;
      21783: inst = 32'h244c8000;
      21784: inst = 32'h24428800;
      21785: inst = 32'h8620000;
      21786: inst = 32'h2a0e0003;
      21787: inst = 32'h294f000a;
      21788: inst = 32'h11200000;
      21789: inst = 32'hd205521;
      21790: inst = 32'h13e00000;
      21791: inst = 32'hfe0a9fb;
      21792: inst = 32'h5be00000;
      21793: inst = 32'h244c8000;
      21794: inst = 32'h24428800;
      21795: inst = 32'h8620000;
      21796: inst = 32'h2a0e0004;
      21797: inst = 32'h294f000a;
      21798: inst = 32'h11200000;
      21799: inst = 32'hd20552b;
      21800: inst = 32'h13e00000;
      21801: inst = 32'hfe0a9fb;
      21802: inst = 32'h5be00000;
      21803: inst = 32'h244c8000;
      21804: inst = 32'h24428800;
      21805: inst = 32'h8620000;
      21806: inst = 32'h2a0e0005;
      21807: inst = 32'h294f000a;
      21808: inst = 32'h11200000;
      21809: inst = 32'hd205535;
      21810: inst = 32'h13e00000;
      21811: inst = 32'hfe0a9fb;
      21812: inst = 32'h5be00000;
      21813: inst = 32'h244c8000;
      21814: inst = 32'h24428800;
      21815: inst = 32'h8620000;
      21816: inst = 32'h2a0e0006;
      21817: inst = 32'h294f000a;
      21818: inst = 32'h11200000;
      21819: inst = 32'hd20553f;
      21820: inst = 32'h13e00000;
      21821: inst = 32'hfe0a9fb;
      21822: inst = 32'h5be00000;
      21823: inst = 32'h244c8000;
      21824: inst = 32'h24428800;
      21825: inst = 32'h8620000;
      21826: inst = 32'h2a0e0007;
      21827: inst = 32'h294f000a;
      21828: inst = 32'h11200000;
      21829: inst = 32'hd205549;
      21830: inst = 32'h13e00000;
      21831: inst = 32'hfe0a9fb;
      21832: inst = 32'h5be00000;
      21833: inst = 32'h244c8000;
      21834: inst = 32'h24428800;
      21835: inst = 32'h8620000;
      21836: inst = 32'hc60d42c;
      21837: inst = 32'h2a0e0003;
      21838: inst = 32'h294f000b;
      21839: inst = 32'h11200000;
      21840: inst = 32'hd205554;
      21841: inst = 32'h13e00000;
      21842: inst = 32'hfe0a9fb;
      21843: inst = 32'h5be00000;
      21844: inst = 32'h244c8000;
      21845: inst = 32'h24428800;
      21846: inst = 32'h8620000;
      21847: inst = 32'h2a0e0006;
      21848: inst = 32'h294f000b;
      21849: inst = 32'h11200000;
      21850: inst = 32'hd20555e;
      21851: inst = 32'h13e00000;
      21852: inst = 32'hfe0a9fb;
      21853: inst = 32'h5be00000;
      21854: inst = 32'h244c8000;
      21855: inst = 32'h24428800;
      21856: inst = 32'h8620000;
      21857: inst = 32'h13e00000;
      21858: inst = 32'hfe06108;
      21859: inst = 32'h5be00000;
      21860: inst = 32'hc6018c3;
      21861: inst = 32'h2a0e0000;
      21862: inst = 32'h294f0000;
      21863: inst = 32'h11200000;
      21864: inst = 32'hd20556c;
      21865: inst = 32'h13e00000;
      21866: inst = 32'hfe0a9fb;
      21867: inst = 32'h5be00000;
      21868: inst = 32'h244c8000;
      21869: inst = 32'h24428800;
      21870: inst = 32'h8620000;
      21871: inst = 32'h2a0e0001;
      21872: inst = 32'h294f0000;
      21873: inst = 32'h11200000;
      21874: inst = 32'hd205576;
      21875: inst = 32'h13e00000;
      21876: inst = 32'hfe0a9fb;
      21877: inst = 32'h5be00000;
      21878: inst = 32'h244c8000;
      21879: inst = 32'h24428800;
      21880: inst = 32'h8620000;
      21881: inst = 32'h2a0e0002;
      21882: inst = 32'h294f0000;
      21883: inst = 32'h11200000;
      21884: inst = 32'hd205580;
      21885: inst = 32'h13e00000;
      21886: inst = 32'hfe0a9fb;
      21887: inst = 32'h5be00000;
      21888: inst = 32'h244c8000;
      21889: inst = 32'h24428800;
      21890: inst = 32'h8620000;
      21891: inst = 32'h2a0e0003;
      21892: inst = 32'h294f0000;
      21893: inst = 32'h11200000;
      21894: inst = 32'hd20558a;
      21895: inst = 32'h13e00000;
      21896: inst = 32'hfe0a9fb;
      21897: inst = 32'h5be00000;
      21898: inst = 32'h244c8000;
      21899: inst = 32'h24428800;
      21900: inst = 32'h8620000;
      21901: inst = 32'h2a0e0004;
      21902: inst = 32'h294f0000;
      21903: inst = 32'h11200000;
      21904: inst = 32'hd205594;
      21905: inst = 32'h13e00000;
      21906: inst = 32'hfe0a9fb;
      21907: inst = 32'h5be00000;
      21908: inst = 32'h244c8000;
      21909: inst = 32'h24428800;
      21910: inst = 32'h8620000;
      21911: inst = 32'h2a0e0005;
      21912: inst = 32'h294f0000;
      21913: inst = 32'h11200000;
      21914: inst = 32'hd20559e;
      21915: inst = 32'h13e00000;
      21916: inst = 32'hfe0a9fb;
      21917: inst = 32'h5be00000;
      21918: inst = 32'h244c8000;
      21919: inst = 32'h24428800;
      21920: inst = 32'h8620000;
      21921: inst = 32'h2a0e0006;
      21922: inst = 32'h294f0000;
      21923: inst = 32'h11200000;
      21924: inst = 32'hd2055a8;
      21925: inst = 32'h13e00000;
      21926: inst = 32'hfe0a9fb;
      21927: inst = 32'h5be00000;
      21928: inst = 32'h244c8000;
      21929: inst = 32'h24428800;
      21930: inst = 32'h8620000;
      21931: inst = 32'h2a0e0007;
      21932: inst = 32'h294f0000;
      21933: inst = 32'h11200000;
      21934: inst = 32'hd2055b2;
      21935: inst = 32'h13e00000;
      21936: inst = 32'hfe0a9fb;
      21937: inst = 32'h5be00000;
      21938: inst = 32'h244c8000;
      21939: inst = 32'h24428800;
      21940: inst = 32'h8620000;
      21941: inst = 32'h2a0e0008;
      21942: inst = 32'h294f0000;
      21943: inst = 32'h11200000;
      21944: inst = 32'hd2055bc;
      21945: inst = 32'h13e00000;
      21946: inst = 32'hfe0a9fb;
      21947: inst = 32'h5be00000;
      21948: inst = 32'h244c8000;
      21949: inst = 32'h24428800;
      21950: inst = 32'h8620000;
      21951: inst = 32'h2a0e0009;
      21952: inst = 32'h294f0000;
      21953: inst = 32'h11200000;
      21954: inst = 32'hd2055c6;
      21955: inst = 32'h13e00000;
      21956: inst = 32'hfe0a9fb;
      21957: inst = 32'h5be00000;
      21958: inst = 32'h244c8000;
      21959: inst = 32'h24428800;
      21960: inst = 32'h8620000;
      21961: inst = 32'h2a0e0000;
      21962: inst = 32'h294f0001;
      21963: inst = 32'h11200000;
      21964: inst = 32'hd2055d0;
      21965: inst = 32'h13e00000;
      21966: inst = 32'hfe0a9fb;
      21967: inst = 32'h5be00000;
      21968: inst = 32'h244c8000;
      21969: inst = 32'h24428800;
      21970: inst = 32'h8620000;
      21971: inst = 32'h2a0e0001;
      21972: inst = 32'h294f0001;
      21973: inst = 32'h11200000;
      21974: inst = 32'hd2055da;
      21975: inst = 32'h13e00000;
      21976: inst = 32'hfe0a9fb;
      21977: inst = 32'h5be00000;
      21978: inst = 32'h244c8000;
      21979: inst = 32'h24428800;
      21980: inst = 32'h8620000;
      21981: inst = 32'h2a0e0002;
      21982: inst = 32'h294f0001;
      21983: inst = 32'h11200000;
      21984: inst = 32'hd2055e4;
      21985: inst = 32'h13e00000;
      21986: inst = 32'hfe0a9fb;
      21987: inst = 32'h5be00000;
      21988: inst = 32'h244c8000;
      21989: inst = 32'h24428800;
      21990: inst = 32'h8620000;
      21991: inst = 32'h2a0e0003;
      21992: inst = 32'h294f0001;
      21993: inst = 32'h11200000;
      21994: inst = 32'hd2055ee;
      21995: inst = 32'h13e00000;
      21996: inst = 32'hfe0a9fb;
      21997: inst = 32'h5be00000;
      21998: inst = 32'h244c8000;
      21999: inst = 32'h24428800;
      22000: inst = 32'h8620000;
      22001: inst = 32'h2a0e0004;
      22002: inst = 32'h294f0001;
      22003: inst = 32'h11200000;
      22004: inst = 32'hd2055f8;
      22005: inst = 32'h13e00000;
      22006: inst = 32'hfe0a9fb;
      22007: inst = 32'h5be00000;
      22008: inst = 32'h244c8000;
      22009: inst = 32'h24428800;
      22010: inst = 32'h8620000;
      22011: inst = 32'h2a0e0005;
      22012: inst = 32'h294f0001;
      22013: inst = 32'h11200000;
      22014: inst = 32'hd205602;
      22015: inst = 32'h13e00000;
      22016: inst = 32'hfe0a9fb;
      22017: inst = 32'h5be00000;
      22018: inst = 32'h244c8000;
      22019: inst = 32'h24428800;
      22020: inst = 32'h8620000;
      22021: inst = 32'h2a0e0006;
      22022: inst = 32'h294f0001;
      22023: inst = 32'h11200000;
      22024: inst = 32'hd20560c;
      22025: inst = 32'h13e00000;
      22026: inst = 32'hfe0a9fb;
      22027: inst = 32'h5be00000;
      22028: inst = 32'h244c8000;
      22029: inst = 32'h24428800;
      22030: inst = 32'h8620000;
      22031: inst = 32'h2a0e0007;
      22032: inst = 32'h294f0001;
      22033: inst = 32'h11200000;
      22034: inst = 32'hd205616;
      22035: inst = 32'h13e00000;
      22036: inst = 32'hfe0a9fb;
      22037: inst = 32'h5be00000;
      22038: inst = 32'h244c8000;
      22039: inst = 32'h24428800;
      22040: inst = 32'h8620000;
      22041: inst = 32'h2a0e0008;
      22042: inst = 32'h294f0001;
      22043: inst = 32'h11200000;
      22044: inst = 32'hd205620;
      22045: inst = 32'h13e00000;
      22046: inst = 32'hfe0a9fb;
      22047: inst = 32'h5be00000;
      22048: inst = 32'h244c8000;
      22049: inst = 32'h24428800;
      22050: inst = 32'h8620000;
      22051: inst = 32'h2a0e0009;
      22052: inst = 32'h294f0001;
      22053: inst = 32'h11200000;
      22054: inst = 32'hd20562a;
      22055: inst = 32'h13e00000;
      22056: inst = 32'hfe0a9fb;
      22057: inst = 32'h5be00000;
      22058: inst = 32'h244c8000;
      22059: inst = 32'h24428800;
      22060: inst = 32'h8620000;
      22061: inst = 32'h2a0e0000;
      22062: inst = 32'h294f0002;
      22063: inst = 32'h11200000;
      22064: inst = 32'hd205634;
      22065: inst = 32'h13e00000;
      22066: inst = 32'hfe0a9fb;
      22067: inst = 32'h5be00000;
      22068: inst = 32'h244c8000;
      22069: inst = 32'h24428800;
      22070: inst = 32'h8620000;
      22071: inst = 32'h2a0e0001;
      22072: inst = 32'h294f0002;
      22073: inst = 32'h11200000;
      22074: inst = 32'hd20563e;
      22075: inst = 32'h13e00000;
      22076: inst = 32'hfe0a9fb;
      22077: inst = 32'h5be00000;
      22078: inst = 32'h244c8000;
      22079: inst = 32'h24428800;
      22080: inst = 32'h8620000;
      22081: inst = 32'h2a0e0002;
      22082: inst = 32'h294f0002;
      22083: inst = 32'h11200000;
      22084: inst = 32'hd205648;
      22085: inst = 32'h13e00000;
      22086: inst = 32'hfe0a9fb;
      22087: inst = 32'h5be00000;
      22088: inst = 32'h244c8000;
      22089: inst = 32'h24428800;
      22090: inst = 32'h8620000;
      22091: inst = 32'h2a0e0003;
      22092: inst = 32'h294f0002;
      22093: inst = 32'h11200000;
      22094: inst = 32'hd205652;
      22095: inst = 32'h13e00000;
      22096: inst = 32'hfe0a9fb;
      22097: inst = 32'h5be00000;
      22098: inst = 32'h244c8000;
      22099: inst = 32'h24428800;
      22100: inst = 32'h8620000;
      22101: inst = 32'h2a0e0004;
      22102: inst = 32'h294f0002;
      22103: inst = 32'h11200000;
      22104: inst = 32'hd20565c;
      22105: inst = 32'h13e00000;
      22106: inst = 32'hfe0a9fb;
      22107: inst = 32'h5be00000;
      22108: inst = 32'h244c8000;
      22109: inst = 32'h24428800;
      22110: inst = 32'h8620000;
      22111: inst = 32'h2a0e0005;
      22112: inst = 32'h294f0002;
      22113: inst = 32'h11200000;
      22114: inst = 32'hd205666;
      22115: inst = 32'h13e00000;
      22116: inst = 32'hfe0a9fb;
      22117: inst = 32'h5be00000;
      22118: inst = 32'h244c8000;
      22119: inst = 32'h24428800;
      22120: inst = 32'h8620000;
      22121: inst = 32'h2a0e0006;
      22122: inst = 32'h294f0002;
      22123: inst = 32'h11200000;
      22124: inst = 32'hd205670;
      22125: inst = 32'h13e00000;
      22126: inst = 32'hfe0a9fb;
      22127: inst = 32'h5be00000;
      22128: inst = 32'h244c8000;
      22129: inst = 32'h24428800;
      22130: inst = 32'h8620000;
      22131: inst = 32'h2a0e0007;
      22132: inst = 32'h294f0002;
      22133: inst = 32'h11200000;
      22134: inst = 32'hd20567a;
      22135: inst = 32'h13e00000;
      22136: inst = 32'hfe0a9fb;
      22137: inst = 32'h5be00000;
      22138: inst = 32'h244c8000;
      22139: inst = 32'h24428800;
      22140: inst = 32'h8620000;
      22141: inst = 32'h2a0e0008;
      22142: inst = 32'h294f0002;
      22143: inst = 32'h11200000;
      22144: inst = 32'hd205684;
      22145: inst = 32'h13e00000;
      22146: inst = 32'hfe0a9fb;
      22147: inst = 32'h5be00000;
      22148: inst = 32'h244c8000;
      22149: inst = 32'h24428800;
      22150: inst = 32'h8620000;
      22151: inst = 32'h2a0e0009;
      22152: inst = 32'h294f0002;
      22153: inst = 32'h11200000;
      22154: inst = 32'hd20568e;
      22155: inst = 32'h13e00000;
      22156: inst = 32'hfe0a9fb;
      22157: inst = 32'h5be00000;
      22158: inst = 32'h244c8000;
      22159: inst = 32'h24428800;
      22160: inst = 32'h8620000;
      22161: inst = 32'h2a0e0000;
      22162: inst = 32'h294f0003;
      22163: inst = 32'h11200000;
      22164: inst = 32'hd205698;
      22165: inst = 32'h13e00000;
      22166: inst = 32'hfe0a9fb;
      22167: inst = 32'h5be00000;
      22168: inst = 32'h244c8000;
      22169: inst = 32'h24428800;
      22170: inst = 32'h8620000;
      22171: inst = 32'h2a0e0001;
      22172: inst = 32'h294f0003;
      22173: inst = 32'h11200000;
      22174: inst = 32'hd2056a2;
      22175: inst = 32'h13e00000;
      22176: inst = 32'hfe0a9fb;
      22177: inst = 32'h5be00000;
      22178: inst = 32'h244c8000;
      22179: inst = 32'h24428800;
      22180: inst = 32'h8620000;
      22181: inst = 32'h2a0e0002;
      22182: inst = 32'h294f0003;
      22183: inst = 32'h11200000;
      22184: inst = 32'hd2056ac;
      22185: inst = 32'h13e00000;
      22186: inst = 32'hfe0a9fb;
      22187: inst = 32'h5be00000;
      22188: inst = 32'h244c8000;
      22189: inst = 32'h24428800;
      22190: inst = 32'h8620000;
      22191: inst = 32'h2a0e0003;
      22192: inst = 32'h294f0003;
      22193: inst = 32'h11200000;
      22194: inst = 32'hd2056b6;
      22195: inst = 32'h13e00000;
      22196: inst = 32'hfe0a9fb;
      22197: inst = 32'h5be00000;
      22198: inst = 32'h244c8000;
      22199: inst = 32'h24428800;
      22200: inst = 32'h8620000;
      22201: inst = 32'h2a0e0004;
      22202: inst = 32'h294f0003;
      22203: inst = 32'h11200000;
      22204: inst = 32'hd2056c0;
      22205: inst = 32'h13e00000;
      22206: inst = 32'hfe0a9fb;
      22207: inst = 32'h5be00000;
      22208: inst = 32'h244c8000;
      22209: inst = 32'h24428800;
      22210: inst = 32'h8620000;
      22211: inst = 32'h2a0e0005;
      22212: inst = 32'h294f0003;
      22213: inst = 32'h11200000;
      22214: inst = 32'hd2056ca;
      22215: inst = 32'h13e00000;
      22216: inst = 32'hfe0a9fb;
      22217: inst = 32'h5be00000;
      22218: inst = 32'h244c8000;
      22219: inst = 32'h24428800;
      22220: inst = 32'h8620000;
      22221: inst = 32'h2a0e0006;
      22222: inst = 32'h294f0003;
      22223: inst = 32'h11200000;
      22224: inst = 32'hd2056d4;
      22225: inst = 32'h13e00000;
      22226: inst = 32'hfe0a9fb;
      22227: inst = 32'h5be00000;
      22228: inst = 32'h244c8000;
      22229: inst = 32'h24428800;
      22230: inst = 32'h8620000;
      22231: inst = 32'h2a0e0007;
      22232: inst = 32'h294f0003;
      22233: inst = 32'h11200000;
      22234: inst = 32'hd2056de;
      22235: inst = 32'h13e00000;
      22236: inst = 32'hfe0a9fb;
      22237: inst = 32'h5be00000;
      22238: inst = 32'h244c8000;
      22239: inst = 32'h24428800;
      22240: inst = 32'h8620000;
      22241: inst = 32'h2a0e0008;
      22242: inst = 32'h294f0003;
      22243: inst = 32'h11200000;
      22244: inst = 32'hd2056e8;
      22245: inst = 32'h13e00000;
      22246: inst = 32'hfe0a9fb;
      22247: inst = 32'h5be00000;
      22248: inst = 32'h244c8000;
      22249: inst = 32'h24428800;
      22250: inst = 32'h8620000;
      22251: inst = 32'h2a0e0009;
      22252: inst = 32'h294f0003;
      22253: inst = 32'h11200000;
      22254: inst = 32'hd2056f2;
      22255: inst = 32'h13e00000;
      22256: inst = 32'hfe0a9fb;
      22257: inst = 32'h5be00000;
      22258: inst = 32'h244c8000;
      22259: inst = 32'h24428800;
      22260: inst = 32'h8620000;
      22261: inst = 32'h2a0e0000;
      22262: inst = 32'h294f0004;
      22263: inst = 32'h11200000;
      22264: inst = 32'hd2056fc;
      22265: inst = 32'h13e00000;
      22266: inst = 32'hfe0a9fb;
      22267: inst = 32'h5be00000;
      22268: inst = 32'h244c8000;
      22269: inst = 32'h24428800;
      22270: inst = 32'h8620000;
      22271: inst = 32'h2a0e0001;
      22272: inst = 32'h294f0004;
      22273: inst = 32'h11200000;
      22274: inst = 32'hd205706;
      22275: inst = 32'h13e00000;
      22276: inst = 32'hfe0a9fb;
      22277: inst = 32'h5be00000;
      22278: inst = 32'h244c8000;
      22279: inst = 32'h24428800;
      22280: inst = 32'h8620000;
      22281: inst = 32'h2a0e0002;
      22282: inst = 32'h294f0004;
      22283: inst = 32'h11200000;
      22284: inst = 32'hd205710;
      22285: inst = 32'h13e00000;
      22286: inst = 32'hfe0a9fb;
      22287: inst = 32'h5be00000;
      22288: inst = 32'h244c8000;
      22289: inst = 32'h24428800;
      22290: inst = 32'h8620000;
      22291: inst = 32'h2a0e0003;
      22292: inst = 32'h294f0004;
      22293: inst = 32'h11200000;
      22294: inst = 32'hd20571a;
      22295: inst = 32'h13e00000;
      22296: inst = 32'hfe0a9fb;
      22297: inst = 32'h5be00000;
      22298: inst = 32'h244c8000;
      22299: inst = 32'h24428800;
      22300: inst = 32'h8620000;
      22301: inst = 32'h2a0e0004;
      22302: inst = 32'h294f0004;
      22303: inst = 32'h11200000;
      22304: inst = 32'hd205724;
      22305: inst = 32'h13e00000;
      22306: inst = 32'hfe0a9fb;
      22307: inst = 32'h5be00000;
      22308: inst = 32'h244c8000;
      22309: inst = 32'h24428800;
      22310: inst = 32'h8620000;
      22311: inst = 32'h2a0e0005;
      22312: inst = 32'h294f0004;
      22313: inst = 32'h11200000;
      22314: inst = 32'hd20572e;
      22315: inst = 32'h13e00000;
      22316: inst = 32'hfe0a9fb;
      22317: inst = 32'h5be00000;
      22318: inst = 32'h244c8000;
      22319: inst = 32'h24428800;
      22320: inst = 32'h8620000;
      22321: inst = 32'h2a0e0006;
      22322: inst = 32'h294f0004;
      22323: inst = 32'h11200000;
      22324: inst = 32'hd205738;
      22325: inst = 32'h13e00000;
      22326: inst = 32'hfe0a9fb;
      22327: inst = 32'h5be00000;
      22328: inst = 32'h244c8000;
      22329: inst = 32'h24428800;
      22330: inst = 32'h8620000;
      22331: inst = 32'h2a0e0007;
      22332: inst = 32'h294f0004;
      22333: inst = 32'h11200000;
      22334: inst = 32'hd205742;
      22335: inst = 32'h13e00000;
      22336: inst = 32'hfe0a9fb;
      22337: inst = 32'h5be00000;
      22338: inst = 32'h244c8000;
      22339: inst = 32'h24428800;
      22340: inst = 32'h8620000;
      22341: inst = 32'h2a0e0008;
      22342: inst = 32'h294f0004;
      22343: inst = 32'h11200000;
      22344: inst = 32'hd20574c;
      22345: inst = 32'h13e00000;
      22346: inst = 32'hfe0a9fb;
      22347: inst = 32'h5be00000;
      22348: inst = 32'h244c8000;
      22349: inst = 32'h24428800;
      22350: inst = 32'h8620000;
      22351: inst = 32'h2a0e0009;
      22352: inst = 32'h294f0004;
      22353: inst = 32'h11200000;
      22354: inst = 32'hd205756;
      22355: inst = 32'h13e00000;
      22356: inst = 32'hfe0a9fb;
      22357: inst = 32'h5be00000;
      22358: inst = 32'h244c8000;
      22359: inst = 32'h24428800;
      22360: inst = 32'h8620000;
      22361: inst = 32'h2a0e0000;
      22362: inst = 32'h294f0005;
      22363: inst = 32'h11200000;
      22364: inst = 32'hd205760;
      22365: inst = 32'h13e00000;
      22366: inst = 32'hfe0a9fb;
      22367: inst = 32'h5be00000;
      22368: inst = 32'h244c8000;
      22369: inst = 32'h24428800;
      22370: inst = 32'h8620000;
      22371: inst = 32'h2a0e0001;
      22372: inst = 32'h294f0005;
      22373: inst = 32'h11200000;
      22374: inst = 32'hd20576a;
      22375: inst = 32'h13e00000;
      22376: inst = 32'hfe0a9fb;
      22377: inst = 32'h5be00000;
      22378: inst = 32'h244c8000;
      22379: inst = 32'h24428800;
      22380: inst = 32'h8620000;
      22381: inst = 32'h2a0e0002;
      22382: inst = 32'h294f0005;
      22383: inst = 32'h11200000;
      22384: inst = 32'hd205774;
      22385: inst = 32'h13e00000;
      22386: inst = 32'hfe0a9fb;
      22387: inst = 32'h5be00000;
      22388: inst = 32'h244c8000;
      22389: inst = 32'h24428800;
      22390: inst = 32'h8620000;
      22391: inst = 32'h2a0e0003;
      22392: inst = 32'h294f0005;
      22393: inst = 32'h11200000;
      22394: inst = 32'hd20577e;
      22395: inst = 32'h13e00000;
      22396: inst = 32'hfe0a9fb;
      22397: inst = 32'h5be00000;
      22398: inst = 32'h244c8000;
      22399: inst = 32'h24428800;
      22400: inst = 32'h8620000;
      22401: inst = 32'h2a0e0004;
      22402: inst = 32'h294f0005;
      22403: inst = 32'h11200000;
      22404: inst = 32'hd205788;
      22405: inst = 32'h13e00000;
      22406: inst = 32'hfe0a9fb;
      22407: inst = 32'h5be00000;
      22408: inst = 32'h244c8000;
      22409: inst = 32'h24428800;
      22410: inst = 32'h8620000;
      22411: inst = 32'h2a0e0005;
      22412: inst = 32'h294f0005;
      22413: inst = 32'h11200000;
      22414: inst = 32'hd205792;
      22415: inst = 32'h13e00000;
      22416: inst = 32'hfe0a9fb;
      22417: inst = 32'h5be00000;
      22418: inst = 32'h244c8000;
      22419: inst = 32'h24428800;
      22420: inst = 32'h8620000;
      22421: inst = 32'h2a0e0006;
      22422: inst = 32'h294f0005;
      22423: inst = 32'h11200000;
      22424: inst = 32'hd20579c;
      22425: inst = 32'h13e00000;
      22426: inst = 32'hfe0a9fb;
      22427: inst = 32'h5be00000;
      22428: inst = 32'h244c8000;
      22429: inst = 32'h24428800;
      22430: inst = 32'h8620000;
      22431: inst = 32'h2a0e0007;
      22432: inst = 32'h294f0005;
      22433: inst = 32'h11200000;
      22434: inst = 32'hd2057a6;
      22435: inst = 32'h13e00000;
      22436: inst = 32'hfe0a9fb;
      22437: inst = 32'h5be00000;
      22438: inst = 32'h244c8000;
      22439: inst = 32'h24428800;
      22440: inst = 32'h8620000;
      22441: inst = 32'h2a0e0008;
      22442: inst = 32'h294f0005;
      22443: inst = 32'h11200000;
      22444: inst = 32'hd2057b0;
      22445: inst = 32'h13e00000;
      22446: inst = 32'hfe0a9fb;
      22447: inst = 32'h5be00000;
      22448: inst = 32'h244c8000;
      22449: inst = 32'h24428800;
      22450: inst = 32'h8620000;
      22451: inst = 32'h2a0e0009;
      22452: inst = 32'h294f0005;
      22453: inst = 32'h11200000;
      22454: inst = 32'hd2057ba;
      22455: inst = 32'h13e00000;
      22456: inst = 32'hfe0a9fb;
      22457: inst = 32'h5be00000;
      22458: inst = 32'h244c8000;
      22459: inst = 32'h24428800;
      22460: inst = 32'h8620000;
      22461: inst = 32'h2a0e0000;
      22462: inst = 32'h294f0006;
      22463: inst = 32'h11200000;
      22464: inst = 32'hd2057c4;
      22465: inst = 32'h13e00000;
      22466: inst = 32'hfe0a9fb;
      22467: inst = 32'h5be00000;
      22468: inst = 32'h244c8000;
      22469: inst = 32'h24428800;
      22470: inst = 32'h8620000;
      22471: inst = 32'h2a0e0001;
      22472: inst = 32'h294f0006;
      22473: inst = 32'h11200000;
      22474: inst = 32'hd2057ce;
      22475: inst = 32'h13e00000;
      22476: inst = 32'hfe0a9fb;
      22477: inst = 32'h5be00000;
      22478: inst = 32'h244c8000;
      22479: inst = 32'h24428800;
      22480: inst = 32'h8620000;
      22481: inst = 32'h2a0e0002;
      22482: inst = 32'h294f0006;
      22483: inst = 32'h11200000;
      22484: inst = 32'hd2057d8;
      22485: inst = 32'h13e00000;
      22486: inst = 32'hfe0a9fb;
      22487: inst = 32'h5be00000;
      22488: inst = 32'h244c8000;
      22489: inst = 32'h24428800;
      22490: inst = 32'h8620000;
      22491: inst = 32'h2a0e0003;
      22492: inst = 32'h294f0006;
      22493: inst = 32'h11200000;
      22494: inst = 32'hd2057e2;
      22495: inst = 32'h13e00000;
      22496: inst = 32'hfe0a9fb;
      22497: inst = 32'h5be00000;
      22498: inst = 32'h244c8000;
      22499: inst = 32'h24428800;
      22500: inst = 32'h8620000;
      22501: inst = 32'h2a0e0004;
      22502: inst = 32'h294f0006;
      22503: inst = 32'h11200000;
      22504: inst = 32'hd2057ec;
      22505: inst = 32'h13e00000;
      22506: inst = 32'hfe0a9fb;
      22507: inst = 32'h5be00000;
      22508: inst = 32'h244c8000;
      22509: inst = 32'h24428800;
      22510: inst = 32'h8620000;
      22511: inst = 32'h2a0e0005;
      22512: inst = 32'h294f0006;
      22513: inst = 32'h11200000;
      22514: inst = 32'hd2057f6;
      22515: inst = 32'h13e00000;
      22516: inst = 32'hfe0a9fb;
      22517: inst = 32'h5be00000;
      22518: inst = 32'h244c8000;
      22519: inst = 32'h24428800;
      22520: inst = 32'h8620000;
      22521: inst = 32'h2a0e0006;
      22522: inst = 32'h294f0006;
      22523: inst = 32'h11200000;
      22524: inst = 32'hd205800;
      22525: inst = 32'h13e00000;
      22526: inst = 32'hfe0a9fb;
      22527: inst = 32'h5be00000;
      22528: inst = 32'h244c8000;
      22529: inst = 32'h24428800;
      22530: inst = 32'h8620000;
      22531: inst = 32'h2a0e0007;
      22532: inst = 32'h294f0006;
      22533: inst = 32'h11200000;
      22534: inst = 32'hd20580a;
      22535: inst = 32'h13e00000;
      22536: inst = 32'hfe0a9fb;
      22537: inst = 32'h5be00000;
      22538: inst = 32'h244c8000;
      22539: inst = 32'h24428800;
      22540: inst = 32'h8620000;
      22541: inst = 32'h2a0e0008;
      22542: inst = 32'h294f0006;
      22543: inst = 32'h11200000;
      22544: inst = 32'hd205814;
      22545: inst = 32'h13e00000;
      22546: inst = 32'hfe0a9fb;
      22547: inst = 32'h5be00000;
      22548: inst = 32'h244c8000;
      22549: inst = 32'h24428800;
      22550: inst = 32'h8620000;
      22551: inst = 32'h2a0e0009;
      22552: inst = 32'h294f0006;
      22553: inst = 32'h11200000;
      22554: inst = 32'hd20581e;
      22555: inst = 32'h13e00000;
      22556: inst = 32'hfe0a9fb;
      22557: inst = 32'h5be00000;
      22558: inst = 32'h244c8000;
      22559: inst = 32'h24428800;
      22560: inst = 32'h8620000;
      22561: inst = 32'hc60f4ce;
      22562: inst = 32'h2a0e0001;
      22563: inst = 32'h294f0007;
      22564: inst = 32'h11200000;
      22565: inst = 32'hd205829;
      22566: inst = 32'h13e00000;
      22567: inst = 32'hfe0a9fb;
      22568: inst = 32'h5be00000;
      22569: inst = 32'h244c8000;
      22570: inst = 32'h24428800;
      22571: inst = 32'h8620000;
      22572: inst = 32'h2a0e0008;
      22573: inst = 32'h294f0007;
      22574: inst = 32'h11200000;
      22575: inst = 32'hd205833;
      22576: inst = 32'h13e00000;
      22577: inst = 32'hfe0a9fb;
      22578: inst = 32'h5be00000;
      22579: inst = 32'h244c8000;
      22580: inst = 32'h24428800;
      22581: inst = 32'h8620000;
      22582: inst = 32'h2a0e0001;
      22583: inst = 32'h294f0008;
      22584: inst = 32'h11200000;
      22585: inst = 32'hd20583d;
      22586: inst = 32'h13e00000;
      22587: inst = 32'hfe0a9fb;
      22588: inst = 32'h5be00000;
      22589: inst = 32'h244c8000;
      22590: inst = 32'h24428800;
      22591: inst = 32'h8620000;
      22592: inst = 32'h2a0e0008;
      22593: inst = 32'h294f0008;
      22594: inst = 32'h11200000;
      22595: inst = 32'hd205847;
      22596: inst = 32'h13e00000;
      22597: inst = 32'hfe0a9fb;
      22598: inst = 32'h5be00000;
      22599: inst = 32'h244c8000;
      22600: inst = 32'h24428800;
      22601: inst = 32'h8620000;
      22602: inst = 32'hc607841;
      22603: inst = 32'h2a0e0002;
      22604: inst = 32'h294f0007;
      22605: inst = 32'h11200000;
      22606: inst = 32'hd205852;
      22607: inst = 32'h13e00000;
      22608: inst = 32'hfe0a9fb;
      22609: inst = 32'h5be00000;
      22610: inst = 32'h244c8000;
      22611: inst = 32'h24428800;
      22612: inst = 32'h8620000;
      22613: inst = 32'h2a0e0003;
      22614: inst = 32'h294f0007;
      22615: inst = 32'h11200000;
      22616: inst = 32'hd20585c;
      22617: inst = 32'h13e00000;
      22618: inst = 32'hfe0a9fb;
      22619: inst = 32'h5be00000;
      22620: inst = 32'h244c8000;
      22621: inst = 32'h24428800;
      22622: inst = 32'h8620000;
      22623: inst = 32'h2a0e0004;
      22624: inst = 32'h294f0007;
      22625: inst = 32'h11200000;
      22626: inst = 32'hd205866;
      22627: inst = 32'h13e00000;
      22628: inst = 32'hfe0a9fb;
      22629: inst = 32'h5be00000;
      22630: inst = 32'h244c8000;
      22631: inst = 32'h24428800;
      22632: inst = 32'h8620000;
      22633: inst = 32'h2a0e0005;
      22634: inst = 32'h294f0007;
      22635: inst = 32'h11200000;
      22636: inst = 32'hd205870;
      22637: inst = 32'h13e00000;
      22638: inst = 32'hfe0a9fb;
      22639: inst = 32'h5be00000;
      22640: inst = 32'h244c8000;
      22641: inst = 32'h24428800;
      22642: inst = 32'h8620000;
      22643: inst = 32'h2a0e0006;
      22644: inst = 32'h294f0007;
      22645: inst = 32'h11200000;
      22646: inst = 32'hd20587a;
      22647: inst = 32'h13e00000;
      22648: inst = 32'hfe0a9fb;
      22649: inst = 32'h5be00000;
      22650: inst = 32'h244c8000;
      22651: inst = 32'h24428800;
      22652: inst = 32'h8620000;
      22653: inst = 32'h2a0e0007;
      22654: inst = 32'h294f0007;
      22655: inst = 32'h11200000;
      22656: inst = 32'hd205884;
      22657: inst = 32'h13e00000;
      22658: inst = 32'hfe0a9fb;
      22659: inst = 32'h5be00000;
      22660: inst = 32'h244c8000;
      22661: inst = 32'h24428800;
      22662: inst = 32'h8620000;
      22663: inst = 32'h2a0e0002;
      22664: inst = 32'h294f0008;
      22665: inst = 32'h11200000;
      22666: inst = 32'hd20588e;
      22667: inst = 32'h13e00000;
      22668: inst = 32'hfe0a9fb;
      22669: inst = 32'h5be00000;
      22670: inst = 32'h244c8000;
      22671: inst = 32'h24428800;
      22672: inst = 32'h8620000;
      22673: inst = 32'h2a0e0003;
      22674: inst = 32'h294f0008;
      22675: inst = 32'h11200000;
      22676: inst = 32'hd205898;
      22677: inst = 32'h13e00000;
      22678: inst = 32'hfe0a9fb;
      22679: inst = 32'h5be00000;
      22680: inst = 32'h244c8000;
      22681: inst = 32'h24428800;
      22682: inst = 32'h8620000;
      22683: inst = 32'h2a0e0004;
      22684: inst = 32'h294f0008;
      22685: inst = 32'h11200000;
      22686: inst = 32'hd2058a2;
      22687: inst = 32'h13e00000;
      22688: inst = 32'hfe0a9fb;
      22689: inst = 32'h5be00000;
      22690: inst = 32'h244c8000;
      22691: inst = 32'h24428800;
      22692: inst = 32'h8620000;
      22693: inst = 32'h2a0e0005;
      22694: inst = 32'h294f0008;
      22695: inst = 32'h11200000;
      22696: inst = 32'hd2058ac;
      22697: inst = 32'h13e00000;
      22698: inst = 32'hfe0a9fb;
      22699: inst = 32'h5be00000;
      22700: inst = 32'h244c8000;
      22701: inst = 32'h24428800;
      22702: inst = 32'h8620000;
      22703: inst = 32'h2a0e0006;
      22704: inst = 32'h294f0008;
      22705: inst = 32'h11200000;
      22706: inst = 32'hd2058b6;
      22707: inst = 32'h13e00000;
      22708: inst = 32'hfe0a9fb;
      22709: inst = 32'h5be00000;
      22710: inst = 32'h244c8000;
      22711: inst = 32'h24428800;
      22712: inst = 32'h8620000;
      22713: inst = 32'h2a0e0007;
      22714: inst = 32'h294f0008;
      22715: inst = 32'h11200000;
      22716: inst = 32'hd2058c0;
      22717: inst = 32'h13e00000;
      22718: inst = 32'hfe0a9fb;
      22719: inst = 32'h5be00000;
      22720: inst = 32'h244c8000;
      22721: inst = 32'h24428800;
      22722: inst = 32'h8620000;
      22723: inst = 32'h2a0e0002;
      22724: inst = 32'h294f0009;
      22725: inst = 32'h11200000;
      22726: inst = 32'hd2058ca;
      22727: inst = 32'h13e00000;
      22728: inst = 32'hfe0a9fb;
      22729: inst = 32'h5be00000;
      22730: inst = 32'h244c8000;
      22731: inst = 32'h24428800;
      22732: inst = 32'h8620000;
      22733: inst = 32'h2a0e0003;
      22734: inst = 32'h294f0009;
      22735: inst = 32'h11200000;
      22736: inst = 32'hd2058d4;
      22737: inst = 32'h13e00000;
      22738: inst = 32'hfe0a9fb;
      22739: inst = 32'h5be00000;
      22740: inst = 32'h244c8000;
      22741: inst = 32'h24428800;
      22742: inst = 32'h8620000;
      22743: inst = 32'h2a0e0004;
      22744: inst = 32'h294f0009;
      22745: inst = 32'h11200000;
      22746: inst = 32'hd2058de;
      22747: inst = 32'h13e00000;
      22748: inst = 32'hfe0a9fb;
      22749: inst = 32'h5be00000;
      22750: inst = 32'h244c8000;
      22751: inst = 32'h24428800;
      22752: inst = 32'h8620000;
      22753: inst = 32'h2a0e0005;
      22754: inst = 32'h294f0009;
      22755: inst = 32'h11200000;
      22756: inst = 32'hd2058e8;
      22757: inst = 32'h13e00000;
      22758: inst = 32'hfe0a9fb;
      22759: inst = 32'h5be00000;
      22760: inst = 32'h244c8000;
      22761: inst = 32'h24428800;
      22762: inst = 32'h8620000;
      22763: inst = 32'h2a0e0006;
      22764: inst = 32'h294f0009;
      22765: inst = 32'h11200000;
      22766: inst = 32'hd2058f2;
      22767: inst = 32'h13e00000;
      22768: inst = 32'hfe0a9fb;
      22769: inst = 32'h5be00000;
      22770: inst = 32'h244c8000;
      22771: inst = 32'h24428800;
      22772: inst = 32'h8620000;
      22773: inst = 32'h2a0e0007;
      22774: inst = 32'h294f0009;
      22775: inst = 32'h11200000;
      22776: inst = 32'hd2058fc;
      22777: inst = 32'h13e00000;
      22778: inst = 32'hfe0a9fb;
      22779: inst = 32'h5be00000;
      22780: inst = 32'h244c8000;
      22781: inst = 32'h24428800;
      22782: inst = 32'h8620000;
      22783: inst = 32'hc6010ac;
      22784: inst = 32'h2a0e0002;
      22785: inst = 32'h294f000a;
      22786: inst = 32'h11200000;
      22787: inst = 32'hd205907;
      22788: inst = 32'h13e00000;
      22789: inst = 32'hfe0a9fb;
      22790: inst = 32'h5be00000;
      22791: inst = 32'h244c8000;
      22792: inst = 32'h24428800;
      22793: inst = 32'h8620000;
      22794: inst = 32'h2a0e0003;
      22795: inst = 32'h294f000a;
      22796: inst = 32'h11200000;
      22797: inst = 32'hd205911;
      22798: inst = 32'h13e00000;
      22799: inst = 32'hfe0a9fb;
      22800: inst = 32'h5be00000;
      22801: inst = 32'h244c8000;
      22802: inst = 32'h24428800;
      22803: inst = 32'h8620000;
      22804: inst = 32'h2a0e0004;
      22805: inst = 32'h294f000a;
      22806: inst = 32'h11200000;
      22807: inst = 32'hd20591b;
      22808: inst = 32'h13e00000;
      22809: inst = 32'hfe0a9fb;
      22810: inst = 32'h5be00000;
      22811: inst = 32'h244c8000;
      22812: inst = 32'h24428800;
      22813: inst = 32'h8620000;
      22814: inst = 32'h2a0e0005;
      22815: inst = 32'h294f000a;
      22816: inst = 32'h11200000;
      22817: inst = 32'hd205925;
      22818: inst = 32'h13e00000;
      22819: inst = 32'hfe0a9fb;
      22820: inst = 32'h5be00000;
      22821: inst = 32'h244c8000;
      22822: inst = 32'h24428800;
      22823: inst = 32'h8620000;
      22824: inst = 32'h2a0e0006;
      22825: inst = 32'h294f000a;
      22826: inst = 32'h11200000;
      22827: inst = 32'hd20592f;
      22828: inst = 32'h13e00000;
      22829: inst = 32'hfe0a9fb;
      22830: inst = 32'h5be00000;
      22831: inst = 32'h244c8000;
      22832: inst = 32'h24428800;
      22833: inst = 32'h8620000;
      22834: inst = 32'h2a0e0007;
      22835: inst = 32'h294f000a;
      22836: inst = 32'h11200000;
      22837: inst = 32'hd205939;
      22838: inst = 32'h13e00000;
      22839: inst = 32'hfe0a9fb;
      22840: inst = 32'h5be00000;
      22841: inst = 32'h244c8000;
      22842: inst = 32'h24428800;
      22843: inst = 32'h8620000;
      22844: inst = 32'hc60d42c;
      22845: inst = 32'h2a0e0003;
      22846: inst = 32'h294f000b;
      22847: inst = 32'h11200000;
      22848: inst = 32'hd205944;
      22849: inst = 32'h13e00000;
      22850: inst = 32'hfe0a9fb;
      22851: inst = 32'h5be00000;
      22852: inst = 32'h244c8000;
      22853: inst = 32'h24428800;
      22854: inst = 32'h8620000;
      22855: inst = 32'h2a0e0006;
      22856: inst = 32'h294f000b;
      22857: inst = 32'h11200000;
      22858: inst = 32'hd20594e;
      22859: inst = 32'h13e00000;
      22860: inst = 32'hfe0a9fb;
      22861: inst = 32'h5be00000;
      22862: inst = 32'h244c8000;
      22863: inst = 32'h24428800;
      22864: inst = 32'h8620000;
      22865: inst = 32'h13e00000;
      22866: inst = 32'hfe06108;
      22867: inst = 32'h5be00000;
      22868: inst = 32'hc6018c3;
      22869: inst = 32'h2a0e0000;
      22870: inst = 32'h294f0000;
      22871: inst = 32'h11200000;
      22872: inst = 32'hd20595c;
      22873: inst = 32'h13e00000;
      22874: inst = 32'hfe0a9fb;
      22875: inst = 32'h5be00000;
      22876: inst = 32'h244c8000;
      22877: inst = 32'h24428800;
      22878: inst = 32'h8620000;
      22879: inst = 32'h2a0e0001;
      22880: inst = 32'h294f0000;
      22881: inst = 32'h11200000;
      22882: inst = 32'hd205966;
      22883: inst = 32'h13e00000;
      22884: inst = 32'hfe0a9fb;
      22885: inst = 32'h5be00000;
      22886: inst = 32'h244c8000;
      22887: inst = 32'h24428800;
      22888: inst = 32'h8620000;
      22889: inst = 32'h2a0e0002;
      22890: inst = 32'h294f0000;
      22891: inst = 32'h11200000;
      22892: inst = 32'hd205970;
      22893: inst = 32'h13e00000;
      22894: inst = 32'hfe0a9fb;
      22895: inst = 32'h5be00000;
      22896: inst = 32'h244c8000;
      22897: inst = 32'h24428800;
      22898: inst = 32'h8620000;
      22899: inst = 32'h2a0e0003;
      22900: inst = 32'h294f0000;
      22901: inst = 32'h11200000;
      22902: inst = 32'hd20597a;
      22903: inst = 32'h13e00000;
      22904: inst = 32'hfe0a9fb;
      22905: inst = 32'h5be00000;
      22906: inst = 32'h244c8000;
      22907: inst = 32'h24428800;
      22908: inst = 32'h8620000;
      22909: inst = 32'h2a0e0004;
      22910: inst = 32'h294f0000;
      22911: inst = 32'h11200000;
      22912: inst = 32'hd205984;
      22913: inst = 32'h13e00000;
      22914: inst = 32'hfe0a9fb;
      22915: inst = 32'h5be00000;
      22916: inst = 32'h244c8000;
      22917: inst = 32'h24428800;
      22918: inst = 32'h8620000;
      22919: inst = 32'h2a0e0005;
      22920: inst = 32'h294f0000;
      22921: inst = 32'h11200000;
      22922: inst = 32'hd20598e;
      22923: inst = 32'h13e00000;
      22924: inst = 32'hfe0a9fb;
      22925: inst = 32'h5be00000;
      22926: inst = 32'h244c8000;
      22927: inst = 32'h24428800;
      22928: inst = 32'h8620000;
      22929: inst = 32'h2a0e0006;
      22930: inst = 32'h294f0000;
      22931: inst = 32'h11200000;
      22932: inst = 32'hd205998;
      22933: inst = 32'h13e00000;
      22934: inst = 32'hfe0a9fb;
      22935: inst = 32'h5be00000;
      22936: inst = 32'h244c8000;
      22937: inst = 32'h24428800;
      22938: inst = 32'h8620000;
      22939: inst = 32'h2a0e0007;
      22940: inst = 32'h294f0000;
      22941: inst = 32'h11200000;
      22942: inst = 32'hd2059a2;
      22943: inst = 32'h13e00000;
      22944: inst = 32'hfe0a9fb;
      22945: inst = 32'h5be00000;
      22946: inst = 32'h244c8000;
      22947: inst = 32'h24428800;
      22948: inst = 32'h8620000;
      22949: inst = 32'h2a0e0008;
      22950: inst = 32'h294f0000;
      22951: inst = 32'h11200000;
      22952: inst = 32'hd2059ac;
      22953: inst = 32'h13e00000;
      22954: inst = 32'hfe0a9fb;
      22955: inst = 32'h5be00000;
      22956: inst = 32'h244c8000;
      22957: inst = 32'h24428800;
      22958: inst = 32'h8620000;
      22959: inst = 32'h2a0e0009;
      22960: inst = 32'h294f0000;
      22961: inst = 32'h11200000;
      22962: inst = 32'hd2059b6;
      22963: inst = 32'h13e00000;
      22964: inst = 32'hfe0a9fb;
      22965: inst = 32'h5be00000;
      22966: inst = 32'h244c8000;
      22967: inst = 32'h24428800;
      22968: inst = 32'h8620000;
      22969: inst = 32'h2a0e0000;
      22970: inst = 32'h294f0001;
      22971: inst = 32'h11200000;
      22972: inst = 32'hd2059c0;
      22973: inst = 32'h13e00000;
      22974: inst = 32'hfe0a9fb;
      22975: inst = 32'h5be00000;
      22976: inst = 32'h244c8000;
      22977: inst = 32'h24428800;
      22978: inst = 32'h8620000;
      22979: inst = 32'h2a0e0001;
      22980: inst = 32'h294f0001;
      22981: inst = 32'h11200000;
      22982: inst = 32'hd2059ca;
      22983: inst = 32'h13e00000;
      22984: inst = 32'hfe0a9fb;
      22985: inst = 32'h5be00000;
      22986: inst = 32'h244c8000;
      22987: inst = 32'h24428800;
      22988: inst = 32'h8620000;
      22989: inst = 32'h2a0e0002;
      22990: inst = 32'h294f0001;
      22991: inst = 32'h11200000;
      22992: inst = 32'hd2059d4;
      22993: inst = 32'h13e00000;
      22994: inst = 32'hfe0a9fb;
      22995: inst = 32'h5be00000;
      22996: inst = 32'h244c8000;
      22997: inst = 32'h24428800;
      22998: inst = 32'h8620000;
      22999: inst = 32'h2a0e0003;
      23000: inst = 32'h294f0001;
      23001: inst = 32'h11200000;
      23002: inst = 32'hd2059de;
      23003: inst = 32'h13e00000;
      23004: inst = 32'hfe0a9fb;
      23005: inst = 32'h5be00000;
      23006: inst = 32'h244c8000;
      23007: inst = 32'h24428800;
      23008: inst = 32'h8620000;
      23009: inst = 32'h2a0e0004;
      23010: inst = 32'h294f0001;
      23011: inst = 32'h11200000;
      23012: inst = 32'hd2059e8;
      23013: inst = 32'h13e00000;
      23014: inst = 32'hfe0a9fb;
      23015: inst = 32'h5be00000;
      23016: inst = 32'h244c8000;
      23017: inst = 32'h24428800;
      23018: inst = 32'h8620000;
      23019: inst = 32'h2a0e0005;
      23020: inst = 32'h294f0001;
      23021: inst = 32'h11200000;
      23022: inst = 32'hd2059f2;
      23023: inst = 32'h13e00000;
      23024: inst = 32'hfe0a9fb;
      23025: inst = 32'h5be00000;
      23026: inst = 32'h244c8000;
      23027: inst = 32'h24428800;
      23028: inst = 32'h8620000;
      23029: inst = 32'h2a0e0006;
      23030: inst = 32'h294f0001;
      23031: inst = 32'h11200000;
      23032: inst = 32'hd2059fc;
      23033: inst = 32'h13e00000;
      23034: inst = 32'hfe0a9fb;
      23035: inst = 32'h5be00000;
      23036: inst = 32'h244c8000;
      23037: inst = 32'h24428800;
      23038: inst = 32'h8620000;
      23039: inst = 32'h2a0e0007;
      23040: inst = 32'h294f0001;
      23041: inst = 32'h11200000;
      23042: inst = 32'hd205a06;
      23043: inst = 32'h13e00000;
      23044: inst = 32'hfe0a9fb;
      23045: inst = 32'h5be00000;
      23046: inst = 32'h244c8000;
      23047: inst = 32'h24428800;
      23048: inst = 32'h8620000;
      23049: inst = 32'h2a0e0008;
      23050: inst = 32'h294f0001;
      23051: inst = 32'h11200000;
      23052: inst = 32'hd205a10;
      23053: inst = 32'h13e00000;
      23054: inst = 32'hfe0a9fb;
      23055: inst = 32'h5be00000;
      23056: inst = 32'h244c8000;
      23057: inst = 32'h24428800;
      23058: inst = 32'h8620000;
      23059: inst = 32'h2a0e0009;
      23060: inst = 32'h294f0001;
      23061: inst = 32'h11200000;
      23062: inst = 32'hd205a1a;
      23063: inst = 32'h13e00000;
      23064: inst = 32'hfe0a9fb;
      23065: inst = 32'h5be00000;
      23066: inst = 32'h244c8000;
      23067: inst = 32'h24428800;
      23068: inst = 32'h8620000;
      23069: inst = 32'h2a0e0000;
      23070: inst = 32'h294f0002;
      23071: inst = 32'h11200000;
      23072: inst = 32'hd205a24;
      23073: inst = 32'h13e00000;
      23074: inst = 32'hfe0a9fb;
      23075: inst = 32'h5be00000;
      23076: inst = 32'h244c8000;
      23077: inst = 32'h24428800;
      23078: inst = 32'h8620000;
      23079: inst = 32'h2a0e0001;
      23080: inst = 32'h294f0002;
      23081: inst = 32'h11200000;
      23082: inst = 32'hd205a2e;
      23083: inst = 32'h13e00000;
      23084: inst = 32'hfe0a9fb;
      23085: inst = 32'h5be00000;
      23086: inst = 32'h244c8000;
      23087: inst = 32'h24428800;
      23088: inst = 32'h8620000;
      23089: inst = 32'h2a0e0000;
      23090: inst = 32'h294f0003;
      23091: inst = 32'h11200000;
      23092: inst = 32'hd205a38;
      23093: inst = 32'h13e00000;
      23094: inst = 32'hfe0a9fb;
      23095: inst = 32'h5be00000;
      23096: inst = 32'h244c8000;
      23097: inst = 32'h24428800;
      23098: inst = 32'h8620000;
      23099: inst = 32'h2a0e0008;
      23100: inst = 32'h294f0003;
      23101: inst = 32'h11200000;
      23102: inst = 32'hd205a42;
      23103: inst = 32'h13e00000;
      23104: inst = 32'hfe0a9fb;
      23105: inst = 32'h5be00000;
      23106: inst = 32'h244c8000;
      23107: inst = 32'h24428800;
      23108: inst = 32'h8620000;
      23109: inst = 32'h2a0e0000;
      23110: inst = 32'h294f0004;
      23111: inst = 32'h11200000;
      23112: inst = 32'hd205a4c;
      23113: inst = 32'h13e00000;
      23114: inst = 32'hfe0a9fb;
      23115: inst = 32'h5be00000;
      23116: inst = 32'h244c8000;
      23117: inst = 32'h24428800;
      23118: inst = 32'h8620000;
      23119: inst = 32'h2a0e0008;
      23120: inst = 32'h294f0004;
      23121: inst = 32'h11200000;
      23122: inst = 32'hd205a56;
      23123: inst = 32'h13e00000;
      23124: inst = 32'hfe0a9fb;
      23125: inst = 32'h5be00000;
      23126: inst = 32'h244c8000;
      23127: inst = 32'h24428800;
      23128: inst = 32'h8620000;
      23129: inst = 32'h2a0e0000;
      23130: inst = 32'h294f0005;
      23131: inst = 32'h11200000;
      23132: inst = 32'hd205a60;
      23133: inst = 32'h13e00000;
      23134: inst = 32'hfe0a9fb;
      23135: inst = 32'h5be00000;
      23136: inst = 32'h244c8000;
      23137: inst = 32'h24428800;
      23138: inst = 32'h8620000;
      23139: inst = 32'h2a0e0001;
      23140: inst = 32'h294f0005;
      23141: inst = 32'h11200000;
      23142: inst = 32'hd205a6a;
      23143: inst = 32'h13e00000;
      23144: inst = 32'hfe0a9fb;
      23145: inst = 32'h5be00000;
      23146: inst = 32'h244c8000;
      23147: inst = 32'h24428800;
      23148: inst = 32'h8620000;
      23149: inst = 32'h2a0e0000;
      23150: inst = 32'h294f0006;
      23151: inst = 32'h11200000;
      23152: inst = 32'hd205a74;
      23153: inst = 32'h13e00000;
      23154: inst = 32'hfe0a9fb;
      23155: inst = 32'h5be00000;
      23156: inst = 32'h244c8000;
      23157: inst = 32'h24428800;
      23158: inst = 32'h8620000;
      23159: inst = 32'h2a0e0001;
      23160: inst = 32'h294f0006;
      23161: inst = 32'h11200000;
      23162: inst = 32'hd205a7e;
      23163: inst = 32'h13e00000;
      23164: inst = 32'hfe0a9fb;
      23165: inst = 32'h5be00000;
      23166: inst = 32'h244c8000;
      23167: inst = 32'h24428800;
      23168: inst = 32'h8620000;
      23169: inst = 32'hc60d42c;
      23170: inst = 32'h2a0e0002;
      23171: inst = 32'h294f0002;
      23172: inst = 32'h11200000;
      23173: inst = 32'hd205a89;
      23174: inst = 32'h13e00000;
      23175: inst = 32'hfe0a9fb;
      23176: inst = 32'h5be00000;
      23177: inst = 32'h244c8000;
      23178: inst = 32'h24428800;
      23179: inst = 32'h8620000;
      23180: inst = 32'h2a0e0003;
      23181: inst = 32'h294f0002;
      23182: inst = 32'h11200000;
      23183: inst = 32'hd205a93;
      23184: inst = 32'h13e00000;
      23185: inst = 32'hfe0a9fb;
      23186: inst = 32'h5be00000;
      23187: inst = 32'h244c8000;
      23188: inst = 32'h24428800;
      23189: inst = 32'h8620000;
      23190: inst = 32'h2a0e0004;
      23191: inst = 32'h294f0002;
      23192: inst = 32'h11200000;
      23193: inst = 32'hd205a9d;
      23194: inst = 32'h13e00000;
      23195: inst = 32'hfe0a9fb;
      23196: inst = 32'h5be00000;
      23197: inst = 32'h244c8000;
      23198: inst = 32'h24428800;
      23199: inst = 32'h8620000;
      23200: inst = 32'h2a0e0005;
      23201: inst = 32'h294f0002;
      23202: inst = 32'h11200000;
      23203: inst = 32'hd205aa7;
      23204: inst = 32'h13e00000;
      23205: inst = 32'hfe0a9fb;
      23206: inst = 32'h5be00000;
      23207: inst = 32'h244c8000;
      23208: inst = 32'h24428800;
      23209: inst = 32'h8620000;
      23210: inst = 32'h2a0e0006;
      23211: inst = 32'h294f0002;
      23212: inst = 32'h11200000;
      23213: inst = 32'hd205ab1;
      23214: inst = 32'h13e00000;
      23215: inst = 32'hfe0a9fb;
      23216: inst = 32'h5be00000;
      23217: inst = 32'h244c8000;
      23218: inst = 32'h24428800;
      23219: inst = 32'h8620000;
      23220: inst = 32'h2a0e0007;
      23221: inst = 32'h294f0002;
      23222: inst = 32'h11200000;
      23223: inst = 32'hd205abb;
      23224: inst = 32'h13e00000;
      23225: inst = 32'hfe0a9fb;
      23226: inst = 32'h5be00000;
      23227: inst = 32'h244c8000;
      23228: inst = 32'h24428800;
      23229: inst = 32'h8620000;
      23230: inst = 32'h2a0e0008;
      23231: inst = 32'h294f0002;
      23232: inst = 32'h11200000;
      23233: inst = 32'hd205ac5;
      23234: inst = 32'h13e00000;
      23235: inst = 32'hfe0a9fb;
      23236: inst = 32'h5be00000;
      23237: inst = 32'h244c8000;
      23238: inst = 32'h24428800;
      23239: inst = 32'h8620000;
      23240: inst = 32'h2a0e0009;
      23241: inst = 32'h294f0002;
      23242: inst = 32'h11200000;
      23243: inst = 32'hd205acf;
      23244: inst = 32'h13e00000;
      23245: inst = 32'hfe0a9fb;
      23246: inst = 32'h5be00000;
      23247: inst = 32'h244c8000;
      23248: inst = 32'h24428800;
      23249: inst = 32'h8620000;
      23250: inst = 32'h2a0e0002;
      23251: inst = 32'h294f0005;
      23252: inst = 32'h11200000;
      23253: inst = 32'hd205ad9;
      23254: inst = 32'h13e00000;
      23255: inst = 32'hfe0a9fb;
      23256: inst = 32'h5be00000;
      23257: inst = 32'h244c8000;
      23258: inst = 32'h24428800;
      23259: inst = 32'h8620000;
      23260: inst = 32'h2a0e0002;
      23261: inst = 32'h294f0006;
      23262: inst = 32'h11200000;
      23263: inst = 32'hd205ae3;
      23264: inst = 32'h13e00000;
      23265: inst = 32'hfe0a9fb;
      23266: inst = 32'h5be00000;
      23267: inst = 32'h244c8000;
      23268: inst = 32'h24428800;
      23269: inst = 32'h8620000;
      23270: inst = 32'h2a0e0003;
      23271: inst = 32'h294f000b;
      23272: inst = 32'h11200000;
      23273: inst = 32'hd205aed;
      23274: inst = 32'h13e00000;
      23275: inst = 32'hfe0a9fb;
      23276: inst = 32'h5be00000;
      23277: inst = 32'h244c8000;
      23278: inst = 32'h24428800;
      23279: inst = 32'h8620000;
      23280: inst = 32'h2a0e0006;
      23281: inst = 32'h294f000b;
      23282: inst = 32'h11200000;
      23283: inst = 32'hd205af7;
      23284: inst = 32'h13e00000;
      23285: inst = 32'hfe0a9fb;
      23286: inst = 32'h5be00000;
      23287: inst = 32'h244c8000;
      23288: inst = 32'h24428800;
      23289: inst = 32'h8620000;
      23290: inst = 32'hc60f4ce;
      23291: inst = 32'h2a0e0001;
      23292: inst = 32'h294f0003;
      23293: inst = 32'h11200000;
      23294: inst = 32'hd205b02;
      23295: inst = 32'h13e00000;
      23296: inst = 32'hfe0a9fb;
      23297: inst = 32'h5be00000;
      23298: inst = 32'h244c8000;
      23299: inst = 32'h24428800;
      23300: inst = 32'h8620000;
      23301: inst = 32'h2a0e0002;
      23302: inst = 32'h294f0003;
      23303: inst = 32'h11200000;
      23304: inst = 32'hd205b0c;
      23305: inst = 32'h13e00000;
      23306: inst = 32'hfe0a9fb;
      23307: inst = 32'h5be00000;
      23308: inst = 32'h244c8000;
      23309: inst = 32'h24428800;
      23310: inst = 32'h8620000;
      23311: inst = 32'h2a0e0003;
      23312: inst = 32'h294f0003;
      23313: inst = 32'h11200000;
      23314: inst = 32'hd205b16;
      23315: inst = 32'h13e00000;
      23316: inst = 32'hfe0a9fb;
      23317: inst = 32'h5be00000;
      23318: inst = 32'h244c8000;
      23319: inst = 32'h24428800;
      23320: inst = 32'h8620000;
      23321: inst = 32'h2a0e0004;
      23322: inst = 32'h294f0003;
      23323: inst = 32'h11200000;
      23324: inst = 32'hd205b20;
      23325: inst = 32'h13e00000;
      23326: inst = 32'hfe0a9fb;
      23327: inst = 32'h5be00000;
      23328: inst = 32'h244c8000;
      23329: inst = 32'h24428800;
      23330: inst = 32'h8620000;
      23331: inst = 32'h2a0e0005;
      23332: inst = 32'h294f0003;
      23333: inst = 32'h11200000;
      23334: inst = 32'hd205b2a;
      23335: inst = 32'h13e00000;
      23336: inst = 32'hfe0a9fb;
      23337: inst = 32'h5be00000;
      23338: inst = 32'h244c8000;
      23339: inst = 32'h24428800;
      23340: inst = 32'h8620000;
      23341: inst = 32'h2a0e0006;
      23342: inst = 32'h294f0003;
      23343: inst = 32'h11200000;
      23344: inst = 32'hd205b34;
      23345: inst = 32'h13e00000;
      23346: inst = 32'hfe0a9fb;
      23347: inst = 32'h5be00000;
      23348: inst = 32'h244c8000;
      23349: inst = 32'h24428800;
      23350: inst = 32'h8620000;
      23351: inst = 32'h2a0e0007;
      23352: inst = 32'h294f0003;
      23353: inst = 32'h11200000;
      23354: inst = 32'hd205b3e;
      23355: inst = 32'h13e00000;
      23356: inst = 32'hfe0a9fb;
      23357: inst = 32'h5be00000;
      23358: inst = 32'h244c8000;
      23359: inst = 32'h24428800;
      23360: inst = 32'h8620000;
      23361: inst = 32'h2a0e0009;
      23362: inst = 32'h294f0003;
      23363: inst = 32'h11200000;
      23364: inst = 32'hd205b48;
      23365: inst = 32'h13e00000;
      23366: inst = 32'hfe0a9fb;
      23367: inst = 32'h5be00000;
      23368: inst = 32'h244c8000;
      23369: inst = 32'h24428800;
      23370: inst = 32'h8620000;
      23371: inst = 32'h2a0e0001;
      23372: inst = 32'h294f0004;
      23373: inst = 32'h11200000;
      23374: inst = 32'hd205b52;
      23375: inst = 32'h13e00000;
      23376: inst = 32'hfe0a9fb;
      23377: inst = 32'h5be00000;
      23378: inst = 32'h244c8000;
      23379: inst = 32'h24428800;
      23380: inst = 32'h8620000;
      23381: inst = 32'h2a0e0002;
      23382: inst = 32'h294f0004;
      23383: inst = 32'h11200000;
      23384: inst = 32'hd205b5c;
      23385: inst = 32'h13e00000;
      23386: inst = 32'hfe0a9fb;
      23387: inst = 32'h5be00000;
      23388: inst = 32'h244c8000;
      23389: inst = 32'h24428800;
      23390: inst = 32'h8620000;
      23391: inst = 32'h2a0e0003;
      23392: inst = 32'h294f0004;
      23393: inst = 32'h11200000;
      23394: inst = 32'hd205b66;
      23395: inst = 32'h13e00000;
      23396: inst = 32'hfe0a9fb;
      23397: inst = 32'h5be00000;
      23398: inst = 32'h244c8000;
      23399: inst = 32'h24428800;
      23400: inst = 32'h8620000;
      23401: inst = 32'h2a0e0004;
      23402: inst = 32'h294f0004;
      23403: inst = 32'h11200000;
      23404: inst = 32'hd205b70;
      23405: inst = 32'h13e00000;
      23406: inst = 32'hfe0a9fb;
      23407: inst = 32'h5be00000;
      23408: inst = 32'h244c8000;
      23409: inst = 32'h24428800;
      23410: inst = 32'h8620000;
      23411: inst = 32'h2a0e0005;
      23412: inst = 32'h294f0004;
      23413: inst = 32'h11200000;
      23414: inst = 32'hd205b7a;
      23415: inst = 32'h13e00000;
      23416: inst = 32'hfe0a9fb;
      23417: inst = 32'h5be00000;
      23418: inst = 32'h244c8000;
      23419: inst = 32'h24428800;
      23420: inst = 32'h8620000;
      23421: inst = 32'h2a0e0006;
      23422: inst = 32'h294f0004;
      23423: inst = 32'h11200000;
      23424: inst = 32'hd205b84;
      23425: inst = 32'h13e00000;
      23426: inst = 32'hfe0a9fb;
      23427: inst = 32'h5be00000;
      23428: inst = 32'h244c8000;
      23429: inst = 32'h24428800;
      23430: inst = 32'h8620000;
      23431: inst = 32'h2a0e0007;
      23432: inst = 32'h294f0004;
      23433: inst = 32'h11200000;
      23434: inst = 32'hd205b8e;
      23435: inst = 32'h13e00000;
      23436: inst = 32'hfe0a9fb;
      23437: inst = 32'h5be00000;
      23438: inst = 32'h244c8000;
      23439: inst = 32'h24428800;
      23440: inst = 32'h8620000;
      23441: inst = 32'h2a0e0009;
      23442: inst = 32'h294f0004;
      23443: inst = 32'h11200000;
      23444: inst = 32'hd205b98;
      23445: inst = 32'h13e00000;
      23446: inst = 32'hfe0a9fb;
      23447: inst = 32'h5be00000;
      23448: inst = 32'h244c8000;
      23449: inst = 32'h24428800;
      23450: inst = 32'h8620000;
      23451: inst = 32'h2a0e0003;
      23452: inst = 32'h294f0005;
      23453: inst = 32'h11200000;
      23454: inst = 32'hd205ba2;
      23455: inst = 32'h13e00000;
      23456: inst = 32'hfe0a9fb;
      23457: inst = 32'h5be00000;
      23458: inst = 32'h244c8000;
      23459: inst = 32'h24428800;
      23460: inst = 32'h8620000;
      23461: inst = 32'h2a0e0004;
      23462: inst = 32'h294f0005;
      23463: inst = 32'h11200000;
      23464: inst = 32'hd205bac;
      23465: inst = 32'h13e00000;
      23466: inst = 32'hfe0a9fb;
      23467: inst = 32'h5be00000;
      23468: inst = 32'h244c8000;
      23469: inst = 32'h24428800;
      23470: inst = 32'h8620000;
      23471: inst = 32'h2a0e0005;
      23472: inst = 32'h294f0005;
      23473: inst = 32'h11200000;
      23474: inst = 32'hd205bb6;
      23475: inst = 32'h13e00000;
      23476: inst = 32'hfe0a9fb;
      23477: inst = 32'h5be00000;
      23478: inst = 32'h244c8000;
      23479: inst = 32'h24428800;
      23480: inst = 32'h8620000;
      23481: inst = 32'h2a0e0006;
      23482: inst = 32'h294f0005;
      23483: inst = 32'h11200000;
      23484: inst = 32'hd205bc0;
      23485: inst = 32'h13e00000;
      23486: inst = 32'hfe0a9fb;
      23487: inst = 32'h5be00000;
      23488: inst = 32'h244c8000;
      23489: inst = 32'h24428800;
      23490: inst = 32'h8620000;
      23491: inst = 32'h2a0e0007;
      23492: inst = 32'h294f0005;
      23493: inst = 32'h11200000;
      23494: inst = 32'hd205bca;
      23495: inst = 32'h13e00000;
      23496: inst = 32'hfe0a9fb;
      23497: inst = 32'h5be00000;
      23498: inst = 32'h244c8000;
      23499: inst = 32'h24428800;
      23500: inst = 32'h8620000;
      23501: inst = 32'h2a0e0008;
      23502: inst = 32'h294f0005;
      23503: inst = 32'h11200000;
      23504: inst = 32'hd205bd4;
      23505: inst = 32'h13e00000;
      23506: inst = 32'hfe0a9fb;
      23507: inst = 32'h5be00000;
      23508: inst = 32'h244c8000;
      23509: inst = 32'h24428800;
      23510: inst = 32'h8620000;
      23511: inst = 32'h2a0e0009;
      23512: inst = 32'h294f0005;
      23513: inst = 32'h11200000;
      23514: inst = 32'hd205bde;
      23515: inst = 32'h13e00000;
      23516: inst = 32'hfe0a9fb;
      23517: inst = 32'h5be00000;
      23518: inst = 32'h244c8000;
      23519: inst = 32'h24428800;
      23520: inst = 32'h8620000;
      23521: inst = 32'h2a0e0003;
      23522: inst = 32'h294f0006;
      23523: inst = 32'h11200000;
      23524: inst = 32'hd205be8;
      23525: inst = 32'h13e00000;
      23526: inst = 32'hfe0a9fb;
      23527: inst = 32'h5be00000;
      23528: inst = 32'h244c8000;
      23529: inst = 32'h24428800;
      23530: inst = 32'h8620000;
      23531: inst = 32'h2a0e0004;
      23532: inst = 32'h294f0006;
      23533: inst = 32'h11200000;
      23534: inst = 32'hd205bf2;
      23535: inst = 32'h13e00000;
      23536: inst = 32'hfe0a9fb;
      23537: inst = 32'h5be00000;
      23538: inst = 32'h244c8000;
      23539: inst = 32'h24428800;
      23540: inst = 32'h8620000;
      23541: inst = 32'h2a0e0005;
      23542: inst = 32'h294f0006;
      23543: inst = 32'h11200000;
      23544: inst = 32'hd205bfc;
      23545: inst = 32'h13e00000;
      23546: inst = 32'hfe0a9fb;
      23547: inst = 32'h5be00000;
      23548: inst = 32'h244c8000;
      23549: inst = 32'h24428800;
      23550: inst = 32'h8620000;
      23551: inst = 32'h2a0e0006;
      23552: inst = 32'h294f0006;
      23553: inst = 32'h11200000;
      23554: inst = 32'hd205c06;
      23555: inst = 32'h13e00000;
      23556: inst = 32'hfe0a9fb;
      23557: inst = 32'h5be00000;
      23558: inst = 32'h244c8000;
      23559: inst = 32'h24428800;
      23560: inst = 32'h8620000;
      23561: inst = 32'h2a0e0007;
      23562: inst = 32'h294f0006;
      23563: inst = 32'h11200000;
      23564: inst = 32'hd205c10;
      23565: inst = 32'h13e00000;
      23566: inst = 32'hfe0a9fb;
      23567: inst = 32'h5be00000;
      23568: inst = 32'h244c8000;
      23569: inst = 32'h24428800;
      23570: inst = 32'h8620000;
      23571: inst = 32'h2a0e0008;
      23572: inst = 32'h294f0006;
      23573: inst = 32'h11200000;
      23574: inst = 32'hd205c1a;
      23575: inst = 32'h13e00000;
      23576: inst = 32'hfe0a9fb;
      23577: inst = 32'h5be00000;
      23578: inst = 32'h244c8000;
      23579: inst = 32'h24428800;
      23580: inst = 32'h8620000;
      23581: inst = 32'h2a0e0009;
      23582: inst = 32'h294f0006;
      23583: inst = 32'h11200000;
      23584: inst = 32'hd205c24;
      23585: inst = 32'h13e00000;
      23586: inst = 32'hfe0a9fb;
      23587: inst = 32'h5be00000;
      23588: inst = 32'h244c8000;
      23589: inst = 32'h24428800;
      23590: inst = 32'h8620000;
      23591: inst = 32'h2a0e0004;
      23592: inst = 32'h294f0008;
      23593: inst = 32'h11200000;
      23594: inst = 32'hd205c2e;
      23595: inst = 32'h13e00000;
      23596: inst = 32'hfe0a9fb;
      23597: inst = 32'h5be00000;
      23598: inst = 32'h244c8000;
      23599: inst = 32'h24428800;
      23600: inst = 32'h8620000;
      23601: inst = 32'h2a0e0008;
      23602: inst = 32'h294f0008;
      23603: inst = 32'h11200000;
      23604: inst = 32'hd205c38;
      23605: inst = 32'h13e00000;
      23606: inst = 32'hfe0a9fb;
      23607: inst = 32'h5be00000;
      23608: inst = 32'h244c8000;
      23609: inst = 32'h24428800;
      23610: inst = 32'h8620000;
      23611: inst = 32'h2a0e0004;
      23612: inst = 32'h294f0009;
      23613: inst = 32'h11200000;
      23614: inst = 32'hd205c42;
      23615: inst = 32'h13e00000;
      23616: inst = 32'hfe0a9fb;
      23617: inst = 32'h5be00000;
      23618: inst = 32'h244c8000;
      23619: inst = 32'h24428800;
      23620: inst = 32'h8620000;
      23621: inst = 32'hc607841;
      23622: inst = 32'h2a0e0002;
      23623: inst = 32'h294f0007;
      23624: inst = 32'h11200000;
      23625: inst = 32'hd205c4d;
      23626: inst = 32'h13e00000;
      23627: inst = 32'hfe0a9fb;
      23628: inst = 32'h5be00000;
      23629: inst = 32'h244c8000;
      23630: inst = 32'h24428800;
      23631: inst = 32'h8620000;
      23632: inst = 32'h2a0e0002;
      23633: inst = 32'h294f0008;
      23634: inst = 32'h11200000;
      23635: inst = 32'hd205c57;
      23636: inst = 32'h13e00000;
      23637: inst = 32'hfe0a9fb;
      23638: inst = 32'h5be00000;
      23639: inst = 32'h244c8000;
      23640: inst = 32'h24428800;
      23641: inst = 32'h8620000;
      23642: inst = 32'hc60a000;
      23643: inst = 32'h2a0e0003;
      23644: inst = 32'h294f0007;
      23645: inst = 32'h11200000;
      23646: inst = 32'hd205c62;
      23647: inst = 32'h13e00000;
      23648: inst = 32'hfe0a9fb;
      23649: inst = 32'h5be00000;
      23650: inst = 32'h244c8000;
      23651: inst = 32'h24428800;
      23652: inst = 32'h8620000;
      23653: inst = 32'h2a0e0004;
      23654: inst = 32'h294f0007;
      23655: inst = 32'h11200000;
      23656: inst = 32'hd205c6c;
      23657: inst = 32'h13e00000;
      23658: inst = 32'hfe0a9fb;
      23659: inst = 32'h5be00000;
      23660: inst = 32'h244c8000;
      23661: inst = 32'h24428800;
      23662: inst = 32'h8620000;
      23663: inst = 32'h2a0e0005;
      23664: inst = 32'h294f0007;
      23665: inst = 32'h11200000;
      23666: inst = 32'hd205c76;
      23667: inst = 32'h13e00000;
      23668: inst = 32'hfe0a9fb;
      23669: inst = 32'h5be00000;
      23670: inst = 32'h244c8000;
      23671: inst = 32'h24428800;
      23672: inst = 32'h8620000;
      23673: inst = 32'h2a0e0006;
      23674: inst = 32'h294f0007;
      23675: inst = 32'h11200000;
      23676: inst = 32'hd205c80;
      23677: inst = 32'h13e00000;
      23678: inst = 32'hfe0a9fb;
      23679: inst = 32'h5be00000;
      23680: inst = 32'h244c8000;
      23681: inst = 32'h24428800;
      23682: inst = 32'h8620000;
      23683: inst = 32'h2a0e0007;
      23684: inst = 32'h294f0007;
      23685: inst = 32'h11200000;
      23686: inst = 32'hd205c8a;
      23687: inst = 32'h13e00000;
      23688: inst = 32'hfe0a9fb;
      23689: inst = 32'h5be00000;
      23690: inst = 32'h244c8000;
      23691: inst = 32'h24428800;
      23692: inst = 32'h8620000;
      23693: inst = 32'h2a0e0003;
      23694: inst = 32'h294f0008;
      23695: inst = 32'h11200000;
      23696: inst = 32'hd205c94;
      23697: inst = 32'h13e00000;
      23698: inst = 32'hfe0a9fb;
      23699: inst = 32'h5be00000;
      23700: inst = 32'h244c8000;
      23701: inst = 32'h24428800;
      23702: inst = 32'h8620000;
      23703: inst = 32'h2a0e0005;
      23704: inst = 32'h294f0008;
      23705: inst = 32'h11200000;
      23706: inst = 32'hd205c9e;
      23707: inst = 32'h13e00000;
      23708: inst = 32'hfe0a9fb;
      23709: inst = 32'h5be00000;
      23710: inst = 32'h244c8000;
      23711: inst = 32'h24428800;
      23712: inst = 32'h8620000;
      23713: inst = 32'h2a0e0006;
      23714: inst = 32'h294f0008;
      23715: inst = 32'h11200000;
      23716: inst = 32'hd205ca8;
      23717: inst = 32'h13e00000;
      23718: inst = 32'hfe0a9fb;
      23719: inst = 32'h5be00000;
      23720: inst = 32'h244c8000;
      23721: inst = 32'h24428800;
      23722: inst = 32'h8620000;
      23723: inst = 32'h2a0e0007;
      23724: inst = 32'h294f0008;
      23725: inst = 32'h11200000;
      23726: inst = 32'hd205cb2;
      23727: inst = 32'h13e00000;
      23728: inst = 32'hfe0a9fb;
      23729: inst = 32'h5be00000;
      23730: inst = 32'h244c8000;
      23731: inst = 32'h24428800;
      23732: inst = 32'h8620000;
      23733: inst = 32'h2a0e0002;
      23734: inst = 32'h294f0009;
      23735: inst = 32'h11200000;
      23736: inst = 32'hd205cbc;
      23737: inst = 32'h13e00000;
      23738: inst = 32'hfe0a9fb;
      23739: inst = 32'h5be00000;
      23740: inst = 32'h244c8000;
      23741: inst = 32'h24428800;
      23742: inst = 32'h8620000;
      23743: inst = 32'h2a0e0003;
      23744: inst = 32'h294f0009;
      23745: inst = 32'h11200000;
      23746: inst = 32'hd205cc6;
      23747: inst = 32'h13e00000;
      23748: inst = 32'hfe0a9fb;
      23749: inst = 32'h5be00000;
      23750: inst = 32'h244c8000;
      23751: inst = 32'h24428800;
      23752: inst = 32'h8620000;
      23753: inst = 32'h2a0e0005;
      23754: inst = 32'h294f0009;
      23755: inst = 32'h11200000;
      23756: inst = 32'hd205cd0;
      23757: inst = 32'h13e00000;
      23758: inst = 32'hfe0a9fb;
      23759: inst = 32'h5be00000;
      23760: inst = 32'h244c8000;
      23761: inst = 32'h24428800;
      23762: inst = 32'h8620000;
      23763: inst = 32'h2a0e0006;
      23764: inst = 32'h294f0009;
      23765: inst = 32'h11200000;
      23766: inst = 32'hd205cda;
      23767: inst = 32'h13e00000;
      23768: inst = 32'hfe0a9fb;
      23769: inst = 32'h5be00000;
      23770: inst = 32'h244c8000;
      23771: inst = 32'h24428800;
      23772: inst = 32'h8620000;
      23773: inst = 32'h2a0e0007;
      23774: inst = 32'h294f0009;
      23775: inst = 32'h11200000;
      23776: inst = 32'hd205ce4;
      23777: inst = 32'h13e00000;
      23778: inst = 32'hfe0a9fb;
      23779: inst = 32'h5be00000;
      23780: inst = 32'h244c8000;
      23781: inst = 32'h24428800;
      23782: inst = 32'h8620000;
      23783: inst = 32'hc6010ac;
      23784: inst = 32'h2a0e0002;
      23785: inst = 32'h294f000a;
      23786: inst = 32'h11200000;
      23787: inst = 32'hd205cef;
      23788: inst = 32'h13e00000;
      23789: inst = 32'hfe0a9fb;
      23790: inst = 32'h5be00000;
      23791: inst = 32'h244c8000;
      23792: inst = 32'h24428800;
      23793: inst = 32'h8620000;
      23794: inst = 32'h2a0e0003;
      23795: inst = 32'h294f000a;
      23796: inst = 32'h11200000;
      23797: inst = 32'hd205cf9;
      23798: inst = 32'h13e00000;
      23799: inst = 32'hfe0a9fb;
      23800: inst = 32'h5be00000;
      23801: inst = 32'h244c8000;
      23802: inst = 32'h24428800;
      23803: inst = 32'h8620000;
      23804: inst = 32'h2a0e0004;
      23805: inst = 32'h294f000a;
      23806: inst = 32'h11200000;
      23807: inst = 32'hd205d03;
      23808: inst = 32'h13e00000;
      23809: inst = 32'hfe0a9fb;
      23810: inst = 32'h5be00000;
      23811: inst = 32'h244c8000;
      23812: inst = 32'h24428800;
      23813: inst = 32'h8620000;
      23814: inst = 32'h2a0e0005;
      23815: inst = 32'h294f000a;
      23816: inst = 32'h11200000;
      23817: inst = 32'hd205d0d;
      23818: inst = 32'h13e00000;
      23819: inst = 32'hfe0a9fb;
      23820: inst = 32'h5be00000;
      23821: inst = 32'h244c8000;
      23822: inst = 32'h24428800;
      23823: inst = 32'h8620000;
      23824: inst = 32'h2a0e0006;
      23825: inst = 32'h294f000a;
      23826: inst = 32'h11200000;
      23827: inst = 32'hd205d17;
      23828: inst = 32'h13e00000;
      23829: inst = 32'hfe0a9fb;
      23830: inst = 32'h5be00000;
      23831: inst = 32'h244c8000;
      23832: inst = 32'h24428800;
      23833: inst = 32'h8620000;
      23834: inst = 32'h2a0e0007;
      23835: inst = 32'h294f000a;
      23836: inst = 32'h11200000;
      23837: inst = 32'hd205d21;
      23838: inst = 32'h13e00000;
      23839: inst = 32'hfe0a9fb;
      23840: inst = 32'h5be00000;
      23841: inst = 32'h244c8000;
      23842: inst = 32'h24428800;
      23843: inst = 32'h8620000;
      23844: inst = 32'h13e00000;
      23845: inst = 32'hfe05d2b;
      23846: inst = 32'h20200003;
      23847: inst = 32'h5be00000;
      23848: inst = 32'h13e00000;
      23849: inst = 32'hfe06108;
      23850: inst = 32'h5be00000;
      23851: inst = 32'h13e00000;
      23852: inst = 32'hfe06108;
      23853: inst = 32'h5be00000;
      23854: inst = 32'hc6018c3;
      23855: inst = 32'h2a0e000a;
      23856: inst = 32'h294f0000;
      23857: inst = 32'h11200000;
      23858: inst = 32'hd205d36;
      23859: inst = 32'h13e00000;
      23860: inst = 32'hfe0a9fb;
      23861: inst = 32'h5be00000;
      23862: inst = 32'h244c8000;
      23863: inst = 32'h24428800;
      23864: inst = 32'h8620000;
      23865: inst = 32'h2a0e0009;
      23866: inst = 32'h294f0000;
      23867: inst = 32'h11200000;
      23868: inst = 32'hd205d40;
      23869: inst = 32'h13e00000;
      23870: inst = 32'hfe0a9fb;
      23871: inst = 32'h5be00000;
      23872: inst = 32'h244c8000;
      23873: inst = 32'h24428800;
      23874: inst = 32'h8620000;
      23875: inst = 32'h2a0e0008;
      23876: inst = 32'h294f0000;
      23877: inst = 32'h11200000;
      23878: inst = 32'hd205d4a;
      23879: inst = 32'h13e00000;
      23880: inst = 32'hfe0a9fb;
      23881: inst = 32'h5be00000;
      23882: inst = 32'h244c8000;
      23883: inst = 32'h24428800;
      23884: inst = 32'h8620000;
      23885: inst = 32'h2a0e0007;
      23886: inst = 32'h294f0000;
      23887: inst = 32'h11200000;
      23888: inst = 32'hd205d54;
      23889: inst = 32'h13e00000;
      23890: inst = 32'hfe0a9fb;
      23891: inst = 32'h5be00000;
      23892: inst = 32'h244c8000;
      23893: inst = 32'h24428800;
      23894: inst = 32'h8620000;
      23895: inst = 32'h2a0e0006;
      23896: inst = 32'h294f0000;
      23897: inst = 32'h11200000;
      23898: inst = 32'hd205d5e;
      23899: inst = 32'h13e00000;
      23900: inst = 32'hfe0a9fb;
      23901: inst = 32'h5be00000;
      23902: inst = 32'h244c8000;
      23903: inst = 32'h24428800;
      23904: inst = 32'h8620000;
      23905: inst = 32'h2a0e0005;
      23906: inst = 32'h294f0000;
      23907: inst = 32'h11200000;
      23908: inst = 32'hd205d68;
      23909: inst = 32'h13e00000;
      23910: inst = 32'hfe0a9fb;
      23911: inst = 32'h5be00000;
      23912: inst = 32'h244c8000;
      23913: inst = 32'h24428800;
      23914: inst = 32'h8620000;
      23915: inst = 32'h2a0e0004;
      23916: inst = 32'h294f0000;
      23917: inst = 32'h11200000;
      23918: inst = 32'hd205d72;
      23919: inst = 32'h13e00000;
      23920: inst = 32'hfe0a9fb;
      23921: inst = 32'h5be00000;
      23922: inst = 32'h244c8000;
      23923: inst = 32'h24428800;
      23924: inst = 32'h8620000;
      23925: inst = 32'h2a0e0003;
      23926: inst = 32'h294f0000;
      23927: inst = 32'h11200000;
      23928: inst = 32'hd205d7c;
      23929: inst = 32'h13e00000;
      23930: inst = 32'hfe0a9fb;
      23931: inst = 32'h5be00000;
      23932: inst = 32'h244c8000;
      23933: inst = 32'h24428800;
      23934: inst = 32'h8620000;
      23935: inst = 32'h2a0e0002;
      23936: inst = 32'h294f0000;
      23937: inst = 32'h11200000;
      23938: inst = 32'hd205d86;
      23939: inst = 32'h13e00000;
      23940: inst = 32'hfe0a9fb;
      23941: inst = 32'h5be00000;
      23942: inst = 32'h244c8000;
      23943: inst = 32'h24428800;
      23944: inst = 32'h8620000;
      23945: inst = 32'h2a0e0001;
      23946: inst = 32'h294f0000;
      23947: inst = 32'h11200000;
      23948: inst = 32'hd205d90;
      23949: inst = 32'h13e00000;
      23950: inst = 32'hfe0a9fb;
      23951: inst = 32'h5be00000;
      23952: inst = 32'h244c8000;
      23953: inst = 32'h24428800;
      23954: inst = 32'h8620000;
      23955: inst = 32'h2a0e000a;
      23956: inst = 32'h294f0001;
      23957: inst = 32'h11200000;
      23958: inst = 32'hd205d9a;
      23959: inst = 32'h13e00000;
      23960: inst = 32'hfe0a9fb;
      23961: inst = 32'h5be00000;
      23962: inst = 32'h244c8000;
      23963: inst = 32'h24428800;
      23964: inst = 32'h8620000;
      23965: inst = 32'h2a0e0009;
      23966: inst = 32'h294f0001;
      23967: inst = 32'h11200000;
      23968: inst = 32'hd205da4;
      23969: inst = 32'h13e00000;
      23970: inst = 32'hfe0a9fb;
      23971: inst = 32'h5be00000;
      23972: inst = 32'h244c8000;
      23973: inst = 32'h24428800;
      23974: inst = 32'h8620000;
      23975: inst = 32'h2a0e0008;
      23976: inst = 32'h294f0001;
      23977: inst = 32'h11200000;
      23978: inst = 32'hd205dae;
      23979: inst = 32'h13e00000;
      23980: inst = 32'hfe0a9fb;
      23981: inst = 32'h5be00000;
      23982: inst = 32'h244c8000;
      23983: inst = 32'h24428800;
      23984: inst = 32'h8620000;
      23985: inst = 32'h2a0e0007;
      23986: inst = 32'h294f0001;
      23987: inst = 32'h11200000;
      23988: inst = 32'hd205db8;
      23989: inst = 32'h13e00000;
      23990: inst = 32'hfe0a9fb;
      23991: inst = 32'h5be00000;
      23992: inst = 32'h244c8000;
      23993: inst = 32'h24428800;
      23994: inst = 32'h8620000;
      23995: inst = 32'h2a0e0006;
      23996: inst = 32'h294f0001;
      23997: inst = 32'h11200000;
      23998: inst = 32'hd205dc2;
      23999: inst = 32'h13e00000;
      24000: inst = 32'hfe0a9fb;
      24001: inst = 32'h5be00000;
      24002: inst = 32'h244c8000;
      24003: inst = 32'h24428800;
      24004: inst = 32'h8620000;
      24005: inst = 32'h2a0e0005;
      24006: inst = 32'h294f0001;
      24007: inst = 32'h11200000;
      24008: inst = 32'hd205dcc;
      24009: inst = 32'h13e00000;
      24010: inst = 32'hfe0a9fb;
      24011: inst = 32'h5be00000;
      24012: inst = 32'h244c8000;
      24013: inst = 32'h24428800;
      24014: inst = 32'h8620000;
      24015: inst = 32'h2a0e0004;
      24016: inst = 32'h294f0001;
      24017: inst = 32'h11200000;
      24018: inst = 32'hd205dd6;
      24019: inst = 32'h13e00000;
      24020: inst = 32'hfe0a9fb;
      24021: inst = 32'h5be00000;
      24022: inst = 32'h244c8000;
      24023: inst = 32'h24428800;
      24024: inst = 32'h8620000;
      24025: inst = 32'h2a0e0003;
      24026: inst = 32'h294f0001;
      24027: inst = 32'h11200000;
      24028: inst = 32'hd205de0;
      24029: inst = 32'h13e00000;
      24030: inst = 32'hfe0a9fb;
      24031: inst = 32'h5be00000;
      24032: inst = 32'h244c8000;
      24033: inst = 32'h24428800;
      24034: inst = 32'h8620000;
      24035: inst = 32'h2a0e0002;
      24036: inst = 32'h294f0001;
      24037: inst = 32'h11200000;
      24038: inst = 32'hd205dea;
      24039: inst = 32'h13e00000;
      24040: inst = 32'hfe0a9fb;
      24041: inst = 32'h5be00000;
      24042: inst = 32'h244c8000;
      24043: inst = 32'h24428800;
      24044: inst = 32'h8620000;
      24045: inst = 32'h2a0e0001;
      24046: inst = 32'h294f0001;
      24047: inst = 32'h11200000;
      24048: inst = 32'hd205df4;
      24049: inst = 32'h13e00000;
      24050: inst = 32'hfe0a9fb;
      24051: inst = 32'h5be00000;
      24052: inst = 32'h244c8000;
      24053: inst = 32'h24428800;
      24054: inst = 32'h8620000;
      24055: inst = 32'h2a0e000a;
      24056: inst = 32'h294f0002;
      24057: inst = 32'h11200000;
      24058: inst = 32'hd205dfe;
      24059: inst = 32'h13e00000;
      24060: inst = 32'hfe0a9fb;
      24061: inst = 32'h5be00000;
      24062: inst = 32'h244c8000;
      24063: inst = 32'h24428800;
      24064: inst = 32'h8620000;
      24065: inst = 32'h2a0e0009;
      24066: inst = 32'h294f0002;
      24067: inst = 32'h11200000;
      24068: inst = 32'hd205e08;
      24069: inst = 32'h13e00000;
      24070: inst = 32'hfe0a9fb;
      24071: inst = 32'h5be00000;
      24072: inst = 32'h244c8000;
      24073: inst = 32'h24428800;
      24074: inst = 32'h8620000;
      24075: inst = 32'h2a0e000a;
      24076: inst = 32'h294f0003;
      24077: inst = 32'h11200000;
      24078: inst = 32'hd205e12;
      24079: inst = 32'h13e00000;
      24080: inst = 32'hfe0a9fb;
      24081: inst = 32'h5be00000;
      24082: inst = 32'h244c8000;
      24083: inst = 32'h24428800;
      24084: inst = 32'h8620000;
      24085: inst = 32'h2a0e0002;
      24086: inst = 32'h294f0003;
      24087: inst = 32'h11200000;
      24088: inst = 32'hd205e1c;
      24089: inst = 32'h13e00000;
      24090: inst = 32'hfe0a9fb;
      24091: inst = 32'h5be00000;
      24092: inst = 32'h244c8000;
      24093: inst = 32'h24428800;
      24094: inst = 32'h8620000;
      24095: inst = 32'h2a0e000a;
      24096: inst = 32'h294f0004;
      24097: inst = 32'h11200000;
      24098: inst = 32'hd205e26;
      24099: inst = 32'h13e00000;
      24100: inst = 32'hfe0a9fb;
      24101: inst = 32'h5be00000;
      24102: inst = 32'h244c8000;
      24103: inst = 32'h24428800;
      24104: inst = 32'h8620000;
      24105: inst = 32'h2a0e0002;
      24106: inst = 32'h294f0004;
      24107: inst = 32'h11200000;
      24108: inst = 32'hd205e30;
      24109: inst = 32'h13e00000;
      24110: inst = 32'hfe0a9fb;
      24111: inst = 32'h5be00000;
      24112: inst = 32'h244c8000;
      24113: inst = 32'h24428800;
      24114: inst = 32'h8620000;
      24115: inst = 32'h2a0e000a;
      24116: inst = 32'h294f0005;
      24117: inst = 32'h11200000;
      24118: inst = 32'hd205e3a;
      24119: inst = 32'h13e00000;
      24120: inst = 32'hfe0a9fb;
      24121: inst = 32'h5be00000;
      24122: inst = 32'h244c8000;
      24123: inst = 32'h24428800;
      24124: inst = 32'h8620000;
      24125: inst = 32'h2a0e0009;
      24126: inst = 32'h294f0005;
      24127: inst = 32'h11200000;
      24128: inst = 32'hd205e44;
      24129: inst = 32'h13e00000;
      24130: inst = 32'hfe0a9fb;
      24131: inst = 32'h5be00000;
      24132: inst = 32'h244c8000;
      24133: inst = 32'h24428800;
      24134: inst = 32'h8620000;
      24135: inst = 32'h2a0e000a;
      24136: inst = 32'h294f0006;
      24137: inst = 32'h11200000;
      24138: inst = 32'hd205e4e;
      24139: inst = 32'h13e00000;
      24140: inst = 32'hfe0a9fb;
      24141: inst = 32'h5be00000;
      24142: inst = 32'h244c8000;
      24143: inst = 32'h24428800;
      24144: inst = 32'h8620000;
      24145: inst = 32'h2a0e0009;
      24146: inst = 32'h294f0006;
      24147: inst = 32'h11200000;
      24148: inst = 32'hd205e58;
      24149: inst = 32'h13e00000;
      24150: inst = 32'hfe0a9fb;
      24151: inst = 32'h5be00000;
      24152: inst = 32'h244c8000;
      24153: inst = 32'h24428800;
      24154: inst = 32'h8620000;
      24155: inst = 32'hc60d42c;
      24156: inst = 32'h2a0e0008;
      24157: inst = 32'h294f0002;
      24158: inst = 32'h11200000;
      24159: inst = 32'hd205e63;
      24160: inst = 32'h13e00000;
      24161: inst = 32'hfe0a9fb;
      24162: inst = 32'h5be00000;
      24163: inst = 32'h244c8000;
      24164: inst = 32'h24428800;
      24165: inst = 32'h8620000;
      24166: inst = 32'h2a0e0007;
      24167: inst = 32'h294f0002;
      24168: inst = 32'h11200000;
      24169: inst = 32'hd205e6d;
      24170: inst = 32'h13e00000;
      24171: inst = 32'hfe0a9fb;
      24172: inst = 32'h5be00000;
      24173: inst = 32'h244c8000;
      24174: inst = 32'h24428800;
      24175: inst = 32'h8620000;
      24176: inst = 32'h2a0e0006;
      24177: inst = 32'h294f0002;
      24178: inst = 32'h11200000;
      24179: inst = 32'hd205e77;
      24180: inst = 32'h13e00000;
      24181: inst = 32'hfe0a9fb;
      24182: inst = 32'h5be00000;
      24183: inst = 32'h244c8000;
      24184: inst = 32'h24428800;
      24185: inst = 32'h8620000;
      24186: inst = 32'h2a0e0005;
      24187: inst = 32'h294f0002;
      24188: inst = 32'h11200000;
      24189: inst = 32'hd205e81;
      24190: inst = 32'h13e00000;
      24191: inst = 32'hfe0a9fb;
      24192: inst = 32'h5be00000;
      24193: inst = 32'h244c8000;
      24194: inst = 32'h24428800;
      24195: inst = 32'h8620000;
      24196: inst = 32'h2a0e0004;
      24197: inst = 32'h294f0002;
      24198: inst = 32'h11200000;
      24199: inst = 32'hd205e8b;
      24200: inst = 32'h13e00000;
      24201: inst = 32'hfe0a9fb;
      24202: inst = 32'h5be00000;
      24203: inst = 32'h244c8000;
      24204: inst = 32'h24428800;
      24205: inst = 32'h8620000;
      24206: inst = 32'h2a0e0003;
      24207: inst = 32'h294f0002;
      24208: inst = 32'h11200000;
      24209: inst = 32'hd205e95;
      24210: inst = 32'h13e00000;
      24211: inst = 32'hfe0a9fb;
      24212: inst = 32'h5be00000;
      24213: inst = 32'h244c8000;
      24214: inst = 32'h24428800;
      24215: inst = 32'h8620000;
      24216: inst = 32'h2a0e0002;
      24217: inst = 32'h294f0002;
      24218: inst = 32'h11200000;
      24219: inst = 32'hd205e9f;
      24220: inst = 32'h13e00000;
      24221: inst = 32'hfe0a9fb;
      24222: inst = 32'h5be00000;
      24223: inst = 32'h244c8000;
      24224: inst = 32'h24428800;
      24225: inst = 32'h8620000;
      24226: inst = 32'h2a0e0001;
      24227: inst = 32'h294f0002;
      24228: inst = 32'h11200000;
      24229: inst = 32'hd205ea9;
      24230: inst = 32'h13e00000;
      24231: inst = 32'hfe0a9fb;
      24232: inst = 32'h5be00000;
      24233: inst = 32'h244c8000;
      24234: inst = 32'h24428800;
      24235: inst = 32'h8620000;
      24236: inst = 32'h2a0e0008;
      24237: inst = 32'h294f0005;
      24238: inst = 32'h11200000;
      24239: inst = 32'hd205eb3;
      24240: inst = 32'h13e00000;
      24241: inst = 32'hfe0a9fb;
      24242: inst = 32'h5be00000;
      24243: inst = 32'h244c8000;
      24244: inst = 32'h24428800;
      24245: inst = 32'h8620000;
      24246: inst = 32'h2a0e0008;
      24247: inst = 32'h294f0006;
      24248: inst = 32'h11200000;
      24249: inst = 32'hd205ebd;
      24250: inst = 32'h13e00000;
      24251: inst = 32'hfe0a9fb;
      24252: inst = 32'h5be00000;
      24253: inst = 32'h244c8000;
      24254: inst = 32'h24428800;
      24255: inst = 32'h8620000;
      24256: inst = 32'h2a0e0007;
      24257: inst = 32'h294f000b;
      24258: inst = 32'h11200000;
      24259: inst = 32'hd205ec7;
      24260: inst = 32'h13e00000;
      24261: inst = 32'hfe0a9fb;
      24262: inst = 32'h5be00000;
      24263: inst = 32'h244c8000;
      24264: inst = 32'h24428800;
      24265: inst = 32'h8620000;
      24266: inst = 32'h2a0e0004;
      24267: inst = 32'h294f000b;
      24268: inst = 32'h11200000;
      24269: inst = 32'hd205ed1;
      24270: inst = 32'h13e00000;
      24271: inst = 32'hfe0a9fb;
      24272: inst = 32'h5be00000;
      24273: inst = 32'h244c8000;
      24274: inst = 32'h24428800;
      24275: inst = 32'h8620000;
      24276: inst = 32'hc60f4ce;
      24277: inst = 32'h2a0e0009;
      24278: inst = 32'h294f0003;
      24279: inst = 32'h11200000;
      24280: inst = 32'hd205edc;
      24281: inst = 32'h13e00000;
      24282: inst = 32'hfe0a9fb;
      24283: inst = 32'h5be00000;
      24284: inst = 32'h244c8000;
      24285: inst = 32'h24428800;
      24286: inst = 32'h8620000;
      24287: inst = 32'h2a0e0008;
      24288: inst = 32'h294f0003;
      24289: inst = 32'h11200000;
      24290: inst = 32'hd205ee6;
      24291: inst = 32'h13e00000;
      24292: inst = 32'hfe0a9fb;
      24293: inst = 32'h5be00000;
      24294: inst = 32'h244c8000;
      24295: inst = 32'h24428800;
      24296: inst = 32'h8620000;
      24297: inst = 32'h2a0e0007;
      24298: inst = 32'h294f0003;
      24299: inst = 32'h11200000;
      24300: inst = 32'hd205ef0;
      24301: inst = 32'h13e00000;
      24302: inst = 32'hfe0a9fb;
      24303: inst = 32'h5be00000;
      24304: inst = 32'h244c8000;
      24305: inst = 32'h24428800;
      24306: inst = 32'h8620000;
      24307: inst = 32'h2a0e0006;
      24308: inst = 32'h294f0003;
      24309: inst = 32'h11200000;
      24310: inst = 32'hd205efa;
      24311: inst = 32'h13e00000;
      24312: inst = 32'hfe0a9fb;
      24313: inst = 32'h5be00000;
      24314: inst = 32'h244c8000;
      24315: inst = 32'h24428800;
      24316: inst = 32'h8620000;
      24317: inst = 32'h2a0e0005;
      24318: inst = 32'h294f0003;
      24319: inst = 32'h11200000;
      24320: inst = 32'hd205f04;
      24321: inst = 32'h13e00000;
      24322: inst = 32'hfe0a9fb;
      24323: inst = 32'h5be00000;
      24324: inst = 32'h244c8000;
      24325: inst = 32'h24428800;
      24326: inst = 32'h8620000;
      24327: inst = 32'h2a0e0004;
      24328: inst = 32'h294f0003;
      24329: inst = 32'h11200000;
      24330: inst = 32'hd205f0e;
      24331: inst = 32'h13e00000;
      24332: inst = 32'hfe0a9fb;
      24333: inst = 32'h5be00000;
      24334: inst = 32'h244c8000;
      24335: inst = 32'h24428800;
      24336: inst = 32'h8620000;
      24337: inst = 32'h2a0e0003;
      24338: inst = 32'h294f0003;
      24339: inst = 32'h11200000;
      24340: inst = 32'hd205f18;
      24341: inst = 32'h13e00000;
      24342: inst = 32'hfe0a9fb;
      24343: inst = 32'h5be00000;
      24344: inst = 32'h244c8000;
      24345: inst = 32'h24428800;
      24346: inst = 32'h8620000;
      24347: inst = 32'h2a0e0001;
      24348: inst = 32'h294f0003;
      24349: inst = 32'h11200000;
      24350: inst = 32'hd205f22;
      24351: inst = 32'h13e00000;
      24352: inst = 32'hfe0a9fb;
      24353: inst = 32'h5be00000;
      24354: inst = 32'h244c8000;
      24355: inst = 32'h24428800;
      24356: inst = 32'h8620000;
      24357: inst = 32'h2a0e0009;
      24358: inst = 32'h294f0004;
      24359: inst = 32'h11200000;
      24360: inst = 32'hd205f2c;
      24361: inst = 32'h13e00000;
      24362: inst = 32'hfe0a9fb;
      24363: inst = 32'h5be00000;
      24364: inst = 32'h244c8000;
      24365: inst = 32'h24428800;
      24366: inst = 32'h8620000;
      24367: inst = 32'h2a0e0008;
      24368: inst = 32'h294f0004;
      24369: inst = 32'h11200000;
      24370: inst = 32'hd205f36;
      24371: inst = 32'h13e00000;
      24372: inst = 32'hfe0a9fb;
      24373: inst = 32'h5be00000;
      24374: inst = 32'h244c8000;
      24375: inst = 32'h24428800;
      24376: inst = 32'h8620000;
      24377: inst = 32'h2a0e0007;
      24378: inst = 32'h294f0004;
      24379: inst = 32'h11200000;
      24380: inst = 32'hd205f40;
      24381: inst = 32'h13e00000;
      24382: inst = 32'hfe0a9fb;
      24383: inst = 32'h5be00000;
      24384: inst = 32'h244c8000;
      24385: inst = 32'h24428800;
      24386: inst = 32'h8620000;
      24387: inst = 32'h2a0e0006;
      24388: inst = 32'h294f0004;
      24389: inst = 32'h11200000;
      24390: inst = 32'hd205f4a;
      24391: inst = 32'h13e00000;
      24392: inst = 32'hfe0a9fb;
      24393: inst = 32'h5be00000;
      24394: inst = 32'h244c8000;
      24395: inst = 32'h24428800;
      24396: inst = 32'h8620000;
      24397: inst = 32'h2a0e0005;
      24398: inst = 32'h294f0004;
      24399: inst = 32'h11200000;
      24400: inst = 32'hd205f54;
      24401: inst = 32'h13e00000;
      24402: inst = 32'hfe0a9fb;
      24403: inst = 32'h5be00000;
      24404: inst = 32'h244c8000;
      24405: inst = 32'h24428800;
      24406: inst = 32'h8620000;
      24407: inst = 32'h2a0e0004;
      24408: inst = 32'h294f0004;
      24409: inst = 32'h11200000;
      24410: inst = 32'hd205f5e;
      24411: inst = 32'h13e00000;
      24412: inst = 32'hfe0a9fb;
      24413: inst = 32'h5be00000;
      24414: inst = 32'h244c8000;
      24415: inst = 32'h24428800;
      24416: inst = 32'h8620000;
      24417: inst = 32'h2a0e0003;
      24418: inst = 32'h294f0004;
      24419: inst = 32'h11200000;
      24420: inst = 32'hd205f68;
      24421: inst = 32'h13e00000;
      24422: inst = 32'hfe0a9fb;
      24423: inst = 32'h5be00000;
      24424: inst = 32'h244c8000;
      24425: inst = 32'h24428800;
      24426: inst = 32'h8620000;
      24427: inst = 32'h2a0e0001;
      24428: inst = 32'h294f0004;
      24429: inst = 32'h11200000;
      24430: inst = 32'hd205f72;
      24431: inst = 32'h13e00000;
      24432: inst = 32'hfe0a9fb;
      24433: inst = 32'h5be00000;
      24434: inst = 32'h244c8000;
      24435: inst = 32'h24428800;
      24436: inst = 32'h8620000;
      24437: inst = 32'h2a0e0007;
      24438: inst = 32'h294f0005;
      24439: inst = 32'h11200000;
      24440: inst = 32'hd205f7c;
      24441: inst = 32'h13e00000;
      24442: inst = 32'hfe0a9fb;
      24443: inst = 32'h5be00000;
      24444: inst = 32'h244c8000;
      24445: inst = 32'h24428800;
      24446: inst = 32'h8620000;
      24447: inst = 32'h2a0e0006;
      24448: inst = 32'h294f0005;
      24449: inst = 32'h11200000;
      24450: inst = 32'hd205f86;
      24451: inst = 32'h13e00000;
      24452: inst = 32'hfe0a9fb;
      24453: inst = 32'h5be00000;
      24454: inst = 32'h244c8000;
      24455: inst = 32'h24428800;
      24456: inst = 32'h8620000;
      24457: inst = 32'h2a0e0005;
      24458: inst = 32'h294f0005;
      24459: inst = 32'h11200000;
      24460: inst = 32'hd205f90;
      24461: inst = 32'h13e00000;
      24462: inst = 32'hfe0a9fb;
      24463: inst = 32'h5be00000;
      24464: inst = 32'h244c8000;
      24465: inst = 32'h24428800;
      24466: inst = 32'h8620000;
      24467: inst = 32'h2a0e0004;
      24468: inst = 32'h294f0005;
      24469: inst = 32'h11200000;
      24470: inst = 32'hd205f9a;
      24471: inst = 32'h13e00000;
      24472: inst = 32'hfe0a9fb;
      24473: inst = 32'h5be00000;
      24474: inst = 32'h244c8000;
      24475: inst = 32'h24428800;
      24476: inst = 32'h8620000;
      24477: inst = 32'h2a0e0003;
      24478: inst = 32'h294f0005;
      24479: inst = 32'h11200000;
      24480: inst = 32'hd205fa4;
      24481: inst = 32'h13e00000;
      24482: inst = 32'hfe0a9fb;
      24483: inst = 32'h5be00000;
      24484: inst = 32'h244c8000;
      24485: inst = 32'h24428800;
      24486: inst = 32'h8620000;
      24487: inst = 32'h2a0e0002;
      24488: inst = 32'h294f0005;
      24489: inst = 32'h11200000;
      24490: inst = 32'hd205fae;
      24491: inst = 32'h13e00000;
      24492: inst = 32'hfe0a9fb;
      24493: inst = 32'h5be00000;
      24494: inst = 32'h244c8000;
      24495: inst = 32'h24428800;
      24496: inst = 32'h8620000;
      24497: inst = 32'h2a0e0001;
      24498: inst = 32'h294f0005;
      24499: inst = 32'h11200000;
      24500: inst = 32'hd205fb8;
      24501: inst = 32'h13e00000;
      24502: inst = 32'hfe0a9fb;
      24503: inst = 32'h5be00000;
      24504: inst = 32'h244c8000;
      24505: inst = 32'h24428800;
      24506: inst = 32'h8620000;
      24507: inst = 32'h2a0e0007;
      24508: inst = 32'h294f0006;
      24509: inst = 32'h11200000;
      24510: inst = 32'hd205fc2;
      24511: inst = 32'h13e00000;
      24512: inst = 32'hfe0a9fb;
      24513: inst = 32'h5be00000;
      24514: inst = 32'h244c8000;
      24515: inst = 32'h24428800;
      24516: inst = 32'h8620000;
      24517: inst = 32'h2a0e0006;
      24518: inst = 32'h294f0006;
      24519: inst = 32'h11200000;
      24520: inst = 32'hd205fcc;
      24521: inst = 32'h13e00000;
      24522: inst = 32'hfe0a9fb;
      24523: inst = 32'h5be00000;
      24524: inst = 32'h244c8000;
      24525: inst = 32'h24428800;
      24526: inst = 32'h8620000;
      24527: inst = 32'h2a0e0005;
      24528: inst = 32'h294f0006;
      24529: inst = 32'h11200000;
      24530: inst = 32'hd205fd6;
      24531: inst = 32'h13e00000;
      24532: inst = 32'hfe0a9fb;
      24533: inst = 32'h5be00000;
      24534: inst = 32'h244c8000;
      24535: inst = 32'h24428800;
      24536: inst = 32'h8620000;
      24537: inst = 32'h2a0e0004;
      24538: inst = 32'h294f0006;
      24539: inst = 32'h11200000;
      24540: inst = 32'hd205fe0;
      24541: inst = 32'h13e00000;
      24542: inst = 32'hfe0a9fb;
      24543: inst = 32'h5be00000;
      24544: inst = 32'h244c8000;
      24545: inst = 32'h24428800;
      24546: inst = 32'h8620000;
      24547: inst = 32'h2a0e0003;
      24548: inst = 32'h294f0006;
      24549: inst = 32'h11200000;
      24550: inst = 32'hd205fea;
      24551: inst = 32'h13e00000;
      24552: inst = 32'hfe0a9fb;
      24553: inst = 32'h5be00000;
      24554: inst = 32'h244c8000;
      24555: inst = 32'h24428800;
      24556: inst = 32'h8620000;
      24557: inst = 32'h2a0e0002;
      24558: inst = 32'h294f0006;
      24559: inst = 32'h11200000;
      24560: inst = 32'hd205ff4;
      24561: inst = 32'h13e00000;
      24562: inst = 32'hfe0a9fb;
      24563: inst = 32'h5be00000;
      24564: inst = 32'h244c8000;
      24565: inst = 32'h24428800;
      24566: inst = 32'h8620000;
      24567: inst = 32'h2a0e0001;
      24568: inst = 32'h294f0006;
      24569: inst = 32'h11200000;
      24570: inst = 32'hd205ffe;
      24571: inst = 32'h13e00000;
      24572: inst = 32'hfe0a9fb;
      24573: inst = 32'h5be00000;
      24574: inst = 32'h244c8000;
      24575: inst = 32'h24428800;
      24576: inst = 32'h8620000;
      24577: inst = 32'h2a0e0006;
      24578: inst = 32'h294f0008;
      24579: inst = 32'h11200000;
      24580: inst = 32'hd206008;
      24581: inst = 32'h13e00000;
      24582: inst = 32'hfe0a9fb;
      24583: inst = 32'h5be00000;
      24584: inst = 32'h244c8000;
      24585: inst = 32'h24428800;
      24586: inst = 32'h8620000;
      24587: inst = 32'h2a0e0002;
      24588: inst = 32'h294f0008;
      24589: inst = 32'h11200000;
      24590: inst = 32'hd206012;
      24591: inst = 32'h13e00000;
      24592: inst = 32'hfe0a9fb;
      24593: inst = 32'h5be00000;
      24594: inst = 32'h244c8000;
      24595: inst = 32'h24428800;
      24596: inst = 32'h8620000;
      24597: inst = 32'h2a0e0006;
      24598: inst = 32'h294f0009;
      24599: inst = 32'h11200000;
      24600: inst = 32'hd20601c;
      24601: inst = 32'h13e00000;
      24602: inst = 32'hfe0a9fb;
      24603: inst = 32'h5be00000;
      24604: inst = 32'h244c8000;
      24605: inst = 32'h24428800;
      24606: inst = 32'h8620000;
      24607: inst = 32'hc607841;
      24608: inst = 32'h2a0e0008;
      24609: inst = 32'h294f0007;
      24610: inst = 32'h11200000;
      24611: inst = 32'hd206027;
      24612: inst = 32'h13e00000;
      24613: inst = 32'hfe0a9fb;
      24614: inst = 32'h5be00000;
      24615: inst = 32'h244c8000;
      24616: inst = 32'h24428800;
      24617: inst = 32'h8620000;
      24618: inst = 32'h2a0e0008;
      24619: inst = 32'h294f0008;
      24620: inst = 32'h11200000;
      24621: inst = 32'hd206031;
      24622: inst = 32'h13e00000;
      24623: inst = 32'hfe0a9fb;
      24624: inst = 32'h5be00000;
      24625: inst = 32'h244c8000;
      24626: inst = 32'h24428800;
      24627: inst = 32'h8620000;
      24628: inst = 32'hc60a000;
      24629: inst = 32'h2a0e0007;
      24630: inst = 32'h294f0007;
      24631: inst = 32'h11200000;
      24632: inst = 32'hd20603c;
      24633: inst = 32'h13e00000;
      24634: inst = 32'hfe0a9fb;
      24635: inst = 32'h5be00000;
      24636: inst = 32'h244c8000;
      24637: inst = 32'h24428800;
      24638: inst = 32'h8620000;
      24639: inst = 32'h2a0e0006;
      24640: inst = 32'h294f0007;
      24641: inst = 32'h11200000;
      24642: inst = 32'hd206046;
      24643: inst = 32'h13e00000;
      24644: inst = 32'hfe0a9fb;
      24645: inst = 32'h5be00000;
      24646: inst = 32'h244c8000;
      24647: inst = 32'h24428800;
      24648: inst = 32'h8620000;
      24649: inst = 32'h2a0e0005;
      24650: inst = 32'h294f0007;
      24651: inst = 32'h11200000;
      24652: inst = 32'hd206050;
      24653: inst = 32'h13e00000;
      24654: inst = 32'hfe0a9fb;
      24655: inst = 32'h5be00000;
      24656: inst = 32'h244c8000;
      24657: inst = 32'h24428800;
      24658: inst = 32'h8620000;
      24659: inst = 32'h2a0e0004;
      24660: inst = 32'h294f0007;
      24661: inst = 32'h11200000;
      24662: inst = 32'hd20605a;
      24663: inst = 32'h13e00000;
      24664: inst = 32'hfe0a9fb;
      24665: inst = 32'h5be00000;
      24666: inst = 32'h244c8000;
      24667: inst = 32'h24428800;
      24668: inst = 32'h8620000;
      24669: inst = 32'h2a0e0003;
      24670: inst = 32'h294f0007;
      24671: inst = 32'h11200000;
      24672: inst = 32'hd206064;
      24673: inst = 32'h13e00000;
      24674: inst = 32'hfe0a9fb;
      24675: inst = 32'h5be00000;
      24676: inst = 32'h244c8000;
      24677: inst = 32'h24428800;
      24678: inst = 32'h8620000;
      24679: inst = 32'h2a0e0007;
      24680: inst = 32'h294f0008;
      24681: inst = 32'h11200000;
      24682: inst = 32'hd20606e;
      24683: inst = 32'h13e00000;
      24684: inst = 32'hfe0a9fb;
      24685: inst = 32'h5be00000;
      24686: inst = 32'h244c8000;
      24687: inst = 32'h24428800;
      24688: inst = 32'h8620000;
      24689: inst = 32'h2a0e0005;
      24690: inst = 32'h294f0008;
      24691: inst = 32'h11200000;
      24692: inst = 32'hd206078;
      24693: inst = 32'h13e00000;
      24694: inst = 32'hfe0a9fb;
      24695: inst = 32'h5be00000;
      24696: inst = 32'h244c8000;
      24697: inst = 32'h24428800;
      24698: inst = 32'h8620000;
      24699: inst = 32'h2a0e0004;
      24700: inst = 32'h294f0008;
      24701: inst = 32'h11200000;
      24702: inst = 32'hd206082;
      24703: inst = 32'h13e00000;
      24704: inst = 32'hfe0a9fb;
      24705: inst = 32'h5be00000;
      24706: inst = 32'h244c8000;
      24707: inst = 32'h24428800;
      24708: inst = 32'h8620000;
      24709: inst = 32'h2a0e0003;
      24710: inst = 32'h294f0008;
      24711: inst = 32'h11200000;
      24712: inst = 32'hd20608c;
      24713: inst = 32'h13e00000;
      24714: inst = 32'hfe0a9fb;
      24715: inst = 32'h5be00000;
      24716: inst = 32'h244c8000;
      24717: inst = 32'h24428800;
      24718: inst = 32'h8620000;
      24719: inst = 32'h2a0e0008;
      24720: inst = 32'h294f0009;
      24721: inst = 32'h11200000;
      24722: inst = 32'hd206096;
      24723: inst = 32'h13e00000;
      24724: inst = 32'hfe0a9fb;
      24725: inst = 32'h5be00000;
      24726: inst = 32'h244c8000;
      24727: inst = 32'h24428800;
      24728: inst = 32'h8620000;
      24729: inst = 32'h2a0e0007;
      24730: inst = 32'h294f0009;
      24731: inst = 32'h11200000;
      24732: inst = 32'hd2060a0;
      24733: inst = 32'h13e00000;
      24734: inst = 32'hfe0a9fb;
      24735: inst = 32'h5be00000;
      24736: inst = 32'h244c8000;
      24737: inst = 32'h24428800;
      24738: inst = 32'h8620000;
      24739: inst = 32'h2a0e0005;
      24740: inst = 32'h294f0009;
      24741: inst = 32'h11200000;
      24742: inst = 32'hd2060aa;
      24743: inst = 32'h13e00000;
      24744: inst = 32'hfe0a9fb;
      24745: inst = 32'h5be00000;
      24746: inst = 32'h244c8000;
      24747: inst = 32'h24428800;
      24748: inst = 32'h8620000;
      24749: inst = 32'h2a0e0004;
      24750: inst = 32'h294f0009;
      24751: inst = 32'h11200000;
      24752: inst = 32'hd2060b4;
      24753: inst = 32'h13e00000;
      24754: inst = 32'hfe0a9fb;
      24755: inst = 32'h5be00000;
      24756: inst = 32'h244c8000;
      24757: inst = 32'h24428800;
      24758: inst = 32'h8620000;
      24759: inst = 32'h2a0e0003;
      24760: inst = 32'h294f0009;
      24761: inst = 32'h11200000;
      24762: inst = 32'hd2060be;
      24763: inst = 32'h13e00000;
      24764: inst = 32'hfe0a9fb;
      24765: inst = 32'h5be00000;
      24766: inst = 32'h244c8000;
      24767: inst = 32'h24428800;
      24768: inst = 32'h8620000;
      24769: inst = 32'hc6010ac;
      24770: inst = 32'h2a0e0008;
      24771: inst = 32'h294f000a;
      24772: inst = 32'h11200000;
      24773: inst = 32'hd2060c9;
      24774: inst = 32'h13e00000;
      24775: inst = 32'hfe0a9fb;
      24776: inst = 32'h5be00000;
      24777: inst = 32'h244c8000;
      24778: inst = 32'h24428800;
      24779: inst = 32'h8620000;
      24780: inst = 32'h2a0e0007;
      24781: inst = 32'h294f000a;
      24782: inst = 32'h11200000;
      24783: inst = 32'hd2060d3;
      24784: inst = 32'h13e00000;
      24785: inst = 32'hfe0a9fb;
      24786: inst = 32'h5be00000;
      24787: inst = 32'h244c8000;
      24788: inst = 32'h24428800;
      24789: inst = 32'h8620000;
      24790: inst = 32'h2a0e0006;
      24791: inst = 32'h294f000a;
      24792: inst = 32'h11200000;
      24793: inst = 32'hd2060dd;
      24794: inst = 32'h13e00000;
      24795: inst = 32'hfe0a9fb;
      24796: inst = 32'h5be00000;
      24797: inst = 32'h244c8000;
      24798: inst = 32'h24428800;
      24799: inst = 32'h8620000;
      24800: inst = 32'h2a0e0005;
      24801: inst = 32'h294f000a;
      24802: inst = 32'h11200000;
      24803: inst = 32'hd2060e7;
      24804: inst = 32'h13e00000;
      24805: inst = 32'hfe0a9fb;
      24806: inst = 32'h5be00000;
      24807: inst = 32'h244c8000;
      24808: inst = 32'h24428800;
      24809: inst = 32'h8620000;
      24810: inst = 32'h2a0e0004;
      24811: inst = 32'h294f000a;
      24812: inst = 32'h11200000;
      24813: inst = 32'hd2060f1;
      24814: inst = 32'h13e00000;
      24815: inst = 32'hfe0a9fb;
      24816: inst = 32'h5be00000;
      24817: inst = 32'h244c8000;
      24818: inst = 32'h24428800;
      24819: inst = 32'h8620000;
      24820: inst = 32'h2a0e0003;
      24821: inst = 32'h294f000a;
      24822: inst = 32'h11200000;
      24823: inst = 32'hd2060fb;
      24824: inst = 32'h13e00000;
      24825: inst = 32'hfe0a9fb;
      24826: inst = 32'h5be00000;
      24827: inst = 32'h244c8000;
      24828: inst = 32'h24428800;
      24829: inst = 32'h8620000;
      24830: inst = 32'h13e00000;
      24831: inst = 32'hfe06105;
      24832: inst = 32'h20200001;
      24833: inst = 32'h5be00000;
      24834: inst = 32'h13e00000;
      24835: inst = 32'hfe06108;
      24836: inst = 32'h5be00000;
      24837: inst = 32'h13e00000;
      24838: inst = 32'hfe06108;
      24839: inst = 32'h5be00000;
      24840: inst = 32'h58000000;
      24841: inst = 32'h10408000;
      24842: inst = 32'hc400002;
      24843: inst = 32'h4420000;
      24844: inst = 32'h10600000;
      24845: inst = 32'hc600010;
      24846: inst = 32'h38421800;
      24847: inst = 32'h4042000f;
      24848: inst = 32'h1c40000f;
      24849: inst = 32'h58000000;
      24850: inst = 32'h58200000;
      24851: inst = 32'hc206b50;
      24852: inst = 32'h10408000;
      24853: inst = 32'hc403fe0;
      24854: inst = 32'h8220000;
      24855: inst = 32'h10408000;
      24856: inst = 32'hc403fe1;
      24857: inst = 32'h8220000;
      24858: inst = 32'h10408000;
      24859: inst = 32'hc403fe2;
      24860: inst = 32'h8220000;
      24861: inst = 32'h10408000;
      24862: inst = 32'hc403ff5;
      24863: inst = 32'h8220000;
      24864: inst = 32'h10408000;
      24865: inst = 32'hc403ff8;
      24866: inst = 32'h8220000;
      24867: inst = 32'h10408000;
      24868: inst = 32'hc403ff9;
      24869: inst = 32'h8220000;
      24870: inst = 32'h10408000;
      24871: inst = 32'hc403ffd;
      24872: inst = 32'h8220000;
      24873: inst = 32'h10408000;
      24874: inst = 32'hc403ffe;
      24875: inst = 32'h8220000;
      24876: inst = 32'h10408000;
      24877: inst = 32'hc403fff;
      24878: inst = 32'h8220000;
      24879: inst = 32'h10408000;
      24880: inst = 32'hc404000;
      24881: inst = 32'h8220000;
      24882: inst = 32'h10408000;
      24883: inst = 32'hc404001;
      24884: inst = 32'h8220000;
      24885: inst = 32'h10408000;
      24886: inst = 32'hc404002;
      24887: inst = 32'h8220000;
      24888: inst = 32'h10408000;
      24889: inst = 32'hc404003;
      24890: inst = 32'h8220000;
      24891: inst = 32'h10408000;
      24892: inst = 32'hc404004;
      24893: inst = 32'h8220000;
      24894: inst = 32'h10408000;
      24895: inst = 32'hc404005;
      24896: inst = 32'h8220000;
      24897: inst = 32'h10408000;
      24898: inst = 32'hc404006;
      24899: inst = 32'h8220000;
      24900: inst = 32'h10408000;
      24901: inst = 32'hc404007;
      24902: inst = 32'h8220000;
      24903: inst = 32'h10408000;
      24904: inst = 32'hc404008;
      24905: inst = 32'h8220000;
      24906: inst = 32'h10408000;
      24907: inst = 32'hc404009;
      24908: inst = 32'h8220000;
      24909: inst = 32'h10408000;
      24910: inst = 32'hc40400a;
      24911: inst = 32'h8220000;
      24912: inst = 32'h10408000;
      24913: inst = 32'hc40400b;
      24914: inst = 32'h8220000;
      24915: inst = 32'h10408000;
      24916: inst = 32'hc40400c;
      24917: inst = 32'h8220000;
      24918: inst = 32'h10408000;
      24919: inst = 32'hc40400d;
      24920: inst = 32'h8220000;
      24921: inst = 32'h10408000;
      24922: inst = 32'hc40400e;
      24923: inst = 32'h8220000;
      24924: inst = 32'h10408000;
      24925: inst = 32'hc40400f;
      24926: inst = 32'h8220000;
      24927: inst = 32'h10408000;
      24928: inst = 32'hc404010;
      24929: inst = 32'h8220000;
      24930: inst = 32'h10408000;
      24931: inst = 32'hc404011;
      24932: inst = 32'h8220000;
      24933: inst = 32'h10408000;
      24934: inst = 32'hc404012;
      24935: inst = 32'h8220000;
      24936: inst = 32'h10408000;
      24937: inst = 32'hc404013;
      24938: inst = 32'h8220000;
      24939: inst = 32'h10408000;
      24940: inst = 32'hc404014;
      24941: inst = 32'h8220000;
      24942: inst = 32'h10408000;
      24943: inst = 32'hc404015;
      24944: inst = 32'h8220000;
      24945: inst = 32'h10408000;
      24946: inst = 32'hc404016;
      24947: inst = 32'h8220000;
      24948: inst = 32'h10408000;
      24949: inst = 32'hc404017;
      24950: inst = 32'h8220000;
      24951: inst = 32'h10408000;
      24952: inst = 32'hc404018;
      24953: inst = 32'h8220000;
      24954: inst = 32'h10408000;
      24955: inst = 32'hc404019;
      24956: inst = 32'h8220000;
      24957: inst = 32'h10408000;
      24958: inst = 32'hc40401a;
      24959: inst = 32'h8220000;
      24960: inst = 32'h10408000;
      24961: inst = 32'hc40401b;
      24962: inst = 32'h8220000;
      24963: inst = 32'h10408000;
      24964: inst = 32'hc40401c;
      24965: inst = 32'h8220000;
      24966: inst = 32'h10408000;
      24967: inst = 32'hc40401d;
      24968: inst = 32'h8220000;
      24969: inst = 32'h10408000;
      24970: inst = 32'hc40401e;
      24971: inst = 32'h8220000;
      24972: inst = 32'h10408000;
      24973: inst = 32'hc40401f;
      24974: inst = 32'h8220000;
      24975: inst = 32'h10408000;
      24976: inst = 32'hc404020;
      24977: inst = 32'h8220000;
      24978: inst = 32'h10408000;
      24979: inst = 32'hc404021;
      24980: inst = 32'h8220000;
      24981: inst = 32'h10408000;
      24982: inst = 32'hc404022;
      24983: inst = 32'h8220000;
      24984: inst = 32'h10408000;
      24985: inst = 32'hc404023;
      24986: inst = 32'h8220000;
      24987: inst = 32'h10408000;
      24988: inst = 32'hc404024;
      24989: inst = 32'h8220000;
      24990: inst = 32'h10408000;
      24991: inst = 32'hc404025;
      24992: inst = 32'h8220000;
      24993: inst = 32'h10408000;
      24994: inst = 32'hc404026;
      24995: inst = 32'h8220000;
      24996: inst = 32'h10408000;
      24997: inst = 32'hc404027;
      24998: inst = 32'h8220000;
      24999: inst = 32'h10408000;
      25000: inst = 32'hc404028;
      25001: inst = 32'h8220000;
      25002: inst = 32'h10408000;
      25003: inst = 32'hc404029;
      25004: inst = 32'h8220000;
      25005: inst = 32'h10408000;
      25006: inst = 32'hc40402a;
      25007: inst = 32'h8220000;
      25008: inst = 32'h10408000;
      25009: inst = 32'hc40402b;
      25010: inst = 32'h8220000;
      25011: inst = 32'h10408000;
      25012: inst = 32'hc40402c;
      25013: inst = 32'h8220000;
      25014: inst = 32'h10408000;
      25015: inst = 32'hc40402d;
      25016: inst = 32'h8220000;
      25017: inst = 32'h10408000;
      25018: inst = 32'hc40402e;
      25019: inst = 32'h8220000;
      25020: inst = 32'h10408000;
      25021: inst = 32'hc40402f;
      25022: inst = 32'h8220000;
      25023: inst = 32'h10408000;
      25024: inst = 32'hc404030;
      25025: inst = 32'h8220000;
      25026: inst = 32'h10408000;
      25027: inst = 32'hc404031;
      25028: inst = 32'h8220000;
      25029: inst = 32'h10408000;
      25030: inst = 32'hc404032;
      25031: inst = 32'h8220000;
      25032: inst = 32'h10408000;
      25033: inst = 32'hc404033;
      25034: inst = 32'h8220000;
      25035: inst = 32'h10408000;
      25036: inst = 32'hc404034;
      25037: inst = 32'h8220000;
      25038: inst = 32'h10408000;
      25039: inst = 32'hc404035;
      25040: inst = 32'h8220000;
      25041: inst = 32'h10408000;
      25042: inst = 32'hc404036;
      25043: inst = 32'h8220000;
      25044: inst = 32'h10408000;
      25045: inst = 32'hc404037;
      25046: inst = 32'h8220000;
      25047: inst = 32'h10408000;
      25048: inst = 32'hc404038;
      25049: inst = 32'h8220000;
      25050: inst = 32'h10408000;
      25051: inst = 32'hc404039;
      25052: inst = 32'h8220000;
      25053: inst = 32'h10408000;
      25054: inst = 32'hc40403a;
      25055: inst = 32'h8220000;
      25056: inst = 32'h10408000;
      25057: inst = 32'hc40403b;
      25058: inst = 32'h8220000;
      25059: inst = 32'h10408000;
      25060: inst = 32'hc40403c;
      25061: inst = 32'h8220000;
      25062: inst = 32'h10408000;
      25063: inst = 32'hc40403d;
      25064: inst = 32'h8220000;
      25065: inst = 32'h10408000;
      25066: inst = 32'hc40403e;
      25067: inst = 32'h8220000;
      25068: inst = 32'h10408000;
      25069: inst = 32'hc40403f;
      25070: inst = 32'h8220000;
      25071: inst = 32'h10408000;
      25072: inst = 32'hc404040;
      25073: inst = 32'h8220000;
      25074: inst = 32'h10408000;
      25075: inst = 32'hc404041;
      25076: inst = 32'h8220000;
      25077: inst = 32'h10408000;
      25078: inst = 32'hc404042;
      25079: inst = 32'h8220000;
      25080: inst = 32'h10408000;
      25081: inst = 32'hc404054;
      25082: inst = 32'h8220000;
      25083: inst = 32'h10408000;
      25084: inst = 32'hc404057;
      25085: inst = 32'h8220000;
      25086: inst = 32'h10408000;
      25087: inst = 32'hc404058;
      25088: inst = 32'h8220000;
      25089: inst = 32'h10408000;
      25090: inst = 32'hc40405c;
      25091: inst = 32'h8220000;
      25092: inst = 32'h10408000;
      25093: inst = 32'hc40405d;
      25094: inst = 32'h8220000;
      25095: inst = 32'h10408000;
      25096: inst = 32'hc40405e;
      25097: inst = 32'h8220000;
      25098: inst = 32'h10408000;
      25099: inst = 32'hc40405f;
      25100: inst = 32'h8220000;
      25101: inst = 32'h10408000;
      25102: inst = 32'hc404060;
      25103: inst = 32'h8220000;
      25104: inst = 32'h10408000;
      25105: inst = 32'hc404061;
      25106: inst = 32'h8220000;
      25107: inst = 32'h10408000;
      25108: inst = 32'hc404062;
      25109: inst = 32'h8220000;
      25110: inst = 32'h10408000;
      25111: inst = 32'hc404063;
      25112: inst = 32'h8220000;
      25113: inst = 32'h10408000;
      25114: inst = 32'hc404064;
      25115: inst = 32'h8220000;
      25116: inst = 32'h10408000;
      25117: inst = 32'hc404065;
      25118: inst = 32'h8220000;
      25119: inst = 32'h10408000;
      25120: inst = 32'hc404066;
      25121: inst = 32'h8220000;
      25122: inst = 32'h10408000;
      25123: inst = 32'hc404067;
      25124: inst = 32'h8220000;
      25125: inst = 32'h10408000;
      25126: inst = 32'hc404068;
      25127: inst = 32'h8220000;
      25128: inst = 32'h10408000;
      25129: inst = 32'hc404069;
      25130: inst = 32'h8220000;
      25131: inst = 32'h10408000;
      25132: inst = 32'hc40406a;
      25133: inst = 32'h8220000;
      25134: inst = 32'h10408000;
      25135: inst = 32'hc40406b;
      25136: inst = 32'h8220000;
      25137: inst = 32'h10408000;
      25138: inst = 32'hc40406c;
      25139: inst = 32'h8220000;
      25140: inst = 32'h10408000;
      25141: inst = 32'hc40406d;
      25142: inst = 32'h8220000;
      25143: inst = 32'h10408000;
      25144: inst = 32'hc40406e;
      25145: inst = 32'h8220000;
      25146: inst = 32'h10408000;
      25147: inst = 32'hc40406f;
      25148: inst = 32'h8220000;
      25149: inst = 32'h10408000;
      25150: inst = 32'hc404070;
      25151: inst = 32'h8220000;
      25152: inst = 32'h10408000;
      25153: inst = 32'hc404071;
      25154: inst = 32'h8220000;
      25155: inst = 32'h10408000;
      25156: inst = 32'hc404072;
      25157: inst = 32'h8220000;
      25158: inst = 32'h10408000;
      25159: inst = 32'hc404073;
      25160: inst = 32'h8220000;
      25161: inst = 32'h10408000;
      25162: inst = 32'hc404074;
      25163: inst = 32'h8220000;
      25164: inst = 32'h10408000;
      25165: inst = 32'hc404075;
      25166: inst = 32'h8220000;
      25167: inst = 32'h10408000;
      25168: inst = 32'hc404076;
      25169: inst = 32'h8220000;
      25170: inst = 32'h10408000;
      25171: inst = 32'hc404077;
      25172: inst = 32'h8220000;
      25173: inst = 32'h10408000;
      25174: inst = 32'hc404078;
      25175: inst = 32'h8220000;
      25176: inst = 32'h10408000;
      25177: inst = 32'hc404079;
      25178: inst = 32'h8220000;
      25179: inst = 32'h10408000;
      25180: inst = 32'hc40407a;
      25181: inst = 32'h8220000;
      25182: inst = 32'h10408000;
      25183: inst = 32'hc40407b;
      25184: inst = 32'h8220000;
      25185: inst = 32'h10408000;
      25186: inst = 32'hc40407c;
      25187: inst = 32'h8220000;
      25188: inst = 32'h10408000;
      25189: inst = 32'hc40407d;
      25190: inst = 32'h8220000;
      25191: inst = 32'h10408000;
      25192: inst = 32'hc40407e;
      25193: inst = 32'h8220000;
      25194: inst = 32'h10408000;
      25195: inst = 32'hc40407f;
      25196: inst = 32'h8220000;
      25197: inst = 32'h10408000;
      25198: inst = 32'hc404080;
      25199: inst = 32'h8220000;
      25200: inst = 32'h10408000;
      25201: inst = 32'hc404081;
      25202: inst = 32'h8220000;
      25203: inst = 32'h10408000;
      25204: inst = 32'hc404082;
      25205: inst = 32'h8220000;
      25206: inst = 32'h10408000;
      25207: inst = 32'hc404083;
      25208: inst = 32'h8220000;
      25209: inst = 32'h10408000;
      25210: inst = 32'hc404084;
      25211: inst = 32'h8220000;
      25212: inst = 32'h10408000;
      25213: inst = 32'hc404085;
      25214: inst = 32'h8220000;
      25215: inst = 32'h10408000;
      25216: inst = 32'hc404086;
      25217: inst = 32'h8220000;
      25218: inst = 32'h10408000;
      25219: inst = 32'hc404087;
      25220: inst = 32'h8220000;
      25221: inst = 32'h10408000;
      25222: inst = 32'hc404088;
      25223: inst = 32'h8220000;
      25224: inst = 32'h10408000;
      25225: inst = 32'hc404089;
      25226: inst = 32'h8220000;
      25227: inst = 32'h10408000;
      25228: inst = 32'hc40408a;
      25229: inst = 32'h8220000;
      25230: inst = 32'h10408000;
      25231: inst = 32'hc40408b;
      25232: inst = 32'h8220000;
      25233: inst = 32'h10408000;
      25234: inst = 32'hc40408c;
      25235: inst = 32'h8220000;
      25236: inst = 32'h10408000;
      25237: inst = 32'hc40408d;
      25238: inst = 32'h8220000;
      25239: inst = 32'h10408000;
      25240: inst = 32'hc40408e;
      25241: inst = 32'h8220000;
      25242: inst = 32'h10408000;
      25243: inst = 32'hc40408f;
      25244: inst = 32'h8220000;
      25245: inst = 32'h10408000;
      25246: inst = 32'hc404090;
      25247: inst = 32'h8220000;
      25248: inst = 32'h10408000;
      25249: inst = 32'hc404091;
      25250: inst = 32'h8220000;
      25251: inst = 32'h10408000;
      25252: inst = 32'hc404092;
      25253: inst = 32'h8220000;
      25254: inst = 32'h10408000;
      25255: inst = 32'hc404093;
      25256: inst = 32'h8220000;
      25257: inst = 32'h10408000;
      25258: inst = 32'hc404094;
      25259: inst = 32'h8220000;
      25260: inst = 32'h10408000;
      25261: inst = 32'hc404095;
      25262: inst = 32'h8220000;
      25263: inst = 32'h10408000;
      25264: inst = 32'hc404096;
      25265: inst = 32'h8220000;
      25266: inst = 32'h10408000;
      25267: inst = 32'hc404097;
      25268: inst = 32'h8220000;
      25269: inst = 32'h10408000;
      25270: inst = 32'hc404098;
      25271: inst = 32'h8220000;
      25272: inst = 32'h10408000;
      25273: inst = 32'hc404099;
      25274: inst = 32'h8220000;
      25275: inst = 32'h10408000;
      25276: inst = 32'hc40409a;
      25277: inst = 32'h8220000;
      25278: inst = 32'h10408000;
      25279: inst = 32'hc40409b;
      25280: inst = 32'h8220000;
      25281: inst = 32'h10408000;
      25282: inst = 32'hc40409c;
      25283: inst = 32'h8220000;
      25284: inst = 32'h10408000;
      25285: inst = 32'hc40409d;
      25286: inst = 32'h8220000;
      25287: inst = 32'h10408000;
      25288: inst = 32'hc40409e;
      25289: inst = 32'h8220000;
      25290: inst = 32'h10408000;
      25291: inst = 32'hc40409f;
      25292: inst = 32'h8220000;
      25293: inst = 32'h10408000;
      25294: inst = 32'hc4040a0;
      25295: inst = 32'h8220000;
      25296: inst = 32'h10408000;
      25297: inst = 32'hc4040a1;
      25298: inst = 32'h8220000;
      25299: inst = 32'h10408000;
      25300: inst = 32'hc4040a2;
      25301: inst = 32'h8220000;
      25302: inst = 32'h10408000;
      25303: inst = 32'hc4040af;
      25304: inst = 32'h8220000;
      25305: inst = 32'h10408000;
      25306: inst = 32'hc4040b2;
      25307: inst = 32'h8220000;
      25308: inst = 32'h10408000;
      25309: inst = 32'hc4040b7;
      25310: inst = 32'h8220000;
      25311: inst = 32'h10408000;
      25312: inst = 32'hc4040b8;
      25313: inst = 32'h8220000;
      25314: inst = 32'h10408000;
      25315: inst = 32'hc4040bb;
      25316: inst = 32'h8220000;
      25317: inst = 32'h10408000;
      25318: inst = 32'hc4040bc;
      25319: inst = 32'h8220000;
      25320: inst = 32'h10408000;
      25321: inst = 32'hc4040bd;
      25322: inst = 32'h8220000;
      25323: inst = 32'h10408000;
      25324: inst = 32'hc4040be;
      25325: inst = 32'h8220000;
      25326: inst = 32'h10408000;
      25327: inst = 32'hc4040bf;
      25328: inst = 32'h8220000;
      25329: inst = 32'h10408000;
      25330: inst = 32'hc4040c0;
      25331: inst = 32'h8220000;
      25332: inst = 32'h10408000;
      25333: inst = 32'hc4040c1;
      25334: inst = 32'h8220000;
      25335: inst = 32'h10408000;
      25336: inst = 32'hc4040c2;
      25337: inst = 32'h8220000;
      25338: inst = 32'h10408000;
      25339: inst = 32'hc4040c3;
      25340: inst = 32'h8220000;
      25341: inst = 32'h10408000;
      25342: inst = 32'hc4040c4;
      25343: inst = 32'h8220000;
      25344: inst = 32'h10408000;
      25345: inst = 32'hc4040c5;
      25346: inst = 32'h8220000;
      25347: inst = 32'h10408000;
      25348: inst = 32'hc4040c6;
      25349: inst = 32'h8220000;
      25350: inst = 32'h10408000;
      25351: inst = 32'hc4040c7;
      25352: inst = 32'h8220000;
      25353: inst = 32'h10408000;
      25354: inst = 32'hc4040c8;
      25355: inst = 32'h8220000;
      25356: inst = 32'h10408000;
      25357: inst = 32'hc4040c9;
      25358: inst = 32'h8220000;
      25359: inst = 32'h10408000;
      25360: inst = 32'hc4040ca;
      25361: inst = 32'h8220000;
      25362: inst = 32'h10408000;
      25363: inst = 32'hc4040cb;
      25364: inst = 32'h8220000;
      25365: inst = 32'h10408000;
      25366: inst = 32'hc4040cc;
      25367: inst = 32'h8220000;
      25368: inst = 32'h10408000;
      25369: inst = 32'hc4040cd;
      25370: inst = 32'h8220000;
      25371: inst = 32'h10408000;
      25372: inst = 32'hc4040ce;
      25373: inst = 32'h8220000;
      25374: inst = 32'h10408000;
      25375: inst = 32'hc4040cf;
      25376: inst = 32'h8220000;
      25377: inst = 32'h10408000;
      25378: inst = 32'hc4040d0;
      25379: inst = 32'h8220000;
      25380: inst = 32'h10408000;
      25381: inst = 32'hc4040d1;
      25382: inst = 32'h8220000;
      25383: inst = 32'h10408000;
      25384: inst = 32'hc4040d2;
      25385: inst = 32'h8220000;
      25386: inst = 32'h10408000;
      25387: inst = 32'hc4040d3;
      25388: inst = 32'h8220000;
      25389: inst = 32'h10408000;
      25390: inst = 32'hc4040d4;
      25391: inst = 32'h8220000;
      25392: inst = 32'h10408000;
      25393: inst = 32'hc4040d5;
      25394: inst = 32'h8220000;
      25395: inst = 32'h10408000;
      25396: inst = 32'hc4040d6;
      25397: inst = 32'h8220000;
      25398: inst = 32'h10408000;
      25399: inst = 32'hc4040d7;
      25400: inst = 32'h8220000;
      25401: inst = 32'h10408000;
      25402: inst = 32'hc4040d8;
      25403: inst = 32'h8220000;
      25404: inst = 32'h10408000;
      25405: inst = 32'hc4040d9;
      25406: inst = 32'h8220000;
      25407: inst = 32'h10408000;
      25408: inst = 32'hc4040da;
      25409: inst = 32'h8220000;
      25410: inst = 32'h10408000;
      25411: inst = 32'hc4040db;
      25412: inst = 32'h8220000;
      25413: inst = 32'h10408000;
      25414: inst = 32'hc4040dc;
      25415: inst = 32'h8220000;
      25416: inst = 32'h10408000;
      25417: inst = 32'hc4040dd;
      25418: inst = 32'h8220000;
      25419: inst = 32'h10408000;
      25420: inst = 32'hc4040de;
      25421: inst = 32'h8220000;
      25422: inst = 32'h10408000;
      25423: inst = 32'hc4040df;
      25424: inst = 32'h8220000;
      25425: inst = 32'h10408000;
      25426: inst = 32'hc4040e0;
      25427: inst = 32'h8220000;
      25428: inst = 32'h10408000;
      25429: inst = 32'hc4040e1;
      25430: inst = 32'h8220000;
      25431: inst = 32'h10408000;
      25432: inst = 32'hc4040e2;
      25433: inst = 32'h8220000;
      25434: inst = 32'h10408000;
      25435: inst = 32'hc4040e3;
      25436: inst = 32'h8220000;
      25437: inst = 32'h10408000;
      25438: inst = 32'hc4040e4;
      25439: inst = 32'h8220000;
      25440: inst = 32'h10408000;
      25441: inst = 32'hc4040e5;
      25442: inst = 32'h8220000;
      25443: inst = 32'h10408000;
      25444: inst = 32'hc4040e6;
      25445: inst = 32'h8220000;
      25446: inst = 32'h10408000;
      25447: inst = 32'hc4040e7;
      25448: inst = 32'h8220000;
      25449: inst = 32'h10408000;
      25450: inst = 32'hc4040e8;
      25451: inst = 32'h8220000;
      25452: inst = 32'h10408000;
      25453: inst = 32'hc4040e9;
      25454: inst = 32'h8220000;
      25455: inst = 32'h10408000;
      25456: inst = 32'hc4040ea;
      25457: inst = 32'h8220000;
      25458: inst = 32'h10408000;
      25459: inst = 32'hc4040eb;
      25460: inst = 32'h8220000;
      25461: inst = 32'h10408000;
      25462: inst = 32'hc4040ec;
      25463: inst = 32'h8220000;
      25464: inst = 32'h10408000;
      25465: inst = 32'hc4040ed;
      25466: inst = 32'h8220000;
      25467: inst = 32'h10408000;
      25468: inst = 32'hc4040ee;
      25469: inst = 32'h8220000;
      25470: inst = 32'h10408000;
      25471: inst = 32'hc4040ef;
      25472: inst = 32'h8220000;
      25473: inst = 32'h10408000;
      25474: inst = 32'hc4040f0;
      25475: inst = 32'h8220000;
      25476: inst = 32'h10408000;
      25477: inst = 32'hc4040f1;
      25478: inst = 32'h8220000;
      25479: inst = 32'h10408000;
      25480: inst = 32'hc4040f2;
      25481: inst = 32'h8220000;
      25482: inst = 32'h10408000;
      25483: inst = 32'hc4040f3;
      25484: inst = 32'h8220000;
      25485: inst = 32'h10408000;
      25486: inst = 32'hc4040f4;
      25487: inst = 32'h8220000;
      25488: inst = 32'h10408000;
      25489: inst = 32'hc4040f5;
      25490: inst = 32'h8220000;
      25491: inst = 32'h10408000;
      25492: inst = 32'hc4040f6;
      25493: inst = 32'h8220000;
      25494: inst = 32'h10408000;
      25495: inst = 32'hc4040f7;
      25496: inst = 32'h8220000;
      25497: inst = 32'h10408000;
      25498: inst = 32'hc4040f8;
      25499: inst = 32'h8220000;
      25500: inst = 32'h10408000;
      25501: inst = 32'hc4040f9;
      25502: inst = 32'h8220000;
      25503: inst = 32'h10408000;
      25504: inst = 32'hc4040fa;
      25505: inst = 32'h8220000;
      25506: inst = 32'h10408000;
      25507: inst = 32'hc4040fb;
      25508: inst = 32'h8220000;
      25509: inst = 32'h10408000;
      25510: inst = 32'hc4040fc;
      25511: inst = 32'h8220000;
      25512: inst = 32'h10408000;
      25513: inst = 32'hc4040fd;
      25514: inst = 32'h8220000;
      25515: inst = 32'h10408000;
      25516: inst = 32'hc4040fe;
      25517: inst = 32'h8220000;
      25518: inst = 32'h10408000;
      25519: inst = 32'hc4040ff;
      25520: inst = 32'h8220000;
      25521: inst = 32'h10408000;
      25522: inst = 32'hc404100;
      25523: inst = 32'h8220000;
      25524: inst = 32'h10408000;
      25525: inst = 32'hc404101;
      25526: inst = 32'h8220000;
      25527: inst = 32'h10408000;
      25528: inst = 32'hc404102;
      25529: inst = 32'h8220000;
      25530: inst = 32'h10408000;
      25531: inst = 32'hc40414c;
      25532: inst = 32'h8220000;
      25533: inst = 32'h10408000;
      25534: inst = 32'hc40414d;
      25535: inst = 32'h8220000;
      25536: inst = 32'h10408000;
      25537: inst = 32'hc40414e;
      25538: inst = 32'h8220000;
      25539: inst = 32'h10408000;
      25540: inst = 32'hc40415d;
      25541: inst = 32'h8220000;
      25542: inst = 32'h10408000;
      25543: inst = 32'hc40415e;
      25544: inst = 32'h8220000;
      25545: inst = 32'h10408000;
      25546: inst = 32'hc40415f;
      25547: inst = 32'h8220000;
      25548: inst = 32'h10408000;
      25549: inst = 32'hc404160;
      25550: inst = 32'h8220000;
      25551: inst = 32'h10408000;
      25552: inst = 32'hc404161;
      25553: inst = 32'h8220000;
      25554: inst = 32'h10408000;
      25555: inst = 32'hc404162;
      25556: inst = 32'h8220000;
      25557: inst = 32'h10408000;
      25558: inst = 32'hc4041ac;
      25559: inst = 32'h8220000;
      25560: inst = 32'h10408000;
      25561: inst = 32'hc4041ad;
      25562: inst = 32'h8220000;
      25563: inst = 32'h10408000;
      25564: inst = 32'hc4041ae;
      25565: inst = 32'h8220000;
      25566: inst = 32'h10408000;
      25567: inst = 32'hc4041bd;
      25568: inst = 32'h8220000;
      25569: inst = 32'h10408000;
      25570: inst = 32'hc4041be;
      25571: inst = 32'h8220000;
      25572: inst = 32'h10408000;
      25573: inst = 32'hc4041bf;
      25574: inst = 32'h8220000;
      25575: inst = 32'h10408000;
      25576: inst = 32'hc4041c0;
      25577: inst = 32'h8220000;
      25578: inst = 32'h10408000;
      25579: inst = 32'hc4041c1;
      25580: inst = 32'h8220000;
      25581: inst = 32'h10408000;
      25582: inst = 32'hc4041c2;
      25583: inst = 32'h8220000;
      25584: inst = 32'h10408000;
      25585: inst = 32'hc40420c;
      25586: inst = 32'h8220000;
      25587: inst = 32'h10408000;
      25588: inst = 32'hc40420d;
      25589: inst = 32'h8220000;
      25590: inst = 32'h10408000;
      25591: inst = 32'hc40420e;
      25592: inst = 32'h8220000;
      25593: inst = 32'h10408000;
      25594: inst = 32'hc40421d;
      25595: inst = 32'h8220000;
      25596: inst = 32'h10408000;
      25597: inst = 32'hc40421e;
      25598: inst = 32'h8220000;
      25599: inst = 32'h10408000;
      25600: inst = 32'hc40421f;
      25601: inst = 32'h8220000;
      25602: inst = 32'h10408000;
      25603: inst = 32'hc404220;
      25604: inst = 32'h8220000;
      25605: inst = 32'h10408000;
      25606: inst = 32'hc404221;
      25607: inst = 32'h8220000;
      25608: inst = 32'h10408000;
      25609: inst = 32'hc404222;
      25610: inst = 32'h8220000;
      25611: inst = 32'h10408000;
      25612: inst = 32'hc40426c;
      25613: inst = 32'h8220000;
      25614: inst = 32'h10408000;
      25615: inst = 32'hc40426d;
      25616: inst = 32'h8220000;
      25617: inst = 32'h10408000;
      25618: inst = 32'hc40426e;
      25619: inst = 32'h8220000;
      25620: inst = 32'h10408000;
      25621: inst = 32'hc40427d;
      25622: inst = 32'h8220000;
      25623: inst = 32'h10408000;
      25624: inst = 32'hc40427e;
      25625: inst = 32'h8220000;
      25626: inst = 32'h10408000;
      25627: inst = 32'hc40427f;
      25628: inst = 32'h8220000;
      25629: inst = 32'h10408000;
      25630: inst = 32'hc404280;
      25631: inst = 32'h8220000;
      25632: inst = 32'h10408000;
      25633: inst = 32'hc404281;
      25634: inst = 32'h8220000;
      25635: inst = 32'h10408000;
      25636: inst = 32'hc404282;
      25637: inst = 32'h8220000;
      25638: inst = 32'h10408000;
      25639: inst = 32'hc4042cc;
      25640: inst = 32'h8220000;
      25641: inst = 32'h10408000;
      25642: inst = 32'hc4042cd;
      25643: inst = 32'h8220000;
      25644: inst = 32'h10408000;
      25645: inst = 32'hc4042ce;
      25646: inst = 32'h8220000;
      25647: inst = 32'h10408000;
      25648: inst = 32'hc4042dd;
      25649: inst = 32'h8220000;
      25650: inst = 32'h10408000;
      25651: inst = 32'hc4042de;
      25652: inst = 32'h8220000;
      25653: inst = 32'h10408000;
      25654: inst = 32'hc4042df;
      25655: inst = 32'h8220000;
      25656: inst = 32'h10408000;
      25657: inst = 32'hc4042e0;
      25658: inst = 32'h8220000;
      25659: inst = 32'h10408000;
      25660: inst = 32'hc4042e1;
      25661: inst = 32'h8220000;
      25662: inst = 32'h10408000;
      25663: inst = 32'hc4042e2;
      25664: inst = 32'h8220000;
      25665: inst = 32'h10408000;
      25666: inst = 32'hc40432c;
      25667: inst = 32'h8220000;
      25668: inst = 32'h10408000;
      25669: inst = 32'hc40432d;
      25670: inst = 32'h8220000;
      25671: inst = 32'h10408000;
      25672: inst = 32'hc40432e;
      25673: inst = 32'h8220000;
      25674: inst = 32'h10408000;
      25675: inst = 32'hc40433d;
      25676: inst = 32'h8220000;
      25677: inst = 32'h10408000;
      25678: inst = 32'hc40433e;
      25679: inst = 32'h8220000;
      25680: inst = 32'h10408000;
      25681: inst = 32'hc40433f;
      25682: inst = 32'h8220000;
      25683: inst = 32'h10408000;
      25684: inst = 32'hc404340;
      25685: inst = 32'h8220000;
      25686: inst = 32'h10408000;
      25687: inst = 32'hc404341;
      25688: inst = 32'h8220000;
      25689: inst = 32'h10408000;
      25690: inst = 32'hc404342;
      25691: inst = 32'h8220000;
      25692: inst = 32'h10408000;
      25693: inst = 32'hc40438c;
      25694: inst = 32'h8220000;
      25695: inst = 32'h10408000;
      25696: inst = 32'hc40438d;
      25697: inst = 32'h8220000;
      25698: inst = 32'h10408000;
      25699: inst = 32'hc40438e;
      25700: inst = 32'h8220000;
      25701: inst = 32'h10408000;
      25702: inst = 32'hc40439d;
      25703: inst = 32'h8220000;
      25704: inst = 32'h10408000;
      25705: inst = 32'hc40439e;
      25706: inst = 32'h8220000;
      25707: inst = 32'h10408000;
      25708: inst = 32'hc40439f;
      25709: inst = 32'h8220000;
      25710: inst = 32'h10408000;
      25711: inst = 32'hc4043a0;
      25712: inst = 32'h8220000;
      25713: inst = 32'h10408000;
      25714: inst = 32'hc4043a1;
      25715: inst = 32'h8220000;
      25716: inst = 32'h10408000;
      25717: inst = 32'hc4043a2;
      25718: inst = 32'h8220000;
      25719: inst = 32'h10408000;
      25720: inst = 32'hc4043ec;
      25721: inst = 32'h8220000;
      25722: inst = 32'h10408000;
      25723: inst = 32'hc4043ed;
      25724: inst = 32'h8220000;
      25725: inst = 32'h10408000;
      25726: inst = 32'hc4043ee;
      25727: inst = 32'h8220000;
      25728: inst = 32'h10408000;
      25729: inst = 32'hc4043fd;
      25730: inst = 32'h8220000;
      25731: inst = 32'h10408000;
      25732: inst = 32'hc4043fe;
      25733: inst = 32'h8220000;
      25734: inst = 32'h10408000;
      25735: inst = 32'hc4043ff;
      25736: inst = 32'h8220000;
      25737: inst = 32'h10408000;
      25738: inst = 32'hc404400;
      25739: inst = 32'h8220000;
      25740: inst = 32'h10408000;
      25741: inst = 32'hc404401;
      25742: inst = 32'h8220000;
      25743: inst = 32'h10408000;
      25744: inst = 32'hc404402;
      25745: inst = 32'h8220000;
      25746: inst = 32'h10408000;
      25747: inst = 32'hc40444c;
      25748: inst = 32'h8220000;
      25749: inst = 32'h10408000;
      25750: inst = 32'hc40444d;
      25751: inst = 32'h8220000;
      25752: inst = 32'h10408000;
      25753: inst = 32'hc40444e;
      25754: inst = 32'h8220000;
      25755: inst = 32'h10408000;
      25756: inst = 32'hc40445d;
      25757: inst = 32'h8220000;
      25758: inst = 32'h10408000;
      25759: inst = 32'hc40445e;
      25760: inst = 32'h8220000;
      25761: inst = 32'h10408000;
      25762: inst = 32'hc40445f;
      25763: inst = 32'h8220000;
      25764: inst = 32'h10408000;
      25765: inst = 32'hc404460;
      25766: inst = 32'h8220000;
      25767: inst = 32'h10408000;
      25768: inst = 32'hc404461;
      25769: inst = 32'h8220000;
      25770: inst = 32'h10408000;
      25771: inst = 32'hc404462;
      25772: inst = 32'h8220000;
      25773: inst = 32'h10408000;
      25774: inst = 32'hc4044ac;
      25775: inst = 32'h8220000;
      25776: inst = 32'h10408000;
      25777: inst = 32'hc4044ad;
      25778: inst = 32'h8220000;
      25779: inst = 32'h10408000;
      25780: inst = 32'hc4044ae;
      25781: inst = 32'h8220000;
      25782: inst = 32'h10408000;
      25783: inst = 32'hc4044bd;
      25784: inst = 32'h8220000;
      25785: inst = 32'h10408000;
      25786: inst = 32'hc4044be;
      25787: inst = 32'h8220000;
      25788: inst = 32'h10408000;
      25789: inst = 32'hc4044bf;
      25790: inst = 32'h8220000;
      25791: inst = 32'h10408000;
      25792: inst = 32'hc4044c0;
      25793: inst = 32'h8220000;
      25794: inst = 32'h10408000;
      25795: inst = 32'hc4044c1;
      25796: inst = 32'h8220000;
      25797: inst = 32'h10408000;
      25798: inst = 32'hc4044c2;
      25799: inst = 32'h8220000;
      25800: inst = 32'h10408000;
      25801: inst = 32'hc40450c;
      25802: inst = 32'h8220000;
      25803: inst = 32'h10408000;
      25804: inst = 32'hc40450d;
      25805: inst = 32'h8220000;
      25806: inst = 32'h10408000;
      25807: inst = 32'hc40450e;
      25808: inst = 32'h8220000;
      25809: inst = 32'h10408000;
      25810: inst = 32'hc40451d;
      25811: inst = 32'h8220000;
      25812: inst = 32'h10408000;
      25813: inst = 32'hc40451e;
      25814: inst = 32'h8220000;
      25815: inst = 32'h10408000;
      25816: inst = 32'hc40451f;
      25817: inst = 32'h8220000;
      25818: inst = 32'h10408000;
      25819: inst = 32'hc404520;
      25820: inst = 32'h8220000;
      25821: inst = 32'h10408000;
      25822: inst = 32'hc404521;
      25823: inst = 32'h8220000;
      25824: inst = 32'h10408000;
      25825: inst = 32'hc404522;
      25826: inst = 32'h8220000;
      25827: inst = 32'h10408000;
      25828: inst = 32'hc40456c;
      25829: inst = 32'h8220000;
      25830: inst = 32'h10408000;
      25831: inst = 32'hc40456d;
      25832: inst = 32'h8220000;
      25833: inst = 32'h10408000;
      25834: inst = 32'hc40456e;
      25835: inst = 32'h8220000;
      25836: inst = 32'h10408000;
      25837: inst = 32'hc40457d;
      25838: inst = 32'h8220000;
      25839: inst = 32'h10408000;
      25840: inst = 32'hc40457e;
      25841: inst = 32'h8220000;
      25842: inst = 32'h10408000;
      25843: inst = 32'hc40457f;
      25844: inst = 32'h8220000;
      25845: inst = 32'h10408000;
      25846: inst = 32'hc404580;
      25847: inst = 32'h8220000;
      25848: inst = 32'h10408000;
      25849: inst = 32'hc404581;
      25850: inst = 32'h8220000;
      25851: inst = 32'h10408000;
      25852: inst = 32'hc404582;
      25853: inst = 32'h8220000;
      25854: inst = 32'h10408000;
      25855: inst = 32'hc4045cc;
      25856: inst = 32'h8220000;
      25857: inst = 32'h10408000;
      25858: inst = 32'hc4045cd;
      25859: inst = 32'h8220000;
      25860: inst = 32'h10408000;
      25861: inst = 32'hc4045ce;
      25862: inst = 32'h8220000;
      25863: inst = 32'h10408000;
      25864: inst = 32'hc4045dd;
      25865: inst = 32'h8220000;
      25866: inst = 32'h10408000;
      25867: inst = 32'hc4045de;
      25868: inst = 32'h8220000;
      25869: inst = 32'h10408000;
      25870: inst = 32'hc4045df;
      25871: inst = 32'h8220000;
      25872: inst = 32'h10408000;
      25873: inst = 32'hc4045e0;
      25874: inst = 32'h8220000;
      25875: inst = 32'h10408000;
      25876: inst = 32'hc4045e1;
      25877: inst = 32'h8220000;
      25878: inst = 32'h10408000;
      25879: inst = 32'hc4045e2;
      25880: inst = 32'h8220000;
      25881: inst = 32'h10408000;
      25882: inst = 32'hc40462c;
      25883: inst = 32'h8220000;
      25884: inst = 32'h10408000;
      25885: inst = 32'hc40462d;
      25886: inst = 32'h8220000;
      25887: inst = 32'h10408000;
      25888: inst = 32'hc40462e;
      25889: inst = 32'h8220000;
      25890: inst = 32'h10408000;
      25891: inst = 32'hc40463d;
      25892: inst = 32'h8220000;
      25893: inst = 32'h10408000;
      25894: inst = 32'hc40463e;
      25895: inst = 32'h8220000;
      25896: inst = 32'h10408000;
      25897: inst = 32'hc40463f;
      25898: inst = 32'h8220000;
      25899: inst = 32'h10408000;
      25900: inst = 32'hc404640;
      25901: inst = 32'h8220000;
      25902: inst = 32'h10408000;
      25903: inst = 32'hc404641;
      25904: inst = 32'h8220000;
      25905: inst = 32'h10408000;
      25906: inst = 32'hc404642;
      25907: inst = 32'h8220000;
      25908: inst = 32'h10408000;
      25909: inst = 32'hc40464e;
      25910: inst = 32'h8220000;
      25911: inst = 32'h10408000;
      25912: inst = 32'hc40464f;
      25913: inst = 32'h8220000;
      25914: inst = 32'h10408000;
      25915: inst = 32'hc404650;
      25916: inst = 32'h8220000;
      25917: inst = 32'h10408000;
      25918: inst = 32'hc404651;
      25919: inst = 32'h8220000;
      25920: inst = 32'h10408000;
      25921: inst = 32'hc404652;
      25922: inst = 32'h8220000;
      25923: inst = 32'h10408000;
      25924: inst = 32'hc404653;
      25925: inst = 32'h8220000;
      25926: inst = 32'h10408000;
      25927: inst = 32'hc404654;
      25928: inst = 32'h8220000;
      25929: inst = 32'h10408000;
      25930: inst = 32'hc404655;
      25931: inst = 32'h8220000;
      25932: inst = 32'h10408000;
      25933: inst = 32'hc404656;
      25934: inst = 32'h8220000;
      25935: inst = 32'h10408000;
      25936: inst = 32'hc404657;
      25937: inst = 32'h8220000;
      25938: inst = 32'h10408000;
      25939: inst = 32'hc404658;
      25940: inst = 32'h8220000;
      25941: inst = 32'h10408000;
      25942: inst = 32'hc404659;
      25943: inst = 32'h8220000;
      25944: inst = 32'h10408000;
      25945: inst = 32'hc40465a;
      25946: inst = 32'h8220000;
      25947: inst = 32'h10408000;
      25948: inst = 32'hc40465b;
      25949: inst = 32'h8220000;
      25950: inst = 32'h10408000;
      25951: inst = 32'hc40465c;
      25952: inst = 32'h8220000;
      25953: inst = 32'h10408000;
      25954: inst = 32'hc40465d;
      25955: inst = 32'h8220000;
      25956: inst = 32'h10408000;
      25957: inst = 32'hc40465e;
      25958: inst = 32'h8220000;
      25959: inst = 32'h10408000;
      25960: inst = 32'hc40465f;
      25961: inst = 32'h8220000;
      25962: inst = 32'h10408000;
      25963: inst = 32'hc404660;
      25964: inst = 32'h8220000;
      25965: inst = 32'h10408000;
      25966: inst = 32'hc404661;
      25967: inst = 32'h8220000;
      25968: inst = 32'h10408000;
      25969: inst = 32'hc404662;
      25970: inst = 32'h8220000;
      25971: inst = 32'h10408000;
      25972: inst = 32'hc404663;
      25973: inst = 32'h8220000;
      25974: inst = 32'h10408000;
      25975: inst = 32'hc404664;
      25976: inst = 32'h8220000;
      25977: inst = 32'h10408000;
      25978: inst = 32'hc404665;
      25979: inst = 32'h8220000;
      25980: inst = 32'h10408000;
      25981: inst = 32'hc404666;
      25982: inst = 32'h8220000;
      25983: inst = 32'h10408000;
      25984: inst = 32'hc404667;
      25985: inst = 32'h8220000;
      25986: inst = 32'h10408000;
      25987: inst = 32'hc404668;
      25988: inst = 32'h8220000;
      25989: inst = 32'h10408000;
      25990: inst = 32'hc404669;
      25991: inst = 32'h8220000;
      25992: inst = 32'h10408000;
      25993: inst = 32'hc40466e;
      25994: inst = 32'h8220000;
      25995: inst = 32'h10408000;
      25996: inst = 32'hc40466f;
      25997: inst = 32'h8220000;
      25998: inst = 32'h10408000;
      25999: inst = 32'hc404673;
      26000: inst = 32'h8220000;
      26001: inst = 32'h10408000;
      26002: inst = 32'hc404676;
      26003: inst = 32'h8220000;
      26004: inst = 32'h10408000;
      26005: inst = 32'hc40468c;
      26006: inst = 32'h8220000;
      26007: inst = 32'h10408000;
      26008: inst = 32'hc40468d;
      26009: inst = 32'h8220000;
      26010: inst = 32'h10408000;
      26011: inst = 32'hc40468e;
      26012: inst = 32'h8220000;
      26013: inst = 32'h10408000;
      26014: inst = 32'hc40469d;
      26015: inst = 32'h8220000;
      26016: inst = 32'h10408000;
      26017: inst = 32'hc40469e;
      26018: inst = 32'h8220000;
      26019: inst = 32'h10408000;
      26020: inst = 32'hc40469f;
      26021: inst = 32'h8220000;
      26022: inst = 32'h10408000;
      26023: inst = 32'hc4046a0;
      26024: inst = 32'h8220000;
      26025: inst = 32'h10408000;
      26026: inst = 32'hc4046a1;
      26027: inst = 32'h8220000;
      26028: inst = 32'h10408000;
      26029: inst = 32'hc4046a2;
      26030: inst = 32'h8220000;
      26031: inst = 32'h10408000;
      26032: inst = 32'hc4046ae;
      26033: inst = 32'h8220000;
      26034: inst = 32'h10408000;
      26035: inst = 32'hc4046af;
      26036: inst = 32'h8220000;
      26037: inst = 32'h10408000;
      26038: inst = 32'hc4046b0;
      26039: inst = 32'h8220000;
      26040: inst = 32'h10408000;
      26041: inst = 32'hc4046b1;
      26042: inst = 32'h8220000;
      26043: inst = 32'h10408000;
      26044: inst = 32'hc4046b2;
      26045: inst = 32'h8220000;
      26046: inst = 32'h10408000;
      26047: inst = 32'hc4046b3;
      26048: inst = 32'h8220000;
      26049: inst = 32'h10408000;
      26050: inst = 32'hc4046b4;
      26051: inst = 32'h8220000;
      26052: inst = 32'h10408000;
      26053: inst = 32'hc4046b5;
      26054: inst = 32'h8220000;
      26055: inst = 32'h10408000;
      26056: inst = 32'hc4046b6;
      26057: inst = 32'h8220000;
      26058: inst = 32'h10408000;
      26059: inst = 32'hc4046b7;
      26060: inst = 32'h8220000;
      26061: inst = 32'h10408000;
      26062: inst = 32'hc4046b8;
      26063: inst = 32'h8220000;
      26064: inst = 32'h10408000;
      26065: inst = 32'hc4046b9;
      26066: inst = 32'h8220000;
      26067: inst = 32'h10408000;
      26068: inst = 32'hc4046ba;
      26069: inst = 32'h8220000;
      26070: inst = 32'h10408000;
      26071: inst = 32'hc4046bb;
      26072: inst = 32'h8220000;
      26073: inst = 32'h10408000;
      26074: inst = 32'hc4046bc;
      26075: inst = 32'h8220000;
      26076: inst = 32'h10408000;
      26077: inst = 32'hc4046bd;
      26078: inst = 32'h8220000;
      26079: inst = 32'h10408000;
      26080: inst = 32'hc4046be;
      26081: inst = 32'h8220000;
      26082: inst = 32'h10408000;
      26083: inst = 32'hc4046bf;
      26084: inst = 32'h8220000;
      26085: inst = 32'h10408000;
      26086: inst = 32'hc4046c0;
      26087: inst = 32'h8220000;
      26088: inst = 32'h10408000;
      26089: inst = 32'hc4046c1;
      26090: inst = 32'h8220000;
      26091: inst = 32'h10408000;
      26092: inst = 32'hc4046c2;
      26093: inst = 32'h8220000;
      26094: inst = 32'h10408000;
      26095: inst = 32'hc4046c3;
      26096: inst = 32'h8220000;
      26097: inst = 32'h10408000;
      26098: inst = 32'hc4046c4;
      26099: inst = 32'h8220000;
      26100: inst = 32'h10408000;
      26101: inst = 32'hc4046c5;
      26102: inst = 32'h8220000;
      26103: inst = 32'h10408000;
      26104: inst = 32'hc4046c6;
      26105: inst = 32'h8220000;
      26106: inst = 32'h10408000;
      26107: inst = 32'hc4046c7;
      26108: inst = 32'h8220000;
      26109: inst = 32'h10408000;
      26110: inst = 32'hc4046c8;
      26111: inst = 32'h8220000;
      26112: inst = 32'h10408000;
      26113: inst = 32'hc4046c9;
      26114: inst = 32'h8220000;
      26115: inst = 32'h10408000;
      26116: inst = 32'hc4046ce;
      26117: inst = 32'h8220000;
      26118: inst = 32'h10408000;
      26119: inst = 32'hc4046cf;
      26120: inst = 32'h8220000;
      26121: inst = 32'h10408000;
      26122: inst = 32'hc4046d0;
      26123: inst = 32'h8220000;
      26124: inst = 32'h10408000;
      26125: inst = 32'hc4046d1;
      26126: inst = 32'h8220000;
      26127: inst = 32'h10408000;
      26128: inst = 32'hc4046d6;
      26129: inst = 32'h8220000;
      26130: inst = 32'h10408000;
      26131: inst = 32'hc4046ec;
      26132: inst = 32'h8220000;
      26133: inst = 32'h10408000;
      26134: inst = 32'hc4046ed;
      26135: inst = 32'h8220000;
      26136: inst = 32'h10408000;
      26137: inst = 32'hc4046ee;
      26138: inst = 32'h8220000;
      26139: inst = 32'h10408000;
      26140: inst = 32'hc4046fd;
      26141: inst = 32'h8220000;
      26142: inst = 32'h10408000;
      26143: inst = 32'hc4046fe;
      26144: inst = 32'h8220000;
      26145: inst = 32'h10408000;
      26146: inst = 32'hc4046ff;
      26147: inst = 32'h8220000;
      26148: inst = 32'h10408000;
      26149: inst = 32'hc404700;
      26150: inst = 32'h8220000;
      26151: inst = 32'h10408000;
      26152: inst = 32'hc404701;
      26153: inst = 32'h8220000;
      26154: inst = 32'h10408000;
      26155: inst = 32'hc404702;
      26156: inst = 32'h8220000;
      26157: inst = 32'h10408000;
      26158: inst = 32'hc40470e;
      26159: inst = 32'h8220000;
      26160: inst = 32'h10408000;
      26161: inst = 32'hc40470f;
      26162: inst = 32'h8220000;
      26163: inst = 32'h10408000;
      26164: inst = 32'hc404710;
      26165: inst = 32'h8220000;
      26166: inst = 32'h10408000;
      26167: inst = 32'hc404711;
      26168: inst = 32'h8220000;
      26169: inst = 32'h10408000;
      26170: inst = 32'hc404712;
      26171: inst = 32'h8220000;
      26172: inst = 32'h10408000;
      26173: inst = 32'hc404713;
      26174: inst = 32'h8220000;
      26175: inst = 32'h10408000;
      26176: inst = 32'hc404714;
      26177: inst = 32'h8220000;
      26178: inst = 32'h10408000;
      26179: inst = 32'hc404715;
      26180: inst = 32'h8220000;
      26181: inst = 32'h10408000;
      26182: inst = 32'hc404716;
      26183: inst = 32'h8220000;
      26184: inst = 32'h10408000;
      26185: inst = 32'hc404717;
      26186: inst = 32'h8220000;
      26187: inst = 32'h10408000;
      26188: inst = 32'hc404718;
      26189: inst = 32'h8220000;
      26190: inst = 32'h10408000;
      26191: inst = 32'hc404719;
      26192: inst = 32'h8220000;
      26193: inst = 32'h10408000;
      26194: inst = 32'hc40471a;
      26195: inst = 32'h8220000;
      26196: inst = 32'h10408000;
      26197: inst = 32'hc40471b;
      26198: inst = 32'h8220000;
      26199: inst = 32'h10408000;
      26200: inst = 32'hc40471c;
      26201: inst = 32'h8220000;
      26202: inst = 32'h10408000;
      26203: inst = 32'hc40471d;
      26204: inst = 32'h8220000;
      26205: inst = 32'h10408000;
      26206: inst = 32'hc40471e;
      26207: inst = 32'h8220000;
      26208: inst = 32'h10408000;
      26209: inst = 32'hc40471f;
      26210: inst = 32'h8220000;
      26211: inst = 32'h10408000;
      26212: inst = 32'hc404720;
      26213: inst = 32'h8220000;
      26214: inst = 32'h10408000;
      26215: inst = 32'hc404721;
      26216: inst = 32'h8220000;
      26217: inst = 32'h10408000;
      26218: inst = 32'hc404722;
      26219: inst = 32'h8220000;
      26220: inst = 32'h10408000;
      26221: inst = 32'hc404723;
      26222: inst = 32'h8220000;
      26223: inst = 32'h10408000;
      26224: inst = 32'hc404724;
      26225: inst = 32'h8220000;
      26226: inst = 32'h10408000;
      26227: inst = 32'hc404725;
      26228: inst = 32'h8220000;
      26229: inst = 32'h10408000;
      26230: inst = 32'hc404726;
      26231: inst = 32'h8220000;
      26232: inst = 32'h10408000;
      26233: inst = 32'hc404727;
      26234: inst = 32'h8220000;
      26235: inst = 32'h10408000;
      26236: inst = 32'hc404728;
      26237: inst = 32'h8220000;
      26238: inst = 32'h10408000;
      26239: inst = 32'hc404729;
      26240: inst = 32'h8220000;
      26241: inst = 32'h10408000;
      26242: inst = 32'hc40472a;
      26243: inst = 32'h8220000;
      26244: inst = 32'h10408000;
      26245: inst = 32'hc40472f;
      26246: inst = 32'h8220000;
      26247: inst = 32'h10408000;
      26248: inst = 32'hc404736;
      26249: inst = 32'h8220000;
      26250: inst = 32'h10408000;
      26251: inst = 32'hc404737;
      26252: inst = 32'h8220000;
      26253: inst = 32'h10408000;
      26254: inst = 32'hc404738;
      26255: inst = 32'h8220000;
      26256: inst = 32'h10408000;
      26257: inst = 32'hc40474c;
      26258: inst = 32'h8220000;
      26259: inst = 32'h10408000;
      26260: inst = 32'hc40474d;
      26261: inst = 32'h8220000;
      26262: inst = 32'h10408000;
      26263: inst = 32'hc40474e;
      26264: inst = 32'h8220000;
      26265: inst = 32'h10408000;
      26266: inst = 32'hc40475d;
      26267: inst = 32'h8220000;
      26268: inst = 32'h10408000;
      26269: inst = 32'hc40475e;
      26270: inst = 32'h8220000;
      26271: inst = 32'h10408000;
      26272: inst = 32'hc40475f;
      26273: inst = 32'h8220000;
      26274: inst = 32'h10408000;
      26275: inst = 32'hc404760;
      26276: inst = 32'h8220000;
      26277: inst = 32'h10408000;
      26278: inst = 32'hc404761;
      26279: inst = 32'h8220000;
      26280: inst = 32'h10408000;
      26281: inst = 32'hc404762;
      26282: inst = 32'h8220000;
      26283: inst = 32'h10408000;
      26284: inst = 32'hc40476e;
      26285: inst = 32'h8220000;
      26286: inst = 32'h10408000;
      26287: inst = 32'hc40476f;
      26288: inst = 32'h8220000;
      26289: inst = 32'h10408000;
      26290: inst = 32'hc404770;
      26291: inst = 32'h8220000;
      26292: inst = 32'h10408000;
      26293: inst = 32'hc4047ac;
      26294: inst = 32'h8220000;
      26295: inst = 32'h10408000;
      26296: inst = 32'hc4047ad;
      26297: inst = 32'h8220000;
      26298: inst = 32'h10408000;
      26299: inst = 32'hc4047ae;
      26300: inst = 32'h8220000;
      26301: inst = 32'h10408000;
      26302: inst = 32'hc4047bd;
      26303: inst = 32'h8220000;
      26304: inst = 32'h10408000;
      26305: inst = 32'hc4047be;
      26306: inst = 32'h8220000;
      26307: inst = 32'h10408000;
      26308: inst = 32'hc4047bf;
      26309: inst = 32'h8220000;
      26310: inst = 32'h10408000;
      26311: inst = 32'hc4047c0;
      26312: inst = 32'h8220000;
      26313: inst = 32'h10408000;
      26314: inst = 32'hc4047c1;
      26315: inst = 32'h8220000;
      26316: inst = 32'h10408000;
      26317: inst = 32'hc4047c2;
      26318: inst = 32'h8220000;
      26319: inst = 32'h10408000;
      26320: inst = 32'hc4047ce;
      26321: inst = 32'h8220000;
      26322: inst = 32'h10408000;
      26323: inst = 32'hc4047cf;
      26324: inst = 32'h8220000;
      26325: inst = 32'h10408000;
      26326: inst = 32'hc4047d0;
      26327: inst = 32'h8220000;
      26328: inst = 32'h10408000;
      26329: inst = 32'hc40480c;
      26330: inst = 32'h8220000;
      26331: inst = 32'h10408000;
      26332: inst = 32'hc40480d;
      26333: inst = 32'h8220000;
      26334: inst = 32'h10408000;
      26335: inst = 32'hc40480e;
      26336: inst = 32'h8220000;
      26337: inst = 32'h10408000;
      26338: inst = 32'hc40481d;
      26339: inst = 32'h8220000;
      26340: inst = 32'h10408000;
      26341: inst = 32'hc40481e;
      26342: inst = 32'h8220000;
      26343: inst = 32'h10408000;
      26344: inst = 32'hc40481f;
      26345: inst = 32'h8220000;
      26346: inst = 32'h10408000;
      26347: inst = 32'hc404820;
      26348: inst = 32'h8220000;
      26349: inst = 32'h10408000;
      26350: inst = 32'hc404821;
      26351: inst = 32'h8220000;
      26352: inst = 32'h10408000;
      26353: inst = 32'hc404822;
      26354: inst = 32'h8220000;
      26355: inst = 32'h10408000;
      26356: inst = 32'hc40482e;
      26357: inst = 32'h8220000;
      26358: inst = 32'h10408000;
      26359: inst = 32'hc40482f;
      26360: inst = 32'h8220000;
      26361: inst = 32'h10408000;
      26362: inst = 32'hc404830;
      26363: inst = 32'h8220000;
      26364: inst = 32'h10408000;
      26365: inst = 32'hc40486c;
      26366: inst = 32'h8220000;
      26367: inst = 32'h10408000;
      26368: inst = 32'hc40486d;
      26369: inst = 32'h8220000;
      26370: inst = 32'h10408000;
      26371: inst = 32'hc40486e;
      26372: inst = 32'h8220000;
      26373: inst = 32'h10408000;
      26374: inst = 32'hc40487d;
      26375: inst = 32'h8220000;
      26376: inst = 32'h10408000;
      26377: inst = 32'hc40487e;
      26378: inst = 32'h8220000;
      26379: inst = 32'h10408000;
      26380: inst = 32'hc40487f;
      26381: inst = 32'h8220000;
      26382: inst = 32'h10408000;
      26383: inst = 32'hc404880;
      26384: inst = 32'h8220000;
      26385: inst = 32'h10408000;
      26386: inst = 32'hc404881;
      26387: inst = 32'h8220000;
      26388: inst = 32'h10408000;
      26389: inst = 32'hc404882;
      26390: inst = 32'h8220000;
      26391: inst = 32'h10408000;
      26392: inst = 32'hc40488e;
      26393: inst = 32'h8220000;
      26394: inst = 32'h10408000;
      26395: inst = 32'hc40488f;
      26396: inst = 32'h8220000;
      26397: inst = 32'h10408000;
      26398: inst = 32'hc404890;
      26399: inst = 32'h8220000;
      26400: inst = 32'h10408000;
      26401: inst = 32'hc4048cc;
      26402: inst = 32'h8220000;
      26403: inst = 32'h10408000;
      26404: inst = 32'hc4048cd;
      26405: inst = 32'h8220000;
      26406: inst = 32'h10408000;
      26407: inst = 32'hc4048ce;
      26408: inst = 32'h8220000;
      26409: inst = 32'h10408000;
      26410: inst = 32'hc4048dd;
      26411: inst = 32'h8220000;
      26412: inst = 32'h10408000;
      26413: inst = 32'hc4048de;
      26414: inst = 32'h8220000;
      26415: inst = 32'h10408000;
      26416: inst = 32'hc4048df;
      26417: inst = 32'h8220000;
      26418: inst = 32'h10408000;
      26419: inst = 32'hc4048e0;
      26420: inst = 32'h8220000;
      26421: inst = 32'h10408000;
      26422: inst = 32'hc4048e1;
      26423: inst = 32'h8220000;
      26424: inst = 32'h10408000;
      26425: inst = 32'hc4048e2;
      26426: inst = 32'h8220000;
      26427: inst = 32'h10408000;
      26428: inst = 32'hc4048ee;
      26429: inst = 32'h8220000;
      26430: inst = 32'h10408000;
      26431: inst = 32'hc4048ef;
      26432: inst = 32'h8220000;
      26433: inst = 32'h10408000;
      26434: inst = 32'hc4048f0;
      26435: inst = 32'h8220000;
      26436: inst = 32'h10408000;
      26437: inst = 32'hc40492c;
      26438: inst = 32'h8220000;
      26439: inst = 32'h10408000;
      26440: inst = 32'hc40492d;
      26441: inst = 32'h8220000;
      26442: inst = 32'h10408000;
      26443: inst = 32'hc40492e;
      26444: inst = 32'h8220000;
      26445: inst = 32'h10408000;
      26446: inst = 32'hc40493d;
      26447: inst = 32'h8220000;
      26448: inst = 32'h10408000;
      26449: inst = 32'hc40493e;
      26450: inst = 32'h8220000;
      26451: inst = 32'h10408000;
      26452: inst = 32'hc40493f;
      26453: inst = 32'h8220000;
      26454: inst = 32'h10408000;
      26455: inst = 32'hc404940;
      26456: inst = 32'h8220000;
      26457: inst = 32'h10408000;
      26458: inst = 32'hc404941;
      26459: inst = 32'h8220000;
      26460: inst = 32'h10408000;
      26461: inst = 32'hc404942;
      26462: inst = 32'h8220000;
      26463: inst = 32'h10408000;
      26464: inst = 32'hc40494e;
      26465: inst = 32'h8220000;
      26466: inst = 32'h10408000;
      26467: inst = 32'hc40494f;
      26468: inst = 32'h8220000;
      26469: inst = 32'h10408000;
      26470: inst = 32'hc404950;
      26471: inst = 32'h8220000;
      26472: inst = 32'h10408000;
      26473: inst = 32'hc404986;
      26474: inst = 32'h8220000;
      26475: inst = 32'h10408000;
      26476: inst = 32'hc404987;
      26477: inst = 32'h8220000;
      26478: inst = 32'h10408000;
      26479: inst = 32'hc404988;
      26480: inst = 32'h8220000;
      26481: inst = 32'h10408000;
      26482: inst = 32'hc404989;
      26483: inst = 32'h8220000;
      26484: inst = 32'h10408000;
      26485: inst = 32'hc40498a;
      26486: inst = 32'h8220000;
      26487: inst = 32'h10408000;
      26488: inst = 32'hc40498b;
      26489: inst = 32'h8220000;
      26490: inst = 32'h10408000;
      26491: inst = 32'hc40498c;
      26492: inst = 32'h8220000;
      26493: inst = 32'h10408000;
      26494: inst = 32'hc40498d;
      26495: inst = 32'h8220000;
      26496: inst = 32'h10408000;
      26497: inst = 32'hc40498e;
      26498: inst = 32'h8220000;
      26499: inst = 32'h10408000;
      26500: inst = 32'hc40499d;
      26501: inst = 32'h8220000;
      26502: inst = 32'h10408000;
      26503: inst = 32'hc40499e;
      26504: inst = 32'h8220000;
      26505: inst = 32'h10408000;
      26506: inst = 32'hc40499f;
      26507: inst = 32'h8220000;
      26508: inst = 32'h10408000;
      26509: inst = 32'hc4049a0;
      26510: inst = 32'h8220000;
      26511: inst = 32'h10408000;
      26512: inst = 32'hc4049a1;
      26513: inst = 32'h8220000;
      26514: inst = 32'h10408000;
      26515: inst = 32'hc4049a2;
      26516: inst = 32'h8220000;
      26517: inst = 32'h10408000;
      26518: inst = 32'hc4049ae;
      26519: inst = 32'h8220000;
      26520: inst = 32'h10408000;
      26521: inst = 32'hc4049af;
      26522: inst = 32'h8220000;
      26523: inst = 32'h10408000;
      26524: inst = 32'hc4049b0;
      26525: inst = 32'h8220000;
      26526: inst = 32'h10408000;
      26527: inst = 32'hc4049e6;
      26528: inst = 32'h8220000;
      26529: inst = 32'h10408000;
      26530: inst = 32'hc4049e7;
      26531: inst = 32'h8220000;
      26532: inst = 32'h10408000;
      26533: inst = 32'hc4049e8;
      26534: inst = 32'h8220000;
      26535: inst = 32'h10408000;
      26536: inst = 32'hc4049e9;
      26537: inst = 32'h8220000;
      26538: inst = 32'h10408000;
      26539: inst = 32'hc4049ea;
      26540: inst = 32'h8220000;
      26541: inst = 32'h10408000;
      26542: inst = 32'hc4049eb;
      26543: inst = 32'h8220000;
      26544: inst = 32'h10408000;
      26545: inst = 32'hc4049ec;
      26546: inst = 32'h8220000;
      26547: inst = 32'h10408000;
      26548: inst = 32'hc4049ed;
      26549: inst = 32'h8220000;
      26550: inst = 32'h10408000;
      26551: inst = 32'hc4049ee;
      26552: inst = 32'h8220000;
      26553: inst = 32'h10408000;
      26554: inst = 32'hc4049fd;
      26555: inst = 32'h8220000;
      26556: inst = 32'h10408000;
      26557: inst = 32'hc4049fe;
      26558: inst = 32'h8220000;
      26559: inst = 32'h10408000;
      26560: inst = 32'hc4049ff;
      26561: inst = 32'h8220000;
      26562: inst = 32'h10408000;
      26563: inst = 32'hc404a00;
      26564: inst = 32'h8220000;
      26565: inst = 32'h10408000;
      26566: inst = 32'hc404a01;
      26567: inst = 32'h8220000;
      26568: inst = 32'h10408000;
      26569: inst = 32'hc404a02;
      26570: inst = 32'h8220000;
      26571: inst = 32'h10408000;
      26572: inst = 32'hc404a0e;
      26573: inst = 32'h8220000;
      26574: inst = 32'h10408000;
      26575: inst = 32'hc404a0f;
      26576: inst = 32'h8220000;
      26577: inst = 32'h10408000;
      26578: inst = 32'hc404a10;
      26579: inst = 32'h8220000;
      26580: inst = 32'h10408000;
      26581: inst = 32'hc404a46;
      26582: inst = 32'h8220000;
      26583: inst = 32'h10408000;
      26584: inst = 32'hc404a47;
      26585: inst = 32'h8220000;
      26586: inst = 32'h10408000;
      26587: inst = 32'hc404a48;
      26588: inst = 32'h8220000;
      26589: inst = 32'h10408000;
      26590: inst = 32'hc404a49;
      26591: inst = 32'h8220000;
      26592: inst = 32'h10408000;
      26593: inst = 32'hc404a4a;
      26594: inst = 32'h8220000;
      26595: inst = 32'h10408000;
      26596: inst = 32'hc404a4b;
      26597: inst = 32'h8220000;
      26598: inst = 32'h10408000;
      26599: inst = 32'hc404a4c;
      26600: inst = 32'h8220000;
      26601: inst = 32'h10408000;
      26602: inst = 32'hc404a4d;
      26603: inst = 32'h8220000;
      26604: inst = 32'h10408000;
      26605: inst = 32'hc404a4e;
      26606: inst = 32'h8220000;
      26607: inst = 32'h10408000;
      26608: inst = 32'hc404a5d;
      26609: inst = 32'h8220000;
      26610: inst = 32'h10408000;
      26611: inst = 32'hc404a5e;
      26612: inst = 32'h8220000;
      26613: inst = 32'h10408000;
      26614: inst = 32'hc404a5f;
      26615: inst = 32'h8220000;
      26616: inst = 32'h10408000;
      26617: inst = 32'hc404a60;
      26618: inst = 32'h8220000;
      26619: inst = 32'h10408000;
      26620: inst = 32'hc404a61;
      26621: inst = 32'h8220000;
      26622: inst = 32'h10408000;
      26623: inst = 32'hc404a62;
      26624: inst = 32'h8220000;
      26625: inst = 32'h10408000;
      26626: inst = 32'hc404a6e;
      26627: inst = 32'h8220000;
      26628: inst = 32'h10408000;
      26629: inst = 32'hc404a6f;
      26630: inst = 32'h8220000;
      26631: inst = 32'h10408000;
      26632: inst = 32'hc404a70;
      26633: inst = 32'h8220000;
      26634: inst = 32'h10408000;
      26635: inst = 32'hc404abd;
      26636: inst = 32'h8220000;
      26637: inst = 32'h10408000;
      26638: inst = 32'hc404abe;
      26639: inst = 32'h8220000;
      26640: inst = 32'h10408000;
      26641: inst = 32'hc404abf;
      26642: inst = 32'h8220000;
      26643: inst = 32'h10408000;
      26644: inst = 32'hc404ac0;
      26645: inst = 32'h8220000;
      26646: inst = 32'h10408000;
      26647: inst = 32'hc404ac1;
      26648: inst = 32'h8220000;
      26649: inst = 32'h10408000;
      26650: inst = 32'hc404ac2;
      26651: inst = 32'h8220000;
      26652: inst = 32'h10408000;
      26653: inst = 32'hc404ace;
      26654: inst = 32'h8220000;
      26655: inst = 32'h10408000;
      26656: inst = 32'hc404acf;
      26657: inst = 32'h8220000;
      26658: inst = 32'h10408000;
      26659: inst = 32'hc404ad0;
      26660: inst = 32'h8220000;
      26661: inst = 32'h10408000;
      26662: inst = 32'hc404b1d;
      26663: inst = 32'h8220000;
      26664: inst = 32'h10408000;
      26665: inst = 32'hc404b1e;
      26666: inst = 32'h8220000;
      26667: inst = 32'h10408000;
      26668: inst = 32'hc404b1f;
      26669: inst = 32'h8220000;
      26670: inst = 32'h10408000;
      26671: inst = 32'hc404b20;
      26672: inst = 32'h8220000;
      26673: inst = 32'h10408000;
      26674: inst = 32'hc404b21;
      26675: inst = 32'h8220000;
      26676: inst = 32'h10408000;
      26677: inst = 32'hc404b22;
      26678: inst = 32'h8220000;
      26679: inst = 32'h10408000;
      26680: inst = 32'hc404b23;
      26681: inst = 32'h8220000;
      26682: inst = 32'h10408000;
      26683: inst = 32'hc404b24;
      26684: inst = 32'h8220000;
      26685: inst = 32'h10408000;
      26686: inst = 32'hc404b25;
      26687: inst = 32'h8220000;
      26688: inst = 32'h10408000;
      26689: inst = 32'hc404b26;
      26690: inst = 32'h8220000;
      26691: inst = 32'h10408000;
      26692: inst = 32'hc404b27;
      26693: inst = 32'h8220000;
      26694: inst = 32'h10408000;
      26695: inst = 32'hc404b28;
      26696: inst = 32'h8220000;
      26697: inst = 32'h10408000;
      26698: inst = 32'hc404b29;
      26699: inst = 32'h8220000;
      26700: inst = 32'h10408000;
      26701: inst = 32'hc404b2a;
      26702: inst = 32'h8220000;
      26703: inst = 32'h10408000;
      26704: inst = 32'hc404b2b;
      26705: inst = 32'h8220000;
      26706: inst = 32'h10408000;
      26707: inst = 32'hc404b2c;
      26708: inst = 32'h8220000;
      26709: inst = 32'h10408000;
      26710: inst = 32'hc404b2d;
      26711: inst = 32'h8220000;
      26712: inst = 32'h10408000;
      26713: inst = 32'hc404b2e;
      26714: inst = 32'h8220000;
      26715: inst = 32'h10408000;
      26716: inst = 32'hc404b2f;
      26717: inst = 32'h8220000;
      26718: inst = 32'h10408000;
      26719: inst = 32'hc404b30;
      26720: inst = 32'h8220000;
      26721: inst = 32'h10408000;
      26722: inst = 32'hc404b7d;
      26723: inst = 32'h8220000;
      26724: inst = 32'h10408000;
      26725: inst = 32'hc404b7e;
      26726: inst = 32'h8220000;
      26727: inst = 32'h10408000;
      26728: inst = 32'hc404b7f;
      26729: inst = 32'h8220000;
      26730: inst = 32'h10408000;
      26731: inst = 32'hc404b80;
      26732: inst = 32'h8220000;
      26733: inst = 32'h10408000;
      26734: inst = 32'hc404b81;
      26735: inst = 32'h8220000;
      26736: inst = 32'h10408000;
      26737: inst = 32'hc404b82;
      26738: inst = 32'h8220000;
      26739: inst = 32'h10408000;
      26740: inst = 32'hc404b83;
      26741: inst = 32'h8220000;
      26742: inst = 32'h10408000;
      26743: inst = 32'hc404b84;
      26744: inst = 32'h8220000;
      26745: inst = 32'h10408000;
      26746: inst = 32'hc404b85;
      26747: inst = 32'h8220000;
      26748: inst = 32'h10408000;
      26749: inst = 32'hc404b86;
      26750: inst = 32'h8220000;
      26751: inst = 32'h10408000;
      26752: inst = 32'hc404b87;
      26753: inst = 32'h8220000;
      26754: inst = 32'h10408000;
      26755: inst = 32'hc404b88;
      26756: inst = 32'h8220000;
      26757: inst = 32'h10408000;
      26758: inst = 32'hc404b89;
      26759: inst = 32'h8220000;
      26760: inst = 32'h10408000;
      26761: inst = 32'hc404b8a;
      26762: inst = 32'h8220000;
      26763: inst = 32'h10408000;
      26764: inst = 32'hc404b8b;
      26765: inst = 32'h8220000;
      26766: inst = 32'h10408000;
      26767: inst = 32'hc404b8c;
      26768: inst = 32'h8220000;
      26769: inst = 32'h10408000;
      26770: inst = 32'hc404b8d;
      26771: inst = 32'h8220000;
      26772: inst = 32'h10408000;
      26773: inst = 32'hc404b8e;
      26774: inst = 32'h8220000;
      26775: inst = 32'h10408000;
      26776: inst = 32'hc404b8f;
      26777: inst = 32'h8220000;
      26778: inst = 32'h10408000;
      26779: inst = 32'hc404b90;
      26780: inst = 32'h8220000;
      26781: inst = 32'h10408000;
      26782: inst = 32'hc404bdd;
      26783: inst = 32'h8220000;
      26784: inst = 32'h10408000;
      26785: inst = 32'hc404bde;
      26786: inst = 32'h8220000;
      26787: inst = 32'h10408000;
      26788: inst = 32'hc404bdf;
      26789: inst = 32'h8220000;
      26790: inst = 32'h10408000;
      26791: inst = 32'hc404be0;
      26792: inst = 32'h8220000;
      26793: inst = 32'h10408000;
      26794: inst = 32'hc404be1;
      26795: inst = 32'h8220000;
      26796: inst = 32'h10408000;
      26797: inst = 32'hc404be2;
      26798: inst = 32'h8220000;
      26799: inst = 32'h10408000;
      26800: inst = 32'hc404be3;
      26801: inst = 32'h8220000;
      26802: inst = 32'h10408000;
      26803: inst = 32'hc404be4;
      26804: inst = 32'h8220000;
      26805: inst = 32'h10408000;
      26806: inst = 32'hc404be5;
      26807: inst = 32'h8220000;
      26808: inst = 32'h10408000;
      26809: inst = 32'hc404be6;
      26810: inst = 32'h8220000;
      26811: inst = 32'h10408000;
      26812: inst = 32'hc404be7;
      26813: inst = 32'h8220000;
      26814: inst = 32'h10408000;
      26815: inst = 32'hc404be8;
      26816: inst = 32'h8220000;
      26817: inst = 32'h10408000;
      26818: inst = 32'hc404be9;
      26819: inst = 32'h8220000;
      26820: inst = 32'h10408000;
      26821: inst = 32'hc404bea;
      26822: inst = 32'h8220000;
      26823: inst = 32'h10408000;
      26824: inst = 32'hc404beb;
      26825: inst = 32'h8220000;
      26826: inst = 32'h10408000;
      26827: inst = 32'hc404bec;
      26828: inst = 32'h8220000;
      26829: inst = 32'h10408000;
      26830: inst = 32'hc404bed;
      26831: inst = 32'h8220000;
      26832: inst = 32'h10408000;
      26833: inst = 32'hc404bee;
      26834: inst = 32'h8220000;
      26835: inst = 32'h10408000;
      26836: inst = 32'hc404bef;
      26837: inst = 32'h8220000;
      26838: inst = 32'h10408000;
      26839: inst = 32'hc404bf0;
      26840: inst = 32'h8220000;
      26841: inst = 32'h10408000;
      26842: inst = 32'hc404c3d;
      26843: inst = 32'h8220000;
      26844: inst = 32'h10408000;
      26845: inst = 32'hc404c3e;
      26846: inst = 32'h8220000;
      26847: inst = 32'h10408000;
      26848: inst = 32'hc404c3f;
      26849: inst = 32'h8220000;
      26850: inst = 32'h10408000;
      26851: inst = 32'hc404c40;
      26852: inst = 32'h8220000;
      26853: inst = 32'h10408000;
      26854: inst = 32'hc404c41;
      26855: inst = 32'h8220000;
      26856: inst = 32'h10408000;
      26857: inst = 32'hc404c42;
      26858: inst = 32'h8220000;
      26859: inst = 32'h10408000;
      26860: inst = 32'hc404c9d;
      26861: inst = 32'h8220000;
      26862: inst = 32'h10408000;
      26863: inst = 32'hc404c9e;
      26864: inst = 32'h8220000;
      26865: inst = 32'h10408000;
      26866: inst = 32'hc404c9f;
      26867: inst = 32'h8220000;
      26868: inst = 32'h10408000;
      26869: inst = 32'hc404ca0;
      26870: inst = 32'h8220000;
      26871: inst = 32'h10408000;
      26872: inst = 32'hc404ca1;
      26873: inst = 32'h8220000;
      26874: inst = 32'h10408000;
      26875: inst = 32'hc404ca2;
      26876: inst = 32'h8220000;
      26877: inst = 32'h10408000;
      26878: inst = 32'hc404cfd;
      26879: inst = 32'h8220000;
      26880: inst = 32'h10408000;
      26881: inst = 32'hc404cfe;
      26882: inst = 32'h8220000;
      26883: inst = 32'h10408000;
      26884: inst = 32'hc404cff;
      26885: inst = 32'h8220000;
      26886: inst = 32'h10408000;
      26887: inst = 32'hc404d00;
      26888: inst = 32'h8220000;
      26889: inst = 32'h10408000;
      26890: inst = 32'hc404d01;
      26891: inst = 32'h8220000;
      26892: inst = 32'h10408000;
      26893: inst = 32'hc404d02;
      26894: inst = 32'h8220000;
      26895: inst = 32'h10408000;
      26896: inst = 32'hc404d25;
      26897: inst = 32'h8220000;
      26898: inst = 32'h10408000;
      26899: inst = 32'hc404d26;
      26900: inst = 32'h8220000;
      26901: inst = 32'h10408000;
      26902: inst = 32'hc404d27;
      26903: inst = 32'h8220000;
      26904: inst = 32'h10408000;
      26905: inst = 32'hc404d28;
      26906: inst = 32'h8220000;
      26907: inst = 32'h10408000;
      26908: inst = 32'hc404d29;
      26909: inst = 32'h8220000;
      26910: inst = 32'h10408000;
      26911: inst = 32'hc404d2a;
      26912: inst = 32'h8220000;
      26913: inst = 32'h10408000;
      26914: inst = 32'hc404d2b;
      26915: inst = 32'h8220000;
      26916: inst = 32'h10408000;
      26917: inst = 32'hc404d2c;
      26918: inst = 32'h8220000;
      26919: inst = 32'h10408000;
      26920: inst = 32'hc404d2d;
      26921: inst = 32'h8220000;
      26922: inst = 32'h10408000;
      26923: inst = 32'hc404d2e;
      26924: inst = 32'h8220000;
      26925: inst = 32'h10408000;
      26926: inst = 32'hc404d2f;
      26927: inst = 32'h8220000;
      26928: inst = 32'h10408000;
      26929: inst = 32'hc404d30;
      26930: inst = 32'h8220000;
      26931: inst = 32'h10408000;
      26932: inst = 32'hc404d31;
      26933: inst = 32'h8220000;
      26934: inst = 32'h10408000;
      26935: inst = 32'hc404d32;
      26936: inst = 32'h8220000;
      26937: inst = 32'h10408000;
      26938: inst = 32'hc404d33;
      26939: inst = 32'h8220000;
      26940: inst = 32'h10408000;
      26941: inst = 32'hc404d34;
      26942: inst = 32'h8220000;
      26943: inst = 32'h10408000;
      26944: inst = 32'hc404d35;
      26945: inst = 32'h8220000;
      26946: inst = 32'h10408000;
      26947: inst = 32'hc404d36;
      26948: inst = 32'h8220000;
      26949: inst = 32'h10408000;
      26950: inst = 32'hc404d37;
      26951: inst = 32'h8220000;
      26952: inst = 32'h10408000;
      26953: inst = 32'hc404d38;
      26954: inst = 32'h8220000;
      26955: inst = 32'h10408000;
      26956: inst = 32'hc404d39;
      26957: inst = 32'h8220000;
      26958: inst = 32'h10408000;
      26959: inst = 32'hc404d3a;
      26960: inst = 32'h8220000;
      26961: inst = 32'h10408000;
      26962: inst = 32'hc404d5d;
      26963: inst = 32'h8220000;
      26964: inst = 32'h10408000;
      26965: inst = 32'hc404d5e;
      26966: inst = 32'h8220000;
      26967: inst = 32'h10408000;
      26968: inst = 32'hc404d5f;
      26969: inst = 32'h8220000;
      26970: inst = 32'h10408000;
      26971: inst = 32'hc404d60;
      26972: inst = 32'h8220000;
      26973: inst = 32'h10408000;
      26974: inst = 32'hc404d61;
      26975: inst = 32'h8220000;
      26976: inst = 32'h10408000;
      26977: inst = 32'hc404d62;
      26978: inst = 32'h8220000;
      26979: inst = 32'h10408000;
      26980: inst = 32'hc404d85;
      26981: inst = 32'h8220000;
      26982: inst = 32'h10408000;
      26983: inst = 32'hc404d86;
      26984: inst = 32'h8220000;
      26985: inst = 32'h10408000;
      26986: inst = 32'hc404d87;
      26987: inst = 32'h8220000;
      26988: inst = 32'h10408000;
      26989: inst = 32'hc404d88;
      26990: inst = 32'h8220000;
      26991: inst = 32'h10408000;
      26992: inst = 32'hc404d89;
      26993: inst = 32'h8220000;
      26994: inst = 32'h10408000;
      26995: inst = 32'hc404d8a;
      26996: inst = 32'h8220000;
      26997: inst = 32'h10408000;
      26998: inst = 32'hc404d8b;
      26999: inst = 32'h8220000;
      27000: inst = 32'h10408000;
      27001: inst = 32'hc404d8c;
      27002: inst = 32'h8220000;
      27003: inst = 32'h10408000;
      27004: inst = 32'hc404d8d;
      27005: inst = 32'h8220000;
      27006: inst = 32'h10408000;
      27007: inst = 32'hc404d8e;
      27008: inst = 32'h8220000;
      27009: inst = 32'h10408000;
      27010: inst = 32'hc404d8f;
      27011: inst = 32'h8220000;
      27012: inst = 32'h10408000;
      27013: inst = 32'hc404d90;
      27014: inst = 32'h8220000;
      27015: inst = 32'h10408000;
      27016: inst = 32'hc404d91;
      27017: inst = 32'h8220000;
      27018: inst = 32'h10408000;
      27019: inst = 32'hc404d92;
      27020: inst = 32'h8220000;
      27021: inst = 32'h10408000;
      27022: inst = 32'hc404d93;
      27023: inst = 32'h8220000;
      27024: inst = 32'h10408000;
      27025: inst = 32'hc404d94;
      27026: inst = 32'h8220000;
      27027: inst = 32'h10408000;
      27028: inst = 32'hc404d95;
      27029: inst = 32'h8220000;
      27030: inst = 32'h10408000;
      27031: inst = 32'hc404d96;
      27032: inst = 32'h8220000;
      27033: inst = 32'h10408000;
      27034: inst = 32'hc404d97;
      27035: inst = 32'h8220000;
      27036: inst = 32'h10408000;
      27037: inst = 32'hc404d98;
      27038: inst = 32'h8220000;
      27039: inst = 32'h10408000;
      27040: inst = 32'hc404d99;
      27041: inst = 32'h8220000;
      27042: inst = 32'h10408000;
      27043: inst = 32'hc404d9a;
      27044: inst = 32'h8220000;
      27045: inst = 32'h10408000;
      27046: inst = 32'hc404dbd;
      27047: inst = 32'h8220000;
      27048: inst = 32'h10408000;
      27049: inst = 32'hc404dbe;
      27050: inst = 32'h8220000;
      27051: inst = 32'h10408000;
      27052: inst = 32'hc404dbf;
      27053: inst = 32'h8220000;
      27054: inst = 32'h10408000;
      27055: inst = 32'hc404dc0;
      27056: inst = 32'h8220000;
      27057: inst = 32'h10408000;
      27058: inst = 32'hc404dc1;
      27059: inst = 32'h8220000;
      27060: inst = 32'h10408000;
      27061: inst = 32'hc404dc2;
      27062: inst = 32'h8220000;
      27063: inst = 32'h10408000;
      27064: inst = 32'hc404de5;
      27065: inst = 32'h8220000;
      27066: inst = 32'h10408000;
      27067: inst = 32'hc404de6;
      27068: inst = 32'h8220000;
      27069: inst = 32'h10408000;
      27070: inst = 32'hc404de7;
      27071: inst = 32'h8220000;
      27072: inst = 32'h10408000;
      27073: inst = 32'hc404de8;
      27074: inst = 32'h8220000;
      27075: inst = 32'h10408000;
      27076: inst = 32'hc404de9;
      27077: inst = 32'h8220000;
      27078: inst = 32'h10408000;
      27079: inst = 32'hc404dea;
      27080: inst = 32'h8220000;
      27081: inst = 32'h10408000;
      27082: inst = 32'hc404deb;
      27083: inst = 32'h8220000;
      27084: inst = 32'h10408000;
      27085: inst = 32'hc404dec;
      27086: inst = 32'h8220000;
      27087: inst = 32'h10408000;
      27088: inst = 32'hc404ded;
      27089: inst = 32'h8220000;
      27090: inst = 32'h10408000;
      27091: inst = 32'hc404dee;
      27092: inst = 32'h8220000;
      27093: inst = 32'h10408000;
      27094: inst = 32'hc404def;
      27095: inst = 32'h8220000;
      27096: inst = 32'h10408000;
      27097: inst = 32'hc404df0;
      27098: inst = 32'h8220000;
      27099: inst = 32'h10408000;
      27100: inst = 32'hc404df1;
      27101: inst = 32'h8220000;
      27102: inst = 32'h10408000;
      27103: inst = 32'hc404df2;
      27104: inst = 32'h8220000;
      27105: inst = 32'h10408000;
      27106: inst = 32'hc404df3;
      27107: inst = 32'h8220000;
      27108: inst = 32'h10408000;
      27109: inst = 32'hc404df4;
      27110: inst = 32'h8220000;
      27111: inst = 32'h10408000;
      27112: inst = 32'hc404df5;
      27113: inst = 32'h8220000;
      27114: inst = 32'h10408000;
      27115: inst = 32'hc404df6;
      27116: inst = 32'h8220000;
      27117: inst = 32'h10408000;
      27118: inst = 32'hc404df7;
      27119: inst = 32'h8220000;
      27120: inst = 32'h10408000;
      27121: inst = 32'hc404df8;
      27122: inst = 32'h8220000;
      27123: inst = 32'h10408000;
      27124: inst = 32'hc404df9;
      27125: inst = 32'h8220000;
      27126: inst = 32'h10408000;
      27127: inst = 32'hc404dfa;
      27128: inst = 32'h8220000;
      27129: inst = 32'h10408000;
      27130: inst = 32'hc404e1d;
      27131: inst = 32'h8220000;
      27132: inst = 32'h10408000;
      27133: inst = 32'hc404e1e;
      27134: inst = 32'h8220000;
      27135: inst = 32'h10408000;
      27136: inst = 32'hc404e1f;
      27137: inst = 32'h8220000;
      27138: inst = 32'h10408000;
      27139: inst = 32'hc404e20;
      27140: inst = 32'h8220000;
      27141: inst = 32'h10408000;
      27142: inst = 32'hc404e21;
      27143: inst = 32'h8220000;
      27144: inst = 32'h10408000;
      27145: inst = 32'hc404e22;
      27146: inst = 32'h8220000;
      27147: inst = 32'h10408000;
      27148: inst = 32'hc404e58;
      27149: inst = 32'h8220000;
      27150: inst = 32'h10408000;
      27151: inst = 32'hc404e59;
      27152: inst = 32'h8220000;
      27153: inst = 32'h10408000;
      27154: inst = 32'hc404e5a;
      27155: inst = 32'h8220000;
      27156: inst = 32'h10408000;
      27157: inst = 32'hc404e7d;
      27158: inst = 32'h8220000;
      27159: inst = 32'h10408000;
      27160: inst = 32'hc404e7e;
      27161: inst = 32'h8220000;
      27162: inst = 32'h10408000;
      27163: inst = 32'hc404e7f;
      27164: inst = 32'h8220000;
      27165: inst = 32'h10408000;
      27166: inst = 32'hc404e80;
      27167: inst = 32'h8220000;
      27168: inst = 32'h10408000;
      27169: inst = 32'hc404e81;
      27170: inst = 32'h8220000;
      27171: inst = 32'h10408000;
      27172: inst = 32'hc404e82;
      27173: inst = 32'h8220000;
      27174: inst = 32'h10408000;
      27175: inst = 32'hc404eb8;
      27176: inst = 32'h8220000;
      27177: inst = 32'h10408000;
      27178: inst = 32'hc404eb9;
      27179: inst = 32'h8220000;
      27180: inst = 32'h10408000;
      27181: inst = 32'hc404eba;
      27182: inst = 32'h8220000;
      27183: inst = 32'h10408000;
      27184: inst = 32'hc404edd;
      27185: inst = 32'h8220000;
      27186: inst = 32'h10408000;
      27187: inst = 32'hc404ede;
      27188: inst = 32'h8220000;
      27189: inst = 32'h10408000;
      27190: inst = 32'hc404edf;
      27191: inst = 32'h8220000;
      27192: inst = 32'h10408000;
      27193: inst = 32'hc404ee0;
      27194: inst = 32'h8220000;
      27195: inst = 32'h10408000;
      27196: inst = 32'hc404ee1;
      27197: inst = 32'h8220000;
      27198: inst = 32'h10408000;
      27199: inst = 32'hc404ee2;
      27200: inst = 32'h8220000;
      27201: inst = 32'h10408000;
      27202: inst = 32'hc404f18;
      27203: inst = 32'h8220000;
      27204: inst = 32'h10408000;
      27205: inst = 32'hc404f19;
      27206: inst = 32'h8220000;
      27207: inst = 32'h10408000;
      27208: inst = 32'hc404f1a;
      27209: inst = 32'h8220000;
      27210: inst = 32'h10408000;
      27211: inst = 32'hc404f3d;
      27212: inst = 32'h8220000;
      27213: inst = 32'h10408000;
      27214: inst = 32'hc404f3e;
      27215: inst = 32'h8220000;
      27216: inst = 32'h10408000;
      27217: inst = 32'hc404f3f;
      27218: inst = 32'h8220000;
      27219: inst = 32'h10408000;
      27220: inst = 32'hc404f40;
      27221: inst = 32'h8220000;
      27222: inst = 32'h10408000;
      27223: inst = 32'hc404f41;
      27224: inst = 32'h8220000;
      27225: inst = 32'h10408000;
      27226: inst = 32'hc404f42;
      27227: inst = 32'h8220000;
      27228: inst = 32'h10408000;
      27229: inst = 32'hc404f78;
      27230: inst = 32'h8220000;
      27231: inst = 32'h10408000;
      27232: inst = 32'hc404f79;
      27233: inst = 32'h8220000;
      27234: inst = 32'h10408000;
      27235: inst = 32'hc404f7a;
      27236: inst = 32'h8220000;
      27237: inst = 32'h10408000;
      27238: inst = 32'hc404f9d;
      27239: inst = 32'h8220000;
      27240: inst = 32'h10408000;
      27241: inst = 32'hc404f9e;
      27242: inst = 32'h8220000;
      27243: inst = 32'h10408000;
      27244: inst = 32'hc404f9f;
      27245: inst = 32'h8220000;
      27246: inst = 32'h10408000;
      27247: inst = 32'hc404fa0;
      27248: inst = 32'h8220000;
      27249: inst = 32'h10408000;
      27250: inst = 32'hc404fa1;
      27251: inst = 32'h8220000;
      27252: inst = 32'h10408000;
      27253: inst = 32'hc404fa2;
      27254: inst = 32'h8220000;
      27255: inst = 32'h10408000;
      27256: inst = 32'hc404fd8;
      27257: inst = 32'h8220000;
      27258: inst = 32'h10408000;
      27259: inst = 32'hc404fd9;
      27260: inst = 32'h8220000;
      27261: inst = 32'h10408000;
      27262: inst = 32'hc404fda;
      27263: inst = 32'h8220000;
      27264: inst = 32'h10408000;
      27265: inst = 32'hc404ffd;
      27266: inst = 32'h8220000;
      27267: inst = 32'h10408000;
      27268: inst = 32'hc404ffe;
      27269: inst = 32'h8220000;
      27270: inst = 32'h10408000;
      27271: inst = 32'hc404fff;
      27272: inst = 32'h8220000;
      27273: inst = 32'h10408000;
      27274: inst = 32'hc405000;
      27275: inst = 32'h8220000;
      27276: inst = 32'h10408000;
      27277: inst = 32'hc405001;
      27278: inst = 32'h8220000;
      27279: inst = 32'h10408000;
      27280: inst = 32'hc405002;
      27281: inst = 32'h8220000;
      27282: inst = 32'h10408000;
      27283: inst = 32'hc405038;
      27284: inst = 32'h8220000;
      27285: inst = 32'h10408000;
      27286: inst = 32'hc405039;
      27287: inst = 32'h8220000;
      27288: inst = 32'h10408000;
      27289: inst = 32'hc40503a;
      27290: inst = 32'h8220000;
      27291: inst = 32'h10408000;
      27292: inst = 32'hc40505d;
      27293: inst = 32'h8220000;
      27294: inst = 32'h10408000;
      27295: inst = 32'hc40505e;
      27296: inst = 32'h8220000;
      27297: inst = 32'h10408000;
      27298: inst = 32'hc40505f;
      27299: inst = 32'h8220000;
      27300: inst = 32'h10408000;
      27301: inst = 32'hc405060;
      27302: inst = 32'h8220000;
      27303: inst = 32'h10408000;
      27304: inst = 32'hc405061;
      27305: inst = 32'h8220000;
      27306: inst = 32'h10408000;
      27307: inst = 32'hc405062;
      27308: inst = 32'h8220000;
      27309: inst = 32'h10408000;
      27310: inst = 32'hc405098;
      27311: inst = 32'h8220000;
      27312: inst = 32'h10408000;
      27313: inst = 32'hc405099;
      27314: inst = 32'h8220000;
      27315: inst = 32'h10408000;
      27316: inst = 32'hc40509a;
      27317: inst = 32'h8220000;
      27318: inst = 32'h10408000;
      27319: inst = 32'hc40509b;
      27320: inst = 32'h8220000;
      27321: inst = 32'h10408000;
      27322: inst = 32'hc40509c;
      27323: inst = 32'h8220000;
      27324: inst = 32'h10408000;
      27325: inst = 32'hc40509d;
      27326: inst = 32'h8220000;
      27327: inst = 32'h10408000;
      27328: inst = 32'hc40509e;
      27329: inst = 32'h8220000;
      27330: inst = 32'h10408000;
      27331: inst = 32'hc40509f;
      27332: inst = 32'h8220000;
      27333: inst = 32'h10408000;
      27334: inst = 32'hc4050a0;
      27335: inst = 32'h8220000;
      27336: inst = 32'h10408000;
      27337: inst = 32'hc4050a1;
      27338: inst = 32'h8220000;
      27339: inst = 32'h10408000;
      27340: inst = 32'hc4050a2;
      27341: inst = 32'h8220000;
      27342: inst = 32'h10408000;
      27343: inst = 32'hc4050a3;
      27344: inst = 32'h8220000;
      27345: inst = 32'h10408000;
      27346: inst = 32'hc4050a4;
      27347: inst = 32'h8220000;
      27348: inst = 32'h10408000;
      27349: inst = 32'hc4050a5;
      27350: inst = 32'h8220000;
      27351: inst = 32'h10408000;
      27352: inst = 32'hc4050a6;
      27353: inst = 32'h8220000;
      27354: inst = 32'h10408000;
      27355: inst = 32'hc4050a7;
      27356: inst = 32'h8220000;
      27357: inst = 32'h10408000;
      27358: inst = 32'hc4050a8;
      27359: inst = 32'h8220000;
      27360: inst = 32'h10408000;
      27361: inst = 32'hc4050a9;
      27362: inst = 32'h8220000;
      27363: inst = 32'h10408000;
      27364: inst = 32'hc4050aa;
      27365: inst = 32'h8220000;
      27366: inst = 32'h10408000;
      27367: inst = 32'hc4050ab;
      27368: inst = 32'h8220000;
      27369: inst = 32'h10408000;
      27370: inst = 32'hc4050ac;
      27371: inst = 32'h8220000;
      27372: inst = 32'h10408000;
      27373: inst = 32'hc4050ad;
      27374: inst = 32'h8220000;
      27375: inst = 32'h10408000;
      27376: inst = 32'hc4050ae;
      27377: inst = 32'h8220000;
      27378: inst = 32'h10408000;
      27379: inst = 32'hc4050af;
      27380: inst = 32'h8220000;
      27381: inst = 32'h10408000;
      27382: inst = 32'hc4050b0;
      27383: inst = 32'h8220000;
      27384: inst = 32'h10408000;
      27385: inst = 32'hc4050b1;
      27386: inst = 32'h8220000;
      27387: inst = 32'h10408000;
      27388: inst = 32'hc4050b2;
      27389: inst = 32'h8220000;
      27390: inst = 32'h10408000;
      27391: inst = 32'hc4050b3;
      27392: inst = 32'h8220000;
      27393: inst = 32'h10408000;
      27394: inst = 32'hc4050b4;
      27395: inst = 32'h8220000;
      27396: inst = 32'h10408000;
      27397: inst = 32'hc4050b5;
      27398: inst = 32'h8220000;
      27399: inst = 32'h10408000;
      27400: inst = 32'hc4050b6;
      27401: inst = 32'h8220000;
      27402: inst = 32'h10408000;
      27403: inst = 32'hc4050b7;
      27404: inst = 32'h8220000;
      27405: inst = 32'h10408000;
      27406: inst = 32'hc4050b8;
      27407: inst = 32'h8220000;
      27408: inst = 32'h10408000;
      27409: inst = 32'hc4050b9;
      27410: inst = 32'h8220000;
      27411: inst = 32'h10408000;
      27412: inst = 32'hc4050ba;
      27413: inst = 32'h8220000;
      27414: inst = 32'h10408000;
      27415: inst = 32'hc4050bb;
      27416: inst = 32'h8220000;
      27417: inst = 32'h10408000;
      27418: inst = 32'hc4050bc;
      27419: inst = 32'h8220000;
      27420: inst = 32'h10408000;
      27421: inst = 32'hc4050bd;
      27422: inst = 32'h8220000;
      27423: inst = 32'h10408000;
      27424: inst = 32'hc4050be;
      27425: inst = 32'h8220000;
      27426: inst = 32'h10408000;
      27427: inst = 32'hc4050bf;
      27428: inst = 32'h8220000;
      27429: inst = 32'h10408000;
      27430: inst = 32'hc4050c0;
      27431: inst = 32'h8220000;
      27432: inst = 32'h10408000;
      27433: inst = 32'hc4050c1;
      27434: inst = 32'h8220000;
      27435: inst = 32'h10408000;
      27436: inst = 32'hc4050c2;
      27437: inst = 32'h8220000;
      27438: inst = 32'h10408000;
      27439: inst = 32'hc4050f8;
      27440: inst = 32'h8220000;
      27441: inst = 32'h10408000;
      27442: inst = 32'hc4050f9;
      27443: inst = 32'h8220000;
      27444: inst = 32'h10408000;
      27445: inst = 32'hc4050fa;
      27446: inst = 32'h8220000;
      27447: inst = 32'h10408000;
      27448: inst = 32'hc4050fb;
      27449: inst = 32'h8220000;
      27450: inst = 32'h10408000;
      27451: inst = 32'hc4050fc;
      27452: inst = 32'h8220000;
      27453: inst = 32'h10408000;
      27454: inst = 32'hc4050fd;
      27455: inst = 32'h8220000;
      27456: inst = 32'h10408000;
      27457: inst = 32'hc4050fe;
      27458: inst = 32'h8220000;
      27459: inst = 32'h10408000;
      27460: inst = 32'hc4050ff;
      27461: inst = 32'h8220000;
      27462: inst = 32'h10408000;
      27463: inst = 32'hc405100;
      27464: inst = 32'h8220000;
      27465: inst = 32'h10408000;
      27466: inst = 32'hc405101;
      27467: inst = 32'h8220000;
      27468: inst = 32'h10408000;
      27469: inst = 32'hc405102;
      27470: inst = 32'h8220000;
      27471: inst = 32'h10408000;
      27472: inst = 32'hc405103;
      27473: inst = 32'h8220000;
      27474: inst = 32'h10408000;
      27475: inst = 32'hc405104;
      27476: inst = 32'h8220000;
      27477: inst = 32'h10408000;
      27478: inst = 32'hc405105;
      27479: inst = 32'h8220000;
      27480: inst = 32'h10408000;
      27481: inst = 32'hc405106;
      27482: inst = 32'h8220000;
      27483: inst = 32'h10408000;
      27484: inst = 32'hc405107;
      27485: inst = 32'h8220000;
      27486: inst = 32'h10408000;
      27487: inst = 32'hc405108;
      27488: inst = 32'h8220000;
      27489: inst = 32'h10408000;
      27490: inst = 32'hc405109;
      27491: inst = 32'h8220000;
      27492: inst = 32'h10408000;
      27493: inst = 32'hc40510a;
      27494: inst = 32'h8220000;
      27495: inst = 32'h10408000;
      27496: inst = 32'hc40510b;
      27497: inst = 32'h8220000;
      27498: inst = 32'h10408000;
      27499: inst = 32'hc40510c;
      27500: inst = 32'h8220000;
      27501: inst = 32'h10408000;
      27502: inst = 32'hc40510d;
      27503: inst = 32'h8220000;
      27504: inst = 32'h10408000;
      27505: inst = 32'hc40510e;
      27506: inst = 32'h8220000;
      27507: inst = 32'h10408000;
      27508: inst = 32'hc40510f;
      27509: inst = 32'h8220000;
      27510: inst = 32'h10408000;
      27511: inst = 32'hc405110;
      27512: inst = 32'h8220000;
      27513: inst = 32'h10408000;
      27514: inst = 32'hc405111;
      27515: inst = 32'h8220000;
      27516: inst = 32'h10408000;
      27517: inst = 32'hc405112;
      27518: inst = 32'h8220000;
      27519: inst = 32'h10408000;
      27520: inst = 32'hc405113;
      27521: inst = 32'h8220000;
      27522: inst = 32'h10408000;
      27523: inst = 32'hc405114;
      27524: inst = 32'h8220000;
      27525: inst = 32'h10408000;
      27526: inst = 32'hc405115;
      27527: inst = 32'h8220000;
      27528: inst = 32'h10408000;
      27529: inst = 32'hc405116;
      27530: inst = 32'h8220000;
      27531: inst = 32'h10408000;
      27532: inst = 32'hc405117;
      27533: inst = 32'h8220000;
      27534: inst = 32'h10408000;
      27535: inst = 32'hc405118;
      27536: inst = 32'h8220000;
      27537: inst = 32'h10408000;
      27538: inst = 32'hc405119;
      27539: inst = 32'h8220000;
      27540: inst = 32'h10408000;
      27541: inst = 32'hc40511a;
      27542: inst = 32'h8220000;
      27543: inst = 32'h10408000;
      27544: inst = 32'hc40511b;
      27545: inst = 32'h8220000;
      27546: inst = 32'h10408000;
      27547: inst = 32'hc40511c;
      27548: inst = 32'h8220000;
      27549: inst = 32'h10408000;
      27550: inst = 32'hc40511d;
      27551: inst = 32'h8220000;
      27552: inst = 32'h10408000;
      27553: inst = 32'hc40511e;
      27554: inst = 32'h8220000;
      27555: inst = 32'h10408000;
      27556: inst = 32'hc40511f;
      27557: inst = 32'h8220000;
      27558: inst = 32'h10408000;
      27559: inst = 32'hc405120;
      27560: inst = 32'h8220000;
      27561: inst = 32'h10408000;
      27562: inst = 32'hc405121;
      27563: inst = 32'h8220000;
      27564: inst = 32'h10408000;
      27565: inst = 32'hc405122;
      27566: inst = 32'h8220000;
      27567: inst = 32'h10408000;
      27568: inst = 32'hc405136;
      27569: inst = 32'h8220000;
      27570: inst = 32'h10408000;
      27571: inst = 32'hc405137;
      27572: inst = 32'h8220000;
      27573: inst = 32'h10408000;
      27574: inst = 32'hc405138;
      27575: inst = 32'h8220000;
      27576: inst = 32'h10408000;
      27577: inst = 32'hc405158;
      27578: inst = 32'h8220000;
      27579: inst = 32'h10408000;
      27580: inst = 32'hc405159;
      27581: inst = 32'h8220000;
      27582: inst = 32'h10408000;
      27583: inst = 32'hc40515a;
      27584: inst = 32'h8220000;
      27585: inst = 32'h10408000;
      27586: inst = 32'hc40515b;
      27587: inst = 32'h8220000;
      27588: inst = 32'h10408000;
      27589: inst = 32'hc40515c;
      27590: inst = 32'h8220000;
      27591: inst = 32'h10408000;
      27592: inst = 32'hc40515d;
      27593: inst = 32'h8220000;
      27594: inst = 32'h10408000;
      27595: inst = 32'hc40515e;
      27596: inst = 32'h8220000;
      27597: inst = 32'h10408000;
      27598: inst = 32'hc40515f;
      27599: inst = 32'h8220000;
      27600: inst = 32'h10408000;
      27601: inst = 32'hc405160;
      27602: inst = 32'h8220000;
      27603: inst = 32'h10408000;
      27604: inst = 32'hc405161;
      27605: inst = 32'h8220000;
      27606: inst = 32'h10408000;
      27607: inst = 32'hc405162;
      27608: inst = 32'h8220000;
      27609: inst = 32'h10408000;
      27610: inst = 32'hc405163;
      27611: inst = 32'h8220000;
      27612: inst = 32'h10408000;
      27613: inst = 32'hc405164;
      27614: inst = 32'h8220000;
      27615: inst = 32'h10408000;
      27616: inst = 32'hc405165;
      27617: inst = 32'h8220000;
      27618: inst = 32'h10408000;
      27619: inst = 32'hc405166;
      27620: inst = 32'h8220000;
      27621: inst = 32'h10408000;
      27622: inst = 32'hc405167;
      27623: inst = 32'h8220000;
      27624: inst = 32'h10408000;
      27625: inst = 32'hc405168;
      27626: inst = 32'h8220000;
      27627: inst = 32'h10408000;
      27628: inst = 32'hc405169;
      27629: inst = 32'h8220000;
      27630: inst = 32'h10408000;
      27631: inst = 32'hc40516a;
      27632: inst = 32'h8220000;
      27633: inst = 32'h10408000;
      27634: inst = 32'hc40516b;
      27635: inst = 32'h8220000;
      27636: inst = 32'h10408000;
      27637: inst = 32'hc40516c;
      27638: inst = 32'h8220000;
      27639: inst = 32'h10408000;
      27640: inst = 32'hc40516d;
      27641: inst = 32'h8220000;
      27642: inst = 32'h10408000;
      27643: inst = 32'hc40516e;
      27644: inst = 32'h8220000;
      27645: inst = 32'h10408000;
      27646: inst = 32'hc40516f;
      27647: inst = 32'h8220000;
      27648: inst = 32'h10408000;
      27649: inst = 32'hc405170;
      27650: inst = 32'h8220000;
      27651: inst = 32'h10408000;
      27652: inst = 32'hc405171;
      27653: inst = 32'h8220000;
      27654: inst = 32'h10408000;
      27655: inst = 32'hc405172;
      27656: inst = 32'h8220000;
      27657: inst = 32'h10408000;
      27658: inst = 32'hc405173;
      27659: inst = 32'h8220000;
      27660: inst = 32'h10408000;
      27661: inst = 32'hc405174;
      27662: inst = 32'h8220000;
      27663: inst = 32'h10408000;
      27664: inst = 32'hc405175;
      27665: inst = 32'h8220000;
      27666: inst = 32'h10408000;
      27667: inst = 32'hc405176;
      27668: inst = 32'h8220000;
      27669: inst = 32'h10408000;
      27670: inst = 32'hc405177;
      27671: inst = 32'h8220000;
      27672: inst = 32'h10408000;
      27673: inst = 32'hc405178;
      27674: inst = 32'h8220000;
      27675: inst = 32'h10408000;
      27676: inst = 32'hc405179;
      27677: inst = 32'h8220000;
      27678: inst = 32'h10408000;
      27679: inst = 32'hc40517a;
      27680: inst = 32'h8220000;
      27681: inst = 32'h10408000;
      27682: inst = 32'hc40517b;
      27683: inst = 32'h8220000;
      27684: inst = 32'h10408000;
      27685: inst = 32'hc40517c;
      27686: inst = 32'h8220000;
      27687: inst = 32'h10408000;
      27688: inst = 32'hc40517d;
      27689: inst = 32'h8220000;
      27690: inst = 32'h10408000;
      27691: inst = 32'hc40517e;
      27692: inst = 32'h8220000;
      27693: inst = 32'h10408000;
      27694: inst = 32'hc40517f;
      27695: inst = 32'h8220000;
      27696: inst = 32'h10408000;
      27697: inst = 32'hc405180;
      27698: inst = 32'h8220000;
      27699: inst = 32'h10408000;
      27700: inst = 32'hc405181;
      27701: inst = 32'h8220000;
      27702: inst = 32'h10408000;
      27703: inst = 32'hc405182;
      27704: inst = 32'h8220000;
      27705: inst = 32'h10408000;
      27706: inst = 32'hc405196;
      27707: inst = 32'h8220000;
      27708: inst = 32'h10408000;
      27709: inst = 32'hc405197;
      27710: inst = 32'h8220000;
      27711: inst = 32'h10408000;
      27712: inst = 32'hc405198;
      27713: inst = 32'h8220000;
      27714: inst = 32'h10408000;
      27715: inst = 32'hc4051dd;
      27716: inst = 32'h8220000;
      27717: inst = 32'h10408000;
      27718: inst = 32'hc4051de;
      27719: inst = 32'h8220000;
      27720: inst = 32'h10408000;
      27721: inst = 32'hc4051df;
      27722: inst = 32'h8220000;
      27723: inst = 32'h10408000;
      27724: inst = 32'hc4051e0;
      27725: inst = 32'h8220000;
      27726: inst = 32'h10408000;
      27727: inst = 32'hc4051e1;
      27728: inst = 32'h8220000;
      27729: inst = 32'h10408000;
      27730: inst = 32'hc4051e2;
      27731: inst = 32'h8220000;
      27732: inst = 32'h10408000;
      27733: inst = 32'hc4051f6;
      27734: inst = 32'h8220000;
      27735: inst = 32'h10408000;
      27736: inst = 32'hc4051f7;
      27737: inst = 32'h8220000;
      27738: inst = 32'h10408000;
      27739: inst = 32'hc4051f8;
      27740: inst = 32'h8220000;
      27741: inst = 32'h10408000;
      27742: inst = 32'hc40523d;
      27743: inst = 32'h8220000;
      27744: inst = 32'h10408000;
      27745: inst = 32'hc40523e;
      27746: inst = 32'h8220000;
      27747: inst = 32'h10408000;
      27748: inst = 32'hc40523f;
      27749: inst = 32'h8220000;
      27750: inst = 32'h10408000;
      27751: inst = 32'hc405240;
      27752: inst = 32'h8220000;
      27753: inst = 32'h10408000;
      27754: inst = 32'hc405241;
      27755: inst = 32'h8220000;
      27756: inst = 32'h10408000;
      27757: inst = 32'hc405242;
      27758: inst = 32'h8220000;
      27759: inst = 32'h10408000;
      27760: inst = 32'hc405256;
      27761: inst = 32'h8220000;
      27762: inst = 32'h10408000;
      27763: inst = 32'hc405257;
      27764: inst = 32'h8220000;
      27765: inst = 32'h10408000;
      27766: inst = 32'hc405258;
      27767: inst = 32'h8220000;
      27768: inst = 32'h10408000;
      27769: inst = 32'hc40529d;
      27770: inst = 32'h8220000;
      27771: inst = 32'h10408000;
      27772: inst = 32'hc40529e;
      27773: inst = 32'h8220000;
      27774: inst = 32'h10408000;
      27775: inst = 32'hc40529f;
      27776: inst = 32'h8220000;
      27777: inst = 32'h10408000;
      27778: inst = 32'hc4052a0;
      27779: inst = 32'h8220000;
      27780: inst = 32'h10408000;
      27781: inst = 32'hc4052a1;
      27782: inst = 32'h8220000;
      27783: inst = 32'h10408000;
      27784: inst = 32'hc4052a2;
      27785: inst = 32'h8220000;
      27786: inst = 32'h10408000;
      27787: inst = 32'hc4052b6;
      27788: inst = 32'h8220000;
      27789: inst = 32'h10408000;
      27790: inst = 32'hc4052b7;
      27791: inst = 32'h8220000;
      27792: inst = 32'h10408000;
      27793: inst = 32'hc4052b8;
      27794: inst = 32'h8220000;
      27795: inst = 32'h10408000;
      27796: inst = 32'hc4052fd;
      27797: inst = 32'h8220000;
      27798: inst = 32'h10408000;
      27799: inst = 32'hc4052fe;
      27800: inst = 32'h8220000;
      27801: inst = 32'h10408000;
      27802: inst = 32'hc4052ff;
      27803: inst = 32'h8220000;
      27804: inst = 32'h10408000;
      27805: inst = 32'hc405300;
      27806: inst = 32'h8220000;
      27807: inst = 32'h10408000;
      27808: inst = 32'hc405301;
      27809: inst = 32'h8220000;
      27810: inst = 32'h10408000;
      27811: inst = 32'hc405302;
      27812: inst = 32'h8220000;
      27813: inst = 32'h10408000;
      27814: inst = 32'hc405316;
      27815: inst = 32'h8220000;
      27816: inst = 32'h10408000;
      27817: inst = 32'hc405317;
      27818: inst = 32'h8220000;
      27819: inst = 32'h10408000;
      27820: inst = 32'hc405318;
      27821: inst = 32'h8220000;
      27822: inst = 32'h10408000;
      27823: inst = 32'hc40535d;
      27824: inst = 32'h8220000;
      27825: inst = 32'h10408000;
      27826: inst = 32'hc40535e;
      27827: inst = 32'h8220000;
      27828: inst = 32'h10408000;
      27829: inst = 32'hc40535f;
      27830: inst = 32'h8220000;
      27831: inst = 32'h10408000;
      27832: inst = 32'hc405360;
      27833: inst = 32'h8220000;
      27834: inst = 32'h10408000;
      27835: inst = 32'hc405361;
      27836: inst = 32'h8220000;
      27837: inst = 32'h10408000;
      27838: inst = 32'hc405362;
      27839: inst = 32'h8220000;
      27840: inst = 32'h10408000;
      27841: inst = 32'hc405376;
      27842: inst = 32'h8220000;
      27843: inst = 32'h10408000;
      27844: inst = 32'hc405377;
      27845: inst = 32'h8220000;
      27846: inst = 32'h10408000;
      27847: inst = 32'hc405378;
      27848: inst = 32'h8220000;
      27849: inst = 32'h10408000;
      27850: inst = 32'hc4053bd;
      27851: inst = 32'h8220000;
      27852: inst = 32'h10408000;
      27853: inst = 32'hc4053be;
      27854: inst = 32'h8220000;
      27855: inst = 32'h10408000;
      27856: inst = 32'hc4053bf;
      27857: inst = 32'h8220000;
      27858: inst = 32'h10408000;
      27859: inst = 32'hc4053c0;
      27860: inst = 32'h8220000;
      27861: inst = 32'h10408000;
      27862: inst = 32'hc4053c1;
      27863: inst = 32'h8220000;
      27864: inst = 32'h10408000;
      27865: inst = 32'hc4053c2;
      27866: inst = 32'h8220000;
      27867: inst = 32'h10408000;
      27868: inst = 32'hc4053d6;
      27869: inst = 32'h8220000;
      27870: inst = 32'h10408000;
      27871: inst = 32'hc4053d7;
      27872: inst = 32'h8220000;
      27873: inst = 32'h10408000;
      27874: inst = 32'hc4053d8;
      27875: inst = 32'h8220000;
      27876: inst = 32'h10408000;
      27877: inst = 32'hc40541d;
      27878: inst = 32'h8220000;
      27879: inst = 32'h10408000;
      27880: inst = 32'hc40541e;
      27881: inst = 32'h8220000;
      27882: inst = 32'h10408000;
      27883: inst = 32'hc40541f;
      27884: inst = 32'h8220000;
      27885: inst = 32'h10408000;
      27886: inst = 32'hc405420;
      27887: inst = 32'h8220000;
      27888: inst = 32'h10408000;
      27889: inst = 32'hc405421;
      27890: inst = 32'h8220000;
      27891: inst = 32'h10408000;
      27892: inst = 32'hc405422;
      27893: inst = 32'h8220000;
      27894: inst = 32'h10408000;
      27895: inst = 32'hc405436;
      27896: inst = 32'h8220000;
      27897: inst = 32'h10408000;
      27898: inst = 32'hc405437;
      27899: inst = 32'h8220000;
      27900: inst = 32'h10408000;
      27901: inst = 32'hc405438;
      27902: inst = 32'h8220000;
      27903: inst = 32'h10408000;
      27904: inst = 32'hc405439;
      27905: inst = 32'h8220000;
      27906: inst = 32'h10408000;
      27907: inst = 32'hc40543a;
      27908: inst = 32'h8220000;
      27909: inst = 32'h10408000;
      27910: inst = 32'hc40543b;
      27911: inst = 32'h8220000;
      27912: inst = 32'h10408000;
      27913: inst = 32'hc40543c;
      27914: inst = 32'h8220000;
      27915: inst = 32'h10408000;
      27916: inst = 32'hc40543d;
      27917: inst = 32'h8220000;
      27918: inst = 32'h10408000;
      27919: inst = 32'hc40543e;
      27920: inst = 32'h8220000;
      27921: inst = 32'h10408000;
      27922: inst = 32'hc40543f;
      27923: inst = 32'h8220000;
      27924: inst = 32'h10408000;
      27925: inst = 32'hc405440;
      27926: inst = 32'h8220000;
      27927: inst = 32'h10408000;
      27928: inst = 32'hc405441;
      27929: inst = 32'h8220000;
      27930: inst = 32'h10408000;
      27931: inst = 32'hc405442;
      27932: inst = 32'h8220000;
      27933: inst = 32'h10408000;
      27934: inst = 32'hc405443;
      27935: inst = 32'h8220000;
      27936: inst = 32'h10408000;
      27937: inst = 32'hc405444;
      27938: inst = 32'h8220000;
      27939: inst = 32'h10408000;
      27940: inst = 32'hc405445;
      27941: inst = 32'h8220000;
      27942: inst = 32'h10408000;
      27943: inst = 32'hc405446;
      27944: inst = 32'h8220000;
      27945: inst = 32'h10408000;
      27946: inst = 32'hc405447;
      27947: inst = 32'h8220000;
      27948: inst = 32'h10408000;
      27949: inst = 32'hc405448;
      27950: inst = 32'h8220000;
      27951: inst = 32'h10408000;
      27952: inst = 32'hc405449;
      27953: inst = 32'h8220000;
      27954: inst = 32'h10408000;
      27955: inst = 32'hc40547d;
      27956: inst = 32'h8220000;
      27957: inst = 32'h10408000;
      27958: inst = 32'hc40547e;
      27959: inst = 32'h8220000;
      27960: inst = 32'h10408000;
      27961: inst = 32'hc40547f;
      27962: inst = 32'h8220000;
      27963: inst = 32'h10408000;
      27964: inst = 32'hc405480;
      27965: inst = 32'h8220000;
      27966: inst = 32'h10408000;
      27967: inst = 32'hc405481;
      27968: inst = 32'h8220000;
      27969: inst = 32'h10408000;
      27970: inst = 32'hc405482;
      27971: inst = 32'h8220000;
      27972: inst = 32'h10408000;
      27973: inst = 32'hc405496;
      27974: inst = 32'h8220000;
      27975: inst = 32'h10408000;
      27976: inst = 32'hc405497;
      27977: inst = 32'h8220000;
      27978: inst = 32'h10408000;
      27979: inst = 32'hc405498;
      27980: inst = 32'h8220000;
      27981: inst = 32'h10408000;
      27982: inst = 32'hc405499;
      27983: inst = 32'h8220000;
      27984: inst = 32'h10408000;
      27985: inst = 32'hc40549a;
      27986: inst = 32'h8220000;
      27987: inst = 32'h10408000;
      27988: inst = 32'hc40549b;
      27989: inst = 32'h8220000;
      27990: inst = 32'h10408000;
      27991: inst = 32'hc40549c;
      27992: inst = 32'h8220000;
      27993: inst = 32'h10408000;
      27994: inst = 32'hc40549d;
      27995: inst = 32'h8220000;
      27996: inst = 32'h10408000;
      27997: inst = 32'hc40549e;
      27998: inst = 32'h8220000;
      27999: inst = 32'h10408000;
      28000: inst = 32'hc40549f;
      28001: inst = 32'h8220000;
      28002: inst = 32'h10408000;
      28003: inst = 32'hc4054a0;
      28004: inst = 32'h8220000;
      28005: inst = 32'h10408000;
      28006: inst = 32'hc4054a1;
      28007: inst = 32'h8220000;
      28008: inst = 32'h10408000;
      28009: inst = 32'hc4054a2;
      28010: inst = 32'h8220000;
      28011: inst = 32'h10408000;
      28012: inst = 32'hc4054a3;
      28013: inst = 32'h8220000;
      28014: inst = 32'h10408000;
      28015: inst = 32'hc4054a4;
      28016: inst = 32'h8220000;
      28017: inst = 32'h10408000;
      28018: inst = 32'hc4054a5;
      28019: inst = 32'h8220000;
      28020: inst = 32'h10408000;
      28021: inst = 32'hc4054a6;
      28022: inst = 32'h8220000;
      28023: inst = 32'h10408000;
      28024: inst = 32'hc4054a7;
      28025: inst = 32'h8220000;
      28026: inst = 32'h10408000;
      28027: inst = 32'hc4054a8;
      28028: inst = 32'h8220000;
      28029: inst = 32'h10408000;
      28030: inst = 32'hc4054a9;
      28031: inst = 32'h8220000;
      28032: inst = 32'h10408000;
      28033: inst = 32'hc4054dd;
      28034: inst = 32'h8220000;
      28035: inst = 32'h10408000;
      28036: inst = 32'hc4054de;
      28037: inst = 32'h8220000;
      28038: inst = 32'h10408000;
      28039: inst = 32'hc4054df;
      28040: inst = 32'h8220000;
      28041: inst = 32'h10408000;
      28042: inst = 32'hc4054e0;
      28043: inst = 32'h8220000;
      28044: inst = 32'h10408000;
      28045: inst = 32'hc4054e1;
      28046: inst = 32'h8220000;
      28047: inst = 32'h10408000;
      28048: inst = 32'hc4054e2;
      28049: inst = 32'h8220000;
      28050: inst = 32'h10408000;
      28051: inst = 32'hc4054f6;
      28052: inst = 32'h8220000;
      28053: inst = 32'h10408000;
      28054: inst = 32'hc4054f7;
      28055: inst = 32'h8220000;
      28056: inst = 32'h10408000;
      28057: inst = 32'hc4054f8;
      28058: inst = 32'h8220000;
      28059: inst = 32'h10408000;
      28060: inst = 32'hc4054f9;
      28061: inst = 32'h8220000;
      28062: inst = 32'h10408000;
      28063: inst = 32'hc4054fa;
      28064: inst = 32'h8220000;
      28065: inst = 32'h10408000;
      28066: inst = 32'hc4054fb;
      28067: inst = 32'h8220000;
      28068: inst = 32'h10408000;
      28069: inst = 32'hc4054fc;
      28070: inst = 32'h8220000;
      28071: inst = 32'h10408000;
      28072: inst = 32'hc4054fd;
      28073: inst = 32'h8220000;
      28074: inst = 32'h10408000;
      28075: inst = 32'hc4054fe;
      28076: inst = 32'h8220000;
      28077: inst = 32'h10408000;
      28078: inst = 32'hc4054ff;
      28079: inst = 32'h8220000;
      28080: inst = 32'h10408000;
      28081: inst = 32'hc405500;
      28082: inst = 32'h8220000;
      28083: inst = 32'h10408000;
      28084: inst = 32'hc405501;
      28085: inst = 32'h8220000;
      28086: inst = 32'h10408000;
      28087: inst = 32'hc405502;
      28088: inst = 32'h8220000;
      28089: inst = 32'h10408000;
      28090: inst = 32'hc405503;
      28091: inst = 32'h8220000;
      28092: inst = 32'h10408000;
      28093: inst = 32'hc405504;
      28094: inst = 32'h8220000;
      28095: inst = 32'h10408000;
      28096: inst = 32'hc405505;
      28097: inst = 32'h8220000;
      28098: inst = 32'h10408000;
      28099: inst = 32'hc405506;
      28100: inst = 32'h8220000;
      28101: inst = 32'h10408000;
      28102: inst = 32'hc405507;
      28103: inst = 32'h8220000;
      28104: inst = 32'h10408000;
      28105: inst = 32'hc405508;
      28106: inst = 32'h8220000;
      28107: inst = 32'h10408000;
      28108: inst = 32'hc405509;
      28109: inst = 32'h8220000;
      28110: inst = 32'h10408000;
      28111: inst = 32'hc40553d;
      28112: inst = 32'h8220000;
      28113: inst = 32'h10408000;
      28114: inst = 32'hc40553e;
      28115: inst = 32'h8220000;
      28116: inst = 32'h10408000;
      28117: inst = 32'hc40553f;
      28118: inst = 32'h8220000;
      28119: inst = 32'h10408000;
      28120: inst = 32'hc405540;
      28121: inst = 32'h8220000;
      28122: inst = 32'h10408000;
      28123: inst = 32'hc405541;
      28124: inst = 32'h8220000;
      28125: inst = 32'h10408000;
      28126: inst = 32'hc405542;
      28127: inst = 32'h8220000;
      28128: inst = 32'h10408000;
      28129: inst = 32'hc405556;
      28130: inst = 32'h8220000;
      28131: inst = 32'h10408000;
      28132: inst = 32'hc405557;
      28133: inst = 32'h8220000;
      28134: inst = 32'h10408000;
      28135: inst = 32'hc405558;
      28136: inst = 32'h8220000;
      28137: inst = 32'h10408000;
      28138: inst = 32'hc40559d;
      28139: inst = 32'h8220000;
      28140: inst = 32'h10408000;
      28141: inst = 32'hc40559e;
      28142: inst = 32'h8220000;
      28143: inst = 32'h10408000;
      28144: inst = 32'hc40559f;
      28145: inst = 32'h8220000;
      28146: inst = 32'h10408000;
      28147: inst = 32'hc4055a0;
      28148: inst = 32'h8220000;
      28149: inst = 32'h10408000;
      28150: inst = 32'hc4055a1;
      28151: inst = 32'h8220000;
      28152: inst = 32'h10408000;
      28153: inst = 32'hc4055a2;
      28154: inst = 32'h8220000;
      28155: inst = 32'h10408000;
      28156: inst = 32'hc4055b6;
      28157: inst = 32'h8220000;
      28158: inst = 32'h10408000;
      28159: inst = 32'hc4055b7;
      28160: inst = 32'h8220000;
      28161: inst = 32'h10408000;
      28162: inst = 32'hc4055b8;
      28163: inst = 32'h8220000;
      28164: inst = 32'h10408000;
      28165: inst = 32'hc4055fd;
      28166: inst = 32'h8220000;
      28167: inst = 32'h10408000;
      28168: inst = 32'hc4055fe;
      28169: inst = 32'h8220000;
      28170: inst = 32'h10408000;
      28171: inst = 32'hc4055ff;
      28172: inst = 32'h8220000;
      28173: inst = 32'h10408000;
      28174: inst = 32'hc405600;
      28175: inst = 32'h8220000;
      28176: inst = 32'h10408000;
      28177: inst = 32'hc405601;
      28178: inst = 32'h8220000;
      28179: inst = 32'h10408000;
      28180: inst = 32'hc405602;
      28181: inst = 32'h8220000;
      28182: inst = 32'h10408000;
      28183: inst = 32'hc405616;
      28184: inst = 32'h8220000;
      28185: inst = 32'h10408000;
      28186: inst = 32'hc405617;
      28187: inst = 32'h8220000;
      28188: inst = 32'h10408000;
      28189: inst = 32'hc405618;
      28190: inst = 32'h8220000;
      28191: inst = 32'h10408000;
      28192: inst = 32'hc40565d;
      28193: inst = 32'h8220000;
      28194: inst = 32'h10408000;
      28195: inst = 32'hc40565e;
      28196: inst = 32'h8220000;
      28197: inst = 32'h10408000;
      28198: inst = 32'hc40565f;
      28199: inst = 32'h8220000;
      28200: inst = 32'h10408000;
      28201: inst = 32'hc405660;
      28202: inst = 32'h8220000;
      28203: inst = 32'h10408000;
      28204: inst = 32'hc405661;
      28205: inst = 32'h8220000;
      28206: inst = 32'h10408000;
      28207: inst = 32'hc405662;
      28208: inst = 32'h8220000;
      28209: inst = 32'h10408000;
      28210: inst = 32'hc405676;
      28211: inst = 32'h8220000;
      28212: inst = 32'h10408000;
      28213: inst = 32'hc405677;
      28214: inst = 32'h8220000;
      28215: inst = 32'h10408000;
      28216: inst = 32'hc405678;
      28217: inst = 32'h8220000;
      28218: inst = 32'h10408000;
      28219: inst = 32'hc4056b7;
      28220: inst = 32'h8220000;
      28221: inst = 32'h10408000;
      28222: inst = 32'hc4056b8;
      28223: inst = 32'h8220000;
      28224: inst = 32'h10408000;
      28225: inst = 32'hc4056b9;
      28226: inst = 32'h8220000;
      28227: inst = 32'h10408000;
      28228: inst = 32'hc4056bd;
      28229: inst = 32'h8220000;
      28230: inst = 32'h10408000;
      28231: inst = 32'hc4056be;
      28232: inst = 32'h8220000;
      28233: inst = 32'h10408000;
      28234: inst = 32'hc4056bf;
      28235: inst = 32'h8220000;
      28236: inst = 32'h10408000;
      28237: inst = 32'hc4056c0;
      28238: inst = 32'h8220000;
      28239: inst = 32'h10408000;
      28240: inst = 32'hc4056c1;
      28241: inst = 32'h8220000;
      28242: inst = 32'h10408000;
      28243: inst = 32'hc4056c2;
      28244: inst = 32'h8220000;
      28245: inst = 32'h10408000;
      28246: inst = 32'hc4056c3;
      28247: inst = 32'h8220000;
      28248: inst = 32'h10408000;
      28249: inst = 32'hc4056c4;
      28250: inst = 32'h8220000;
      28251: inst = 32'h10408000;
      28252: inst = 32'hc4056c5;
      28253: inst = 32'h8220000;
      28254: inst = 32'h10408000;
      28255: inst = 32'hc4056c6;
      28256: inst = 32'h8220000;
      28257: inst = 32'h10408000;
      28258: inst = 32'hc4056c7;
      28259: inst = 32'h8220000;
      28260: inst = 32'h10408000;
      28261: inst = 32'hc4056c8;
      28262: inst = 32'h8220000;
      28263: inst = 32'h10408000;
      28264: inst = 32'hc4056c9;
      28265: inst = 32'h8220000;
      28266: inst = 32'h10408000;
      28267: inst = 32'hc4056d4;
      28268: inst = 32'h8220000;
      28269: inst = 32'h10408000;
      28270: inst = 32'hc4056d5;
      28271: inst = 32'h8220000;
      28272: inst = 32'h10408000;
      28273: inst = 32'hc4056d6;
      28274: inst = 32'h8220000;
      28275: inst = 32'h10408000;
      28276: inst = 32'hc4056d7;
      28277: inst = 32'h8220000;
      28278: inst = 32'h10408000;
      28279: inst = 32'hc4056d8;
      28280: inst = 32'h8220000;
      28281: inst = 32'h10408000;
      28282: inst = 32'hc4056d9;
      28283: inst = 32'h8220000;
      28284: inst = 32'h10408000;
      28285: inst = 32'hc4056da;
      28286: inst = 32'h8220000;
      28287: inst = 32'h10408000;
      28288: inst = 32'hc4056db;
      28289: inst = 32'h8220000;
      28290: inst = 32'h10408000;
      28291: inst = 32'hc4056dc;
      28292: inst = 32'h8220000;
      28293: inst = 32'h10408000;
      28294: inst = 32'hc4056dd;
      28295: inst = 32'h8220000;
      28296: inst = 32'h10408000;
      28297: inst = 32'hc4056de;
      28298: inst = 32'h8220000;
      28299: inst = 32'h10408000;
      28300: inst = 32'hc4056df;
      28301: inst = 32'h8220000;
      28302: inst = 32'h10408000;
      28303: inst = 32'hc4056e0;
      28304: inst = 32'h8220000;
      28305: inst = 32'h10408000;
      28306: inst = 32'hc4056e1;
      28307: inst = 32'h8220000;
      28308: inst = 32'h10408000;
      28309: inst = 32'hc4056e2;
      28310: inst = 32'h8220000;
      28311: inst = 32'h10408000;
      28312: inst = 32'hc4056e3;
      28313: inst = 32'h8220000;
      28314: inst = 32'h10408000;
      28315: inst = 32'hc4056e4;
      28316: inst = 32'h8220000;
      28317: inst = 32'h10408000;
      28318: inst = 32'hc4056e5;
      28319: inst = 32'h8220000;
      28320: inst = 32'h10408000;
      28321: inst = 32'hc4056e6;
      28322: inst = 32'h8220000;
      28323: inst = 32'h10408000;
      28324: inst = 32'hc4056e7;
      28325: inst = 32'h8220000;
      28326: inst = 32'h10408000;
      28327: inst = 32'hc4056e8;
      28328: inst = 32'h8220000;
      28329: inst = 32'h10408000;
      28330: inst = 32'hc4056e9;
      28331: inst = 32'h8220000;
      28332: inst = 32'h10408000;
      28333: inst = 32'hc4056ea;
      28334: inst = 32'h8220000;
      28335: inst = 32'h10408000;
      28336: inst = 32'hc4056eb;
      28337: inst = 32'h8220000;
      28338: inst = 32'h10408000;
      28339: inst = 32'hc4056ec;
      28340: inst = 32'h8220000;
      28341: inst = 32'h10408000;
      28342: inst = 32'hc4056ed;
      28343: inst = 32'h8220000;
      28344: inst = 32'h10408000;
      28345: inst = 32'hc4056ee;
      28346: inst = 32'h8220000;
      28347: inst = 32'h10408000;
      28348: inst = 32'hc4056ef;
      28349: inst = 32'h8220000;
      28350: inst = 32'h10408000;
      28351: inst = 32'hc4056f0;
      28352: inst = 32'h8220000;
      28353: inst = 32'h10408000;
      28354: inst = 32'hc4056f1;
      28355: inst = 32'h8220000;
      28356: inst = 32'h10408000;
      28357: inst = 32'hc4056f2;
      28358: inst = 32'h8220000;
      28359: inst = 32'h10408000;
      28360: inst = 32'hc4056f3;
      28361: inst = 32'h8220000;
      28362: inst = 32'h10408000;
      28363: inst = 32'hc4056f4;
      28364: inst = 32'h8220000;
      28365: inst = 32'h10408000;
      28366: inst = 32'hc4056f5;
      28367: inst = 32'h8220000;
      28368: inst = 32'h10408000;
      28369: inst = 32'hc4056f6;
      28370: inst = 32'h8220000;
      28371: inst = 32'h10408000;
      28372: inst = 32'hc4056f7;
      28373: inst = 32'h8220000;
      28374: inst = 32'h10408000;
      28375: inst = 32'hc4056f8;
      28376: inst = 32'h8220000;
      28377: inst = 32'h10408000;
      28378: inst = 32'hc4056f9;
      28379: inst = 32'h8220000;
      28380: inst = 32'h10408000;
      28381: inst = 32'hc4056fa;
      28382: inst = 32'h8220000;
      28383: inst = 32'h10408000;
      28384: inst = 32'hc4056fb;
      28385: inst = 32'h8220000;
      28386: inst = 32'h10408000;
      28387: inst = 32'hc4056fc;
      28388: inst = 32'h8220000;
      28389: inst = 32'h10408000;
      28390: inst = 32'hc4056fd;
      28391: inst = 32'h8220000;
      28392: inst = 32'h10408000;
      28393: inst = 32'hc405701;
      28394: inst = 32'h8220000;
      28395: inst = 32'h10408000;
      28396: inst = 32'hc405702;
      28397: inst = 32'h8220000;
      28398: inst = 32'h10408000;
      28399: inst = 32'hc405703;
      28400: inst = 32'h8220000;
      28401: inst = 32'h10408000;
      28402: inst = 32'hc405704;
      28403: inst = 32'h8220000;
      28404: inst = 32'h10408000;
      28405: inst = 32'hc405705;
      28406: inst = 32'h8220000;
      28407: inst = 32'h10408000;
      28408: inst = 32'hc405706;
      28409: inst = 32'h8220000;
      28410: inst = 32'h10408000;
      28411: inst = 32'hc405707;
      28412: inst = 32'h8220000;
      28413: inst = 32'h10408000;
      28414: inst = 32'hc405708;
      28415: inst = 32'h8220000;
      28416: inst = 32'h10408000;
      28417: inst = 32'hc405709;
      28418: inst = 32'h8220000;
      28419: inst = 32'h10408000;
      28420: inst = 32'hc40570a;
      28421: inst = 32'h8220000;
      28422: inst = 32'h10408000;
      28423: inst = 32'hc40570b;
      28424: inst = 32'h8220000;
      28425: inst = 32'h10408000;
      28426: inst = 32'hc40570c;
      28427: inst = 32'h8220000;
      28428: inst = 32'h10408000;
      28429: inst = 32'hc40570d;
      28430: inst = 32'h8220000;
      28431: inst = 32'h10408000;
      28432: inst = 32'hc40570e;
      28433: inst = 32'h8220000;
      28434: inst = 32'h10408000;
      28435: inst = 32'hc40570f;
      28436: inst = 32'h8220000;
      28437: inst = 32'h10408000;
      28438: inst = 32'hc405710;
      28439: inst = 32'h8220000;
      28440: inst = 32'h10408000;
      28441: inst = 32'hc405717;
      28442: inst = 32'h8220000;
      28443: inst = 32'h10408000;
      28444: inst = 32'hc405718;
      28445: inst = 32'h8220000;
      28446: inst = 32'h10408000;
      28447: inst = 32'hc405719;
      28448: inst = 32'h8220000;
      28449: inst = 32'h10408000;
      28450: inst = 32'hc40571d;
      28451: inst = 32'h8220000;
      28452: inst = 32'h10408000;
      28453: inst = 32'hc40571e;
      28454: inst = 32'h8220000;
      28455: inst = 32'h10408000;
      28456: inst = 32'hc40571f;
      28457: inst = 32'h8220000;
      28458: inst = 32'h10408000;
      28459: inst = 32'hc405720;
      28460: inst = 32'h8220000;
      28461: inst = 32'h10408000;
      28462: inst = 32'hc405721;
      28463: inst = 32'h8220000;
      28464: inst = 32'h10408000;
      28465: inst = 32'hc405722;
      28466: inst = 32'h8220000;
      28467: inst = 32'h10408000;
      28468: inst = 32'hc405723;
      28469: inst = 32'h8220000;
      28470: inst = 32'h10408000;
      28471: inst = 32'hc405724;
      28472: inst = 32'h8220000;
      28473: inst = 32'h10408000;
      28474: inst = 32'hc405725;
      28475: inst = 32'h8220000;
      28476: inst = 32'h10408000;
      28477: inst = 32'hc405726;
      28478: inst = 32'h8220000;
      28479: inst = 32'h10408000;
      28480: inst = 32'hc405727;
      28481: inst = 32'h8220000;
      28482: inst = 32'h10408000;
      28483: inst = 32'hc405728;
      28484: inst = 32'h8220000;
      28485: inst = 32'h10408000;
      28486: inst = 32'hc405729;
      28487: inst = 32'h8220000;
      28488: inst = 32'h10408000;
      28489: inst = 32'hc40572a;
      28490: inst = 32'h8220000;
      28491: inst = 32'h10408000;
      28492: inst = 32'hc40572b;
      28493: inst = 32'h8220000;
      28494: inst = 32'h10408000;
      28495: inst = 32'hc40572c;
      28496: inst = 32'h8220000;
      28497: inst = 32'h10408000;
      28498: inst = 32'hc40572d;
      28499: inst = 32'h8220000;
      28500: inst = 32'h10408000;
      28501: inst = 32'hc40572e;
      28502: inst = 32'h8220000;
      28503: inst = 32'h10408000;
      28504: inst = 32'hc40572f;
      28505: inst = 32'h8220000;
      28506: inst = 32'h10408000;
      28507: inst = 32'hc405730;
      28508: inst = 32'h8220000;
      28509: inst = 32'h10408000;
      28510: inst = 32'hc405731;
      28511: inst = 32'h8220000;
      28512: inst = 32'h10408000;
      28513: inst = 32'hc405732;
      28514: inst = 32'h8220000;
      28515: inst = 32'h10408000;
      28516: inst = 32'hc405733;
      28517: inst = 32'h8220000;
      28518: inst = 32'h10408000;
      28519: inst = 32'hc405734;
      28520: inst = 32'h8220000;
      28521: inst = 32'h10408000;
      28522: inst = 32'hc405735;
      28523: inst = 32'h8220000;
      28524: inst = 32'h10408000;
      28525: inst = 32'hc405736;
      28526: inst = 32'h8220000;
      28527: inst = 32'h10408000;
      28528: inst = 32'hc405737;
      28529: inst = 32'h8220000;
      28530: inst = 32'h10408000;
      28531: inst = 32'hc405738;
      28532: inst = 32'h8220000;
      28533: inst = 32'h10408000;
      28534: inst = 32'hc405739;
      28535: inst = 32'h8220000;
      28536: inst = 32'h10408000;
      28537: inst = 32'hc40573a;
      28538: inst = 32'h8220000;
      28539: inst = 32'h10408000;
      28540: inst = 32'hc40573b;
      28541: inst = 32'h8220000;
      28542: inst = 32'h10408000;
      28543: inst = 32'hc40573c;
      28544: inst = 32'h8220000;
      28545: inst = 32'h10408000;
      28546: inst = 32'hc40573d;
      28547: inst = 32'h8220000;
      28548: inst = 32'h10408000;
      28549: inst = 32'hc40573e;
      28550: inst = 32'h8220000;
      28551: inst = 32'h10408000;
      28552: inst = 32'hc40573f;
      28553: inst = 32'h8220000;
      28554: inst = 32'h10408000;
      28555: inst = 32'hc405740;
      28556: inst = 32'h8220000;
      28557: inst = 32'h10408000;
      28558: inst = 32'hc405741;
      28559: inst = 32'h8220000;
      28560: inst = 32'h10408000;
      28561: inst = 32'hc405742;
      28562: inst = 32'h8220000;
      28563: inst = 32'h10408000;
      28564: inst = 32'hc405743;
      28565: inst = 32'h8220000;
      28566: inst = 32'h10408000;
      28567: inst = 32'hc405744;
      28568: inst = 32'h8220000;
      28569: inst = 32'h10408000;
      28570: inst = 32'hc405745;
      28571: inst = 32'h8220000;
      28572: inst = 32'h10408000;
      28573: inst = 32'hc405746;
      28574: inst = 32'h8220000;
      28575: inst = 32'h10408000;
      28576: inst = 32'hc405747;
      28577: inst = 32'h8220000;
      28578: inst = 32'h10408000;
      28579: inst = 32'hc405748;
      28580: inst = 32'h8220000;
      28581: inst = 32'h10408000;
      28582: inst = 32'hc405749;
      28583: inst = 32'h8220000;
      28584: inst = 32'h10408000;
      28585: inst = 32'hc40574a;
      28586: inst = 32'h8220000;
      28587: inst = 32'h10408000;
      28588: inst = 32'hc40574b;
      28589: inst = 32'h8220000;
      28590: inst = 32'h10408000;
      28591: inst = 32'hc40574c;
      28592: inst = 32'h8220000;
      28593: inst = 32'h10408000;
      28594: inst = 32'hc40574d;
      28595: inst = 32'h8220000;
      28596: inst = 32'h10408000;
      28597: inst = 32'hc40574e;
      28598: inst = 32'h8220000;
      28599: inst = 32'h10408000;
      28600: inst = 32'hc40574f;
      28601: inst = 32'h8220000;
      28602: inst = 32'h10408000;
      28603: inst = 32'hc405750;
      28604: inst = 32'h8220000;
      28605: inst = 32'h10408000;
      28606: inst = 32'hc405751;
      28607: inst = 32'h8220000;
      28608: inst = 32'h10408000;
      28609: inst = 32'hc405752;
      28610: inst = 32'h8220000;
      28611: inst = 32'h10408000;
      28612: inst = 32'hc405753;
      28613: inst = 32'h8220000;
      28614: inst = 32'h10408000;
      28615: inst = 32'hc405754;
      28616: inst = 32'h8220000;
      28617: inst = 32'h10408000;
      28618: inst = 32'hc405755;
      28619: inst = 32'h8220000;
      28620: inst = 32'h10408000;
      28621: inst = 32'hc405756;
      28622: inst = 32'h8220000;
      28623: inst = 32'h10408000;
      28624: inst = 32'hc405757;
      28625: inst = 32'h8220000;
      28626: inst = 32'h10408000;
      28627: inst = 32'hc405758;
      28628: inst = 32'h8220000;
      28629: inst = 32'h10408000;
      28630: inst = 32'hc405759;
      28631: inst = 32'h8220000;
      28632: inst = 32'h10408000;
      28633: inst = 32'hc40575a;
      28634: inst = 32'h8220000;
      28635: inst = 32'h10408000;
      28636: inst = 32'hc40575b;
      28637: inst = 32'h8220000;
      28638: inst = 32'h10408000;
      28639: inst = 32'hc40575c;
      28640: inst = 32'h8220000;
      28641: inst = 32'h10408000;
      28642: inst = 32'hc40575d;
      28643: inst = 32'h8220000;
      28644: inst = 32'h10408000;
      28645: inst = 32'hc40575e;
      28646: inst = 32'h8220000;
      28647: inst = 32'h10408000;
      28648: inst = 32'hc405761;
      28649: inst = 32'h8220000;
      28650: inst = 32'h10408000;
      28651: inst = 32'hc405762;
      28652: inst = 32'h8220000;
      28653: inst = 32'h10408000;
      28654: inst = 32'hc405763;
      28655: inst = 32'h8220000;
      28656: inst = 32'h10408000;
      28657: inst = 32'hc405764;
      28658: inst = 32'h8220000;
      28659: inst = 32'h10408000;
      28660: inst = 32'hc405765;
      28661: inst = 32'h8220000;
      28662: inst = 32'h10408000;
      28663: inst = 32'hc405766;
      28664: inst = 32'h8220000;
      28665: inst = 32'h10408000;
      28666: inst = 32'hc405767;
      28667: inst = 32'h8220000;
      28668: inst = 32'h10408000;
      28669: inst = 32'hc405768;
      28670: inst = 32'h8220000;
      28671: inst = 32'h10408000;
      28672: inst = 32'hc405769;
      28673: inst = 32'h8220000;
      28674: inst = 32'h10408000;
      28675: inst = 32'hc40576a;
      28676: inst = 32'h8220000;
      28677: inst = 32'h10408000;
      28678: inst = 32'hc40576b;
      28679: inst = 32'h8220000;
      28680: inst = 32'h10408000;
      28681: inst = 32'hc40576c;
      28682: inst = 32'h8220000;
      28683: inst = 32'h10408000;
      28684: inst = 32'hc40576d;
      28685: inst = 32'h8220000;
      28686: inst = 32'h10408000;
      28687: inst = 32'hc40576e;
      28688: inst = 32'h8220000;
      28689: inst = 32'h10408000;
      28690: inst = 32'hc40576f;
      28691: inst = 32'h8220000;
      28692: inst = 32'h10408000;
      28693: inst = 32'hc405770;
      28694: inst = 32'h8220000;
      28695: inst = 32'h10408000;
      28696: inst = 32'hc40577d;
      28697: inst = 32'h8220000;
      28698: inst = 32'h10408000;
      28699: inst = 32'hc40577e;
      28700: inst = 32'h8220000;
      28701: inst = 32'h10408000;
      28702: inst = 32'hc40577f;
      28703: inst = 32'h8220000;
      28704: inst = 32'h10408000;
      28705: inst = 32'hc405780;
      28706: inst = 32'h8220000;
      28707: inst = 32'h10408000;
      28708: inst = 32'hc405781;
      28709: inst = 32'h8220000;
      28710: inst = 32'h10408000;
      28711: inst = 32'hc405782;
      28712: inst = 32'h8220000;
      28713: inst = 32'h10408000;
      28714: inst = 32'hc405783;
      28715: inst = 32'h8220000;
      28716: inst = 32'h10408000;
      28717: inst = 32'hc405784;
      28718: inst = 32'h8220000;
      28719: inst = 32'h10408000;
      28720: inst = 32'hc405785;
      28721: inst = 32'h8220000;
      28722: inst = 32'h10408000;
      28723: inst = 32'hc405786;
      28724: inst = 32'h8220000;
      28725: inst = 32'h10408000;
      28726: inst = 32'hc405787;
      28727: inst = 32'h8220000;
      28728: inst = 32'h10408000;
      28729: inst = 32'hc405788;
      28730: inst = 32'h8220000;
      28731: inst = 32'h10408000;
      28732: inst = 32'hc405789;
      28733: inst = 32'h8220000;
      28734: inst = 32'h10408000;
      28735: inst = 32'hc40578a;
      28736: inst = 32'h8220000;
      28737: inst = 32'h10408000;
      28738: inst = 32'hc40578b;
      28739: inst = 32'h8220000;
      28740: inst = 32'h10408000;
      28741: inst = 32'hc40578c;
      28742: inst = 32'h8220000;
      28743: inst = 32'h10408000;
      28744: inst = 32'hc40578d;
      28745: inst = 32'h8220000;
      28746: inst = 32'h10408000;
      28747: inst = 32'hc40578e;
      28748: inst = 32'h8220000;
      28749: inst = 32'h10408000;
      28750: inst = 32'hc40578f;
      28751: inst = 32'h8220000;
      28752: inst = 32'h10408000;
      28753: inst = 32'hc405790;
      28754: inst = 32'h8220000;
      28755: inst = 32'h10408000;
      28756: inst = 32'hc405791;
      28757: inst = 32'h8220000;
      28758: inst = 32'h10408000;
      28759: inst = 32'hc405792;
      28760: inst = 32'h8220000;
      28761: inst = 32'h10408000;
      28762: inst = 32'hc405793;
      28763: inst = 32'h8220000;
      28764: inst = 32'h10408000;
      28765: inst = 32'hc405794;
      28766: inst = 32'h8220000;
      28767: inst = 32'h10408000;
      28768: inst = 32'hc405795;
      28769: inst = 32'h8220000;
      28770: inst = 32'h10408000;
      28771: inst = 32'hc405796;
      28772: inst = 32'h8220000;
      28773: inst = 32'h10408000;
      28774: inst = 32'hc405797;
      28775: inst = 32'h8220000;
      28776: inst = 32'h10408000;
      28777: inst = 32'hc405798;
      28778: inst = 32'h8220000;
      28779: inst = 32'h10408000;
      28780: inst = 32'hc405799;
      28781: inst = 32'h8220000;
      28782: inst = 32'h10408000;
      28783: inst = 32'hc40579a;
      28784: inst = 32'h8220000;
      28785: inst = 32'h10408000;
      28786: inst = 32'hc40579b;
      28787: inst = 32'h8220000;
      28788: inst = 32'h10408000;
      28789: inst = 32'hc40579c;
      28790: inst = 32'h8220000;
      28791: inst = 32'h10408000;
      28792: inst = 32'hc40579d;
      28793: inst = 32'h8220000;
      28794: inst = 32'h10408000;
      28795: inst = 32'hc40579e;
      28796: inst = 32'h8220000;
      28797: inst = 32'h10408000;
      28798: inst = 32'hc40579f;
      28799: inst = 32'h8220000;
      28800: inst = 32'h10408000;
      28801: inst = 32'hc4057a0;
      28802: inst = 32'h8220000;
      28803: inst = 32'h10408000;
      28804: inst = 32'hc4057a1;
      28805: inst = 32'h8220000;
      28806: inst = 32'h10408000;
      28807: inst = 32'hc4057a2;
      28808: inst = 32'h8220000;
      28809: inst = 32'h10408000;
      28810: inst = 32'hc4057a3;
      28811: inst = 32'h8220000;
      28812: inst = 32'h10408000;
      28813: inst = 32'hc4057a4;
      28814: inst = 32'h8220000;
      28815: inst = 32'h10408000;
      28816: inst = 32'hc4057a5;
      28817: inst = 32'h8220000;
      28818: inst = 32'h10408000;
      28819: inst = 32'hc4057a6;
      28820: inst = 32'h8220000;
      28821: inst = 32'h10408000;
      28822: inst = 32'hc4057a7;
      28823: inst = 32'h8220000;
      28824: inst = 32'h10408000;
      28825: inst = 32'hc4057a8;
      28826: inst = 32'h8220000;
      28827: inst = 32'h10408000;
      28828: inst = 32'hc4057a9;
      28829: inst = 32'h8220000;
      28830: inst = 32'h10408000;
      28831: inst = 32'hc4057aa;
      28832: inst = 32'h8220000;
      28833: inst = 32'h10408000;
      28834: inst = 32'hc4057ab;
      28835: inst = 32'h8220000;
      28836: inst = 32'h10408000;
      28837: inst = 32'hc4057ac;
      28838: inst = 32'h8220000;
      28839: inst = 32'h10408000;
      28840: inst = 32'hc4057ad;
      28841: inst = 32'h8220000;
      28842: inst = 32'h10408000;
      28843: inst = 32'hc4057ae;
      28844: inst = 32'h8220000;
      28845: inst = 32'h10408000;
      28846: inst = 32'hc4057af;
      28847: inst = 32'h8220000;
      28848: inst = 32'h10408000;
      28849: inst = 32'hc4057b0;
      28850: inst = 32'h8220000;
      28851: inst = 32'h10408000;
      28852: inst = 32'hc4057b1;
      28853: inst = 32'h8220000;
      28854: inst = 32'h10408000;
      28855: inst = 32'hc4057b2;
      28856: inst = 32'h8220000;
      28857: inst = 32'h10408000;
      28858: inst = 32'hc4057b3;
      28859: inst = 32'h8220000;
      28860: inst = 32'h10408000;
      28861: inst = 32'hc4057b4;
      28862: inst = 32'h8220000;
      28863: inst = 32'h10408000;
      28864: inst = 32'hc4057b5;
      28865: inst = 32'h8220000;
      28866: inst = 32'h10408000;
      28867: inst = 32'hc4057b6;
      28868: inst = 32'h8220000;
      28869: inst = 32'h10408000;
      28870: inst = 32'hc4057b7;
      28871: inst = 32'h8220000;
      28872: inst = 32'h10408000;
      28873: inst = 32'hc4057b8;
      28874: inst = 32'h8220000;
      28875: inst = 32'h10408000;
      28876: inst = 32'hc4057b9;
      28877: inst = 32'h8220000;
      28878: inst = 32'h10408000;
      28879: inst = 32'hc4057ba;
      28880: inst = 32'h8220000;
      28881: inst = 32'h10408000;
      28882: inst = 32'hc4057bb;
      28883: inst = 32'h8220000;
      28884: inst = 32'h10408000;
      28885: inst = 32'hc4057bc;
      28886: inst = 32'h8220000;
      28887: inst = 32'h10408000;
      28888: inst = 32'hc4057bd;
      28889: inst = 32'h8220000;
      28890: inst = 32'h10408000;
      28891: inst = 32'hc4057be;
      28892: inst = 32'h8220000;
      28893: inst = 32'h10408000;
      28894: inst = 32'hc4057c1;
      28895: inst = 32'h8220000;
      28896: inst = 32'h10408000;
      28897: inst = 32'hc4057c2;
      28898: inst = 32'h8220000;
      28899: inst = 32'h10408000;
      28900: inst = 32'hc4057c3;
      28901: inst = 32'h8220000;
      28902: inst = 32'h10408000;
      28903: inst = 32'hc4057c4;
      28904: inst = 32'h8220000;
      28905: inst = 32'h10408000;
      28906: inst = 32'hc4057c5;
      28907: inst = 32'h8220000;
      28908: inst = 32'h10408000;
      28909: inst = 32'hc4057c6;
      28910: inst = 32'h8220000;
      28911: inst = 32'h10408000;
      28912: inst = 32'hc4057c7;
      28913: inst = 32'h8220000;
      28914: inst = 32'h10408000;
      28915: inst = 32'hc4057c8;
      28916: inst = 32'h8220000;
      28917: inst = 32'h10408000;
      28918: inst = 32'hc4057c9;
      28919: inst = 32'h8220000;
      28920: inst = 32'h10408000;
      28921: inst = 32'hc4057ca;
      28922: inst = 32'h8220000;
      28923: inst = 32'h10408000;
      28924: inst = 32'hc4057cb;
      28925: inst = 32'h8220000;
      28926: inst = 32'h10408000;
      28927: inst = 32'hc4057cc;
      28928: inst = 32'h8220000;
      28929: inst = 32'h10408000;
      28930: inst = 32'hc4057cd;
      28931: inst = 32'h8220000;
      28932: inst = 32'h10408000;
      28933: inst = 32'hc4057ce;
      28934: inst = 32'h8220000;
      28935: inst = 32'h10408000;
      28936: inst = 32'hc4057cf;
      28937: inst = 32'h8220000;
      28938: inst = 32'h10408000;
      28939: inst = 32'hc4057d0;
      28940: inst = 32'h8220000;
      28941: inst = 32'h10408000;
      28942: inst = 32'hc4057dd;
      28943: inst = 32'h8220000;
      28944: inst = 32'h10408000;
      28945: inst = 32'hc4057de;
      28946: inst = 32'h8220000;
      28947: inst = 32'h10408000;
      28948: inst = 32'hc4057df;
      28949: inst = 32'h8220000;
      28950: inst = 32'hc20eeb6;
      28951: inst = 32'h10408000;
      28952: inst = 32'hc403fe3;
      28953: inst = 32'h8220000;
      28954: inst = 32'h10408000;
      28955: inst = 32'hc404043;
      28956: inst = 32'h8220000;
      28957: inst = 32'h10408000;
      28958: inst = 32'hc4040a3;
      28959: inst = 32'h8220000;
      28960: inst = 32'h10408000;
      28961: inst = 32'hc404103;
      28962: inst = 32'h8220000;
      28963: inst = 32'h10408000;
      28964: inst = 32'hc40410e;
      28965: inst = 32'h8220000;
      28966: inst = 32'h10408000;
      28967: inst = 32'hc40410f;
      28968: inst = 32'h8220000;
      28969: inst = 32'h10408000;
      28970: inst = 32'hc404110;
      28971: inst = 32'h8220000;
      28972: inst = 32'h10408000;
      28973: inst = 32'hc404111;
      28974: inst = 32'h8220000;
      28975: inst = 32'h10408000;
      28976: inst = 32'hc404112;
      28977: inst = 32'h8220000;
      28978: inst = 32'h10408000;
      28979: inst = 32'hc404115;
      28980: inst = 32'h8220000;
      28981: inst = 32'h10408000;
      28982: inst = 32'hc404118;
      28983: inst = 32'h8220000;
      28984: inst = 32'h10408000;
      28985: inst = 32'hc404119;
      28986: inst = 32'h8220000;
      28987: inst = 32'h10408000;
      28988: inst = 32'hc40411a;
      28989: inst = 32'h8220000;
      28990: inst = 32'h10408000;
      28991: inst = 32'hc40411b;
      28992: inst = 32'h8220000;
      28993: inst = 32'h10408000;
      28994: inst = 32'hc40411c;
      28995: inst = 32'h8220000;
      28996: inst = 32'h10408000;
      28997: inst = 32'hc40411d;
      28998: inst = 32'h8220000;
      28999: inst = 32'h10408000;
      29000: inst = 32'hc40411e;
      29001: inst = 32'h8220000;
      29002: inst = 32'h10408000;
      29003: inst = 32'hc40411f;
      29004: inst = 32'h8220000;
      29005: inst = 32'h10408000;
      29006: inst = 32'hc404120;
      29007: inst = 32'h8220000;
      29008: inst = 32'h10408000;
      29009: inst = 32'hc404121;
      29010: inst = 32'h8220000;
      29011: inst = 32'h10408000;
      29012: inst = 32'hc404122;
      29013: inst = 32'h8220000;
      29014: inst = 32'h10408000;
      29015: inst = 32'hc404123;
      29016: inst = 32'h8220000;
      29017: inst = 32'h10408000;
      29018: inst = 32'hc404124;
      29019: inst = 32'h8220000;
      29020: inst = 32'h10408000;
      29021: inst = 32'hc404125;
      29022: inst = 32'h8220000;
      29023: inst = 32'h10408000;
      29024: inst = 32'hc404126;
      29025: inst = 32'h8220000;
      29026: inst = 32'h10408000;
      29027: inst = 32'hc404127;
      29028: inst = 32'h8220000;
      29029: inst = 32'h10408000;
      29030: inst = 32'hc404128;
      29031: inst = 32'h8220000;
      29032: inst = 32'h10408000;
      29033: inst = 32'hc404129;
      29034: inst = 32'h8220000;
      29035: inst = 32'h10408000;
      29036: inst = 32'hc40412a;
      29037: inst = 32'h8220000;
      29038: inst = 32'h10408000;
      29039: inst = 32'hc40412b;
      29040: inst = 32'h8220000;
      29041: inst = 32'h10408000;
      29042: inst = 32'hc40412c;
      29043: inst = 32'h8220000;
      29044: inst = 32'h10408000;
      29045: inst = 32'hc40412d;
      29046: inst = 32'h8220000;
      29047: inst = 32'h10408000;
      29048: inst = 32'hc40412e;
      29049: inst = 32'h8220000;
      29050: inst = 32'h10408000;
      29051: inst = 32'hc40412f;
      29052: inst = 32'h8220000;
      29053: inst = 32'h10408000;
      29054: inst = 32'hc404130;
      29055: inst = 32'h8220000;
      29056: inst = 32'h10408000;
      29057: inst = 32'hc404131;
      29058: inst = 32'h8220000;
      29059: inst = 32'h10408000;
      29060: inst = 32'hc404132;
      29061: inst = 32'h8220000;
      29062: inst = 32'h10408000;
      29063: inst = 32'hc404133;
      29064: inst = 32'h8220000;
      29065: inst = 32'h10408000;
      29066: inst = 32'hc404134;
      29067: inst = 32'h8220000;
      29068: inst = 32'h10408000;
      29069: inst = 32'hc404135;
      29070: inst = 32'h8220000;
      29071: inst = 32'h10408000;
      29072: inst = 32'hc404136;
      29073: inst = 32'h8220000;
      29074: inst = 32'h10408000;
      29075: inst = 32'hc404137;
      29076: inst = 32'h8220000;
      29077: inst = 32'h10408000;
      29078: inst = 32'hc404138;
      29079: inst = 32'h8220000;
      29080: inst = 32'h10408000;
      29081: inst = 32'hc404139;
      29082: inst = 32'h8220000;
      29083: inst = 32'h10408000;
      29084: inst = 32'hc40413a;
      29085: inst = 32'h8220000;
      29086: inst = 32'h10408000;
      29087: inst = 32'hc40413b;
      29088: inst = 32'h8220000;
      29089: inst = 32'h10408000;
      29090: inst = 32'hc40413c;
      29091: inst = 32'h8220000;
      29092: inst = 32'h10408000;
      29093: inst = 32'hc40413d;
      29094: inst = 32'h8220000;
      29095: inst = 32'h10408000;
      29096: inst = 32'hc40413e;
      29097: inst = 32'h8220000;
      29098: inst = 32'h10408000;
      29099: inst = 32'hc40413f;
      29100: inst = 32'h8220000;
      29101: inst = 32'h10408000;
      29102: inst = 32'hc404140;
      29103: inst = 32'h8220000;
      29104: inst = 32'h10408000;
      29105: inst = 32'hc404141;
      29106: inst = 32'h8220000;
      29107: inst = 32'h10408000;
      29108: inst = 32'hc404142;
      29109: inst = 32'h8220000;
      29110: inst = 32'h10408000;
      29111: inst = 32'hc404143;
      29112: inst = 32'h8220000;
      29113: inst = 32'h10408000;
      29114: inst = 32'hc404144;
      29115: inst = 32'h8220000;
      29116: inst = 32'h10408000;
      29117: inst = 32'hc404145;
      29118: inst = 32'h8220000;
      29119: inst = 32'h10408000;
      29120: inst = 32'hc404146;
      29121: inst = 32'h8220000;
      29122: inst = 32'h10408000;
      29123: inst = 32'hc404147;
      29124: inst = 32'h8220000;
      29125: inst = 32'h10408000;
      29126: inst = 32'hc404148;
      29127: inst = 32'h8220000;
      29128: inst = 32'h10408000;
      29129: inst = 32'hc404149;
      29130: inst = 32'h8220000;
      29131: inst = 32'h10408000;
      29132: inst = 32'hc40414a;
      29133: inst = 32'h8220000;
      29134: inst = 32'h10408000;
      29135: inst = 32'hc40414b;
      29136: inst = 32'h8220000;
      29137: inst = 32'h10408000;
      29138: inst = 32'hc40414f;
      29139: inst = 32'h8220000;
      29140: inst = 32'h10408000;
      29141: inst = 32'hc404150;
      29142: inst = 32'h8220000;
      29143: inst = 32'h10408000;
      29144: inst = 32'hc404163;
      29145: inst = 32'h8220000;
      29146: inst = 32'h10408000;
      29147: inst = 32'hc40416e;
      29148: inst = 32'h8220000;
      29149: inst = 32'h10408000;
      29150: inst = 32'hc40416f;
      29151: inst = 32'h8220000;
      29152: inst = 32'h10408000;
      29153: inst = 32'hc404170;
      29154: inst = 32'h8220000;
      29155: inst = 32'h10408000;
      29156: inst = 32'hc404171;
      29157: inst = 32'h8220000;
      29158: inst = 32'h10408000;
      29159: inst = 32'hc404172;
      29160: inst = 32'h8220000;
      29161: inst = 32'h10408000;
      29162: inst = 32'hc404173;
      29163: inst = 32'h8220000;
      29164: inst = 32'h10408000;
      29165: inst = 32'hc404174;
      29166: inst = 32'h8220000;
      29167: inst = 32'h10408000;
      29168: inst = 32'hc404175;
      29169: inst = 32'h8220000;
      29170: inst = 32'h10408000;
      29171: inst = 32'hc404178;
      29172: inst = 32'h8220000;
      29173: inst = 32'h10408000;
      29174: inst = 32'hc404179;
      29175: inst = 32'h8220000;
      29176: inst = 32'h10408000;
      29177: inst = 32'hc40417a;
      29178: inst = 32'h8220000;
      29179: inst = 32'h10408000;
      29180: inst = 32'hc40417c;
      29181: inst = 32'h8220000;
      29182: inst = 32'h10408000;
      29183: inst = 32'hc40417d;
      29184: inst = 32'h8220000;
      29185: inst = 32'h10408000;
      29186: inst = 32'hc40417e;
      29187: inst = 32'h8220000;
      29188: inst = 32'h10408000;
      29189: inst = 32'hc40417f;
      29190: inst = 32'h8220000;
      29191: inst = 32'h10408000;
      29192: inst = 32'hc404180;
      29193: inst = 32'h8220000;
      29194: inst = 32'h10408000;
      29195: inst = 32'hc404181;
      29196: inst = 32'h8220000;
      29197: inst = 32'h10408000;
      29198: inst = 32'hc404182;
      29199: inst = 32'h8220000;
      29200: inst = 32'h10408000;
      29201: inst = 32'hc404183;
      29202: inst = 32'h8220000;
      29203: inst = 32'h10408000;
      29204: inst = 32'hc404184;
      29205: inst = 32'h8220000;
      29206: inst = 32'h10408000;
      29207: inst = 32'hc404185;
      29208: inst = 32'h8220000;
      29209: inst = 32'h10408000;
      29210: inst = 32'hc404186;
      29211: inst = 32'h8220000;
      29212: inst = 32'h10408000;
      29213: inst = 32'hc404187;
      29214: inst = 32'h8220000;
      29215: inst = 32'h10408000;
      29216: inst = 32'hc404188;
      29217: inst = 32'h8220000;
      29218: inst = 32'h10408000;
      29219: inst = 32'hc404189;
      29220: inst = 32'h8220000;
      29221: inst = 32'h10408000;
      29222: inst = 32'hc40418a;
      29223: inst = 32'h8220000;
      29224: inst = 32'h10408000;
      29225: inst = 32'hc40418b;
      29226: inst = 32'h8220000;
      29227: inst = 32'h10408000;
      29228: inst = 32'hc40418c;
      29229: inst = 32'h8220000;
      29230: inst = 32'h10408000;
      29231: inst = 32'hc40418d;
      29232: inst = 32'h8220000;
      29233: inst = 32'h10408000;
      29234: inst = 32'hc40418e;
      29235: inst = 32'h8220000;
      29236: inst = 32'h10408000;
      29237: inst = 32'hc40418f;
      29238: inst = 32'h8220000;
      29239: inst = 32'h10408000;
      29240: inst = 32'hc404190;
      29241: inst = 32'h8220000;
      29242: inst = 32'h10408000;
      29243: inst = 32'hc404191;
      29244: inst = 32'h8220000;
      29245: inst = 32'h10408000;
      29246: inst = 32'hc404192;
      29247: inst = 32'h8220000;
      29248: inst = 32'h10408000;
      29249: inst = 32'hc404193;
      29250: inst = 32'h8220000;
      29251: inst = 32'h10408000;
      29252: inst = 32'hc404194;
      29253: inst = 32'h8220000;
      29254: inst = 32'h10408000;
      29255: inst = 32'hc404195;
      29256: inst = 32'h8220000;
      29257: inst = 32'h10408000;
      29258: inst = 32'hc404196;
      29259: inst = 32'h8220000;
      29260: inst = 32'h10408000;
      29261: inst = 32'hc404197;
      29262: inst = 32'h8220000;
      29263: inst = 32'h10408000;
      29264: inst = 32'hc404198;
      29265: inst = 32'h8220000;
      29266: inst = 32'h10408000;
      29267: inst = 32'hc404199;
      29268: inst = 32'h8220000;
      29269: inst = 32'h10408000;
      29270: inst = 32'hc40419a;
      29271: inst = 32'h8220000;
      29272: inst = 32'h10408000;
      29273: inst = 32'hc40419b;
      29274: inst = 32'h8220000;
      29275: inst = 32'h10408000;
      29276: inst = 32'hc40419c;
      29277: inst = 32'h8220000;
      29278: inst = 32'h10408000;
      29279: inst = 32'hc40419d;
      29280: inst = 32'h8220000;
      29281: inst = 32'h10408000;
      29282: inst = 32'hc40419e;
      29283: inst = 32'h8220000;
      29284: inst = 32'h10408000;
      29285: inst = 32'hc40419f;
      29286: inst = 32'h8220000;
      29287: inst = 32'h10408000;
      29288: inst = 32'hc4041a0;
      29289: inst = 32'h8220000;
      29290: inst = 32'h10408000;
      29291: inst = 32'hc4041a1;
      29292: inst = 32'h8220000;
      29293: inst = 32'h10408000;
      29294: inst = 32'hc4041a2;
      29295: inst = 32'h8220000;
      29296: inst = 32'h10408000;
      29297: inst = 32'hc4041a3;
      29298: inst = 32'h8220000;
      29299: inst = 32'h10408000;
      29300: inst = 32'hc4041a4;
      29301: inst = 32'h8220000;
      29302: inst = 32'h10408000;
      29303: inst = 32'hc4041a5;
      29304: inst = 32'h8220000;
      29305: inst = 32'h10408000;
      29306: inst = 32'hc4041a6;
      29307: inst = 32'h8220000;
      29308: inst = 32'h10408000;
      29309: inst = 32'hc4041a7;
      29310: inst = 32'h8220000;
      29311: inst = 32'h10408000;
      29312: inst = 32'hc4041a8;
      29313: inst = 32'h8220000;
      29314: inst = 32'h10408000;
      29315: inst = 32'hc4041a9;
      29316: inst = 32'h8220000;
      29317: inst = 32'h10408000;
      29318: inst = 32'hc4041aa;
      29319: inst = 32'h8220000;
      29320: inst = 32'h10408000;
      29321: inst = 32'hc4041ab;
      29322: inst = 32'h8220000;
      29323: inst = 32'h10408000;
      29324: inst = 32'hc4041af;
      29325: inst = 32'h8220000;
      29326: inst = 32'h10408000;
      29327: inst = 32'hc4041b5;
      29328: inst = 32'h8220000;
      29329: inst = 32'h10408000;
      29330: inst = 32'hc4041c3;
      29331: inst = 32'h8220000;
      29332: inst = 32'h10408000;
      29333: inst = 32'hc4041cd;
      29334: inst = 32'h8220000;
      29335: inst = 32'h10408000;
      29336: inst = 32'hc4041ce;
      29337: inst = 32'h8220000;
      29338: inst = 32'h10408000;
      29339: inst = 32'hc4041cf;
      29340: inst = 32'h8220000;
      29341: inst = 32'h10408000;
      29342: inst = 32'hc4041d2;
      29343: inst = 32'h8220000;
      29344: inst = 32'h10408000;
      29345: inst = 32'hc4041d3;
      29346: inst = 32'h8220000;
      29347: inst = 32'h10408000;
      29348: inst = 32'hc4041d4;
      29349: inst = 32'h8220000;
      29350: inst = 32'h10408000;
      29351: inst = 32'hc4041d5;
      29352: inst = 32'h8220000;
      29353: inst = 32'h10408000;
      29354: inst = 32'hc4041d9;
      29355: inst = 32'h8220000;
      29356: inst = 32'h10408000;
      29357: inst = 32'hc4041da;
      29358: inst = 32'h8220000;
      29359: inst = 32'h10408000;
      29360: inst = 32'hc4041dd;
      29361: inst = 32'h8220000;
      29362: inst = 32'h10408000;
      29363: inst = 32'hc4041de;
      29364: inst = 32'h8220000;
      29365: inst = 32'h10408000;
      29366: inst = 32'hc4041df;
      29367: inst = 32'h8220000;
      29368: inst = 32'h10408000;
      29369: inst = 32'hc4041e0;
      29370: inst = 32'h8220000;
      29371: inst = 32'h10408000;
      29372: inst = 32'hc4041e1;
      29373: inst = 32'h8220000;
      29374: inst = 32'h10408000;
      29375: inst = 32'hc4041e2;
      29376: inst = 32'h8220000;
      29377: inst = 32'h10408000;
      29378: inst = 32'hc4041e3;
      29379: inst = 32'h8220000;
      29380: inst = 32'h10408000;
      29381: inst = 32'hc4041e4;
      29382: inst = 32'h8220000;
      29383: inst = 32'h10408000;
      29384: inst = 32'hc4041e5;
      29385: inst = 32'h8220000;
      29386: inst = 32'h10408000;
      29387: inst = 32'hc4041e6;
      29388: inst = 32'h8220000;
      29389: inst = 32'h10408000;
      29390: inst = 32'hc4041e7;
      29391: inst = 32'h8220000;
      29392: inst = 32'h10408000;
      29393: inst = 32'hc4041e8;
      29394: inst = 32'h8220000;
      29395: inst = 32'h10408000;
      29396: inst = 32'hc4041e9;
      29397: inst = 32'h8220000;
      29398: inst = 32'h10408000;
      29399: inst = 32'hc4041ea;
      29400: inst = 32'h8220000;
      29401: inst = 32'h10408000;
      29402: inst = 32'hc4041eb;
      29403: inst = 32'h8220000;
      29404: inst = 32'h10408000;
      29405: inst = 32'hc4041ec;
      29406: inst = 32'h8220000;
      29407: inst = 32'h10408000;
      29408: inst = 32'hc4041ed;
      29409: inst = 32'h8220000;
      29410: inst = 32'h10408000;
      29411: inst = 32'hc4041ee;
      29412: inst = 32'h8220000;
      29413: inst = 32'h10408000;
      29414: inst = 32'hc4041ef;
      29415: inst = 32'h8220000;
      29416: inst = 32'h10408000;
      29417: inst = 32'hc4041f0;
      29418: inst = 32'h8220000;
      29419: inst = 32'h10408000;
      29420: inst = 32'hc4041f1;
      29421: inst = 32'h8220000;
      29422: inst = 32'h10408000;
      29423: inst = 32'hc4041f2;
      29424: inst = 32'h8220000;
      29425: inst = 32'h10408000;
      29426: inst = 32'hc4041f3;
      29427: inst = 32'h8220000;
      29428: inst = 32'h10408000;
      29429: inst = 32'hc4041f4;
      29430: inst = 32'h8220000;
      29431: inst = 32'h10408000;
      29432: inst = 32'hc4041f5;
      29433: inst = 32'h8220000;
      29434: inst = 32'h10408000;
      29435: inst = 32'hc4041f6;
      29436: inst = 32'h8220000;
      29437: inst = 32'h10408000;
      29438: inst = 32'hc4041f7;
      29439: inst = 32'h8220000;
      29440: inst = 32'h10408000;
      29441: inst = 32'hc4041f8;
      29442: inst = 32'h8220000;
      29443: inst = 32'h10408000;
      29444: inst = 32'hc4041f9;
      29445: inst = 32'h8220000;
      29446: inst = 32'h10408000;
      29447: inst = 32'hc4041fa;
      29448: inst = 32'h8220000;
      29449: inst = 32'h10408000;
      29450: inst = 32'hc4041fb;
      29451: inst = 32'h8220000;
      29452: inst = 32'h10408000;
      29453: inst = 32'hc4041fc;
      29454: inst = 32'h8220000;
      29455: inst = 32'h10408000;
      29456: inst = 32'hc4041fd;
      29457: inst = 32'h8220000;
      29458: inst = 32'h10408000;
      29459: inst = 32'hc4041fe;
      29460: inst = 32'h8220000;
      29461: inst = 32'h10408000;
      29462: inst = 32'hc4041ff;
      29463: inst = 32'h8220000;
      29464: inst = 32'h10408000;
      29465: inst = 32'hc404200;
      29466: inst = 32'h8220000;
      29467: inst = 32'h10408000;
      29468: inst = 32'hc404201;
      29469: inst = 32'h8220000;
      29470: inst = 32'h10408000;
      29471: inst = 32'hc404202;
      29472: inst = 32'h8220000;
      29473: inst = 32'h10408000;
      29474: inst = 32'hc404203;
      29475: inst = 32'h8220000;
      29476: inst = 32'h10408000;
      29477: inst = 32'hc404204;
      29478: inst = 32'h8220000;
      29479: inst = 32'h10408000;
      29480: inst = 32'hc404205;
      29481: inst = 32'h8220000;
      29482: inst = 32'h10408000;
      29483: inst = 32'hc404206;
      29484: inst = 32'h8220000;
      29485: inst = 32'h10408000;
      29486: inst = 32'hc404207;
      29487: inst = 32'h8220000;
      29488: inst = 32'h10408000;
      29489: inst = 32'hc404208;
      29490: inst = 32'h8220000;
      29491: inst = 32'h10408000;
      29492: inst = 32'hc404209;
      29493: inst = 32'h8220000;
      29494: inst = 32'h10408000;
      29495: inst = 32'hc40420a;
      29496: inst = 32'h8220000;
      29497: inst = 32'h10408000;
      29498: inst = 32'hc40420b;
      29499: inst = 32'h8220000;
      29500: inst = 32'h10408000;
      29501: inst = 32'hc40420f;
      29502: inst = 32'h8220000;
      29503: inst = 32'h10408000;
      29504: inst = 32'hc404214;
      29505: inst = 32'h8220000;
      29506: inst = 32'h10408000;
      29507: inst = 32'hc404223;
      29508: inst = 32'h8220000;
      29509: inst = 32'h10408000;
      29510: inst = 32'hc40422d;
      29511: inst = 32'h8220000;
      29512: inst = 32'h10408000;
      29513: inst = 32'hc40422e;
      29514: inst = 32'h8220000;
      29515: inst = 32'h10408000;
      29516: inst = 32'hc404232;
      29517: inst = 32'h8220000;
      29518: inst = 32'h10408000;
      29519: inst = 32'hc404233;
      29520: inst = 32'h8220000;
      29521: inst = 32'h10408000;
      29522: inst = 32'hc404234;
      29523: inst = 32'h8220000;
      29524: inst = 32'h10408000;
      29525: inst = 32'hc404235;
      29526: inst = 32'h8220000;
      29527: inst = 32'h10408000;
      29528: inst = 32'hc404236;
      29529: inst = 32'h8220000;
      29530: inst = 32'h10408000;
      29531: inst = 32'hc404237;
      29532: inst = 32'h8220000;
      29533: inst = 32'h10408000;
      29534: inst = 32'hc404238;
      29535: inst = 32'h8220000;
      29536: inst = 32'h10408000;
      29537: inst = 32'hc404239;
      29538: inst = 32'h8220000;
      29539: inst = 32'h10408000;
      29540: inst = 32'hc40423a;
      29541: inst = 32'h8220000;
      29542: inst = 32'h10408000;
      29543: inst = 32'hc40423d;
      29544: inst = 32'h8220000;
      29545: inst = 32'h10408000;
      29546: inst = 32'hc40423e;
      29547: inst = 32'h8220000;
      29548: inst = 32'h10408000;
      29549: inst = 32'hc40423f;
      29550: inst = 32'h8220000;
      29551: inst = 32'h10408000;
      29552: inst = 32'hc404240;
      29553: inst = 32'h8220000;
      29554: inst = 32'h10408000;
      29555: inst = 32'hc404241;
      29556: inst = 32'h8220000;
      29557: inst = 32'h10408000;
      29558: inst = 32'hc404242;
      29559: inst = 32'h8220000;
      29560: inst = 32'h10408000;
      29561: inst = 32'hc404243;
      29562: inst = 32'h8220000;
      29563: inst = 32'h10408000;
      29564: inst = 32'hc404244;
      29565: inst = 32'h8220000;
      29566: inst = 32'h10408000;
      29567: inst = 32'hc404245;
      29568: inst = 32'h8220000;
      29569: inst = 32'h10408000;
      29570: inst = 32'hc404246;
      29571: inst = 32'h8220000;
      29572: inst = 32'h10408000;
      29573: inst = 32'hc404247;
      29574: inst = 32'h8220000;
      29575: inst = 32'h10408000;
      29576: inst = 32'hc404248;
      29577: inst = 32'h8220000;
      29578: inst = 32'h10408000;
      29579: inst = 32'hc404249;
      29580: inst = 32'h8220000;
      29581: inst = 32'h10408000;
      29582: inst = 32'hc40424a;
      29583: inst = 32'h8220000;
      29584: inst = 32'h10408000;
      29585: inst = 32'hc40424b;
      29586: inst = 32'h8220000;
      29587: inst = 32'h10408000;
      29588: inst = 32'hc40424c;
      29589: inst = 32'h8220000;
      29590: inst = 32'h10408000;
      29591: inst = 32'hc40424d;
      29592: inst = 32'h8220000;
      29593: inst = 32'h10408000;
      29594: inst = 32'hc40424e;
      29595: inst = 32'h8220000;
      29596: inst = 32'h10408000;
      29597: inst = 32'hc40424f;
      29598: inst = 32'h8220000;
      29599: inst = 32'h10408000;
      29600: inst = 32'hc404250;
      29601: inst = 32'h8220000;
      29602: inst = 32'h10408000;
      29603: inst = 32'hc404251;
      29604: inst = 32'h8220000;
      29605: inst = 32'h10408000;
      29606: inst = 32'hc404252;
      29607: inst = 32'h8220000;
      29608: inst = 32'h10408000;
      29609: inst = 32'hc404253;
      29610: inst = 32'h8220000;
      29611: inst = 32'h10408000;
      29612: inst = 32'hc404254;
      29613: inst = 32'h8220000;
      29614: inst = 32'h10408000;
      29615: inst = 32'hc404255;
      29616: inst = 32'h8220000;
      29617: inst = 32'h10408000;
      29618: inst = 32'hc404256;
      29619: inst = 32'h8220000;
      29620: inst = 32'h10408000;
      29621: inst = 32'hc404257;
      29622: inst = 32'h8220000;
      29623: inst = 32'h10408000;
      29624: inst = 32'hc404258;
      29625: inst = 32'h8220000;
      29626: inst = 32'h10408000;
      29627: inst = 32'hc404259;
      29628: inst = 32'h8220000;
      29629: inst = 32'h10408000;
      29630: inst = 32'hc40425a;
      29631: inst = 32'h8220000;
      29632: inst = 32'h10408000;
      29633: inst = 32'hc40425b;
      29634: inst = 32'h8220000;
      29635: inst = 32'h10408000;
      29636: inst = 32'hc40425c;
      29637: inst = 32'h8220000;
      29638: inst = 32'h10408000;
      29639: inst = 32'hc40425d;
      29640: inst = 32'h8220000;
      29641: inst = 32'h10408000;
      29642: inst = 32'hc40425e;
      29643: inst = 32'h8220000;
      29644: inst = 32'h10408000;
      29645: inst = 32'hc40425f;
      29646: inst = 32'h8220000;
      29647: inst = 32'h10408000;
      29648: inst = 32'hc404260;
      29649: inst = 32'h8220000;
      29650: inst = 32'h10408000;
      29651: inst = 32'hc404261;
      29652: inst = 32'h8220000;
      29653: inst = 32'h10408000;
      29654: inst = 32'hc404262;
      29655: inst = 32'h8220000;
      29656: inst = 32'h10408000;
      29657: inst = 32'hc404263;
      29658: inst = 32'h8220000;
      29659: inst = 32'h10408000;
      29660: inst = 32'hc404264;
      29661: inst = 32'h8220000;
      29662: inst = 32'h10408000;
      29663: inst = 32'hc404265;
      29664: inst = 32'h8220000;
      29665: inst = 32'h10408000;
      29666: inst = 32'hc404266;
      29667: inst = 32'h8220000;
      29668: inst = 32'h10408000;
      29669: inst = 32'hc404267;
      29670: inst = 32'h8220000;
      29671: inst = 32'h10408000;
      29672: inst = 32'hc404268;
      29673: inst = 32'h8220000;
      29674: inst = 32'h10408000;
      29675: inst = 32'hc404269;
      29676: inst = 32'h8220000;
      29677: inst = 32'h10408000;
      29678: inst = 32'hc40426a;
      29679: inst = 32'h8220000;
      29680: inst = 32'h10408000;
      29681: inst = 32'hc40426b;
      29682: inst = 32'h8220000;
      29683: inst = 32'h10408000;
      29684: inst = 32'hc40426f;
      29685: inst = 32'h8220000;
      29686: inst = 32'h10408000;
      29687: inst = 32'hc404283;
      29688: inst = 32'h8220000;
      29689: inst = 32'h10408000;
      29690: inst = 32'hc40428d;
      29691: inst = 32'h8220000;
      29692: inst = 32'h10408000;
      29693: inst = 32'hc40428e;
      29694: inst = 32'h8220000;
      29695: inst = 32'h10408000;
      29696: inst = 32'hc404291;
      29697: inst = 32'h8220000;
      29698: inst = 32'h10408000;
      29699: inst = 32'hc404292;
      29700: inst = 32'h8220000;
      29701: inst = 32'h10408000;
      29702: inst = 32'hc404293;
      29703: inst = 32'h8220000;
      29704: inst = 32'h10408000;
      29705: inst = 32'hc404294;
      29706: inst = 32'h8220000;
      29707: inst = 32'h10408000;
      29708: inst = 32'hc404295;
      29709: inst = 32'h8220000;
      29710: inst = 32'h10408000;
      29711: inst = 32'hc404296;
      29712: inst = 32'h8220000;
      29713: inst = 32'h10408000;
      29714: inst = 32'hc404297;
      29715: inst = 32'h8220000;
      29716: inst = 32'h10408000;
      29717: inst = 32'hc404298;
      29718: inst = 32'h8220000;
      29719: inst = 32'h10408000;
      29720: inst = 32'hc404299;
      29721: inst = 32'h8220000;
      29722: inst = 32'h10408000;
      29723: inst = 32'hc40429a;
      29724: inst = 32'h8220000;
      29725: inst = 32'h10408000;
      29726: inst = 32'hc40429d;
      29727: inst = 32'h8220000;
      29728: inst = 32'h10408000;
      29729: inst = 32'hc40429e;
      29730: inst = 32'h8220000;
      29731: inst = 32'h10408000;
      29732: inst = 32'hc40429f;
      29733: inst = 32'h8220000;
      29734: inst = 32'h10408000;
      29735: inst = 32'hc4042a0;
      29736: inst = 32'h8220000;
      29737: inst = 32'h10408000;
      29738: inst = 32'hc4042a1;
      29739: inst = 32'h8220000;
      29740: inst = 32'h10408000;
      29741: inst = 32'hc4042a2;
      29742: inst = 32'h8220000;
      29743: inst = 32'h10408000;
      29744: inst = 32'hc4042a3;
      29745: inst = 32'h8220000;
      29746: inst = 32'h10408000;
      29747: inst = 32'hc4042a4;
      29748: inst = 32'h8220000;
      29749: inst = 32'h10408000;
      29750: inst = 32'hc4042a5;
      29751: inst = 32'h8220000;
      29752: inst = 32'h10408000;
      29753: inst = 32'hc4042a6;
      29754: inst = 32'h8220000;
      29755: inst = 32'h10408000;
      29756: inst = 32'hc4042a7;
      29757: inst = 32'h8220000;
      29758: inst = 32'h10408000;
      29759: inst = 32'hc4042a8;
      29760: inst = 32'h8220000;
      29761: inst = 32'h10408000;
      29762: inst = 32'hc4042a9;
      29763: inst = 32'h8220000;
      29764: inst = 32'h10408000;
      29765: inst = 32'hc4042aa;
      29766: inst = 32'h8220000;
      29767: inst = 32'h10408000;
      29768: inst = 32'hc4042ab;
      29769: inst = 32'h8220000;
      29770: inst = 32'h10408000;
      29771: inst = 32'hc4042ac;
      29772: inst = 32'h8220000;
      29773: inst = 32'h10408000;
      29774: inst = 32'hc4042ad;
      29775: inst = 32'h8220000;
      29776: inst = 32'h10408000;
      29777: inst = 32'hc4042ae;
      29778: inst = 32'h8220000;
      29779: inst = 32'h10408000;
      29780: inst = 32'hc4042af;
      29781: inst = 32'h8220000;
      29782: inst = 32'h10408000;
      29783: inst = 32'hc4042b0;
      29784: inst = 32'h8220000;
      29785: inst = 32'h10408000;
      29786: inst = 32'hc4042b1;
      29787: inst = 32'h8220000;
      29788: inst = 32'h10408000;
      29789: inst = 32'hc4042b2;
      29790: inst = 32'h8220000;
      29791: inst = 32'h10408000;
      29792: inst = 32'hc4042b3;
      29793: inst = 32'h8220000;
      29794: inst = 32'h10408000;
      29795: inst = 32'hc4042b4;
      29796: inst = 32'h8220000;
      29797: inst = 32'h10408000;
      29798: inst = 32'hc4042b5;
      29799: inst = 32'h8220000;
      29800: inst = 32'h10408000;
      29801: inst = 32'hc4042b6;
      29802: inst = 32'h8220000;
      29803: inst = 32'h10408000;
      29804: inst = 32'hc4042b7;
      29805: inst = 32'h8220000;
      29806: inst = 32'h10408000;
      29807: inst = 32'hc4042b8;
      29808: inst = 32'h8220000;
      29809: inst = 32'h10408000;
      29810: inst = 32'hc4042b9;
      29811: inst = 32'h8220000;
      29812: inst = 32'h10408000;
      29813: inst = 32'hc4042ba;
      29814: inst = 32'h8220000;
      29815: inst = 32'h10408000;
      29816: inst = 32'hc4042bb;
      29817: inst = 32'h8220000;
      29818: inst = 32'h10408000;
      29819: inst = 32'hc4042bc;
      29820: inst = 32'h8220000;
      29821: inst = 32'h10408000;
      29822: inst = 32'hc4042bd;
      29823: inst = 32'h8220000;
      29824: inst = 32'h10408000;
      29825: inst = 32'hc4042be;
      29826: inst = 32'h8220000;
      29827: inst = 32'h10408000;
      29828: inst = 32'hc4042bf;
      29829: inst = 32'h8220000;
      29830: inst = 32'h10408000;
      29831: inst = 32'hc4042c0;
      29832: inst = 32'h8220000;
      29833: inst = 32'h10408000;
      29834: inst = 32'hc4042c1;
      29835: inst = 32'h8220000;
      29836: inst = 32'h10408000;
      29837: inst = 32'hc4042c2;
      29838: inst = 32'h8220000;
      29839: inst = 32'h10408000;
      29840: inst = 32'hc4042c3;
      29841: inst = 32'h8220000;
      29842: inst = 32'h10408000;
      29843: inst = 32'hc4042c4;
      29844: inst = 32'h8220000;
      29845: inst = 32'h10408000;
      29846: inst = 32'hc4042c5;
      29847: inst = 32'h8220000;
      29848: inst = 32'h10408000;
      29849: inst = 32'hc4042c6;
      29850: inst = 32'h8220000;
      29851: inst = 32'h10408000;
      29852: inst = 32'hc4042c7;
      29853: inst = 32'h8220000;
      29854: inst = 32'h10408000;
      29855: inst = 32'hc4042c8;
      29856: inst = 32'h8220000;
      29857: inst = 32'h10408000;
      29858: inst = 32'hc4042c9;
      29859: inst = 32'h8220000;
      29860: inst = 32'h10408000;
      29861: inst = 32'hc4042ca;
      29862: inst = 32'h8220000;
      29863: inst = 32'h10408000;
      29864: inst = 32'hc4042cb;
      29865: inst = 32'h8220000;
      29866: inst = 32'h10408000;
      29867: inst = 32'hc4042cf;
      29868: inst = 32'h8220000;
      29869: inst = 32'h10408000;
      29870: inst = 32'hc4042d3;
      29871: inst = 32'h8220000;
      29872: inst = 32'h10408000;
      29873: inst = 32'hc4042da;
      29874: inst = 32'h8220000;
      29875: inst = 32'h10408000;
      29876: inst = 32'hc4042db;
      29877: inst = 32'h8220000;
      29878: inst = 32'h10408000;
      29879: inst = 32'hc4042e3;
      29880: inst = 32'h8220000;
      29881: inst = 32'h10408000;
      29882: inst = 32'hc4042ed;
      29883: inst = 32'h8220000;
      29884: inst = 32'h10408000;
      29885: inst = 32'hc4042ee;
      29886: inst = 32'h8220000;
      29887: inst = 32'h10408000;
      29888: inst = 32'hc4042ef;
      29889: inst = 32'h8220000;
      29890: inst = 32'h10408000;
      29891: inst = 32'hc4042f0;
      29892: inst = 32'h8220000;
      29893: inst = 32'h10408000;
      29894: inst = 32'hc4042f1;
      29895: inst = 32'h8220000;
      29896: inst = 32'h10408000;
      29897: inst = 32'hc4042f2;
      29898: inst = 32'h8220000;
      29899: inst = 32'h10408000;
      29900: inst = 32'hc4042f3;
      29901: inst = 32'h8220000;
      29902: inst = 32'h10408000;
      29903: inst = 32'hc4042f4;
      29904: inst = 32'h8220000;
      29905: inst = 32'h10408000;
      29906: inst = 32'hc4042f5;
      29907: inst = 32'h8220000;
      29908: inst = 32'h10408000;
      29909: inst = 32'hc4042f6;
      29910: inst = 32'h8220000;
      29911: inst = 32'h10408000;
      29912: inst = 32'hc4042f7;
      29913: inst = 32'h8220000;
      29914: inst = 32'h10408000;
      29915: inst = 32'hc4042f8;
      29916: inst = 32'h8220000;
      29917: inst = 32'h10408000;
      29918: inst = 32'hc4042f9;
      29919: inst = 32'h8220000;
      29920: inst = 32'h10408000;
      29921: inst = 32'hc4042fa;
      29922: inst = 32'h8220000;
      29923: inst = 32'h10408000;
      29924: inst = 32'hc4042fb;
      29925: inst = 32'h8220000;
      29926: inst = 32'h10408000;
      29927: inst = 32'hc4042fc;
      29928: inst = 32'h8220000;
      29929: inst = 32'h10408000;
      29930: inst = 32'hc4042fd;
      29931: inst = 32'h8220000;
      29932: inst = 32'h10408000;
      29933: inst = 32'hc4042fe;
      29934: inst = 32'h8220000;
      29935: inst = 32'h10408000;
      29936: inst = 32'hc4042ff;
      29937: inst = 32'h8220000;
      29938: inst = 32'h10408000;
      29939: inst = 32'hc404300;
      29940: inst = 32'h8220000;
      29941: inst = 32'h10408000;
      29942: inst = 32'hc404301;
      29943: inst = 32'h8220000;
      29944: inst = 32'h10408000;
      29945: inst = 32'hc404302;
      29946: inst = 32'h8220000;
      29947: inst = 32'h10408000;
      29948: inst = 32'hc404303;
      29949: inst = 32'h8220000;
      29950: inst = 32'h10408000;
      29951: inst = 32'hc404304;
      29952: inst = 32'h8220000;
      29953: inst = 32'h10408000;
      29954: inst = 32'hc404305;
      29955: inst = 32'h8220000;
      29956: inst = 32'h10408000;
      29957: inst = 32'hc404306;
      29958: inst = 32'h8220000;
      29959: inst = 32'h10408000;
      29960: inst = 32'hc404307;
      29961: inst = 32'h8220000;
      29962: inst = 32'h10408000;
      29963: inst = 32'hc404308;
      29964: inst = 32'h8220000;
      29965: inst = 32'h10408000;
      29966: inst = 32'hc404309;
      29967: inst = 32'h8220000;
      29968: inst = 32'h10408000;
      29969: inst = 32'hc40430a;
      29970: inst = 32'h8220000;
      29971: inst = 32'h10408000;
      29972: inst = 32'hc40430b;
      29973: inst = 32'h8220000;
      29974: inst = 32'h10408000;
      29975: inst = 32'hc40430c;
      29976: inst = 32'h8220000;
      29977: inst = 32'h10408000;
      29978: inst = 32'hc40430d;
      29979: inst = 32'h8220000;
      29980: inst = 32'h10408000;
      29981: inst = 32'hc40430e;
      29982: inst = 32'h8220000;
      29983: inst = 32'h10408000;
      29984: inst = 32'hc40430f;
      29985: inst = 32'h8220000;
      29986: inst = 32'h10408000;
      29987: inst = 32'hc404310;
      29988: inst = 32'h8220000;
      29989: inst = 32'h10408000;
      29990: inst = 32'hc404311;
      29991: inst = 32'h8220000;
      29992: inst = 32'h10408000;
      29993: inst = 32'hc404312;
      29994: inst = 32'h8220000;
      29995: inst = 32'h10408000;
      29996: inst = 32'hc404313;
      29997: inst = 32'h8220000;
      29998: inst = 32'h10408000;
      29999: inst = 32'hc404314;
      30000: inst = 32'h8220000;
      30001: inst = 32'h10408000;
      30002: inst = 32'hc404315;
      30003: inst = 32'h8220000;
      30004: inst = 32'h10408000;
      30005: inst = 32'hc404316;
      30006: inst = 32'h8220000;
      30007: inst = 32'h10408000;
      30008: inst = 32'hc404317;
      30009: inst = 32'h8220000;
      30010: inst = 32'h10408000;
      30011: inst = 32'hc404318;
      30012: inst = 32'h8220000;
      30013: inst = 32'h10408000;
      30014: inst = 32'hc404319;
      30015: inst = 32'h8220000;
      30016: inst = 32'h10408000;
      30017: inst = 32'hc40431a;
      30018: inst = 32'h8220000;
      30019: inst = 32'h10408000;
      30020: inst = 32'hc40431b;
      30021: inst = 32'h8220000;
      30022: inst = 32'h10408000;
      30023: inst = 32'hc40431c;
      30024: inst = 32'h8220000;
      30025: inst = 32'h10408000;
      30026: inst = 32'hc40431d;
      30027: inst = 32'h8220000;
      30028: inst = 32'h10408000;
      30029: inst = 32'hc40431e;
      30030: inst = 32'h8220000;
      30031: inst = 32'h10408000;
      30032: inst = 32'hc40431f;
      30033: inst = 32'h8220000;
      30034: inst = 32'h10408000;
      30035: inst = 32'hc404320;
      30036: inst = 32'h8220000;
      30037: inst = 32'h10408000;
      30038: inst = 32'hc404321;
      30039: inst = 32'h8220000;
      30040: inst = 32'h10408000;
      30041: inst = 32'hc404322;
      30042: inst = 32'h8220000;
      30043: inst = 32'h10408000;
      30044: inst = 32'hc404323;
      30045: inst = 32'h8220000;
      30046: inst = 32'h10408000;
      30047: inst = 32'hc404324;
      30048: inst = 32'h8220000;
      30049: inst = 32'h10408000;
      30050: inst = 32'hc404325;
      30051: inst = 32'h8220000;
      30052: inst = 32'h10408000;
      30053: inst = 32'hc404326;
      30054: inst = 32'h8220000;
      30055: inst = 32'h10408000;
      30056: inst = 32'hc404327;
      30057: inst = 32'h8220000;
      30058: inst = 32'h10408000;
      30059: inst = 32'hc404328;
      30060: inst = 32'h8220000;
      30061: inst = 32'h10408000;
      30062: inst = 32'hc404329;
      30063: inst = 32'h8220000;
      30064: inst = 32'h10408000;
      30065: inst = 32'hc40432a;
      30066: inst = 32'h8220000;
      30067: inst = 32'h10408000;
      30068: inst = 32'hc40432b;
      30069: inst = 32'h8220000;
      30070: inst = 32'h10408000;
      30071: inst = 32'hc40432f;
      30072: inst = 32'h8220000;
      30073: inst = 32'h10408000;
      30074: inst = 32'hc404330;
      30075: inst = 32'h8220000;
      30076: inst = 32'h10408000;
      30077: inst = 32'hc404333;
      30078: inst = 32'h8220000;
      30079: inst = 32'h10408000;
      30080: inst = 32'hc404334;
      30081: inst = 32'h8220000;
      30082: inst = 32'h10408000;
      30083: inst = 32'hc404343;
      30084: inst = 32'h8220000;
      30085: inst = 32'h10408000;
      30086: inst = 32'hc40434d;
      30087: inst = 32'h8220000;
      30088: inst = 32'h10408000;
      30089: inst = 32'hc40434e;
      30090: inst = 32'h8220000;
      30091: inst = 32'h10408000;
      30092: inst = 32'hc40434f;
      30093: inst = 32'h8220000;
      30094: inst = 32'h10408000;
      30095: inst = 32'hc404350;
      30096: inst = 32'h8220000;
      30097: inst = 32'h10408000;
      30098: inst = 32'hc404351;
      30099: inst = 32'h8220000;
      30100: inst = 32'h10408000;
      30101: inst = 32'hc404352;
      30102: inst = 32'h8220000;
      30103: inst = 32'h10408000;
      30104: inst = 32'hc404353;
      30105: inst = 32'h8220000;
      30106: inst = 32'h10408000;
      30107: inst = 32'hc404354;
      30108: inst = 32'h8220000;
      30109: inst = 32'h10408000;
      30110: inst = 32'hc404355;
      30111: inst = 32'h8220000;
      30112: inst = 32'h10408000;
      30113: inst = 32'hc404356;
      30114: inst = 32'h8220000;
      30115: inst = 32'h10408000;
      30116: inst = 32'hc404357;
      30117: inst = 32'h8220000;
      30118: inst = 32'h10408000;
      30119: inst = 32'hc404358;
      30120: inst = 32'h8220000;
      30121: inst = 32'h10408000;
      30122: inst = 32'hc404359;
      30123: inst = 32'h8220000;
      30124: inst = 32'h10408000;
      30125: inst = 32'hc40435a;
      30126: inst = 32'h8220000;
      30127: inst = 32'h10408000;
      30128: inst = 32'hc40435b;
      30129: inst = 32'h8220000;
      30130: inst = 32'h10408000;
      30131: inst = 32'hc40435c;
      30132: inst = 32'h8220000;
      30133: inst = 32'h10408000;
      30134: inst = 32'hc40435d;
      30135: inst = 32'h8220000;
      30136: inst = 32'h10408000;
      30137: inst = 32'hc40435e;
      30138: inst = 32'h8220000;
      30139: inst = 32'h10408000;
      30140: inst = 32'hc40435f;
      30141: inst = 32'h8220000;
      30142: inst = 32'h10408000;
      30143: inst = 32'hc404360;
      30144: inst = 32'h8220000;
      30145: inst = 32'h10408000;
      30146: inst = 32'hc404361;
      30147: inst = 32'h8220000;
      30148: inst = 32'h10408000;
      30149: inst = 32'hc404362;
      30150: inst = 32'h8220000;
      30151: inst = 32'h10408000;
      30152: inst = 32'hc404363;
      30153: inst = 32'h8220000;
      30154: inst = 32'h10408000;
      30155: inst = 32'hc404364;
      30156: inst = 32'h8220000;
      30157: inst = 32'h10408000;
      30158: inst = 32'hc404365;
      30159: inst = 32'h8220000;
      30160: inst = 32'h10408000;
      30161: inst = 32'hc404366;
      30162: inst = 32'h8220000;
      30163: inst = 32'h10408000;
      30164: inst = 32'hc404367;
      30165: inst = 32'h8220000;
      30166: inst = 32'h10408000;
      30167: inst = 32'hc404368;
      30168: inst = 32'h8220000;
      30169: inst = 32'h10408000;
      30170: inst = 32'hc404369;
      30171: inst = 32'h8220000;
      30172: inst = 32'h10408000;
      30173: inst = 32'hc40436a;
      30174: inst = 32'h8220000;
      30175: inst = 32'h10408000;
      30176: inst = 32'hc40436b;
      30177: inst = 32'h8220000;
      30178: inst = 32'h10408000;
      30179: inst = 32'hc40436c;
      30180: inst = 32'h8220000;
      30181: inst = 32'h10408000;
      30182: inst = 32'hc40436d;
      30183: inst = 32'h8220000;
      30184: inst = 32'h10408000;
      30185: inst = 32'hc40436e;
      30186: inst = 32'h8220000;
      30187: inst = 32'h10408000;
      30188: inst = 32'hc40436f;
      30189: inst = 32'h8220000;
      30190: inst = 32'h10408000;
      30191: inst = 32'hc404370;
      30192: inst = 32'h8220000;
      30193: inst = 32'h10408000;
      30194: inst = 32'hc404371;
      30195: inst = 32'h8220000;
      30196: inst = 32'h10408000;
      30197: inst = 32'hc404372;
      30198: inst = 32'h8220000;
      30199: inst = 32'h10408000;
      30200: inst = 32'hc404373;
      30201: inst = 32'h8220000;
      30202: inst = 32'h10408000;
      30203: inst = 32'hc404374;
      30204: inst = 32'h8220000;
      30205: inst = 32'h10408000;
      30206: inst = 32'hc404375;
      30207: inst = 32'h8220000;
      30208: inst = 32'h10408000;
      30209: inst = 32'hc404376;
      30210: inst = 32'h8220000;
      30211: inst = 32'h10408000;
      30212: inst = 32'hc404377;
      30213: inst = 32'h8220000;
      30214: inst = 32'h10408000;
      30215: inst = 32'hc404378;
      30216: inst = 32'h8220000;
      30217: inst = 32'h10408000;
      30218: inst = 32'hc404379;
      30219: inst = 32'h8220000;
      30220: inst = 32'h10408000;
      30221: inst = 32'hc40437a;
      30222: inst = 32'h8220000;
      30223: inst = 32'h10408000;
      30224: inst = 32'hc40437b;
      30225: inst = 32'h8220000;
      30226: inst = 32'h10408000;
      30227: inst = 32'hc40437c;
      30228: inst = 32'h8220000;
      30229: inst = 32'h10408000;
      30230: inst = 32'hc40437d;
      30231: inst = 32'h8220000;
      30232: inst = 32'h10408000;
      30233: inst = 32'hc40437e;
      30234: inst = 32'h8220000;
      30235: inst = 32'h10408000;
      30236: inst = 32'hc40437f;
      30237: inst = 32'h8220000;
      30238: inst = 32'h10408000;
      30239: inst = 32'hc404380;
      30240: inst = 32'h8220000;
      30241: inst = 32'h10408000;
      30242: inst = 32'hc404381;
      30243: inst = 32'h8220000;
      30244: inst = 32'h10408000;
      30245: inst = 32'hc404382;
      30246: inst = 32'h8220000;
      30247: inst = 32'h10408000;
      30248: inst = 32'hc404383;
      30249: inst = 32'h8220000;
      30250: inst = 32'h10408000;
      30251: inst = 32'hc404384;
      30252: inst = 32'h8220000;
      30253: inst = 32'h10408000;
      30254: inst = 32'hc404385;
      30255: inst = 32'h8220000;
      30256: inst = 32'h10408000;
      30257: inst = 32'hc404386;
      30258: inst = 32'h8220000;
      30259: inst = 32'h10408000;
      30260: inst = 32'hc404387;
      30261: inst = 32'h8220000;
      30262: inst = 32'h10408000;
      30263: inst = 32'hc404388;
      30264: inst = 32'h8220000;
      30265: inst = 32'h10408000;
      30266: inst = 32'hc404389;
      30267: inst = 32'h8220000;
      30268: inst = 32'h10408000;
      30269: inst = 32'hc40438a;
      30270: inst = 32'h8220000;
      30271: inst = 32'h10408000;
      30272: inst = 32'hc40438b;
      30273: inst = 32'h8220000;
      30274: inst = 32'h10408000;
      30275: inst = 32'hc40438f;
      30276: inst = 32'h8220000;
      30277: inst = 32'h10408000;
      30278: inst = 32'hc404390;
      30279: inst = 32'h8220000;
      30280: inst = 32'h10408000;
      30281: inst = 32'hc4043a3;
      30282: inst = 32'h8220000;
      30283: inst = 32'h10408000;
      30284: inst = 32'hc4043ad;
      30285: inst = 32'h8220000;
      30286: inst = 32'h10408000;
      30287: inst = 32'hc4043ae;
      30288: inst = 32'h8220000;
      30289: inst = 32'h10408000;
      30290: inst = 32'hc4043af;
      30291: inst = 32'h8220000;
      30292: inst = 32'h10408000;
      30293: inst = 32'hc4043b0;
      30294: inst = 32'h8220000;
      30295: inst = 32'h10408000;
      30296: inst = 32'hc4043b1;
      30297: inst = 32'h8220000;
      30298: inst = 32'h10408000;
      30299: inst = 32'hc4043b2;
      30300: inst = 32'h8220000;
      30301: inst = 32'h10408000;
      30302: inst = 32'hc4043b3;
      30303: inst = 32'h8220000;
      30304: inst = 32'h10408000;
      30305: inst = 32'hc4043b4;
      30306: inst = 32'h8220000;
      30307: inst = 32'h10408000;
      30308: inst = 32'hc4043b5;
      30309: inst = 32'h8220000;
      30310: inst = 32'h10408000;
      30311: inst = 32'hc4043b6;
      30312: inst = 32'h8220000;
      30313: inst = 32'h10408000;
      30314: inst = 32'hc4043b7;
      30315: inst = 32'h8220000;
      30316: inst = 32'h10408000;
      30317: inst = 32'hc4043b8;
      30318: inst = 32'h8220000;
      30319: inst = 32'h10408000;
      30320: inst = 32'hc4043b9;
      30321: inst = 32'h8220000;
      30322: inst = 32'h10408000;
      30323: inst = 32'hc4043ba;
      30324: inst = 32'h8220000;
      30325: inst = 32'h10408000;
      30326: inst = 32'hc4043bb;
      30327: inst = 32'h8220000;
      30328: inst = 32'h10408000;
      30329: inst = 32'hc4043bc;
      30330: inst = 32'h8220000;
      30331: inst = 32'h10408000;
      30332: inst = 32'hc4043bd;
      30333: inst = 32'h8220000;
      30334: inst = 32'h10408000;
      30335: inst = 32'hc4043be;
      30336: inst = 32'h8220000;
      30337: inst = 32'h10408000;
      30338: inst = 32'hc4043bf;
      30339: inst = 32'h8220000;
      30340: inst = 32'h10408000;
      30341: inst = 32'hc4043c0;
      30342: inst = 32'h8220000;
      30343: inst = 32'h10408000;
      30344: inst = 32'hc4043c1;
      30345: inst = 32'h8220000;
      30346: inst = 32'h10408000;
      30347: inst = 32'hc4043c2;
      30348: inst = 32'h8220000;
      30349: inst = 32'h10408000;
      30350: inst = 32'hc4043c3;
      30351: inst = 32'h8220000;
      30352: inst = 32'h10408000;
      30353: inst = 32'hc4043c4;
      30354: inst = 32'h8220000;
      30355: inst = 32'h10408000;
      30356: inst = 32'hc4043c5;
      30357: inst = 32'h8220000;
      30358: inst = 32'h10408000;
      30359: inst = 32'hc4043c6;
      30360: inst = 32'h8220000;
      30361: inst = 32'h10408000;
      30362: inst = 32'hc4043c7;
      30363: inst = 32'h8220000;
      30364: inst = 32'h10408000;
      30365: inst = 32'hc4043c8;
      30366: inst = 32'h8220000;
      30367: inst = 32'h10408000;
      30368: inst = 32'hc4043c9;
      30369: inst = 32'h8220000;
      30370: inst = 32'h10408000;
      30371: inst = 32'hc4043ca;
      30372: inst = 32'h8220000;
      30373: inst = 32'h10408000;
      30374: inst = 32'hc4043cb;
      30375: inst = 32'h8220000;
      30376: inst = 32'h10408000;
      30377: inst = 32'hc4043cc;
      30378: inst = 32'h8220000;
      30379: inst = 32'h10408000;
      30380: inst = 32'hc4043cd;
      30381: inst = 32'h8220000;
      30382: inst = 32'h10408000;
      30383: inst = 32'hc4043ce;
      30384: inst = 32'h8220000;
      30385: inst = 32'h10408000;
      30386: inst = 32'hc4043cf;
      30387: inst = 32'h8220000;
      30388: inst = 32'h10408000;
      30389: inst = 32'hc4043d0;
      30390: inst = 32'h8220000;
      30391: inst = 32'h10408000;
      30392: inst = 32'hc4043d1;
      30393: inst = 32'h8220000;
      30394: inst = 32'h10408000;
      30395: inst = 32'hc4043d2;
      30396: inst = 32'h8220000;
      30397: inst = 32'h10408000;
      30398: inst = 32'hc4043d3;
      30399: inst = 32'h8220000;
      30400: inst = 32'h10408000;
      30401: inst = 32'hc4043d4;
      30402: inst = 32'h8220000;
      30403: inst = 32'h10408000;
      30404: inst = 32'hc4043d5;
      30405: inst = 32'h8220000;
      30406: inst = 32'h10408000;
      30407: inst = 32'hc4043d6;
      30408: inst = 32'h8220000;
      30409: inst = 32'h10408000;
      30410: inst = 32'hc4043d7;
      30411: inst = 32'h8220000;
      30412: inst = 32'h10408000;
      30413: inst = 32'hc4043d8;
      30414: inst = 32'h8220000;
      30415: inst = 32'h10408000;
      30416: inst = 32'hc4043d9;
      30417: inst = 32'h8220000;
      30418: inst = 32'h10408000;
      30419: inst = 32'hc4043da;
      30420: inst = 32'h8220000;
      30421: inst = 32'h10408000;
      30422: inst = 32'hc4043db;
      30423: inst = 32'h8220000;
      30424: inst = 32'h10408000;
      30425: inst = 32'hc4043dc;
      30426: inst = 32'h8220000;
      30427: inst = 32'h10408000;
      30428: inst = 32'hc4043dd;
      30429: inst = 32'h8220000;
      30430: inst = 32'h10408000;
      30431: inst = 32'hc4043de;
      30432: inst = 32'h8220000;
      30433: inst = 32'h10408000;
      30434: inst = 32'hc4043df;
      30435: inst = 32'h8220000;
      30436: inst = 32'h10408000;
      30437: inst = 32'hc4043e0;
      30438: inst = 32'h8220000;
      30439: inst = 32'h10408000;
      30440: inst = 32'hc4043e1;
      30441: inst = 32'h8220000;
      30442: inst = 32'h10408000;
      30443: inst = 32'hc4043e2;
      30444: inst = 32'h8220000;
      30445: inst = 32'h10408000;
      30446: inst = 32'hc4043e3;
      30447: inst = 32'h8220000;
      30448: inst = 32'h10408000;
      30449: inst = 32'hc4043e4;
      30450: inst = 32'h8220000;
      30451: inst = 32'h10408000;
      30452: inst = 32'hc4043e5;
      30453: inst = 32'h8220000;
      30454: inst = 32'h10408000;
      30455: inst = 32'hc4043e6;
      30456: inst = 32'h8220000;
      30457: inst = 32'h10408000;
      30458: inst = 32'hc4043e7;
      30459: inst = 32'h8220000;
      30460: inst = 32'h10408000;
      30461: inst = 32'hc4043e8;
      30462: inst = 32'h8220000;
      30463: inst = 32'h10408000;
      30464: inst = 32'hc4043e9;
      30465: inst = 32'h8220000;
      30466: inst = 32'h10408000;
      30467: inst = 32'hc4043ea;
      30468: inst = 32'h8220000;
      30469: inst = 32'h10408000;
      30470: inst = 32'hc4043eb;
      30471: inst = 32'h8220000;
      30472: inst = 32'h10408000;
      30473: inst = 32'hc4043ef;
      30474: inst = 32'h8220000;
      30475: inst = 32'h10408000;
      30476: inst = 32'hc4043f9;
      30477: inst = 32'h8220000;
      30478: inst = 32'h10408000;
      30479: inst = 32'hc404403;
      30480: inst = 32'h8220000;
      30481: inst = 32'h10408000;
      30482: inst = 32'hc404404;
      30483: inst = 32'h8220000;
      30484: inst = 32'h10408000;
      30485: inst = 32'hc404405;
      30486: inst = 32'h8220000;
      30487: inst = 32'h10408000;
      30488: inst = 32'hc404406;
      30489: inst = 32'h8220000;
      30490: inst = 32'h10408000;
      30491: inst = 32'hc404407;
      30492: inst = 32'h8220000;
      30493: inst = 32'h10408000;
      30494: inst = 32'hc404408;
      30495: inst = 32'h8220000;
      30496: inst = 32'h10408000;
      30497: inst = 32'hc404409;
      30498: inst = 32'h8220000;
      30499: inst = 32'h10408000;
      30500: inst = 32'hc40440a;
      30501: inst = 32'h8220000;
      30502: inst = 32'h10408000;
      30503: inst = 32'hc40440b;
      30504: inst = 32'h8220000;
      30505: inst = 32'h10408000;
      30506: inst = 32'hc40440c;
      30507: inst = 32'h8220000;
      30508: inst = 32'h10408000;
      30509: inst = 32'hc40440d;
      30510: inst = 32'h8220000;
      30511: inst = 32'h10408000;
      30512: inst = 32'hc40440e;
      30513: inst = 32'h8220000;
      30514: inst = 32'h10408000;
      30515: inst = 32'hc40440f;
      30516: inst = 32'h8220000;
      30517: inst = 32'h10408000;
      30518: inst = 32'hc404410;
      30519: inst = 32'h8220000;
      30520: inst = 32'h10408000;
      30521: inst = 32'hc404411;
      30522: inst = 32'h8220000;
      30523: inst = 32'h10408000;
      30524: inst = 32'hc404412;
      30525: inst = 32'h8220000;
      30526: inst = 32'h10408000;
      30527: inst = 32'hc404413;
      30528: inst = 32'h8220000;
      30529: inst = 32'h10408000;
      30530: inst = 32'hc404414;
      30531: inst = 32'h8220000;
      30532: inst = 32'h10408000;
      30533: inst = 32'hc404415;
      30534: inst = 32'h8220000;
      30535: inst = 32'h10408000;
      30536: inst = 32'hc404416;
      30537: inst = 32'h8220000;
      30538: inst = 32'h10408000;
      30539: inst = 32'hc404417;
      30540: inst = 32'h8220000;
      30541: inst = 32'h10408000;
      30542: inst = 32'hc404418;
      30543: inst = 32'h8220000;
      30544: inst = 32'h10408000;
      30545: inst = 32'hc404419;
      30546: inst = 32'h8220000;
      30547: inst = 32'h10408000;
      30548: inst = 32'hc40441a;
      30549: inst = 32'h8220000;
      30550: inst = 32'h10408000;
      30551: inst = 32'hc40441b;
      30552: inst = 32'h8220000;
      30553: inst = 32'h10408000;
      30554: inst = 32'hc40441c;
      30555: inst = 32'h8220000;
      30556: inst = 32'h10408000;
      30557: inst = 32'hc40441d;
      30558: inst = 32'h8220000;
      30559: inst = 32'h10408000;
      30560: inst = 32'hc40441e;
      30561: inst = 32'h8220000;
      30562: inst = 32'h10408000;
      30563: inst = 32'hc40441f;
      30564: inst = 32'h8220000;
      30565: inst = 32'h10408000;
      30566: inst = 32'hc404420;
      30567: inst = 32'h8220000;
      30568: inst = 32'h10408000;
      30569: inst = 32'hc404421;
      30570: inst = 32'h8220000;
      30571: inst = 32'h10408000;
      30572: inst = 32'hc404422;
      30573: inst = 32'h8220000;
      30574: inst = 32'h10408000;
      30575: inst = 32'hc404423;
      30576: inst = 32'h8220000;
      30577: inst = 32'h10408000;
      30578: inst = 32'hc404424;
      30579: inst = 32'h8220000;
      30580: inst = 32'h10408000;
      30581: inst = 32'hc404425;
      30582: inst = 32'h8220000;
      30583: inst = 32'h10408000;
      30584: inst = 32'hc404426;
      30585: inst = 32'h8220000;
      30586: inst = 32'h10408000;
      30587: inst = 32'hc404427;
      30588: inst = 32'h8220000;
      30589: inst = 32'h10408000;
      30590: inst = 32'hc404428;
      30591: inst = 32'h8220000;
      30592: inst = 32'h10408000;
      30593: inst = 32'hc404429;
      30594: inst = 32'h8220000;
      30595: inst = 32'h10408000;
      30596: inst = 32'hc40442a;
      30597: inst = 32'h8220000;
      30598: inst = 32'h10408000;
      30599: inst = 32'hc40442b;
      30600: inst = 32'h8220000;
      30601: inst = 32'h10408000;
      30602: inst = 32'hc40442c;
      30603: inst = 32'h8220000;
      30604: inst = 32'h10408000;
      30605: inst = 32'hc40442d;
      30606: inst = 32'h8220000;
      30607: inst = 32'h10408000;
      30608: inst = 32'hc40442e;
      30609: inst = 32'h8220000;
      30610: inst = 32'h10408000;
      30611: inst = 32'hc40442f;
      30612: inst = 32'h8220000;
      30613: inst = 32'h10408000;
      30614: inst = 32'hc404430;
      30615: inst = 32'h8220000;
      30616: inst = 32'h10408000;
      30617: inst = 32'hc404431;
      30618: inst = 32'h8220000;
      30619: inst = 32'h10408000;
      30620: inst = 32'hc404432;
      30621: inst = 32'h8220000;
      30622: inst = 32'h10408000;
      30623: inst = 32'hc404433;
      30624: inst = 32'h8220000;
      30625: inst = 32'h10408000;
      30626: inst = 32'hc404434;
      30627: inst = 32'h8220000;
      30628: inst = 32'h10408000;
      30629: inst = 32'hc404435;
      30630: inst = 32'h8220000;
      30631: inst = 32'h10408000;
      30632: inst = 32'hc404436;
      30633: inst = 32'h8220000;
      30634: inst = 32'h10408000;
      30635: inst = 32'hc404437;
      30636: inst = 32'h8220000;
      30637: inst = 32'h10408000;
      30638: inst = 32'hc404438;
      30639: inst = 32'h8220000;
      30640: inst = 32'h10408000;
      30641: inst = 32'hc404439;
      30642: inst = 32'h8220000;
      30643: inst = 32'h10408000;
      30644: inst = 32'hc40443a;
      30645: inst = 32'h8220000;
      30646: inst = 32'h10408000;
      30647: inst = 32'hc40443b;
      30648: inst = 32'h8220000;
      30649: inst = 32'h10408000;
      30650: inst = 32'hc40443c;
      30651: inst = 32'h8220000;
      30652: inst = 32'h10408000;
      30653: inst = 32'hc40443d;
      30654: inst = 32'h8220000;
      30655: inst = 32'h10408000;
      30656: inst = 32'hc40443e;
      30657: inst = 32'h8220000;
      30658: inst = 32'h10408000;
      30659: inst = 32'hc40443f;
      30660: inst = 32'h8220000;
      30661: inst = 32'h10408000;
      30662: inst = 32'hc404440;
      30663: inst = 32'h8220000;
      30664: inst = 32'h10408000;
      30665: inst = 32'hc404441;
      30666: inst = 32'h8220000;
      30667: inst = 32'h10408000;
      30668: inst = 32'hc404442;
      30669: inst = 32'h8220000;
      30670: inst = 32'h10408000;
      30671: inst = 32'hc404443;
      30672: inst = 32'h8220000;
      30673: inst = 32'h10408000;
      30674: inst = 32'hc404444;
      30675: inst = 32'h8220000;
      30676: inst = 32'h10408000;
      30677: inst = 32'hc404445;
      30678: inst = 32'h8220000;
      30679: inst = 32'h10408000;
      30680: inst = 32'hc404446;
      30681: inst = 32'h8220000;
      30682: inst = 32'h10408000;
      30683: inst = 32'hc404447;
      30684: inst = 32'h8220000;
      30685: inst = 32'h10408000;
      30686: inst = 32'hc404448;
      30687: inst = 32'h8220000;
      30688: inst = 32'h10408000;
      30689: inst = 32'hc404449;
      30690: inst = 32'h8220000;
      30691: inst = 32'h10408000;
      30692: inst = 32'hc40444a;
      30693: inst = 32'h8220000;
      30694: inst = 32'h10408000;
      30695: inst = 32'hc40444b;
      30696: inst = 32'h8220000;
      30697: inst = 32'h10408000;
      30698: inst = 32'hc40444f;
      30699: inst = 32'h8220000;
      30700: inst = 32'h10408000;
      30701: inst = 32'hc404455;
      30702: inst = 32'h8220000;
      30703: inst = 32'h10408000;
      30704: inst = 32'hc404463;
      30705: inst = 32'h8220000;
      30706: inst = 32'h10408000;
      30707: inst = 32'hc404464;
      30708: inst = 32'h8220000;
      30709: inst = 32'h10408000;
      30710: inst = 32'hc404465;
      30711: inst = 32'h8220000;
      30712: inst = 32'h10408000;
      30713: inst = 32'hc404466;
      30714: inst = 32'h8220000;
      30715: inst = 32'h10408000;
      30716: inst = 32'hc404467;
      30717: inst = 32'h8220000;
      30718: inst = 32'h10408000;
      30719: inst = 32'hc404468;
      30720: inst = 32'h8220000;
      30721: inst = 32'h10408000;
      30722: inst = 32'hc404469;
      30723: inst = 32'h8220000;
      30724: inst = 32'h10408000;
      30725: inst = 32'hc40446a;
      30726: inst = 32'h8220000;
      30727: inst = 32'h10408000;
      30728: inst = 32'hc40446b;
      30729: inst = 32'h8220000;
      30730: inst = 32'h10408000;
      30731: inst = 32'hc40446c;
      30732: inst = 32'h8220000;
      30733: inst = 32'h10408000;
      30734: inst = 32'hc40446d;
      30735: inst = 32'h8220000;
      30736: inst = 32'h10408000;
      30737: inst = 32'hc40446e;
      30738: inst = 32'h8220000;
      30739: inst = 32'h10408000;
      30740: inst = 32'hc40446f;
      30741: inst = 32'h8220000;
      30742: inst = 32'h10408000;
      30743: inst = 32'hc404470;
      30744: inst = 32'h8220000;
      30745: inst = 32'h10408000;
      30746: inst = 32'hc404471;
      30747: inst = 32'h8220000;
      30748: inst = 32'h10408000;
      30749: inst = 32'hc404472;
      30750: inst = 32'h8220000;
      30751: inst = 32'h10408000;
      30752: inst = 32'hc404473;
      30753: inst = 32'h8220000;
      30754: inst = 32'h10408000;
      30755: inst = 32'hc404474;
      30756: inst = 32'h8220000;
      30757: inst = 32'h10408000;
      30758: inst = 32'hc404475;
      30759: inst = 32'h8220000;
      30760: inst = 32'h10408000;
      30761: inst = 32'hc404476;
      30762: inst = 32'h8220000;
      30763: inst = 32'h10408000;
      30764: inst = 32'hc404477;
      30765: inst = 32'h8220000;
      30766: inst = 32'h10408000;
      30767: inst = 32'hc404478;
      30768: inst = 32'h8220000;
      30769: inst = 32'h10408000;
      30770: inst = 32'hc404479;
      30771: inst = 32'h8220000;
      30772: inst = 32'h10408000;
      30773: inst = 32'hc40447a;
      30774: inst = 32'h8220000;
      30775: inst = 32'h10408000;
      30776: inst = 32'hc40447b;
      30777: inst = 32'h8220000;
      30778: inst = 32'h10408000;
      30779: inst = 32'hc40447c;
      30780: inst = 32'h8220000;
      30781: inst = 32'h10408000;
      30782: inst = 32'hc40447d;
      30783: inst = 32'h8220000;
      30784: inst = 32'h10408000;
      30785: inst = 32'hc40447e;
      30786: inst = 32'h8220000;
      30787: inst = 32'h10408000;
      30788: inst = 32'hc40447f;
      30789: inst = 32'h8220000;
      30790: inst = 32'h10408000;
      30791: inst = 32'hc404480;
      30792: inst = 32'h8220000;
      30793: inst = 32'h10408000;
      30794: inst = 32'hc404481;
      30795: inst = 32'h8220000;
      30796: inst = 32'h10408000;
      30797: inst = 32'hc404482;
      30798: inst = 32'h8220000;
      30799: inst = 32'h10408000;
      30800: inst = 32'hc404483;
      30801: inst = 32'h8220000;
      30802: inst = 32'h10408000;
      30803: inst = 32'hc404484;
      30804: inst = 32'h8220000;
      30805: inst = 32'h10408000;
      30806: inst = 32'hc404485;
      30807: inst = 32'h8220000;
      30808: inst = 32'h10408000;
      30809: inst = 32'hc404486;
      30810: inst = 32'h8220000;
      30811: inst = 32'h10408000;
      30812: inst = 32'hc404487;
      30813: inst = 32'h8220000;
      30814: inst = 32'h10408000;
      30815: inst = 32'hc404488;
      30816: inst = 32'h8220000;
      30817: inst = 32'h10408000;
      30818: inst = 32'hc404489;
      30819: inst = 32'h8220000;
      30820: inst = 32'h10408000;
      30821: inst = 32'hc40448a;
      30822: inst = 32'h8220000;
      30823: inst = 32'h10408000;
      30824: inst = 32'hc40448b;
      30825: inst = 32'h8220000;
      30826: inst = 32'h10408000;
      30827: inst = 32'hc40448c;
      30828: inst = 32'h8220000;
      30829: inst = 32'h10408000;
      30830: inst = 32'hc40448d;
      30831: inst = 32'h8220000;
      30832: inst = 32'h10408000;
      30833: inst = 32'hc40448e;
      30834: inst = 32'h8220000;
      30835: inst = 32'h10408000;
      30836: inst = 32'hc40448f;
      30837: inst = 32'h8220000;
      30838: inst = 32'h10408000;
      30839: inst = 32'hc404490;
      30840: inst = 32'h8220000;
      30841: inst = 32'h10408000;
      30842: inst = 32'hc404491;
      30843: inst = 32'h8220000;
      30844: inst = 32'h10408000;
      30845: inst = 32'hc404492;
      30846: inst = 32'h8220000;
      30847: inst = 32'h10408000;
      30848: inst = 32'hc404493;
      30849: inst = 32'h8220000;
      30850: inst = 32'h10408000;
      30851: inst = 32'hc404494;
      30852: inst = 32'h8220000;
      30853: inst = 32'h10408000;
      30854: inst = 32'hc404495;
      30855: inst = 32'h8220000;
      30856: inst = 32'h10408000;
      30857: inst = 32'hc404496;
      30858: inst = 32'h8220000;
      30859: inst = 32'h10408000;
      30860: inst = 32'hc404497;
      30861: inst = 32'h8220000;
      30862: inst = 32'h10408000;
      30863: inst = 32'hc404498;
      30864: inst = 32'h8220000;
      30865: inst = 32'h10408000;
      30866: inst = 32'hc404499;
      30867: inst = 32'h8220000;
      30868: inst = 32'h10408000;
      30869: inst = 32'hc40449a;
      30870: inst = 32'h8220000;
      30871: inst = 32'h10408000;
      30872: inst = 32'hc40449b;
      30873: inst = 32'h8220000;
      30874: inst = 32'h10408000;
      30875: inst = 32'hc40449c;
      30876: inst = 32'h8220000;
      30877: inst = 32'h10408000;
      30878: inst = 32'hc40449d;
      30879: inst = 32'h8220000;
      30880: inst = 32'h10408000;
      30881: inst = 32'hc40449e;
      30882: inst = 32'h8220000;
      30883: inst = 32'h10408000;
      30884: inst = 32'hc40449f;
      30885: inst = 32'h8220000;
      30886: inst = 32'h10408000;
      30887: inst = 32'hc4044a0;
      30888: inst = 32'h8220000;
      30889: inst = 32'h10408000;
      30890: inst = 32'hc4044a1;
      30891: inst = 32'h8220000;
      30892: inst = 32'h10408000;
      30893: inst = 32'hc4044a2;
      30894: inst = 32'h8220000;
      30895: inst = 32'h10408000;
      30896: inst = 32'hc4044a3;
      30897: inst = 32'h8220000;
      30898: inst = 32'h10408000;
      30899: inst = 32'hc4044a4;
      30900: inst = 32'h8220000;
      30901: inst = 32'h10408000;
      30902: inst = 32'hc4044a5;
      30903: inst = 32'h8220000;
      30904: inst = 32'h10408000;
      30905: inst = 32'hc4044a6;
      30906: inst = 32'h8220000;
      30907: inst = 32'h10408000;
      30908: inst = 32'hc4044a7;
      30909: inst = 32'h8220000;
      30910: inst = 32'h10408000;
      30911: inst = 32'hc4044a8;
      30912: inst = 32'h8220000;
      30913: inst = 32'h10408000;
      30914: inst = 32'hc4044a9;
      30915: inst = 32'h8220000;
      30916: inst = 32'h10408000;
      30917: inst = 32'hc4044aa;
      30918: inst = 32'h8220000;
      30919: inst = 32'h10408000;
      30920: inst = 32'hc4044ab;
      30921: inst = 32'h8220000;
      30922: inst = 32'h10408000;
      30923: inst = 32'hc4044af;
      30924: inst = 32'h8220000;
      30925: inst = 32'h10408000;
      30926: inst = 32'hc4044b0;
      30927: inst = 32'h8220000;
      30928: inst = 32'h10408000;
      30929: inst = 32'hc4044b1;
      30930: inst = 32'h8220000;
      30931: inst = 32'h10408000;
      30932: inst = 32'hc4044b2;
      30933: inst = 32'h8220000;
      30934: inst = 32'h10408000;
      30935: inst = 32'hc4044b7;
      30936: inst = 32'h8220000;
      30937: inst = 32'h10408000;
      30938: inst = 32'hc4044c3;
      30939: inst = 32'h8220000;
      30940: inst = 32'h10408000;
      30941: inst = 32'hc4044c4;
      30942: inst = 32'h8220000;
      30943: inst = 32'h10408000;
      30944: inst = 32'hc4044c5;
      30945: inst = 32'h8220000;
      30946: inst = 32'h10408000;
      30947: inst = 32'hc4044c6;
      30948: inst = 32'h8220000;
      30949: inst = 32'h10408000;
      30950: inst = 32'hc4044c7;
      30951: inst = 32'h8220000;
      30952: inst = 32'h10408000;
      30953: inst = 32'hc4044c8;
      30954: inst = 32'h8220000;
      30955: inst = 32'h10408000;
      30956: inst = 32'hc4044c9;
      30957: inst = 32'h8220000;
      30958: inst = 32'h10408000;
      30959: inst = 32'hc4044ca;
      30960: inst = 32'h8220000;
      30961: inst = 32'h10408000;
      30962: inst = 32'hc4044cb;
      30963: inst = 32'h8220000;
      30964: inst = 32'h10408000;
      30965: inst = 32'hc4044cc;
      30966: inst = 32'h8220000;
      30967: inst = 32'h10408000;
      30968: inst = 32'hc4044cd;
      30969: inst = 32'h8220000;
      30970: inst = 32'h10408000;
      30971: inst = 32'hc4044ce;
      30972: inst = 32'h8220000;
      30973: inst = 32'h10408000;
      30974: inst = 32'hc4044cf;
      30975: inst = 32'h8220000;
      30976: inst = 32'h10408000;
      30977: inst = 32'hc4044d0;
      30978: inst = 32'h8220000;
      30979: inst = 32'h10408000;
      30980: inst = 32'hc4044d1;
      30981: inst = 32'h8220000;
      30982: inst = 32'h10408000;
      30983: inst = 32'hc4044d2;
      30984: inst = 32'h8220000;
      30985: inst = 32'h10408000;
      30986: inst = 32'hc4044d3;
      30987: inst = 32'h8220000;
      30988: inst = 32'h10408000;
      30989: inst = 32'hc4044d4;
      30990: inst = 32'h8220000;
      30991: inst = 32'h10408000;
      30992: inst = 32'hc4044d5;
      30993: inst = 32'h8220000;
      30994: inst = 32'h10408000;
      30995: inst = 32'hc4044d6;
      30996: inst = 32'h8220000;
      30997: inst = 32'h10408000;
      30998: inst = 32'hc4044d7;
      30999: inst = 32'h8220000;
      31000: inst = 32'h10408000;
      31001: inst = 32'hc4044d8;
      31002: inst = 32'h8220000;
      31003: inst = 32'h10408000;
      31004: inst = 32'hc4044d9;
      31005: inst = 32'h8220000;
      31006: inst = 32'h10408000;
      31007: inst = 32'hc4044da;
      31008: inst = 32'h8220000;
      31009: inst = 32'h10408000;
      31010: inst = 32'hc4044db;
      31011: inst = 32'h8220000;
      31012: inst = 32'h10408000;
      31013: inst = 32'hc4044dc;
      31014: inst = 32'h8220000;
      31015: inst = 32'h10408000;
      31016: inst = 32'hc4044dd;
      31017: inst = 32'h8220000;
      31018: inst = 32'h10408000;
      31019: inst = 32'hc4044de;
      31020: inst = 32'h8220000;
      31021: inst = 32'h10408000;
      31022: inst = 32'hc4044df;
      31023: inst = 32'h8220000;
      31024: inst = 32'h10408000;
      31025: inst = 32'hc4044e0;
      31026: inst = 32'h8220000;
      31027: inst = 32'h10408000;
      31028: inst = 32'hc4044e1;
      31029: inst = 32'h8220000;
      31030: inst = 32'h10408000;
      31031: inst = 32'hc4044e2;
      31032: inst = 32'h8220000;
      31033: inst = 32'h10408000;
      31034: inst = 32'hc4044e3;
      31035: inst = 32'h8220000;
      31036: inst = 32'h10408000;
      31037: inst = 32'hc4044e4;
      31038: inst = 32'h8220000;
      31039: inst = 32'h10408000;
      31040: inst = 32'hc4044e5;
      31041: inst = 32'h8220000;
      31042: inst = 32'h10408000;
      31043: inst = 32'hc4044e6;
      31044: inst = 32'h8220000;
      31045: inst = 32'h10408000;
      31046: inst = 32'hc4044e7;
      31047: inst = 32'h8220000;
      31048: inst = 32'h10408000;
      31049: inst = 32'hc4044e8;
      31050: inst = 32'h8220000;
      31051: inst = 32'h10408000;
      31052: inst = 32'hc4044e9;
      31053: inst = 32'h8220000;
      31054: inst = 32'h10408000;
      31055: inst = 32'hc4044ea;
      31056: inst = 32'h8220000;
      31057: inst = 32'h10408000;
      31058: inst = 32'hc4044eb;
      31059: inst = 32'h8220000;
      31060: inst = 32'h10408000;
      31061: inst = 32'hc4044ec;
      31062: inst = 32'h8220000;
      31063: inst = 32'h10408000;
      31064: inst = 32'hc4044ed;
      31065: inst = 32'h8220000;
      31066: inst = 32'h10408000;
      31067: inst = 32'hc4044ee;
      31068: inst = 32'h8220000;
      31069: inst = 32'h10408000;
      31070: inst = 32'hc4044ef;
      31071: inst = 32'h8220000;
      31072: inst = 32'h10408000;
      31073: inst = 32'hc4044f0;
      31074: inst = 32'h8220000;
      31075: inst = 32'h10408000;
      31076: inst = 32'hc4044f1;
      31077: inst = 32'h8220000;
      31078: inst = 32'h10408000;
      31079: inst = 32'hc4044f2;
      31080: inst = 32'h8220000;
      31081: inst = 32'h10408000;
      31082: inst = 32'hc4044f3;
      31083: inst = 32'h8220000;
      31084: inst = 32'h10408000;
      31085: inst = 32'hc4044f4;
      31086: inst = 32'h8220000;
      31087: inst = 32'h10408000;
      31088: inst = 32'hc4044f5;
      31089: inst = 32'h8220000;
      31090: inst = 32'h10408000;
      31091: inst = 32'hc4044f6;
      31092: inst = 32'h8220000;
      31093: inst = 32'h10408000;
      31094: inst = 32'hc4044f7;
      31095: inst = 32'h8220000;
      31096: inst = 32'h10408000;
      31097: inst = 32'hc4044f8;
      31098: inst = 32'h8220000;
      31099: inst = 32'h10408000;
      31100: inst = 32'hc4044f9;
      31101: inst = 32'h8220000;
      31102: inst = 32'h10408000;
      31103: inst = 32'hc4044fa;
      31104: inst = 32'h8220000;
      31105: inst = 32'h10408000;
      31106: inst = 32'hc4044fb;
      31107: inst = 32'h8220000;
      31108: inst = 32'h10408000;
      31109: inst = 32'hc4044fc;
      31110: inst = 32'h8220000;
      31111: inst = 32'h10408000;
      31112: inst = 32'hc4044fd;
      31113: inst = 32'h8220000;
      31114: inst = 32'h10408000;
      31115: inst = 32'hc4044fe;
      31116: inst = 32'h8220000;
      31117: inst = 32'h10408000;
      31118: inst = 32'hc4044ff;
      31119: inst = 32'h8220000;
      31120: inst = 32'h10408000;
      31121: inst = 32'hc404500;
      31122: inst = 32'h8220000;
      31123: inst = 32'h10408000;
      31124: inst = 32'hc404501;
      31125: inst = 32'h8220000;
      31126: inst = 32'h10408000;
      31127: inst = 32'hc404502;
      31128: inst = 32'h8220000;
      31129: inst = 32'h10408000;
      31130: inst = 32'hc404503;
      31131: inst = 32'h8220000;
      31132: inst = 32'h10408000;
      31133: inst = 32'hc404504;
      31134: inst = 32'h8220000;
      31135: inst = 32'h10408000;
      31136: inst = 32'hc404505;
      31137: inst = 32'h8220000;
      31138: inst = 32'h10408000;
      31139: inst = 32'hc404506;
      31140: inst = 32'h8220000;
      31141: inst = 32'h10408000;
      31142: inst = 32'hc404507;
      31143: inst = 32'h8220000;
      31144: inst = 32'h10408000;
      31145: inst = 32'hc404508;
      31146: inst = 32'h8220000;
      31147: inst = 32'h10408000;
      31148: inst = 32'hc404509;
      31149: inst = 32'h8220000;
      31150: inst = 32'h10408000;
      31151: inst = 32'hc40450a;
      31152: inst = 32'h8220000;
      31153: inst = 32'h10408000;
      31154: inst = 32'hc40450b;
      31155: inst = 32'h8220000;
      31156: inst = 32'h10408000;
      31157: inst = 32'hc40450f;
      31158: inst = 32'h8220000;
      31159: inst = 32'h10408000;
      31160: inst = 32'hc404512;
      31161: inst = 32'h8220000;
      31162: inst = 32'h10408000;
      31163: inst = 32'hc404513;
      31164: inst = 32'h8220000;
      31165: inst = 32'h10408000;
      31166: inst = 32'hc404523;
      31167: inst = 32'h8220000;
      31168: inst = 32'h10408000;
      31169: inst = 32'hc404524;
      31170: inst = 32'h8220000;
      31171: inst = 32'h10408000;
      31172: inst = 32'hc404525;
      31173: inst = 32'h8220000;
      31174: inst = 32'h10408000;
      31175: inst = 32'hc404526;
      31176: inst = 32'h8220000;
      31177: inst = 32'h10408000;
      31178: inst = 32'hc404527;
      31179: inst = 32'h8220000;
      31180: inst = 32'h10408000;
      31181: inst = 32'hc404528;
      31182: inst = 32'h8220000;
      31183: inst = 32'h10408000;
      31184: inst = 32'hc404529;
      31185: inst = 32'h8220000;
      31186: inst = 32'h10408000;
      31187: inst = 32'hc40452a;
      31188: inst = 32'h8220000;
      31189: inst = 32'h10408000;
      31190: inst = 32'hc40452b;
      31191: inst = 32'h8220000;
      31192: inst = 32'h10408000;
      31193: inst = 32'hc40452c;
      31194: inst = 32'h8220000;
      31195: inst = 32'h10408000;
      31196: inst = 32'hc40452d;
      31197: inst = 32'h8220000;
      31198: inst = 32'h10408000;
      31199: inst = 32'hc40452e;
      31200: inst = 32'h8220000;
      31201: inst = 32'h10408000;
      31202: inst = 32'hc40452f;
      31203: inst = 32'h8220000;
      31204: inst = 32'h10408000;
      31205: inst = 32'hc404530;
      31206: inst = 32'h8220000;
      31207: inst = 32'h10408000;
      31208: inst = 32'hc404531;
      31209: inst = 32'h8220000;
      31210: inst = 32'h10408000;
      31211: inst = 32'hc404532;
      31212: inst = 32'h8220000;
      31213: inst = 32'h10408000;
      31214: inst = 32'hc404533;
      31215: inst = 32'h8220000;
      31216: inst = 32'h10408000;
      31217: inst = 32'hc404534;
      31218: inst = 32'h8220000;
      31219: inst = 32'h10408000;
      31220: inst = 32'hc404535;
      31221: inst = 32'h8220000;
      31222: inst = 32'h10408000;
      31223: inst = 32'hc404536;
      31224: inst = 32'h8220000;
      31225: inst = 32'h10408000;
      31226: inst = 32'hc404537;
      31227: inst = 32'h8220000;
      31228: inst = 32'h10408000;
      31229: inst = 32'hc404538;
      31230: inst = 32'h8220000;
      31231: inst = 32'h10408000;
      31232: inst = 32'hc404539;
      31233: inst = 32'h8220000;
      31234: inst = 32'h10408000;
      31235: inst = 32'hc40453a;
      31236: inst = 32'h8220000;
      31237: inst = 32'h10408000;
      31238: inst = 32'hc40453b;
      31239: inst = 32'h8220000;
      31240: inst = 32'h10408000;
      31241: inst = 32'hc40453c;
      31242: inst = 32'h8220000;
      31243: inst = 32'h10408000;
      31244: inst = 32'hc40453d;
      31245: inst = 32'h8220000;
      31246: inst = 32'h10408000;
      31247: inst = 32'hc40453e;
      31248: inst = 32'h8220000;
      31249: inst = 32'h10408000;
      31250: inst = 32'hc40453f;
      31251: inst = 32'h8220000;
      31252: inst = 32'h10408000;
      31253: inst = 32'hc404540;
      31254: inst = 32'h8220000;
      31255: inst = 32'h10408000;
      31256: inst = 32'hc404541;
      31257: inst = 32'h8220000;
      31258: inst = 32'h10408000;
      31259: inst = 32'hc404542;
      31260: inst = 32'h8220000;
      31261: inst = 32'h10408000;
      31262: inst = 32'hc404543;
      31263: inst = 32'h8220000;
      31264: inst = 32'h10408000;
      31265: inst = 32'hc404544;
      31266: inst = 32'h8220000;
      31267: inst = 32'h10408000;
      31268: inst = 32'hc404545;
      31269: inst = 32'h8220000;
      31270: inst = 32'h10408000;
      31271: inst = 32'hc404546;
      31272: inst = 32'h8220000;
      31273: inst = 32'h10408000;
      31274: inst = 32'hc404547;
      31275: inst = 32'h8220000;
      31276: inst = 32'h10408000;
      31277: inst = 32'hc404548;
      31278: inst = 32'h8220000;
      31279: inst = 32'h10408000;
      31280: inst = 32'hc404549;
      31281: inst = 32'h8220000;
      31282: inst = 32'h10408000;
      31283: inst = 32'hc40454a;
      31284: inst = 32'h8220000;
      31285: inst = 32'h10408000;
      31286: inst = 32'hc40454b;
      31287: inst = 32'h8220000;
      31288: inst = 32'h10408000;
      31289: inst = 32'hc40454c;
      31290: inst = 32'h8220000;
      31291: inst = 32'h10408000;
      31292: inst = 32'hc40454d;
      31293: inst = 32'h8220000;
      31294: inst = 32'h10408000;
      31295: inst = 32'hc40454e;
      31296: inst = 32'h8220000;
      31297: inst = 32'h10408000;
      31298: inst = 32'hc40454f;
      31299: inst = 32'h8220000;
      31300: inst = 32'h10408000;
      31301: inst = 32'hc404550;
      31302: inst = 32'h8220000;
      31303: inst = 32'h10408000;
      31304: inst = 32'hc404551;
      31305: inst = 32'h8220000;
      31306: inst = 32'h10408000;
      31307: inst = 32'hc404552;
      31308: inst = 32'h8220000;
      31309: inst = 32'h10408000;
      31310: inst = 32'hc404553;
      31311: inst = 32'h8220000;
      31312: inst = 32'h10408000;
      31313: inst = 32'hc404554;
      31314: inst = 32'h8220000;
      31315: inst = 32'h10408000;
      31316: inst = 32'hc404555;
      31317: inst = 32'h8220000;
      31318: inst = 32'h10408000;
      31319: inst = 32'hc404556;
      31320: inst = 32'h8220000;
      31321: inst = 32'h10408000;
      31322: inst = 32'hc404557;
      31323: inst = 32'h8220000;
      31324: inst = 32'h10408000;
      31325: inst = 32'hc404558;
      31326: inst = 32'h8220000;
      31327: inst = 32'h10408000;
      31328: inst = 32'hc404559;
      31329: inst = 32'h8220000;
      31330: inst = 32'h10408000;
      31331: inst = 32'hc40455a;
      31332: inst = 32'h8220000;
      31333: inst = 32'h10408000;
      31334: inst = 32'hc40455b;
      31335: inst = 32'h8220000;
      31336: inst = 32'h10408000;
      31337: inst = 32'hc40455c;
      31338: inst = 32'h8220000;
      31339: inst = 32'h10408000;
      31340: inst = 32'hc40455d;
      31341: inst = 32'h8220000;
      31342: inst = 32'h10408000;
      31343: inst = 32'hc40455e;
      31344: inst = 32'h8220000;
      31345: inst = 32'h10408000;
      31346: inst = 32'hc40455f;
      31347: inst = 32'h8220000;
      31348: inst = 32'h10408000;
      31349: inst = 32'hc404560;
      31350: inst = 32'h8220000;
      31351: inst = 32'h10408000;
      31352: inst = 32'hc404561;
      31353: inst = 32'h8220000;
      31354: inst = 32'h10408000;
      31355: inst = 32'hc404562;
      31356: inst = 32'h8220000;
      31357: inst = 32'h10408000;
      31358: inst = 32'hc404563;
      31359: inst = 32'h8220000;
      31360: inst = 32'h10408000;
      31361: inst = 32'hc404564;
      31362: inst = 32'h8220000;
      31363: inst = 32'h10408000;
      31364: inst = 32'hc404565;
      31365: inst = 32'h8220000;
      31366: inst = 32'h10408000;
      31367: inst = 32'hc404566;
      31368: inst = 32'h8220000;
      31369: inst = 32'h10408000;
      31370: inst = 32'hc404567;
      31371: inst = 32'h8220000;
      31372: inst = 32'h10408000;
      31373: inst = 32'hc404568;
      31374: inst = 32'h8220000;
      31375: inst = 32'h10408000;
      31376: inst = 32'hc404569;
      31377: inst = 32'h8220000;
      31378: inst = 32'h10408000;
      31379: inst = 32'hc40456a;
      31380: inst = 32'h8220000;
      31381: inst = 32'h10408000;
      31382: inst = 32'hc40456b;
      31383: inst = 32'h8220000;
      31384: inst = 32'h10408000;
      31385: inst = 32'hc40456f;
      31386: inst = 32'h8220000;
      31387: inst = 32'h10408000;
      31388: inst = 32'hc40457a;
      31389: inst = 32'h8220000;
      31390: inst = 32'h10408000;
      31391: inst = 32'hc40457b;
      31392: inst = 32'h8220000;
      31393: inst = 32'h10408000;
      31394: inst = 32'hc40457c;
      31395: inst = 32'h8220000;
      31396: inst = 32'h10408000;
      31397: inst = 32'hc404583;
      31398: inst = 32'h8220000;
      31399: inst = 32'h10408000;
      31400: inst = 32'hc404584;
      31401: inst = 32'h8220000;
      31402: inst = 32'h10408000;
      31403: inst = 32'hc404585;
      31404: inst = 32'h8220000;
      31405: inst = 32'h10408000;
      31406: inst = 32'hc404586;
      31407: inst = 32'h8220000;
      31408: inst = 32'h10408000;
      31409: inst = 32'hc404587;
      31410: inst = 32'h8220000;
      31411: inst = 32'h10408000;
      31412: inst = 32'hc404588;
      31413: inst = 32'h8220000;
      31414: inst = 32'h10408000;
      31415: inst = 32'hc404589;
      31416: inst = 32'h8220000;
      31417: inst = 32'h10408000;
      31418: inst = 32'hc40458a;
      31419: inst = 32'h8220000;
      31420: inst = 32'h10408000;
      31421: inst = 32'hc40458b;
      31422: inst = 32'h8220000;
      31423: inst = 32'h10408000;
      31424: inst = 32'hc40458c;
      31425: inst = 32'h8220000;
      31426: inst = 32'h10408000;
      31427: inst = 32'hc40458d;
      31428: inst = 32'h8220000;
      31429: inst = 32'h10408000;
      31430: inst = 32'hc40458e;
      31431: inst = 32'h8220000;
      31432: inst = 32'h10408000;
      31433: inst = 32'hc40458f;
      31434: inst = 32'h8220000;
      31435: inst = 32'h10408000;
      31436: inst = 32'hc404590;
      31437: inst = 32'h8220000;
      31438: inst = 32'h10408000;
      31439: inst = 32'hc404591;
      31440: inst = 32'h8220000;
      31441: inst = 32'h10408000;
      31442: inst = 32'hc404592;
      31443: inst = 32'h8220000;
      31444: inst = 32'h10408000;
      31445: inst = 32'hc404593;
      31446: inst = 32'h8220000;
      31447: inst = 32'h10408000;
      31448: inst = 32'hc404594;
      31449: inst = 32'h8220000;
      31450: inst = 32'h10408000;
      31451: inst = 32'hc404595;
      31452: inst = 32'h8220000;
      31453: inst = 32'h10408000;
      31454: inst = 32'hc404596;
      31455: inst = 32'h8220000;
      31456: inst = 32'h10408000;
      31457: inst = 32'hc404597;
      31458: inst = 32'h8220000;
      31459: inst = 32'h10408000;
      31460: inst = 32'hc404598;
      31461: inst = 32'h8220000;
      31462: inst = 32'h10408000;
      31463: inst = 32'hc404599;
      31464: inst = 32'h8220000;
      31465: inst = 32'h10408000;
      31466: inst = 32'hc40459a;
      31467: inst = 32'h8220000;
      31468: inst = 32'h10408000;
      31469: inst = 32'hc40459b;
      31470: inst = 32'h8220000;
      31471: inst = 32'h10408000;
      31472: inst = 32'hc40459c;
      31473: inst = 32'h8220000;
      31474: inst = 32'h10408000;
      31475: inst = 32'hc40459d;
      31476: inst = 32'h8220000;
      31477: inst = 32'h10408000;
      31478: inst = 32'hc40459e;
      31479: inst = 32'h8220000;
      31480: inst = 32'h10408000;
      31481: inst = 32'hc40459f;
      31482: inst = 32'h8220000;
      31483: inst = 32'h10408000;
      31484: inst = 32'hc4045a0;
      31485: inst = 32'h8220000;
      31486: inst = 32'h10408000;
      31487: inst = 32'hc4045a1;
      31488: inst = 32'h8220000;
      31489: inst = 32'h10408000;
      31490: inst = 32'hc4045a2;
      31491: inst = 32'h8220000;
      31492: inst = 32'h10408000;
      31493: inst = 32'hc4045a3;
      31494: inst = 32'h8220000;
      31495: inst = 32'h10408000;
      31496: inst = 32'hc4045a4;
      31497: inst = 32'h8220000;
      31498: inst = 32'h10408000;
      31499: inst = 32'hc4045a5;
      31500: inst = 32'h8220000;
      31501: inst = 32'h10408000;
      31502: inst = 32'hc4045a6;
      31503: inst = 32'h8220000;
      31504: inst = 32'h10408000;
      31505: inst = 32'hc4045a7;
      31506: inst = 32'h8220000;
      31507: inst = 32'h10408000;
      31508: inst = 32'hc4045a8;
      31509: inst = 32'h8220000;
      31510: inst = 32'h10408000;
      31511: inst = 32'hc4045a9;
      31512: inst = 32'h8220000;
      31513: inst = 32'h10408000;
      31514: inst = 32'hc4045aa;
      31515: inst = 32'h8220000;
      31516: inst = 32'h10408000;
      31517: inst = 32'hc4045ab;
      31518: inst = 32'h8220000;
      31519: inst = 32'h10408000;
      31520: inst = 32'hc4045ac;
      31521: inst = 32'h8220000;
      31522: inst = 32'h10408000;
      31523: inst = 32'hc4045ad;
      31524: inst = 32'h8220000;
      31525: inst = 32'h10408000;
      31526: inst = 32'hc4045ae;
      31527: inst = 32'h8220000;
      31528: inst = 32'h10408000;
      31529: inst = 32'hc4045af;
      31530: inst = 32'h8220000;
      31531: inst = 32'h10408000;
      31532: inst = 32'hc4045b0;
      31533: inst = 32'h8220000;
      31534: inst = 32'h10408000;
      31535: inst = 32'hc4045b1;
      31536: inst = 32'h8220000;
      31537: inst = 32'h10408000;
      31538: inst = 32'hc4045b2;
      31539: inst = 32'h8220000;
      31540: inst = 32'h10408000;
      31541: inst = 32'hc4045b3;
      31542: inst = 32'h8220000;
      31543: inst = 32'h10408000;
      31544: inst = 32'hc4045b4;
      31545: inst = 32'h8220000;
      31546: inst = 32'h10408000;
      31547: inst = 32'hc4045b5;
      31548: inst = 32'h8220000;
      31549: inst = 32'h10408000;
      31550: inst = 32'hc4045b6;
      31551: inst = 32'h8220000;
      31552: inst = 32'h10408000;
      31553: inst = 32'hc4045b7;
      31554: inst = 32'h8220000;
      31555: inst = 32'h10408000;
      31556: inst = 32'hc4045b8;
      31557: inst = 32'h8220000;
      31558: inst = 32'h10408000;
      31559: inst = 32'hc4045b9;
      31560: inst = 32'h8220000;
      31561: inst = 32'h10408000;
      31562: inst = 32'hc4045ba;
      31563: inst = 32'h8220000;
      31564: inst = 32'h10408000;
      31565: inst = 32'hc4045bb;
      31566: inst = 32'h8220000;
      31567: inst = 32'h10408000;
      31568: inst = 32'hc4045bc;
      31569: inst = 32'h8220000;
      31570: inst = 32'h10408000;
      31571: inst = 32'hc4045bd;
      31572: inst = 32'h8220000;
      31573: inst = 32'h10408000;
      31574: inst = 32'hc4045be;
      31575: inst = 32'h8220000;
      31576: inst = 32'h10408000;
      31577: inst = 32'hc4045bf;
      31578: inst = 32'h8220000;
      31579: inst = 32'h10408000;
      31580: inst = 32'hc4045c0;
      31581: inst = 32'h8220000;
      31582: inst = 32'h10408000;
      31583: inst = 32'hc4045c1;
      31584: inst = 32'h8220000;
      31585: inst = 32'h10408000;
      31586: inst = 32'hc4045c2;
      31587: inst = 32'h8220000;
      31588: inst = 32'h10408000;
      31589: inst = 32'hc4045c3;
      31590: inst = 32'h8220000;
      31591: inst = 32'h10408000;
      31592: inst = 32'hc4045c4;
      31593: inst = 32'h8220000;
      31594: inst = 32'h10408000;
      31595: inst = 32'hc4045c5;
      31596: inst = 32'h8220000;
      31597: inst = 32'h10408000;
      31598: inst = 32'hc4045c6;
      31599: inst = 32'h8220000;
      31600: inst = 32'h10408000;
      31601: inst = 32'hc4045c7;
      31602: inst = 32'h8220000;
      31603: inst = 32'h10408000;
      31604: inst = 32'hc4045c8;
      31605: inst = 32'h8220000;
      31606: inst = 32'h10408000;
      31607: inst = 32'hc4045c9;
      31608: inst = 32'h8220000;
      31609: inst = 32'h10408000;
      31610: inst = 32'hc4045ca;
      31611: inst = 32'h8220000;
      31612: inst = 32'h10408000;
      31613: inst = 32'hc4045cb;
      31614: inst = 32'h8220000;
      31615: inst = 32'h10408000;
      31616: inst = 32'hc4045cf;
      31617: inst = 32'h8220000;
      31618: inst = 32'h10408000;
      31619: inst = 32'hc4045d0;
      31620: inst = 32'h8220000;
      31621: inst = 32'h10408000;
      31622: inst = 32'hc4045d4;
      31623: inst = 32'h8220000;
      31624: inst = 32'h10408000;
      31625: inst = 32'hc4045d5;
      31626: inst = 32'h8220000;
      31627: inst = 32'h10408000;
      31628: inst = 32'hc4045d6;
      31629: inst = 32'h8220000;
      31630: inst = 32'h10408000;
      31631: inst = 32'hc4045d7;
      31632: inst = 32'h8220000;
      31633: inst = 32'h10408000;
      31634: inst = 32'hc4045da;
      31635: inst = 32'h8220000;
      31636: inst = 32'h10408000;
      31637: inst = 32'hc4045db;
      31638: inst = 32'h8220000;
      31639: inst = 32'h10408000;
      31640: inst = 32'hc4045e3;
      31641: inst = 32'h8220000;
      31642: inst = 32'h10408000;
      31643: inst = 32'hc4045e4;
      31644: inst = 32'h8220000;
      31645: inst = 32'h10408000;
      31646: inst = 32'hc4045e5;
      31647: inst = 32'h8220000;
      31648: inst = 32'h10408000;
      31649: inst = 32'hc4045e6;
      31650: inst = 32'h8220000;
      31651: inst = 32'h10408000;
      31652: inst = 32'hc4045e7;
      31653: inst = 32'h8220000;
      31654: inst = 32'h10408000;
      31655: inst = 32'hc4045e8;
      31656: inst = 32'h8220000;
      31657: inst = 32'h10408000;
      31658: inst = 32'hc4045e9;
      31659: inst = 32'h8220000;
      31660: inst = 32'h10408000;
      31661: inst = 32'hc4045ea;
      31662: inst = 32'h8220000;
      31663: inst = 32'h10408000;
      31664: inst = 32'hc4045eb;
      31665: inst = 32'h8220000;
      31666: inst = 32'h10408000;
      31667: inst = 32'hc4045ec;
      31668: inst = 32'h8220000;
      31669: inst = 32'h10408000;
      31670: inst = 32'hc4045ed;
      31671: inst = 32'h8220000;
      31672: inst = 32'h10408000;
      31673: inst = 32'hc4045ee;
      31674: inst = 32'h8220000;
      31675: inst = 32'h10408000;
      31676: inst = 32'hc4045ef;
      31677: inst = 32'h8220000;
      31678: inst = 32'h10408000;
      31679: inst = 32'hc4045f0;
      31680: inst = 32'h8220000;
      31681: inst = 32'h10408000;
      31682: inst = 32'hc4045f1;
      31683: inst = 32'h8220000;
      31684: inst = 32'h10408000;
      31685: inst = 32'hc4045f2;
      31686: inst = 32'h8220000;
      31687: inst = 32'h10408000;
      31688: inst = 32'hc4045f3;
      31689: inst = 32'h8220000;
      31690: inst = 32'h10408000;
      31691: inst = 32'hc4045f4;
      31692: inst = 32'h8220000;
      31693: inst = 32'h10408000;
      31694: inst = 32'hc4045f5;
      31695: inst = 32'h8220000;
      31696: inst = 32'h10408000;
      31697: inst = 32'hc4045f6;
      31698: inst = 32'h8220000;
      31699: inst = 32'h10408000;
      31700: inst = 32'hc4045f7;
      31701: inst = 32'h8220000;
      31702: inst = 32'h10408000;
      31703: inst = 32'hc4045f8;
      31704: inst = 32'h8220000;
      31705: inst = 32'h10408000;
      31706: inst = 32'hc4045f9;
      31707: inst = 32'h8220000;
      31708: inst = 32'h10408000;
      31709: inst = 32'hc4045fa;
      31710: inst = 32'h8220000;
      31711: inst = 32'h10408000;
      31712: inst = 32'hc4045fb;
      31713: inst = 32'h8220000;
      31714: inst = 32'h10408000;
      31715: inst = 32'hc4045fc;
      31716: inst = 32'h8220000;
      31717: inst = 32'h10408000;
      31718: inst = 32'hc4045fd;
      31719: inst = 32'h8220000;
      31720: inst = 32'h10408000;
      31721: inst = 32'hc4045fe;
      31722: inst = 32'h8220000;
      31723: inst = 32'h10408000;
      31724: inst = 32'hc4045ff;
      31725: inst = 32'h8220000;
      31726: inst = 32'h10408000;
      31727: inst = 32'hc404600;
      31728: inst = 32'h8220000;
      31729: inst = 32'h10408000;
      31730: inst = 32'hc404601;
      31731: inst = 32'h8220000;
      31732: inst = 32'h10408000;
      31733: inst = 32'hc404602;
      31734: inst = 32'h8220000;
      31735: inst = 32'h10408000;
      31736: inst = 32'hc404603;
      31737: inst = 32'h8220000;
      31738: inst = 32'h10408000;
      31739: inst = 32'hc404604;
      31740: inst = 32'h8220000;
      31741: inst = 32'h10408000;
      31742: inst = 32'hc404605;
      31743: inst = 32'h8220000;
      31744: inst = 32'h10408000;
      31745: inst = 32'hc404606;
      31746: inst = 32'h8220000;
      31747: inst = 32'h10408000;
      31748: inst = 32'hc404607;
      31749: inst = 32'h8220000;
      31750: inst = 32'h10408000;
      31751: inst = 32'hc404608;
      31752: inst = 32'h8220000;
      31753: inst = 32'h10408000;
      31754: inst = 32'hc404609;
      31755: inst = 32'h8220000;
      31756: inst = 32'h10408000;
      31757: inst = 32'hc40460a;
      31758: inst = 32'h8220000;
      31759: inst = 32'h10408000;
      31760: inst = 32'hc40460b;
      31761: inst = 32'h8220000;
      31762: inst = 32'h10408000;
      31763: inst = 32'hc40460c;
      31764: inst = 32'h8220000;
      31765: inst = 32'h10408000;
      31766: inst = 32'hc40460d;
      31767: inst = 32'h8220000;
      31768: inst = 32'h10408000;
      31769: inst = 32'hc40460e;
      31770: inst = 32'h8220000;
      31771: inst = 32'h10408000;
      31772: inst = 32'hc40460f;
      31773: inst = 32'h8220000;
      31774: inst = 32'h10408000;
      31775: inst = 32'hc404610;
      31776: inst = 32'h8220000;
      31777: inst = 32'h10408000;
      31778: inst = 32'hc404611;
      31779: inst = 32'h8220000;
      31780: inst = 32'h10408000;
      31781: inst = 32'hc404612;
      31782: inst = 32'h8220000;
      31783: inst = 32'h10408000;
      31784: inst = 32'hc404613;
      31785: inst = 32'h8220000;
      31786: inst = 32'h10408000;
      31787: inst = 32'hc404614;
      31788: inst = 32'h8220000;
      31789: inst = 32'h10408000;
      31790: inst = 32'hc404615;
      31791: inst = 32'h8220000;
      31792: inst = 32'h10408000;
      31793: inst = 32'hc404616;
      31794: inst = 32'h8220000;
      31795: inst = 32'h10408000;
      31796: inst = 32'hc404617;
      31797: inst = 32'h8220000;
      31798: inst = 32'h10408000;
      31799: inst = 32'hc404618;
      31800: inst = 32'h8220000;
      31801: inst = 32'h10408000;
      31802: inst = 32'hc404619;
      31803: inst = 32'h8220000;
      31804: inst = 32'h10408000;
      31805: inst = 32'hc40461a;
      31806: inst = 32'h8220000;
      31807: inst = 32'h10408000;
      31808: inst = 32'hc40461b;
      31809: inst = 32'h8220000;
      31810: inst = 32'h10408000;
      31811: inst = 32'hc40461c;
      31812: inst = 32'h8220000;
      31813: inst = 32'h10408000;
      31814: inst = 32'hc40461d;
      31815: inst = 32'h8220000;
      31816: inst = 32'h10408000;
      31817: inst = 32'hc40461e;
      31818: inst = 32'h8220000;
      31819: inst = 32'h10408000;
      31820: inst = 32'hc40461f;
      31821: inst = 32'h8220000;
      31822: inst = 32'h10408000;
      31823: inst = 32'hc404620;
      31824: inst = 32'h8220000;
      31825: inst = 32'h10408000;
      31826: inst = 32'hc404621;
      31827: inst = 32'h8220000;
      31828: inst = 32'h10408000;
      31829: inst = 32'hc404622;
      31830: inst = 32'h8220000;
      31831: inst = 32'h10408000;
      31832: inst = 32'hc404623;
      31833: inst = 32'h8220000;
      31834: inst = 32'h10408000;
      31835: inst = 32'hc404624;
      31836: inst = 32'h8220000;
      31837: inst = 32'h10408000;
      31838: inst = 32'hc404625;
      31839: inst = 32'h8220000;
      31840: inst = 32'h10408000;
      31841: inst = 32'hc404626;
      31842: inst = 32'h8220000;
      31843: inst = 32'h10408000;
      31844: inst = 32'hc404627;
      31845: inst = 32'h8220000;
      31846: inst = 32'h10408000;
      31847: inst = 32'hc404628;
      31848: inst = 32'h8220000;
      31849: inst = 32'h10408000;
      31850: inst = 32'hc404629;
      31851: inst = 32'h8220000;
      31852: inst = 32'h10408000;
      31853: inst = 32'hc40462a;
      31854: inst = 32'h8220000;
      31855: inst = 32'h10408000;
      31856: inst = 32'hc40462b;
      31857: inst = 32'h8220000;
      31858: inst = 32'h10408000;
      31859: inst = 32'hc40462f;
      31860: inst = 32'h8220000;
      31861: inst = 32'h10408000;
      31862: inst = 32'hc404630;
      31863: inst = 32'h8220000;
      31864: inst = 32'h10408000;
      31865: inst = 32'hc404631;
      31866: inst = 32'h8220000;
      31867: inst = 32'h10408000;
      31868: inst = 32'hc404632;
      31869: inst = 32'h8220000;
      31870: inst = 32'h10408000;
      31871: inst = 32'hc404633;
      31872: inst = 32'h8220000;
      31873: inst = 32'h10408000;
      31874: inst = 32'hc404634;
      31875: inst = 32'h8220000;
      31876: inst = 32'h10408000;
      31877: inst = 32'hc404635;
      31878: inst = 32'h8220000;
      31879: inst = 32'h10408000;
      31880: inst = 32'hc404636;
      31881: inst = 32'h8220000;
      31882: inst = 32'h10408000;
      31883: inst = 32'hc404637;
      31884: inst = 32'h8220000;
      31885: inst = 32'h10408000;
      31886: inst = 32'hc404638;
      31887: inst = 32'h8220000;
      31888: inst = 32'h10408000;
      31889: inst = 32'hc404639;
      31890: inst = 32'h8220000;
      31891: inst = 32'h10408000;
      31892: inst = 32'hc40463a;
      31893: inst = 32'h8220000;
      31894: inst = 32'h10408000;
      31895: inst = 32'hc40463b;
      31896: inst = 32'h8220000;
      31897: inst = 32'h10408000;
      31898: inst = 32'hc40463c;
      31899: inst = 32'h8220000;
      31900: inst = 32'h10408000;
      31901: inst = 32'hc404643;
      31902: inst = 32'h8220000;
      31903: inst = 32'h10408000;
      31904: inst = 32'hc404644;
      31905: inst = 32'h8220000;
      31906: inst = 32'h10408000;
      31907: inst = 32'hc404645;
      31908: inst = 32'h8220000;
      31909: inst = 32'h10408000;
      31910: inst = 32'hc404646;
      31911: inst = 32'h8220000;
      31912: inst = 32'h10408000;
      31913: inst = 32'hc404647;
      31914: inst = 32'h8220000;
      31915: inst = 32'h10408000;
      31916: inst = 32'hc404648;
      31917: inst = 32'h8220000;
      31918: inst = 32'h10408000;
      31919: inst = 32'hc404649;
      31920: inst = 32'h8220000;
      31921: inst = 32'h10408000;
      31922: inst = 32'hc40464a;
      31923: inst = 32'h8220000;
      31924: inst = 32'h10408000;
      31925: inst = 32'hc40464b;
      31926: inst = 32'h8220000;
      31927: inst = 32'h10408000;
      31928: inst = 32'hc40464c;
      31929: inst = 32'h8220000;
      31930: inst = 32'h10408000;
      31931: inst = 32'hc40464d;
      31932: inst = 32'h8220000;
      31933: inst = 32'h10408000;
      31934: inst = 32'hc40467a;
      31935: inst = 32'h8220000;
      31936: inst = 32'h10408000;
      31937: inst = 32'hc40467b;
      31938: inst = 32'h8220000;
      31939: inst = 32'h10408000;
      31940: inst = 32'hc40467c;
      31941: inst = 32'h8220000;
      31942: inst = 32'h10408000;
      31943: inst = 32'hc40467d;
      31944: inst = 32'h8220000;
      31945: inst = 32'h10408000;
      31946: inst = 32'hc40467e;
      31947: inst = 32'h8220000;
      31948: inst = 32'h10408000;
      31949: inst = 32'hc40467f;
      31950: inst = 32'h8220000;
      31951: inst = 32'h10408000;
      31952: inst = 32'hc404680;
      31953: inst = 32'h8220000;
      31954: inst = 32'h10408000;
      31955: inst = 32'hc404681;
      31956: inst = 32'h8220000;
      31957: inst = 32'h10408000;
      31958: inst = 32'hc404682;
      31959: inst = 32'h8220000;
      31960: inst = 32'h10408000;
      31961: inst = 32'hc404683;
      31962: inst = 32'h8220000;
      31963: inst = 32'h10408000;
      31964: inst = 32'hc404684;
      31965: inst = 32'h8220000;
      31966: inst = 32'h10408000;
      31967: inst = 32'hc404685;
      31968: inst = 32'h8220000;
      31969: inst = 32'h10408000;
      31970: inst = 32'hc404686;
      31971: inst = 32'h8220000;
      31972: inst = 32'h10408000;
      31973: inst = 32'hc404687;
      31974: inst = 32'h8220000;
      31975: inst = 32'h10408000;
      31976: inst = 32'hc404688;
      31977: inst = 32'h8220000;
      31978: inst = 32'h10408000;
      31979: inst = 32'hc404689;
      31980: inst = 32'h8220000;
      31981: inst = 32'h10408000;
      31982: inst = 32'hc40468a;
      31983: inst = 32'h8220000;
      31984: inst = 32'h10408000;
      31985: inst = 32'hc40468b;
      31986: inst = 32'h8220000;
      31987: inst = 32'h10408000;
      31988: inst = 32'hc40468f;
      31989: inst = 32'h8220000;
      31990: inst = 32'h10408000;
      31991: inst = 32'hc404690;
      31992: inst = 32'h8220000;
      31993: inst = 32'h10408000;
      31994: inst = 32'hc404691;
      31995: inst = 32'h8220000;
      31996: inst = 32'h10408000;
      31997: inst = 32'hc404692;
      31998: inst = 32'h8220000;
      31999: inst = 32'h10408000;
      32000: inst = 32'hc404693;
      32001: inst = 32'h8220000;
      32002: inst = 32'h10408000;
      32003: inst = 32'hc404694;
      32004: inst = 32'h8220000;
      32005: inst = 32'h10408000;
      32006: inst = 32'hc404695;
      32007: inst = 32'h8220000;
      32008: inst = 32'h10408000;
      32009: inst = 32'hc404696;
      32010: inst = 32'h8220000;
      32011: inst = 32'h10408000;
      32012: inst = 32'hc404697;
      32013: inst = 32'h8220000;
      32014: inst = 32'h10408000;
      32015: inst = 32'hc404698;
      32016: inst = 32'h8220000;
      32017: inst = 32'h10408000;
      32018: inst = 32'hc404699;
      32019: inst = 32'h8220000;
      32020: inst = 32'h10408000;
      32021: inst = 32'hc40469a;
      32022: inst = 32'h8220000;
      32023: inst = 32'h10408000;
      32024: inst = 32'hc40469b;
      32025: inst = 32'h8220000;
      32026: inst = 32'h10408000;
      32027: inst = 32'hc40469c;
      32028: inst = 32'h8220000;
      32029: inst = 32'h10408000;
      32030: inst = 32'hc4046a3;
      32031: inst = 32'h8220000;
      32032: inst = 32'h10408000;
      32033: inst = 32'hc4046a4;
      32034: inst = 32'h8220000;
      32035: inst = 32'h10408000;
      32036: inst = 32'hc4046a5;
      32037: inst = 32'h8220000;
      32038: inst = 32'h10408000;
      32039: inst = 32'hc4046a6;
      32040: inst = 32'h8220000;
      32041: inst = 32'h10408000;
      32042: inst = 32'hc4046a7;
      32043: inst = 32'h8220000;
      32044: inst = 32'h10408000;
      32045: inst = 32'hc4046a8;
      32046: inst = 32'h8220000;
      32047: inst = 32'h10408000;
      32048: inst = 32'hc4046a9;
      32049: inst = 32'h8220000;
      32050: inst = 32'h10408000;
      32051: inst = 32'hc4046aa;
      32052: inst = 32'h8220000;
      32053: inst = 32'h10408000;
      32054: inst = 32'hc4046ab;
      32055: inst = 32'h8220000;
      32056: inst = 32'h10408000;
      32057: inst = 32'hc4046ac;
      32058: inst = 32'h8220000;
      32059: inst = 32'h10408000;
      32060: inst = 32'hc4046ad;
      32061: inst = 32'h8220000;
      32062: inst = 32'h10408000;
      32063: inst = 32'hc4046da;
      32064: inst = 32'h8220000;
      32065: inst = 32'h10408000;
      32066: inst = 32'hc4046db;
      32067: inst = 32'h8220000;
      32068: inst = 32'h10408000;
      32069: inst = 32'hc4046dc;
      32070: inst = 32'h8220000;
      32071: inst = 32'h10408000;
      32072: inst = 32'hc4046dd;
      32073: inst = 32'h8220000;
      32074: inst = 32'h10408000;
      32075: inst = 32'hc4046de;
      32076: inst = 32'h8220000;
      32077: inst = 32'h10408000;
      32078: inst = 32'hc4046df;
      32079: inst = 32'h8220000;
      32080: inst = 32'h10408000;
      32081: inst = 32'hc4046e0;
      32082: inst = 32'h8220000;
      32083: inst = 32'h10408000;
      32084: inst = 32'hc4046e1;
      32085: inst = 32'h8220000;
      32086: inst = 32'h10408000;
      32087: inst = 32'hc4046e2;
      32088: inst = 32'h8220000;
      32089: inst = 32'h10408000;
      32090: inst = 32'hc4046e3;
      32091: inst = 32'h8220000;
      32092: inst = 32'h10408000;
      32093: inst = 32'hc4046e4;
      32094: inst = 32'h8220000;
      32095: inst = 32'h10408000;
      32096: inst = 32'hc4046e5;
      32097: inst = 32'h8220000;
      32098: inst = 32'h10408000;
      32099: inst = 32'hc4046e6;
      32100: inst = 32'h8220000;
      32101: inst = 32'h10408000;
      32102: inst = 32'hc4046e7;
      32103: inst = 32'h8220000;
      32104: inst = 32'h10408000;
      32105: inst = 32'hc4046e8;
      32106: inst = 32'h8220000;
      32107: inst = 32'h10408000;
      32108: inst = 32'hc4046e9;
      32109: inst = 32'h8220000;
      32110: inst = 32'h10408000;
      32111: inst = 32'hc4046ea;
      32112: inst = 32'h8220000;
      32113: inst = 32'h10408000;
      32114: inst = 32'hc4046eb;
      32115: inst = 32'h8220000;
      32116: inst = 32'h10408000;
      32117: inst = 32'hc4046ef;
      32118: inst = 32'h8220000;
      32119: inst = 32'h10408000;
      32120: inst = 32'hc4046f0;
      32121: inst = 32'h8220000;
      32122: inst = 32'h10408000;
      32123: inst = 32'hc4046f1;
      32124: inst = 32'h8220000;
      32125: inst = 32'h10408000;
      32126: inst = 32'hc4046f2;
      32127: inst = 32'h8220000;
      32128: inst = 32'h10408000;
      32129: inst = 32'hc4046f3;
      32130: inst = 32'h8220000;
      32131: inst = 32'h10408000;
      32132: inst = 32'hc4046f4;
      32133: inst = 32'h8220000;
      32134: inst = 32'h10408000;
      32135: inst = 32'hc4046f5;
      32136: inst = 32'h8220000;
      32137: inst = 32'h10408000;
      32138: inst = 32'hc4046f6;
      32139: inst = 32'h8220000;
      32140: inst = 32'h10408000;
      32141: inst = 32'hc4046f7;
      32142: inst = 32'h8220000;
      32143: inst = 32'h10408000;
      32144: inst = 32'hc4046f8;
      32145: inst = 32'h8220000;
      32146: inst = 32'h10408000;
      32147: inst = 32'hc4046f9;
      32148: inst = 32'h8220000;
      32149: inst = 32'h10408000;
      32150: inst = 32'hc4046fa;
      32151: inst = 32'h8220000;
      32152: inst = 32'h10408000;
      32153: inst = 32'hc4046fb;
      32154: inst = 32'h8220000;
      32155: inst = 32'h10408000;
      32156: inst = 32'hc4046fc;
      32157: inst = 32'h8220000;
      32158: inst = 32'h10408000;
      32159: inst = 32'hc404703;
      32160: inst = 32'h8220000;
      32161: inst = 32'h10408000;
      32162: inst = 32'hc404704;
      32163: inst = 32'h8220000;
      32164: inst = 32'h10408000;
      32165: inst = 32'hc404705;
      32166: inst = 32'h8220000;
      32167: inst = 32'h10408000;
      32168: inst = 32'hc404706;
      32169: inst = 32'h8220000;
      32170: inst = 32'h10408000;
      32171: inst = 32'hc404707;
      32172: inst = 32'h8220000;
      32173: inst = 32'h10408000;
      32174: inst = 32'hc404708;
      32175: inst = 32'h8220000;
      32176: inst = 32'h10408000;
      32177: inst = 32'hc404709;
      32178: inst = 32'h8220000;
      32179: inst = 32'h10408000;
      32180: inst = 32'hc40470a;
      32181: inst = 32'h8220000;
      32182: inst = 32'h10408000;
      32183: inst = 32'hc40470b;
      32184: inst = 32'h8220000;
      32185: inst = 32'h10408000;
      32186: inst = 32'hc40470c;
      32187: inst = 32'h8220000;
      32188: inst = 32'h10408000;
      32189: inst = 32'hc40470d;
      32190: inst = 32'h8220000;
      32191: inst = 32'h10408000;
      32192: inst = 32'hc40473a;
      32193: inst = 32'h8220000;
      32194: inst = 32'h10408000;
      32195: inst = 32'hc40473b;
      32196: inst = 32'h8220000;
      32197: inst = 32'h10408000;
      32198: inst = 32'hc40473c;
      32199: inst = 32'h8220000;
      32200: inst = 32'h10408000;
      32201: inst = 32'hc40473d;
      32202: inst = 32'h8220000;
      32203: inst = 32'h10408000;
      32204: inst = 32'hc40473e;
      32205: inst = 32'h8220000;
      32206: inst = 32'h10408000;
      32207: inst = 32'hc40473f;
      32208: inst = 32'h8220000;
      32209: inst = 32'h10408000;
      32210: inst = 32'hc404740;
      32211: inst = 32'h8220000;
      32212: inst = 32'h10408000;
      32213: inst = 32'hc404741;
      32214: inst = 32'h8220000;
      32215: inst = 32'h10408000;
      32216: inst = 32'hc404742;
      32217: inst = 32'h8220000;
      32218: inst = 32'h10408000;
      32219: inst = 32'hc404743;
      32220: inst = 32'h8220000;
      32221: inst = 32'h10408000;
      32222: inst = 32'hc404744;
      32223: inst = 32'h8220000;
      32224: inst = 32'h10408000;
      32225: inst = 32'hc404745;
      32226: inst = 32'h8220000;
      32227: inst = 32'h10408000;
      32228: inst = 32'hc404746;
      32229: inst = 32'h8220000;
      32230: inst = 32'h10408000;
      32231: inst = 32'hc404747;
      32232: inst = 32'h8220000;
      32233: inst = 32'h10408000;
      32234: inst = 32'hc404748;
      32235: inst = 32'h8220000;
      32236: inst = 32'h10408000;
      32237: inst = 32'hc404749;
      32238: inst = 32'h8220000;
      32239: inst = 32'h10408000;
      32240: inst = 32'hc40474a;
      32241: inst = 32'h8220000;
      32242: inst = 32'h10408000;
      32243: inst = 32'hc40474b;
      32244: inst = 32'h8220000;
      32245: inst = 32'h10408000;
      32246: inst = 32'hc40474f;
      32247: inst = 32'h8220000;
      32248: inst = 32'h10408000;
      32249: inst = 32'hc404750;
      32250: inst = 32'h8220000;
      32251: inst = 32'h10408000;
      32252: inst = 32'hc404751;
      32253: inst = 32'h8220000;
      32254: inst = 32'h10408000;
      32255: inst = 32'hc404752;
      32256: inst = 32'h8220000;
      32257: inst = 32'h10408000;
      32258: inst = 32'hc404753;
      32259: inst = 32'h8220000;
      32260: inst = 32'h10408000;
      32261: inst = 32'hc404754;
      32262: inst = 32'h8220000;
      32263: inst = 32'h10408000;
      32264: inst = 32'hc404755;
      32265: inst = 32'h8220000;
      32266: inst = 32'h10408000;
      32267: inst = 32'hc404756;
      32268: inst = 32'h8220000;
      32269: inst = 32'h10408000;
      32270: inst = 32'hc404757;
      32271: inst = 32'h8220000;
      32272: inst = 32'h10408000;
      32273: inst = 32'hc404758;
      32274: inst = 32'h8220000;
      32275: inst = 32'h10408000;
      32276: inst = 32'hc404759;
      32277: inst = 32'h8220000;
      32278: inst = 32'h10408000;
      32279: inst = 32'hc40475a;
      32280: inst = 32'h8220000;
      32281: inst = 32'h10408000;
      32282: inst = 32'hc40475b;
      32283: inst = 32'h8220000;
      32284: inst = 32'h10408000;
      32285: inst = 32'hc40475c;
      32286: inst = 32'h8220000;
      32287: inst = 32'h10408000;
      32288: inst = 32'hc404763;
      32289: inst = 32'h8220000;
      32290: inst = 32'h10408000;
      32291: inst = 32'hc404764;
      32292: inst = 32'h8220000;
      32293: inst = 32'h10408000;
      32294: inst = 32'hc404765;
      32295: inst = 32'h8220000;
      32296: inst = 32'h10408000;
      32297: inst = 32'hc404766;
      32298: inst = 32'h8220000;
      32299: inst = 32'h10408000;
      32300: inst = 32'hc404767;
      32301: inst = 32'h8220000;
      32302: inst = 32'h10408000;
      32303: inst = 32'hc404768;
      32304: inst = 32'h8220000;
      32305: inst = 32'h10408000;
      32306: inst = 32'hc404769;
      32307: inst = 32'h8220000;
      32308: inst = 32'h10408000;
      32309: inst = 32'hc40476a;
      32310: inst = 32'h8220000;
      32311: inst = 32'h10408000;
      32312: inst = 32'hc40476b;
      32313: inst = 32'h8220000;
      32314: inst = 32'h10408000;
      32315: inst = 32'hc40476c;
      32316: inst = 32'h8220000;
      32317: inst = 32'h10408000;
      32318: inst = 32'hc40476d;
      32319: inst = 32'h8220000;
      32320: inst = 32'h10408000;
      32321: inst = 32'hc404771;
      32322: inst = 32'h8220000;
      32323: inst = 32'h10408000;
      32324: inst = 32'hc404772;
      32325: inst = 32'h8220000;
      32326: inst = 32'h10408000;
      32327: inst = 32'hc404773;
      32328: inst = 32'h8220000;
      32329: inst = 32'h10408000;
      32330: inst = 32'hc404774;
      32331: inst = 32'h8220000;
      32332: inst = 32'h10408000;
      32333: inst = 32'hc404775;
      32334: inst = 32'h8220000;
      32335: inst = 32'h10408000;
      32336: inst = 32'hc404776;
      32337: inst = 32'h8220000;
      32338: inst = 32'h10408000;
      32339: inst = 32'hc404777;
      32340: inst = 32'h8220000;
      32341: inst = 32'h10408000;
      32342: inst = 32'hc404778;
      32343: inst = 32'h8220000;
      32344: inst = 32'h10408000;
      32345: inst = 32'hc404779;
      32346: inst = 32'h8220000;
      32347: inst = 32'h10408000;
      32348: inst = 32'hc40477a;
      32349: inst = 32'h8220000;
      32350: inst = 32'h10408000;
      32351: inst = 32'hc40477b;
      32352: inst = 32'h8220000;
      32353: inst = 32'h10408000;
      32354: inst = 32'hc40477c;
      32355: inst = 32'h8220000;
      32356: inst = 32'h10408000;
      32357: inst = 32'hc40477d;
      32358: inst = 32'h8220000;
      32359: inst = 32'h10408000;
      32360: inst = 32'hc40477e;
      32361: inst = 32'h8220000;
      32362: inst = 32'h10408000;
      32363: inst = 32'hc40477f;
      32364: inst = 32'h8220000;
      32365: inst = 32'h10408000;
      32366: inst = 32'hc404780;
      32367: inst = 32'h8220000;
      32368: inst = 32'h10408000;
      32369: inst = 32'hc404781;
      32370: inst = 32'h8220000;
      32371: inst = 32'h10408000;
      32372: inst = 32'hc404782;
      32373: inst = 32'h8220000;
      32374: inst = 32'h10408000;
      32375: inst = 32'hc404783;
      32376: inst = 32'h8220000;
      32377: inst = 32'h10408000;
      32378: inst = 32'hc404784;
      32379: inst = 32'h8220000;
      32380: inst = 32'h10408000;
      32381: inst = 32'hc404785;
      32382: inst = 32'h8220000;
      32383: inst = 32'h10408000;
      32384: inst = 32'hc404786;
      32385: inst = 32'h8220000;
      32386: inst = 32'h10408000;
      32387: inst = 32'hc404787;
      32388: inst = 32'h8220000;
      32389: inst = 32'h10408000;
      32390: inst = 32'hc404788;
      32391: inst = 32'h8220000;
      32392: inst = 32'h10408000;
      32393: inst = 32'hc404789;
      32394: inst = 32'h8220000;
      32395: inst = 32'h10408000;
      32396: inst = 32'hc40478a;
      32397: inst = 32'h8220000;
      32398: inst = 32'h10408000;
      32399: inst = 32'hc404795;
      32400: inst = 32'h8220000;
      32401: inst = 32'h10408000;
      32402: inst = 32'hc404796;
      32403: inst = 32'h8220000;
      32404: inst = 32'h10408000;
      32405: inst = 32'hc404797;
      32406: inst = 32'h8220000;
      32407: inst = 32'h10408000;
      32408: inst = 32'hc404799;
      32409: inst = 32'h8220000;
      32410: inst = 32'h10408000;
      32411: inst = 32'hc40479a;
      32412: inst = 32'h8220000;
      32413: inst = 32'h10408000;
      32414: inst = 32'hc40479b;
      32415: inst = 32'h8220000;
      32416: inst = 32'h10408000;
      32417: inst = 32'hc40479c;
      32418: inst = 32'h8220000;
      32419: inst = 32'h10408000;
      32420: inst = 32'hc40479d;
      32421: inst = 32'h8220000;
      32422: inst = 32'h10408000;
      32423: inst = 32'hc40479e;
      32424: inst = 32'h8220000;
      32425: inst = 32'h10408000;
      32426: inst = 32'hc40479f;
      32427: inst = 32'h8220000;
      32428: inst = 32'h10408000;
      32429: inst = 32'hc4047a0;
      32430: inst = 32'h8220000;
      32431: inst = 32'h10408000;
      32432: inst = 32'hc4047a1;
      32433: inst = 32'h8220000;
      32434: inst = 32'h10408000;
      32435: inst = 32'hc4047a2;
      32436: inst = 32'h8220000;
      32437: inst = 32'h10408000;
      32438: inst = 32'hc4047a3;
      32439: inst = 32'h8220000;
      32440: inst = 32'h10408000;
      32441: inst = 32'hc4047a4;
      32442: inst = 32'h8220000;
      32443: inst = 32'h10408000;
      32444: inst = 32'hc4047a5;
      32445: inst = 32'h8220000;
      32446: inst = 32'h10408000;
      32447: inst = 32'hc4047a6;
      32448: inst = 32'h8220000;
      32449: inst = 32'h10408000;
      32450: inst = 32'hc4047a7;
      32451: inst = 32'h8220000;
      32452: inst = 32'h10408000;
      32453: inst = 32'hc4047a8;
      32454: inst = 32'h8220000;
      32455: inst = 32'h10408000;
      32456: inst = 32'hc4047a9;
      32457: inst = 32'h8220000;
      32458: inst = 32'h10408000;
      32459: inst = 32'hc4047aa;
      32460: inst = 32'h8220000;
      32461: inst = 32'h10408000;
      32462: inst = 32'hc4047ab;
      32463: inst = 32'h8220000;
      32464: inst = 32'h10408000;
      32465: inst = 32'hc4047af;
      32466: inst = 32'h8220000;
      32467: inst = 32'h10408000;
      32468: inst = 32'hc4047b0;
      32469: inst = 32'h8220000;
      32470: inst = 32'h10408000;
      32471: inst = 32'hc4047b1;
      32472: inst = 32'h8220000;
      32473: inst = 32'h10408000;
      32474: inst = 32'hc4047b2;
      32475: inst = 32'h8220000;
      32476: inst = 32'h10408000;
      32477: inst = 32'hc4047b3;
      32478: inst = 32'h8220000;
      32479: inst = 32'h10408000;
      32480: inst = 32'hc4047b4;
      32481: inst = 32'h8220000;
      32482: inst = 32'h10408000;
      32483: inst = 32'hc4047b5;
      32484: inst = 32'h8220000;
      32485: inst = 32'h10408000;
      32486: inst = 32'hc4047b6;
      32487: inst = 32'h8220000;
      32488: inst = 32'h10408000;
      32489: inst = 32'hc4047b7;
      32490: inst = 32'h8220000;
      32491: inst = 32'h10408000;
      32492: inst = 32'hc4047b8;
      32493: inst = 32'h8220000;
      32494: inst = 32'h10408000;
      32495: inst = 32'hc4047b9;
      32496: inst = 32'h8220000;
      32497: inst = 32'h10408000;
      32498: inst = 32'hc4047ba;
      32499: inst = 32'h8220000;
      32500: inst = 32'h10408000;
      32501: inst = 32'hc4047bb;
      32502: inst = 32'h8220000;
      32503: inst = 32'h10408000;
      32504: inst = 32'hc4047bc;
      32505: inst = 32'h8220000;
      32506: inst = 32'h10408000;
      32507: inst = 32'hc4047c3;
      32508: inst = 32'h8220000;
      32509: inst = 32'h10408000;
      32510: inst = 32'hc4047c4;
      32511: inst = 32'h8220000;
      32512: inst = 32'h10408000;
      32513: inst = 32'hc4047c5;
      32514: inst = 32'h8220000;
      32515: inst = 32'h10408000;
      32516: inst = 32'hc4047c6;
      32517: inst = 32'h8220000;
      32518: inst = 32'h10408000;
      32519: inst = 32'hc4047c7;
      32520: inst = 32'h8220000;
      32521: inst = 32'h10408000;
      32522: inst = 32'hc4047c8;
      32523: inst = 32'h8220000;
      32524: inst = 32'h10408000;
      32525: inst = 32'hc4047c9;
      32526: inst = 32'h8220000;
      32527: inst = 32'h10408000;
      32528: inst = 32'hc4047ca;
      32529: inst = 32'h8220000;
      32530: inst = 32'h10408000;
      32531: inst = 32'hc4047cb;
      32532: inst = 32'h8220000;
      32533: inst = 32'h10408000;
      32534: inst = 32'hc4047cc;
      32535: inst = 32'h8220000;
      32536: inst = 32'h10408000;
      32537: inst = 32'hc4047cd;
      32538: inst = 32'h8220000;
      32539: inst = 32'h10408000;
      32540: inst = 32'hc4047d1;
      32541: inst = 32'h8220000;
      32542: inst = 32'h10408000;
      32543: inst = 32'hc4047d2;
      32544: inst = 32'h8220000;
      32545: inst = 32'h10408000;
      32546: inst = 32'hc4047d3;
      32547: inst = 32'h8220000;
      32548: inst = 32'h10408000;
      32549: inst = 32'hc4047d4;
      32550: inst = 32'h8220000;
      32551: inst = 32'h10408000;
      32552: inst = 32'hc4047d5;
      32553: inst = 32'h8220000;
      32554: inst = 32'h10408000;
      32555: inst = 32'hc4047d6;
      32556: inst = 32'h8220000;
      32557: inst = 32'h10408000;
      32558: inst = 32'hc4047d7;
      32559: inst = 32'h8220000;
      32560: inst = 32'h10408000;
      32561: inst = 32'hc4047d8;
      32562: inst = 32'h8220000;
      32563: inst = 32'h10408000;
      32564: inst = 32'hc4047d9;
      32565: inst = 32'h8220000;
      32566: inst = 32'h10408000;
      32567: inst = 32'hc4047da;
      32568: inst = 32'h8220000;
      32569: inst = 32'h10408000;
      32570: inst = 32'hc4047db;
      32571: inst = 32'h8220000;
      32572: inst = 32'h10408000;
      32573: inst = 32'hc4047dc;
      32574: inst = 32'h8220000;
      32575: inst = 32'h10408000;
      32576: inst = 32'hc4047dd;
      32577: inst = 32'h8220000;
      32578: inst = 32'h10408000;
      32579: inst = 32'hc4047de;
      32580: inst = 32'h8220000;
      32581: inst = 32'h10408000;
      32582: inst = 32'hc4047df;
      32583: inst = 32'h8220000;
      32584: inst = 32'h10408000;
      32585: inst = 32'hc4047e0;
      32586: inst = 32'h8220000;
      32587: inst = 32'h10408000;
      32588: inst = 32'hc4047e1;
      32589: inst = 32'h8220000;
      32590: inst = 32'h10408000;
      32591: inst = 32'hc4047e2;
      32592: inst = 32'h8220000;
      32593: inst = 32'h10408000;
      32594: inst = 32'hc4047e3;
      32595: inst = 32'h8220000;
      32596: inst = 32'h10408000;
      32597: inst = 32'hc4047e4;
      32598: inst = 32'h8220000;
      32599: inst = 32'h10408000;
      32600: inst = 32'hc4047e5;
      32601: inst = 32'h8220000;
      32602: inst = 32'h10408000;
      32603: inst = 32'hc4047e6;
      32604: inst = 32'h8220000;
      32605: inst = 32'h10408000;
      32606: inst = 32'hc4047e7;
      32607: inst = 32'h8220000;
      32608: inst = 32'h10408000;
      32609: inst = 32'hc4047e8;
      32610: inst = 32'h8220000;
      32611: inst = 32'h10408000;
      32612: inst = 32'hc4047e9;
      32613: inst = 32'h8220000;
      32614: inst = 32'h10408000;
      32615: inst = 32'hc4047ea;
      32616: inst = 32'h8220000;
      32617: inst = 32'h10408000;
      32618: inst = 32'hc4047ee;
      32619: inst = 32'h8220000;
      32620: inst = 32'h10408000;
      32621: inst = 32'hc4047ef;
      32622: inst = 32'h8220000;
      32623: inst = 32'h10408000;
      32624: inst = 32'hc4047f6;
      32625: inst = 32'h8220000;
      32626: inst = 32'h10408000;
      32627: inst = 32'hc4047f7;
      32628: inst = 32'h8220000;
      32629: inst = 32'h10408000;
      32630: inst = 32'hc4047fa;
      32631: inst = 32'h8220000;
      32632: inst = 32'h10408000;
      32633: inst = 32'hc4047fb;
      32634: inst = 32'h8220000;
      32635: inst = 32'h10408000;
      32636: inst = 32'hc4047fc;
      32637: inst = 32'h8220000;
      32638: inst = 32'h10408000;
      32639: inst = 32'hc4047fd;
      32640: inst = 32'h8220000;
      32641: inst = 32'h10408000;
      32642: inst = 32'hc4047fe;
      32643: inst = 32'h8220000;
      32644: inst = 32'h10408000;
      32645: inst = 32'hc4047ff;
      32646: inst = 32'h8220000;
      32647: inst = 32'h10408000;
      32648: inst = 32'hc404800;
      32649: inst = 32'h8220000;
      32650: inst = 32'h10408000;
      32651: inst = 32'hc404801;
      32652: inst = 32'h8220000;
      32653: inst = 32'h10408000;
      32654: inst = 32'hc404802;
      32655: inst = 32'h8220000;
      32656: inst = 32'h10408000;
      32657: inst = 32'hc404803;
      32658: inst = 32'h8220000;
      32659: inst = 32'h10408000;
      32660: inst = 32'hc404804;
      32661: inst = 32'h8220000;
      32662: inst = 32'h10408000;
      32663: inst = 32'hc404805;
      32664: inst = 32'h8220000;
      32665: inst = 32'h10408000;
      32666: inst = 32'hc404806;
      32667: inst = 32'h8220000;
      32668: inst = 32'h10408000;
      32669: inst = 32'hc404807;
      32670: inst = 32'h8220000;
      32671: inst = 32'h10408000;
      32672: inst = 32'hc404808;
      32673: inst = 32'h8220000;
      32674: inst = 32'h10408000;
      32675: inst = 32'hc404809;
      32676: inst = 32'h8220000;
      32677: inst = 32'h10408000;
      32678: inst = 32'hc40480a;
      32679: inst = 32'h8220000;
      32680: inst = 32'h10408000;
      32681: inst = 32'hc40480b;
      32682: inst = 32'h8220000;
      32683: inst = 32'h10408000;
      32684: inst = 32'hc40480f;
      32685: inst = 32'h8220000;
      32686: inst = 32'h10408000;
      32687: inst = 32'hc404810;
      32688: inst = 32'h8220000;
      32689: inst = 32'h10408000;
      32690: inst = 32'hc404811;
      32691: inst = 32'h8220000;
      32692: inst = 32'h10408000;
      32693: inst = 32'hc404812;
      32694: inst = 32'h8220000;
      32695: inst = 32'h10408000;
      32696: inst = 32'hc404813;
      32697: inst = 32'h8220000;
      32698: inst = 32'h10408000;
      32699: inst = 32'hc404814;
      32700: inst = 32'h8220000;
      32701: inst = 32'h10408000;
      32702: inst = 32'hc404815;
      32703: inst = 32'h8220000;
      32704: inst = 32'h10408000;
      32705: inst = 32'hc404816;
      32706: inst = 32'h8220000;
      32707: inst = 32'h10408000;
      32708: inst = 32'hc404817;
      32709: inst = 32'h8220000;
      32710: inst = 32'h10408000;
      32711: inst = 32'hc404818;
      32712: inst = 32'h8220000;
      32713: inst = 32'h10408000;
      32714: inst = 32'hc404819;
      32715: inst = 32'h8220000;
      32716: inst = 32'h10408000;
      32717: inst = 32'hc40481a;
      32718: inst = 32'h8220000;
      32719: inst = 32'h10408000;
      32720: inst = 32'hc40481b;
      32721: inst = 32'h8220000;
      32722: inst = 32'h10408000;
      32723: inst = 32'hc40481c;
      32724: inst = 32'h8220000;
      32725: inst = 32'h10408000;
      32726: inst = 32'hc404823;
      32727: inst = 32'h8220000;
      32728: inst = 32'h10408000;
      32729: inst = 32'hc404824;
      32730: inst = 32'h8220000;
      32731: inst = 32'h10408000;
      32732: inst = 32'hc404825;
      32733: inst = 32'h8220000;
      32734: inst = 32'h10408000;
      32735: inst = 32'hc404826;
      32736: inst = 32'h8220000;
      32737: inst = 32'h10408000;
      32738: inst = 32'hc404827;
      32739: inst = 32'h8220000;
      32740: inst = 32'h10408000;
      32741: inst = 32'hc404828;
      32742: inst = 32'h8220000;
      32743: inst = 32'h10408000;
      32744: inst = 32'hc404829;
      32745: inst = 32'h8220000;
      32746: inst = 32'h10408000;
      32747: inst = 32'hc40482a;
      32748: inst = 32'h8220000;
      32749: inst = 32'h10408000;
      32750: inst = 32'hc40482b;
      32751: inst = 32'h8220000;
      32752: inst = 32'h10408000;
      32753: inst = 32'hc40482c;
      32754: inst = 32'h8220000;
      32755: inst = 32'h10408000;
      32756: inst = 32'hc40482d;
      32757: inst = 32'h8220000;
      32758: inst = 32'h10408000;
      32759: inst = 32'hc404831;
      32760: inst = 32'h8220000;
      32761: inst = 32'h10408000;
      32762: inst = 32'hc404832;
      32763: inst = 32'h8220000;
      32764: inst = 32'h10408000;
      32765: inst = 32'hc404833;
      32766: inst = 32'h8220000;
      32767: inst = 32'h10408000;
      32768: inst = 32'hc404834;
      32769: inst = 32'h8220000;
      32770: inst = 32'h10408000;
      32771: inst = 32'hc404835;
      32772: inst = 32'h8220000;
      32773: inst = 32'h10408000;
      32774: inst = 32'hc404836;
      32775: inst = 32'h8220000;
      32776: inst = 32'h10408000;
      32777: inst = 32'hc404837;
      32778: inst = 32'h8220000;
      32779: inst = 32'h10408000;
      32780: inst = 32'hc404838;
      32781: inst = 32'h8220000;
      32782: inst = 32'h10408000;
      32783: inst = 32'hc404839;
      32784: inst = 32'h8220000;
      32785: inst = 32'h10408000;
      32786: inst = 32'hc40483a;
      32787: inst = 32'h8220000;
      32788: inst = 32'h10408000;
      32789: inst = 32'hc40483b;
      32790: inst = 32'h8220000;
      32791: inst = 32'h10408000;
      32792: inst = 32'hc40483c;
      32793: inst = 32'h8220000;
      32794: inst = 32'h10408000;
      32795: inst = 32'hc40483d;
      32796: inst = 32'h8220000;
      32797: inst = 32'h10408000;
      32798: inst = 32'hc40483e;
      32799: inst = 32'h8220000;
      32800: inst = 32'h10408000;
      32801: inst = 32'hc40483f;
      32802: inst = 32'h8220000;
      32803: inst = 32'h10408000;
      32804: inst = 32'hc404840;
      32805: inst = 32'h8220000;
      32806: inst = 32'h10408000;
      32807: inst = 32'hc404841;
      32808: inst = 32'h8220000;
      32809: inst = 32'h10408000;
      32810: inst = 32'hc404842;
      32811: inst = 32'h8220000;
      32812: inst = 32'h10408000;
      32813: inst = 32'hc404843;
      32814: inst = 32'h8220000;
      32815: inst = 32'h10408000;
      32816: inst = 32'hc404844;
      32817: inst = 32'h8220000;
      32818: inst = 32'h10408000;
      32819: inst = 32'hc404845;
      32820: inst = 32'h8220000;
      32821: inst = 32'h10408000;
      32822: inst = 32'hc404846;
      32823: inst = 32'h8220000;
      32824: inst = 32'h10408000;
      32825: inst = 32'hc404847;
      32826: inst = 32'h8220000;
      32827: inst = 32'h10408000;
      32828: inst = 32'hc404848;
      32829: inst = 32'h8220000;
      32830: inst = 32'h10408000;
      32831: inst = 32'hc404849;
      32832: inst = 32'h8220000;
      32833: inst = 32'h10408000;
      32834: inst = 32'hc40484a;
      32835: inst = 32'h8220000;
      32836: inst = 32'h10408000;
      32837: inst = 32'hc40484b;
      32838: inst = 32'h8220000;
      32839: inst = 32'h10408000;
      32840: inst = 32'hc40484c;
      32841: inst = 32'h8220000;
      32842: inst = 32'h10408000;
      32843: inst = 32'hc40484d;
      32844: inst = 32'h8220000;
      32845: inst = 32'h10408000;
      32846: inst = 32'hc40484e;
      32847: inst = 32'h8220000;
      32848: inst = 32'h10408000;
      32849: inst = 32'hc40484f;
      32850: inst = 32'h8220000;
      32851: inst = 32'h10408000;
      32852: inst = 32'hc404850;
      32853: inst = 32'h8220000;
      32854: inst = 32'h10408000;
      32855: inst = 32'hc404851;
      32856: inst = 32'h8220000;
      32857: inst = 32'h10408000;
      32858: inst = 32'hc404852;
      32859: inst = 32'h8220000;
      32860: inst = 32'h10408000;
      32861: inst = 32'hc404853;
      32862: inst = 32'h8220000;
      32863: inst = 32'h10408000;
      32864: inst = 32'hc40485a;
      32865: inst = 32'h8220000;
      32866: inst = 32'h10408000;
      32867: inst = 32'hc40485b;
      32868: inst = 32'h8220000;
      32869: inst = 32'h10408000;
      32870: inst = 32'hc40485c;
      32871: inst = 32'h8220000;
      32872: inst = 32'h10408000;
      32873: inst = 32'hc40485d;
      32874: inst = 32'h8220000;
      32875: inst = 32'h10408000;
      32876: inst = 32'hc40485e;
      32877: inst = 32'h8220000;
      32878: inst = 32'h10408000;
      32879: inst = 32'hc40485f;
      32880: inst = 32'h8220000;
      32881: inst = 32'h10408000;
      32882: inst = 32'hc404860;
      32883: inst = 32'h8220000;
      32884: inst = 32'h10408000;
      32885: inst = 32'hc404861;
      32886: inst = 32'h8220000;
      32887: inst = 32'h10408000;
      32888: inst = 32'hc404862;
      32889: inst = 32'h8220000;
      32890: inst = 32'h10408000;
      32891: inst = 32'hc404863;
      32892: inst = 32'h8220000;
      32893: inst = 32'h10408000;
      32894: inst = 32'hc404864;
      32895: inst = 32'h8220000;
      32896: inst = 32'h10408000;
      32897: inst = 32'hc404865;
      32898: inst = 32'h8220000;
      32899: inst = 32'h10408000;
      32900: inst = 32'hc404866;
      32901: inst = 32'h8220000;
      32902: inst = 32'h10408000;
      32903: inst = 32'hc404867;
      32904: inst = 32'h8220000;
      32905: inst = 32'h10408000;
      32906: inst = 32'hc404868;
      32907: inst = 32'h8220000;
      32908: inst = 32'h10408000;
      32909: inst = 32'hc404869;
      32910: inst = 32'h8220000;
      32911: inst = 32'h10408000;
      32912: inst = 32'hc40486a;
      32913: inst = 32'h8220000;
      32914: inst = 32'h10408000;
      32915: inst = 32'hc40486b;
      32916: inst = 32'h8220000;
      32917: inst = 32'h10408000;
      32918: inst = 32'hc40486f;
      32919: inst = 32'h8220000;
      32920: inst = 32'h10408000;
      32921: inst = 32'hc404870;
      32922: inst = 32'h8220000;
      32923: inst = 32'h10408000;
      32924: inst = 32'hc404871;
      32925: inst = 32'h8220000;
      32926: inst = 32'h10408000;
      32927: inst = 32'hc404872;
      32928: inst = 32'h8220000;
      32929: inst = 32'h10408000;
      32930: inst = 32'hc404873;
      32931: inst = 32'h8220000;
      32932: inst = 32'h10408000;
      32933: inst = 32'hc404874;
      32934: inst = 32'h8220000;
      32935: inst = 32'h10408000;
      32936: inst = 32'hc404875;
      32937: inst = 32'h8220000;
      32938: inst = 32'h10408000;
      32939: inst = 32'hc404876;
      32940: inst = 32'h8220000;
      32941: inst = 32'h10408000;
      32942: inst = 32'hc404877;
      32943: inst = 32'h8220000;
      32944: inst = 32'h10408000;
      32945: inst = 32'hc404878;
      32946: inst = 32'h8220000;
      32947: inst = 32'h10408000;
      32948: inst = 32'hc404879;
      32949: inst = 32'h8220000;
      32950: inst = 32'h10408000;
      32951: inst = 32'hc40487a;
      32952: inst = 32'h8220000;
      32953: inst = 32'h10408000;
      32954: inst = 32'hc40487b;
      32955: inst = 32'h8220000;
      32956: inst = 32'h10408000;
      32957: inst = 32'hc40487c;
      32958: inst = 32'h8220000;
      32959: inst = 32'h10408000;
      32960: inst = 32'hc404883;
      32961: inst = 32'h8220000;
      32962: inst = 32'h10408000;
      32963: inst = 32'hc404884;
      32964: inst = 32'h8220000;
      32965: inst = 32'h10408000;
      32966: inst = 32'hc404885;
      32967: inst = 32'h8220000;
      32968: inst = 32'h10408000;
      32969: inst = 32'hc404886;
      32970: inst = 32'h8220000;
      32971: inst = 32'h10408000;
      32972: inst = 32'hc404887;
      32973: inst = 32'h8220000;
      32974: inst = 32'h10408000;
      32975: inst = 32'hc404888;
      32976: inst = 32'h8220000;
      32977: inst = 32'h10408000;
      32978: inst = 32'hc404889;
      32979: inst = 32'h8220000;
      32980: inst = 32'h10408000;
      32981: inst = 32'hc40488a;
      32982: inst = 32'h8220000;
      32983: inst = 32'h10408000;
      32984: inst = 32'hc40488b;
      32985: inst = 32'h8220000;
      32986: inst = 32'h10408000;
      32987: inst = 32'hc40488c;
      32988: inst = 32'h8220000;
      32989: inst = 32'h10408000;
      32990: inst = 32'hc40488d;
      32991: inst = 32'h8220000;
      32992: inst = 32'h10408000;
      32993: inst = 32'hc404891;
      32994: inst = 32'h8220000;
      32995: inst = 32'h10408000;
      32996: inst = 32'hc404892;
      32997: inst = 32'h8220000;
      32998: inst = 32'h10408000;
      32999: inst = 32'hc404893;
      33000: inst = 32'h8220000;
      33001: inst = 32'h10408000;
      33002: inst = 32'hc404894;
      33003: inst = 32'h8220000;
      33004: inst = 32'h10408000;
      33005: inst = 32'hc404895;
      33006: inst = 32'h8220000;
      33007: inst = 32'h10408000;
      33008: inst = 32'hc404896;
      33009: inst = 32'h8220000;
      33010: inst = 32'h10408000;
      33011: inst = 32'hc404897;
      33012: inst = 32'h8220000;
      33013: inst = 32'h10408000;
      33014: inst = 32'hc404898;
      33015: inst = 32'h8220000;
      33016: inst = 32'h10408000;
      33017: inst = 32'hc404899;
      33018: inst = 32'h8220000;
      33019: inst = 32'h10408000;
      33020: inst = 32'hc40489a;
      33021: inst = 32'h8220000;
      33022: inst = 32'h10408000;
      33023: inst = 32'hc40489b;
      33024: inst = 32'h8220000;
      33025: inst = 32'h10408000;
      33026: inst = 32'hc40489c;
      33027: inst = 32'h8220000;
      33028: inst = 32'h10408000;
      33029: inst = 32'hc40489d;
      33030: inst = 32'h8220000;
      33031: inst = 32'h10408000;
      33032: inst = 32'hc40489e;
      33033: inst = 32'h8220000;
      33034: inst = 32'h10408000;
      33035: inst = 32'hc40489f;
      33036: inst = 32'h8220000;
      33037: inst = 32'h10408000;
      33038: inst = 32'hc4048a0;
      33039: inst = 32'h8220000;
      33040: inst = 32'h10408000;
      33041: inst = 32'hc4048a1;
      33042: inst = 32'h8220000;
      33043: inst = 32'h10408000;
      33044: inst = 32'hc4048a2;
      33045: inst = 32'h8220000;
      33046: inst = 32'h10408000;
      33047: inst = 32'hc4048a3;
      33048: inst = 32'h8220000;
      33049: inst = 32'h10408000;
      33050: inst = 32'hc4048a4;
      33051: inst = 32'h8220000;
      33052: inst = 32'h10408000;
      33053: inst = 32'hc4048a5;
      33054: inst = 32'h8220000;
      33055: inst = 32'h10408000;
      33056: inst = 32'hc4048a6;
      33057: inst = 32'h8220000;
      33058: inst = 32'h10408000;
      33059: inst = 32'hc4048a7;
      33060: inst = 32'h8220000;
      33061: inst = 32'h10408000;
      33062: inst = 32'hc4048a8;
      33063: inst = 32'h8220000;
      33064: inst = 32'h10408000;
      33065: inst = 32'hc4048a9;
      33066: inst = 32'h8220000;
      33067: inst = 32'h10408000;
      33068: inst = 32'hc4048aa;
      33069: inst = 32'h8220000;
      33070: inst = 32'h10408000;
      33071: inst = 32'hc4048ab;
      33072: inst = 32'h8220000;
      33073: inst = 32'h10408000;
      33074: inst = 32'hc4048ac;
      33075: inst = 32'h8220000;
      33076: inst = 32'h10408000;
      33077: inst = 32'hc4048ad;
      33078: inst = 32'h8220000;
      33079: inst = 32'h10408000;
      33080: inst = 32'hc4048ae;
      33081: inst = 32'h8220000;
      33082: inst = 32'h10408000;
      33083: inst = 32'hc4048af;
      33084: inst = 32'h8220000;
      33085: inst = 32'h10408000;
      33086: inst = 32'hc4048b0;
      33087: inst = 32'h8220000;
      33088: inst = 32'h10408000;
      33089: inst = 32'hc4048b1;
      33090: inst = 32'h8220000;
      33091: inst = 32'h10408000;
      33092: inst = 32'hc4048b2;
      33093: inst = 32'h8220000;
      33094: inst = 32'h10408000;
      33095: inst = 32'hc4048b3;
      33096: inst = 32'h8220000;
      33097: inst = 32'h10408000;
      33098: inst = 32'hc4048ba;
      33099: inst = 32'h8220000;
      33100: inst = 32'h10408000;
      33101: inst = 32'hc4048bb;
      33102: inst = 32'h8220000;
      33103: inst = 32'h10408000;
      33104: inst = 32'hc4048bc;
      33105: inst = 32'h8220000;
      33106: inst = 32'h10408000;
      33107: inst = 32'hc4048bd;
      33108: inst = 32'h8220000;
      33109: inst = 32'h10408000;
      33110: inst = 32'hc4048be;
      33111: inst = 32'h8220000;
      33112: inst = 32'h10408000;
      33113: inst = 32'hc4048bf;
      33114: inst = 32'h8220000;
      33115: inst = 32'h10408000;
      33116: inst = 32'hc4048c0;
      33117: inst = 32'h8220000;
      33118: inst = 32'h10408000;
      33119: inst = 32'hc4048c1;
      33120: inst = 32'h8220000;
      33121: inst = 32'h10408000;
      33122: inst = 32'hc4048c2;
      33123: inst = 32'h8220000;
      33124: inst = 32'h10408000;
      33125: inst = 32'hc4048c3;
      33126: inst = 32'h8220000;
      33127: inst = 32'h10408000;
      33128: inst = 32'hc4048c4;
      33129: inst = 32'h8220000;
      33130: inst = 32'h10408000;
      33131: inst = 32'hc4048c5;
      33132: inst = 32'h8220000;
      33133: inst = 32'h10408000;
      33134: inst = 32'hc4048c6;
      33135: inst = 32'h8220000;
      33136: inst = 32'h10408000;
      33137: inst = 32'hc4048c7;
      33138: inst = 32'h8220000;
      33139: inst = 32'h10408000;
      33140: inst = 32'hc4048c8;
      33141: inst = 32'h8220000;
      33142: inst = 32'h10408000;
      33143: inst = 32'hc4048c9;
      33144: inst = 32'h8220000;
      33145: inst = 32'h10408000;
      33146: inst = 32'hc4048ca;
      33147: inst = 32'h8220000;
      33148: inst = 32'h10408000;
      33149: inst = 32'hc4048cb;
      33150: inst = 32'h8220000;
      33151: inst = 32'h10408000;
      33152: inst = 32'hc4048cf;
      33153: inst = 32'h8220000;
      33154: inst = 32'h10408000;
      33155: inst = 32'hc4048d0;
      33156: inst = 32'h8220000;
      33157: inst = 32'h10408000;
      33158: inst = 32'hc4048d1;
      33159: inst = 32'h8220000;
      33160: inst = 32'h10408000;
      33161: inst = 32'hc4048d2;
      33162: inst = 32'h8220000;
      33163: inst = 32'h10408000;
      33164: inst = 32'hc4048d3;
      33165: inst = 32'h8220000;
      33166: inst = 32'h10408000;
      33167: inst = 32'hc4048d4;
      33168: inst = 32'h8220000;
      33169: inst = 32'h10408000;
      33170: inst = 32'hc4048d5;
      33171: inst = 32'h8220000;
      33172: inst = 32'h10408000;
      33173: inst = 32'hc4048d6;
      33174: inst = 32'h8220000;
      33175: inst = 32'h10408000;
      33176: inst = 32'hc4048d7;
      33177: inst = 32'h8220000;
      33178: inst = 32'h10408000;
      33179: inst = 32'hc4048d8;
      33180: inst = 32'h8220000;
      33181: inst = 32'h10408000;
      33182: inst = 32'hc4048d9;
      33183: inst = 32'h8220000;
      33184: inst = 32'h10408000;
      33185: inst = 32'hc4048da;
      33186: inst = 32'h8220000;
      33187: inst = 32'h10408000;
      33188: inst = 32'hc4048db;
      33189: inst = 32'h8220000;
      33190: inst = 32'h10408000;
      33191: inst = 32'hc4048dc;
      33192: inst = 32'h8220000;
      33193: inst = 32'h10408000;
      33194: inst = 32'hc4048e3;
      33195: inst = 32'h8220000;
      33196: inst = 32'h10408000;
      33197: inst = 32'hc4048e4;
      33198: inst = 32'h8220000;
      33199: inst = 32'h10408000;
      33200: inst = 32'hc4048e5;
      33201: inst = 32'h8220000;
      33202: inst = 32'h10408000;
      33203: inst = 32'hc4048e6;
      33204: inst = 32'h8220000;
      33205: inst = 32'h10408000;
      33206: inst = 32'hc4048e7;
      33207: inst = 32'h8220000;
      33208: inst = 32'h10408000;
      33209: inst = 32'hc4048e8;
      33210: inst = 32'h8220000;
      33211: inst = 32'h10408000;
      33212: inst = 32'hc4048e9;
      33213: inst = 32'h8220000;
      33214: inst = 32'h10408000;
      33215: inst = 32'hc4048ea;
      33216: inst = 32'h8220000;
      33217: inst = 32'h10408000;
      33218: inst = 32'hc4048eb;
      33219: inst = 32'h8220000;
      33220: inst = 32'h10408000;
      33221: inst = 32'hc4048ec;
      33222: inst = 32'h8220000;
      33223: inst = 32'h10408000;
      33224: inst = 32'hc4048ed;
      33225: inst = 32'h8220000;
      33226: inst = 32'h10408000;
      33227: inst = 32'hc4048f1;
      33228: inst = 32'h8220000;
      33229: inst = 32'h10408000;
      33230: inst = 32'hc4048f2;
      33231: inst = 32'h8220000;
      33232: inst = 32'h10408000;
      33233: inst = 32'hc4048f3;
      33234: inst = 32'h8220000;
      33235: inst = 32'h10408000;
      33236: inst = 32'hc4048f4;
      33237: inst = 32'h8220000;
      33238: inst = 32'h10408000;
      33239: inst = 32'hc4048f5;
      33240: inst = 32'h8220000;
      33241: inst = 32'h10408000;
      33242: inst = 32'hc4048f6;
      33243: inst = 32'h8220000;
      33244: inst = 32'h10408000;
      33245: inst = 32'hc4048f7;
      33246: inst = 32'h8220000;
      33247: inst = 32'h10408000;
      33248: inst = 32'hc4048f8;
      33249: inst = 32'h8220000;
      33250: inst = 32'h10408000;
      33251: inst = 32'hc4048f9;
      33252: inst = 32'h8220000;
      33253: inst = 32'h10408000;
      33254: inst = 32'hc4048fa;
      33255: inst = 32'h8220000;
      33256: inst = 32'h10408000;
      33257: inst = 32'hc4048fb;
      33258: inst = 32'h8220000;
      33259: inst = 32'h10408000;
      33260: inst = 32'hc4048fc;
      33261: inst = 32'h8220000;
      33262: inst = 32'h10408000;
      33263: inst = 32'hc4048fd;
      33264: inst = 32'h8220000;
      33265: inst = 32'h10408000;
      33266: inst = 32'hc4048fe;
      33267: inst = 32'h8220000;
      33268: inst = 32'h10408000;
      33269: inst = 32'hc4048ff;
      33270: inst = 32'h8220000;
      33271: inst = 32'h10408000;
      33272: inst = 32'hc404900;
      33273: inst = 32'h8220000;
      33274: inst = 32'h10408000;
      33275: inst = 32'hc404901;
      33276: inst = 32'h8220000;
      33277: inst = 32'h10408000;
      33278: inst = 32'hc404902;
      33279: inst = 32'h8220000;
      33280: inst = 32'h10408000;
      33281: inst = 32'hc404903;
      33282: inst = 32'h8220000;
      33283: inst = 32'h10408000;
      33284: inst = 32'hc404904;
      33285: inst = 32'h8220000;
      33286: inst = 32'h10408000;
      33287: inst = 32'hc404905;
      33288: inst = 32'h8220000;
      33289: inst = 32'h10408000;
      33290: inst = 32'hc404906;
      33291: inst = 32'h8220000;
      33292: inst = 32'h10408000;
      33293: inst = 32'hc404907;
      33294: inst = 32'h8220000;
      33295: inst = 32'h10408000;
      33296: inst = 32'hc404908;
      33297: inst = 32'h8220000;
      33298: inst = 32'h10408000;
      33299: inst = 32'hc404909;
      33300: inst = 32'h8220000;
      33301: inst = 32'h10408000;
      33302: inst = 32'hc40490a;
      33303: inst = 32'h8220000;
      33304: inst = 32'h10408000;
      33305: inst = 32'hc40490b;
      33306: inst = 32'h8220000;
      33307: inst = 32'h10408000;
      33308: inst = 32'hc40490c;
      33309: inst = 32'h8220000;
      33310: inst = 32'h10408000;
      33311: inst = 32'hc40490d;
      33312: inst = 32'h8220000;
      33313: inst = 32'h10408000;
      33314: inst = 32'hc40490e;
      33315: inst = 32'h8220000;
      33316: inst = 32'h10408000;
      33317: inst = 32'hc40490f;
      33318: inst = 32'h8220000;
      33319: inst = 32'h10408000;
      33320: inst = 32'hc404910;
      33321: inst = 32'h8220000;
      33322: inst = 32'h10408000;
      33323: inst = 32'hc404911;
      33324: inst = 32'h8220000;
      33325: inst = 32'h10408000;
      33326: inst = 32'hc404912;
      33327: inst = 32'h8220000;
      33328: inst = 32'h10408000;
      33329: inst = 32'hc404913;
      33330: inst = 32'h8220000;
      33331: inst = 32'h10408000;
      33332: inst = 32'hc404916;
      33333: inst = 32'h8220000;
      33334: inst = 32'h10408000;
      33335: inst = 32'hc40491a;
      33336: inst = 32'h8220000;
      33337: inst = 32'h10408000;
      33338: inst = 32'hc40491b;
      33339: inst = 32'h8220000;
      33340: inst = 32'h10408000;
      33341: inst = 32'hc40491c;
      33342: inst = 32'h8220000;
      33343: inst = 32'h10408000;
      33344: inst = 32'hc40491d;
      33345: inst = 32'h8220000;
      33346: inst = 32'h10408000;
      33347: inst = 32'hc40491e;
      33348: inst = 32'h8220000;
      33349: inst = 32'h10408000;
      33350: inst = 32'hc40491f;
      33351: inst = 32'h8220000;
      33352: inst = 32'h10408000;
      33353: inst = 32'hc404920;
      33354: inst = 32'h8220000;
      33355: inst = 32'h10408000;
      33356: inst = 32'hc404921;
      33357: inst = 32'h8220000;
      33358: inst = 32'h10408000;
      33359: inst = 32'hc404922;
      33360: inst = 32'h8220000;
      33361: inst = 32'h10408000;
      33362: inst = 32'hc404923;
      33363: inst = 32'h8220000;
      33364: inst = 32'h10408000;
      33365: inst = 32'hc404924;
      33366: inst = 32'h8220000;
      33367: inst = 32'h10408000;
      33368: inst = 32'hc404925;
      33369: inst = 32'h8220000;
      33370: inst = 32'h10408000;
      33371: inst = 32'hc404926;
      33372: inst = 32'h8220000;
      33373: inst = 32'h10408000;
      33374: inst = 32'hc404927;
      33375: inst = 32'h8220000;
      33376: inst = 32'h10408000;
      33377: inst = 32'hc404928;
      33378: inst = 32'h8220000;
      33379: inst = 32'h10408000;
      33380: inst = 32'hc404929;
      33381: inst = 32'h8220000;
      33382: inst = 32'h10408000;
      33383: inst = 32'hc40492a;
      33384: inst = 32'h8220000;
      33385: inst = 32'h10408000;
      33386: inst = 32'hc40492b;
      33387: inst = 32'h8220000;
      33388: inst = 32'h10408000;
      33389: inst = 32'hc40492f;
      33390: inst = 32'h8220000;
      33391: inst = 32'h10408000;
      33392: inst = 32'hc404930;
      33393: inst = 32'h8220000;
      33394: inst = 32'h10408000;
      33395: inst = 32'hc404931;
      33396: inst = 32'h8220000;
      33397: inst = 32'h10408000;
      33398: inst = 32'hc404932;
      33399: inst = 32'h8220000;
      33400: inst = 32'h10408000;
      33401: inst = 32'hc404933;
      33402: inst = 32'h8220000;
      33403: inst = 32'h10408000;
      33404: inst = 32'hc404934;
      33405: inst = 32'h8220000;
      33406: inst = 32'h10408000;
      33407: inst = 32'hc404935;
      33408: inst = 32'h8220000;
      33409: inst = 32'h10408000;
      33410: inst = 32'hc404936;
      33411: inst = 32'h8220000;
      33412: inst = 32'h10408000;
      33413: inst = 32'hc404937;
      33414: inst = 32'h8220000;
      33415: inst = 32'h10408000;
      33416: inst = 32'hc404938;
      33417: inst = 32'h8220000;
      33418: inst = 32'h10408000;
      33419: inst = 32'hc404939;
      33420: inst = 32'h8220000;
      33421: inst = 32'h10408000;
      33422: inst = 32'hc40493a;
      33423: inst = 32'h8220000;
      33424: inst = 32'h10408000;
      33425: inst = 32'hc40493b;
      33426: inst = 32'h8220000;
      33427: inst = 32'h10408000;
      33428: inst = 32'hc40493c;
      33429: inst = 32'h8220000;
      33430: inst = 32'h10408000;
      33431: inst = 32'hc404943;
      33432: inst = 32'h8220000;
      33433: inst = 32'h10408000;
      33434: inst = 32'hc404944;
      33435: inst = 32'h8220000;
      33436: inst = 32'h10408000;
      33437: inst = 32'hc404945;
      33438: inst = 32'h8220000;
      33439: inst = 32'h10408000;
      33440: inst = 32'hc404946;
      33441: inst = 32'h8220000;
      33442: inst = 32'h10408000;
      33443: inst = 32'hc404947;
      33444: inst = 32'h8220000;
      33445: inst = 32'h10408000;
      33446: inst = 32'hc404948;
      33447: inst = 32'h8220000;
      33448: inst = 32'h10408000;
      33449: inst = 32'hc404949;
      33450: inst = 32'h8220000;
      33451: inst = 32'h10408000;
      33452: inst = 32'hc40494a;
      33453: inst = 32'h8220000;
      33454: inst = 32'h10408000;
      33455: inst = 32'hc40494b;
      33456: inst = 32'h8220000;
      33457: inst = 32'h10408000;
      33458: inst = 32'hc40494c;
      33459: inst = 32'h8220000;
      33460: inst = 32'h10408000;
      33461: inst = 32'hc40494d;
      33462: inst = 32'h8220000;
      33463: inst = 32'h10408000;
      33464: inst = 32'hc404951;
      33465: inst = 32'h8220000;
      33466: inst = 32'h10408000;
      33467: inst = 32'hc404952;
      33468: inst = 32'h8220000;
      33469: inst = 32'h10408000;
      33470: inst = 32'hc404953;
      33471: inst = 32'h8220000;
      33472: inst = 32'h10408000;
      33473: inst = 32'hc404954;
      33474: inst = 32'h8220000;
      33475: inst = 32'h10408000;
      33476: inst = 32'hc404955;
      33477: inst = 32'h8220000;
      33478: inst = 32'h10408000;
      33479: inst = 32'hc404956;
      33480: inst = 32'h8220000;
      33481: inst = 32'h10408000;
      33482: inst = 32'hc404957;
      33483: inst = 32'h8220000;
      33484: inst = 32'h10408000;
      33485: inst = 32'hc404958;
      33486: inst = 32'h8220000;
      33487: inst = 32'h10408000;
      33488: inst = 32'hc404959;
      33489: inst = 32'h8220000;
      33490: inst = 32'h10408000;
      33491: inst = 32'hc40495a;
      33492: inst = 32'h8220000;
      33493: inst = 32'h10408000;
      33494: inst = 32'hc40495b;
      33495: inst = 32'h8220000;
      33496: inst = 32'h10408000;
      33497: inst = 32'hc40495c;
      33498: inst = 32'h8220000;
      33499: inst = 32'h10408000;
      33500: inst = 32'hc40495d;
      33501: inst = 32'h8220000;
      33502: inst = 32'h10408000;
      33503: inst = 32'hc40495e;
      33504: inst = 32'h8220000;
      33505: inst = 32'h10408000;
      33506: inst = 32'hc40495f;
      33507: inst = 32'h8220000;
      33508: inst = 32'h10408000;
      33509: inst = 32'hc404960;
      33510: inst = 32'h8220000;
      33511: inst = 32'h10408000;
      33512: inst = 32'hc404961;
      33513: inst = 32'h8220000;
      33514: inst = 32'h10408000;
      33515: inst = 32'hc404962;
      33516: inst = 32'h8220000;
      33517: inst = 32'h10408000;
      33518: inst = 32'hc404963;
      33519: inst = 32'h8220000;
      33520: inst = 32'h10408000;
      33521: inst = 32'hc404964;
      33522: inst = 32'h8220000;
      33523: inst = 32'h10408000;
      33524: inst = 32'hc404965;
      33525: inst = 32'h8220000;
      33526: inst = 32'h10408000;
      33527: inst = 32'hc404966;
      33528: inst = 32'h8220000;
      33529: inst = 32'h10408000;
      33530: inst = 32'hc404967;
      33531: inst = 32'h8220000;
      33532: inst = 32'h10408000;
      33533: inst = 32'hc404968;
      33534: inst = 32'h8220000;
      33535: inst = 32'h10408000;
      33536: inst = 32'hc404969;
      33537: inst = 32'h8220000;
      33538: inst = 32'h10408000;
      33539: inst = 32'hc40496a;
      33540: inst = 32'h8220000;
      33541: inst = 32'h10408000;
      33542: inst = 32'hc40496b;
      33543: inst = 32'h8220000;
      33544: inst = 32'h10408000;
      33545: inst = 32'hc40496c;
      33546: inst = 32'h8220000;
      33547: inst = 32'h10408000;
      33548: inst = 32'hc40496d;
      33549: inst = 32'h8220000;
      33550: inst = 32'h10408000;
      33551: inst = 32'hc40496e;
      33552: inst = 32'h8220000;
      33553: inst = 32'h10408000;
      33554: inst = 32'hc40496f;
      33555: inst = 32'h8220000;
      33556: inst = 32'h10408000;
      33557: inst = 32'hc404970;
      33558: inst = 32'h8220000;
      33559: inst = 32'h10408000;
      33560: inst = 32'hc404971;
      33561: inst = 32'h8220000;
      33562: inst = 32'h10408000;
      33563: inst = 32'hc404972;
      33564: inst = 32'h8220000;
      33565: inst = 32'h10408000;
      33566: inst = 32'hc404973;
      33567: inst = 32'h8220000;
      33568: inst = 32'h10408000;
      33569: inst = 32'hc404974;
      33570: inst = 32'h8220000;
      33571: inst = 32'h10408000;
      33572: inst = 32'hc404975;
      33573: inst = 32'h8220000;
      33574: inst = 32'h10408000;
      33575: inst = 32'hc404976;
      33576: inst = 32'h8220000;
      33577: inst = 32'h10408000;
      33578: inst = 32'hc404977;
      33579: inst = 32'h8220000;
      33580: inst = 32'h10408000;
      33581: inst = 32'hc404978;
      33582: inst = 32'h8220000;
      33583: inst = 32'h10408000;
      33584: inst = 32'hc404979;
      33585: inst = 32'h8220000;
      33586: inst = 32'h10408000;
      33587: inst = 32'hc40497a;
      33588: inst = 32'h8220000;
      33589: inst = 32'h10408000;
      33590: inst = 32'hc40497b;
      33591: inst = 32'h8220000;
      33592: inst = 32'h10408000;
      33593: inst = 32'hc40497c;
      33594: inst = 32'h8220000;
      33595: inst = 32'h10408000;
      33596: inst = 32'hc40497d;
      33597: inst = 32'h8220000;
      33598: inst = 32'h10408000;
      33599: inst = 32'hc40497e;
      33600: inst = 32'h8220000;
      33601: inst = 32'h10408000;
      33602: inst = 32'hc40497f;
      33603: inst = 32'h8220000;
      33604: inst = 32'h10408000;
      33605: inst = 32'hc404980;
      33606: inst = 32'h8220000;
      33607: inst = 32'h10408000;
      33608: inst = 32'hc404981;
      33609: inst = 32'h8220000;
      33610: inst = 32'h10408000;
      33611: inst = 32'hc404982;
      33612: inst = 32'h8220000;
      33613: inst = 32'h10408000;
      33614: inst = 32'hc404983;
      33615: inst = 32'h8220000;
      33616: inst = 32'h10408000;
      33617: inst = 32'hc404984;
      33618: inst = 32'h8220000;
      33619: inst = 32'h10408000;
      33620: inst = 32'hc404985;
      33621: inst = 32'h8220000;
      33622: inst = 32'h10408000;
      33623: inst = 32'hc40498f;
      33624: inst = 32'h8220000;
      33625: inst = 32'h10408000;
      33626: inst = 32'hc404990;
      33627: inst = 32'h8220000;
      33628: inst = 32'h10408000;
      33629: inst = 32'hc404991;
      33630: inst = 32'h8220000;
      33631: inst = 32'h10408000;
      33632: inst = 32'hc404992;
      33633: inst = 32'h8220000;
      33634: inst = 32'h10408000;
      33635: inst = 32'hc404993;
      33636: inst = 32'h8220000;
      33637: inst = 32'h10408000;
      33638: inst = 32'hc404994;
      33639: inst = 32'h8220000;
      33640: inst = 32'h10408000;
      33641: inst = 32'hc404995;
      33642: inst = 32'h8220000;
      33643: inst = 32'h10408000;
      33644: inst = 32'hc404996;
      33645: inst = 32'h8220000;
      33646: inst = 32'h10408000;
      33647: inst = 32'hc404997;
      33648: inst = 32'h8220000;
      33649: inst = 32'h10408000;
      33650: inst = 32'hc404998;
      33651: inst = 32'h8220000;
      33652: inst = 32'h10408000;
      33653: inst = 32'hc404999;
      33654: inst = 32'h8220000;
      33655: inst = 32'h10408000;
      33656: inst = 32'hc40499a;
      33657: inst = 32'h8220000;
      33658: inst = 32'h10408000;
      33659: inst = 32'hc40499b;
      33660: inst = 32'h8220000;
      33661: inst = 32'h10408000;
      33662: inst = 32'hc40499c;
      33663: inst = 32'h8220000;
      33664: inst = 32'h10408000;
      33665: inst = 32'hc4049a3;
      33666: inst = 32'h8220000;
      33667: inst = 32'h10408000;
      33668: inst = 32'hc4049a4;
      33669: inst = 32'h8220000;
      33670: inst = 32'h10408000;
      33671: inst = 32'hc4049a5;
      33672: inst = 32'h8220000;
      33673: inst = 32'h10408000;
      33674: inst = 32'hc4049a6;
      33675: inst = 32'h8220000;
      33676: inst = 32'h10408000;
      33677: inst = 32'hc4049a7;
      33678: inst = 32'h8220000;
      33679: inst = 32'h10408000;
      33680: inst = 32'hc4049a8;
      33681: inst = 32'h8220000;
      33682: inst = 32'h10408000;
      33683: inst = 32'hc4049a9;
      33684: inst = 32'h8220000;
      33685: inst = 32'h10408000;
      33686: inst = 32'hc4049aa;
      33687: inst = 32'h8220000;
      33688: inst = 32'h10408000;
      33689: inst = 32'hc4049ab;
      33690: inst = 32'h8220000;
      33691: inst = 32'h10408000;
      33692: inst = 32'hc4049ac;
      33693: inst = 32'h8220000;
      33694: inst = 32'h10408000;
      33695: inst = 32'hc4049ad;
      33696: inst = 32'h8220000;
      33697: inst = 32'h10408000;
      33698: inst = 32'hc4049b1;
      33699: inst = 32'h8220000;
      33700: inst = 32'h10408000;
      33701: inst = 32'hc4049b2;
      33702: inst = 32'h8220000;
      33703: inst = 32'h10408000;
      33704: inst = 32'hc4049b3;
      33705: inst = 32'h8220000;
      33706: inst = 32'h10408000;
      33707: inst = 32'hc4049b4;
      33708: inst = 32'h8220000;
      33709: inst = 32'h10408000;
      33710: inst = 32'hc4049b5;
      33711: inst = 32'h8220000;
      33712: inst = 32'h10408000;
      33713: inst = 32'hc4049b6;
      33714: inst = 32'h8220000;
      33715: inst = 32'h10408000;
      33716: inst = 32'hc4049b7;
      33717: inst = 32'h8220000;
      33718: inst = 32'h10408000;
      33719: inst = 32'hc4049b8;
      33720: inst = 32'h8220000;
      33721: inst = 32'h10408000;
      33722: inst = 32'hc4049b9;
      33723: inst = 32'h8220000;
      33724: inst = 32'h10408000;
      33725: inst = 32'hc4049ba;
      33726: inst = 32'h8220000;
      33727: inst = 32'h10408000;
      33728: inst = 32'hc4049bb;
      33729: inst = 32'h8220000;
      33730: inst = 32'h10408000;
      33731: inst = 32'hc4049bc;
      33732: inst = 32'h8220000;
      33733: inst = 32'h10408000;
      33734: inst = 32'hc4049bd;
      33735: inst = 32'h8220000;
      33736: inst = 32'h10408000;
      33737: inst = 32'hc4049be;
      33738: inst = 32'h8220000;
      33739: inst = 32'h10408000;
      33740: inst = 32'hc4049bf;
      33741: inst = 32'h8220000;
      33742: inst = 32'h10408000;
      33743: inst = 32'hc4049c0;
      33744: inst = 32'h8220000;
      33745: inst = 32'h10408000;
      33746: inst = 32'hc4049c1;
      33747: inst = 32'h8220000;
      33748: inst = 32'h10408000;
      33749: inst = 32'hc4049c2;
      33750: inst = 32'h8220000;
      33751: inst = 32'h10408000;
      33752: inst = 32'hc4049c3;
      33753: inst = 32'h8220000;
      33754: inst = 32'h10408000;
      33755: inst = 32'hc4049c4;
      33756: inst = 32'h8220000;
      33757: inst = 32'h10408000;
      33758: inst = 32'hc4049c5;
      33759: inst = 32'h8220000;
      33760: inst = 32'h10408000;
      33761: inst = 32'hc4049c6;
      33762: inst = 32'h8220000;
      33763: inst = 32'h10408000;
      33764: inst = 32'hc4049c7;
      33765: inst = 32'h8220000;
      33766: inst = 32'h10408000;
      33767: inst = 32'hc4049c8;
      33768: inst = 32'h8220000;
      33769: inst = 32'h10408000;
      33770: inst = 32'hc4049c9;
      33771: inst = 32'h8220000;
      33772: inst = 32'h10408000;
      33773: inst = 32'hc4049ca;
      33774: inst = 32'h8220000;
      33775: inst = 32'h10408000;
      33776: inst = 32'hc4049cb;
      33777: inst = 32'h8220000;
      33778: inst = 32'h10408000;
      33779: inst = 32'hc4049cc;
      33780: inst = 32'h8220000;
      33781: inst = 32'h10408000;
      33782: inst = 32'hc4049cd;
      33783: inst = 32'h8220000;
      33784: inst = 32'h10408000;
      33785: inst = 32'hc4049ce;
      33786: inst = 32'h8220000;
      33787: inst = 32'h10408000;
      33788: inst = 32'hc4049cf;
      33789: inst = 32'h8220000;
      33790: inst = 32'h10408000;
      33791: inst = 32'hc4049d0;
      33792: inst = 32'h8220000;
      33793: inst = 32'h10408000;
      33794: inst = 32'hc4049d1;
      33795: inst = 32'h8220000;
      33796: inst = 32'h10408000;
      33797: inst = 32'hc4049d2;
      33798: inst = 32'h8220000;
      33799: inst = 32'h10408000;
      33800: inst = 32'hc4049d3;
      33801: inst = 32'h8220000;
      33802: inst = 32'h10408000;
      33803: inst = 32'hc4049d4;
      33804: inst = 32'h8220000;
      33805: inst = 32'h10408000;
      33806: inst = 32'hc4049d5;
      33807: inst = 32'h8220000;
      33808: inst = 32'h10408000;
      33809: inst = 32'hc4049d6;
      33810: inst = 32'h8220000;
      33811: inst = 32'h10408000;
      33812: inst = 32'hc4049d7;
      33813: inst = 32'h8220000;
      33814: inst = 32'h10408000;
      33815: inst = 32'hc4049d8;
      33816: inst = 32'h8220000;
      33817: inst = 32'h10408000;
      33818: inst = 32'hc4049d9;
      33819: inst = 32'h8220000;
      33820: inst = 32'h10408000;
      33821: inst = 32'hc4049da;
      33822: inst = 32'h8220000;
      33823: inst = 32'h10408000;
      33824: inst = 32'hc4049db;
      33825: inst = 32'h8220000;
      33826: inst = 32'h10408000;
      33827: inst = 32'hc4049dc;
      33828: inst = 32'h8220000;
      33829: inst = 32'h10408000;
      33830: inst = 32'hc4049dd;
      33831: inst = 32'h8220000;
      33832: inst = 32'h10408000;
      33833: inst = 32'hc4049de;
      33834: inst = 32'h8220000;
      33835: inst = 32'h10408000;
      33836: inst = 32'hc4049df;
      33837: inst = 32'h8220000;
      33838: inst = 32'h10408000;
      33839: inst = 32'hc4049e0;
      33840: inst = 32'h8220000;
      33841: inst = 32'h10408000;
      33842: inst = 32'hc4049e1;
      33843: inst = 32'h8220000;
      33844: inst = 32'h10408000;
      33845: inst = 32'hc4049e2;
      33846: inst = 32'h8220000;
      33847: inst = 32'h10408000;
      33848: inst = 32'hc4049e3;
      33849: inst = 32'h8220000;
      33850: inst = 32'h10408000;
      33851: inst = 32'hc4049e4;
      33852: inst = 32'h8220000;
      33853: inst = 32'h10408000;
      33854: inst = 32'hc4049e5;
      33855: inst = 32'h8220000;
      33856: inst = 32'h10408000;
      33857: inst = 32'hc4049ef;
      33858: inst = 32'h8220000;
      33859: inst = 32'h10408000;
      33860: inst = 32'hc4049f0;
      33861: inst = 32'h8220000;
      33862: inst = 32'h10408000;
      33863: inst = 32'hc4049f1;
      33864: inst = 32'h8220000;
      33865: inst = 32'h10408000;
      33866: inst = 32'hc4049f2;
      33867: inst = 32'h8220000;
      33868: inst = 32'h10408000;
      33869: inst = 32'hc4049f3;
      33870: inst = 32'h8220000;
      33871: inst = 32'h10408000;
      33872: inst = 32'hc4049f4;
      33873: inst = 32'h8220000;
      33874: inst = 32'h10408000;
      33875: inst = 32'hc4049f5;
      33876: inst = 32'h8220000;
      33877: inst = 32'h10408000;
      33878: inst = 32'hc4049f6;
      33879: inst = 32'h8220000;
      33880: inst = 32'h10408000;
      33881: inst = 32'hc4049f7;
      33882: inst = 32'h8220000;
      33883: inst = 32'h10408000;
      33884: inst = 32'hc4049f8;
      33885: inst = 32'h8220000;
      33886: inst = 32'h10408000;
      33887: inst = 32'hc4049f9;
      33888: inst = 32'h8220000;
      33889: inst = 32'h10408000;
      33890: inst = 32'hc4049fa;
      33891: inst = 32'h8220000;
      33892: inst = 32'h10408000;
      33893: inst = 32'hc4049fb;
      33894: inst = 32'h8220000;
      33895: inst = 32'h10408000;
      33896: inst = 32'hc4049fc;
      33897: inst = 32'h8220000;
      33898: inst = 32'h10408000;
      33899: inst = 32'hc404a03;
      33900: inst = 32'h8220000;
      33901: inst = 32'h10408000;
      33902: inst = 32'hc404a04;
      33903: inst = 32'h8220000;
      33904: inst = 32'h10408000;
      33905: inst = 32'hc404a05;
      33906: inst = 32'h8220000;
      33907: inst = 32'h10408000;
      33908: inst = 32'hc404a06;
      33909: inst = 32'h8220000;
      33910: inst = 32'h10408000;
      33911: inst = 32'hc404a07;
      33912: inst = 32'h8220000;
      33913: inst = 32'h10408000;
      33914: inst = 32'hc404a08;
      33915: inst = 32'h8220000;
      33916: inst = 32'h10408000;
      33917: inst = 32'hc404a09;
      33918: inst = 32'h8220000;
      33919: inst = 32'h10408000;
      33920: inst = 32'hc404a0a;
      33921: inst = 32'h8220000;
      33922: inst = 32'h10408000;
      33923: inst = 32'hc404a0b;
      33924: inst = 32'h8220000;
      33925: inst = 32'h10408000;
      33926: inst = 32'hc404a0c;
      33927: inst = 32'h8220000;
      33928: inst = 32'h10408000;
      33929: inst = 32'hc404a0d;
      33930: inst = 32'h8220000;
      33931: inst = 32'h10408000;
      33932: inst = 32'hc404a11;
      33933: inst = 32'h8220000;
      33934: inst = 32'h10408000;
      33935: inst = 32'hc404a12;
      33936: inst = 32'h8220000;
      33937: inst = 32'h10408000;
      33938: inst = 32'hc404a13;
      33939: inst = 32'h8220000;
      33940: inst = 32'h10408000;
      33941: inst = 32'hc404a14;
      33942: inst = 32'h8220000;
      33943: inst = 32'h10408000;
      33944: inst = 32'hc404a15;
      33945: inst = 32'h8220000;
      33946: inst = 32'h10408000;
      33947: inst = 32'hc404a16;
      33948: inst = 32'h8220000;
      33949: inst = 32'h10408000;
      33950: inst = 32'hc404a17;
      33951: inst = 32'h8220000;
      33952: inst = 32'h10408000;
      33953: inst = 32'hc404a18;
      33954: inst = 32'h8220000;
      33955: inst = 32'h10408000;
      33956: inst = 32'hc404a19;
      33957: inst = 32'h8220000;
      33958: inst = 32'h10408000;
      33959: inst = 32'hc404a1a;
      33960: inst = 32'h8220000;
      33961: inst = 32'h10408000;
      33962: inst = 32'hc404a1b;
      33963: inst = 32'h8220000;
      33964: inst = 32'h10408000;
      33965: inst = 32'hc404a1c;
      33966: inst = 32'h8220000;
      33967: inst = 32'h10408000;
      33968: inst = 32'hc404a1d;
      33969: inst = 32'h8220000;
      33970: inst = 32'h10408000;
      33971: inst = 32'hc404a1e;
      33972: inst = 32'h8220000;
      33973: inst = 32'h10408000;
      33974: inst = 32'hc404a1f;
      33975: inst = 32'h8220000;
      33976: inst = 32'h10408000;
      33977: inst = 32'hc404a20;
      33978: inst = 32'h8220000;
      33979: inst = 32'h10408000;
      33980: inst = 32'hc404a21;
      33981: inst = 32'h8220000;
      33982: inst = 32'h10408000;
      33983: inst = 32'hc404a22;
      33984: inst = 32'h8220000;
      33985: inst = 32'h10408000;
      33986: inst = 32'hc404a23;
      33987: inst = 32'h8220000;
      33988: inst = 32'h10408000;
      33989: inst = 32'hc404a24;
      33990: inst = 32'h8220000;
      33991: inst = 32'h10408000;
      33992: inst = 32'hc404a25;
      33993: inst = 32'h8220000;
      33994: inst = 32'h10408000;
      33995: inst = 32'hc404a26;
      33996: inst = 32'h8220000;
      33997: inst = 32'h10408000;
      33998: inst = 32'hc404a27;
      33999: inst = 32'h8220000;
      34000: inst = 32'h10408000;
      34001: inst = 32'hc404a28;
      34002: inst = 32'h8220000;
      34003: inst = 32'h10408000;
      34004: inst = 32'hc404a29;
      34005: inst = 32'h8220000;
      34006: inst = 32'h10408000;
      34007: inst = 32'hc404a2a;
      34008: inst = 32'h8220000;
      34009: inst = 32'h10408000;
      34010: inst = 32'hc404a2b;
      34011: inst = 32'h8220000;
      34012: inst = 32'h10408000;
      34013: inst = 32'hc404a2c;
      34014: inst = 32'h8220000;
      34015: inst = 32'h10408000;
      34016: inst = 32'hc404a2d;
      34017: inst = 32'h8220000;
      34018: inst = 32'h10408000;
      34019: inst = 32'hc404a2e;
      34020: inst = 32'h8220000;
      34021: inst = 32'h10408000;
      34022: inst = 32'hc404a2f;
      34023: inst = 32'h8220000;
      34024: inst = 32'h10408000;
      34025: inst = 32'hc404a30;
      34026: inst = 32'h8220000;
      34027: inst = 32'h10408000;
      34028: inst = 32'hc404a31;
      34029: inst = 32'h8220000;
      34030: inst = 32'h10408000;
      34031: inst = 32'hc404a32;
      34032: inst = 32'h8220000;
      34033: inst = 32'h10408000;
      34034: inst = 32'hc404a33;
      34035: inst = 32'h8220000;
      34036: inst = 32'h10408000;
      34037: inst = 32'hc404a34;
      34038: inst = 32'h8220000;
      34039: inst = 32'h10408000;
      34040: inst = 32'hc404a35;
      34041: inst = 32'h8220000;
      34042: inst = 32'h10408000;
      34043: inst = 32'hc404a36;
      34044: inst = 32'h8220000;
      34045: inst = 32'h10408000;
      34046: inst = 32'hc404a37;
      34047: inst = 32'h8220000;
      34048: inst = 32'h10408000;
      34049: inst = 32'hc404a38;
      34050: inst = 32'h8220000;
      34051: inst = 32'h10408000;
      34052: inst = 32'hc404a39;
      34053: inst = 32'h8220000;
      34054: inst = 32'h10408000;
      34055: inst = 32'hc404a3a;
      34056: inst = 32'h8220000;
      34057: inst = 32'h10408000;
      34058: inst = 32'hc404a3b;
      34059: inst = 32'h8220000;
      34060: inst = 32'h10408000;
      34061: inst = 32'hc404a3c;
      34062: inst = 32'h8220000;
      34063: inst = 32'h10408000;
      34064: inst = 32'hc404a3d;
      34065: inst = 32'h8220000;
      34066: inst = 32'h10408000;
      34067: inst = 32'hc404a3e;
      34068: inst = 32'h8220000;
      34069: inst = 32'h10408000;
      34070: inst = 32'hc404a3f;
      34071: inst = 32'h8220000;
      34072: inst = 32'h10408000;
      34073: inst = 32'hc404a40;
      34074: inst = 32'h8220000;
      34075: inst = 32'h10408000;
      34076: inst = 32'hc404a41;
      34077: inst = 32'h8220000;
      34078: inst = 32'h10408000;
      34079: inst = 32'hc404a42;
      34080: inst = 32'h8220000;
      34081: inst = 32'h10408000;
      34082: inst = 32'hc404a43;
      34083: inst = 32'h8220000;
      34084: inst = 32'h10408000;
      34085: inst = 32'hc404a44;
      34086: inst = 32'h8220000;
      34087: inst = 32'h10408000;
      34088: inst = 32'hc404a45;
      34089: inst = 32'h8220000;
      34090: inst = 32'h10408000;
      34091: inst = 32'hc404a4f;
      34092: inst = 32'h8220000;
      34093: inst = 32'h10408000;
      34094: inst = 32'hc404a50;
      34095: inst = 32'h8220000;
      34096: inst = 32'h10408000;
      34097: inst = 32'hc404a51;
      34098: inst = 32'h8220000;
      34099: inst = 32'h10408000;
      34100: inst = 32'hc404a52;
      34101: inst = 32'h8220000;
      34102: inst = 32'h10408000;
      34103: inst = 32'hc404a53;
      34104: inst = 32'h8220000;
      34105: inst = 32'h10408000;
      34106: inst = 32'hc404a54;
      34107: inst = 32'h8220000;
      34108: inst = 32'h10408000;
      34109: inst = 32'hc404a55;
      34110: inst = 32'h8220000;
      34111: inst = 32'h10408000;
      34112: inst = 32'hc404a56;
      34113: inst = 32'h8220000;
      34114: inst = 32'h10408000;
      34115: inst = 32'hc404a57;
      34116: inst = 32'h8220000;
      34117: inst = 32'h10408000;
      34118: inst = 32'hc404a58;
      34119: inst = 32'h8220000;
      34120: inst = 32'h10408000;
      34121: inst = 32'hc404a59;
      34122: inst = 32'h8220000;
      34123: inst = 32'h10408000;
      34124: inst = 32'hc404a5a;
      34125: inst = 32'h8220000;
      34126: inst = 32'h10408000;
      34127: inst = 32'hc404a5b;
      34128: inst = 32'h8220000;
      34129: inst = 32'h10408000;
      34130: inst = 32'hc404a5c;
      34131: inst = 32'h8220000;
      34132: inst = 32'h10408000;
      34133: inst = 32'hc404a63;
      34134: inst = 32'h8220000;
      34135: inst = 32'h10408000;
      34136: inst = 32'hc404a64;
      34137: inst = 32'h8220000;
      34138: inst = 32'h10408000;
      34139: inst = 32'hc404a65;
      34140: inst = 32'h8220000;
      34141: inst = 32'h10408000;
      34142: inst = 32'hc404a66;
      34143: inst = 32'h8220000;
      34144: inst = 32'h10408000;
      34145: inst = 32'hc404a67;
      34146: inst = 32'h8220000;
      34147: inst = 32'h10408000;
      34148: inst = 32'hc404a68;
      34149: inst = 32'h8220000;
      34150: inst = 32'h10408000;
      34151: inst = 32'hc404a69;
      34152: inst = 32'h8220000;
      34153: inst = 32'h10408000;
      34154: inst = 32'hc404a6a;
      34155: inst = 32'h8220000;
      34156: inst = 32'h10408000;
      34157: inst = 32'hc404a6b;
      34158: inst = 32'h8220000;
      34159: inst = 32'h10408000;
      34160: inst = 32'hc404a6c;
      34161: inst = 32'h8220000;
      34162: inst = 32'h10408000;
      34163: inst = 32'hc404a6d;
      34164: inst = 32'h8220000;
      34165: inst = 32'h10408000;
      34166: inst = 32'hc404a71;
      34167: inst = 32'h8220000;
      34168: inst = 32'h10408000;
      34169: inst = 32'hc404a72;
      34170: inst = 32'h8220000;
      34171: inst = 32'h10408000;
      34172: inst = 32'hc404a73;
      34173: inst = 32'h8220000;
      34174: inst = 32'h10408000;
      34175: inst = 32'hc404a74;
      34176: inst = 32'h8220000;
      34177: inst = 32'h10408000;
      34178: inst = 32'hc404a75;
      34179: inst = 32'h8220000;
      34180: inst = 32'h10408000;
      34181: inst = 32'hc404a76;
      34182: inst = 32'h8220000;
      34183: inst = 32'h10408000;
      34184: inst = 32'hc404a77;
      34185: inst = 32'h8220000;
      34186: inst = 32'h10408000;
      34187: inst = 32'hc404a78;
      34188: inst = 32'h8220000;
      34189: inst = 32'h10408000;
      34190: inst = 32'hc404a79;
      34191: inst = 32'h8220000;
      34192: inst = 32'h10408000;
      34193: inst = 32'hc404a7a;
      34194: inst = 32'h8220000;
      34195: inst = 32'h10408000;
      34196: inst = 32'hc404a7b;
      34197: inst = 32'h8220000;
      34198: inst = 32'h10408000;
      34199: inst = 32'hc404a7c;
      34200: inst = 32'h8220000;
      34201: inst = 32'h10408000;
      34202: inst = 32'hc404a7d;
      34203: inst = 32'h8220000;
      34204: inst = 32'h10408000;
      34205: inst = 32'hc404a7e;
      34206: inst = 32'h8220000;
      34207: inst = 32'h10408000;
      34208: inst = 32'hc404a7f;
      34209: inst = 32'h8220000;
      34210: inst = 32'h10408000;
      34211: inst = 32'hc404a80;
      34212: inst = 32'h8220000;
      34213: inst = 32'h10408000;
      34214: inst = 32'hc404a81;
      34215: inst = 32'h8220000;
      34216: inst = 32'h10408000;
      34217: inst = 32'hc404a82;
      34218: inst = 32'h8220000;
      34219: inst = 32'h10408000;
      34220: inst = 32'hc404a83;
      34221: inst = 32'h8220000;
      34222: inst = 32'h10408000;
      34223: inst = 32'hc404a84;
      34224: inst = 32'h8220000;
      34225: inst = 32'h10408000;
      34226: inst = 32'hc404a85;
      34227: inst = 32'h8220000;
      34228: inst = 32'h10408000;
      34229: inst = 32'hc404a86;
      34230: inst = 32'h8220000;
      34231: inst = 32'h10408000;
      34232: inst = 32'hc404a87;
      34233: inst = 32'h8220000;
      34234: inst = 32'h10408000;
      34235: inst = 32'hc404a88;
      34236: inst = 32'h8220000;
      34237: inst = 32'h10408000;
      34238: inst = 32'hc404a89;
      34239: inst = 32'h8220000;
      34240: inst = 32'h10408000;
      34241: inst = 32'hc404a8a;
      34242: inst = 32'h8220000;
      34243: inst = 32'h10408000;
      34244: inst = 32'hc404a8b;
      34245: inst = 32'h8220000;
      34246: inst = 32'h10408000;
      34247: inst = 32'hc404a8c;
      34248: inst = 32'h8220000;
      34249: inst = 32'h10408000;
      34250: inst = 32'hc404a8d;
      34251: inst = 32'h8220000;
      34252: inst = 32'h10408000;
      34253: inst = 32'hc404a8e;
      34254: inst = 32'h8220000;
      34255: inst = 32'h10408000;
      34256: inst = 32'hc404a8f;
      34257: inst = 32'h8220000;
      34258: inst = 32'h10408000;
      34259: inst = 32'hc404a90;
      34260: inst = 32'h8220000;
      34261: inst = 32'h10408000;
      34262: inst = 32'hc404a91;
      34263: inst = 32'h8220000;
      34264: inst = 32'h10408000;
      34265: inst = 32'hc404a92;
      34266: inst = 32'h8220000;
      34267: inst = 32'h10408000;
      34268: inst = 32'hc404a93;
      34269: inst = 32'h8220000;
      34270: inst = 32'h10408000;
      34271: inst = 32'hc404a94;
      34272: inst = 32'h8220000;
      34273: inst = 32'h10408000;
      34274: inst = 32'hc404a95;
      34275: inst = 32'h8220000;
      34276: inst = 32'h10408000;
      34277: inst = 32'hc404a96;
      34278: inst = 32'h8220000;
      34279: inst = 32'h10408000;
      34280: inst = 32'hc404a97;
      34281: inst = 32'h8220000;
      34282: inst = 32'h10408000;
      34283: inst = 32'hc404a98;
      34284: inst = 32'h8220000;
      34285: inst = 32'h10408000;
      34286: inst = 32'hc404a99;
      34287: inst = 32'h8220000;
      34288: inst = 32'h10408000;
      34289: inst = 32'hc404a9a;
      34290: inst = 32'h8220000;
      34291: inst = 32'h10408000;
      34292: inst = 32'hc404a9b;
      34293: inst = 32'h8220000;
      34294: inst = 32'h10408000;
      34295: inst = 32'hc404a9c;
      34296: inst = 32'h8220000;
      34297: inst = 32'h10408000;
      34298: inst = 32'hc404a9d;
      34299: inst = 32'h8220000;
      34300: inst = 32'h10408000;
      34301: inst = 32'hc404a9e;
      34302: inst = 32'h8220000;
      34303: inst = 32'h10408000;
      34304: inst = 32'hc404a9f;
      34305: inst = 32'h8220000;
      34306: inst = 32'h10408000;
      34307: inst = 32'hc404aa0;
      34308: inst = 32'h8220000;
      34309: inst = 32'h10408000;
      34310: inst = 32'hc404aa1;
      34311: inst = 32'h8220000;
      34312: inst = 32'h10408000;
      34313: inst = 32'hc404aa2;
      34314: inst = 32'h8220000;
      34315: inst = 32'h10408000;
      34316: inst = 32'hc404aa3;
      34317: inst = 32'h8220000;
      34318: inst = 32'h10408000;
      34319: inst = 32'hc404aa4;
      34320: inst = 32'h8220000;
      34321: inst = 32'h10408000;
      34322: inst = 32'hc404aa5;
      34323: inst = 32'h8220000;
      34324: inst = 32'h10408000;
      34325: inst = 32'hc404aa6;
      34326: inst = 32'h8220000;
      34327: inst = 32'h10408000;
      34328: inst = 32'hc404aa7;
      34329: inst = 32'h8220000;
      34330: inst = 32'h10408000;
      34331: inst = 32'hc404aa8;
      34332: inst = 32'h8220000;
      34333: inst = 32'h10408000;
      34334: inst = 32'hc404aa9;
      34335: inst = 32'h8220000;
      34336: inst = 32'h10408000;
      34337: inst = 32'hc404aaa;
      34338: inst = 32'h8220000;
      34339: inst = 32'h10408000;
      34340: inst = 32'hc404aab;
      34341: inst = 32'h8220000;
      34342: inst = 32'h10408000;
      34343: inst = 32'hc404aac;
      34344: inst = 32'h8220000;
      34345: inst = 32'h10408000;
      34346: inst = 32'hc404aad;
      34347: inst = 32'h8220000;
      34348: inst = 32'h10408000;
      34349: inst = 32'hc404aae;
      34350: inst = 32'h8220000;
      34351: inst = 32'h10408000;
      34352: inst = 32'hc404aaf;
      34353: inst = 32'h8220000;
      34354: inst = 32'h10408000;
      34355: inst = 32'hc404ab0;
      34356: inst = 32'h8220000;
      34357: inst = 32'h10408000;
      34358: inst = 32'hc404ab1;
      34359: inst = 32'h8220000;
      34360: inst = 32'h10408000;
      34361: inst = 32'hc404ab2;
      34362: inst = 32'h8220000;
      34363: inst = 32'h10408000;
      34364: inst = 32'hc404ab3;
      34365: inst = 32'h8220000;
      34366: inst = 32'h10408000;
      34367: inst = 32'hc404ab4;
      34368: inst = 32'h8220000;
      34369: inst = 32'h10408000;
      34370: inst = 32'hc404ab5;
      34371: inst = 32'h8220000;
      34372: inst = 32'h10408000;
      34373: inst = 32'hc404ab6;
      34374: inst = 32'h8220000;
      34375: inst = 32'h10408000;
      34376: inst = 32'hc404ab7;
      34377: inst = 32'h8220000;
      34378: inst = 32'h10408000;
      34379: inst = 32'hc404ab8;
      34380: inst = 32'h8220000;
      34381: inst = 32'h10408000;
      34382: inst = 32'hc404ab9;
      34383: inst = 32'h8220000;
      34384: inst = 32'h10408000;
      34385: inst = 32'hc404aba;
      34386: inst = 32'h8220000;
      34387: inst = 32'h10408000;
      34388: inst = 32'hc404abb;
      34389: inst = 32'h8220000;
      34390: inst = 32'h10408000;
      34391: inst = 32'hc404abc;
      34392: inst = 32'h8220000;
      34393: inst = 32'h10408000;
      34394: inst = 32'hc404ac3;
      34395: inst = 32'h8220000;
      34396: inst = 32'h10408000;
      34397: inst = 32'hc404ac4;
      34398: inst = 32'h8220000;
      34399: inst = 32'h10408000;
      34400: inst = 32'hc404ac5;
      34401: inst = 32'h8220000;
      34402: inst = 32'h10408000;
      34403: inst = 32'hc404ac6;
      34404: inst = 32'h8220000;
      34405: inst = 32'h10408000;
      34406: inst = 32'hc404ac7;
      34407: inst = 32'h8220000;
      34408: inst = 32'h10408000;
      34409: inst = 32'hc404ac8;
      34410: inst = 32'h8220000;
      34411: inst = 32'h10408000;
      34412: inst = 32'hc404ac9;
      34413: inst = 32'h8220000;
      34414: inst = 32'h10408000;
      34415: inst = 32'hc404aca;
      34416: inst = 32'h8220000;
      34417: inst = 32'h10408000;
      34418: inst = 32'hc404acb;
      34419: inst = 32'h8220000;
      34420: inst = 32'h10408000;
      34421: inst = 32'hc404acc;
      34422: inst = 32'h8220000;
      34423: inst = 32'h10408000;
      34424: inst = 32'hc404acd;
      34425: inst = 32'h8220000;
      34426: inst = 32'h10408000;
      34427: inst = 32'hc404ad1;
      34428: inst = 32'h8220000;
      34429: inst = 32'h10408000;
      34430: inst = 32'hc404ad2;
      34431: inst = 32'h8220000;
      34432: inst = 32'h10408000;
      34433: inst = 32'hc404ad3;
      34434: inst = 32'h8220000;
      34435: inst = 32'h10408000;
      34436: inst = 32'hc404ad4;
      34437: inst = 32'h8220000;
      34438: inst = 32'h10408000;
      34439: inst = 32'hc404ad5;
      34440: inst = 32'h8220000;
      34441: inst = 32'h10408000;
      34442: inst = 32'hc404ad6;
      34443: inst = 32'h8220000;
      34444: inst = 32'h10408000;
      34445: inst = 32'hc404ad7;
      34446: inst = 32'h8220000;
      34447: inst = 32'h10408000;
      34448: inst = 32'hc404ad8;
      34449: inst = 32'h8220000;
      34450: inst = 32'h10408000;
      34451: inst = 32'hc404ad9;
      34452: inst = 32'h8220000;
      34453: inst = 32'h10408000;
      34454: inst = 32'hc404ada;
      34455: inst = 32'h8220000;
      34456: inst = 32'h10408000;
      34457: inst = 32'hc404adb;
      34458: inst = 32'h8220000;
      34459: inst = 32'h10408000;
      34460: inst = 32'hc404adc;
      34461: inst = 32'h8220000;
      34462: inst = 32'h10408000;
      34463: inst = 32'hc404add;
      34464: inst = 32'h8220000;
      34465: inst = 32'h10408000;
      34466: inst = 32'hc404ade;
      34467: inst = 32'h8220000;
      34468: inst = 32'h10408000;
      34469: inst = 32'hc404adf;
      34470: inst = 32'h8220000;
      34471: inst = 32'h10408000;
      34472: inst = 32'hc404ae0;
      34473: inst = 32'h8220000;
      34474: inst = 32'h10408000;
      34475: inst = 32'hc404ae1;
      34476: inst = 32'h8220000;
      34477: inst = 32'h10408000;
      34478: inst = 32'hc404ae2;
      34479: inst = 32'h8220000;
      34480: inst = 32'h10408000;
      34481: inst = 32'hc404ae3;
      34482: inst = 32'h8220000;
      34483: inst = 32'h10408000;
      34484: inst = 32'hc404ae4;
      34485: inst = 32'h8220000;
      34486: inst = 32'h10408000;
      34487: inst = 32'hc404ae5;
      34488: inst = 32'h8220000;
      34489: inst = 32'h10408000;
      34490: inst = 32'hc404ae6;
      34491: inst = 32'h8220000;
      34492: inst = 32'h10408000;
      34493: inst = 32'hc404ae7;
      34494: inst = 32'h8220000;
      34495: inst = 32'h10408000;
      34496: inst = 32'hc404ae8;
      34497: inst = 32'h8220000;
      34498: inst = 32'h10408000;
      34499: inst = 32'hc404ae9;
      34500: inst = 32'h8220000;
      34501: inst = 32'h10408000;
      34502: inst = 32'hc404aea;
      34503: inst = 32'h8220000;
      34504: inst = 32'h10408000;
      34505: inst = 32'hc404aeb;
      34506: inst = 32'h8220000;
      34507: inst = 32'h10408000;
      34508: inst = 32'hc404aec;
      34509: inst = 32'h8220000;
      34510: inst = 32'h10408000;
      34511: inst = 32'hc404aed;
      34512: inst = 32'h8220000;
      34513: inst = 32'h10408000;
      34514: inst = 32'hc404aee;
      34515: inst = 32'h8220000;
      34516: inst = 32'h10408000;
      34517: inst = 32'hc404aef;
      34518: inst = 32'h8220000;
      34519: inst = 32'h10408000;
      34520: inst = 32'hc404af0;
      34521: inst = 32'h8220000;
      34522: inst = 32'h10408000;
      34523: inst = 32'hc404af1;
      34524: inst = 32'h8220000;
      34525: inst = 32'h10408000;
      34526: inst = 32'hc404af2;
      34527: inst = 32'h8220000;
      34528: inst = 32'h10408000;
      34529: inst = 32'hc404af3;
      34530: inst = 32'h8220000;
      34531: inst = 32'h10408000;
      34532: inst = 32'hc404af4;
      34533: inst = 32'h8220000;
      34534: inst = 32'h10408000;
      34535: inst = 32'hc404af5;
      34536: inst = 32'h8220000;
      34537: inst = 32'h10408000;
      34538: inst = 32'hc404af6;
      34539: inst = 32'h8220000;
      34540: inst = 32'h10408000;
      34541: inst = 32'hc404af7;
      34542: inst = 32'h8220000;
      34543: inst = 32'h10408000;
      34544: inst = 32'hc404af8;
      34545: inst = 32'h8220000;
      34546: inst = 32'h10408000;
      34547: inst = 32'hc404af9;
      34548: inst = 32'h8220000;
      34549: inst = 32'h10408000;
      34550: inst = 32'hc404afa;
      34551: inst = 32'h8220000;
      34552: inst = 32'h10408000;
      34553: inst = 32'hc404afb;
      34554: inst = 32'h8220000;
      34555: inst = 32'h10408000;
      34556: inst = 32'hc404afc;
      34557: inst = 32'h8220000;
      34558: inst = 32'h10408000;
      34559: inst = 32'hc404afd;
      34560: inst = 32'h8220000;
      34561: inst = 32'h10408000;
      34562: inst = 32'hc404afe;
      34563: inst = 32'h8220000;
      34564: inst = 32'h10408000;
      34565: inst = 32'hc404aff;
      34566: inst = 32'h8220000;
      34567: inst = 32'h10408000;
      34568: inst = 32'hc404b00;
      34569: inst = 32'h8220000;
      34570: inst = 32'h10408000;
      34571: inst = 32'hc404b01;
      34572: inst = 32'h8220000;
      34573: inst = 32'h10408000;
      34574: inst = 32'hc404b02;
      34575: inst = 32'h8220000;
      34576: inst = 32'h10408000;
      34577: inst = 32'hc404b03;
      34578: inst = 32'h8220000;
      34579: inst = 32'h10408000;
      34580: inst = 32'hc404b04;
      34581: inst = 32'h8220000;
      34582: inst = 32'h10408000;
      34583: inst = 32'hc404b05;
      34584: inst = 32'h8220000;
      34585: inst = 32'h10408000;
      34586: inst = 32'hc404b06;
      34587: inst = 32'h8220000;
      34588: inst = 32'h10408000;
      34589: inst = 32'hc404b07;
      34590: inst = 32'h8220000;
      34591: inst = 32'h10408000;
      34592: inst = 32'hc404b08;
      34593: inst = 32'h8220000;
      34594: inst = 32'h10408000;
      34595: inst = 32'hc404b09;
      34596: inst = 32'h8220000;
      34597: inst = 32'h10408000;
      34598: inst = 32'hc404b0a;
      34599: inst = 32'h8220000;
      34600: inst = 32'h10408000;
      34601: inst = 32'hc404b0b;
      34602: inst = 32'h8220000;
      34603: inst = 32'h10408000;
      34604: inst = 32'hc404b0c;
      34605: inst = 32'h8220000;
      34606: inst = 32'h10408000;
      34607: inst = 32'hc404b0d;
      34608: inst = 32'h8220000;
      34609: inst = 32'h10408000;
      34610: inst = 32'hc404b0e;
      34611: inst = 32'h8220000;
      34612: inst = 32'h10408000;
      34613: inst = 32'hc404b0f;
      34614: inst = 32'h8220000;
      34615: inst = 32'h10408000;
      34616: inst = 32'hc404b10;
      34617: inst = 32'h8220000;
      34618: inst = 32'h10408000;
      34619: inst = 32'hc404b11;
      34620: inst = 32'h8220000;
      34621: inst = 32'h10408000;
      34622: inst = 32'hc404b12;
      34623: inst = 32'h8220000;
      34624: inst = 32'h10408000;
      34625: inst = 32'hc404b13;
      34626: inst = 32'h8220000;
      34627: inst = 32'h10408000;
      34628: inst = 32'hc404b14;
      34629: inst = 32'h8220000;
      34630: inst = 32'h10408000;
      34631: inst = 32'hc404b15;
      34632: inst = 32'h8220000;
      34633: inst = 32'h10408000;
      34634: inst = 32'hc404b16;
      34635: inst = 32'h8220000;
      34636: inst = 32'h10408000;
      34637: inst = 32'hc404b17;
      34638: inst = 32'h8220000;
      34639: inst = 32'h10408000;
      34640: inst = 32'hc404b18;
      34641: inst = 32'h8220000;
      34642: inst = 32'h10408000;
      34643: inst = 32'hc404b19;
      34644: inst = 32'h8220000;
      34645: inst = 32'h10408000;
      34646: inst = 32'hc404b1a;
      34647: inst = 32'h8220000;
      34648: inst = 32'h10408000;
      34649: inst = 32'hc404b1b;
      34650: inst = 32'h8220000;
      34651: inst = 32'h10408000;
      34652: inst = 32'hc404b1c;
      34653: inst = 32'h8220000;
      34654: inst = 32'h10408000;
      34655: inst = 32'hc404b31;
      34656: inst = 32'h8220000;
      34657: inst = 32'h10408000;
      34658: inst = 32'hc404b32;
      34659: inst = 32'h8220000;
      34660: inst = 32'h10408000;
      34661: inst = 32'hc404b33;
      34662: inst = 32'h8220000;
      34663: inst = 32'h10408000;
      34664: inst = 32'hc404b34;
      34665: inst = 32'h8220000;
      34666: inst = 32'h10408000;
      34667: inst = 32'hc404b35;
      34668: inst = 32'h8220000;
      34669: inst = 32'h10408000;
      34670: inst = 32'hc404b36;
      34671: inst = 32'h8220000;
      34672: inst = 32'h10408000;
      34673: inst = 32'hc404b37;
      34674: inst = 32'h8220000;
      34675: inst = 32'h10408000;
      34676: inst = 32'hc404b38;
      34677: inst = 32'h8220000;
      34678: inst = 32'h10408000;
      34679: inst = 32'hc404b39;
      34680: inst = 32'h8220000;
      34681: inst = 32'h10408000;
      34682: inst = 32'hc404b3a;
      34683: inst = 32'h8220000;
      34684: inst = 32'h10408000;
      34685: inst = 32'hc404b3b;
      34686: inst = 32'h8220000;
      34687: inst = 32'h10408000;
      34688: inst = 32'hc404b3c;
      34689: inst = 32'h8220000;
      34690: inst = 32'h10408000;
      34691: inst = 32'hc404b3d;
      34692: inst = 32'h8220000;
      34693: inst = 32'h10408000;
      34694: inst = 32'hc404b3e;
      34695: inst = 32'h8220000;
      34696: inst = 32'h10408000;
      34697: inst = 32'hc404b3f;
      34698: inst = 32'h8220000;
      34699: inst = 32'h10408000;
      34700: inst = 32'hc404b40;
      34701: inst = 32'h8220000;
      34702: inst = 32'h10408000;
      34703: inst = 32'hc404b41;
      34704: inst = 32'h8220000;
      34705: inst = 32'h10408000;
      34706: inst = 32'hc404b42;
      34707: inst = 32'h8220000;
      34708: inst = 32'h10408000;
      34709: inst = 32'hc404b43;
      34710: inst = 32'h8220000;
      34711: inst = 32'h10408000;
      34712: inst = 32'hc404b44;
      34713: inst = 32'h8220000;
      34714: inst = 32'h10408000;
      34715: inst = 32'hc404b45;
      34716: inst = 32'h8220000;
      34717: inst = 32'h10408000;
      34718: inst = 32'hc404b46;
      34719: inst = 32'h8220000;
      34720: inst = 32'h10408000;
      34721: inst = 32'hc404b47;
      34722: inst = 32'h8220000;
      34723: inst = 32'h10408000;
      34724: inst = 32'hc404b48;
      34725: inst = 32'h8220000;
      34726: inst = 32'h10408000;
      34727: inst = 32'hc404b49;
      34728: inst = 32'h8220000;
      34729: inst = 32'h10408000;
      34730: inst = 32'hc404b4a;
      34731: inst = 32'h8220000;
      34732: inst = 32'h10408000;
      34733: inst = 32'hc404b4b;
      34734: inst = 32'h8220000;
      34735: inst = 32'h10408000;
      34736: inst = 32'hc404b4c;
      34737: inst = 32'h8220000;
      34738: inst = 32'h10408000;
      34739: inst = 32'hc404b4d;
      34740: inst = 32'h8220000;
      34741: inst = 32'h10408000;
      34742: inst = 32'hc404b4e;
      34743: inst = 32'h8220000;
      34744: inst = 32'h10408000;
      34745: inst = 32'hc404b4f;
      34746: inst = 32'h8220000;
      34747: inst = 32'h10408000;
      34748: inst = 32'hc404b50;
      34749: inst = 32'h8220000;
      34750: inst = 32'h10408000;
      34751: inst = 32'hc404b51;
      34752: inst = 32'h8220000;
      34753: inst = 32'h10408000;
      34754: inst = 32'hc404b52;
      34755: inst = 32'h8220000;
      34756: inst = 32'h10408000;
      34757: inst = 32'hc404b53;
      34758: inst = 32'h8220000;
      34759: inst = 32'h10408000;
      34760: inst = 32'hc404b54;
      34761: inst = 32'h8220000;
      34762: inst = 32'h10408000;
      34763: inst = 32'hc404b55;
      34764: inst = 32'h8220000;
      34765: inst = 32'h10408000;
      34766: inst = 32'hc404b56;
      34767: inst = 32'h8220000;
      34768: inst = 32'h10408000;
      34769: inst = 32'hc404b57;
      34770: inst = 32'h8220000;
      34771: inst = 32'h10408000;
      34772: inst = 32'hc404b58;
      34773: inst = 32'h8220000;
      34774: inst = 32'h10408000;
      34775: inst = 32'hc404b59;
      34776: inst = 32'h8220000;
      34777: inst = 32'h10408000;
      34778: inst = 32'hc404b5a;
      34779: inst = 32'h8220000;
      34780: inst = 32'h10408000;
      34781: inst = 32'hc404b5b;
      34782: inst = 32'h8220000;
      34783: inst = 32'h10408000;
      34784: inst = 32'hc404b5c;
      34785: inst = 32'h8220000;
      34786: inst = 32'h10408000;
      34787: inst = 32'hc404b5d;
      34788: inst = 32'h8220000;
      34789: inst = 32'h10408000;
      34790: inst = 32'hc404b5e;
      34791: inst = 32'h8220000;
      34792: inst = 32'h10408000;
      34793: inst = 32'hc404b5f;
      34794: inst = 32'h8220000;
      34795: inst = 32'h10408000;
      34796: inst = 32'hc404b60;
      34797: inst = 32'h8220000;
      34798: inst = 32'h10408000;
      34799: inst = 32'hc404b61;
      34800: inst = 32'h8220000;
      34801: inst = 32'h10408000;
      34802: inst = 32'hc404b62;
      34803: inst = 32'h8220000;
      34804: inst = 32'h10408000;
      34805: inst = 32'hc404b63;
      34806: inst = 32'h8220000;
      34807: inst = 32'h10408000;
      34808: inst = 32'hc404b64;
      34809: inst = 32'h8220000;
      34810: inst = 32'h10408000;
      34811: inst = 32'hc404b65;
      34812: inst = 32'h8220000;
      34813: inst = 32'h10408000;
      34814: inst = 32'hc404b66;
      34815: inst = 32'h8220000;
      34816: inst = 32'h10408000;
      34817: inst = 32'hc404b67;
      34818: inst = 32'h8220000;
      34819: inst = 32'h10408000;
      34820: inst = 32'hc404b68;
      34821: inst = 32'h8220000;
      34822: inst = 32'h10408000;
      34823: inst = 32'hc404b69;
      34824: inst = 32'h8220000;
      34825: inst = 32'h10408000;
      34826: inst = 32'hc404b6a;
      34827: inst = 32'h8220000;
      34828: inst = 32'h10408000;
      34829: inst = 32'hc404b6b;
      34830: inst = 32'h8220000;
      34831: inst = 32'h10408000;
      34832: inst = 32'hc404b6c;
      34833: inst = 32'h8220000;
      34834: inst = 32'h10408000;
      34835: inst = 32'hc404b6d;
      34836: inst = 32'h8220000;
      34837: inst = 32'h10408000;
      34838: inst = 32'hc404b6e;
      34839: inst = 32'h8220000;
      34840: inst = 32'h10408000;
      34841: inst = 32'hc404b6f;
      34842: inst = 32'h8220000;
      34843: inst = 32'h10408000;
      34844: inst = 32'hc404b70;
      34845: inst = 32'h8220000;
      34846: inst = 32'h10408000;
      34847: inst = 32'hc404b71;
      34848: inst = 32'h8220000;
      34849: inst = 32'h10408000;
      34850: inst = 32'hc404b72;
      34851: inst = 32'h8220000;
      34852: inst = 32'h10408000;
      34853: inst = 32'hc404b73;
      34854: inst = 32'h8220000;
      34855: inst = 32'h10408000;
      34856: inst = 32'hc404b74;
      34857: inst = 32'h8220000;
      34858: inst = 32'h10408000;
      34859: inst = 32'hc404b75;
      34860: inst = 32'h8220000;
      34861: inst = 32'h10408000;
      34862: inst = 32'hc404b76;
      34863: inst = 32'h8220000;
      34864: inst = 32'h10408000;
      34865: inst = 32'hc404b77;
      34866: inst = 32'h8220000;
      34867: inst = 32'h10408000;
      34868: inst = 32'hc404b78;
      34869: inst = 32'h8220000;
      34870: inst = 32'h10408000;
      34871: inst = 32'hc404b79;
      34872: inst = 32'h8220000;
      34873: inst = 32'h10408000;
      34874: inst = 32'hc404b7a;
      34875: inst = 32'h8220000;
      34876: inst = 32'h10408000;
      34877: inst = 32'hc404b7b;
      34878: inst = 32'h8220000;
      34879: inst = 32'h10408000;
      34880: inst = 32'hc404b7c;
      34881: inst = 32'h8220000;
      34882: inst = 32'h10408000;
      34883: inst = 32'hc404b91;
      34884: inst = 32'h8220000;
      34885: inst = 32'h10408000;
      34886: inst = 32'hc404b92;
      34887: inst = 32'h8220000;
      34888: inst = 32'h10408000;
      34889: inst = 32'hc404b93;
      34890: inst = 32'h8220000;
      34891: inst = 32'h10408000;
      34892: inst = 32'hc404b94;
      34893: inst = 32'h8220000;
      34894: inst = 32'h10408000;
      34895: inst = 32'hc404b95;
      34896: inst = 32'h8220000;
      34897: inst = 32'h10408000;
      34898: inst = 32'hc404b96;
      34899: inst = 32'h8220000;
      34900: inst = 32'h10408000;
      34901: inst = 32'hc404b97;
      34902: inst = 32'h8220000;
      34903: inst = 32'h10408000;
      34904: inst = 32'hc404b98;
      34905: inst = 32'h8220000;
      34906: inst = 32'h10408000;
      34907: inst = 32'hc404b99;
      34908: inst = 32'h8220000;
      34909: inst = 32'h10408000;
      34910: inst = 32'hc404b9a;
      34911: inst = 32'h8220000;
      34912: inst = 32'h10408000;
      34913: inst = 32'hc404b9b;
      34914: inst = 32'h8220000;
      34915: inst = 32'h10408000;
      34916: inst = 32'hc404b9c;
      34917: inst = 32'h8220000;
      34918: inst = 32'h10408000;
      34919: inst = 32'hc404b9d;
      34920: inst = 32'h8220000;
      34921: inst = 32'h10408000;
      34922: inst = 32'hc404b9e;
      34923: inst = 32'h8220000;
      34924: inst = 32'h10408000;
      34925: inst = 32'hc404b9f;
      34926: inst = 32'h8220000;
      34927: inst = 32'h10408000;
      34928: inst = 32'hc404ba0;
      34929: inst = 32'h8220000;
      34930: inst = 32'h10408000;
      34931: inst = 32'hc404ba1;
      34932: inst = 32'h8220000;
      34933: inst = 32'h10408000;
      34934: inst = 32'hc404ba2;
      34935: inst = 32'h8220000;
      34936: inst = 32'h10408000;
      34937: inst = 32'hc404ba3;
      34938: inst = 32'h8220000;
      34939: inst = 32'h10408000;
      34940: inst = 32'hc404ba4;
      34941: inst = 32'h8220000;
      34942: inst = 32'h10408000;
      34943: inst = 32'hc404ba5;
      34944: inst = 32'h8220000;
      34945: inst = 32'h10408000;
      34946: inst = 32'hc404ba6;
      34947: inst = 32'h8220000;
      34948: inst = 32'h10408000;
      34949: inst = 32'hc404ba7;
      34950: inst = 32'h8220000;
      34951: inst = 32'h10408000;
      34952: inst = 32'hc404ba8;
      34953: inst = 32'h8220000;
      34954: inst = 32'h10408000;
      34955: inst = 32'hc404ba9;
      34956: inst = 32'h8220000;
      34957: inst = 32'h10408000;
      34958: inst = 32'hc404baa;
      34959: inst = 32'h8220000;
      34960: inst = 32'h10408000;
      34961: inst = 32'hc404bab;
      34962: inst = 32'h8220000;
      34963: inst = 32'h10408000;
      34964: inst = 32'hc404bac;
      34965: inst = 32'h8220000;
      34966: inst = 32'h10408000;
      34967: inst = 32'hc404bad;
      34968: inst = 32'h8220000;
      34969: inst = 32'h10408000;
      34970: inst = 32'hc404bae;
      34971: inst = 32'h8220000;
      34972: inst = 32'h10408000;
      34973: inst = 32'hc404baf;
      34974: inst = 32'h8220000;
      34975: inst = 32'h10408000;
      34976: inst = 32'hc404bb0;
      34977: inst = 32'h8220000;
      34978: inst = 32'h10408000;
      34979: inst = 32'hc404bb1;
      34980: inst = 32'h8220000;
      34981: inst = 32'h10408000;
      34982: inst = 32'hc404bb2;
      34983: inst = 32'h8220000;
      34984: inst = 32'h10408000;
      34985: inst = 32'hc404bb3;
      34986: inst = 32'h8220000;
      34987: inst = 32'h10408000;
      34988: inst = 32'hc404bb4;
      34989: inst = 32'h8220000;
      34990: inst = 32'h10408000;
      34991: inst = 32'hc404bb5;
      34992: inst = 32'h8220000;
      34993: inst = 32'h10408000;
      34994: inst = 32'hc404bb6;
      34995: inst = 32'h8220000;
      34996: inst = 32'h10408000;
      34997: inst = 32'hc404bb7;
      34998: inst = 32'h8220000;
      34999: inst = 32'h10408000;
      35000: inst = 32'hc404bb8;
      35001: inst = 32'h8220000;
      35002: inst = 32'h10408000;
      35003: inst = 32'hc404bb9;
      35004: inst = 32'h8220000;
      35005: inst = 32'h10408000;
      35006: inst = 32'hc404bba;
      35007: inst = 32'h8220000;
      35008: inst = 32'h10408000;
      35009: inst = 32'hc404bbb;
      35010: inst = 32'h8220000;
      35011: inst = 32'h10408000;
      35012: inst = 32'hc404bbc;
      35013: inst = 32'h8220000;
      35014: inst = 32'h10408000;
      35015: inst = 32'hc404bbd;
      35016: inst = 32'h8220000;
      35017: inst = 32'h10408000;
      35018: inst = 32'hc404bbe;
      35019: inst = 32'h8220000;
      35020: inst = 32'h10408000;
      35021: inst = 32'hc404bbf;
      35022: inst = 32'h8220000;
      35023: inst = 32'h10408000;
      35024: inst = 32'hc404bc0;
      35025: inst = 32'h8220000;
      35026: inst = 32'h10408000;
      35027: inst = 32'hc404bc1;
      35028: inst = 32'h8220000;
      35029: inst = 32'h10408000;
      35030: inst = 32'hc404bc2;
      35031: inst = 32'h8220000;
      35032: inst = 32'h10408000;
      35033: inst = 32'hc404bc3;
      35034: inst = 32'h8220000;
      35035: inst = 32'h10408000;
      35036: inst = 32'hc404bc4;
      35037: inst = 32'h8220000;
      35038: inst = 32'h10408000;
      35039: inst = 32'hc404bc5;
      35040: inst = 32'h8220000;
      35041: inst = 32'h10408000;
      35042: inst = 32'hc404bc6;
      35043: inst = 32'h8220000;
      35044: inst = 32'h10408000;
      35045: inst = 32'hc404bc7;
      35046: inst = 32'h8220000;
      35047: inst = 32'h10408000;
      35048: inst = 32'hc404bc8;
      35049: inst = 32'h8220000;
      35050: inst = 32'h10408000;
      35051: inst = 32'hc404bc9;
      35052: inst = 32'h8220000;
      35053: inst = 32'h10408000;
      35054: inst = 32'hc404bca;
      35055: inst = 32'h8220000;
      35056: inst = 32'h10408000;
      35057: inst = 32'hc404bcb;
      35058: inst = 32'h8220000;
      35059: inst = 32'h10408000;
      35060: inst = 32'hc404bcc;
      35061: inst = 32'h8220000;
      35062: inst = 32'h10408000;
      35063: inst = 32'hc404bcd;
      35064: inst = 32'h8220000;
      35065: inst = 32'h10408000;
      35066: inst = 32'hc404bce;
      35067: inst = 32'h8220000;
      35068: inst = 32'h10408000;
      35069: inst = 32'hc404bcf;
      35070: inst = 32'h8220000;
      35071: inst = 32'h10408000;
      35072: inst = 32'hc404bd0;
      35073: inst = 32'h8220000;
      35074: inst = 32'h10408000;
      35075: inst = 32'hc404bd1;
      35076: inst = 32'h8220000;
      35077: inst = 32'h10408000;
      35078: inst = 32'hc404bd2;
      35079: inst = 32'h8220000;
      35080: inst = 32'h10408000;
      35081: inst = 32'hc404bd3;
      35082: inst = 32'h8220000;
      35083: inst = 32'h10408000;
      35084: inst = 32'hc404bd4;
      35085: inst = 32'h8220000;
      35086: inst = 32'h10408000;
      35087: inst = 32'hc404bd5;
      35088: inst = 32'h8220000;
      35089: inst = 32'h10408000;
      35090: inst = 32'hc404bd6;
      35091: inst = 32'h8220000;
      35092: inst = 32'h10408000;
      35093: inst = 32'hc404bd7;
      35094: inst = 32'h8220000;
      35095: inst = 32'h10408000;
      35096: inst = 32'hc404bd8;
      35097: inst = 32'h8220000;
      35098: inst = 32'h10408000;
      35099: inst = 32'hc404bd9;
      35100: inst = 32'h8220000;
      35101: inst = 32'h10408000;
      35102: inst = 32'hc404bda;
      35103: inst = 32'h8220000;
      35104: inst = 32'h10408000;
      35105: inst = 32'hc404bdb;
      35106: inst = 32'h8220000;
      35107: inst = 32'h10408000;
      35108: inst = 32'hc404bdc;
      35109: inst = 32'h8220000;
      35110: inst = 32'h10408000;
      35111: inst = 32'hc404bf1;
      35112: inst = 32'h8220000;
      35113: inst = 32'h10408000;
      35114: inst = 32'hc404bf2;
      35115: inst = 32'h8220000;
      35116: inst = 32'h10408000;
      35117: inst = 32'hc404bf3;
      35118: inst = 32'h8220000;
      35119: inst = 32'h10408000;
      35120: inst = 32'hc404bf4;
      35121: inst = 32'h8220000;
      35122: inst = 32'h10408000;
      35123: inst = 32'hc404bf5;
      35124: inst = 32'h8220000;
      35125: inst = 32'h10408000;
      35126: inst = 32'hc404bf6;
      35127: inst = 32'h8220000;
      35128: inst = 32'h10408000;
      35129: inst = 32'hc404bf7;
      35130: inst = 32'h8220000;
      35131: inst = 32'h10408000;
      35132: inst = 32'hc404bf8;
      35133: inst = 32'h8220000;
      35134: inst = 32'h10408000;
      35135: inst = 32'hc404bf9;
      35136: inst = 32'h8220000;
      35137: inst = 32'h10408000;
      35138: inst = 32'hc404bfa;
      35139: inst = 32'h8220000;
      35140: inst = 32'h10408000;
      35141: inst = 32'hc404bfb;
      35142: inst = 32'h8220000;
      35143: inst = 32'h10408000;
      35144: inst = 32'hc404bfc;
      35145: inst = 32'h8220000;
      35146: inst = 32'h10408000;
      35147: inst = 32'hc404bfd;
      35148: inst = 32'h8220000;
      35149: inst = 32'h10408000;
      35150: inst = 32'hc404bfe;
      35151: inst = 32'h8220000;
      35152: inst = 32'h10408000;
      35153: inst = 32'hc404bff;
      35154: inst = 32'h8220000;
      35155: inst = 32'h10408000;
      35156: inst = 32'hc404c00;
      35157: inst = 32'h8220000;
      35158: inst = 32'h10408000;
      35159: inst = 32'hc404c01;
      35160: inst = 32'h8220000;
      35161: inst = 32'h10408000;
      35162: inst = 32'hc404c02;
      35163: inst = 32'h8220000;
      35164: inst = 32'h10408000;
      35165: inst = 32'hc404c03;
      35166: inst = 32'h8220000;
      35167: inst = 32'h10408000;
      35168: inst = 32'hc404c04;
      35169: inst = 32'h8220000;
      35170: inst = 32'h10408000;
      35171: inst = 32'hc404c05;
      35172: inst = 32'h8220000;
      35173: inst = 32'h10408000;
      35174: inst = 32'hc404c06;
      35175: inst = 32'h8220000;
      35176: inst = 32'h10408000;
      35177: inst = 32'hc404c07;
      35178: inst = 32'h8220000;
      35179: inst = 32'h10408000;
      35180: inst = 32'hc404c08;
      35181: inst = 32'h8220000;
      35182: inst = 32'h10408000;
      35183: inst = 32'hc404c09;
      35184: inst = 32'h8220000;
      35185: inst = 32'h10408000;
      35186: inst = 32'hc404c0a;
      35187: inst = 32'h8220000;
      35188: inst = 32'h10408000;
      35189: inst = 32'hc404c0b;
      35190: inst = 32'h8220000;
      35191: inst = 32'h10408000;
      35192: inst = 32'hc404c0c;
      35193: inst = 32'h8220000;
      35194: inst = 32'h10408000;
      35195: inst = 32'hc404c0d;
      35196: inst = 32'h8220000;
      35197: inst = 32'h10408000;
      35198: inst = 32'hc404c0e;
      35199: inst = 32'h8220000;
      35200: inst = 32'h10408000;
      35201: inst = 32'hc404c0f;
      35202: inst = 32'h8220000;
      35203: inst = 32'h10408000;
      35204: inst = 32'hc404c10;
      35205: inst = 32'h8220000;
      35206: inst = 32'h10408000;
      35207: inst = 32'hc404c11;
      35208: inst = 32'h8220000;
      35209: inst = 32'h10408000;
      35210: inst = 32'hc404c12;
      35211: inst = 32'h8220000;
      35212: inst = 32'h10408000;
      35213: inst = 32'hc404c13;
      35214: inst = 32'h8220000;
      35215: inst = 32'h10408000;
      35216: inst = 32'hc404c14;
      35217: inst = 32'h8220000;
      35218: inst = 32'h10408000;
      35219: inst = 32'hc404c15;
      35220: inst = 32'h8220000;
      35221: inst = 32'h10408000;
      35222: inst = 32'hc404c16;
      35223: inst = 32'h8220000;
      35224: inst = 32'h10408000;
      35225: inst = 32'hc404c17;
      35226: inst = 32'h8220000;
      35227: inst = 32'h10408000;
      35228: inst = 32'hc404c18;
      35229: inst = 32'h8220000;
      35230: inst = 32'h10408000;
      35231: inst = 32'hc404c19;
      35232: inst = 32'h8220000;
      35233: inst = 32'h10408000;
      35234: inst = 32'hc404c1a;
      35235: inst = 32'h8220000;
      35236: inst = 32'h10408000;
      35237: inst = 32'hc404c1b;
      35238: inst = 32'h8220000;
      35239: inst = 32'h10408000;
      35240: inst = 32'hc404c1c;
      35241: inst = 32'h8220000;
      35242: inst = 32'h10408000;
      35243: inst = 32'hc404c1d;
      35244: inst = 32'h8220000;
      35245: inst = 32'h10408000;
      35246: inst = 32'hc404c1e;
      35247: inst = 32'h8220000;
      35248: inst = 32'h10408000;
      35249: inst = 32'hc404c1f;
      35250: inst = 32'h8220000;
      35251: inst = 32'h10408000;
      35252: inst = 32'hc404c20;
      35253: inst = 32'h8220000;
      35254: inst = 32'h10408000;
      35255: inst = 32'hc404c21;
      35256: inst = 32'h8220000;
      35257: inst = 32'h10408000;
      35258: inst = 32'hc404c22;
      35259: inst = 32'h8220000;
      35260: inst = 32'h10408000;
      35261: inst = 32'hc404c23;
      35262: inst = 32'h8220000;
      35263: inst = 32'h10408000;
      35264: inst = 32'hc404c24;
      35265: inst = 32'h8220000;
      35266: inst = 32'h10408000;
      35267: inst = 32'hc404c25;
      35268: inst = 32'h8220000;
      35269: inst = 32'h10408000;
      35270: inst = 32'hc404c26;
      35271: inst = 32'h8220000;
      35272: inst = 32'h10408000;
      35273: inst = 32'hc404c27;
      35274: inst = 32'h8220000;
      35275: inst = 32'h10408000;
      35276: inst = 32'hc404c28;
      35277: inst = 32'h8220000;
      35278: inst = 32'h10408000;
      35279: inst = 32'hc404c29;
      35280: inst = 32'h8220000;
      35281: inst = 32'h10408000;
      35282: inst = 32'hc404c2a;
      35283: inst = 32'h8220000;
      35284: inst = 32'h10408000;
      35285: inst = 32'hc404c2b;
      35286: inst = 32'h8220000;
      35287: inst = 32'h10408000;
      35288: inst = 32'hc404c2c;
      35289: inst = 32'h8220000;
      35290: inst = 32'h10408000;
      35291: inst = 32'hc404c2d;
      35292: inst = 32'h8220000;
      35293: inst = 32'h10408000;
      35294: inst = 32'hc404c2e;
      35295: inst = 32'h8220000;
      35296: inst = 32'h10408000;
      35297: inst = 32'hc404c2f;
      35298: inst = 32'h8220000;
      35299: inst = 32'h10408000;
      35300: inst = 32'hc404c30;
      35301: inst = 32'h8220000;
      35302: inst = 32'h10408000;
      35303: inst = 32'hc404c31;
      35304: inst = 32'h8220000;
      35305: inst = 32'h10408000;
      35306: inst = 32'hc404c32;
      35307: inst = 32'h8220000;
      35308: inst = 32'h10408000;
      35309: inst = 32'hc404c33;
      35310: inst = 32'h8220000;
      35311: inst = 32'h10408000;
      35312: inst = 32'hc404c34;
      35313: inst = 32'h8220000;
      35314: inst = 32'h10408000;
      35315: inst = 32'hc404c35;
      35316: inst = 32'h8220000;
      35317: inst = 32'h10408000;
      35318: inst = 32'hc404c36;
      35319: inst = 32'h8220000;
      35320: inst = 32'h10408000;
      35321: inst = 32'hc404c37;
      35322: inst = 32'h8220000;
      35323: inst = 32'h10408000;
      35324: inst = 32'hc404c38;
      35325: inst = 32'h8220000;
      35326: inst = 32'h10408000;
      35327: inst = 32'hc404c39;
      35328: inst = 32'h8220000;
      35329: inst = 32'h10408000;
      35330: inst = 32'hc404c3a;
      35331: inst = 32'h8220000;
      35332: inst = 32'h10408000;
      35333: inst = 32'hc404c3b;
      35334: inst = 32'h8220000;
      35335: inst = 32'h10408000;
      35336: inst = 32'hc404c3c;
      35337: inst = 32'h8220000;
      35338: inst = 32'h10408000;
      35339: inst = 32'hc404c43;
      35340: inst = 32'h8220000;
      35341: inst = 32'h10408000;
      35342: inst = 32'hc404c44;
      35343: inst = 32'h8220000;
      35344: inst = 32'h10408000;
      35345: inst = 32'hc404c45;
      35346: inst = 32'h8220000;
      35347: inst = 32'h10408000;
      35348: inst = 32'hc404c46;
      35349: inst = 32'h8220000;
      35350: inst = 32'h10408000;
      35351: inst = 32'hc404c47;
      35352: inst = 32'h8220000;
      35353: inst = 32'h10408000;
      35354: inst = 32'hc404c48;
      35355: inst = 32'h8220000;
      35356: inst = 32'h10408000;
      35357: inst = 32'hc404c49;
      35358: inst = 32'h8220000;
      35359: inst = 32'h10408000;
      35360: inst = 32'hc404c4a;
      35361: inst = 32'h8220000;
      35362: inst = 32'h10408000;
      35363: inst = 32'hc404c4b;
      35364: inst = 32'h8220000;
      35365: inst = 32'h10408000;
      35366: inst = 32'hc404c4c;
      35367: inst = 32'h8220000;
      35368: inst = 32'h10408000;
      35369: inst = 32'hc404c4d;
      35370: inst = 32'h8220000;
      35371: inst = 32'h10408000;
      35372: inst = 32'hc404c4e;
      35373: inst = 32'h8220000;
      35374: inst = 32'h10408000;
      35375: inst = 32'hc404c4f;
      35376: inst = 32'h8220000;
      35377: inst = 32'h10408000;
      35378: inst = 32'hc404c50;
      35379: inst = 32'h8220000;
      35380: inst = 32'h10408000;
      35381: inst = 32'hc404c51;
      35382: inst = 32'h8220000;
      35383: inst = 32'h10408000;
      35384: inst = 32'hc404c52;
      35385: inst = 32'h8220000;
      35386: inst = 32'h10408000;
      35387: inst = 32'hc404c53;
      35388: inst = 32'h8220000;
      35389: inst = 32'h10408000;
      35390: inst = 32'hc404c54;
      35391: inst = 32'h8220000;
      35392: inst = 32'h10408000;
      35393: inst = 32'hc404c55;
      35394: inst = 32'h8220000;
      35395: inst = 32'h10408000;
      35396: inst = 32'hc404c56;
      35397: inst = 32'h8220000;
      35398: inst = 32'h10408000;
      35399: inst = 32'hc404c57;
      35400: inst = 32'h8220000;
      35401: inst = 32'h10408000;
      35402: inst = 32'hc404c58;
      35403: inst = 32'h8220000;
      35404: inst = 32'h10408000;
      35405: inst = 32'hc404c59;
      35406: inst = 32'h8220000;
      35407: inst = 32'h10408000;
      35408: inst = 32'hc404c5a;
      35409: inst = 32'h8220000;
      35410: inst = 32'h10408000;
      35411: inst = 32'hc404c5b;
      35412: inst = 32'h8220000;
      35413: inst = 32'h10408000;
      35414: inst = 32'hc404c5c;
      35415: inst = 32'h8220000;
      35416: inst = 32'h10408000;
      35417: inst = 32'hc404c5d;
      35418: inst = 32'h8220000;
      35419: inst = 32'h10408000;
      35420: inst = 32'hc404c5e;
      35421: inst = 32'h8220000;
      35422: inst = 32'h10408000;
      35423: inst = 32'hc404c5f;
      35424: inst = 32'h8220000;
      35425: inst = 32'h10408000;
      35426: inst = 32'hc404c60;
      35427: inst = 32'h8220000;
      35428: inst = 32'h10408000;
      35429: inst = 32'hc404c61;
      35430: inst = 32'h8220000;
      35431: inst = 32'h10408000;
      35432: inst = 32'hc404c62;
      35433: inst = 32'h8220000;
      35434: inst = 32'h10408000;
      35435: inst = 32'hc404c63;
      35436: inst = 32'h8220000;
      35437: inst = 32'h10408000;
      35438: inst = 32'hc404c64;
      35439: inst = 32'h8220000;
      35440: inst = 32'h10408000;
      35441: inst = 32'hc404c65;
      35442: inst = 32'h8220000;
      35443: inst = 32'h10408000;
      35444: inst = 32'hc404c66;
      35445: inst = 32'h8220000;
      35446: inst = 32'h10408000;
      35447: inst = 32'hc404c67;
      35448: inst = 32'h8220000;
      35449: inst = 32'h10408000;
      35450: inst = 32'hc404c68;
      35451: inst = 32'h8220000;
      35452: inst = 32'h10408000;
      35453: inst = 32'hc404c69;
      35454: inst = 32'h8220000;
      35455: inst = 32'h10408000;
      35456: inst = 32'hc404c6a;
      35457: inst = 32'h8220000;
      35458: inst = 32'h10408000;
      35459: inst = 32'hc404c6b;
      35460: inst = 32'h8220000;
      35461: inst = 32'h10408000;
      35462: inst = 32'hc404c6c;
      35463: inst = 32'h8220000;
      35464: inst = 32'h10408000;
      35465: inst = 32'hc404c6d;
      35466: inst = 32'h8220000;
      35467: inst = 32'h10408000;
      35468: inst = 32'hc404c6e;
      35469: inst = 32'h8220000;
      35470: inst = 32'h10408000;
      35471: inst = 32'hc404c6f;
      35472: inst = 32'h8220000;
      35473: inst = 32'h10408000;
      35474: inst = 32'hc404c70;
      35475: inst = 32'h8220000;
      35476: inst = 32'h10408000;
      35477: inst = 32'hc404c71;
      35478: inst = 32'h8220000;
      35479: inst = 32'h10408000;
      35480: inst = 32'hc404c72;
      35481: inst = 32'h8220000;
      35482: inst = 32'h10408000;
      35483: inst = 32'hc404c73;
      35484: inst = 32'h8220000;
      35485: inst = 32'h10408000;
      35486: inst = 32'hc404c74;
      35487: inst = 32'h8220000;
      35488: inst = 32'h10408000;
      35489: inst = 32'hc404c75;
      35490: inst = 32'h8220000;
      35491: inst = 32'h10408000;
      35492: inst = 32'hc404c76;
      35493: inst = 32'h8220000;
      35494: inst = 32'h10408000;
      35495: inst = 32'hc404c77;
      35496: inst = 32'h8220000;
      35497: inst = 32'h10408000;
      35498: inst = 32'hc404c78;
      35499: inst = 32'h8220000;
      35500: inst = 32'h10408000;
      35501: inst = 32'hc404c79;
      35502: inst = 32'h8220000;
      35503: inst = 32'h10408000;
      35504: inst = 32'hc404c7a;
      35505: inst = 32'h8220000;
      35506: inst = 32'h10408000;
      35507: inst = 32'hc404c7b;
      35508: inst = 32'h8220000;
      35509: inst = 32'h10408000;
      35510: inst = 32'hc404c7c;
      35511: inst = 32'h8220000;
      35512: inst = 32'h10408000;
      35513: inst = 32'hc404c7d;
      35514: inst = 32'h8220000;
      35515: inst = 32'h10408000;
      35516: inst = 32'hc404c7e;
      35517: inst = 32'h8220000;
      35518: inst = 32'h10408000;
      35519: inst = 32'hc404c7f;
      35520: inst = 32'h8220000;
      35521: inst = 32'h10408000;
      35522: inst = 32'hc404c80;
      35523: inst = 32'h8220000;
      35524: inst = 32'h10408000;
      35525: inst = 32'hc404c81;
      35526: inst = 32'h8220000;
      35527: inst = 32'h10408000;
      35528: inst = 32'hc404c82;
      35529: inst = 32'h8220000;
      35530: inst = 32'h10408000;
      35531: inst = 32'hc404c83;
      35532: inst = 32'h8220000;
      35533: inst = 32'h10408000;
      35534: inst = 32'hc404c84;
      35535: inst = 32'h8220000;
      35536: inst = 32'h10408000;
      35537: inst = 32'hc404c85;
      35538: inst = 32'h8220000;
      35539: inst = 32'h10408000;
      35540: inst = 32'hc404c86;
      35541: inst = 32'h8220000;
      35542: inst = 32'h10408000;
      35543: inst = 32'hc404c87;
      35544: inst = 32'h8220000;
      35545: inst = 32'h10408000;
      35546: inst = 32'hc404c88;
      35547: inst = 32'h8220000;
      35548: inst = 32'h10408000;
      35549: inst = 32'hc404c89;
      35550: inst = 32'h8220000;
      35551: inst = 32'h10408000;
      35552: inst = 32'hc404c8a;
      35553: inst = 32'h8220000;
      35554: inst = 32'h10408000;
      35555: inst = 32'hc404c8b;
      35556: inst = 32'h8220000;
      35557: inst = 32'h10408000;
      35558: inst = 32'hc404c8c;
      35559: inst = 32'h8220000;
      35560: inst = 32'h10408000;
      35561: inst = 32'hc404c8d;
      35562: inst = 32'h8220000;
      35563: inst = 32'h10408000;
      35564: inst = 32'hc404c8e;
      35565: inst = 32'h8220000;
      35566: inst = 32'h10408000;
      35567: inst = 32'hc404c8f;
      35568: inst = 32'h8220000;
      35569: inst = 32'h10408000;
      35570: inst = 32'hc404c90;
      35571: inst = 32'h8220000;
      35572: inst = 32'h10408000;
      35573: inst = 32'hc404c91;
      35574: inst = 32'h8220000;
      35575: inst = 32'h10408000;
      35576: inst = 32'hc404c92;
      35577: inst = 32'h8220000;
      35578: inst = 32'h10408000;
      35579: inst = 32'hc404c93;
      35580: inst = 32'h8220000;
      35581: inst = 32'h10408000;
      35582: inst = 32'hc404c94;
      35583: inst = 32'h8220000;
      35584: inst = 32'h10408000;
      35585: inst = 32'hc404c95;
      35586: inst = 32'h8220000;
      35587: inst = 32'h10408000;
      35588: inst = 32'hc404c96;
      35589: inst = 32'h8220000;
      35590: inst = 32'h10408000;
      35591: inst = 32'hc404c97;
      35592: inst = 32'h8220000;
      35593: inst = 32'h10408000;
      35594: inst = 32'hc404c98;
      35595: inst = 32'h8220000;
      35596: inst = 32'h10408000;
      35597: inst = 32'hc404c99;
      35598: inst = 32'h8220000;
      35599: inst = 32'h10408000;
      35600: inst = 32'hc404c9a;
      35601: inst = 32'h8220000;
      35602: inst = 32'h10408000;
      35603: inst = 32'hc404c9b;
      35604: inst = 32'h8220000;
      35605: inst = 32'h10408000;
      35606: inst = 32'hc404c9c;
      35607: inst = 32'h8220000;
      35608: inst = 32'h10408000;
      35609: inst = 32'hc404ca3;
      35610: inst = 32'h8220000;
      35611: inst = 32'h10408000;
      35612: inst = 32'hc404ca4;
      35613: inst = 32'h8220000;
      35614: inst = 32'h10408000;
      35615: inst = 32'hc404ca5;
      35616: inst = 32'h8220000;
      35617: inst = 32'h10408000;
      35618: inst = 32'hc404ca6;
      35619: inst = 32'h8220000;
      35620: inst = 32'h10408000;
      35621: inst = 32'hc404ca7;
      35622: inst = 32'h8220000;
      35623: inst = 32'h10408000;
      35624: inst = 32'hc404ca8;
      35625: inst = 32'h8220000;
      35626: inst = 32'h10408000;
      35627: inst = 32'hc404ca9;
      35628: inst = 32'h8220000;
      35629: inst = 32'h10408000;
      35630: inst = 32'hc404caa;
      35631: inst = 32'h8220000;
      35632: inst = 32'h10408000;
      35633: inst = 32'hc404cab;
      35634: inst = 32'h8220000;
      35635: inst = 32'h10408000;
      35636: inst = 32'hc404cac;
      35637: inst = 32'h8220000;
      35638: inst = 32'h10408000;
      35639: inst = 32'hc404cad;
      35640: inst = 32'h8220000;
      35641: inst = 32'h10408000;
      35642: inst = 32'hc404cae;
      35643: inst = 32'h8220000;
      35644: inst = 32'h10408000;
      35645: inst = 32'hc404caf;
      35646: inst = 32'h8220000;
      35647: inst = 32'h10408000;
      35648: inst = 32'hc404cb0;
      35649: inst = 32'h8220000;
      35650: inst = 32'h10408000;
      35651: inst = 32'hc404cb1;
      35652: inst = 32'h8220000;
      35653: inst = 32'h10408000;
      35654: inst = 32'hc404cb2;
      35655: inst = 32'h8220000;
      35656: inst = 32'h10408000;
      35657: inst = 32'hc404cb3;
      35658: inst = 32'h8220000;
      35659: inst = 32'h10408000;
      35660: inst = 32'hc404cb4;
      35661: inst = 32'h8220000;
      35662: inst = 32'h10408000;
      35663: inst = 32'hc404cb5;
      35664: inst = 32'h8220000;
      35665: inst = 32'h10408000;
      35666: inst = 32'hc404cb6;
      35667: inst = 32'h8220000;
      35668: inst = 32'h10408000;
      35669: inst = 32'hc404cb7;
      35670: inst = 32'h8220000;
      35671: inst = 32'h10408000;
      35672: inst = 32'hc404cb8;
      35673: inst = 32'h8220000;
      35674: inst = 32'h10408000;
      35675: inst = 32'hc404cb9;
      35676: inst = 32'h8220000;
      35677: inst = 32'h10408000;
      35678: inst = 32'hc404cba;
      35679: inst = 32'h8220000;
      35680: inst = 32'h10408000;
      35681: inst = 32'hc404cbb;
      35682: inst = 32'h8220000;
      35683: inst = 32'h10408000;
      35684: inst = 32'hc404cbc;
      35685: inst = 32'h8220000;
      35686: inst = 32'h10408000;
      35687: inst = 32'hc404cbd;
      35688: inst = 32'h8220000;
      35689: inst = 32'h10408000;
      35690: inst = 32'hc404cbe;
      35691: inst = 32'h8220000;
      35692: inst = 32'h10408000;
      35693: inst = 32'hc404cbf;
      35694: inst = 32'h8220000;
      35695: inst = 32'h10408000;
      35696: inst = 32'hc404cc0;
      35697: inst = 32'h8220000;
      35698: inst = 32'h10408000;
      35699: inst = 32'hc404cc1;
      35700: inst = 32'h8220000;
      35701: inst = 32'h10408000;
      35702: inst = 32'hc404cc2;
      35703: inst = 32'h8220000;
      35704: inst = 32'h10408000;
      35705: inst = 32'hc404cc3;
      35706: inst = 32'h8220000;
      35707: inst = 32'h10408000;
      35708: inst = 32'hc404cc4;
      35709: inst = 32'h8220000;
      35710: inst = 32'h10408000;
      35711: inst = 32'hc404cc5;
      35712: inst = 32'h8220000;
      35713: inst = 32'h10408000;
      35714: inst = 32'hc404cc6;
      35715: inst = 32'h8220000;
      35716: inst = 32'h10408000;
      35717: inst = 32'hc404cc7;
      35718: inst = 32'h8220000;
      35719: inst = 32'h10408000;
      35720: inst = 32'hc404cc8;
      35721: inst = 32'h8220000;
      35722: inst = 32'h10408000;
      35723: inst = 32'hc404cc9;
      35724: inst = 32'h8220000;
      35725: inst = 32'h10408000;
      35726: inst = 32'hc404cca;
      35727: inst = 32'h8220000;
      35728: inst = 32'h10408000;
      35729: inst = 32'hc404ccb;
      35730: inst = 32'h8220000;
      35731: inst = 32'h10408000;
      35732: inst = 32'hc404ccc;
      35733: inst = 32'h8220000;
      35734: inst = 32'h10408000;
      35735: inst = 32'hc404ccd;
      35736: inst = 32'h8220000;
      35737: inst = 32'h10408000;
      35738: inst = 32'hc404cce;
      35739: inst = 32'h8220000;
      35740: inst = 32'h10408000;
      35741: inst = 32'hc404ccf;
      35742: inst = 32'h8220000;
      35743: inst = 32'h10408000;
      35744: inst = 32'hc404cd0;
      35745: inst = 32'h8220000;
      35746: inst = 32'h10408000;
      35747: inst = 32'hc404cd1;
      35748: inst = 32'h8220000;
      35749: inst = 32'h10408000;
      35750: inst = 32'hc404cd2;
      35751: inst = 32'h8220000;
      35752: inst = 32'h10408000;
      35753: inst = 32'hc404cd3;
      35754: inst = 32'h8220000;
      35755: inst = 32'h10408000;
      35756: inst = 32'hc404cd4;
      35757: inst = 32'h8220000;
      35758: inst = 32'h10408000;
      35759: inst = 32'hc404cd5;
      35760: inst = 32'h8220000;
      35761: inst = 32'h10408000;
      35762: inst = 32'hc404cd6;
      35763: inst = 32'h8220000;
      35764: inst = 32'h10408000;
      35765: inst = 32'hc404cd7;
      35766: inst = 32'h8220000;
      35767: inst = 32'h10408000;
      35768: inst = 32'hc404cd8;
      35769: inst = 32'h8220000;
      35770: inst = 32'h10408000;
      35771: inst = 32'hc404cd9;
      35772: inst = 32'h8220000;
      35773: inst = 32'h10408000;
      35774: inst = 32'hc404cda;
      35775: inst = 32'h8220000;
      35776: inst = 32'h10408000;
      35777: inst = 32'hc404cdb;
      35778: inst = 32'h8220000;
      35779: inst = 32'h10408000;
      35780: inst = 32'hc404cdc;
      35781: inst = 32'h8220000;
      35782: inst = 32'h10408000;
      35783: inst = 32'hc404cdd;
      35784: inst = 32'h8220000;
      35785: inst = 32'h10408000;
      35786: inst = 32'hc404cde;
      35787: inst = 32'h8220000;
      35788: inst = 32'h10408000;
      35789: inst = 32'hc404cdf;
      35790: inst = 32'h8220000;
      35791: inst = 32'h10408000;
      35792: inst = 32'hc404ce0;
      35793: inst = 32'h8220000;
      35794: inst = 32'h10408000;
      35795: inst = 32'hc404ce1;
      35796: inst = 32'h8220000;
      35797: inst = 32'h10408000;
      35798: inst = 32'hc404ce2;
      35799: inst = 32'h8220000;
      35800: inst = 32'h10408000;
      35801: inst = 32'hc404ce3;
      35802: inst = 32'h8220000;
      35803: inst = 32'h10408000;
      35804: inst = 32'hc404ce4;
      35805: inst = 32'h8220000;
      35806: inst = 32'h10408000;
      35807: inst = 32'hc404ce5;
      35808: inst = 32'h8220000;
      35809: inst = 32'h10408000;
      35810: inst = 32'hc404ce6;
      35811: inst = 32'h8220000;
      35812: inst = 32'h10408000;
      35813: inst = 32'hc404ce7;
      35814: inst = 32'h8220000;
      35815: inst = 32'h10408000;
      35816: inst = 32'hc404ce8;
      35817: inst = 32'h8220000;
      35818: inst = 32'h10408000;
      35819: inst = 32'hc404ce9;
      35820: inst = 32'h8220000;
      35821: inst = 32'h10408000;
      35822: inst = 32'hc404cea;
      35823: inst = 32'h8220000;
      35824: inst = 32'h10408000;
      35825: inst = 32'hc404ceb;
      35826: inst = 32'h8220000;
      35827: inst = 32'h10408000;
      35828: inst = 32'hc404cec;
      35829: inst = 32'h8220000;
      35830: inst = 32'h10408000;
      35831: inst = 32'hc404ced;
      35832: inst = 32'h8220000;
      35833: inst = 32'h10408000;
      35834: inst = 32'hc404cee;
      35835: inst = 32'h8220000;
      35836: inst = 32'h10408000;
      35837: inst = 32'hc404cef;
      35838: inst = 32'h8220000;
      35839: inst = 32'h10408000;
      35840: inst = 32'hc404cf0;
      35841: inst = 32'h8220000;
      35842: inst = 32'h10408000;
      35843: inst = 32'hc404cf1;
      35844: inst = 32'h8220000;
      35845: inst = 32'h10408000;
      35846: inst = 32'hc404cf2;
      35847: inst = 32'h8220000;
      35848: inst = 32'h10408000;
      35849: inst = 32'hc404cf3;
      35850: inst = 32'h8220000;
      35851: inst = 32'h10408000;
      35852: inst = 32'hc404cf4;
      35853: inst = 32'h8220000;
      35854: inst = 32'h10408000;
      35855: inst = 32'hc404cf5;
      35856: inst = 32'h8220000;
      35857: inst = 32'h10408000;
      35858: inst = 32'hc404cf6;
      35859: inst = 32'h8220000;
      35860: inst = 32'h10408000;
      35861: inst = 32'hc404cf7;
      35862: inst = 32'h8220000;
      35863: inst = 32'h10408000;
      35864: inst = 32'hc404cf8;
      35865: inst = 32'h8220000;
      35866: inst = 32'h10408000;
      35867: inst = 32'hc404cf9;
      35868: inst = 32'h8220000;
      35869: inst = 32'h10408000;
      35870: inst = 32'hc404cfa;
      35871: inst = 32'h8220000;
      35872: inst = 32'h10408000;
      35873: inst = 32'hc404cfb;
      35874: inst = 32'h8220000;
      35875: inst = 32'h10408000;
      35876: inst = 32'hc404cfc;
      35877: inst = 32'h8220000;
      35878: inst = 32'h10408000;
      35879: inst = 32'hc404d03;
      35880: inst = 32'h8220000;
      35881: inst = 32'h10408000;
      35882: inst = 32'hc404d04;
      35883: inst = 32'h8220000;
      35884: inst = 32'h10408000;
      35885: inst = 32'hc404d05;
      35886: inst = 32'h8220000;
      35887: inst = 32'h10408000;
      35888: inst = 32'hc404d06;
      35889: inst = 32'h8220000;
      35890: inst = 32'h10408000;
      35891: inst = 32'hc404d07;
      35892: inst = 32'h8220000;
      35893: inst = 32'h10408000;
      35894: inst = 32'hc404d08;
      35895: inst = 32'h8220000;
      35896: inst = 32'h10408000;
      35897: inst = 32'hc404d09;
      35898: inst = 32'h8220000;
      35899: inst = 32'h10408000;
      35900: inst = 32'hc404d0a;
      35901: inst = 32'h8220000;
      35902: inst = 32'h10408000;
      35903: inst = 32'hc404d0b;
      35904: inst = 32'h8220000;
      35905: inst = 32'h10408000;
      35906: inst = 32'hc404d0c;
      35907: inst = 32'h8220000;
      35908: inst = 32'h10408000;
      35909: inst = 32'hc404d0d;
      35910: inst = 32'h8220000;
      35911: inst = 32'h10408000;
      35912: inst = 32'hc404d0e;
      35913: inst = 32'h8220000;
      35914: inst = 32'h10408000;
      35915: inst = 32'hc404d0f;
      35916: inst = 32'h8220000;
      35917: inst = 32'h10408000;
      35918: inst = 32'hc404d10;
      35919: inst = 32'h8220000;
      35920: inst = 32'h10408000;
      35921: inst = 32'hc404d11;
      35922: inst = 32'h8220000;
      35923: inst = 32'h10408000;
      35924: inst = 32'hc404d12;
      35925: inst = 32'h8220000;
      35926: inst = 32'h10408000;
      35927: inst = 32'hc404d13;
      35928: inst = 32'h8220000;
      35929: inst = 32'h10408000;
      35930: inst = 32'hc404d14;
      35931: inst = 32'h8220000;
      35932: inst = 32'h10408000;
      35933: inst = 32'hc404d15;
      35934: inst = 32'h8220000;
      35935: inst = 32'h10408000;
      35936: inst = 32'hc404d16;
      35937: inst = 32'h8220000;
      35938: inst = 32'h10408000;
      35939: inst = 32'hc404d17;
      35940: inst = 32'h8220000;
      35941: inst = 32'h10408000;
      35942: inst = 32'hc404d18;
      35943: inst = 32'h8220000;
      35944: inst = 32'h10408000;
      35945: inst = 32'hc404d19;
      35946: inst = 32'h8220000;
      35947: inst = 32'h10408000;
      35948: inst = 32'hc404d1a;
      35949: inst = 32'h8220000;
      35950: inst = 32'h10408000;
      35951: inst = 32'hc404d1b;
      35952: inst = 32'h8220000;
      35953: inst = 32'h10408000;
      35954: inst = 32'hc404d1c;
      35955: inst = 32'h8220000;
      35956: inst = 32'h10408000;
      35957: inst = 32'hc404d1d;
      35958: inst = 32'h8220000;
      35959: inst = 32'h10408000;
      35960: inst = 32'hc404d1e;
      35961: inst = 32'h8220000;
      35962: inst = 32'h10408000;
      35963: inst = 32'hc404d1f;
      35964: inst = 32'h8220000;
      35965: inst = 32'h10408000;
      35966: inst = 32'hc404d20;
      35967: inst = 32'h8220000;
      35968: inst = 32'h10408000;
      35969: inst = 32'hc404d21;
      35970: inst = 32'h8220000;
      35971: inst = 32'h10408000;
      35972: inst = 32'hc404d22;
      35973: inst = 32'h8220000;
      35974: inst = 32'h10408000;
      35975: inst = 32'hc404d23;
      35976: inst = 32'h8220000;
      35977: inst = 32'h10408000;
      35978: inst = 32'hc404d24;
      35979: inst = 32'h8220000;
      35980: inst = 32'h10408000;
      35981: inst = 32'hc404d3b;
      35982: inst = 32'h8220000;
      35983: inst = 32'h10408000;
      35984: inst = 32'hc404d3c;
      35985: inst = 32'h8220000;
      35986: inst = 32'h10408000;
      35987: inst = 32'hc404d3d;
      35988: inst = 32'h8220000;
      35989: inst = 32'h10408000;
      35990: inst = 32'hc404d3e;
      35991: inst = 32'h8220000;
      35992: inst = 32'h10408000;
      35993: inst = 32'hc404d3f;
      35994: inst = 32'h8220000;
      35995: inst = 32'h10408000;
      35996: inst = 32'hc404d40;
      35997: inst = 32'h8220000;
      35998: inst = 32'h10408000;
      35999: inst = 32'hc404d41;
      36000: inst = 32'h8220000;
      36001: inst = 32'h10408000;
      36002: inst = 32'hc404d42;
      36003: inst = 32'h8220000;
      36004: inst = 32'h10408000;
      36005: inst = 32'hc404d43;
      36006: inst = 32'h8220000;
      36007: inst = 32'h10408000;
      36008: inst = 32'hc404d44;
      36009: inst = 32'h8220000;
      36010: inst = 32'h10408000;
      36011: inst = 32'hc404d45;
      36012: inst = 32'h8220000;
      36013: inst = 32'h10408000;
      36014: inst = 32'hc404d46;
      36015: inst = 32'h8220000;
      36016: inst = 32'h10408000;
      36017: inst = 32'hc404d47;
      36018: inst = 32'h8220000;
      36019: inst = 32'h10408000;
      36020: inst = 32'hc404d48;
      36021: inst = 32'h8220000;
      36022: inst = 32'h10408000;
      36023: inst = 32'hc404d49;
      36024: inst = 32'h8220000;
      36025: inst = 32'h10408000;
      36026: inst = 32'hc404d4a;
      36027: inst = 32'h8220000;
      36028: inst = 32'h10408000;
      36029: inst = 32'hc404d4b;
      36030: inst = 32'h8220000;
      36031: inst = 32'h10408000;
      36032: inst = 32'hc404d4c;
      36033: inst = 32'h8220000;
      36034: inst = 32'h10408000;
      36035: inst = 32'hc404d4d;
      36036: inst = 32'h8220000;
      36037: inst = 32'h10408000;
      36038: inst = 32'hc404d4e;
      36039: inst = 32'h8220000;
      36040: inst = 32'h10408000;
      36041: inst = 32'hc404d4f;
      36042: inst = 32'h8220000;
      36043: inst = 32'h10408000;
      36044: inst = 32'hc404d50;
      36045: inst = 32'h8220000;
      36046: inst = 32'h10408000;
      36047: inst = 32'hc404d51;
      36048: inst = 32'h8220000;
      36049: inst = 32'h10408000;
      36050: inst = 32'hc404d52;
      36051: inst = 32'h8220000;
      36052: inst = 32'h10408000;
      36053: inst = 32'hc404d53;
      36054: inst = 32'h8220000;
      36055: inst = 32'h10408000;
      36056: inst = 32'hc404d54;
      36057: inst = 32'h8220000;
      36058: inst = 32'h10408000;
      36059: inst = 32'hc404d55;
      36060: inst = 32'h8220000;
      36061: inst = 32'h10408000;
      36062: inst = 32'hc404d56;
      36063: inst = 32'h8220000;
      36064: inst = 32'h10408000;
      36065: inst = 32'hc404d57;
      36066: inst = 32'h8220000;
      36067: inst = 32'h10408000;
      36068: inst = 32'hc404d58;
      36069: inst = 32'h8220000;
      36070: inst = 32'h10408000;
      36071: inst = 32'hc404d59;
      36072: inst = 32'h8220000;
      36073: inst = 32'h10408000;
      36074: inst = 32'hc404d5a;
      36075: inst = 32'h8220000;
      36076: inst = 32'h10408000;
      36077: inst = 32'hc404d5b;
      36078: inst = 32'h8220000;
      36079: inst = 32'h10408000;
      36080: inst = 32'hc404d5c;
      36081: inst = 32'h8220000;
      36082: inst = 32'h10408000;
      36083: inst = 32'hc404d63;
      36084: inst = 32'h8220000;
      36085: inst = 32'h10408000;
      36086: inst = 32'hc404d64;
      36087: inst = 32'h8220000;
      36088: inst = 32'h10408000;
      36089: inst = 32'hc404d65;
      36090: inst = 32'h8220000;
      36091: inst = 32'h10408000;
      36092: inst = 32'hc404d66;
      36093: inst = 32'h8220000;
      36094: inst = 32'h10408000;
      36095: inst = 32'hc404d67;
      36096: inst = 32'h8220000;
      36097: inst = 32'h10408000;
      36098: inst = 32'hc404d68;
      36099: inst = 32'h8220000;
      36100: inst = 32'h10408000;
      36101: inst = 32'hc404d69;
      36102: inst = 32'h8220000;
      36103: inst = 32'h10408000;
      36104: inst = 32'hc404d6a;
      36105: inst = 32'h8220000;
      36106: inst = 32'h10408000;
      36107: inst = 32'hc404d6b;
      36108: inst = 32'h8220000;
      36109: inst = 32'h10408000;
      36110: inst = 32'hc404d6c;
      36111: inst = 32'h8220000;
      36112: inst = 32'h10408000;
      36113: inst = 32'hc404d6d;
      36114: inst = 32'h8220000;
      36115: inst = 32'h10408000;
      36116: inst = 32'hc404d6e;
      36117: inst = 32'h8220000;
      36118: inst = 32'h10408000;
      36119: inst = 32'hc404d6f;
      36120: inst = 32'h8220000;
      36121: inst = 32'h10408000;
      36122: inst = 32'hc404d70;
      36123: inst = 32'h8220000;
      36124: inst = 32'h10408000;
      36125: inst = 32'hc404d71;
      36126: inst = 32'h8220000;
      36127: inst = 32'h10408000;
      36128: inst = 32'hc404d72;
      36129: inst = 32'h8220000;
      36130: inst = 32'h10408000;
      36131: inst = 32'hc404d73;
      36132: inst = 32'h8220000;
      36133: inst = 32'h10408000;
      36134: inst = 32'hc404d74;
      36135: inst = 32'h8220000;
      36136: inst = 32'h10408000;
      36137: inst = 32'hc404d75;
      36138: inst = 32'h8220000;
      36139: inst = 32'h10408000;
      36140: inst = 32'hc404d76;
      36141: inst = 32'h8220000;
      36142: inst = 32'h10408000;
      36143: inst = 32'hc404d77;
      36144: inst = 32'h8220000;
      36145: inst = 32'h10408000;
      36146: inst = 32'hc404d78;
      36147: inst = 32'h8220000;
      36148: inst = 32'h10408000;
      36149: inst = 32'hc404d79;
      36150: inst = 32'h8220000;
      36151: inst = 32'h10408000;
      36152: inst = 32'hc404d7a;
      36153: inst = 32'h8220000;
      36154: inst = 32'h10408000;
      36155: inst = 32'hc404d7b;
      36156: inst = 32'h8220000;
      36157: inst = 32'h10408000;
      36158: inst = 32'hc404d7c;
      36159: inst = 32'h8220000;
      36160: inst = 32'h10408000;
      36161: inst = 32'hc404d7d;
      36162: inst = 32'h8220000;
      36163: inst = 32'h10408000;
      36164: inst = 32'hc404d7e;
      36165: inst = 32'h8220000;
      36166: inst = 32'h10408000;
      36167: inst = 32'hc404d7f;
      36168: inst = 32'h8220000;
      36169: inst = 32'h10408000;
      36170: inst = 32'hc404d80;
      36171: inst = 32'h8220000;
      36172: inst = 32'h10408000;
      36173: inst = 32'hc404d81;
      36174: inst = 32'h8220000;
      36175: inst = 32'h10408000;
      36176: inst = 32'hc404d82;
      36177: inst = 32'h8220000;
      36178: inst = 32'h10408000;
      36179: inst = 32'hc404d83;
      36180: inst = 32'h8220000;
      36181: inst = 32'h10408000;
      36182: inst = 32'hc404d84;
      36183: inst = 32'h8220000;
      36184: inst = 32'h10408000;
      36185: inst = 32'hc404d9b;
      36186: inst = 32'h8220000;
      36187: inst = 32'h10408000;
      36188: inst = 32'hc404d9c;
      36189: inst = 32'h8220000;
      36190: inst = 32'h10408000;
      36191: inst = 32'hc404d9d;
      36192: inst = 32'h8220000;
      36193: inst = 32'h10408000;
      36194: inst = 32'hc404d9e;
      36195: inst = 32'h8220000;
      36196: inst = 32'h10408000;
      36197: inst = 32'hc404d9f;
      36198: inst = 32'h8220000;
      36199: inst = 32'h10408000;
      36200: inst = 32'hc404da0;
      36201: inst = 32'h8220000;
      36202: inst = 32'h10408000;
      36203: inst = 32'hc404da1;
      36204: inst = 32'h8220000;
      36205: inst = 32'h10408000;
      36206: inst = 32'hc404da2;
      36207: inst = 32'h8220000;
      36208: inst = 32'h10408000;
      36209: inst = 32'hc404da3;
      36210: inst = 32'h8220000;
      36211: inst = 32'h10408000;
      36212: inst = 32'hc404da4;
      36213: inst = 32'h8220000;
      36214: inst = 32'h10408000;
      36215: inst = 32'hc404da5;
      36216: inst = 32'h8220000;
      36217: inst = 32'h10408000;
      36218: inst = 32'hc404da6;
      36219: inst = 32'h8220000;
      36220: inst = 32'h10408000;
      36221: inst = 32'hc404da7;
      36222: inst = 32'h8220000;
      36223: inst = 32'h10408000;
      36224: inst = 32'hc404da8;
      36225: inst = 32'h8220000;
      36226: inst = 32'h10408000;
      36227: inst = 32'hc404da9;
      36228: inst = 32'h8220000;
      36229: inst = 32'h10408000;
      36230: inst = 32'hc404daa;
      36231: inst = 32'h8220000;
      36232: inst = 32'h10408000;
      36233: inst = 32'hc404dab;
      36234: inst = 32'h8220000;
      36235: inst = 32'h10408000;
      36236: inst = 32'hc404dac;
      36237: inst = 32'h8220000;
      36238: inst = 32'h10408000;
      36239: inst = 32'hc404dad;
      36240: inst = 32'h8220000;
      36241: inst = 32'h10408000;
      36242: inst = 32'hc404dae;
      36243: inst = 32'h8220000;
      36244: inst = 32'h10408000;
      36245: inst = 32'hc404daf;
      36246: inst = 32'h8220000;
      36247: inst = 32'h10408000;
      36248: inst = 32'hc404db0;
      36249: inst = 32'h8220000;
      36250: inst = 32'h10408000;
      36251: inst = 32'hc404db1;
      36252: inst = 32'h8220000;
      36253: inst = 32'h10408000;
      36254: inst = 32'hc404db2;
      36255: inst = 32'h8220000;
      36256: inst = 32'h10408000;
      36257: inst = 32'hc404db3;
      36258: inst = 32'h8220000;
      36259: inst = 32'h10408000;
      36260: inst = 32'hc404db4;
      36261: inst = 32'h8220000;
      36262: inst = 32'h10408000;
      36263: inst = 32'hc404db5;
      36264: inst = 32'h8220000;
      36265: inst = 32'h10408000;
      36266: inst = 32'hc404db6;
      36267: inst = 32'h8220000;
      36268: inst = 32'h10408000;
      36269: inst = 32'hc404db7;
      36270: inst = 32'h8220000;
      36271: inst = 32'h10408000;
      36272: inst = 32'hc404db8;
      36273: inst = 32'h8220000;
      36274: inst = 32'h10408000;
      36275: inst = 32'hc404db9;
      36276: inst = 32'h8220000;
      36277: inst = 32'h10408000;
      36278: inst = 32'hc404dba;
      36279: inst = 32'h8220000;
      36280: inst = 32'h10408000;
      36281: inst = 32'hc404dbb;
      36282: inst = 32'h8220000;
      36283: inst = 32'h10408000;
      36284: inst = 32'hc404dbc;
      36285: inst = 32'h8220000;
      36286: inst = 32'h10408000;
      36287: inst = 32'hc404dc3;
      36288: inst = 32'h8220000;
      36289: inst = 32'h10408000;
      36290: inst = 32'hc404dc4;
      36291: inst = 32'h8220000;
      36292: inst = 32'h10408000;
      36293: inst = 32'hc404dc5;
      36294: inst = 32'h8220000;
      36295: inst = 32'h10408000;
      36296: inst = 32'hc404dc6;
      36297: inst = 32'h8220000;
      36298: inst = 32'h10408000;
      36299: inst = 32'hc404dc7;
      36300: inst = 32'h8220000;
      36301: inst = 32'h10408000;
      36302: inst = 32'hc404dc8;
      36303: inst = 32'h8220000;
      36304: inst = 32'h10408000;
      36305: inst = 32'hc404dc9;
      36306: inst = 32'h8220000;
      36307: inst = 32'h10408000;
      36308: inst = 32'hc404dca;
      36309: inst = 32'h8220000;
      36310: inst = 32'h10408000;
      36311: inst = 32'hc404dcb;
      36312: inst = 32'h8220000;
      36313: inst = 32'h10408000;
      36314: inst = 32'hc404dcc;
      36315: inst = 32'h8220000;
      36316: inst = 32'h10408000;
      36317: inst = 32'hc404dcd;
      36318: inst = 32'h8220000;
      36319: inst = 32'h10408000;
      36320: inst = 32'hc404dce;
      36321: inst = 32'h8220000;
      36322: inst = 32'h10408000;
      36323: inst = 32'hc404dcf;
      36324: inst = 32'h8220000;
      36325: inst = 32'h10408000;
      36326: inst = 32'hc404dd0;
      36327: inst = 32'h8220000;
      36328: inst = 32'h10408000;
      36329: inst = 32'hc404dd1;
      36330: inst = 32'h8220000;
      36331: inst = 32'h10408000;
      36332: inst = 32'hc404dd2;
      36333: inst = 32'h8220000;
      36334: inst = 32'h10408000;
      36335: inst = 32'hc404dd3;
      36336: inst = 32'h8220000;
      36337: inst = 32'h10408000;
      36338: inst = 32'hc404dd4;
      36339: inst = 32'h8220000;
      36340: inst = 32'h10408000;
      36341: inst = 32'hc404dd5;
      36342: inst = 32'h8220000;
      36343: inst = 32'h10408000;
      36344: inst = 32'hc404dd6;
      36345: inst = 32'h8220000;
      36346: inst = 32'h10408000;
      36347: inst = 32'hc404dd7;
      36348: inst = 32'h8220000;
      36349: inst = 32'h10408000;
      36350: inst = 32'hc404dd8;
      36351: inst = 32'h8220000;
      36352: inst = 32'h10408000;
      36353: inst = 32'hc404dd9;
      36354: inst = 32'h8220000;
      36355: inst = 32'h10408000;
      36356: inst = 32'hc404dda;
      36357: inst = 32'h8220000;
      36358: inst = 32'h10408000;
      36359: inst = 32'hc404ddb;
      36360: inst = 32'h8220000;
      36361: inst = 32'h10408000;
      36362: inst = 32'hc404ddc;
      36363: inst = 32'h8220000;
      36364: inst = 32'h10408000;
      36365: inst = 32'hc404ddd;
      36366: inst = 32'h8220000;
      36367: inst = 32'h10408000;
      36368: inst = 32'hc404dde;
      36369: inst = 32'h8220000;
      36370: inst = 32'h10408000;
      36371: inst = 32'hc404ddf;
      36372: inst = 32'h8220000;
      36373: inst = 32'h10408000;
      36374: inst = 32'hc404de0;
      36375: inst = 32'h8220000;
      36376: inst = 32'h10408000;
      36377: inst = 32'hc404de1;
      36378: inst = 32'h8220000;
      36379: inst = 32'h10408000;
      36380: inst = 32'hc404de2;
      36381: inst = 32'h8220000;
      36382: inst = 32'h10408000;
      36383: inst = 32'hc404de3;
      36384: inst = 32'h8220000;
      36385: inst = 32'h10408000;
      36386: inst = 32'hc404de4;
      36387: inst = 32'h8220000;
      36388: inst = 32'h10408000;
      36389: inst = 32'hc404dfb;
      36390: inst = 32'h8220000;
      36391: inst = 32'h10408000;
      36392: inst = 32'hc404dfc;
      36393: inst = 32'h8220000;
      36394: inst = 32'h10408000;
      36395: inst = 32'hc404dfd;
      36396: inst = 32'h8220000;
      36397: inst = 32'h10408000;
      36398: inst = 32'hc404dfe;
      36399: inst = 32'h8220000;
      36400: inst = 32'h10408000;
      36401: inst = 32'hc404dff;
      36402: inst = 32'h8220000;
      36403: inst = 32'h10408000;
      36404: inst = 32'hc404e00;
      36405: inst = 32'h8220000;
      36406: inst = 32'h10408000;
      36407: inst = 32'hc404e01;
      36408: inst = 32'h8220000;
      36409: inst = 32'h10408000;
      36410: inst = 32'hc404e02;
      36411: inst = 32'h8220000;
      36412: inst = 32'h10408000;
      36413: inst = 32'hc404e03;
      36414: inst = 32'h8220000;
      36415: inst = 32'h10408000;
      36416: inst = 32'hc404e04;
      36417: inst = 32'h8220000;
      36418: inst = 32'h10408000;
      36419: inst = 32'hc404e05;
      36420: inst = 32'h8220000;
      36421: inst = 32'h10408000;
      36422: inst = 32'hc404e06;
      36423: inst = 32'h8220000;
      36424: inst = 32'h10408000;
      36425: inst = 32'hc404e07;
      36426: inst = 32'h8220000;
      36427: inst = 32'h10408000;
      36428: inst = 32'hc404e08;
      36429: inst = 32'h8220000;
      36430: inst = 32'h10408000;
      36431: inst = 32'hc404e09;
      36432: inst = 32'h8220000;
      36433: inst = 32'h10408000;
      36434: inst = 32'hc404e0a;
      36435: inst = 32'h8220000;
      36436: inst = 32'h10408000;
      36437: inst = 32'hc404e0b;
      36438: inst = 32'h8220000;
      36439: inst = 32'h10408000;
      36440: inst = 32'hc404e0c;
      36441: inst = 32'h8220000;
      36442: inst = 32'h10408000;
      36443: inst = 32'hc404e0d;
      36444: inst = 32'h8220000;
      36445: inst = 32'h10408000;
      36446: inst = 32'hc404e0e;
      36447: inst = 32'h8220000;
      36448: inst = 32'h10408000;
      36449: inst = 32'hc404e0f;
      36450: inst = 32'h8220000;
      36451: inst = 32'h10408000;
      36452: inst = 32'hc404e10;
      36453: inst = 32'h8220000;
      36454: inst = 32'h10408000;
      36455: inst = 32'hc404e11;
      36456: inst = 32'h8220000;
      36457: inst = 32'h10408000;
      36458: inst = 32'hc404e12;
      36459: inst = 32'h8220000;
      36460: inst = 32'h10408000;
      36461: inst = 32'hc404e13;
      36462: inst = 32'h8220000;
      36463: inst = 32'h10408000;
      36464: inst = 32'hc404e14;
      36465: inst = 32'h8220000;
      36466: inst = 32'h10408000;
      36467: inst = 32'hc404e15;
      36468: inst = 32'h8220000;
      36469: inst = 32'h10408000;
      36470: inst = 32'hc404e16;
      36471: inst = 32'h8220000;
      36472: inst = 32'h10408000;
      36473: inst = 32'hc404e17;
      36474: inst = 32'h8220000;
      36475: inst = 32'h10408000;
      36476: inst = 32'hc404e18;
      36477: inst = 32'h8220000;
      36478: inst = 32'h10408000;
      36479: inst = 32'hc404e19;
      36480: inst = 32'h8220000;
      36481: inst = 32'h10408000;
      36482: inst = 32'hc404e1a;
      36483: inst = 32'h8220000;
      36484: inst = 32'h10408000;
      36485: inst = 32'hc404e1b;
      36486: inst = 32'h8220000;
      36487: inst = 32'h10408000;
      36488: inst = 32'hc404e1c;
      36489: inst = 32'h8220000;
      36490: inst = 32'h10408000;
      36491: inst = 32'hc404e23;
      36492: inst = 32'h8220000;
      36493: inst = 32'h10408000;
      36494: inst = 32'hc404e24;
      36495: inst = 32'h8220000;
      36496: inst = 32'h10408000;
      36497: inst = 32'hc404e25;
      36498: inst = 32'h8220000;
      36499: inst = 32'h10408000;
      36500: inst = 32'hc404e26;
      36501: inst = 32'h8220000;
      36502: inst = 32'h10408000;
      36503: inst = 32'hc404e27;
      36504: inst = 32'h8220000;
      36505: inst = 32'h10408000;
      36506: inst = 32'hc404e28;
      36507: inst = 32'h8220000;
      36508: inst = 32'h10408000;
      36509: inst = 32'hc404e29;
      36510: inst = 32'h8220000;
      36511: inst = 32'h10408000;
      36512: inst = 32'hc404e2a;
      36513: inst = 32'h8220000;
      36514: inst = 32'h10408000;
      36515: inst = 32'hc404e2b;
      36516: inst = 32'h8220000;
      36517: inst = 32'h10408000;
      36518: inst = 32'hc404e2c;
      36519: inst = 32'h8220000;
      36520: inst = 32'h10408000;
      36521: inst = 32'hc404e2d;
      36522: inst = 32'h8220000;
      36523: inst = 32'h10408000;
      36524: inst = 32'hc404e2e;
      36525: inst = 32'h8220000;
      36526: inst = 32'h10408000;
      36527: inst = 32'hc404e2f;
      36528: inst = 32'h8220000;
      36529: inst = 32'h10408000;
      36530: inst = 32'hc404e30;
      36531: inst = 32'h8220000;
      36532: inst = 32'h10408000;
      36533: inst = 32'hc404e31;
      36534: inst = 32'h8220000;
      36535: inst = 32'h10408000;
      36536: inst = 32'hc404e32;
      36537: inst = 32'h8220000;
      36538: inst = 32'h10408000;
      36539: inst = 32'hc404e33;
      36540: inst = 32'h8220000;
      36541: inst = 32'h10408000;
      36542: inst = 32'hc404e34;
      36543: inst = 32'h8220000;
      36544: inst = 32'h10408000;
      36545: inst = 32'hc404e35;
      36546: inst = 32'h8220000;
      36547: inst = 32'h10408000;
      36548: inst = 32'hc404e36;
      36549: inst = 32'h8220000;
      36550: inst = 32'h10408000;
      36551: inst = 32'hc404e37;
      36552: inst = 32'h8220000;
      36553: inst = 32'h10408000;
      36554: inst = 32'hc404e38;
      36555: inst = 32'h8220000;
      36556: inst = 32'h10408000;
      36557: inst = 32'hc404e39;
      36558: inst = 32'h8220000;
      36559: inst = 32'h10408000;
      36560: inst = 32'hc404e3a;
      36561: inst = 32'h8220000;
      36562: inst = 32'h10408000;
      36563: inst = 32'hc404e3b;
      36564: inst = 32'h8220000;
      36565: inst = 32'h10408000;
      36566: inst = 32'hc404e3c;
      36567: inst = 32'h8220000;
      36568: inst = 32'h10408000;
      36569: inst = 32'hc404e3d;
      36570: inst = 32'h8220000;
      36571: inst = 32'h10408000;
      36572: inst = 32'hc404e3e;
      36573: inst = 32'h8220000;
      36574: inst = 32'h10408000;
      36575: inst = 32'hc404e3f;
      36576: inst = 32'h8220000;
      36577: inst = 32'h10408000;
      36578: inst = 32'hc404e40;
      36579: inst = 32'h8220000;
      36580: inst = 32'h10408000;
      36581: inst = 32'hc404e41;
      36582: inst = 32'h8220000;
      36583: inst = 32'h10408000;
      36584: inst = 32'hc404e42;
      36585: inst = 32'h8220000;
      36586: inst = 32'h10408000;
      36587: inst = 32'hc404e43;
      36588: inst = 32'h8220000;
      36589: inst = 32'h10408000;
      36590: inst = 32'hc404e44;
      36591: inst = 32'h8220000;
      36592: inst = 32'h10408000;
      36593: inst = 32'hc404e45;
      36594: inst = 32'h8220000;
      36595: inst = 32'h10408000;
      36596: inst = 32'hc404e46;
      36597: inst = 32'h8220000;
      36598: inst = 32'h10408000;
      36599: inst = 32'hc404e47;
      36600: inst = 32'h8220000;
      36601: inst = 32'h10408000;
      36602: inst = 32'hc404e48;
      36603: inst = 32'h8220000;
      36604: inst = 32'h10408000;
      36605: inst = 32'hc404e49;
      36606: inst = 32'h8220000;
      36607: inst = 32'h10408000;
      36608: inst = 32'hc404e4a;
      36609: inst = 32'h8220000;
      36610: inst = 32'h10408000;
      36611: inst = 32'hc404e4b;
      36612: inst = 32'h8220000;
      36613: inst = 32'h10408000;
      36614: inst = 32'hc404e4c;
      36615: inst = 32'h8220000;
      36616: inst = 32'h10408000;
      36617: inst = 32'hc404e4d;
      36618: inst = 32'h8220000;
      36619: inst = 32'h10408000;
      36620: inst = 32'hc404e4e;
      36621: inst = 32'h8220000;
      36622: inst = 32'h10408000;
      36623: inst = 32'hc404e4f;
      36624: inst = 32'h8220000;
      36625: inst = 32'h10408000;
      36626: inst = 32'hc404e50;
      36627: inst = 32'h8220000;
      36628: inst = 32'h10408000;
      36629: inst = 32'hc404e51;
      36630: inst = 32'h8220000;
      36631: inst = 32'h10408000;
      36632: inst = 32'hc404e52;
      36633: inst = 32'h8220000;
      36634: inst = 32'h10408000;
      36635: inst = 32'hc404e53;
      36636: inst = 32'h8220000;
      36637: inst = 32'h10408000;
      36638: inst = 32'hc404e54;
      36639: inst = 32'h8220000;
      36640: inst = 32'h10408000;
      36641: inst = 32'hc404e55;
      36642: inst = 32'h8220000;
      36643: inst = 32'h10408000;
      36644: inst = 32'hc404e56;
      36645: inst = 32'h8220000;
      36646: inst = 32'h10408000;
      36647: inst = 32'hc404e57;
      36648: inst = 32'h8220000;
      36649: inst = 32'h10408000;
      36650: inst = 32'hc404e5b;
      36651: inst = 32'h8220000;
      36652: inst = 32'h10408000;
      36653: inst = 32'hc404e5c;
      36654: inst = 32'h8220000;
      36655: inst = 32'h10408000;
      36656: inst = 32'hc404e5d;
      36657: inst = 32'h8220000;
      36658: inst = 32'h10408000;
      36659: inst = 32'hc404e5e;
      36660: inst = 32'h8220000;
      36661: inst = 32'h10408000;
      36662: inst = 32'hc404e5f;
      36663: inst = 32'h8220000;
      36664: inst = 32'h10408000;
      36665: inst = 32'hc404e60;
      36666: inst = 32'h8220000;
      36667: inst = 32'h10408000;
      36668: inst = 32'hc404e61;
      36669: inst = 32'h8220000;
      36670: inst = 32'h10408000;
      36671: inst = 32'hc404e62;
      36672: inst = 32'h8220000;
      36673: inst = 32'h10408000;
      36674: inst = 32'hc404e63;
      36675: inst = 32'h8220000;
      36676: inst = 32'h10408000;
      36677: inst = 32'hc404e64;
      36678: inst = 32'h8220000;
      36679: inst = 32'h10408000;
      36680: inst = 32'hc404e65;
      36681: inst = 32'h8220000;
      36682: inst = 32'h10408000;
      36683: inst = 32'hc404e66;
      36684: inst = 32'h8220000;
      36685: inst = 32'h10408000;
      36686: inst = 32'hc404e67;
      36687: inst = 32'h8220000;
      36688: inst = 32'h10408000;
      36689: inst = 32'hc404e68;
      36690: inst = 32'h8220000;
      36691: inst = 32'h10408000;
      36692: inst = 32'hc404e69;
      36693: inst = 32'h8220000;
      36694: inst = 32'h10408000;
      36695: inst = 32'hc404e6a;
      36696: inst = 32'h8220000;
      36697: inst = 32'h10408000;
      36698: inst = 32'hc404e6b;
      36699: inst = 32'h8220000;
      36700: inst = 32'h10408000;
      36701: inst = 32'hc404e6c;
      36702: inst = 32'h8220000;
      36703: inst = 32'h10408000;
      36704: inst = 32'hc404e6d;
      36705: inst = 32'h8220000;
      36706: inst = 32'h10408000;
      36707: inst = 32'hc404e6e;
      36708: inst = 32'h8220000;
      36709: inst = 32'h10408000;
      36710: inst = 32'hc404e6f;
      36711: inst = 32'h8220000;
      36712: inst = 32'h10408000;
      36713: inst = 32'hc404e70;
      36714: inst = 32'h8220000;
      36715: inst = 32'h10408000;
      36716: inst = 32'hc404e71;
      36717: inst = 32'h8220000;
      36718: inst = 32'h10408000;
      36719: inst = 32'hc404e72;
      36720: inst = 32'h8220000;
      36721: inst = 32'h10408000;
      36722: inst = 32'hc404e73;
      36723: inst = 32'h8220000;
      36724: inst = 32'h10408000;
      36725: inst = 32'hc404e74;
      36726: inst = 32'h8220000;
      36727: inst = 32'h10408000;
      36728: inst = 32'hc404e75;
      36729: inst = 32'h8220000;
      36730: inst = 32'h10408000;
      36731: inst = 32'hc404e76;
      36732: inst = 32'h8220000;
      36733: inst = 32'h10408000;
      36734: inst = 32'hc404e77;
      36735: inst = 32'h8220000;
      36736: inst = 32'h10408000;
      36737: inst = 32'hc404e78;
      36738: inst = 32'h8220000;
      36739: inst = 32'h10408000;
      36740: inst = 32'hc404e79;
      36741: inst = 32'h8220000;
      36742: inst = 32'h10408000;
      36743: inst = 32'hc404e7a;
      36744: inst = 32'h8220000;
      36745: inst = 32'h10408000;
      36746: inst = 32'hc404e7b;
      36747: inst = 32'h8220000;
      36748: inst = 32'h10408000;
      36749: inst = 32'hc404e7c;
      36750: inst = 32'h8220000;
      36751: inst = 32'h10408000;
      36752: inst = 32'hc404e83;
      36753: inst = 32'h8220000;
      36754: inst = 32'h10408000;
      36755: inst = 32'hc404e84;
      36756: inst = 32'h8220000;
      36757: inst = 32'h10408000;
      36758: inst = 32'hc404e85;
      36759: inst = 32'h8220000;
      36760: inst = 32'h10408000;
      36761: inst = 32'hc404e86;
      36762: inst = 32'h8220000;
      36763: inst = 32'h10408000;
      36764: inst = 32'hc404e87;
      36765: inst = 32'h8220000;
      36766: inst = 32'h10408000;
      36767: inst = 32'hc404e88;
      36768: inst = 32'h8220000;
      36769: inst = 32'h10408000;
      36770: inst = 32'hc404e89;
      36771: inst = 32'h8220000;
      36772: inst = 32'h10408000;
      36773: inst = 32'hc404e8a;
      36774: inst = 32'h8220000;
      36775: inst = 32'h10408000;
      36776: inst = 32'hc404e8b;
      36777: inst = 32'h8220000;
      36778: inst = 32'h10408000;
      36779: inst = 32'hc404e8c;
      36780: inst = 32'h8220000;
      36781: inst = 32'h10408000;
      36782: inst = 32'hc404e8d;
      36783: inst = 32'h8220000;
      36784: inst = 32'h10408000;
      36785: inst = 32'hc404e8e;
      36786: inst = 32'h8220000;
      36787: inst = 32'h10408000;
      36788: inst = 32'hc404e8f;
      36789: inst = 32'h8220000;
      36790: inst = 32'h10408000;
      36791: inst = 32'hc404e90;
      36792: inst = 32'h8220000;
      36793: inst = 32'h10408000;
      36794: inst = 32'hc404e91;
      36795: inst = 32'h8220000;
      36796: inst = 32'h10408000;
      36797: inst = 32'hc404e92;
      36798: inst = 32'h8220000;
      36799: inst = 32'h10408000;
      36800: inst = 32'hc404e93;
      36801: inst = 32'h8220000;
      36802: inst = 32'h10408000;
      36803: inst = 32'hc404e94;
      36804: inst = 32'h8220000;
      36805: inst = 32'h10408000;
      36806: inst = 32'hc404e95;
      36807: inst = 32'h8220000;
      36808: inst = 32'h10408000;
      36809: inst = 32'hc404e96;
      36810: inst = 32'h8220000;
      36811: inst = 32'h10408000;
      36812: inst = 32'hc404e97;
      36813: inst = 32'h8220000;
      36814: inst = 32'h10408000;
      36815: inst = 32'hc404e98;
      36816: inst = 32'h8220000;
      36817: inst = 32'h10408000;
      36818: inst = 32'hc404e99;
      36819: inst = 32'h8220000;
      36820: inst = 32'h10408000;
      36821: inst = 32'hc404e9a;
      36822: inst = 32'h8220000;
      36823: inst = 32'h10408000;
      36824: inst = 32'hc404e9b;
      36825: inst = 32'h8220000;
      36826: inst = 32'h10408000;
      36827: inst = 32'hc404e9c;
      36828: inst = 32'h8220000;
      36829: inst = 32'h10408000;
      36830: inst = 32'hc404e9d;
      36831: inst = 32'h8220000;
      36832: inst = 32'h10408000;
      36833: inst = 32'hc404e9e;
      36834: inst = 32'h8220000;
      36835: inst = 32'h10408000;
      36836: inst = 32'hc404e9f;
      36837: inst = 32'h8220000;
      36838: inst = 32'h10408000;
      36839: inst = 32'hc404ea0;
      36840: inst = 32'h8220000;
      36841: inst = 32'h10408000;
      36842: inst = 32'hc404ea1;
      36843: inst = 32'h8220000;
      36844: inst = 32'h10408000;
      36845: inst = 32'hc404ea2;
      36846: inst = 32'h8220000;
      36847: inst = 32'h10408000;
      36848: inst = 32'hc404ea3;
      36849: inst = 32'h8220000;
      36850: inst = 32'h10408000;
      36851: inst = 32'hc404ea4;
      36852: inst = 32'h8220000;
      36853: inst = 32'h10408000;
      36854: inst = 32'hc404ea5;
      36855: inst = 32'h8220000;
      36856: inst = 32'h10408000;
      36857: inst = 32'hc404ea6;
      36858: inst = 32'h8220000;
      36859: inst = 32'h10408000;
      36860: inst = 32'hc404ea7;
      36861: inst = 32'h8220000;
      36862: inst = 32'h10408000;
      36863: inst = 32'hc404ea8;
      36864: inst = 32'h8220000;
      36865: inst = 32'h10408000;
      36866: inst = 32'hc404ea9;
      36867: inst = 32'h8220000;
      36868: inst = 32'h10408000;
      36869: inst = 32'hc404eaa;
      36870: inst = 32'h8220000;
      36871: inst = 32'h10408000;
      36872: inst = 32'hc404eab;
      36873: inst = 32'h8220000;
      36874: inst = 32'h10408000;
      36875: inst = 32'hc404eac;
      36876: inst = 32'h8220000;
      36877: inst = 32'h10408000;
      36878: inst = 32'hc404ead;
      36879: inst = 32'h8220000;
      36880: inst = 32'h10408000;
      36881: inst = 32'hc404eae;
      36882: inst = 32'h8220000;
      36883: inst = 32'h10408000;
      36884: inst = 32'hc404eaf;
      36885: inst = 32'h8220000;
      36886: inst = 32'h10408000;
      36887: inst = 32'hc404eb0;
      36888: inst = 32'h8220000;
      36889: inst = 32'h10408000;
      36890: inst = 32'hc404eb1;
      36891: inst = 32'h8220000;
      36892: inst = 32'h10408000;
      36893: inst = 32'hc404eb2;
      36894: inst = 32'h8220000;
      36895: inst = 32'h10408000;
      36896: inst = 32'hc404eb3;
      36897: inst = 32'h8220000;
      36898: inst = 32'h10408000;
      36899: inst = 32'hc404eb4;
      36900: inst = 32'h8220000;
      36901: inst = 32'h10408000;
      36902: inst = 32'hc404eb5;
      36903: inst = 32'h8220000;
      36904: inst = 32'h10408000;
      36905: inst = 32'hc404eb6;
      36906: inst = 32'h8220000;
      36907: inst = 32'h10408000;
      36908: inst = 32'hc404eb7;
      36909: inst = 32'h8220000;
      36910: inst = 32'h10408000;
      36911: inst = 32'hc404ebb;
      36912: inst = 32'h8220000;
      36913: inst = 32'h10408000;
      36914: inst = 32'hc404ebc;
      36915: inst = 32'h8220000;
      36916: inst = 32'h10408000;
      36917: inst = 32'hc404ebd;
      36918: inst = 32'h8220000;
      36919: inst = 32'h10408000;
      36920: inst = 32'hc404ebe;
      36921: inst = 32'h8220000;
      36922: inst = 32'h10408000;
      36923: inst = 32'hc404ebf;
      36924: inst = 32'h8220000;
      36925: inst = 32'h10408000;
      36926: inst = 32'hc404ec0;
      36927: inst = 32'h8220000;
      36928: inst = 32'h10408000;
      36929: inst = 32'hc404ec1;
      36930: inst = 32'h8220000;
      36931: inst = 32'h10408000;
      36932: inst = 32'hc404ec2;
      36933: inst = 32'h8220000;
      36934: inst = 32'h10408000;
      36935: inst = 32'hc404ec3;
      36936: inst = 32'h8220000;
      36937: inst = 32'h10408000;
      36938: inst = 32'hc404ec4;
      36939: inst = 32'h8220000;
      36940: inst = 32'h10408000;
      36941: inst = 32'hc404ec5;
      36942: inst = 32'h8220000;
      36943: inst = 32'h10408000;
      36944: inst = 32'hc404ec6;
      36945: inst = 32'h8220000;
      36946: inst = 32'h10408000;
      36947: inst = 32'hc404ec7;
      36948: inst = 32'h8220000;
      36949: inst = 32'h10408000;
      36950: inst = 32'hc404ec8;
      36951: inst = 32'h8220000;
      36952: inst = 32'h10408000;
      36953: inst = 32'hc404ec9;
      36954: inst = 32'h8220000;
      36955: inst = 32'h10408000;
      36956: inst = 32'hc404eca;
      36957: inst = 32'h8220000;
      36958: inst = 32'h10408000;
      36959: inst = 32'hc404ecb;
      36960: inst = 32'h8220000;
      36961: inst = 32'h10408000;
      36962: inst = 32'hc404ecc;
      36963: inst = 32'h8220000;
      36964: inst = 32'h10408000;
      36965: inst = 32'hc404ecd;
      36966: inst = 32'h8220000;
      36967: inst = 32'h10408000;
      36968: inst = 32'hc404ece;
      36969: inst = 32'h8220000;
      36970: inst = 32'h10408000;
      36971: inst = 32'hc404ecf;
      36972: inst = 32'h8220000;
      36973: inst = 32'h10408000;
      36974: inst = 32'hc404ed0;
      36975: inst = 32'h8220000;
      36976: inst = 32'h10408000;
      36977: inst = 32'hc404ed1;
      36978: inst = 32'h8220000;
      36979: inst = 32'h10408000;
      36980: inst = 32'hc404ed2;
      36981: inst = 32'h8220000;
      36982: inst = 32'h10408000;
      36983: inst = 32'hc404ed3;
      36984: inst = 32'h8220000;
      36985: inst = 32'h10408000;
      36986: inst = 32'hc404ed4;
      36987: inst = 32'h8220000;
      36988: inst = 32'h10408000;
      36989: inst = 32'hc404ed5;
      36990: inst = 32'h8220000;
      36991: inst = 32'h10408000;
      36992: inst = 32'hc404ed6;
      36993: inst = 32'h8220000;
      36994: inst = 32'h10408000;
      36995: inst = 32'hc404ed7;
      36996: inst = 32'h8220000;
      36997: inst = 32'h10408000;
      36998: inst = 32'hc404ed8;
      36999: inst = 32'h8220000;
      37000: inst = 32'h10408000;
      37001: inst = 32'hc404ed9;
      37002: inst = 32'h8220000;
      37003: inst = 32'h10408000;
      37004: inst = 32'hc404eda;
      37005: inst = 32'h8220000;
      37006: inst = 32'h10408000;
      37007: inst = 32'hc404edb;
      37008: inst = 32'h8220000;
      37009: inst = 32'h10408000;
      37010: inst = 32'hc404edc;
      37011: inst = 32'h8220000;
      37012: inst = 32'h10408000;
      37013: inst = 32'hc404ee3;
      37014: inst = 32'h8220000;
      37015: inst = 32'h10408000;
      37016: inst = 32'hc404ee4;
      37017: inst = 32'h8220000;
      37018: inst = 32'h10408000;
      37019: inst = 32'hc404ee5;
      37020: inst = 32'h8220000;
      37021: inst = 32'h10408000;
      37022: inst = 32'hc404ee6;
      37023: inst = 32'h8220000;
      37024: inst = 32'h10408000;
      37025: inst = 32'hc404ee7;
      37026: inst = 32'h8220000;
      37027: inst = 32'h10408000;
      37028: inst = 32'hc404ee8;
      37029: inst = 32'h8220000;
      37030: inst = 32'h10408000;
      37031: inst = 32'hc404ee9;
      37032: inst = 32'h8220000;
      37033: inst = 32'h10408000;
      37034: inst = 32'hc404eea;
      37035: inst = 32'h8220000;
      37036: inst = 32'h10408000;
      37037: inst = 32'hc404eeb;
      37038: inst = 32'h8220000;
      37039: inst = 32'h10408000;
      37040: inst = 32'hc404eec;
      37041: inst = 32'h8220000;
      37042: inst = 32'h10408000;
      37043: inst = 32'hc404eed;
      37044: inst = 32'h8220000;
      37045: inst = 32'h10408000;
      37046: inst = 32'hc404eee;
      37047: inst = 32'h8220000;
      37048: inst = 32'h10408000;
      37049: inst = 32'hc404eef;
      37050: inst = 32'h8220000;
      37051: inst = 32'h10408000;
      37052: inst = 32'hc404ef0;
      37053: inst = 32'h8220000;
      37054: inst = 32'h10408000;
      37055: inst = 32'hc404ef1;
      37056: inst = 32'h8220000;
      37057: inst = 32'h10408000;
      37058: inst = 32'hc404ef2;
      37059: inst = 32'h8220000;
      37060: inst = 32'h10408000;
      37061: inst = 32'hc404ef3;
      37062: inst = 32'h8220000;
      37063: inst = 32'h10408000;
      37064: inst = 32'hc404ef4;
      37065: inst = 32'h8220000;
      37066: inst = 32'h10408000;
      37067: inst = 32'hc404ef5;
      37068: inst = 32'h8220000;
      37069: inst = 32'h10408000;
      37070: inst = 32'hc404ef6;
      37071: inst = 32'h8220000;
      37072: inst = 32'h10408000;
      37073: inst = 32'hc404ef7;
      37074: inst = 32'h8220000;
      37075: inst = 32'h10408000;
      37076: inst = 32'hc404ef8;
      37077: inst = 32'h8220000;
      37078: inst = 32'h10408000;
      37079: inst = 32'hc404ef9;
      37080: inst = 32'h8220000;
      37081: inst = 32'h10408000;
      37082: inst = 32'hc404efa;
      37083: inst = 32'h8220000;
      37084: inst = 32'h10408000;
      37085: inst = 32'hc404efb;
      37086: inst = 32'h8220000;
      37087: inst = 32'h10408000;
      37088: inst = 32'hc404efc;
      37089: inst = 32'h8220000;
      37090: inst = 32'h10408000;
      37091: inst = 32'hc404efd;
      37092: inst = 32'h8220000;
      37093: inst = 32'h10408000;
      37094: inst = 32'hc404efe;
      37095: inst = 32'h8220000;
      37096: inst = 32'h10408000;
      37097: inst = 32'hc404eff;
      37098: inst = 32'h8220000;
      37099: inst = 32'h10408000;
      37100: inst = 32'hc404f00;
      37101: inst = 32'h8220000;
      37102: inst = 32'h10408000;
      37103: inst = 32'hc404f01;
      37104: inst = 32'h8220000;
      37105: inst = 32'h10408000;
      37106: inst = 32'hc404f02;
      37107: inst = 32'h8220000;
      37108: inst = 32'h10408000;
      37109: inst = 32'hc404f03;
      37110: inst = 32'h8220000;
      37111: inst = 32'h10408000;
      37112: inst = 32'hc404f04;
      37113: inst = 32'h8220000;
      37114: inst = 32'h10408000;
      37115: inst = 32'hc404f05;
      37116: inst = 32'h8220000;
      37117: inst = 32'h10408000;
      37118: inst = 32'hc404f06;
      37119: inst = 32'h8220000;
      37120: inst = 32'h10408000;
      37121: inst = 32'hc404f07;
      37122: inst = 32'h8220000;
      37123: inst = 32'h10408000;
      37124: inst = 32'hc404f08;
      37125: inst = 32'h8220000;
      37126: inst = 32'h10408000;
      37127: inst = 32'hc404f09;
      37128: inst = 32'h8220000;
      37129: inst = 32'h10408000;
      37130: inst = 32'hc404f0a;
      37131: inst = 32'h8220000;
      37132: inst = 32'h10408000;
      37133: inst = 32'hc404f0b;
      37134: inst = 32'h8220000;
      37135: inst = 32'h10408000;
      37136: inst = 32'hc404f0c;
      37137: inst = 32'h8220000;
      37138: inst = 32'h10408000;
      37139: inst = 32'hc404f0d;
      37140: inst = 32'h8220000;
      37141: inst = 32'h10408000;
      37142: inst = 32'hc404f0e;
      37143: inst = 32'h8220000;
      37144: inst = 32'h10408000;
      37145: inst = 32'hc404f0f;
      37146: inst = 32'h8220000;
      37147: inst = 32'h10408000;
      37148: inst = 32'hc404f10;
      37149: inst = 32'h8220000;
      37150: inst = 32'h10408000;
      37151: inst = 32'hc404f11;
      37152: inst = 32'h8220000;
      37153: inst = 32'h10408000;
      37154: inst = 32'hc404f12;
      37155: inst = 32'h8220000;
      37156: inst = 32'h10408000;
      37157: inst = 32'hc404f13;
      37158: inst = 32'h8220000;
      37159: inst = 32'h10408000;
      37160: inst = 32'hc404f14;
      37161: inst = 32'h8220000;
      37162: inst = 32'h10408000;
      37163: inst = 32'hc404f15;
      37164: inst = 32'h8220000;
      37165: inst = 32'h10408000;
      37166: inst = 32'hc404f16;
      37167: inst = 32'h8220000;
      37168: inst = 32'h10408000;
      37169: inst = 32'hc404f17;
      37170: inst = 32'h8220000;
      37171: inst = 32'h10408000;
      37172: inst = 32'hc404f1b;
      37173: inst = 32'h8220000;
      37174: inst = 32'h10408000;
      37175: inst = 32'hc404f1c;
      37176: inst = 32'h8220000;
      37177: inst = 32'h10408000;
      37178: inst = 32'hc404f1d;
      37179: inst = 32'h8220000;
      37180: inst = 32'h10408000;
      37181: inst = 32'hc404f1e;
      37182: inst = 32'h8220000;
      37183: inst = 32'h10408000;
      37184: inst = 32'hc404f1f;
      37185: inst = 32'h8220000;
      37186: inst = 32'h10408000;
      37187: inst = 32'hc404f20;
      37188: inst = 32'h8220000;
      37189: inst = 32'h10408000;
      37190: inst = 32'hc404f21;
      37191: inst = 32'h8220000;
      37192: inst = 32'h10408000;
      37193: inst = 32'hc404f22;
      37194: inst = 32'h8220000;
      37195: inst = 32'h10408000;
      37196: inst = 32'hc404f23;
      37197: inst = 32'h8220000;
      37198: inst = 32'h10408000;
      37199: inst = 32'hc404f24;
      37200: inst = 32'h8220000;
      37201: inst = 32'h10408000;
      37202: inst = 32'hc404f25;
      37203: inst = 32'h8220000;
      37204: inst = 32'h10408000;
      37205: inst = 32'hc404f26;
      37206: inst = 32'h8220000;
      37207: inst = 32'h10408000;
      37208: inst = 32'hc404f27;
      37209: inst = 32'h8220000;
      37210: inst = 32'h10408000;
      37211: inst = 32'hc404f28;
      37212: inst = 32'h8220000;
      37213: inst = 32'h10408000;
      37214: inst = 32'hc404f29;
      37215: inst = 32'h8220000;
      37216: inst = 32'h10408000;
      37217: inst = 32'hc404f2a;
      37218: inst = 32'h8220000;
      37219: inst = 32'h10408000;
      37220: inst = 32'hc404f2b;
      37221: inst = 32'h8220000;
      37222: inst = 32'h10408000;
      37223: inst = 32'hc404f2c;
      37224: inst = 32'h8220000;
      37225: inst = 32'h10408000;
      37226: inst = 32'hc404f2d;
      37227: inst = 32'h8220000;
      37228: inst = 32'h10408000;
      37229: inst = 32'hc404f2e;
      37230: inst = 32'h8220000;
      37231: inst = 32'h10408000;
      37232: inst = 32'hc404f2f;
      37233: inst = 32'h8220000;
      37234: inst = 32'h10408000;
      37235: inst = 32'hc404f30;
      37236: inst = 32'h8220000;
      37237: inst = 32'h10408000;
      37238: inst = 32'hc404f31;
      37239: inst = 32'h8220000;
      37240: inst = 32'h10408000;
      37241: inst = 32'hc404f32;
      37242: inst = 32'h8220000;
      37243: inst = 32'h10408000;
      37244: inst = 32'hc404f33;
      37245: inst = 32'h8220000;
      37246: inst = 32'h10408000;
      37247: inst = 32'hc404f34;
      37248: inst = 32'h8220000;
      37249: inst = 32'h10408000;
      37250: inst = 32'hc404f35;
      37251: inst = 32'h8220000;
      37252: inst = 32'h10408000;
      37253: inst = 32'hc404f36;
      37254: inst = 32'h8220000;
      37255: inst = 32'h10408000;
      37256: inst = 32'hc404f37;
      37257: inst = 32'h8220000;
      37258: inst = 32'h10408000;
      37259: inst = 32'hc404f38;
      37260: inst = 32'h8220000;
      37261: inst = 32'h10408000;
      37262: inst = 32'hc404f39;
      37263: inst = 32'h8220000;
      37264: inst = 32'h10408000;
      37265: inst = 32'hc404f3a;
      37266: inst = 32'h8220000;
      37267: inst = 32'h10408000;
      37268: inst = 32'hc404f3b;
      37269: inst = 32'h8220000;
      37270: inst = 32'h10408000;
      37271: inst = 32'hc404f3c;
      37272: inst = 32'h8220000;
      37273: inst = 32'h10408000;
      37274: inst = 32'hc404f43;
      37275: inst = 32'h8220000;
      37276: inst = 32'h10408000;
      37277: inst = 32'hc404f44;
      37278: inst = 32'h8220000;
      37279: inst = 32'h10408000;
      37280: inst = 32'hc404f45;
      37281: inst = 32'h8220000;
      37282: inst = 32'h10408000;
      37283: inst = 32'hc404f46;
      37284: inst = 32'h8220000;
      37285: inst = 32'h10408000;
      37286: inst = 32'hc404f47;
      37287: inst = 32'h8220000;
      37288: inst = 32'h10408000;
      37289: inst = 32'hc404f48;
      37290: inst = 32'h8220000;
      37291: inst = 32'h10408000;
      37292: inst = 32'hc404f49;
      37293: inst = 32'h8220000;
      37294: inst = 32'h10408000;
      37295: inst = 32'hc404f4a;
      37296: inst = 32'h8220000;
      37297: inst = 32'h10408000;
      37298: inst = 32'hc404f4b;
      37299: inst = 32'h8220000;
      37300: inst = 32'h10408000;
      37301: inst = 32'hc404f4c;
      37302: inst = 32'h8220000;
      37303: inst = 32'h10408000;
      37304: inst = 32'hc404f4d;
      37305: inst = 32'h8220000;
      37306: inst = 32'h10408000;
      37307: inst = 32'hc404f4e;
      37308: inst = 32'h8220000;
      37309: inst = 32'h10408000;
      37310: inst = 32'hc404f4f;
      37311: inst = 32'h8220000;
      37312: inst = 32'h10408000;
      37313: inst = 32'hc404f50;
      37314: inst = 32'h8220000;
      37315: inst = 32'h10408000;
      37316: inst = 32'hc404f51;
      37317: inst = 32'h8220000;
      37318: inst = 32'h10408000;
      37319: inst = 32'hc404f52;
      37320: inst = 32'h8220000;
      37321: inst = 32'h10408000;
      37322: inst = 32'hc404f53;
      37323: inst = 32'h8220000;
      37324: inst = 32'h10408000;
      37325: inst = 32'hc404f54;
      37326: inst = 32'h8220000;
      37327: inst = 32'h10408000;
      37328: inst = 32'hc404f55;
      37329: inst = 32'h8220000;
      37330: inst = 32'h10408000;
      37331: inst = 32'hc404f56;
      37332: inst = 32'h8220000;
      37333: inst = 32'h10408000;
      37334: inst = 32'hc404f57;
      37335: inst = 32'h8220000;
      37336: inst = 32'h10408000;
      37337: inst = 32'hc404f58;
      37338: inst = 32'h8220000;
      37339: inst = 32'h10408000;
      37340: inst = 32'hc404f59;
      37341: inst = 32'h8220000;
      37342: inst = 32'h10408000;
      37343: inst = 32'hc404f5a;
      37344: inst = 32'h8220000;
      37345: inst = 32'h10408000;
      37346: inst = 32'hc404f5b;
      37347: inst = 32'h8220000;
      37348: inst = 32'h10408000;
      37349: inst = 32'hc404f5c;
      37350: inst = 32'h8220000;
      37351: inst = 32'h10408000;
      37352: inst = 32'hc404f5d;
      37353: inst = 32'h8220000;
      37354: inst = 32'h10408000;
      37355: inst = 32'hc404f5e;
      37356: inst = 32'h8220000;
      37357: inst = 32'h10408000;
      37358: inst = 32'hc404f5f;
      37359: inst = 32'h8220000;
      37360: inst = 32'h10408000;
      37361: inst = 32'hc404f60;
      37362: inst = 32'h8220000;
      37363: inst = 32'h10408000;
      37364: inst = 32'hc404f61;
      37365: inst = 32'h8220000;
      37366: inst = 32'h10408000;
      37367: inst = 32'hc404f62;
      37368: inst = 32'h8220000;
      37369: inst = 32'h10408000;
      37370: inst = 32'hc404f63;
      37371: inst = 32'h8220000;
      37372: inst = 32'h10408000;
      37373: inst = 32'hc404f64;
      37374: inst = 32'h8220000;
      37375: inst = 32'h10408000;
      37376: inst = 32'hc404f65;
      37377: inst = 32'h8220000;
      37378: inst = 32'h10408000;
      37379: inst = 32'hc404f66;
      37380: inst = 32'h8220000;
      37381: inst = 32'h10408000;
      37382: inst = 32'hc404f67;
      37383: inst = 32'h8220000;
      37384: inst = 32'h10408000;
      37385: inst = 32'hc404f68;
      37386: inst = 32'h8220000;
      37387: inst = 32'h10408000;
      37388: inst = 32'hc404f69;
      37389: inst = 32'h8220000;
      37390: inst = 32'h10408000;
      37391: inst = 32'hc404f6a;
      37392: inst = 32'h8220000;
      37393: inst = 32'h10408000;
      37394: inst = 32'hc404f6b;
      37395: inst = 32'h8220000;
      37396: inst = 32'h10408000;
      37397: inst = 32'hc404f6c;
      37398: inst = 32'h8220000;
      37399: inst = 32'h10408000;
      37400: inst = 32'hc404f6d;
      37401: inst = 32'h8220000;
      37402: inst = 32'h10408000;
      37403: inst = 32'hc404f6e;
      37404: inst = 32'h8220000;
      37405: inst = 32'h10408000;
      37406: inst = 32'hc404f6f;
      37407: inst = 32'h8220000;
      37408: inst = 32'h10408000;
      37409: inst = 32'hc404f70;
      37410: inst = 32'h8220000;
      37411: inst = 32'h10408000;
      37412: inst = 32'hc404f71;
      37413: inst = 32'h8220000;
      37414: inst = 32'h10408000;
      37415: inst = 32'hc404f72;
      37416: inst = 32'h8220000;
      37417: inst = 32'h10408000;
      37418: inst = 32'hc404f73;
      37419: inst = 32'h8220000;
      37420: inst = 32'h10408000;
      37421: inst = 32'hc404f74;
      37422: inst = 32'h8220000;
      37423: inst = 32'h10408000;
      37424: inst = 32'hc404f75;
      37425: inst = 32'h8220000;
      37426: inst = 32'h10408000;
      37427: inst = 32'hc404f76;
      37428: inst = 32'h8220000;
      37429: inst = 32'h10408000;
      37430: inst = 32'hc404f77;
      37431: inst = 32'h8220000;
      37432: inst = 32'h10408000;
      37433: inst = 32'hc404f7b;
      37434: inst = 32'h8220000;
      37435: inst = 32'h10408000;
      37436: inst = 32'hc404f7c;
      37437: inst = 32'h8220000;
      37438: inst = 32'h10408000;
      37439: inst = 32'hc404f7d;
      37440: inst = 32'h8220000;
      37441: inst = 32'h10408000;
      37442: inst = 32'hc404f7e;
      37443: inst = 32'h8220000;
      37444: inst = 32'h10408000;
      37445: inst = 32'hc404f7f;
      37446: inst = 32'h8220000;
      37447: inst = 32'h10408000;
      37448: inst = 32'hc404f80;
      37449: inst = 32'h8220000;
      37450: inst = 32'h10408000;
      37451: inst = 32'hc404f81;
      37452: inst = 32'h8220000;
      37453: inst = 32'h10408000;
      37454: inst = 32'hc404f82;
      37455: inst = 32'h8220000;
      37456: inst = 32'h10408000;
      37457: inst = 32'hc404f83;
      37458: inst = 32'h8220000;
      37459: inst = 32'h10408000;
      37460: inst = 32'hc404f84;
      37461: inst = 32'h8220000;
      37462: inst = 32'h10408000;
      37463: inst = 32'hc404f85;
      37464: inst = 32'h8220000;
      37465: inst = 32'h10408000;
      37466: inst = 32'hc404f86;
      37467: inst = 32'h8220000;
      37468: inst = 32'h10408000;
      37469: inst = 32'hc404f87;
      37470: inst = 32'h8220000;
      37471: inst = 32'h10408000;
      37472: inst = 32'hc404f88;
      37473: inst = 32'h8220000;
      37474: inst = 32'h10408000;
      37475: inst = 32'hc404f89;
      37476: inst = 32'h8220000;
      37477: inst = 32'h10408000;
      37478: inst = 32'hc404f8a;
      37479: inst = 32'h8220000;
      37480: inst = 32'h10408000;
      37481: inst = 32'hc404f8b;
      37482: inst = 32'h8220000;
      37483: inst = 32'h10408000;
      37484: inst = 32'hc404f8c;
      37485: inst = 32'h8220000;
      37486: inst = 32'h10408000;
      37487: inst = 32'hc404f8d;
      37488: inst = 32'h8220000;
      37489: inst = 32'h10408000;
      37490: inst = 32'hc404f8e;
      37491: inst = 32'h8220000;
      37492: inst = 32'h10408000;
      37493: inst = 32'hc404f8f;
      37494: inst = 32'h8220000;
      37495: inst = 32'h10408000;
      37496: inst = 32'hc404f90;
      37497: inst = 32'h8220000;
      37498: inst = 32'h10408000;
      37499: inst = 32'hc404f91;
      37500: inst = 32'h8220000;
      37501: inst = 32'h10408000;
      37502: inst = 32'hc404f92;
      37503: inst = 32'h8220000;
      37504: inst = 32'h10408000;
      37505: inst = 32'hc404f93;
      37506: inst = 32'h8220000;
      37507: inst = 32'h10408000;
      37508: inst = 32'hc404f94;
      37509: inst = 32'h8220000;
      37510: inst = 32'h10408000;
      37511: inst = 32'hc404f95;
      37512: inst = 32'h8220000;
      37513: inst = 32'h10408000;
      37514: inst = 32'hc404f96;
      37515: inst = 32'h8220000;
      37516: inst = 32'h10408000;
      37517: inst = 32'hc404f97;
      37518: inst = 32'h8220000;
      37519: inst = 32'h10408000;
      37520: inst = 32'hc404f98;
      37521: inst = 32'h8220000;
      37522: inst = 32'h10408000;
      37523: inst = 32'hc404f99;
      37524: inst = 32'h8220000;
      37525: inst = 32'h10408000;
      37526: inst = 32'hc404f9a;
      37527: inst = 32'h8220000;
      37528: inst = 32'h10408000;
      37529: inst = 32'hc404f9b;
      37530: inst = 32'h8220000;
      37531: inst = 32'h10408000;
      37532: inst = 32'hc404f9c;
      37533: inst = 32'h8220000;
      37534: inst = 32'h10408000;
      37535: inst = 32'hc404fa3;
      37536: inst = 32'h8220000;
      37537: inst = 32'h10408000;
      37538: inst = 32'hc404fa4;
      37539: inst = 32'h8220000;
      37540: inst = 32'h10408000;
      37541: inst = 32'hc404fa5;
      37542: inst = 32'h8220000;
      37543: inst = 32'h10408000;
      37544: inst = 32'hc404fa6;
      37545: inst = 32'h8220000;
      37546: inst = 32'h10408000;
      37547: inst = 32'hc404fa7;
      37548: inst = 32'h8220000;
      37549: inst = 32'h10408000;
      37550: inst = 32'hc404fa8;
      37551: inst = 32'h8220000;
      37552: inst = 32'h10408000;
      37553: inst = 32'hc404fa9;
      37554: inst = 32'h8220000;
      37555: inst = 32'h10408000;
      37556: inst = 32'hc404faa;
      37557: inst = 32'h8220000;
      37558: inst = 32'h10408000;
      37559: inst = 32'hc404fab;
      37560: inst = 32'h8220000;
      37561: inst = 32'h10408000;
      37562: inst = 32'hc404fac;
      37563: inst = 32'h8220000;
      37564: inst = 32'h10408000;
      37565: inst = 32'hc404fad;
      37566: inst = 32'h8220000;
      37567: inst = 32'h10408000;
      37568: inst = 32'hc404fae;
      37569: inst = 32'h8220000;
      37570: inst = 32'h10408000;
      37571: inst = 32'hc404faf;
      37572: inst = 32'h8220000;
      37573: inst = 32'h10408000;
      37574: inst = 32'hc404fb0;
      37575: inst = 32'h8220000;
      37576: inst = 32'h10408000;
      37577: inst = 32'hc404fb1;
      37578: inst = 32'h8220000;
      37579: inst = 32'h10408000;
      37580: inst = 32'hc404fb2;
      37581: inst = 32'h8220000;
      37582: inst = 32'h10408000;
      37583: inst = 32'hc404fb3;
      37584: inst = 32'h8220000;
      37585: inst = 32'h10408000;
      37586: inst = 32'hc404fb4;
      37587: inst = 32'h8220000;
      37588: inst = 32'h10408000;
      37589: inst = 32'hc404fb5;
      37590: inst = 32'h8220000;
      37591: inst = 32'h10408000;
      37592: inst = 32'hc404fb6;
      37593: inst = 32'h8220000;
      37594: inst = 32'h10408000;
      37595: inst = 32'hc404fb7;
      37596: inst = 32'h8220000;
      37597: inst = 32'h10408000;
      37598: inst = 32'hc404fb8;
      37599: inst = 32'h8220000;
      37600: inst = 32'h10408000;
      37601: inst = 32'hc404fb9;
      37602: inst = 32'h8220000;
      37603: inst = 32'h10408000;
      37604: inst = 32'hc404fba;
      37605: inst = 32'h8220000;
      37606: inst = 32'h10408000;
      37607: inst = 32'hc404fbb;
      37608: inst = 32'h8220000;
      37609: inst = 32'h10408000;
      37610: inst = 32'hc404fbc;
      37611: inst = 32'h8220000;
      37612: inst = 32'h10408000;
      37613: inst = 32'hc404fbd;
      37614: inst = 32'h8220000;
      37615: inst = 32'h10408000;
      37616: inst = 32'hc404fbe;
      37617: inst = 32'h8220000;
      37618: inst = 32'h10408000;
      37619: inst = 32'hc404fbf;
      37620: inst = 32'h8220000;
      37621: inst = 32'h10408000;
      37622: inst = 32'hc404fc0;
      37623: inst = 32'h8220000;
      37624: inst = 32'h10408000;
      37625: inst = 32'hc404fc1;
      37626: inst = 32'h8220000;
      37627: inst = 32'h10408000;
      37628: inst = 32'hc404fc2;
      37629: inst = 32'h8220000;
      37630: inst = 32'h10408000;
      37631: inst = 32'hc404fc3;
      37632: inst = 32'h8220000;
      37633: inst = 32'h10408000;
      37634: inst = 32'hc404fc4;
      37635: inst = 32'h8220000;
      37636: inst = 32'h10408000;
      37637: inst = 32'hc404fc5;
      37638: inst = 32'h8220000;
      37639: inst = 32'h10408000;
      37640: inst = 32'hc404fc6;
      37641: inst = 32'h8220000;
      37642: inst = 32'h10408000;
      37643: inst = 32'hc404fc7;
      37644: inst = 32'h8220000;
      37645: inst = 32'h10408000;
      37646: inst = 32'hc404fc8;
      37647: inst = 32'h8220000;
      37648: inst = 32'h10408000;
      37649: inst = 32'hc404fc9;
      37650: inst = 32'h8220000;
      37651: inst = 32'h10408000;
      37652: inst = 32'hc404fca;
      37653: inst = 32'h8220000;
      37654: inst = 32'h10408000;
      37655: inst = 32'hc404fcb;
      37656: inst = 32'h8220000;
      37657: inst = 32'h10408000;
      37658: inst = 32'hc404fcc;
      37659: inst = 32'h8220000;
      37660: inst = 32'h10408000;
      37661: inst = 32'hc404fcd;
      37662: inst = 32'h8220000;
      37663: inst = 32'h10408000;
      37664: inst = 32'hc404fce;
      37665: inst = 32'h8220000;
      37666: inst = 32'h10408000;
      37667: inst = 32'hc404fcf;
      37668: inst = 32'h8220000;
      37669: inst = 32'h10408000;
      37670: inst = 32'hc404fd0;
      37671: inst = 32'h8220000;
      37672: inst = 32'h10408000;
      37673: inst = 32'hc404fd1;
      37674: inst = 32'h8220000;
      37675: inst = 32'h10408000;
      37676: inst = 32'hc404fd2;
      37677: inst = 32'h8220000;
      37678: inst = 32'h10408000;
      37679: inst = 32'hc404fd3;
      37680: inst = 32'h8220000;
      37681: inst = 32'h10408000;
      37682: inst = 32'hc404fd4;
      37683: inst = 32'h8220000;
      37684: inst = 32'h10408000;
      37685: inst = 32'hc404fd5;
      37686: inst = 32'h8220000;
      37687: inst = 32'h10408000;
      37688: inst = 32'hc404fd6;
      37689: inst = 32'h8220000;
      37690: inst = 32'h10408000;
      37691: inst = 32'hc404fd7;
      37692: inst = 32'h8220000;
      37693: inst = 32'h10408000;
      37694: inst = 32'hc404fdb;
      37695: inst = 32'h8220000;
      37696: inst = 32'h10408000;
      37697: inst = 32'hc404fdc;
      37698: inst = 32'h8220000;
      37699: inst = 32'h10408000;
      37700: inst = 32'hc404fdd;
      37701: inst = 32'h8220000;
      37702: inst = 32'h10408000;
      37703: inst = 32'hc404fde;
      37704: inst = 32'h8220000;
      37705: inst = 32'h10408000;
      37706: inst = 32'hc404fdf;
      37707: inst = 32'h8220000;
      37708: inst = 32'h10408000;
      37709: inst = 32'hc404fe0;
      37710: inst = 32'h8220000;
      37711: inst = 32'h10408000;
      37712: inst = 32'hc404fe1;
      37713: inst = 32'h8220000;
      37714: inst = 32'h10408000;
      37715: inst = 32'hc404fe2;
      37716: inst = 32'h8220000;
      37717: inst = 32'h10408000;
      37718: inst = 32'hc404fe3;
      37719: inst = 32'h8220000;
      37720: inst = 32'h10408000;
      37721: inst = 32'hc404fe4;
      37722: inst = 32'h8220000;
      37723: inst = 32'h10408000;
      37724: inst = 32'hc404fe5;
      37725: inst = 32'h8220000;
      37726: inst = 32'h10408000;
      37727: inst = 32'hc404fe6;
      37728: inst = 32'h8220000;
      37729: inst = 32'h10408000;
      37730: inst = 32'hc404fe7;
      37731: inst = 32'h8220000;
      37732: inst = 32'h10408000;
      37733: inst = 32'hc404fe8;
      37734: inst = 32'h8220000;
      37735: inst = 32'h10408000;
      37736: inst = 32'hc404fe9;
      37737: inst = 32'h8220000;
      37738: inst = 32'h10408000;
      37739: inst = 32'hc404fea;
      37740: inst = 32'h8220000;
      37741: inst = 32'h10408000;
      37742: inst = 32'hc404feb;
      37743: inst = 32'h8220000;
      37744: inst = 32'h10408000;
      37745: inst = 32'hc404fec;
      37746: inst = 32'h8220000;
      37747: inst = 32'h10408000;
      37748: inst = 32'hc404fed;
      37749: inst = 32'h8220000;
      37750: inst = 32'h10408000;
      37751: inst = 32'hc404fee;
      37752: inst = 32'h8220000;
      37753: inst = 32'h10408000;
      37754: inst = 32'hc404fef;
      37755: inst = 32'h8220000;
      37756: inst = 32'h10408000;
      37757: inst = 32'hc404ff0;
      37758: inst = 32'h8220000;
      37759: inst = 32'h10408000;
      37760: inst = 32'hc404ff1;
      37761: inst = 32'h8220000;
      37762: inst = 32'h10408000;
      37763: inst = 32'hc404ff2;
      37764: inst = 32'h8220000;
      37765: inst = 32'h10408000;
      37766: inst = 32'hc404ff3;
      37767: inst = 32'h8220000;
      37768: inst = 32'h10408000;
      37769: inst = 32'hc404ff4;
      37770: inst = 32'h8220000;
      37771: inst = 32'h10408000;
      37772: inst = 32'hc404ff5;
      37773: inst = 32'h8220000;
      37774: inst = 32'h10408000;
      37775: inst = 32'hc404ff6;
      37776: inst = 32'h8220000;
      37777: inst = 32'h10408000;
      37778: inst = 32'hc404ff7;
      37779: inst = 32'h8220000;
      37780: inst = 32'h10408000;
      37781: inst = 32'hc404ff8;
      37782: inst = 32'h8220000;
      37783: inst = 32'h10408000;
      37784: inst = 32'hc404ff9;
      37785: inst = 32'h8220000;
      37786: inst = 32'h10408000;
      37787: inst = 32'hc404ffa;
      37788: inst = 32'h8220000;
      37789: inst = 32'h10408000;
      37790: inst = 32'hc404ffb;
      37791: inst = 32'h8220000;
      37792: inst = 32'h10408000;
      37793: inst = 32'hc404ffc;
      37794: inst = 32'h8220000;
      37795: inst = 32'h10408000;
      37796: inst = 32'hc405003;
      37797: inst = 32'h8220000;
      37798: inst = 32'h10408000;
      37799: inst = 32'hc405004;
      37800: inst = 32'h8220000;
      37801: inst = 32'h10408000;
      37802: inst = 32'hc405005;
      37803: inst = 32'h8220000;
      37804: inst = 32'h10408000;
      37805: inst = 32'hc405006;
      37806: inst = 32'h8220000;
      37807: inst = 32'h10408000;
      37808: inst = 32'hc405007;
      37809: inst = 32'h8220000;
      37810: inst = 32'h10408000;
      37811: inst = 32'hc405008;
      37812: inst = 32'h8220000;
      37813: inst = 32'h10408000;
      37814: inst = 32'hc405009;
      37815: inst = 32'h8220000;
      37816: inst = 32'h10408000;
      37817: inst = 32'hc40500a;
      37818: inst = 32'h8220000;
      37819: inst = 32'h10408000;
      37820: inst = 32'hc40500b;
      37821: inst = 32'h8220000;
      37822: inst = 32'h10408000;
      37823: inst = 32'hc40500c;
      37824: inst = 32'h8220000;
      37825: inst = 32'h10408000;
      37826: inst = 32'hc40500d;
      37827: inst = 32'h8220000;
      37828: inst = 32'h10408000;
      37829: inst = 32'hc40500e;
      37830: inst = 32'h8220000;
      37831: inst = 32'h10408000;
      37832: inst = 32'hc40500f;
      37833: inst = 32'h8220000;
      37834: inst = 32'h10408000;
      37835: inst = 32'hc405010;
      37836: inst = 32'h8220000;
      37837: inst = 32'h10408000;
      37838: inst = 32'hc405011;
      37839: inst = 32'h8220000;
      37840: inst = 32'h10408000;
      37841: inst = 32'hc405012;
      37842: inst = 32'h8220000;
      37843: inst = 32'h10408000;
      37844: inst = 32'hc405013;
      37845: inst = 32'h8220000;
      37846: inst = 32'h10408000;
      37847: inst = 32'hc405014;
      37848: inst = 32'h8220000;
      37849: inst = 32'h10408000;
      37850: inst = 32'hc405015;
      37851: inst = 32'h8220000;
      37852: inst = 32'h10408000;
      37853: inst = 32'hc405016;
      37854: inst = 32'h8220000;
      37855: inst = 32'h10408000;
      37856: inst = 32'hc405017;
      37857: inst = 32'h8220000;
      37858: inst = 32'h10408000;
      37859: inst = 32'hc405018;
      37860: inst = 32'h8220000;
      37861: inst = 32'h10408000;
      37862: inst = 32'hc405019;
      37863: inst = 32'h8220000;
      37864: inst = 32'h10408000;
      37865: inst = 32'hc40501a;
      37866: inst = 32'h8220000;
      37867: inst = 32'h10408000;
      37868: inst = 32'hc40501b;
      37869: inst = 32'h8220000;
      37870: inst = 32'h10408000;
      37871: inst = 32'hc40501c;
      37872: inst = 32'h8220000;
      37873: inst = 32'h10408000;
      37874: inst = 32'hc40501d;
      37875: inst = 32'h8220000;
      37876: inst = 32'h10408000;
      37877: inst = 32'hc40501e;
      37878: inst = 32'h8220000;
      37879: inst = 32'h10408000;
      37880: inst = 32'hc40501f;
      37881: inst = 32'h8220000;
      37882: inst = 32'h10408000;
      37883: inst = 32'hc405020;
      37884: inst = 32'h8220000;
      37885: inst = 32'h10408000;
      37886: inst = 32'hc405021;
      37887: inst = 32'h8220000;
      37888: inst = 32'h10408000;
      37889: inst = 32'hc405022;
      37890: inst = 32'h8220000;
      37891: inst = 32'h10408000;
      37892: inst = 32'hc405023;
      37893: inst = 32'h8220000;
      37894: inst = 32'h10408000;
      37895: inst = 32'hc405024;
      37896: inst = 32'h8220000;
      37897: inst = 32'h10408000;
      37898: inst = 32'hc405025;
      37899: inst = 32'h8220000;
      37900: inst = 32'h10408000;
      37901: inst = 32'hc405026;
      37902: inst = 32'h8220000;
      37903: inst = 32'h10408000;
      37904: inst = 32'hc405027;
      37905: inst = 32'h8220000;
      37906: inst = 32'h10408000;
      37907: inst = 32'hc405028;
      37908: inst = 32'h8220000;
      37909: inst = 32'h10408000;
      37910: inst = 32'hc405029;
      37911: inst = 32'h8220000;
      37912: inst = 32'h10408000;
      37913: inst = 32'hc40502a;
      37914: inst = 32'h8220000;
      37915: inst = 32'h10408000;
      37916: inst = 32'hc40502b;
      37917: inst = 32'h8220000;
      37918: inst = 32'h10408000;
      37919: inst = 32'hc40502c;
      37920: inst = 32'h8220000;
      37921: inst = 32'h10408000;
      37922: inst = 32'hc40502d;
      37923: inst = 32'h8220000;
      37924: inst = 32'h10408000;
      37925: inst = 32'hc40502e;
      37926: inst = 32'h8220000;
      37927: inst = 32'h10408000;
      37928: inst = 32'hc40502f;
      37929: inst = 32'h8220000;
      37930: inst = 32'h10408000;
      37931: inst = 32'hc405030;
      37932: inst = 32'h8220000;
      37933: inst = 32'h10408000;
      37934: inst = 32'hc405031;
      37935: inst = 32'h8220000;
      37936: inst = 32'h10408000;
      37937: inst = 32'hc405032;
      37938: inst = 32'h8220000;
      37939: inst = 32'h10408000;
      37940: inst = 32'hc405033;
      37941: inst = 32'h8220000;
      37942: inst = 32'h10408000;
      37943: inst = 32'hc405034;
      37944: inst = 32'h8220000;
      37945: inst = 32'h10408000;
      37946: inst = 32'hc405035;
      37947: inst = 32'h8220000;
      37948: inst = 32'h10408000;
      37949: inst = 32'hc405036;
      37950: inst = 32'h8220000;
      37951: inst = 32'h10408000;
      37952: inst = 32'hc405037;
      37953: inst = 32'h8220000;
      37954: inst = 32'h10408000;
      37955: inst = 32'hc40503b;
      37956: inst = 32'h8220000;
      37957: inst = 32'h10408000;
      37958: inst = 32'hc40503c;
      37959: inst = 32'h8220000;
      37960: inst = 32'h10408000;
      37961: inst = 32'hc40503d;
      37962: inst = 32'h8220000;
      37963: inst = 32'h10408000;
      37964: inst = 32'hc40503e;
      37965: inst = 32'h8220000;
      37966: inst = 32'h10408000;
      37967: inst = 32'hc40503f;
      37968: inst = 32'h8220000;
      37969: inst = 32'h10408000;
      37970: inst = 32'hc405040;
      37971: inst = 32'h8220000;
      37972: inst = 32'h10408000;
      37973: inst = 32'hc405041;
      37974: inst = 32'h8220000;
      37975: inst = 32'h10408000;
      37976: inst = 32'hc405042;
      37977: inst = 32'h8220000;
      37978: inst = 32'h10408000;
      37979: inst = 32'hc405043;
      37980: inst = 32'h8220000;
      37981: inst = 32'h10408000;
      37982: inst = 32'hc405044;
      37983: inst = 32'h8220000;
      37984: inst = 32'h10408000;
      37985: inst = 32'hc405045;
      37986: inst = 32'h8220000;
      37987: inst = 32'h10408000;
      37988: inst = 32'hc405046;
      37989: inst = 32'h8220000;
      37990: inst = 32'h10408000;
      37991: inst = 32'hc405047;
      37992: inst = 32'h8220000;
      37993: inst = 32'h10408000;
      37994: inst = 32'hc405048;
      37995: inst = 32'h8220000;
      37996: inst = 32'h10408000;
      37997: inst = 32'hc405049;
      37998: inst = 32'h8220000;
      37999: inst = 32'h10408000;
      38000: inst = 32'hc40504a;
      38001: inst = 32'h8220000;
      38002: inst = 32'h10408000;
      38003: inst = 32'hc40504b;
      38004: inst = 32'h8220000;
      38005: inst = 32'h10408000;
      38006: inst = 32'hc40504c;
      38007: inst = 32'h8220000;
      38008: inst = 32'h10408000;
      38009: inst = 32'hc40504d;
      38010: inst = 32'h8220000;
      38011: inst = 32'h10408000;
      38012: inst = 32'hc40504e;
      38013: inst = 32'h8220000;
      38014: inst = 32'h10408000;
      38015: inst = 32'hc40504f;
      38016: inst = 32'h8220000;
      38017: inst = 32'h10408000;
      38018: inst = 32'hc405050;
      38019: inst = 32'h8220000;
      38020: inst = 32'h10408000;
      38021: inst = 32'hc405051;
      38022: inst = 32'h8220000;
      38023: inst = 32'h10408000;
      38024: inst = 32'hc405052;
      38025: inst = 32'h8220000;
      38026: inst = 32'h10408000;
      38027: inst = 32'hc405053;
      38028: inst = 32'h8220000;
      38029: inst = 32'h10408000;
      38030: inst = 32'hc405054;
      38031: inst = 32'h8220000;
      38032: inst = 32'h10408000;
      38033: inst = 32'hc405055;
      38034: inst = 32'h8220000;
      38035: inst = 32'h10408000;
      38036: inst = 32'hc405056;
      38037: inst = 32'h8220000;
      38038: inst = 32'h10408000;
      38039: inst = 32'hc405057;
      38040: inst = 32'h8220000;
      38041: inst = 32'h10408000;
      38042: inst = 32'hc405058;
      38043: inst = 32'h8220000;
      38044: inst = 32'h10408000;
      38045: inst = 32'hc405059;
      38046: inst = 32'h8220000;
      38047: inst = 32'h10408000;
      38048: inst = 32'hc40505a;
      38049: inst = 32'h8220000;
      38050: inst = 32'h10408000;
      38051: inst = 32'hc40505b;
      38052: inst = 32'h8220000;
      38053: inst = 32'h10408000;
      38054: inst = 32'hc40505c;
      38055: inst = 32'h8220000;
      38056: inst = 32'h10408000;
      38057: inst = 32'hc405063;
      38058: inst = 32'h8220000;
      38059: inst = 32'h10408000;
      38060: inst = 32'hc405064;
      38061: inst = 32'h8220000;
      38062: inst = 32'h10408000;
      38063: inst = 32'hc405065;
      38064: inst = 32'h8220000;
      38065: inst = 32'h10408000;
      38066: inst = 32'hc405066;
      38067: inst = 32'h8220000;
      38068: inst = 32'h10408000;
      38069: inst = 32'hc405067;
      38070: inst = 32'h8220000;
      38071: inst = 32'h10408000;
      38072: inst = 32'hc405068;
      38073: inst = 32'h8220000;
      38074: inst = 32'h10408000;
      38075: inst = 32'hc405069;
      38076: inst = 32'h8220000;
      38077: inst = 32'h10408000;
      38078: inst = 32'hc40506a;
      38079: inst = 32'h8220000;
      38080: inst = 32'h10408000;
      38081: inst = 32'hc40506b;
      38082: inst = 32'h8220000;
      38083: inst = 32'h10408000;
      38084: inst = 32'hc40506c;
      38085: inst = 32'h8220000;
      38086: inst = 32'h10408000;
      38087: inst = 32'hc40506d;
      38088: inst = 32'h8220000;
      38089: inst = 32'h10408000;
      38090: inst = 32'hc40506e;
      38091: inst = 32'h8220000;
      38092: inst = 32'h10408000;
      38093: inst = 32'hc40506f;
      38094: inst = 32'h8220000;
      38095: inst = 32'h10408000;
      38096: inst = 32'hc405070;
      38097: inst = 32'h8220000;
      38098: inst = 32'h10408000;
      38099: inst = 32'hc405071;
      38100: inst = 32'h8220000;
      38101: inst = 32'h10408000;
      38102: inst = 32'hc405072;
      38103: inst = 32'h8220000;
      38104: inst = 32'h10408000;
      38105: inst = 32'hc405073;
      38106: inst = 32'h8220000;
      38107: inst = 32'h10408000;
      38108: inst = 32'hc405074;
      38109: inst = 32'h8220000;
      38110: inst = 32'h10408000;
      38111: inst = 32'hc405075;
      38112: inst = 32'h8220000;
      38113: inst = 32'h10408000;
      38114: inst = 32'hc405076;
      38115: inst = 32'h8220000;
      38116: inst = 32'h10408000;
      38117: inst = 32'hc405077;
      38118: inst = 32'h8220000;
      38119: inst = 32'h10408000;
      38120: inst = 32'hc405078;
      38121: inst = 32'h8220000;
      38122: inst = 32'h10408000;
      38123: inst = 32'hc405079;
      38124: inst = 32'h8220000;
      38125: inst = 32'h10408000;
      38126: inst = 32'hc40507a;
      38127: inst = 32'h8220000;
      38128: inst = 32'h10408000;
      38129: inst = 32'hc40507b;
      38130: inst = 32'h8220000;
      38131: inst = 32'h10408000;
      38132: inst = 32'hc40507c;
      38133: inst = 32'h8220000;
      38134: inst = 32'h10408000;
      38135: inst = 32'hc40507d;
      38136: inst = 32'h8220000;
      38137: inst = 32'h10408000;
      38138: inst = 32'hc40507e;
      38139: inst = 32'h8220000;
      38140: inst = 32'h10408000;
      38141: inst = 32'hc40507f;
      38142: inst = 32'h8220000;
      38143: inst = 32'h10408000;
      38144: inst = 32'hc405080;
      38145: inst = 32'h8220000;
      38146: inst = 32'h10408000;
      38147: inst = 32'hc405081;
      38148: inst = 32'h8220000;
      38149: inst = 32'h10408000;
      38150: inst = 32'hc405082;
      38151: inst = 32'h8220000;
      38152: inst = 32'h10408000;
      38153: inst = 32'hc405083;
      38154: inst = 32'h8220000;
      38155: inst = 32'h10408000;
      38156: inst = 32'hc405084;
      38157: inst = 32'h8220000;
      38158: inst = 32'h10408000;
      38159: inst = 32'hc405085;
      38160: inst = 32'h8220000;
      38161: inst = 32'h10408000;
      38162: inst = 32'hc405086;
      38163: inst = 32'h8220000;
      38164: inst = 32'h10408000;
      38165: inst = 32'hc405087;
      38166: inst = 32'h8220000;
      38167: inst = 32'h10408000;
      38168: inst = 32'hc405088;
      38169: inst = 32'h8220000;
      38170: inst = 32'h10408000;
      38171: inst = 32'hc405089;
      38172: inst = 32'h8220000;
      38173: inst = 32'h10408000;
      38174: inst = 32'hc40508a;
      38175: inst = 32'h8220000;
      38176: inst = 32'h10408000;
      38177: inst = 32'hc40508b;
      38178: inst = 32'h8220000;
      38179: inst = 32'h10408000;
      38180: inst = 32'hc40508c;
      38181: inst = 32'h8220000;
      38182: inst = 32'h10408000;
      38183: inst = 32'hc40508d;
      38184: inst = 32'h8220000;
      38185: inst = 32'h10408000;
      38186: inst = 32'hc40508e;
      38187: inst = 32'h8220000;
      38188: inst = 32'h10408000;
      38189: inst = 32'hc40508f;
      38190: inst = 32'h8220000;
      38191: inst = 32'h10408000;
      38192: inst = 32'hc405090;
      38193: inst = 32'h8220000;
      38194: inst = 32'h10408000;
      38195: inst = 32'hc405091;
      38196: inst = 32'h8220000;
      38197: inst = 32'h10408000;
      38198: inst = 32'hc405092;
      38199: inst = 32'h8220000;
      38200: inst = 32'h10408000;
      38201: inst = 32'hc405093;
      38202: inst = 32'h8220000;
      38203: inst = 32'h10408000;
      38204: inst = 32'hc405094;
      38205: inst = 32'h8220000;
      38206: inst = 32'h10408000;
      38207: inst = 32'hc405095;
      38208: inst = 32'h8220000;
      38209: inst = 32'h10408000;
      38210: inst = 32'hc405096;
      38211: inst = 32'h8220000;
      38212: inst = 32'h10408000;
      38213: inst = 32'hc405097;
      38214: inst = 32'h8220000;
      38215: inst = 32'h10408000;
      38216: inst = 32'hc4050c3;
      38217: inst = 32'h8220000;
      38218: inst = 32'h10408000;
      38219: inst = 32'hc4050c4;
      38220: inst = 32'h8220000;
      38221: inst = 32'h10408000;
      38222: inst = 32'hc4050c5;
      38223: inst = 32'h8220000;
      38224: inst = 32'h10408000;
      38225: inst = 32'hc4050c6;
      38226: inst = 32'h8220000;
      38227: inst = 32'h10408000;
      38228: inst = 32'hc4050c7;
      38229: inst = 32'h8220000;
      38230: inst = 32'h10408000;
      38231: inst = 32'hc4050c8;
      38232: inst = 32'h8220000;
      38233: inst = 32'h10408000;
      38234: inst = 32'hc4050c9;
      38235: inst = 32'h8220000;
      38236: inst = 32'h10408000;
      38237: inst = 32'hc4050ca;
      38238: inst = 32'h8220000;
      38239: inst = 32'h10408000;
      38240: inst = 32'hc4050cb;
      38241: inst = 32'h8220000;
      38242: inst = 32'h10408000;
      38243: inst = 32'hc4050cc;
      38244: inst = 32'h8220000;
      38245: inst = 32'h10408000;
      38246: inst = 32'hc4050cd;
      38247: inst = 32'h8220000;
      38248: inst = 32'h10408000;
      38249: inst = 32'hc4050ce;
      38250: inst = 32'h8220000;
      38251: inst = 32'h10408000;
      38252: inst = 32'hc4050cf;
      38253: inst = 32'h8220000;
      38254: inst = 32'h10408000;
      38255: inst = 32'hc4050d0;
      38256: inst = 32'h8220000;
      38257: inst = 32'h10408000;
      38258: inst = 32'hc4050d1;
      38259: inst = 32'h8220000;
      38260: inst = 32'h10408000;
      38261: inst = 32'hc4050d2;
      38262: inst = 32'h8220000;
      38263: inst = 32'h10408000;
      38264: inst = 32'hc4050d3;
      38265: inst = 32'h8220000;
      38266: inst = 32'h10408000;
      38267: inst = 32'hc4050d4;
      38268: inst = 32'h8220000;
      38269: inst = 32'h10408000;
      38270: inst = 32'hc4050d5;
      38271: inst = 32'h8220000;
      38272: inst = 32'h10408000;
      38273: inst = 32'hc4050d6;
      38274: inst = 32'h8220000;
      38275: inst = 32'h10408000;
      38276: inst = 32'hc4050d7;
      38277: inst = 32'h8220000;
      38278: inst = 32'h10408000;
      38279: inst = 32'hc4050d8;
      38280: inst = 32'h8220000;
      38281: inst = 32'h10408000;
      38282: inst = 32'hc4050d9;
      38283: inst = 32'h8220000;
      38284: inst = 32'h10408000;
      38285: inst = 32'hc4050da;
      38286: inst = 32'h8220000;
      38287: inst = 32'h10408000;
      38288: inst = 32'hc4050db;
      38289: inst = 32'h8220000;
      38290: inst = 32'h10408000;
      38291: inst = 32'hc4050dc;
      38292: inst = 32'h8220000;
      38293: inst = 32'h10408000;
      38294: inst = 32'hc4050dd;
      38295: inst = 32'h8220000;
      38296: inst = 32'h10408000;
      38297: inst = 32'hc4050de;
      38298: inst = 32'h8220000;
      38299: inst = 32'h10408000;
      38300: inst = 32'hc4050df;
      38301: inst = 32'h8220000;
      38302: inst = 32'h10408000;
      38303: inst = 32'hc4050e0;
      38304: inst = 32'h8220000;
      38305: inst = 32'h10408000;
      38306: inst = 32'hc4050e1;
      38307: inst = 32'h8220000;
      38308: inst = 32'h10408000;
      38309: inst = 32'hc4050e2;
      38310: inst = 32'h8220000;
      38311: inst = 32'h10408000;
      38312: inst = 32'hc4050e3;
      38313: inst = 32'h8220000;
      38314: inst = 32'h10408000;
      38315: inst = 32'hc4050e4;
      38316: inst = 32'h8220000;
      38317: inst = 32'h10408000;
      38318: inst = 32'hc4050e5;
      38319: inst = 32'h8220000;
      38320: inst = 32'h10408000;
      38321: inst = 32'hc4050e6;
      38322: inst = 32'h8220000;
      38323: inst = 32'h10408000;
      38324: inst = 32'hc4050e7;
      38325: inst = 32'h8220000;
      38326: inst = 32'h10408000;
      38327: inst = 32'hc4050e8;
      38328: inst = 32'h8220000;
      38329: inst = 32'h10408000;
      38330: inst = 32'hc4050e9;
      38331: inst = 32'h8220000;
      38332: inst = 32'h10408000;
      38333: inst = 32'hc4050ea;
      38334: inst = 32'h8220000;
      38335: inst = 32'h10408000;
      38336: inst = 32'hc4050eb;
      38337: inst = 32'h8220000;
      38338: inst = 32'h10408000;
      38339: inst = 32'hc4050ec;
      38340: inst = 32'h8220000;
      38341: inst = 32'h10408000;
      38342: inst = 32'hc4050ed;
      38343: inst = 32'h8220000;
      38344: inst = 32'h10408000;
      38345: inst = 32'hc4050ee;
      38346: inst = 32'h8220000;
      38347: inst = 32'h10408000;
      38348: inst = 32'hc4050ef;
      38349: inst = 32'h8220000;
      38350: inst = 32'h10408000;
      38351: inst = 32'hc4050f0;
      38352: inst = 32'h8220000;
      38353: inst = 32'h10408000;
      38354: inst = 32'hc4050f1;
      38355: inst = 32'h8220000;
      38356: inst = 32'h10408000;
      38357: inst = 32'hc4050f2;
      38358: inst = 32'h8220000;
      38359: inst = 32'h10408000;
      38360: inst = 32'hc4050f3;
      38361: inst = 32'h8220000;
      38362: inst = 32'h10408000;
      38363: inst = 32'hc4050f4;
      38364: inst = 32'h8220000;
      38365: inst = 32'h10408000;
      38366: inst = 32'hc4050f5;
      38367: inst = 32'h8220000;
      38368: inst = 32'h10408000;
      38369: inst = 32'hc4050f6;
      38370: inst = 32'h8220000;
      38371: inst = 32'h10408000;
      38372: inst = 32'hc4050f7;
      38373: inst = 32'h8220000;
      38374: inst = 32'h10408000;
      38375: inst = 32'hc405123;
      38376: inst = 32'h8220000;
      38377: inst = 32'h10408000;
      38378: inst = 32'hc405124;
      38379: inst = 32'h8220000;
      38380: inst = 32'h10408000;
      38381: inst = 32'hc405125;
      38382: inst = 32'h8220000;
      38383: inst = 32'h10408000;
      38384: inst = 32'hc405126;
      38385: inst = 32'h8220000;
      38386: inst = 32'h10408000;
      38387: inst = 32'hc405127;
      38388: inst = 32'h8220000;
      38389: inst = 32'h10408000;
      38390: inst = 32'hc405128;
      38391: inst = 32'h8220000;
      38392: inst = 32'h10408000;
      38393: inst = 32'hc405129;
      38394: inst = 32'h8220000;
      38395: inst = 32'h10408000;
      38396: inst = 32'hc40512a;
      38397: inst = 32'h8220000;
      38398: inst = 32'h10408000;
      38399: inst = 32'hc40512b;
      38400: inst = 32'h8220000;
      38401: inst = 32'h10408000;
      38402: inst = 32'hc40512c;
      38403: inst = 32'h8220000;
      38404: inst = 32'h10408000;
      38405: inst = 32'hc40512d;
      38406: inst = 32'h8220000;
      38407: inst = 32'h10408000;
      38408: inst = 32'hc40512e;
      38409: inst = 32'h8220000;
      38410: inst = 32'h10408000;
      38411: inst = 32'hc40512f;
      38412: inst = 32'h8220000;
      38413: inst = 32'h10408000;
      38414: inst = 32'hc405130;
      38415: inst = 32'h8220000;
      38416: inst = 32'h10408000;
      38417: inst = 32'hc405131;
      38418: inst = 32'h8220000;
      38419: inst = 32'h10408000;
      38420: inst = 32'hc405132;
      38421: inst = 32'h8220000;
      38422: inst = 32'h10408000;
      38423: inst = 32'hc405133;
      38424: inst = 32'h8220000;
      38425: inst = 32'h10408000;
      38426: inst = 32'hc405134;
      38427: inst = 32'h8220000;
      38428: inst = 32'h10408000;
      38429: inst = 32'hc405135;
      38430: inst = 32'h8220000;
      38431: inst = 32'h10408000;
      38432: inst = 32'hc405139;
      38433: inst = 32'h8220000;
      38434: inst = 32'h10408000;
      38435: inst = 32'hc40513a;
      38436: inst = 32'h8220000;
      38437: inst = 32'h10408000;
      38438: inst = 32'hc40513b;
      38439: inst = 32'h8220000;
      38440: inst = 32'h10408000;
      38441: inst = 32'hc40513c;
      38442: inst = 32'h8220000;
      38443: inst = 32'h10408000;
      38444: inst = 32'hc40513d;
      38445: inst = 32'h8220000;
      38446: inst = 32'h10408000;
      38447: inst = 32'hc40513e;
      38448: inst = 32'h8220000;
      38449: inst = 32'h10408000;
      38450: inst = 32'hc40513f;
      38451: inst = 32'h8220000;
      38452: inst = 32'h10408000;
      38453: inst = 32'hc405140;
      38454: inst = 32'h8220000;
      38455: inst = 32'h10408000;
      38456: inst = 32'hc405141;
      38457: inst = 32'h8220000;
      38458: inst = 32'h10408000;
      38459: inst = 32'hc405142;
      38460: inst = 32'h8220000;
      38461: inst = 32'h10408000;
      38462: inst = 32'hc405143;
      38463: inst = 32'h8220000;
      38464: inst = 32'h10408000;
      38465: inst = 32'hc405144;
      38466: inst = 32'h8220000;
      38467: inst = 32'h10408000;
      38468: inst = 32'hc405145;
      38469: inst = 32'h8220000;
      38470: inst = 32'h10408000;
      38471: inst = 32'hc405146;
      38472: inst = 32'h8220000;
      38473: inst = 32'h10408000;
      38474: inst = 32'hc405147;
      38475: inst = 32'h8220000;
      38476: inst = 32'h10408000;
      38477: inst = 32'hc405148;
      38478: inst = 32'h8220000;
      38479: inst = 32'h10408000;
      38480: inst = 32'hc405149;
      38481: inst = 32'h8220000;
      38482: inst = 32'h10408000;
      38483: inst = 32'hc40514a;
      38484: inst = 32'h8220000;
      38485: inst = 32'h10408000;
      38486: inst = 32'hc40514b;
      38487: inst = 32'h8220000;
      38488: inst = 32'h10408000;
      38489: inst = 32'hc40514c;
      38490: inst = 32'h8220000;
      38491: inst = 32'h10408000;
      38492: inst = 32'hc40514d;
      38493: inst = 32'h8220000;
      38494: inst = 32'h10408000;
      38495: inst = 32'hc40514e;
      38496: inst = 32'h8220000;
      38497: inst = 32'h10408000;
      38498: inst = 32'hc40514f;
      38499: inst = 32'h8220000;
      38500: inst = 32'h10408000;
      38501: inst = 32'hc405150;
      38502: inst = 32'h8220000;
      38503: inst = 32'h10408000;
      38504: inst = 32'hc405151;
      38505: inst = 32'h8220000;
      38506: inst = 32'h10408000;
      38507: inst = 32'hc405152;
      38508: inst = 32'h8220000;
      38509: inst = 32'h10408000;
      38510: inst = 32'hc405153;
      38511: inst = 32'h8220000;
      38512: inst = 32'h10408000;
      38513: inst = 32'hc405154;
      38514: inst = 32'h8220000;
      38515: inst = 32'h10408000;
      38516: inst = 32'hc405155;
      38517: inst = 32'h8220000;
      38518: inst = 32'h10408000;
      38519: inst = 32'hc405156;
      38520: inst = 32'h8220000;
      38521: inst = 32'h10408000;
      38522: inst = 32'hc405157;
      38523: inst = 32'h8220000;
      38524: inst = 32'h10408000;
      38525: inst = 32'hc405183;
      38526: inst = 32'h8220000;
      38527: inst = 32'h10408000;
      38528: inst = 32'hc405184;
      38529: inst = 32'h8220000;
      38530: inst = 32'h10408000;
      38531: inst = 32'hc405185;
      38532: inst = 32'h8220000;
      38533: inst = 32'h10408000;
      38534: inst = 32'hc405186;
      38535: inst = 32'h8220000;
      38536: inst = 32'h10408000;
      38537: inst = 32'hc405187;
      38538: inst = 32'h8220000;
      38539: inst = 32'h10408000;
      38540: inst = 32'hc405188;
      38541: inst = 32'h8220000;
      38542: inst = 32'h10408000;
      38543: inst = 32'hc405189;
      38544: inst = 32'h8220000;
      38545: inst = 32'h10408000;
      38546: inst = 32'hc40518a;
      38547: inst = 32'h8220000;
      38548: inst = 32'h10408000;
      38549: inst = 32'hc40518b;
      38550: inst = 32'h8220000;
      38551: inst = 32'h10408000;
      38552: inst = 32'hc40518c;
      38553: inst = 32'h8220000;
      38554: inst = 32'h10408000;
      38555: inst = 32'hc40518d;
      38556: inst = 32'h8220000;
      38557: inst = 32'h10408000;
      38558: inst = 32'hc40518e;
      38559: inst = 32'h8220000;
      38560: inst = 32'h10408000;
      38561: inst = 32'hc40518f;
      38562: inst = 32'h8220000;
      38563: inst = 32'h10408000;
      38564: inst = 32'hc405190;
      38565: inst = 32'h8220000;
      38566: inst = 32'h10408000;
      38567: inst = 32'hc405191;
      38568: inst = 32'h8220000;
      38569: inst = 32'h10408000;
      38570: inst = 32'hc405192;
      38571: inst = 32'h8220000;
      38572: inst = 32'h10408000;
      38573: inst = 32'hc405193;
      38574: inst = 32'h8220000;
      38575: inst = 32'h10408000;
      38576: inst = 32'hc405194;
      38577: inst = 32'h8220000;
      38578: inst = 32'h10408000;
      38579: inst = 32'hc405195;
      38580: inst = 32'h8220000;
      38581: inst = 32'h10408000;
      38582: inst = 32'hc405199;
      38583: inst = 32'h8220000;
      38584: inst = 32'h10408000;
      38585: inst = 32'hc40519a;
      38586: inst = 32'h8220000;
      38587: inst = 32'h10408000;
      38588: inst = 32'hc40519b;
      38589: inst = 32'h8220000;
      38590: inst = 32'h10408000;
      38591: inst = 32'hc40519c;
      38592: inst = 32'h8220000;
      38593: inst = 32'h10408000;
      38594: inst = 32'hc40519d;
      38595: inst = 32'h8220000;
      38596: inst = 32'h10408000;
      38597: inst = 32'hc40519e;
      38598: inst = 32'h8220000;
      38599: inst = 32'h10408000;
      38600: inst = 32'hc40519f;
      38601: inst = 32'h8220000;
      38602: inst = 32'h10408000;
      38603: inst = 32'hc4051a0;
      38604: inst = 32'h8220000;
      38605: inst = 32'h10408000;
      38606: inst = 32'hc4051a1;
      38607: inst = 32'h8220000;
      38608: inst = 32'h10408000;
      38609: inst = 32'hc4051a2;
      38610: inst = 32'h8220000;
      38611: inst = 32'h10408000;
      38612: inst = 32'hc4051a3;
      38613: inst = 32'h8220000;
      38614: inst = 32'h10408000;
      38615: inst = 32'hc4051a4;
      38616: inst = 32'h8220000;
      38617: inst = 32'h10408000;
      38618: inst = 32'hc4051a5;
      38619: inst = 32'h8220000;
      38620: inst = 32'h10408000;
      38621: inst = 32'hc4051a6;
      38622: inst = 32'h8220000;
      38623: inst = 32'h10408000;
      38624: inst = 32'hc4051a7;
      38625: inst = 32'h8220000;
      38626: inst = 32'h10408000;
      38627: inst = 32'hc4051a8;
      38628: inst = 32'h8220000;
      38629: inst = 32'h10408000;
      38630: inst = 32'hc4051a9;
      38631: inst = 32'h8220000;
      38632: inst = 32'h10408000;
      38633: inst = 32'hc4051aa;
      38634: inst = 32'h8220000;
      38635: inst = 32'h10408000;
      38636: inst = 32'hc4051ab;
      38637: inst = 32'h8220000;
      38638: inst = 32'h10408000;
      38639: inst = 32'hc4051ac;
      38640: inst = 32'h8220000;
      38641: inst = 32'h10408000;
      38642: inst = 32'hc4051ad;
      38643: inst = 32'h8220000;
      38644: inst = 32'h10408000;
      38645: inst = 32'hc4051ae;
      38646: inst = 32'h8220000;
      38647: inst = 32'h10408000;
      38648: inst = 32'hc4051af;
      38649: inst = 32'h8220000;
      38650: inst = 32'h10408000;
      38651: inst = 32'hc4051b0;
      38652: inst = 32'h8220000;
      38653: inst = 32'h10408000;
      38654: inst = 32'hc4051b1;
      38655: inst = 32'h8220000;
      38656: inst = 32'h10408000;
      38657: inst = 32'hc4051b2;
      38658: inst = 32'h8220000;
      38659: inst = 32'h10408000;
      38660: inst = 32'hc4051b3;
      38661: inst = 32'h8220000;
      38662: inst = 32'h10408000;
      38663: inst = 32'hc4051b4;
      38664: inst = 32'h8220000;
      38665: inst = 32'h10408000;
      38666: inst = 32'hc4051b5;
      38667: inst = 32'h8220000;
      38668: inst = 32'h10408000;
      38669: inst = 32'hc4051b6;
      38670: inst = 32'h8220000;
      38671: inst = 32'h10408000;
      38672: inst = 32'hc4051b7;
      38673: inst = 32'h8220000;
      38674: inst = 32'h10408000;
      38675: inst = 32'hc4051b8;
      38676: inst = 32'h8220000;
      38677: inst = 32'h10408000;
      38678: inst = 32'hc4051b9;
      38679: inst = 32'h8220000;
      38680: inst = 32'h10408000;
      38681: inst = 32'hc4051ba;
      38682: inst = 32'h8220000;
      38683: inst = 32'h10408000;
      38684: inst = 32'hc4051bb;
      38685: inst = 32'h8220000;
      38686: inst = 32'h10408000;
      38687: inst = 32'hc4051bc;
      38688: inst = 32'h8220000;
      38689: inst = 32'h10408000;
      38690: inst = 32'hc4051bd;
      38691: inst = 32'h8220000;
      38692: inst = 32'h10408000;
      38693: inst = 32'hc4051be;
      38694: inst = 32'h8220000;
      38695: inst = 32'h10408000;
      38696: inst = 32'hc4051bf;
      38697: inst = 32'h8220000;
      38698: inst = 32'h10408000;
      38699: inst = 32'hc4051c0;
      38700: inst = 32'h8220000;
      38701: inst = 32'h10408000;
      38702: inst = 32'hc4051c1;
      38703: inst = 32'h8220000;
      38704: inst = 32'h10408000;
      38705: inst = 32'hc4051c2;
      38706: inst = 32'h8220000;
      38707: inst = 32'h10408000;
      38708: inst = 32'hc4051c3;
      38709: inst = 32'h8220000;
      38710: inst = 32'h10408000;
      38711: inst = 32'hc4051c4;
      38712: inst = 32'h8220000;
      38713: inst = 32'h10408000;
      38714: inst = 32'hc4051c5;
      38715: inst = 32'h8220000;
      38716: inst = 32'h10408000;
      38717: inst = 32'hc4051c6;
      38718: inst = 32'h8220000;
      38719: inst = 32'h10408000;
      38720: inst = 32'hc4051c7;
      38721: inst = 32'h8220000;
      38722: inst = 32'h10408000;
      38723: inst = 32'hc4051c8;
      38724: inst = 32'h8220000;
      38725: inst = 32'h10408000;
      38726: inst = 32'hc4051c9;
      38727: inst = 32'h8220000;
      38728: inst = 32'h10408000;
      38729: inst = 32'hc4051ca;
      38730: inst = 32'h8220000;
      38731: inst = 32'h10408000;
      38732: inst = 32'hc4051cb;
      38733: inst = 32'h8220000;
      38734: inst = 32'h10408000;
      38735: inst = 32'hc4051cc;
      38736: inst = 32'h8220000;
      38737: inst = 32'h10408000;
      38738: inst = 32'hc4051cd;
      38739: inst = 32'h8220000;
      38740: inst = 32'h10408000;
      38741: inst = 32'hc4051ce;
      38742: inst = 32'h8220000;
      38743: inst = 32'h10408000;
      38744: inst = 32'hc4051cf;
      38745: inst = 32'h8220000;
      38746: inst = 32'h10408000;
      38747: inst = 32'hc4051d0;
      38748: inst = 32'h8220000;
      38749: inst = 32'h10408000;
      38750: inst = 32'hc4051d1;
      38751: inst = 32'h8220000;
      38752: inst = 32'h10408000;
      38753: inst = 32'hc4051d2;
      38754: inst = 32'h8220000;
      38755: inst = 32'h10408000;
      38756: inst = 32'hc4051d3;
      38757: inst = 32'h8220000;
      38758: inst = 32'h10408000;
      38759: inst = 32'hc4051d4;
      38760: inst = 32'h8220000;
      38761: inst = 32'h10408000;
      38762: inst = 32'hc4051d5;
      38763: inst = 32'h8220000;
      38764: inst = 32'h10408000;
      38765: inst = 32'hc4051d6;
      38766: inst = 32'h8220000;
      38767: inst = 32'h10408000;
      38768: inst = 32'hc4051d7;
      38769: inst = 32'h8220000;
      38770: inst = 32'h10408000;
      38771: inst = 32'hc4051d8;
      38772: inst = 32'h8220000;
      38773: inst = 32'h10408000;
      38774: inst = 32'hc4051d9;
      38775: inst = 32'h8220000;
      38776: inst = 32'h10408000;
      38777: inst = 32'hc4051da;
      38778: inst = 32'h8220000;
      38779: inst = 32'h10408000;
      38780: inst = 32'hc4051db;
      38781: inst = 32'h8220000;
      38782: inst = 32'h10408000;
      38783: inst = 32'hc4051dc;
      38784: inst = 32'h8220000;
      38785: inst = 32'h10408000;
      38786: inst = 32'hc4051e3;
      38787: inst = 32'h8220000;
      38788: inst = 32'h10408000;
      38789: inst = 32'hc4051e4;
      38790: inst = 32'h8220000;
      38791: inst = 32'h10408000;
      38792: inst = 32'hc4051e5;
      38793: inst = 32'h8220000;
      38794: inst = 32'h10408000;
      38795: inst = 32'hc4051e6;
      38796: inst = 32'h8220000;
      38797: inst = 32'h10408000;
      38798: inst = 32'hc4051e7;
      38799: inst = 32'h8220000;
      38800: inst = 32'h10408000;
      38801: inst = 32'hc4051e8;
      38802: inst = 32'h8220000;
      38803: inst = 32'h10408000;
      38804: inst = 32'hc4051e9;
      38805: inst = 32'h8220000;
      38806: inst = 32'h10408000;
      38807: inst = 32'hc4051ea;
      38808: inst = 32'h8220000;
      38809: inst = 32'h10408000;
      38810: inst = 32'hc4051eb;
      38811: inst = 32'h8220000;
      38812: inst = 32'h10408000;
      38813: inst = 32'hc4051ec;
      38814: inst = 32'h8220000;
      38815: inst = 32'h10408000;
      38816: inst = 32'hc4051ed;
      38817: inst = 32'h8220000;
      38818: inst = 32'h10408000;
      38819: inst = 32'hc4051ee;
      38820: inst = 32'h8220000;
      38821: inst = 32'h10408000;
      38822: inst = 32'hc4051ef;
      38823: inst = 32'h8220000;
      38824: inst = 32'h10408000;
      38825: inst = 32'hc4051f0;
      38826: inst = 32'h8220000;
      38827: inst = 32'h10408000;
      38828: inst = 32'hc4051f1;
      38829: inst = 32'h8220000;
      38830: inst = 32'h10408000;
      38831: inst = 32'hc4051f2;
      38832: inst = 32'h8220000;
      38833: inst = 32'h10408000;
      38834: inst = 32'hc4051f3;
      38835: inst = 32'h8220000;
      38836: inst = 32'h10408000;
      38837: inst = 32'hc4051f4;
      38838: inst = 32'h8220000;
      38839: inst = 32'h10408000;
      38840: inst = 32'hc4051f5;
      38841: inst = 32'h8220000;
      38842: inst = 32'h10408000;
      38843: inst = 32'hc4051f9;
      38844: inst = 32'h8220000;
      38845: inst = 32'h10408000;
      38846: inst = 32'hc4051fa;
      38847: inst = 32'h8220000;
      38848: inst = 32'h10408000;
      38849: inst = 32'hc4051fb;
      38850: inst = 32'h8220000;
      38851: inst = 32'h10408000;
      38852: inst = 32'hc4051fc;
      38853: inst = 32'h8220000;
      38854: inst = 32'h10408000;
      38855: inst = 32'hc4051fd;
      38856: inst = 32'h8220000;
      38857: inst = 32'h10408000;
      38858: inst = 32'hc4051fe;
      38859: inst = 32'h8220000;
      38860: inst = 32'h10408000;
      38861: inst = 32'hc4051ff;
      38862: inst = 32'h8220000;
      38863: inst = 32'h10408000;
      38864: inst = 32'hc405200;
      38865: inst = 32'h8220000;
      38866: inst = 32'h10408000;
      38867: inst = 32'hc405201;
      38868: inst = 32'h8220000;
      38869: inst = 32'h10408000;
      38870: inst = 32'hc405202;
      38871: inst = 32'h8220000;
      38872: inst = 32'h10408000;
      38873: inst = 32'hc405203;
      38874: inst = 32'h8220000;
      38875: inst = 32'h10408000;
      38876: inst = 32'hc405204;
      38877: inst = 32'h8220000;
      38878: inst = 32'h10408000;
      38879: inst = 32'hc405205;
      38880: inst = 32'h8220000;
      38881: inst = 32'h10408000;
      38882: inst = 32'hc405206;
      38883: inst = 32'h8220000;
      38884: inst = 32'h10408000;
      38885: inst = 32'hc405207;
      38886: inst = 32'h8220000;
      38887: inst = 32'h10408000;
      38888: inst = 32'hc405208;
      38889: inst = 32'h8220000;
      38890: inst = 32'h10408000;
      38891: inst = 32'hc405209;
      38892: inst = 32'h8220000;
      38893: inst = 32'h10408000;
      38894: inst = 32'hc40520a;
      38895: inst = 32'h8220000;
      38896: inst = 32'h10408000;
      38897: inst = 32'hc40520b;
      38898: inst = 32'h8220000;
      38899: inst = 32'h10408000;
      38900: inst = 32'hc40520c;
      38901: inst = 32'h8220000;
      38902: inst = 32'h10408000;
      38903: inst = 32'hc40520d;
      38904: inst = 32'h8220000;
      38905: inst = 32'h10408000;
      38906: inst = 32'hc40520e;
      38907: inst = 32'h8220000;
      38908: inst = 32'h10408000;
      38909: inst = 32'hc40520f;
      38910: inst = 32'h8220000;
      38911: inst = 32'h10408000;
      38912: inst = 32'hc405210;
      38913: inst = 32'h8220000;
      38914: inst = 32'h10408000;
      38915: inst = 32'hc405211;
      38916: inst = 32'h8220000;
      38917: inst = 32'h10408000;
      38918: inst = 32'hc405212;
      38919: inst = 32'h8220000;
      38920: inst = 32'h10408000;
      38921: inst = 32'hc405213;
      38922: inst = 32'h8220000;
      38923: inst = 32'h10408000;
      38924: inst = 32'hc405214;
      38925: inst = 32'h8220000;
      38926: inst = 32'h10408000;
      38927: inst = 32'hc405215;
      38928: inst = 32'h8220000;
      38929: inst = 32'h10408000;
      38930: inst = 32'hc405216;
      38931: inst = 32'h8220000;
      38932: inst = 32'h10408000;
      38933: inst = 32'hc405217;
      38934: inst = 32'h8220000;
      38935: inst = 32'h10408000;
      38936: inst = 32'hc405218;
      38937: inst = 32'h8220000;
      38938: inst = 32'h10408000;
      38939: inst = 32'hc405219;
      38940: inst = 32'h8220000;
      38941: inst = 32'h10408000;
      38942: inst = 32'hc40521a;
      38943: inst = 32'h8220000;
      38944: inst = 32'h10408000;
      38945: inst = 32'hc40521b;
      38946: inst = 32'h8220000;
      38947: inst = 32'h10408000;
      38948: inst = 32'hc40521c;
      38949: inst = 32'h8220000;
      38950: inst = 32'h10408000;
      38951: inst = 32'hc40521d;
      38952: inst = 32'h8220000;
      38953: inst = 32'h10408000;
      38954: inst = 32'hc40521e;
      38955: inst = 32'h8220000;
      38956: inst = 32'h10408000;
      38957: inst = 32'hc40521f;
      38958: inst = 32'h8220000;
      38959: inst = 32'h10408000;
      38960: inst = 32'hc405220;
      38961: inst = 32'h8220000;
      38962: inst = 32'h10408000;
      38963: inst = 32'hc405221;
      38964: inst = 32'h8220000;
      38965: inst = 32'h10408000;
      38966: inst = 32'hc405222;
      38967: inst = 32'h8220000;
      38968: inst = 32'h10408000;
      38969: inst = 32'hc405223;
      38970: inst = 32'h8220000;
      38971: inst = 32'h10408000;
      38972: inst = 32'hc405224;
      38973: inst = 32'h8220000;
      38974: inst = 32'h10408000;
      38975: inst = 32'hc405225;
      38976: inst = 32'h8220000;
      38977: inst = 32'h10408000;
      38978: inst = 32'hc405226;
      38979: inst = 32'h8220000;
      38980: inst = 32'h10408000;
      38981: inst = 32'hc405227;
      38982: inst = 32'h8220000;
      38983: inst = 32'h10408000;
      38984: inst = 32'hc405228;
      38985: inst = 32'h8220000;
      38986: inst = 32'h10408000;
      38987: inst = 32'hc405229;
      38988: inst = 32'h8220000;
      38989: inst = 32'h10408000;
      38990: inst = 32'hc40522a;
      38991: inst = 32'h8220000;
      38992: inst = 32'h10408000;
      38993: inst = 32'hc40522b;
      38994: inst = 32'h8220000;
      38995: inst = 32'h10408000;
      38996: inst = 32'hc40522c;
      38997: inst = 32'h8220000;
      38998: inst = 32'h10408000;
      38999: inst = 32'hc40522d;
      39000: inst = 32'h8220000;
      39001: inst = 32'h10408000;
      39002: inst = 32'hc40522e;
      39003: inst = 32'h8220000;
      39004: inst = 32'h10408000;
      39005: inst = 32'hc40522f;
      39006: inst = 32'h8220000;
      39007: inst = 32'h10408000;
      39008: inst = 32'hc405230;
      39009: inst = 32'h8220000;
      39010: inst = 32'h10408000;
      39011: inst = 32'hc405231;
      39012: inst = 32'h8220000;
      39013: inst = 32'h10408000;
      39014: inst = 32'hc405232;
      39015: inst = 32'h8220000;
      39016: inst = 32'h10408000;
      39017: inst = 32'hc405233;
      39018: inst = 32'h8220000;
      39019: inst = 32'h10408000;
      39020: inst = 32'hc405234;
      39021: inst = 32'h8220000;
      39022: inst = 32'h10408000;
      39023: inst = 32'hc405235;
      39024: inst = 32'h8220000;
      39025: inst = 32'h10408000;
      39026: inst = 32'hc405236;
      39027: inst = 32'h8220000;
      39028: inst = 32'h10408000;
      39029: inst = 32'hc405237;
      39030: inst = 32'h8220000;
      39031: inst = 32'h10408000;
      39032: inst = 32'hc405238;
      39033: inst = 32'h8220000;
      39034: inst = 32'h10408000;
      39035: inst = 32'hc405239;
      39036: inst = 32'h8220000;
      39037: inst = 32'h10408000;
      39038: inst = 32'hc40523a;
      39039: inst = 32'h8220000;
      39040: inst = 32'h10408000;
      39041: inst = 32'hc40523b;
      39042: inst = 32'h8220000;
      39043: inst = 32'h10408000;
      39044: inst = 32'hc40523c;
      39045: inst = 32'h8220000;
      39046: inst = 32'h10408000;
      39047: inst = 32'hc405243;
      39048: inst = 32'h8220000;
      39049: inst = 32'h10408000;
      39050: inst = 32'hc405244;
      39051: inst = 32'h8220000;
      39052: inst = 32'h10408000;
      39053: inst = 32'hc405245;
      39054: inst = 32'h8220000;
      39055: inst = 32'h10408000;
      39056: inst = 32'hc405246;
      39057: inst = 32'h8220000;
      39058: inst = 32'h10408000;
      39059: inst = 32'hc405247;
      39060: inst = 32'h8220000;
      39061: inst = 32'h10408000;
      39062: inst = 32'hc405248;
      39063: inst = 32'h8220000;
      39064: inst = 32'h10408000;
      39065: inst = 32'hc405249;
      39066: inst = 32'h8220000;
      39067: inst = 32'h10408000;
      39068: inst = 32'hc40524a;
      39069: inst = 32'h8220000;
      39070: inst = 32'h10408000;
      39071: inst = 32'hc40524b;
      39072: inst = 32'h8220000;
      39073: inst = 32'h10408000;
      39074: inst = 32'hc40524c;
      39075: inst = 32'h8220000;
      39076: inst = 32'h10408000;
      39077: inst = 32'hc40524d;
      39078: inst = 32'h8220000;
      39079: inst = 32'h10408000;
      39080: inst = 32'hc40524e;
      39081: inst = 32'h8220000;
      39082: inst = 32'h10408000;
      39083: inst = 32'hc40524f;
      39084: inst = 32'h8220000;
      39085: inst = 32'h10408000;
      39086: inst = 32'hc405250;
      39087: inst = 32'h8220000;
      39088: inst = 32'h10408000;
      39089: inst = 32'hc405251;
      39090: inst = 32'h8220000;
      39091: inst = 32'h10408000;
      39092: inst = 32'hc405252;
      39093: inst = 32'h8220000;
      39094: inst = 32'h10408000;
      39095: inst = 32'hc405253;
      39096: inst = 32'h8220000;
      39097: inst = 32'h10408000;
      39098: inst = 32'hc405254;
      39099: inst = 32'h8220000;
      39100: inst = 32'h10408000;
      39101: inst = 32'hc405255;
      39102: inst = 32'h8220000;
      39103: inst = 32'h10408000;
      39104: inst = 32'hc405259;
      39105: inst = 32'h8220000;
      39106: inst = 32'h10408000;
      39107: inst = 32'hc40525a;
      39108: inst = 32'h8220000;
      39109: inst = 32'h10408000;
      39110: inst = 32'hc40525b;
      39111: inst = 32'h8220000;
      39112: inst = 32'h10408000;
      39113: inst = 32'hc40525c;
      39114: inst = 32'h8220000;
      39115: inst = 32'h10408000;
      39116: inst = 32'hc40525d;
      39117: inst = 32'h8220000;
      39118: inst = 32'h10408000;
      39119: inst = 32'hc40525e;
      39120: inst = 32'h8220000;
      39121: inst = 32'h10408000;
      39122: inst = 32'hc40525f;
      39123: inst = 32'h8220000;
      39124: inst = 32'h10408000;
      39125: inst = 32'hc405260;
      39126: inst = 32'h8220000;
      39127: inst = 32'h10408000;
      39128: inst = 32'hc405261;
      39129: inst = 32'h8220000;
      39130: inst = 32'h10408000;
      39131: inst = 32'hc405262;
      39132: inst = 32'h8220000;
      39133: inst = 32'h10408000;
      39134: inst = 32'hc405263;
      39135: inst = 32'h8220000;
      39136: inst = 32'h10408000;
      39137: inst = 32'hc405264;
      39138: inst = 32'h8220000;
      39139: inst = 32'h10408000;
      39140: inst = 32'hc405265;
      39141: inst = 32'h8220000;
      39142: inst = 32'h10408000;
      39143: inst = 32'hc405266;
      39144: inst = 32'h8220000;
      39145: inst = 32'h10408000;
      39146: inst = 32'hc405267;
      39147: inst = 32'h8220000;
      39148: inst = 32'h10408000;
      39149: inst = 32'hc405268;
      39150: inst = 32'h8220000;
      39151: inst = 32'h10408000;
      39152: inst = 32'hc405269;
      39153: inst = 32'h8220000;
      39154: inst = 32'h10408000;
      39155: inst = 32'hc40526a;
      39156: inst = 32'h8220000;
      39157: inst = 32'h10408000;
      39158: inst = 32'hc40526b;
      39159: inst = 32'h8220000;
      39160: inst = 32'h10408000;
      39161: inst = 32'hc40526c;
      39162: inst = 32'h8220000;
      39163: inst = 32'h10408000;
      39164: inst = 32'hc40526d;
      39165: inst = 32'h8220000;
      39166: inst = 32'h10408000;
      39167: inst = 32'hc40526e;
      39168: inst = 32'h8220000;
      39169: inst = 32'h10408000;
      39170: inst = 32'hc40526f;
      39171: inst = 32'h8220000;
      39172: inst = 32'h10408000;
      39173: inst = 32'hc405270;
      39174: inst = 32'h8220000;
      39175: inst = 32'h10408000;
      39176: inst = 32'hc405271;
      39177: inst = 32'h8220000;
      39178: inst = 32'h10408000;
      39179: inst = 32'hc405272;
      39180: inst = 32'h8220000;
      39181: inst = 32'h10408000;
      39182: inst = 32'hc405273;
      39183: inst = 32'h8220000;
      39184: inst = 32'h10408000;
      39185: inst = 32'hc405274;
      39186: inst = 32'h8220000;
      39187: inst = 32'h10408000;
      39188: inst = 32'hc405275;
      39189: inst = 32'h8220000;
      39190: inst = 32'h10408000;
      39191: inst = 32'hc405276;
      39192: inst = 32'h8220000;
      39193: inst = 32'h10408000;
      39194: inst = 32'hc405277;
      39195: inst = 32'h8220000;
      39196: inst = 32'h10408000;
      39197: inst = 32'hc405278;
      39198: inst = 32'h8220000;
      39199: inst = 32'h10408000;
      39200: inst = 32'hc405279;
      39201: inst = 32'h8220000;
      39202: inst = 32'h10408000;
      39203: inst = 32'hc40527a;
      39204: inst = 32'h8220000;
      39205: inst = 32'h10408000;
      39206: inst = 32'hc40527b;
      39207: inst = 32'h8220000;
      39208: inst = 32'h10408000;
      39209: inst = 32'hc40527c;
      39210: inst = 32'h8220000;
      39211: inst = 32'h10408000;
      39212: inst = 32'hc40527d;
      39213: inst = 32'h8220000;
      39214: inst = 32'h10408000;
      39215: inst = 32'hc40527e;
      39216: inst = 32'h8220000;
      39217: inst = 32'h10408000;
      39218: inst = 32'hc40527f;
      39219: inst = 32'h8220000;
      39220: inst = 32'h10408000;
      39221: inst = 32'hc405280;
      39222: inst = 32'h8220000;
      39223: inst = 32'h10408000;
      39224: inst = 32'hc405281;
      39225: inst = 32'h8220000;
      39226: inst = 32'h10408000;
      39227: inst = 32'hc405282;
      39228: inst = 32'h8220000;
      39229: inst = 32'h10408000;
      39230: inst = 32'hc405283;
      39231: inst = 32'h8220000;
      39232: inst = 32'h10408000;
      39233: inst = 32'hc405284;
      39234: inst = 32'h8220000;
      39235: inst = 32'h10408000;
      39236: inst = 32'hc405285;
      39237: inst = 32'h8220000;
      39238: inst = 32'h10408000;
      39239: inst = 32'hc405286;
      39240: inst = 32'h8220000;
      39241: inst = 32'h10408000;
      39242: inst = 32'hc405287;
      39243: inst = 32'h8220000;
      39244: inst = 32'h10408000;
      39245: inst = 32'hc405288;
      39246: inst = 32'h8220000;
      39247: inst = 32'h10408000;
      39248: inst = 32'hc405289;
      39249: inst = 32'h8220000;
      39250: inst = 32'h10408000;
      39251: inst = 32'hc40528a;
      39252: inst = 32'h8220000;
      39253: inst = 32'h10408000;
      39254: inst = 32'hc40528b;
      39255: inst = 32'h8220000;
      39256: inst = 32'h10408000;
      39257: inst = 32'hc40528c;
      39258: inst = 32'h8220000;
      39259: inst = 32'h10408000;
      39260: inst = 32'hc40528d;
      39261: inst = 32'h8220000;
      39262: inst = 32'h10408000;
      39263: inst = 32'hc40528e;
      39264: inst = 32'h8220000;
      39265: inst = 32'h10408000;
      39266: inst = 32'hc40528f;
      39267: inst = 32'h8220000;
      39268: inst = 32'h10408000;
      39269: inst = 32'hc405290;
      39270: inst = 32'h8220000;
      39271: inst = 32'h10408000;
      39272: inst = 32'hc405291;
      39273: inst = 32'h8220000;
      39274: inst = 32'h10408000;
      39275: inst = 32'hc405292;
      39276: inst = 32'h8220000;
      39277: inst = 32'h10408000;
      39278: inst = 32'hc405293;
      39279: inst = 32'h8220000;
      39280: inst = 32'h10408000;
      39281: inst = 32'hc405294;
      39282: inst = 32'h8220000;
      39283: inst = 32'h10408000;
      39284: inst = 32'hc405295;
      39285: inst = 32'h8220000;
      39286: inst = 32'h10408000;
      39287: inst = 32'hc405296;
      39288: inst = 32'h8220000;
      39289: inst = 32'h10408000;
      39290: inst = 32'hc405297;
      39291: inst = 32'h8220000;
      39292: inst = 32'h10408000;
      39293: inst = 32'hc405298;
      39294: inst = 32'h8220000;
      39295: inst = 32'h10408000;
      39296: inst = 32'hc405299;
      39297: inst = 32'h8220000;
      39298: inst = 32'h10408000;
      39299: inst = 32'hc40529a;
      39300: inst = 32'h8220000;
      39301: inst = 32'h10408000;
      39302: inst = 32'hc40529b;
      39303: inst = 32'h8220000;
      39304: inst = 32'h10408000;
      39305: inst = 32'hc40529c;
      39306: inst = 32'h8220000;
      39307: inst = 32'h10408000;
      39308: inst = 32'hc4052a3;
      39309: inst = 32'h8220000;
      39310: inst = 32'h10408000;
      39311: inst = 32'hc4052a4;
      39312: inst = 32'h8220000;
      39313: inst = 32'h10408000;
      39314: inst = 32'hc4052a5;
      39315: inst = 32'h8220000;
      39316: inst = 32'h10408000;
      39317: inst = 32'hc4052a6;
      39318: inst = 32'h8220000;
      39319: inst = 32'h10408000;
      39320: inst = 32'hc4052a7;
      39321: inst = 32'h8220000;
      39322: inst = 32'h10408000;
      39323: inst = 32'hc4052a8;
      39324: inst = 32'h8220000;
      39325: inst = 32'h10408000;
      39326: inst = 32'hc4052a9;
      39327: inst = 32'h8220000;
      39328: inst = 32'h10408000;
      39329: inst = 32'hc4052aa;
      39330: inst = 32'h8220000;
      39331: inst = 32'h10408000;
      39332: inst = 32'hc4052ab;
      39333: inst = 32'h8220000;
      39334: inst = 32'h10408000;
      39335: inst = 32'hc4052ac;
      39336: inst = 32'h8220000;
      39337: inst = 32'h10408000;
      39338: inst = 32'hc4052ad;
      39339: inst = 32'h8220000;
      39340: inst = 32'h10408000;
      39341: inst = 32'hc4052ae;
      39342: inst = 32'h8220000;
      39343: inst = 32'h10408000;
      39344: inst = 32'hc4052af;
      39345: inst = 32'h8220000;
      39346: inst = 32'h10408000;
      39347: inst = 32'hc4052b0;
      39348: inst = 32'h8220000;
      39349: inst = 32'h10408000;
      39350: inst = 32'hc4052b1;
      39351: inst = 32'h8220000;
      39352: inst = 32'h10408000;
      39353: inst = 32'hc4052b2;
      39354: inst = 32'h8220000;
      39355: inst = 32'h10408000;
      39356: inst = 32'hc4052b3;
      39357: inst = 32'h8220000;
      39358: inst = 32'h10408000;
      39359: inst = 32'hc4052b4;
      39360: inst = 32'h8220000;
      39361: inst = 32'h10408000;
      39362: inst = 32'hc4052b5;
      39363: inst = 32'h8220000;
      39364: inst = 32'h10408000;
      39365: inst = 32'hc4052b9;
      39366: inst = 32'h8220000;
      39367: inst = 32'h10408000;
      39368: inst = 32'hc4052ba;
      39369: inst = 32'h8220000;
      39370: inst = 32'h10408000;
      39371: inst = 32'hc4052bb;
      39372: inst = 32'h8220000;
      39373: inst = 32'h10408000;
      39374: inst = 32'hc4052bc;
      39375: inst = 32'h8220000;
      39376: inst = 32'h10408000;
      39377: inst = 32'hc4052bd;
      39378: inst = 32'h8220000;
      39379: inst = 32'h10408000;
      39380: inst = 32'hc4052be;
      39381: inst = 32'h8220000;
      39382: inst = 32'h10408000;
      39383: inst = 32'hc4052bf;
      39384: inst = 32'h8220000;
      39385: inst = 32'h10408000;
      39386: inst = 32'hc4052c0;
      39387: inst = 32'h8220000;
      39388: inst = 32'h10408000;
      39389: inst = 32'hc4052c1;
      39390: inst = 32'h8220000;
      39391: inst = 32'h10408000;
      39392: inst = 32'hc4052c2;
      39393: inst = 32'h8220000;
      39394: inst = 32'h10408000;
      39395: inst = 32'hc4052c3;
      39396: inst = 32'h8220000;
      39397: inst = 32'h10408000;
      39398: inst = 32'hc4052c4;
      39399: inst = 32'h8220000;
      39400: inst = 32'h10408000;
      39401: inst = 32'hc4052c5;
      39402: inst = 32'h8220000;
      39403: inst = 32'h10408000;
      39404: inst = 32'hc4052c6;
      39405: inst = 32'h8220000;
      39406: inst = 32'h10408000;
      39407: inst = 32'hc4052c7;
      39408: inst = 32'h8220000;
      39409: inst = 32'h10408000;
      39410: inst = 32'hc4052c8;
      39411: inst = 32'h8220000;
      39412: inst = 32'h10408000;
      39413: inst = 32'hc4052c9;
      39414: inst = 32'h8220000;
      39415: inst = 32'h10408000;
      39416: inst = 32'hc4052ca;
      39417: inst = 32'h8220000;
      39418: inst = 32'h10408000;
      39419: inst = 32'hc4052cb;
      39420: inst = 32'h8220000;
      39421: inst = 32'h10408000;
      39422: inst = 32'hc4052cc;
      39423: inst = 32'h8220000;
      39424: inst = 32'h10408000;
      39425: inst = 32'hc4052cd;
      39426: inst = 32'h8220000;
      39427: inst = 32'h10408000;
      39428: inst = 32'hc4052ce;
      39429: inst = 32'h8220000;
      39430: inst = 32'h10408000;
      39431: inst = 32'hc4052cf;
      39432: inst = 32'h8220000;
      39433: inst = 32'h10408000;
      39434: inst = 32'hc4052d0;
      39435: inst = 32'h8220000;
      39436: inst = 32'h10408000;
      39437: inst = 32'hc4052d1;
      39438: inst = 32'h8220000;
      39439: inst = 32'h10408000;
      39440: inst = 32'hc4052d2;
      39441: inst = 32'h8220000;
      39442: inst = 32'h10408000;
      39443: inst = 32'hc4052d3;
      39444: inst = 32'h8220000;
      39445: inst = 32'h10408000;
      39446: inst = 32'hc4052d4;
      39447: inst = 32'h8220000;
      39448: inst = 32'h10408000;
      39449: inst = 32'hc4052d5;
      39450: inst = 32'h8220000;
      39451: inst = 32'h10408000;
      39452: inst = 32'hc4052d6;
      39453: inst = 32'h8220000;
      39454: inst = 32'h10408000;
      39455: inst = 32'hc4052d7;
      39456: inst = 32'h8220000;
      39457: inst = 32'h10408000;
      39458: inst = 32'hc4052d8;
      39459: inst = 32'h8220000;
      39460: inst = 32'h10408000;
      39461: inst = 32'hc4052d9;
      39462: inst = 32'h8220000;
      39463: inst = 32'h10408000;
      39464: inst = 32'hc4052da;
      39465: inst = 32'h8220000;
      39466: inst = 32'h10408000;
      39467: inst = 32'hc4052db;
      39468: inst = 32'h8220000;
      39469: inst = 32'h10408000;
      39470: inst = 32'hc4052dc;
      39471: inst = 32'h8220000;
      39472: inst = 32'h10408000;
      39473: inst = 32'hc4052dd;
      39474: inst = 32'h8220000;
      39475: inst = 32'h10408000;
      39476: inst = 32'hc4052de;
      39477: inst = 32'h8220000;
      39478: inst = 32'h10408000;
      39479: inst = 32'hc4052df;
      39480: inst = 32'h8220000;
      39481: inst = 32'h10408000;
      39482: inst = 32'hc4052e0;
      39483: inst = 32'h8220000;
      39484: inst = 32'h10408000;
      39485: inst = 32'hc4052e1;
      39486: inst = 32'h8220000;
      39487: inst = 32'h10408000;
      39488: inst = 32'hc4052e2;
      39489: inst = 32'h8220000;
      39490: inst = 32'h10408000;
      39491: inst = 32'hc4052e3;
      39492: inst = 32'h8220000;
      39493: inst = 32'h10408000;
      39494: inst = 32'hc4052e4;
      39495: inst = 32'h8220000;
      39496: inst = 32'h10408000;
      39497: inst = 32'hc4052e5;
      39498: inst = 32'h8220000;
      39499: inst = 32'h10408000;
      39500: inst = 32'hc4052e6;
      39501: inst = 32'h8220000;
      39502: inst = 32'h10408000;
      39503: inst = 32'hc4052e7;
      39504: inst = 32'h8220000;
      39505: inst = 32'h10408000;
      39506: inst = 32'hc4052e8;
      39507: inst = 32'h8220000;
      39508: inst = 32'h10408000;
      39509: inst = 32'hc4052e9;
      39510: inst = 32'h8220000;
      39511: inst = 32'h10408000;
      39512: inst = 32'hc4052ea;
      39513: inst = 32'h8220000;
      39514: inst = 32'h10408000;
      39515: inst = 32'hc4052eb;
      39516: inst = 32'h8220000;
      39517: inst = 32'h10408000;
      39518: inst = 32'hc4052ec;
      39519: inst = 32'h8220000;
      39520: inst = 32'h10408000;
      39521: inst = 32'hc4052ed;
      39522: inst = 32'h8220000;
      39523: inst = 32'h10408000;
      39524: inst = 32'hc4052ee;
      39525: inst = 32'h8220000;
      39526: inst = 32'h10408000;
      39527: inst = 32'hc4052ef;
      39528: inst = 32'h8220000;
      39529: inst = 32'h10408000;
      39530: inst = 32'hc4052f0;
      39531: inst = 32'h8220000;
      39532: inst = 32'h10408000;
      39533: inst = 32'hc4052f1;
      39534: inst = 32'h8220000;
      39535: inst = 32'h10408000;
      39536: inst = 32'hc4052f2;
      39537: inst = 32'h8220000;
      39538: inst = 32'h10408000;
      39539: inst = 32'hc4052f3;
      39540: inst = 32'h8220000;
      39541: inst = 32'h10408000;
      39542: inst = 32'hc4052f4;
      39543: inst = 32'h8220000;
      39544: inst = 32'h10408000;
      39545: inst = 32'hc4052f5;
      39546: inst = 32'h8220000;
      39547: inst = 32'h10408000;
      39548: inst = 32'hc4052f6;
      39549: inst = 32'h8220000;
      39550: inst = 32'h10408000;
      39551: inst = 32'hc4052f7;
      39552: inst = 32'h8220000;
      39553: inst = 32'h10408000;
      39554: inst = 32'hc4052f8;
      39555: inst = 32'h8220000;
      39556: inst = 32'h10408000;
      39557: inst = 32'hc4052f9;
      39558: inst = 32'h8220000;
      39559: inst = 32'h10408000;
      39560: inst = 32'hc4052fa;
      39561: inst = 32'h8220000;
      39562: inst = 32'h10408000;
      39563: inst = 32'hc4052fb;
      39564: inst = 32'h8220000;
      39565: inst = 32'h10408000;
      39566: inst = 32'hc4052fc;
      39567: inst = 32'h8220000;
      39568: inst = 32'h10408000;
      39569: inst = 32'hc405303;
      39570: inst = 32'h8220000;
      39571: inst = 32'h10408000;
      39572: inst = 32'hc405304;
      39573: inst = 32'h8220000;
      39574: inst = 32'h10408000;
      39575: inst = 32'hc405305;
      39576: inst = 32'h8220000;
      39577: inst = 32'h10408000;
      39578: inst = 32'hc405306;
      39579: inst = 32'h8220000;
      39580: inst = 32'h10408000;
      39581: inst = 32'hc405307;
      39582: inst = 32'h8220000;
      39583: inst = 32'h10408000;
      39584: inst = 32'hc405308;
      39585: inst = 32'h8220000;
      39586: inst = 32'h10408000;
      39587: inst = 32'hc405309;
      39588: inst = 32'h8220000;
      39589: inst = 32'h10408000;
      39590: inst = 32'hc40530a;
      39591: inst = 32'h8220000;
      39592: inst = 32'h10408000;
      39593: inst = 32'hc40530b;
      39594: inst = 32'h8220000;
      39595: inst = 32'h10408000;
      39596: inst = 32'hc40530c;
      39597: inst = 32'h8220000;
      39598: inst = 32'h10408000;
      39599: inst = 32'hc40530d;
      39600: inst = 32'h8220000;
      39601: inst = 32'h10408000;
      39602: inst = 32'hc40530e;
      39603: inst = 32'h8220000;
      39604: inst = 32'h10408000;
      39605: inst = 32'hc40530f;
      39606: inst = 32'h8220000;
      39607: inst = 32'h10408000;
      39608: inst = 32'hc405310;
      39609: inst = 32'h8220000;
      39610: inst = 32'h10408000;
      39611: inst = 32'hc405311;
      39612: inst = 32'h8220000;
      39613: inst = 32'h10408000;
      39614: inst = 32'hc405312;
      39615: inst = 32'h8220000;
      39616: inst = 32'h10408000;
      39617: inst = 32'hc405313;
      39618: inst = 32'h8220000;
      39619: inst = 32'h10408000;
      39620: inst = 32'hc405314;
      39621: inst = 32'h8220000;
      39622: inst = 32'h10408000;
      39623: inst = 32'hc405315;
      39624: inst = 32'h8220000;
      39625: inst = 32'h10408000;
      39626: inst = 32'hc405319;
      39627: inst = 32'h8220000;
      39628: inst = 32'h10408000;
      39629: inst = 32'hc40531a;
      39630: inst = 32'h8220000;
      39631: inst = 32'h10408000;
      39632: inst = 32'hc40531b;
      39633: inst = 32'h8220000;
      39634: inst = 32'h10408000;
      39635: inst = 32'hc40531c;
      39636: inst = 32'h8220000;
      39637: inst = 32'h10408000;
      39638: inst = 32'hc40531d;
      39639: inst = 32'h8220000;
      39640: inst = 32'h10408000;
      39641: inst = 32'hc40531e;
      39642: inst = 32'h8220000;
      39643: inst = 32'h10408000;
      39644: inst = 32'hc40531f;
      39645: inst = 32'h8220000;
      39646: inst = 32'h10408000;
      39647: inst = 32'hc405320;
      39648: inst = 32'h8220000;
      39649: inst = 32'h10408000;
      39650: inst = 32'hc405321;
      39651: inst = 32'h8220000;
      39652: inst = 32'h10408000;
      39653: inst = 32'hc405322;
      39654: inst = 32'h8220000;
      39655: inst = 32'h10408000;
      39656: inst = 32'hc405323;
      39657: inst = 32'h8220000;
      39658: inst = 32'h10408000;
      39659: inst = 32'hc405324;
      39660: inst = 32'h8220000;
      39661: inst = 32'h10408000;
      39662: inst = 32'hc405325;
      39663: inst = 32'h8220000;
      39664: inst = 32'h10408000;
      39665: inst = 32'hc405326;
      39666: inst = 32'h8220000;
      39667: inst = 32'h10408000;
      39668: inst = 32'hc405327;
      39669: inst = 32'h8220000;
      39670: inst = 32'h10408000;
      39671: inst = 32'hc405328;
      39672: inst = 32'h8220000;
      39673: inst = 32'h10408000;
      39674: inst = 32'hc405329;
      39675: inst = 32'h8220000;
      39676: inst = 32'h10408000;
      39677: inst = 32'hc40532a;
      39678: inst = 32'h8220000;
      39679: inst = 32'h10408000;
      39680: inst = 32'hc40532b;
      39681: inst = 32'h8220000;
      39682: inst = 32'h10408000;
      39683: inst = 32'hc40532c;
      39684: inst = 32'h8220000;
      39685: inst = 32'h10408000;
      39686: inst = 32'hc40532d;
      39687: inst = 32'h8220000;
      39688: inst = 32'h10408000;
      39689: inst = 32'hc40532e;
      39690: inst = 32'h8220000;
      39691: inst = 32'h10408000;
      39692: inst = 32'hc40532f;
      39693: inst = 32'h8220000;
      39694: inst = 32'h10408000;
      39695: inst = 32'hc405330;
      39696: inst = 32'h8220000;
      39697: inst = 32'h10408000;
      39698: inst = 32'hc405331;
      39699: inst = 32'h8220000;
      39700: inst = 32'h10408000;
      39701: inst = 32'hc405332;
      39702: inst = 32'h8220000;
      39703: inst = 32'h10408000;
      39704: inst = 32'hc405333;
      39705: inst = 32'h8220000;
      39706: inst = 32'h10408000;
      39707: inst = 32'hc405334;
      39708: inst = 32'h8220000;
      39709: inst = 32'h10408000;
      39710: inst = 32'hc405335;
      39711: inst = 32'h8220000;
      39712: inst = 32'h10408000;
      39713: inst = 32'hc405336;
      39714: inst = 32'h8220000;
      39715: inst = 32'h10408000;
      39716: inst = 32'hc405337;
      39717: inst = 32'h8220000;
      39718: inst = 32'h10408000;
      39719: inst = 32'hc405338;
      39720: inst = 32'h8220000;
      39721: inst = 32'h10408000;
      39722: inst = 32'hc405339;
      39723: inst = 32'h8220000;
      39724: inst = 32'h10408000;
      39725: inst = 32'hc40533a;
      39726: inst = 32'h8220000;
      39727: inst = 32'h10408000;
      39728: inst = 32'hc40533b;
      39729: inst = 32'h8220000;
      39730: inst = 32'h10408000;
      39731: inst = 32'hc40533c;
      39732: inst = 32'h8220000;
      39733: inst = 32'h10408000;
      39734: inst = 32'hc40533d;
      39735: inst = 32'h8220000;
      39736: inst = 32'h10408000;
      39737: inst = 32'hc40533e;
      39738: inst = 32'h8220000;
      39739: inst = 32'h10408000;
      39740: inst = 32'hc40533f;
      39741: inst = 32'h8220000;
      39742: inst = 32'h10408000;
      39743: inst = 32'hc405340;
      39744: inst = 32'h8220000;
      39745: inst = 32'h10408000;
      39746: inst = 32'hc405341;
      39747: inst = 32'h8220000;
      39748: inst = 32'h10408000;
      39749: inst = 32'hc405342;
      39750: inst = 32'h8220000;
      39751: inst = 32'h10408000;
      39752: inst = 32'hc405343;
      39753: inst = 32'h8220000;
      39754: inst = 32'h10408000;
      39755: inst = 32'hc405344;
      39756: inst = 32'h8220000;
      39757: inst = 32'h10408000;
      39758: inst = 32'hc405345;
      39759: inst = 32'h8220000;
      39760: inst = 32'h10408000;
      39761: inst = 32'hc405346;
      39762: inst = 32'h8220000;
      39763: inst = 32'h10408000;
      39764: inst = 32'hc405347;
      39765: inst = 32'h8220000;
      39766: inst = 32'h10408000;
      39767: inst = 32'hc405348;
      39768: inst = 32'h8220000;
      39769: inst = 32'h10408000;
      39770: inst = 32'hc405349;
      39771: inst = 32'h8220000;
      39772: inst = 32'h10408000;
      39773: inst = 32'hc40534a;
      39774: inst = 32'h8220000;
      39775: inst = 32'h10408000;
      39776: inst = 32'hc40534b;
      39777: inst = 32'h8220000;
      39778: inst = 32'h10408000;
      39779: inst = 32'hc40534c;
      39780: inst = 32'h8220000;
      39781: inst = 32'h10408000;
      39782: inst = 32'hc40534d;
      39783: inst = 32'h8220000;
      39784: inst = 32'h10408000;
      39785: inst = 32'hc40534e;
      39786: inst = 32'h8220000;
      39787: inst = 32'h10408000;
      39788: inst = 32'hc40534f;
      39789: inst = 32'h8220000;
      39790: inst = 32'h10408000;
      39791: inst = 32'hc405350;
      39792: inst = 32'h8220000;
      39793: inst = 32'h10408000;
      39794: inst = 32'hc405351;
      39795: inst = 32'h8220000;
      39796: inst = 32'h10408000;
      39797: inst = 32'hc40535c;
      39798: inst = 32'h8220000;
      39799: inst = 32'h10408000;
      39800: inst = 32'hc405363;
      39801: inst = 32'h8220000;
      39802: inst = 32'h10408000;
      39803: inst = 32'hc405364;
      39804: inst = 32'h8220000;
      39805: inst = 32'h10408000;
      39806: inst = 32'hc405365;
      39807: inst = 32'h8220000;
      39808: inst = 32'h10408000;
      39809: inst = 32'hc405366;
      39810: inst = 32'h8220000;
      39811: inst = 32'h10408000;
      39812: inst = 32'hc405367;
      39813: inst = 32'h8220000;
      39814: inst = 32'h10408000;
      39815: inst = 32'hc405368;
      39816: inst = 32'h8220000;
      39817: inst = 32'h10408000;
      39818: inst = 32'hc405369;
      39819: inst = 32'h8220000;
      39820: inst = 32'h10408000;
      39821: inst = 32'hc40536a;
      39822: inst = 32'h8220000;
      39823: inst = 32'h10408000;
      39824: inst = 32'hc40536b;
      39825: inst = 32'h8220000;
      39826: inst = 32'h10408000;
      39827: inst = 32'hc40536c;
      39828: inst = 32'h8220000;
      39829: inst = 32'h10408000;
      39830: inst = 32'hc40536d;
      39831: inst = 32'h8220000;
      39832: inst = 32'h10408000;
      39833: inst = 32'hc40536e;
      39834: inst = 32'h8220000;
      39835: inst = 32'h10408000;
      39836: inst = 32'hc40536f;
      39837: inst = 32'h8220000;
      39838: inst = 32'h10408000;
      39839: inst = 32'hc405370;
      39840: inst = 32'h8220000;
      39841: inst = 32'h10408000;
      39842: inst = 32'hc405371;
      39843: inst = 32'h8220000;
      39844: inst = 32'h10408000;
      39845: inst = 32'hc405372;
      39846: inst = 32'h8220000;
      39847: inst = 32'h10408000;
      39848: inst = 32'hc405373;
      39849: inst = 32'h8220000;
      39850: inst = 32'h10408000;
      39851: inst = 32'hc405374;
      39852: inst = 32'h8220000;
      39853: inst = 32'h10408000;
      39854: inst = 32'hc405375;
      39855: inst = 32'h8220000;
      39856: inst = 32'h10408000;
      39857: inst = 32'hc405379;
      39858: inst = 32'h8220000;
      39859: inst = 32'h10408000;
      39860: inst = 32'hc40537a;
      39861: inst = 32'h8220000;
      39862: inst = 32'h10408000;
      39863: inst = 32'hc40537b;
      39864: inst = 32'h8220000;
      39865: inst = 32'h10408000;
      39866: inst = 32'hc40537c;
      39867: inst = 32'h8220000;
      39868: inst = 32'h10408000;
      39869: inst = 32'hc40537d;
      39870: inst = 32'h8220000;
      39871: inst = 32'h10408000;
      39872: inst = 32'hc40537e;
      39873: inst = 32'h8220000;
      39874: inst = 32'h10408000;
      39875: inst = 32'hc40537f;
      39876: inst = 32'h8220000;
      39877: inst = 32'h10408000;
      39878: inst = 32'hc405380;
      39879: inst = 32'h8220000;
      39880: inst = 32'h10408000;
      39881: inst = 32'hc405381;
      39882: inst = 32'h8220000;
      39883: inst = 32'h10408000;
      39884: inst = 32'hc405382;
      39885: inst = 32'h8220000;
      39886: inst = 32'h10408000;
      39887: inst = 32'hc405383;
      39888: inst = 32'h8220000;
      39889: inst = 32'h10408000;
      39890: inst = 32'hc405384;
      39891: inst = 32'h8220000;
      39892: inst = 32'h10408000;
      39893: inst = 32'hc405385;
      39894: inst = 32'h8220000;
      39895: inst = 32'h10408000;
      39896: inst = 32'hc405386;
      39897: inst = 32'h8220000;
      39898: inst = 32'h10408000;
      39899: inst = 32'hc405387;
      39900: inst = 32'h8220000;
      39901: inst = 32'h10408000;
      39902: inst = 32'hc405388;
      39903: inst = 32'h8220000;
      39904: inst = 32'h10408000;
      39905: inst = 32'hc405389;
      39906: inst = 32'h8220000;
      39907: inst = 32'h10408000;
      39908: inst = 32'hc40538a;
      39909: inst = 32'h8220000;
      39910: inst = 32'h10408000;
      39911: inst = 32'hc40538b;
      39912: inst = 32'h8220000;
      39913: inst = 32'h10408000;
      39914: inst = 32'hc40538c;
      39915: inst = 32'h8220000;
      39916: inst = 32'h10408000;
      39917: inst = 32'hc40538d;
      39918: inst = 32'h8220000;
      39919: inst = 32'h10408000;
      39920: inst = 32'hc40538e;
      39921: inst = 32'h8220000;
      39922: inst = 32'h10408000;
      39923: inst = 32'hc40538f;
      39924: inst = 32'h8220000;
      39925: inst = 32'h10408000;
      39926: inst = 32'hc405390;
      39927: inst = 32'h8220000;
      39928: inst = 32'h10408000;
      39929: inst = 32'hc405391;
      39930: inst = 32'h8220000;
      39931: inst = 32'h10408000;
      39932: inst = 32'hc405392;
      39933: inst = 32'h8220000;
      39934: inst = 32'h10408000;
      39935: inst = 32'hc405393;
      39936: inst = 32'h8220000;
      39937: inst = 32'h10408000;
      39938: inst = 32'hc405394;
      39939: inst = 32'h8220000;
      39940: inst = 32'h10408000;
      39941: inst = 32'hc405395;
      39942: inst = 32'h8220000;
      39943: inst = 32'h10408000;
      39944: inst = 32'hc405396;
      39945: inst = 32'h8220000;
      39946: inst = 32'h10408000;
      39947: inst = 32'hc405397;
      39948: inst = 32'h8220000;
      39949: inst = 32'h10408000;
      39950: inst = 32'hc405398;
      39951: inst = 32'h8220000;
      39952: inst = 32'h10408000;
      39953: inst = 32'hc405399;
      39954: inst = 32'h8220000;
      39955: inst = 32'h10408000;
      39956: inst = 32'hc40539a;
      39957: inst = 32'h8220000;
      39958: inst = 32'h10408000;
      39959: inst = 32'hc40539b;
      39960: inst = 32'h8220000;
      39961: inst = 32'h10408000;
      39962: inst = 32'hc40539c;
      39963: inst = 32'h8220000;
      39964: inst = 32'h10408000;
      39965: inst = 32'hc40539d;
      39966: inst = 32'h8220000;
      39967: inst = 32'h10408000;
      39968: inst = 32'hc40539e;
      39969: inst = 32'h8220000;
      39970: inst = 32'h10408000;
      39971: inst = 32'hc40539f;
      39972: inst = 32'h8220000;
      39973: inst = 32'h10408000;
      39974: inst = 32'hc4053a0;
      39975: inst = 32'h8220000;
      39976: inst = 32'h10408000;
      39977: inst = 32'hc4053a1;
      39978: inst = 32'h8220000;
      39979: inst = 32'h10408000;
      39980: inst = 32'hc4053a2;
      39981: inst = 32'h8220000;
      39982: inst = 32'h10408000;
      39983: inst = 32'hc4053a3;
      39984: inst = 32'h8220000;
      39985: inst = 32'h10408000;
      39986: inst = 32'hc4053a4;
      39987: inst = 32'h8220000;
      39988: inst = 32'h10408000;
      39989: inst = 32'hc4053a5;
      39990: inst = 32'h8220000;
      39991: inst = 32'h10408000;
      39992: inst = 32'hc4053a6;
      39993: inst = 32'h8220000;
      39994: inst = 32'h10408000;
      39995: inst = 32'hc4053a7;
      39996: inst = 32'h8220000;
      39997: inst = 32'h10408000;
      39998: inst = 32'hc4053a8;
      39999: inst = 32'h8220000;
      40000: inst = 32'h10408000;
      40001: inst = 32'hc4053a9;
      40002: inst = 32'h8220000;
      40003: inst = 32'h10408000;
      40004: inst = 32'hc4053aa;
      40005: inst = 32'h8220000;
      40006: inst = 32'h10408000;
      40007: inst = 32'hc4053ab;
      40008: inst = 32'h8220000;
      40009: inst = 32'h10408000;
      40010: inst = 32'hc4053ac;
      40011: inst = 32'h8220000;
      40012: inst = 32'h10408000;
      40013: inst = 32'hc4053ad;
      40014: inst = 32'h8220000;
      40015: inst = 32'h10408000;
      40016: inst = 32'hc4053ae;
      40017: inst = 32'h8220000;
      40018: inst = 32'h10408000;
      40019: inst = 32'hc4053af;
      40020: inst = 32'h8220000;
      40021: inst = 32'h10408000;
      40022: inst = 32'hc4053b0;
      40023: inst = 32'h8220000;
      40024: inst = 32'h10408000;
      40025: inst = 32'hc4053b1;
      40026: inst = 32'h8220000;
      40027: inst = 32'h10408000;
      40028: inst = 32'hc4053bc;
      40029: inst = 32'h8220000;
      40030: inst = 32'h10408000;
      40031: inst = 32'hc4053c3;
      40032: inst = 32'h8220000;
      40033: inst = 32'h10408000;
      40034: inst = 32'hc4053c4;
      40035: inst = 32'h8220000;
      40036: inst = 32'h10408000;
      40037: inst = 32'hc4053c5;
      40038: inst = 32'h8220000;
      40039: inst = 32'h10408000;
      40040: inst = 32'hc4053c6;
      40041: inst = 32'h8220000;
      40042: inst = 32'h10408000;
      40043: inst = 32'hc4053c7;
      40044: inst = 32'h8220000;
      40045: inst = 32'h10408000;
      40046: inst = 32'hc4053cf;
      40047: inst = 32'h8220000;
      40048: inst = 32'h10408000;
      40049: inst = 32'hc4053d0;
      40050: inst = 32'h8220000;
      40051: inst = 32'h10408000;
      40052: inst = 32'hc4053d1;
      40053: inst = 32'h8220000;
      40054: inst = 32'h10408000;
      40055: inst = 32'hc4053d2;
      40056: inst = 32'h8220000;
      40057: inst = 32'h10408000;
      40058: inst = 32'hc4053d3;
      40059: inst = 32'h8220000;
      40060: inst = 32'h10408000;
      40061: inst = 32'hc4053d4;
      40062: inst = 32'h8220000;
      40063: inst = 32'h10408000;
      40064: inst = 32'hc4053d5;
      40065: inst = 32'h8220000;
      40066: inst = 32'h10408000;
      40067: inst = 32'hc4053d9;
      40068: inst = 32'h8220000;
      40069: inst = 32'h10408000;
      40070: inst = 32'hc4053da;
      40071: inst = 32'h8220000;
      40072: inst = 32'h10408000;
      40073: inst = 32'hc4053db;
      40074: inst = 32'h8220000;
      40075: inst = 32'h10408000;
      40076: inst = 32'hc4053dc;
      40077: inst = 32'h8220000;
      40078: inst = 32'h10408000;
      40079: inst = 32'hc4053dd;
      40080: inst = 32'h8220000;
      40081: inst = 32'h10408000;
      40082: inst = 32'hc4053de;
      40083: inst = 32'h8220000;
      40084: inst = 32'h10408000;
      40085: inst = 32'hc4053df;
      40086: inst = 32'h8220000;
      40087: inst = 32'h10408000;
      40088: inst = 32'hc4053e0;
      40089: inst = 32'h8220000;
      40090: inst = 32'h10408000;
      40091: inst = 32'hc4053e1;
      40092: inst = 32'h8220000;
      40093: inst = 32'h10408000;
      40094: inst = 32'hc4053e2;
      40095: inst = 32'h8220000;
      40096: inst = 32'h10408000;
      40097: inst = 32'hc4053e3;
      40098: inst = 32'h8220000;
      40099: inst = 32'h10408000;
      40100: inst = 32'hc4053e4;
      40101: inst = 32'h8220000;
      40102: inst = 32'h10408000;
      40103: inst = 32'hc4053e5;
      40104: inst = 32'h8220000;
      40105: inst = 32'h10408000;
      40106: inst = 32'hc4053e6;
      40107: inst = 32'h8220000;
      40108: inst = 32'h10408000;
      40109: inst = 32'hc4053e7;
      40110: inst = 32'h8220000;
      40111: inst = 32'h10408000;
      40112: inst = 32'hc4053e8;
      40113: inst = 32'h8220000;
      40114: inst = 32'h10408000;
      40115: inst = 32'hc4053e9;
      40116: inst = 32'h8220000;
      40117: inst = 32'h10408000;
      40118: inst = 32'hc4053ea;
      40119: inst = 32'h8220000;
      40120: inst = 32'h10408000;
      40121: inst = 32'hc4053eb;
      40122: inst = 32'h8220000;
      40123: inst = 32'h10408000;
      40124: inst = 32'hc4053ec;
      40125: inst = 32'h8220000;
      40126: inst = 32'h10408000;
      40127: inst = 32'hc4053ed;
      40128: inst = 32'h8220000;
      40129: inst = 32'h10408000;
      40130: inst = 32'hc4053ee;
      40131: inst = 32'h8220000;
      40132: inst = 32'h10408000;
      40133: inst = 32'hc4053ef;
      40134: inst = 32'h8220000;
      40135: inst = 32'h10408000;
      40136: inst = 32'hc4053f0;
      40137: inst = 32'h8220000;
      40138: inst = 32'h10408000;
      40139: inst = 32'hc4053f1;
      40140: inst = 32'h8220000;
      40141: inst = 32'h10408000;
      40142: inst = 32'hc4053f2;
      40143: inst = 32'h8220000;
      40144: inst = 32'h10408000;
      40145: inst = 32'hc4053f3;
      40146: inst = 32'h8220000;
      40147: inst = 32'h10408000;
      40148: inst = 32'hc4053f4;
      40149: inst = 32'h8220000;
      40150: inst = 32'h10408000;
      40151: inst = 32'hc4053f5;
      40152: inst = 32'h8220000;
      40153: inst = 32'h10408000;
      40154: inst = 32'hc4053f6;
      40155: inst = 32'h8220000;
      40156: inst = 32'h10408000;
      40157: inst = 32'hc4053f7;
      40158: inst = 32'h8220000;
      40159: inst = 32'h10408000;
      40160: inst = 32'hc4053f8;
      40161: inst = 32'h8220000;
      40162: inst = 32'h10408000;
      40163: inst = 32'hc4053f9;
      40164: inst = 32'h8220000;
      40165: inst = 32'h10408000;
      40166: inst = 32'hc4053fa;
      40167: inst = 32'h8220000;
      40168: inst = 32'h10408000;
      40169: inst = 32'hc4053fb;
      40170: inst = 32'h8220000;
      40171: inst = 32'h10408000;
      40172: inst = 32'hc4053fc;
      40173: inst = 32'h8220000;
      40174: inst = 32'h10408000;
      40175: inst = 32'hc4053fd;
      40176: inst = 32'h8220000;
      40177: inst = 32'h10408000;
      40178: inst = 32'hc4053fe;
      40179: inst = 32'h8220000;
      40180: inst = 32'h10408000;
      40181: inst = 32'hc4053ff;
      40182: inst = 32'h8220000;
      40183: inst = 32'h10408000;
      40184: inst = 32'hc405400;
      40185: inst = 32'h8220000;
      40186: inst = 32'h10408000;
      40187: inst = 32'hc405401;
      40188: inst = 32'h8220000;
      40189: inst = 32'h10408000;
      40190: inst = 32'hc405402;
      40191: inst = 32'h8220000;
      40192: inst = 32'h10408000;
      40193: inst = 32'hc405403;
      40194: inst = 32'h8220000;
      40195: inst = 32'h10408000;
      40196: inst = 32'hc405404;
      40197: inst = 32'h8220000;
      40198: inst = 32'h10408000;
      40199: inst = 32'hc405405;
      40200: inst = 32'h8220000;
      40201: inst = 32'h10408000;
      40202: inst = 32'hc405406;
      40203: inst = 32'h8220000;
      40204: inst = 32'h10408000;
      40205: inst = 32'hc405407;
      40206: inst = 32'h8220000;
      40207: inst = 32'h10408000;
      40208: inst = 32'hc405408;
      40209: inst = 32'h8220000;
      40210: inst = 32'h10408000;
      40211: inst = 32'hc405409;
      40212: inst = 32'h8220000;
      40213: inst = 32'h10408000;
      40214: inst = 32'hc40540a;
      40215: inst = 32'h8220000;
      40216: inst = 32'h10408000;
      40217: inst = 32'hc40540b;
      40218: inst = 32'h8220000;
      40219: inst = 32'h10408000;
      40220: inst = 32'hc40540c;
      40221: inst = 32'h8220000;
      40222: inst = 32'h10408000;
      40223: inst = 32'hc40540d;
      40224: inst = 32'h8220000;
      40225: inst = 32'h10408000;
      40226: inst = 32'hc40540e;
      40227: inst = 32'h8220000;
      40228: inst = 32'h10408000;
      40229: inst = 32'hc40540f;
      40230: inst = 32'h8220000;
      40231: inst = 32'h10408000;
      40232: inst = 32'hc405410;
      40233: inst = 32'h8220000;
      40234: inst = 32'h10408000;
      40235: inst = 32'hc405411;
      40236: inst = 32'h8220000;
      40237: inst = 32'h10408000;
      40238: inst = 32'hc40541c;
      40239: inst = 32'h8220000;
      40240: inst = 32'h10408000;
      40241: inst = 32'hc405423;
      40242: inst = 32'h8220000;
      40243: inst = 32'h10408000;
      40244: inst = 32'hc405424;
      40245: inst = 32'h8220000;
      40246: inst = 32'h10408000;
      40247: inst = 32'hc405425;
      40248: inst = 32'h8220000;
      40249: inst = 32'h10408000;
      40250: inst = 32'hc405426;
      40251: inst = 32'h8220000;
      40252: inst = 32'h10408000;
      40253: inst = 32'hc405430;
      40254: inst = 32'h8220000;
      40255: inst = 32'h10408000;
      40256: inst = 32'hc405431;
      40257: inst = 32'h8220000;
      40258: inst = 32'h10408000;
      40259: inst = 32'hc405432;
      40260: inst = 32'h8220000;
      40261: inst = 32'h10408000;
      40262: inst = 32'hc405433;
      40263: inst = 32'h8220000;
      40264: inst = 32'h10408000;
      40265: inst = 32'hc405434;
      40266: inst = 32'h8220000;
      40267: inst = 32'h10408000;
      40268: inst = 32'hc405435;
      40269: inst = 32'h8220000;
      40270: inst = 32'h10408000;
      40271: inst = 32'hc40544a;
      40272: inst = 32'h8220000;
      40273: inst = 32'h10408000;
      40274: inst = 32'hc40544b;
      40275: inst = 32'h8220000;
      40276: inst = 32'h10408000;
      40277: inst = 32'hc40544c;
      40278: inst = 32'h8220000;
      40279: inst = 32'h10408000;
      40280: inst = 32'hc40544d;
      40281: inst = 32'h8220000;
      40282: inst = 32'h10408000;
      40283: inst = 32'hc40544e;
      40284: inst = 32'h8220000;
      40285: inst = 32'h10408000;
      40286: inst = 32'hc40544f;
      40287: inst = 32'h8220000;
      40288: inst = 32'h10408000;
      40289: inst = 32'hc405450;
      40290: inst = 32'h8220000;
      40291: inst = 32'h10408000;
      40292: inst = 32'hc405451;
      40293: inst = 32'h8220000;
      40294: inst = 32'h10408000;
      40295: inst = 32'hc405452;
      40296: inst = 32'h8220000;
      40297: inst = 32'h10408000;
      40298: inst = 32'hc405453;
      40299: inst = 32'h8220000;
      40300: inst = 32'h10408000;
      40301: inst = 32'hc405454;
      40302: inst = 32'h8220000;
      40303: inst = 32'h10408000;
      40304: inst = 32'hc405455;
      40305: inst = 32'h8220000;
      40306: inst = 32'h10408000;
      40307: inst = 32'hc405456;
      40308: inst = 32'h8220000;
      40309: inst = 32'h10408000;
      40310: inst = 32'hc405457;
      40311: inst = 32'h8220000;
      40312: inst = 32'h10408000;
      40313: inst = 32'hc405458;
      40314: inst = 32'h8220000;
      40315: inst = 32'h10408000;
      40316: inst = 32'hc405459;
      40317: inst = 32'h8220000;
      40318: inst = 32'h10408000;
      40319: inst = 32'hc40545a;
      40320: inst = 32'h8220000;
      40321: inst = 32'h10408000;
      40322: inst = 32'hc40545b;
      40323: inst = 32'h8220000;
      40324: inst = 32'h10408000;
      40325: inst = 32'hc40545c;
      40326: inst = 32'h8220000;
      40327: inst = 32'h10408000;
      40328: inst = 32'hc40545d;
      40329: inst = 32'h8220000;
      40330: inst = 32'h10408000;
      40331: inst = 32'hc40545e;
      40332: inst = 32'h8220000;
      40333: inst = 32'h10408000;
      40334: inst = 32'hc40545f;
      40335: inst = 32'h8220000;
      40336: inst = 32'h10408000;
      40337: inst = 32'hc405460;
      40338: inst = 32'h8220000;
      40339: inst = 32'h10408000;
      40340: inst = 32'hc405461;
      40341: inst = 32'h8220000;
      40342: inst = 32'h10408000;
      40343: inst = 32'hc405462;
      40344: inst = 32'h8220000;
      40345: inst = 32'h10408000;
      40346: inst = 32'hc405463;
      40347: inst = 32'h8220000;
      40348: inst = 32'h10408000;
      40349: inst = 32'hc405464;
      40350: inst = 32'h8220000;
      40351: inst = 32'h10408000;
      40352: inst = 32'hc405465;
      40353: inst = 32'h8220000;
      40354: inst = 32'h10408000;
      40355: inst = 32'hc405466;
      40356: inst = 32'h8220000;
      40357: inst = 32'h10408000;
      40358: inst = 32'hc405467;
      40359: inst = 32'h8220000;
      40360: inst = 32'h10408000;
      40361: inst = 32'hc405468;
      40362: inst = 32'h8220000;
      40363: inst = 32'h10408000;
      40364: inst = 32'hc405469;
      40365: inst = 32'h8220000;
      40366: inst = 32'h10408000;
      40367: inst = 32'hc40546a;
      40368: inst = 32'h8220000;
      40369: inst = 32'h10408000;
      40370: inst = 32'hc40546b;
      40371: inst = 32'h8220000;
      40372: inst = 32'h10408000;
      40373: inst = 32'hc40546c;
      40374: inst = 32'h8220000;
      40375: inst = 32'h10408000;
      40376: inst = 32'hc40546d;
      40377: inst = 32'h8220000;
      40378: inst = 32'h10408000;
      40379: inst = 32'hc40546e;
      40380: inst = 32'h8220000;
      40381: inst = 32'h10408000;
      40382: inst = 32'hc40546f;
      40383: inst = 32'h8220000;
      40384: inst = 32'h10408000;
      40385: inst = 32'hc405470;
      40386: inst = 32'h8220000;
      40387: inst = 32'h10408000;
      40388: inst = 32'hc405471;
      40389: inst = 32'h8220000;
      40390: inst = 32'h10408000;
      40391: inst = 32'hc40547c;
      40392: inst = 32'h8220000;
      40393: inst = 32'h10408000;
      40394: inst = 32'hc405483;
      40395: inst = 32'h8220000;
      40396: inst = 32'h10408000;
      40397: inst = 32'hc405484;
      40398: inst = 32'h8220000;
      40399: inst = 32'h10408000;
      40400: inst = 32'hc405485;
      40401: inst = 32'h8220000;
      40402: inst = 32'h10408000;
      40403: inst = 32'hc405486;
      40404: inst = 32'h8220000;
      40405: inst = 32'h10408000;
      40406: inst = 32'hc405490;
      40407: inst = 32'h8220000;
      40408: inst = 32'h10408000;
      40409: inst = 32'hc405491;
      40410: inst = 32'h8220000;
      40411: inst = 32'h10408000;
      40412: inst = 32'hc405492;
      40413: inst = 32'h8220000;
      40414: inst = 32'h10408000;
      40415: inst = 32'hc405493;
      40416: inst = 32'h8220000;
      40417: inst = 32'h10408000;
      40418: inst = 32'hc405494;
      40419: inst = 32'h8220000;
      40420: inst = 32'h10408000;
      40421: inst = 32'hc405495;
      40422: inst = 32'h8220000;
      40423: inst = 32'h10408000;
      40424: inst = 32'hc4054aa;
      40425: inst = 32'h8220000;
      40426: inst = 32'h10408000;
      40427: inst = 32'hc4054ab;
      40428: inst = 32'h8220000;
      40429: inst = 32'h10408000;
      40430: inst = 32'hc4054ac;
      40431: inst = 32'h8220000;
      40432: inst = 32'h10408000;
      40433: inst = 32'hc4054ad;
      40434: inst = 32'h8220000;
      40435: inst = 32'h10408000;
      40436: inst = 32'hc4054ae;
      40437: inst = 32'h8220000;
      40438: inst = 32'h10408000;
      40439: inst = 32'hc4054af;
      40440: inst = 32'h8220000;
      40441: inst = 32'h10408000;
      40442: inst = 32'hc4054b0;
      40443: inst = 32'h8220000;
      40444: inst = 32'h10408000;
      40445: inst = 32'hc4054b1;
      40446: inst = 32'h8220000;
      40447: inst = 32'h10408000;
      40448: inst = 32'hc4054b2;
      40449: inst = 32'h8220000;
      40450: inst = 32'h10408000;
      40451: inst = 32'hc4054b3;
      40452: inst = 32'h8220000;
      40453: inst = 32'h10408000;
      40454: inst = 32'hc4054b4;
      40455: inst = 32'h8220000;
      40456: inst = 32'h10408000;
      40457: inst = 32'hc4054b5;
      40458: inst = 32'h8220000;
      40459: inst = 32'h10408000;
      40460: inst = 32'hc4054b6;
      40461: inst = 32'h8220000;
      40462: inst = 32'h10408000;
      40463: inst = 32'hc4054b7;
      40464: inst = 32'h8220000;
      40465: inst = 32'h10408000;
      40466: inst = 32'hc4054b8;
      40467: inst = 32'h8220000;
      40468: inst = 32'h10408000;
      40469: inst = 32'hc4054b9;
      40470: inst = 32'h8220000;
      40471: inst = 32'h10408000;
      40472: inst = 32'hc4054ba;
      40473: inst = 32'h8220000;
      40474: inst = 32'h10408000;
      40475: inst = 32'hc4054bb;
      40476: inst = 32'h8220000;
      40477: inst = 32'h10408000;
      40478: inst = 32'hc4054bc;
      40479: inst = 32'h8220000;
      40480: inst = 32'h10408000;
      40481: inst = 32'hc4054bd;
      40482: inst = 32'h8220000;
      40483: inst = 32'h10408000;
      40484: inst = 32'hc4054be;
      40485: inst = 32'h8220000;
      40486: inst = 32'h10408000;
      40487: inst = 32'hc4054bf;
      40488: inst = 32'h8220000;
      40489: inst = 32'h10408000;
      40490: inst = 32'hc4054c0;
      40491: inst = 32'h8220000;
      40492: inst = 32'h10408000;
      40493: inst = 32'hc4054c1;
      40494: inst = 32'h8220000;
      40495: inst = 32'h10408000;
      40496: inst = 32'hc4054c2;
      40497: inst = 32'h8220000;
      40498: inst = 32'h10408000;
      40499: inst = 32'hc4054c3;
      40500: inst = 32'h8220000;
      40501: inst = 32'h10408000;
      40502: inst = 32'hc4054c4;
      40503: inst = 32'h8220000;
      40504: inst = 32'h10408000;
      40505: inst = 32'hc4054c5;
      40506: inst = 32'h8220000;
      40507: inst = 32'h10408000;
      40508: inst = 32'hc4054c6;
      40509: inst = 32'h8220000;
      40510: inst = 32'h10408000;
      40511: inst = 32'hc4054c7;
      40512: inst = 32'h8220000;
      40513: inst = 32'h10408000;
      40514: inst = 32'hc4054c8;
      40515: inst = 32'h8220000;
      40516: inst = 32'h10408000;
      40517: inst = 32'hc4054c9;
      40518: inst = 32'h8220000;
      40519: inst = 32'h10408000;
      40520: inst = 32'hc4054ca;
      40521: inst = 32'h8220000;
      40522: inst = 32'h10408000;
      40523: inst = 32'hc4054cb;
      40524: inst = 32'h8220000;
      40525: inst = 32'h10408000;
      40526: inst = 32'hc4054cc;
      40527: inst = 32'h8220000;
      40528: inst = 32'h10408000;
      40529: inst = 32'hc4054cd;
      40530: inst = 32'h8220000;
      40531: inst = 32'h10408000;
      40532: inst = 32'hc4054ce;
      40533: inst = 32'h8220000;
      40534: inst = 32'h10408000;
      40535: inst = 32'hc4054cf;
      40536: inst = 32'h8220000;
      40537: inst = 32'h10408000;
      40538: inst = 32'hc4054d0;
      40539: inst = 32'h8220000;
      40540: inst = 32'h10408000;
      40541: inst = 32'hc4054d1;
      40542: inst = 32'h8220000;
      40543: inst = 32'h10408000;
      40544: inst = 32'hc4054dc;
      40545: inst = 32'h8220000;
      40546: inst = 32'h10408000;
      40547: inst = 32'hc4054e3;
      40548: inst = 32'h8220000;
      40549: inst = 32'h10408000;
      40550: inst = 32'hc4054e4;
      40551: inst = 32'h8220000;
      40552: inst = 32'h10408000;
      40553: inst = 32'hc4054e5;
      40554: inst = 32'h8220000;
      40555: inst = 32'h10408000;
      40556: inst = 32'hc4054e6;
      40557: inst = 32'h8220000;
      40558: inst = 32'h10408000;
      40559: inst = 32'hc4054f0;
      40560: inst = 32'h8220000;
      40561: inst = 32'h10408000;
      40562: inst = 32'hc4054f1;
      40563: inst = 32'h8220000;
      40564: inst = 32'h10408000;
      40565: inst = 32'hc4054f2;
      40566: inst = 32'h8220000;
      40567: inst = 32'h10408000;
      40568: inst = 32'hc4054f3;
      40569: inst = 32'h8220000;
      40570: inst = 32'h10408000;
      40571: inst = 32'hc4054f4;
      40572: inst = 32'h8220000;
      40573: inst = 32'h10408000;
      40574: inst = 32'hc4054f5;
      40575: inst = 32'h8220000;
      40576: inst = 32'h10408000;
      40577: inst = 32'hc40550a;
      40578: inst = 32'h8220000;
      40579: inst = 32'h10408000;
      40580: inst = 32'hc40550b;
      40581: inst = 32'h8220000;
      40582: inst = 32'h10408000;
      40583: inst = 32'hc40550c;
      40584: inst = 32'h8220000;
      40585: inst = 32'h10408000;
      40586: inst = 32'hc40550d;
      40587: inst = 32'h8220000;
      40588: inst = 32'h10408000;
      40589: inst = 32'hc40550e;
      40590: inst = 32'h8220000;
      40591: inst = 32'h10408000;
      40592: inst = 32'hc40550f;
      40593: inst = 32'h8220000;
      40594: inst = 32'h10408000;
      40595: inst = 32'hc405510;
      40596: inst = 32'h8220000;
      40597: inst = 32'h10408000;
      40598: inst = 32'hc405511;
      40599: inst = 32'h8220000;
      40600: inst = 32'h10408000;
      40601: inst = 32'hc405512;
      40602: inst = 32'h8220000;
      40603: inst = 32'h10408000;
      40604: inst = 32'hc405513;
      40605: inst = 32'h8220000;
      40606: inst = 32'h10408000;
      40607: inst = 32'hc405514;
      40608: inst = 32'h8220000;
      40609: inst = 32'h10408000;
      40610: inst = 32'hc405515;
      40611: inst = 32'h8220000;
      40612: inst = 32'h10408000;
      40613: inst = 32'hc405516;
      40614: inst = 32'h8220000;
      40615: inst = 32'h10408000;
      40616: inst = 32'hc405517;
      40617: inst = 32'h8220000;
      40618: inst = 32'h10408000;
      40619: inst = 32'hc405518;
      40620: inst = 32'h8220000;
      40621: inst = 32'h10408000;
      40622: inst = 32'hc405519;
      40623: inst = 32'h8220000;
      40624: inst = 32'h10408000;
      40625: inst = 32'hc40551a;
      40626: inst = 32'h8220000;
      40627: inst = 32'h10408000;
      40628: inst = 32'hc40551b;
      40629: inst = 32'h8220000;
      40630: inst = 32'h10408000;
      40631: inst = 32'hc40551c;
      40632: inst = 32'h8220000;
      40633: inst = 32'h10408000;
      40634: inst = 32'hc40551d;
      40635: inst = 32'h8220000;
      40636: inst = 32'h10408000;
      40637: inst = 32'hc40551e;
      40638: inst = 32'h8220000;
      40639: inst = 32'h10408000;
      40640: inst = 32'hc40551f;
      40641: inst = 32'h8220000;
      40642: inst = 32'h10408000;
      40643: inst = 32'hc405520;
      40644: inst = 32'h8220000;
      40645: inst = 32'h10408000;
      40646: inst = 32'hc405521;
      40647: inst = 32'h8220000;
      40648: inst = 32'h10408000;
      40649: inst = 32'hc405522;
      40650: inst = 32'h8220000;
      40651: inst = 32'h10408000;
      40652: inst = 32'hc405523;
      40653: inst = 32'h8220000;
      40654: inst = 32'h10408000;
      40655: inst = 32'hc405524;
      40656: inst = 32'h8220000;
      40657: inst = 32'h10408000;
      40658: inst = 32'hc405525;
      40659: inst = 32'h8220000;
      40660: inst = 32'h10408000;
      40661: inst = 32'hc405526;
      40662: inst = 32'h8220000;
      40663: inst = 32'h10408000;
      40664: inst = 32'hc405527;
      40665: inst = 32'h8220000;
      40666: inst = 32'h10408000;
      40667: inst = 32'hc405528;
      40668: inst = 32'h8220000;
      40669: inst = 32'h10408000;
      40670: inst = 32'hc405529;
      40671: inst = 32'h8220000;
      40672: inst = 32'h10408000;
      40673: inst = 32'hc40552a;
      40674: inst = 32'h8220000;
      40675: inst = 32'h10408000;
      40676: inst = 32'hc40552b;
      40677: inst = 32'h8220000;
      40678: inst = 32'h10408000;
      40679: inst = 32'hc40552c;
      40680: inst = 32'h8220000;
      40681: inst = 32'h10408000;
      40682: inst = 32'hc40552d;
      40683: inst = 32'h8220000;
      40684: inst = 32'h10408000;
      40685: inst = 32'hc40552e;
      40686: inst = 32'h8220000;
      40687: inst = 32'h10408000;
      40688: inst = 32'hc40552f;
      40689: inst = 32'h8220000;
      40690: inst = 32'h10408000;
      40691: inst = 32'hc405530;
      40692: inst = 32'h8220000;
      40693: inst = 32'h10408000;
      40694: inst = 32'hc405531;
      40695: inst = 32'h8220000;
      40696: inst = 32'h10408000;
      40697: inst = 32'hc40553c;
      40698: inst = 32'h8220000;
      40699: inst = 32'h10408000;
      40700: inst = 32'hc405543;
      40701: inst = 32'h8220000;
      40702: inst = 32'h10408000;
      40703: inst = 32'hc405544;
      40704: inst = 32'h8220000;
      40705: inst = 32'h10408000;
      40706: inst = 32'hc405545;
      40707: inst = 32'h8220000;
      40708: inst = 32'h10408000;
      40709: inst = 32'hc405546;
      40710: inst = 32'h8220000;
      40711: inst = 32'h10408000;
      40712: inst = 32'hc405550;
      40713: inst = 32'h8220000;
      40714: inst = 32'h10408000;
      40715: inst = 32'hc405551;
      40716: inst = 32'h8220000;
      40717: inst = 32'h10408000;
      40718: inst = 32'hc405552;
      40719: inst = 32'h8220000;
      40720: inst = 32'h10408000;
      40721: inst = 32'hc405553;
      40722: inst = 32'h8220000;
      40723: inst = 32'h10408000;
      40724: inst = 32'hc405554;
      40725: inst = 32'h8220000;
      40726: inst = 32'h10408000;
      40727: inst = 32'hc405555;
      40728: inst = 32'h8220000;
      40729: inst = 32'h10408000;
      40730: inst = 32'hc405559;
      40731: inst = 32'h8220000;
      40732: inst = 32'h10408000;
      40733: inst = 32'hc40555a;
      40734: inst = 32'h8220000;
      40735: inst = 32'h10408000;
      40736: inst = 32'hc40555b;
      40737: inst = 32'h8220000;
      40738: inst = 32'h10408000;
      40739: inst = 32'hc40555c;
      40740: inst = 32'h8220000;
      40741: inst = 32'h10408000;
      40742: inst = 32'hc40555d;
      40743: inst = 32'h8220000;
      40744: inst = 32'h10408000;
      40745: inst = 32'hc40555e;
      40746: inst = 32'h8220000;
      40747: inst = 32'h10408000;
      40748: inst = 32'hc40555f;
      40749: inst = 32'h8220000;
      40750: inst = 32'h10408000;
      40751: inst = 32'hc405560;
      40752: inst = 32'h8220000;
      40753: inst = 32'h10408000;
      40754: inst = 32'hc405561;
      40755: inst = 32'h8220000;
      40756: inst = 32'h10408000;
      40757: inst = 32'hc405562;
      40758: inst = 32'h8220000;
      40759: inst = 32'h10408000;
      40760: inst = 32'hc405563;
      40761: inst = 32'h8220000;
      40762: inst = 32'h10408000;
      40763: inst = 32'hc405564;
      40764: inst = 32'h8220000;
      40765: inst = 32'h10408000;
      40766: inst = 32'hc405565;
      40767: inst = 32'h8220000;
      40768: inst = 32'h10408000;
      40769: inst = 32'hc405566;
      40770: inst = 32'h8220000;
      40771: inst = 32'h10408000;
      40772: inst = 32'hc405567;
      40773: inst = 32'h8220000;
      40774: inst = 32'h10408000;
      40775: inst = 32'hc405568;
      40776: inst = 32'h8220000;
      40777: inst = 32'h10408000;
      40778: inst = 32'hc405569;
      40779: inst = 32'h8220000;
      40780: inst = 32'h10408000;
      40781: inst = 32'hc40556a;
      40782: inst = 32'h8220000;
      40783: inst = 32'h10408000;
      40784: inst = 32'hc40556b;
      40785: inst = 32'h8220000;
      40786: inst = 32'h10408000;
      40787: inst = 32'hc40556c;
      40788: inst = 32'h8220000;
      40789: inst = 32'h10408000;
      40790: inst = 32'hc40556d;
      40791: inst = 32'h8220000;
      40792: inst = 32'h10408000;
      40793: inst = 32'hc40556e;
      40794: inst = 32'h8220000;
      40795: inst = 32'h10408000;
      40796: inst = 32'hc40556f;
      40797: inst = 32'h8220000;
      40798: inst = 32'h10408000;
      40799: inst = 32'hc405570;
      40800: inst = 32'h8220000;
      40801: inst = 32'h10408000;
      40802: inst = 32'hc405571;
      40803: inst = 32'h8220000;
      40804: inst = 32'h10408000;
      40805: inst = 32'hc405572;
      40806: inst = 32'h8220000;
      40807: inst = 32'h10408000;
      40808: inst = 32'hc405573;
      40809: inst = 32'h8220000;
      40810: inst = 32'h10408000;
      40811: inst = 32'hc405574;
      40812: inst = 32'h8220000;
      40813: inst = 32'h10408000;
      40814: inst = 32'hc405575;
      40815: inst = 32'h8220000;
      40816: inst = 32'h10408000;
      40817: inst = 32'hc405576;
      40818: inst = 32'h8220000;
      40819: inst = 32'h10408000;
      40820: inst = 32'hc405577;
      40821: inst = 32'h8220000;
      40822: inst = 32'h10408000;
      40823: inst = 32'hc405578;
      40824: inst = 32'h8220000;
      40825: inst = 32'h10408000;
      40826: inst = 32'hc405579;
      40827: inst = 32'h8220000;
      40828: inst = 32'h10408000;
      40829: inst = 32'hc40557a;
      40830: inst = 32'h8220000;
      40831: inst = 32'h10408000;
      40832: inst = 32'hc40557b;
      40833: inst = 32'h8220000;
      40834: inst = 32'h10408000;
      40835: inst = 32'hc40557c;
      40836: inst = 32'h8220000;
      40837: inst = 32'h10408000;
      40838: inst = 32'hc40557d;
      40839: inst = 32'h8220000;
      40840: inst = 32'h10408000;
      40841: inst = 32'hc40557e;
      40842: inst = 32'h8220000;
      40843: inst = 32'h10408000;
      40844: inst = 32'hc40557f;
      40845: inst = 32'h8220000;
      40846: inst = 32'h10408000;
      40847: inst = 32'hc405580;
      40848: inst = 32'h8220000;
      40849: inst = 32'h10408000;
      40850: inst = 32'hc405581;
      40851: inst = 32'h8220000;
      40852: inst = 32'h10408000;
      40853: inst = 32'hc405582;
      40854: inst = 32'h8220000;
      40855: inst = 32'h10408000;
      40856: inst = 32'hc405583;
      40857: inst = 32'h8220000;
      40858: inst = 32'h10408000;
      40859: inst = 32'hc405584;
      40860: inst = 32'h8220000;
      40861: inst = 32'h10408000;
      40862: inst = 32'hc405585;
      40863: inst = 32'h8220000;
      40864: inst = 32'h10408000;
      40865: inst = 32'hc405586;
      40866: inst = 32'h8220000;
      40867: inst = 32'h10408000;
      40868: inst = 32'hc405587;
      40869: inst = 32'h8220000;
      40870: inst = 32'h10408000;
      40871: inst = 32'hc405588;
      40872: inst = 32'h8220000;
      40873: inst = 32'h10408000;
      40874: inst = 32'hc405589;
      40875: inst = 32'h8220000;
      40876: inst = 32'h10408000;
      40877: inst = 32'hc40558a;
      40878: inst = 32'h8220000;
      40879: inst = 32'h10408000;
      40880: inst = 32'hc40558b;
      40881: inst = 32'h8220000;
      40882: inst = 32'h10408000;
      40883: inst = 32'hc40558c;
      40884: inst = 32'h8220000;
      40885: inst = 32'h10408000;
      40886: inst = 32'hc40558d;
      40887: inst = 32'h8220000;
      40888: inst = 32'h10408000;
      40889: inst = 32'hc40558e;
      40890: inst = 32'h8220000;
      40891: inst = 32'h10408000;
      40892: inst = 32'hc40558f;
      40893: inst = 32'h8220000;
      40894: inst = 32'h10408000;
      40895: inst = 32'hc405590;
      40896: inst = 32'h8220000;
      40897: inst = 32'h10408000;
      40898: inst = 32'hc405591;
      40899: inst = 32'h8220000;
      40900: inst = 32'h10408000;
      40901: inst = 32'hc40559c;
      40902: inst = 32'h8220000;
      40903: inst = 32'h10408000;
      40904: inst = 32'hc4055a3;
      40905: inst = 32'h8220000;
      40906: inst = 32'h10408000;
      40907: inst = 32'hc4055a4;
      40908: inst = 32'h8220000;
      40909: inst = 32'h10408000;
      40910: inst = 32'hc4055a5;
      40911: inst = 32'h8220000;
      40912: inst = 32'h10408000;
      40913: inst = 32'hc4055a6;
      40914: inst = 32'h8220000;
      40915: inst = 32'h10408000;
      40916: inst = 32'hc4055b0;
      40917: inst = 32'h8220000;
      40918: inst = 32'h10408000;
      40919: inst = 32'hc4055b1;
      40920: inst = 32'h8220000;
      40921: inst = 32'h10408000;
      40922: inst = 32'hc4055b2;
      40923: inst = 32'h8220000;
      40924: inst = 32'h10408000;
      40925: inst = 32'hc4055b3;
      40926: inst = 32'h8220000;
      40927: inst = 32'h10408000;
      40928: inst = 32'hc4055b4;
      40929: inst = 32'h8220000;
      40930: inst = 32'h10408000;
      40931: inst = 32'hc4055b5;
      40932: inst = 32'h8220000;
      40933: inst = 32'h10408000;
      40934: inst = 32'hc4055b9;
      40935: inst = 32'h8220000;
      40936: inst = 32'h10408000;
      40937: inst = 32'hc4055ba;
      40938: inst = 32'h8220000;
      40939: inst = 32'h10408000;
      40940: inst = 32'hc4055bb;
      40941: inst = 32'h8220000;
      40942: inst = 32'h10408000;
      40943: inst = 32'hc4055bc;
      40944: inst = 32'h8220000;
      40945: inst = 32'h10408000;
      40946: inst = 32'hc4055bd;
      40947: inst = 32'h8220000;
      40948: inst = 32'h10408000;
      40949: inst = 32'hc4055be;
      40950: inst = 32'h8220000;
      40951: inst = 32'h10408000;
      40952: inst = 32'hc4055bf;
      40953: inst = 32'h8220000;
      40954: inst = 32'h10408000;
      40955: inst = 32'hc4055c0;
      40956: inst = 32'h8220000;
      40957: inst = 32'h10408000;
      40958: inst = 32'hc4055c1;
      40959: inst = 32'h8220000;
      40960: inst = 32'h10408000;
      40961: inst = 32'hc4055c2;
      40962: inst = 32'h8220000;
      40963: inst = 32'h10408000;
      40964: inst = 32'hc4055c3;
      40965: inst = 32'h8220000;
      40966: inst = 32'h10408000;
      40967: inst = 32'hc4055c4;
      40968: inst = 32'h8220000;
      40969: inst = 32'h10408000;
      40970: inst = 32'hc4055c5;
      40971: inst = 32'h8220000;
      40972: inst = 32'h10408000;
      40973: inst = 32'hc4055c6;
      40974: inst = 32'h8220000;
      40975: inst = 32'h10408000;
      40976: inst = 32'hc4055c7;
      40977: inst = 32'h8220000;
      40978: inst = 32'h10408000;
      40979: inst = 32'hc4055c8;
      40980: inst = 32'h8220000;
      40981: inst = 32'h10408000;
      40982: inst = 32'hc4055c9;
      40983: inst = 32'h8220000;
      40984: inst = 32'h10408000;
      40985: inst = 32'hc4055ca;
      40986: inst = 32'h8220000;
      40987: inst = 32'h10408000;
      40988: inst = 32'hc4055cb;
      40989: inst = 32'h8220000;
      40990: inst = 32'h10408000;
      40991: inst = 32'hc4055cc;
      40992: inst = 32'h8220000;
      40993: inst = 32'h10408000;
      40994: inst = 32'hc4055cd;
      40995: inst = 32'h8220000;
      40996: inst = 32'h10408000;
      40997: inst = 32'hc4055ce;
      40998: inst = 32'h8220000;
      40999: inst = 32'h10408000;
      41000: inst = 32'hc4055cf;
      41001: inst = 32'h8220000;
      41002: inst = 32'h10408000;
      41003: inst = 32'hc4055d0;
      41004: inst = 32'h8220000;
      41005: inst = 32'h10408000;
      41006: inst = 32'hc4055d1;
      41007: inst = 32'h8220000;
      41008: inst = 32'h10408000;
      41009: inst = 32'hc4055d2;
      41010: inst = 32'h8220000;
      41011: inst = 32'h10408000;
      41012: inst = 32'hc4055d3;
      41013: inst = 32'h8220000;
      41014: inst = 32'h10408000;
      41015: inst = 32'hc4055d4;
      41016: inst = 32'h8220000;
      41017: inst = 32'h10408000;
      41018: inst = 32'hc4055d5;
      41019: inst = 32'h8220000;
      41020: inst = 32'h10408000;
      41021: inst = 32'hc4055d6;
      41022: inst = 32'h8220000;
      41023: inst = 32'h10408000;
      41024: inst = 32'hc4055d7;
      41025: inst = 32'h8220000;
      41026: inst = 32'h10408000;
      41027: inst = 32'hc4055d8;
      41028: inst = 32'h8220000;
      41029: inst = 32'h10408000;
      41030: inst = 32'hc4055d9;
      41031: inst = 32'h8220000;
      41032: inst = 32'h10408000;
      41033: inst = 32'hc4055da;
      41034: inst = 32'h8220000;
      41035: inst = 32'h10408000;
      41036: inst = 32'hc4055db;
      41037: inst = 32'h8220000;
      41038: inst = 32'h10408000;
      41039: inst = 32'hc4055dc;
      41040: inst = 32'h8220000;
      41041: inst = 32'h10408000;
      41042: inst = 32'hc4055dd;
      41043: inst = 32'h8220000;
      41044: inst = 32'h10408000;
      41045: inst = 32'hc4055de;
      41046: inst = 32'h8220000;
      41047: inst = 32'h10408000;
      41048: inst = 32'hc4055df;
      41049: inst = 32'h8220000;
      41050: inst = 32'h10408000;
      41051: inst = 32'hc4055e0;
      41052: inst = 32'h8220000;
      41053: inst = 32'h10408000;
      41054: inst = 32'hc4055e1;
      41055: inst = 32'h8220000;
      41056: inst = 32'h10408000;
      41057: inst = 32'hc4055e2;
      41058: inst = 32'h8220000;
      41059: inst = 32'h10408000;
      41060: inst = 32'hc4055e3;
      41061: inst = 32'h8220000;
      41062: inst = 32'h10408000;
      41063: inst = 32'hc4055e4;
      41064: inst = 32'h8220000;
      41065: inst = 32'h10408000;
      41066: inst = 32'hc4055e5;
      41067: inst = 32'h8220000;
      41068: inst = 32'h10408000;
      41069: inst = 32'hc4055e6;
      41070: inst = 32'h8220000;
      41071: inst = 32'h10408000;
      41072: inst = 32'hc4055e7;
      41073: inst = 32'h8220000;
      41074: inst = 32'h10408000;
      41075: inst = 32'hc4055e8;
      41076: inst = 32'h8220000;
      41077: inst = 32'h10408000;
      41078: inst = 32'hc4055e9;
      41079: inst = 32'h8220000;
      41080: inst = 32'h10408000;
      41081: inst = 32'hc4055ea;
      41082: inst = 32'h8220000;
      41083: inst = 32'h10408000;
      41084: inst = 32'hc4055eb;
      41085: inst = 32'h8220000;
      41086: inst = 32'h10408000;
      41087: inst = 32'hc4055ec;
      41088: inst = 32'h8220000;
      41089: inst = 32'h10408000;
      41090: inst = 32'hc4055ed;
      41091: inst = 32'h8220000;
      41092: inst = 32'h10408000;
      41093: inst = 32'hc4055ee;
      41094: inst = 32'h8220000;
      41095: inst = 32'h10408000;
      41096: inst = 32'hc4055ef;
      41097: inst = 32'h8220000;
      41098: inst = 32'h10408000;
      41099: inst = 32'hc4055f0;
      41100: inst = 32'h8220000;
      41101: inst = 32'h10408000;
      41102: inst = 32'hc4055f1;
      41103: inst = 32'h8220000;
      41104: inst = 32'h10408000;
      41105: inst = 32'hc4055fc;
      41106: inst = 32'h8220000;
      41107: inst = 32'h10408000;
      41108: inst = 32'hc405603;
      41109: inst = 32'h8220000;
      41110: inst = 32'h10408000;
      41111: inst = 32'hc405604;
      41112: inst = 32'h8220000;
      41113: inst = 32'h10408000;
      41114: inst = 32'hc405605;
      41115: inst = 32'h8220000;
      41116: inst = 32'h10408000;
      41117: inst = 32'hc405606;
      41118: inst = 32'h8220000;
      41119: inst = 32'h10408000;
      41120: inst = 32'hc405613;
      41121: inst = 32'h8220000;
      41122: inst = 32'h10408000;
      41123: inst = 32'hc405614;
      41124: inst = 32'h8220000;
      41125: inst = 32'h10408000;
      41126: inst = 32'hc405615;
      41127: inst = 32'h8220000;
      41128: inst = 32'h10408000;
      41129: inst = 32'hc405619;
      41130: inst = 32'h8220000;
      41131: inst = 32'h10408000;
      41132: inst = 32'hc40561a;
      41133: inst = 32'h8220000;
      41134: inst = 32'h10408000;
      41135: inst = 32'hc40561b;
      41136: inst = 32'h8220000;
      41137: inst = 32'h10408000;
      41138: inst = 32'hc40561c;
      41139: inst = 32'h8220000;
      41140: inst = 32'h10408000;
      41141: inst = 32'hc40561d;
      41142: inst = 32'h8220000;
      41143: inst = 32'h10408000;
      41144: inst = 32'hc40561e;
      41145: inst = 32'h8220000;
      41146: inst = 32'h10408000;
      41147: inst = 32'hc40561f;
      41148: inst = 32'h8220000;
      41149: inst = 32'h10408000;
      41150: inst = 32'hc405620;
      41151: inst = 32'h8220000;
      41152: inst = 32'h10408000;
      41153: inst = 32'hc405621;
      41154: inst = 32'h8220000;
      41155: inst = 32'h10408000;
      41156: inst = 32'hc405622;
      41157: inst = 32'h8220000;
      41158: inst = 32'h10408000;
      41159: inst = 32'hc405623;
      41160: inst = 32'h8220000;
      41161: inst = 32'h10408000;
      41162: inst = 32'hc405624;
      41163: inst = 32'h8220000;
      41164: inst = 32'h10408000;
      41165: inst = 32'hc405625;
      41166: inst = 32'h8220000;
      41167: inst = 32'h10408000;
      41168: inst = 32'hc405626;
      41169: inst = 32'h8220000;
      41170: inst = 32'h10408000;
      41171: inst = 32'hc405627;
      41172: inst = 32'h8220000;
      41173: inst = 32'h10408000;
      41174: inst = 32'hc405628;
      41175: inst = 32'h8220000;
      41176: inst = 32'h10408000;
      41177: inst = 32'hc405629;
      41178: inst = 32'h8220000;
      41179: inst = 32'h10408000;
      41180: inst = 32'hc40562a;
      41181: inst = 32'h8220000;
      41182: inst = 32'h10408000;
      41183: inst = 32'hc40562b;
      41184: inst = 32'h8220000;
      41185: inst = 32'h10408000;
      41186: inst = 32'hc40562c;
      41187: inst = 32'h8220000;
      41188: inst = 32'h10408000;
      41189: inst = 32'hc40562d;
      41190: inst = 32'h8220000;
      41191: inst = 32'h10408000;
      41192: inst = 32'hc40562e;
      41193: inst = 32'h8220000;
      41194: inst = 32'h10408000;
      41195: inst = 32'hc40562f;
      41196: inst = 32'h8220000;
      41197: inst = 32'h10408000;
      41198: inst = 32'hc405630;
      41199: inst = 32'h8220000;
      41200: inst = 32'h10408000;
      41201: inst = 32'hc405631;
      41202: inst = 32'h8220000;
      41203: inst = 32'h10408000;
      41204: inst = 32'hc405632;
      41205: inst = 32'h8220000;
      41206: inst = 32'h10408000;
      41207: inst = 32'hc405633;
      41208: inst = 32'h8220000;
      41209: inst = 32'h10408000;
      41210: inst = 32'hc405634;
      41211: inst = 32'h8220000;
      41212: inst = 32'h10408000;
      41213: inst = 32'hc405635;
      41214: inst = 32'h8220000;
      41215: inst = 32'h10408000;
      41216: inst = 32'hc405636;
      41217: inst = 32'h8220000;
      41218: inst = 32'h10408000;
      41219: inst = 32'hc405637;
      41220: inst = 32'h8220000;
      41221: inst = 32'h10408000;
      41222: inst = 32'hc405638;
      41223: inst = 32'h8220000;
      41224: inst = 32'h10408000;
      41225: inst = 32'hc405639;
      41226: inst = 32'h8220000;
      41227: inst = 32'h10408000;
      41228: inst = 32'hc40563a;
      41229: inst = 32'h8220000;
      41230: inst = 32'h10408000;
      41231: inst = 32'hc40563b;
      41232: inst = 32'h8220000;
      41233: inst = 32'h10408000;
      41234: inst = 32'hc40563c;
      41235: inst = 32'h8220000;
      41236: inst = 32'h10408000;
      41237: inst = 32'hc40563d;
      41238: inst = 32'h8220000;
      41239: inst = 32'h10408000;
      41240: inst = 32'hc40563e;
      41241: inst = 32'h8220000;
      41242: inst = 32'h10408000;
      41243: inst = 32'hc40563f;
      41244: inst = 32'h8220000;
      41245: inst = 32'h10408000;
      41246: inst = 32'hc405640;
      41247: inst = 32'h8220000;
      41248: inst = 32'h10408000;
      41249: inst = 32'hc405641;
      41250: inst = 32'h8220000;
      41251: inst = 32'h10408000;
      41252: inst = 32'hc405642;
      41253: inst = 32'h8220000;
      41254: inst = 32'h10408000;
      41255: inst = 32'hc405643;
      41256: inst = 32'h8220000;
      41257: inst = 32'h10408000;
      41258: inst = 32'hc405644;
      41259: inst = 32'h8220000;
      41260: inst = 32'h10408000;
      41261: inst = 32'hc405645;
      41262: inst = 32'h8220000;
      41263: inst = 32'h10408000;
      41264: inst = 32'hc405646;
      41265: inst = 32'h8220000;
      41266: inst = 32'h10408000;
      41267: inst = 32'hc405647;
      41268: inst = 32'h8220000;
      41269: inst = 32'h10408000;
      41270: inst = 32'hc405648;
      41271: inst = 32'h8220000;
      41272: inst = 32'h10408000;
      41273: inst = 32'hc405649;
      41274: inst = 32'h8220000;
      41275: inst = 32'h10408000;
      41276: inst = 32'hc40564a;
      41277: inst = 32'h8220000;
      41278: inst = 32'h10408000;
      41279: inst = 32'hc40564b;
      41280: inst = 32'h8220000;
      41281: inst = 32'h10408000;
      41282: inst = 32'hc40564c;
      41283: inst = 32'h8220000;
      41284: inst = 32'h10408000;
      41285: inst = 32'hc40564d;
      41286: inst = 32'h8220000;
      41287: inst = 32'h10408000;
      41288: inst = 32'hc40564e;
      41289: inst = 32'h8220000;
      41290: inst = 32'h10408000;
      41291: inst = 32'hc40564f;
      41292: inst = 32'h8220000;
      41293: inst = 32'h10408000;
      41294: inst = 32'hc405650;
      41295: inst = 32'h8220000;
      41296: inst = 32'h10408000;
      41297: inst = 32'hc405651;
      41298: inst = 32'h8220000;
      41299: inst = 32'h10408000;
      41300: inst = 32'hc40565c;
      41301: inst = 32'h8220000;
      41302: inst = 32'h10408000;
      41303: inst = 32'hc405663;
      41304: inst = 32'h8220000;
      41305: inst = 32'h10408000;
      41306: inst = 32'hc405664;
      41307: inst = 32'h8220000;
      41308: inst = 32'h10408000;
      41309: inst = 32'hc405665;
      41310: inst = 32'h8220000;
      41311: inst = 32'h10408000;
      41312: inst = 32'hc405666;
      41313: inst = 32'h8220000;
      41314: inst = 32'h10408000;
      41315: inst = 32'hc405667;
      41316: inst = 32'h8220000;
      41317: inst = 32'h10408000;
      41318: inst = 32'hc405674;
      41319: inst = 32'h8220000;
      41320: inst = 32'h10408000;
      41321: inst = 32'hc405675;
      41322: inst = 32'h8220000;
      41323: inst = 32'h10408000;
      41324: inst = 32'hc405679;
      41325: inst = 32'h8220000;
      41326: inst = 32'h10408000;
      41327: inst = 32'hc40567a;
      41328: inst = 32'h8220000;
      41329: inst = 32'h10408000;
      41330: inst = 32'hc40567b;
      41331: inst = 32'h8220000;
      41332: inst = 32'h10408000;
      41333: inst = 32'hc40567c;
      41334: inst = 32'h8220000;
      41335: inst = 32'h10408000;
      41336: inst = 32'hc40567d;
      41337: inst = 32'h8220000;
      41338: inst = 32'h10408000;
      41339: inst = 32'hc40567e;
      41340: inst = 32'h8220000;
      41341: inst = 32'h10408000;
      41342: inst = 32'hc40567f;
      41343: inst = 32'h8220000;
      41344: inst = 32'h10408000;
      41345: inst = 32'hc405680;
      41346: inst = 32'h8220000;
      41347: inst = 32'h10408000;
      41348: inst = 32'hc405681;
      41349: inst = 32'h8220000;
      41350: inst = 32'h10408000;
      41351: inst = 32'hc405682;
      41352: inst = 32'h8220000;
      41353: inst = 32'h10408000;
      41354: inst = 32'hc405683;
      41355: inst = 32'h8220000;
      41356: inst = 32'h10408000;
      41357: inst = 32'hc405684;
      41358: inst = 32'h8220000;
      41359: inst = 32'h10408000;
      41360: inst = 32'hc405685;
      41361: inst = 32'h8220000;
      41362: inst = 32'h10408000;
      41363: inst = 32'hc405686;
      41364: inst = 32'h8220000;
      41365: inst = 32'h10408000;
      41366: inst = 32'hc405687;
      41367: inst = 32'h8220000;
      41368: inst = 32'h10408000;
      41369: inst = 32'hc405688;
      41370: inst = 32'h8220000;
      41371: inst = 32'h10408000;
      41372: inst = 32'hc405689;
      41373: inst = 32'h8220000;
      41374: inst = 32'h10408000;
      41375: inst = 32'hc40568a;
      41376: inst = 32'h8220000;
      41377: inst = 32'h10408000;
      41378: inst = 32'hc40568b;
      41379: inst = 32'h8220000;
      41380: inst = 32'h10408000;
      41381: inst = 32'hc40568c;
      41382: inst = 32'h8220000;
      41383: inst = 32'h10408000;
      41384: inst = 32'hc40568d;
      41385: inst = 32'h8220000;
      41386: inst = 32'h10408000;
      41387: inst = 32'hc40568e;
      41388: inst = 32'h8220000;
      41389: inst = 32'h10408000;
      41390: inst = 32'hc40568f;
      41391: inst = 32'h8220000;
      41392: inst = 32'h10408000;
      41393: inst = 32'hc405690;
      41394: inst = 32'h8220000;
      41395: inst = 32'h10408000;
      41396: inst = 32'hc405691;
      41397: inst = 32'h8220000;
      41398: inst = 32'h10408000;
      41399: inst = 32'hc405692;
      41400: inst = 32'h8220000;
      41401: inst = 32'h10408000;
      41402: inst = 32'hc405693;
      41403: inst = 32'h8220000;
      41404: inst = 32'h10408000;
      41405: inst = 32'hc405694;
      41406: inst = 32'h8220000;
      41407: inst = 32'h10408000;
      41408: inst = 32'hc405695;
      41409: inst = 32'h8220000;
      41410: inst = 32'h10408000;
      41411: inst = 32'hc405696;
      41412: inst = 32'h8220000;
      41413: inst = 32'h10408000;
      41414: inst = 32'hc405697;
      41415: inst = 32'h8220000;
      41416: inst = 32'h10408000;
      41417: inst = 32'hc405698;
      41418: inst = 32'h8220000;
      41419: inst = 32'h10408000;
      41420: inst = 32'hc405699;
      41421: inst = 32'h8220000;
      41422: inst = 32'h10408000;
      41423: inst = 32'hc40569a;
      41424: inst = 32'h8220000;
      41425: inst = 32'h10408000;
      41426: inst = 32'hc40569b;
      41427: inst = 32'h8220000;
      41428: inst = 32'h10408000;
      41429: inst = 32'hc40569c;
      41430: inst = 32'h8220000;
      41431: inst = 32'h10408000;
      41432: inst = 32'hc40569d;
      41433: inst = 32'h8220000;
      41434: inst = 32'h10408000;
      41435: inst = 32'hc40569e;
      41436: inst = 32'h8220000;
      41437: inst = 32'h10408000;
      41438: inst = 32'hc40569f;
      41439: inst = 32'h8220000;
      41440: inst = 32'h10408000;
      41441: inst = 32'hc4056a0;
      41442: inst = 32'h8220000;
      41443: inst = 32'h10408000;
      41444: inst = 32'hc4056a1;
      41445: inst = 32'h8220000;
      41446: inst = 32'h10408000;
      41447: inst = 32'hc4056a2;
      41448: inst = 32'h8220000;
      41449: inst = 32'h10408000;
      41450: inst = 32'hc4056a3;
      41451: inst = 32'h8220000;
      41452: inst = 32'h10408000;
      41453: inst = 32'hc4056a4;
      41454: inst = 32'h8220000;
      41455: inst = 32'h10408000;
      41456: inst = 32'hc4056a5;
      41457: inst = 32'h8220000;
      41458: inst = 32'h10408000;
      41459: inst = 32'hc4056a6;
      41460: inst = 32'h8220000;
      41461: inst = 32'h10408000;
      41462: inst = 32'hc4056a7;
      41463: inst = 32'h8220000;
      41464: inst = 32'h10408000;
      41465: inst = 32'hc4056a8;
      41466: inst = 32'h8220000;
      41467: inst = 32'h10408000;
      41468: inst = 32'hc4056a9;
      41469: inst = 32'h8220000;
      41470: inst = 32'h10408000;
      41471: inst = 32'hc4056aa;
      41472: inst = 32'h8220000;
      41473: inst = 32'h10408000;
      41474: inst = 32'hc4056ab;
      41475: inst = 32'h8220000;
      41476: inst = 32'h10408000;
      41477: inst = 32'hc4056ac;
      41478: inst = 32'h8220000;
      41479: inst = 32'h10408000;
      41480: inst = 32'hc4056ad;
      41481: inst = 32'h8220000;
      41482: inst = 32'h10408000;
      41483: inst = 32'hc4056ae;
      41484: inst = 32'h8220000;
      41485: inst = 32'h10408000;
      41486: inst = 32'hc4056af;
      41487: inst = 32'h8220000;
      41488: inst = 32'h10408000;
      41489: inst = 32'hc4056b0;
      41490: inst = 32'h8220000;
      41491: inst = 32'h10408000;
      41492: inst = 32'hc4056b1;
      41493: inst = 32'h8220000;
      41494: inst = 32'h10408000;
      41495: inst = 32'hc4056bc;
      41496: inst = 32'h8220000;
      41497: inst = 32'h10408000;
      41498: inst = 32'hc405711;
      41499: inst = 32'h8220000;
      41500: inst = 32'h10408000;
      41501: inst = 32'hc40571c;
      41502: inst = 32'h8220000;
      41503: inst = 32'h10408000;
      41504: inst = 32'hc405771;
      41505: inst = 32'h8220000;
      41506: inst = 32'h10408000;
      41507: inst = 32'hc40577c;
      41508: inst = 32'h8220000;
      41509: inst = 32'h10408000;
      41510: inst = 32'hc4057d1;
      41511: inst = 32'h8220000;
      41512: inst = 32'h10408000;
      41513: inst = 32'hc4057dc;
      41514: inst = 32'h8220000;
      41515: inst = 32'hc20cba6;
      41516: inst = 32'h10408000;
      41517: inst = 32'hc403fe4;
      41518: inst = 32'h8220000;
      41519: inst = 32'h10408000;
      41520: inst = 32'hc403fec;
      41521: inst = 32'h8220000;
      41522: inst = 32'h10408000;
      41523: inst = 32'hc4040ac;
      41524: inst = 32'h8220000;
      41525: inst = 32'h10408000;
      41526: inst = 32'hc40410c;
      41527: inst = 32'h8220000;
      41528: inst = 32'h10408000;
      41529: inst = 32'hc40416c;
      41530: inst = 32'h8220000;
      41531: inst = 32'h10408000;
      41532: inst = 32'hc4041c4;
      41533: inst = 32'h8220000;
      41534: inst = 32'h10408000;
      41535: inst = 32'hc404224;
      41536: inst = 32'h8220000;
      41537: inst = 32'h10408000;
      41538: inst = 32'hc404284;
      41539: inst = 32'h8220000;
      41540: inst = 32'h10408000;
      41541: inst = 32'hc40428c;
      41542: inst = 32'h8220000;
      41543: inst = 32'h10408000;
      41544: inst = 32'hc4042e4;
      41545: inst = 32'h8220000;
      41546: inst = 32'h10408000;
      41547: inst = 32'hc4042ec;
      41548: inst = 32'h8220000;
      41549: inst = 32'h10408000;
      41550: inst = 32'hc404344;
      41551: inst = 32'h8220000;
      41552: inst = 32'h10408000;
      41553: inst = 32'hc40434c;
      41554: inst = 32'h8220000;
      41555: inst = 32'h10408000;
      41556: inst = 32'hc4054d2;
      41557: inst = 32'h8220000;
      41558: inst = 32'hc20cb44;
      41559: inst = 32'h10408000;
      41560: inst = 32'hc403fe5;
      41561: inst = 32'h8220000;
      41562: inst = 32'h10408000;
      41563: inst = 32'hc403fe6;
      41564: inst = 32'h8220000;
      41565: inst = 32'h10408000;
      41566: inst = 32'hc403fe7;
      41567: inst = 32'h8220000;
      41568: inst = 32'h10408000;
      41569: inst = 32'hc403fe8;
      41570: inst = 32'h8220000;
      41571: inst = 32'h10408000;
      41572: inst = 32'hc403fe9;
      41573: inst = 32'h8220000;
      41574: inst = 32'h10408000;
      41575: inst = 32'hc403fea;
      41576: inst = 32'h8220000;
      41577: inst = 32'h10408000;
      41578: inst = 32'hc403feb;
      41579: inst = 32'h8220000;
      41580: inst = 32'h10408000;
      41581: inst = 32'hc404104;
      41582: inst = 32'h8220000;
      41583: inst = 32'h10408000;
      41584: inst = 32'hc4043a6;
      41585: inst = 32'h8220000;
      41586: inst = 32'h10408000;
      41587: inst = 32'hc4043a7;
      41588: inst = 32'h8220000;
      41589: inst = 32'h10408000;
      41590: inst = 32'hc4043a8;
      41591: inst = 32'h8220000;
      41592: inst = 32'h10408000;
      41593: inst = 32'hc4043a9;
      41594: inst = 32'h8220000;
      41595: inst = 32'h10408000;
      41596: inst = 32'hc4043aa;
      41597: inst = 32'h8220000;
      41598: inst = 32'h10408000;
      41599: inst = 32'hc4043ab;
      41600: inst = 32'h8220000;
      41601: inst = 32'h10408000;
      41602: inst = 32'hc405354;
      41603: inst = 32'h8220000;
      41604: inst = 32'h10408000;
      41605: inst = 32'hc4053b2;
      41606: inst = 32'h8220000;
      41607: inst = 32'h10408000;
      41608: inst = 32'hc405532;
      41609: inst = 32'h8220000;
      41610: inst = 32'hc20a5f0;
      41611: inst = 32'h10408000;
      41612: inst = 32'hc403fed;
      41613: inst = 32'h8220000;
      41614: inst = 32'hc203d29;
      41615: inst = 32'h10408000;
      41616: inst = 32'hc403fee;
      41617: inst = 32'h8220000;
      41618: inst = 32'hc203ca9;
      41619: inst = 32'h10408000;
      41620: inst = 32'hc403fef;
      41621: inst = 32'h8220000;
      41622: inst = 32'hc20448a;
      41623: inst = 32'h10408000;
      41624: inst = 32'hc403ff0;
      41625: inst = 32'h8220000;
      41626: inst = 32'hc20636f;
      41627: inst = 32'h10408000;
      41628: inst = 32'hc403ff1;
      41629: inst = 32'h8220000;
      41630: inst = 32'h10408000;
      41631: inst = 32'hc403ff7;
      41632: inst = 32'h8220000;
      41633: inst = 32'h10408000;
      41634: inst = 32'hc404053;
      41635: inst = 32'h8220000;
      41636: inst = 32'h10408000;
      41637: inst = 32'hc404675;
      41638: inst = 32'h8220000;
      41639: inst = 32'h10408000;
      41640: inst = 32'hc404677;
      41641: inst = 32'h8220000;
      41642: inst = 32'h10408000;
      41643: inst = 32'hc4046ca;
      41644: inst = 32'h8220000;
      41645: inst = 32'h10408000;
      41646: inst = 32'hc4046d5;
      41647: inst = 32'h8220000;
      41648: inst = 32'h10408000;
      41649: inst = 32'hc404732;
      41650: inst = 32'h8220000;
      41651: inst = 32'hc2053ac;
      41652: inst = 32'h10408000;
      41653: inst = 32'hc403ff2;
      41654: inst = 32'h8220000;
      41655: inst = 32'hc203427;
      41656: inst = 32'h10408000;
      41657: inst = 32'hc403ff3;
      41658: inst = 32'h8220000;
      41659: inst = 32'hc20638f;
      41660: inst = 32'h10408000;
      41661: inst = 32'hc403ff4;
      41662: inst = 32'h8220000;
      41663: inst = 32'hc204bac;
      41664: inst = 32'h10408000;
      41665: inst = 32'hc403ff6;
      41666: inst = 32'h8220000;
      41667: inst = 32'h10408000;
      41668: inst = 32'hc40404e;
      41669: inst = 32'h8220000;
      41670: inst = 32'hc204549;
      41671: inst = 32'h10408000;
      41672: inst = 32'hc403ffa;
      41673: inst = 32'h8220000;
      41674: inst = 32'hc20546c;
      41675: inst = 32'h10408000;
      41676: inst = 32'hc403ffb;
      41677: inst = 32'h8220000;
      41678: inst = 32'hc20544d;
      41679: inst = 32'h10408000;
      41680: inst = 32'hc403ffc;
      41681: inst = 32'h8220000;
      41682: inst = 32'hc20cb86;
      41683: inst = 32'h10408000;
      41684: inst = 32'hc404044;
      41685: inst = 32'h8220000;
      41686: inst = 32'hc20dba5;
      41687: inst = 32'h10408000;
      41688: inst = 32'hc404045;
      41689: inst = 32'h8220000;
      41690: inst = 32'h10408000;
      41691: inst = 32'hc4041c6;
      41692: inst = 32'h8220000;
      41693: inst = 32'h10408000;
      41694: inst = 32'hc4041c7;
      41695: inst = 32'h8220000;
      41696: inst = 32'h10408000;
      41697: inst = 32'hc40428a;
      41698: inst = 32'h8220000;
      41699: inst = 32'h10408000;
      41700: inst = 32'hc404345;
      41701: inst = 32'h8220000;
      41702: inst = 32'h10408000;
      41703: inst = 32'hc4053b4;
      41704: inst = 32'h8220000;
      41705: inst = 32'h10408000;
      41706: inst = 32'hc405713;
      41707: inst = 32'h8220000;
      41708: inst = 32'hc20dbc5;
      41709: inst = 32'h10408000;
      41710: inst = 32'hc404046;
      41711: inst = 32'h8220000;
      41712: inst = 32'h10408000;
      41713: inst = 32'hc404047;
      41714: inst = 32'h8220000;
      41715: inst = 32'h10408000;
      41716: inst = 32'hc4040a9;
      41717: inst = 32'h8220000;
      41718: inst = 32'h10408000;
      41719: inst = 32'hc4040aa;
      41720: inst = 32'h8220000;
      41721: inst = 32'h10408000;
      41722: inst = 32'hc4040ab;
      41723: inst = 32'h8220000;
      41724: inst = 32'h10408000;
      41725: inst = 32'hc404109;
      41726: inst = 32'h8220000;
      41727: inst = 32'h10408000;
      41728: inst = 32'hc40410a;
      41729: inst = 32'h8220000;
      41730: inst = 32'h10408000;
      41731: inst = 32'hc40410b;
      41732: inst = 32'h8220000;
      41733: inst = 32'h10408000;
      41734: inst = 32'hc404169;
      41735: inst = 32'h8220000;
      41736: inst = 32'h10408000;
      41737: inst = 32'hc4041c8;
      41738: inst = 32'h8220000;
      41739: inst = 32'h10408000;
      41740: inst = 32'hc4041c9;
      41741: inst = 32'h8220000;
      41742: inst = 32'h10408000;
      41743: inst = 32'hc404226;
      41744: inst = 32'h8220000;
      41745: inst = 32'h10408000;
      41746: inst = 32'hc404227;
      41747: inst = 32'h8220000;
      41748: inst = 32'h10408000;
      41749: inst = 32'hc404228;
      41750: inst = 32'h8220000;
      41751: inst = 32'h10408000;
      41752: inst = 32'hc404286;
      41753: inst = 32'h8220000;
      41754: inst = 32'h10408000;
      41755: inst = 32'hc404287;
      41756: inst = 32'h8220000;
      41757: inst = 32'h10408000;
      41758: inst = 32'hc404288;
      41759: inst = 32'h8220000;
      41760: inst = 32'h10408000;
      41761: inst = 32'hc404289;
      41762: inst = 32'h8220000;
      41763: inst = 32'h10408000;
      41764: inst = 32'hc4042e6;
      41765: inst = 32'h8220000;
      41766: inst = 32'h10408000;
      41767: inst = 32'hc4042e7;
      41768: inst = 32'h8220000;
      41769: inst = 32'h10408000;
      41770: inst = 32'hc4042e8;
      41771: inst = 32'h8220000;
      41772: inst = 32'h10408000;
      41773: inst = 32'hc4042e9;
      41774: inst = 32'h8220000;
      41775: inst = 32'h10408000;
      41776: inst = 32'hc4042ea;
      41777: inst = 32'h8220000;
      41778: inst = 32'h10408000;
      41779: inst = 32'hc4042eb;
      41780: inst = 32'h8220000;
      41781: inst = 32'h10408000;
      41782: inst = 32'hc405594;
      41783: inst = 32'h8220000;
      41784: inst = 32'h10408000;
      41785: inst = 32'hc4055f4;
      41786: inst = 32'h8220000;
      41787: inst = 32'h10408000;
      41788: inst = 32'hc405653;
      41789: inst = 32'h8220000;
      41790: inst = 32'hc20dbc6;
      41791: inst = 32'h10408000;
      41792: inst = 32'hc404048;
      41793: inst = 32'h8220000;
      41794: inst = 32'h10408000;
      41795: inst = 32'hc404049;
      41796: inst = 32'h8220000;
      41797: inst = 32'h10408000;
      41798: inst = 32'hc40404a;
      41799: inst = 32'h8220000;
      41800: inst = 32'h10408000;
      41801: inst = 32'hc404229;
      41802: inst = 32'h8220000;
      41803: inst = 32'h10408000;
      41804: inst = 32'hc404347;
      41805: inst = 32'h8220000;
      41806: inst = 32'h10408000;
      41807: inst = 32'hc404348;
      41808: inst = 32'h8220000;
      41809: inst = 32'h10408000;
      41810: inst = 32'hc404349;
      41811: inst = 32'h8220000;
      41812: inst = 32'h10408000;
      41813: inst = 32'hc40434a;
      41814: inst = 32'h8220000;
      41815: inst = 32'h10408000;
      41816: inst = 32'hc4055f3;
      41817: inst = 32'h8220000;
      41818: inst = 32'hc20e3c6;
      41819: inst = 32'h10408000;
      41820: inst = 32'hc40404b;
      41821: inst = 32'h8220000;
      41822: inst = 32'h10408000;
      41823: inst = 32'hc404346;
      41824: inst = 32'h8220000;
      41825: inst = 32'h10408000;
      41826: inst = 32'hc40434b;
      41827: inst = 32'h8220000;
      41828: inst = 32'h10408000;
      41829: inst = 32'hc405654;
      41830: inst = 32'h8220000;
      41831: inst = 32'hc20cb85;
      41832: inst = 32'h10408000;
      41833: inst = 32'hc40404c;
      41834: inst = 32'h8220000;
      41835: inst = 32'hc206d0b;
      41836: inst = 32'h10408000;
      41837: inst = 32'hc40404d;
      41838: inst = 32'h8220000;
      41839: inst = 32'hc205c2d;
      41840: inst = 32'h10408000;
      41841: inst = 32'hc40404f;
      41842: inst = 32'h8220000;
      41843: inst = 32'hc203d88;
      41844: inst = 32'h10408000;
      41845: inst = 32'hc404050;
      41846: inst = 32'h8220000;
      41847: inst = 32'hc206b6f;
      41848: inst = 32'h10408000;
      41849: inst = 32'hc404051;
      41850: inst = 32'h8220000;
      41851: inst = 32'h10408000;
      41852: inst = 32'hc40466d;
      41853: inst = 32'h8220000;
      41854: inst = 32'h10408000;
      41855: inst = 32'hc4046d7;
      41856: inst = 32'h8220000;
      41857: inst = 32'h10408000;
      41858: inst = 32'hc40472e;
      41859: inst = 32'h8220000;
      41860: inst = 32'hc206b4f;
      41861: inst = 32'h10408000;
      41862: inst = 32'hc404052;
      41863: inst = 32'h8220000;
      41864: inst = 32'h10408000;
      41865: inst = 32'hc4056b6;
      41866: inst = 32'h8220000;
      41867: inst = 32'hc20542d;
      41868: inst = 32'h10408000;
      41869: inst = 32'hc404055;
      41870: inst = 32'h8220000;
      41871: inst = 32'h10408000;
      41872: inst = 32'hc4040b1;
      41873: inst = 32'h8220000;
      41874: inst = 32'hc205bee;
      41875: inst = 32'h10408000;
      41876: inst = 32'hc404056;
      41877: inst = 32'h8220000;
      41878: inst = 32'h10408000;
      41879: inst = 32'hc4040b5;
      41880: inst = 32'h8220000;
      41881: inst = 32'hc2063af;
      41882: inst = 32'h10408000;
      41883: inst = 32'hc404059;
      41884: inst = 32'h8220000;
      41885: inst = 32'hc203d49;
      41886: inst = 32'h10408000;
      41887: inst = 32'hc40405a;
      41888: inst = 32'h8220000;
      41889: inst = 32'hc206b70;
      41890: inst = 32'h10408000;
      41891: inst = 32'hc40405b;
      41892: inst = 32'h8220000;
      41893: inst = 32'h10408000;
      41894: inst = 32'hc404679;
      41895: inst = 32'h8220000;
      41896: inst = 32'h10408000;
      41897: inst = 32'hc40472d;
      41898: inst = 32'h8220000;
      41899: inst = 32'h10408000;
      41900: inst = 32'hc404730;
      41901: inst = 32'h8220000;
      41902: inst = 32'hc20cb64;
      41903: inst = 32'h10408000;
      41904: inst = 32'hc4040a4;
      41905: inst = 32'h8220000;
      41906: inst = 32'h10408000;
      41907: inst = 32'hc404164;
      41908: inst = 32'h8220000;
      41909: inst = 32'hc20dc08;
      41910: inst = 32'h10408000;
      41911: inst = 32'hc4040a5;
      41912: inst = 32'h8220000;
      41913: inst = 32'hc20f77b;
      41914: inst = 32'h10408000;
      41915: inst = 32'hc4040a6;
      41916: inst = 32'h8220000;
      41917: inst = 32'h10408000;
      41918: inst = 32'hc404154;
      41919: inst = 32'h8220000;
      41920: inst = 32'h10408000;
      41921: inst = 32'hc404155;
      41922: inst = 32'h8220000;
      41923: inst = 32'h10408000;
      41924: inst = 32'hc4041b0;
      41925: inst = 32'h8220000;
      41926: inst = 32'h10408000;
      41927: inst = 32'hc4041b7;
      41928: inst = 32'h8220000;
      41929: inst = 32'h10408000;
      41930: inst = 32'hc404274;
      41931: inst = 32'h8220000;
      41932: inst = 32'h10408000;
      41933: inst = 32'hc40427a;
      41934: inst = 32'h8220000;
      41935: inst = 32'h10408000;
      41936: inst = 32'hc404339;
      41937: inst = 32'h8220000;
      41938: inst = 32'h10408000;
      41939: inst = 32'hc4043fa;
      41940: inst = 32'h8220000;
      41941: inst = 32'h10408000;
      41942: inst = 32'hc404453;
      41943: inst = 32'h8220000;
      41944: inst = 32'h10408000;
      41945: inst = 32'hc404458;
      41946: inst = 32'h8220000;
      41947: inst = 32'h10408000;
      41948: inst = 32'hc4044b6;
      41949: inst = 32'h8220000;
      41950: inst = 32'h10408000;
      41951: inst = 32'hc4044ba;
      41952: inst = 32'h8220000;
      41953: inst = 32'h10408000;
      41954: inst = 32'hc404519;
      41955: inst = 32'h8220000;
      41956: inst = 32'h10408000;
      41957: inst = 32'hc4045d3;
      41958: inst = 32'h8220000;
      41959: inst = 32'hc20e48a;
      41960: inst = 32'h10408000;
      41961: inst = 32'hc4040a7;
      41962: inst = 32'h8220000;
      41963: inst = 32'hc20db84;
      41964: inst = 32'h10408000;
      41965: inst = 32'hc4040a8;
      41966: inst = 32'h8220000;
      41967: inst = 32'h10408000;
      41968: inst = 32'hc404108;
      41969: inst = 32'h8220000;
      41970: inst = 32'h10408000;
      41971: inst = 32'hc404168;
      41972: inst = 32'h8220000;
      41973: inst = 32'hc20a5d0;
      41974: inst = 32'h10408000;
      41975: inst = 32'hc4040ad;
      41976: inst = 32'h8220000;
      41977: inst = 32'h10408000;
      41978: inst = 32'hc404231;
      41979: inst = 32'h8220000;
      41980: inst = 32'h10408000;
      41981: inst = 32'hc404290;
      41982: inst = 32'h8220000;
      41983: inst = 32'hc205b6e;
      41984: inst = 32'h10408000;
      41985: inst = 32'hc4040ae;
      41986: inst = 32'h8220000;
      41987: inst = 32'hc204ccb;
      41988: inst = 32'h10408000;
      41989: inst = 32'hc4040b0;
      41990: inst = 32'h8220000;
      41991: inst = 32'h10408000;
      41992: inst = 32'hc4040ba;
      41993: inst = 32'h8220000;
      41994: inst = 32'hc2043aa;
      41995: inst = 32'h10408000;
      41996: inst = 32'hc4040b3;
      41997: inst = 32'h8220000;
      41998: inst = 32'h10408000;
      41999: inst = 32'hc4040b4;
      42000: inst = 32'h8220000;
      42001: inst = 32'hc2063ae;
      42002: inst = 32'h10408000;
      42003: inst = 32'hc4040b6;
      42004: inst = 32'h8220000;
      42005: inst = 32'h10408000;
      42006: inst = 32'hc40466a;
      42007: inst = 32'h8220000;
      42008: inst = 32'h10408000;
      42009: inst = 32'hc4046cd;
      42010: inst = 32'h8220000;
      42011: inst = 32'hc20544c;
      42012: inst = 32'h10408000;
      42013: inst = 32'hc4040b9;
      42014: inst = 32'h8220000;
      42015: inst = 32'h10408000;
      42016: inst = 32'hc4046cc;
      42017: inst = 32'h8220000;
      42018: inst = 32'h10408000;
      42019: inst = 32'hc40472b;
      42020: inst = 32'h8220000;
      42021: inst = 32'hc20dc28;
      42022: inst = 32'h10408000;
      42023: inst = 32'hc404105;
      42024: inst = 32'h8220000;
      42025: inst = 32'h10408000;
      42026: inst = 32'hc405533;
      42027: inst = 32'h8220000;
      42028: inst = 32'hc20ffff;
      42029: inst = 32'h10408000;
      42030: inst = 32'hc404106;
      42031: inst = 32'h8220000;
      42032: inst = 32'h10408000;
      42033: inst = 32'hc40439b;
      42034: inst = 32'h8220000;
      42035: inst = 32'h10408000;
      42036: inst = 32'hc404515;
      42037: inst = 32'h8220000;
      42038: inst = 32'hc20e4cc;
      42039: inst = 32'h10408000;
      42040: inst = 32'hc404107;
      42041: inst = 32'h8220000;
      42042: inst = 32'h10408000;
      42043: inst = 32'hc404167;
      42044: inst = 32'h8220000;
      42045: inst = 32'hc20ce94;
      42046: inst = 32'h10408000;
      42047: inst = 32'hc40410d;
      42048: inst = 32'h8220000;
      42049: inst = 32'hc20c632;
      42050: inst = 32'h10408000;
      42051: inst = 32'hc404113;
      42052: inst = 32'h8220000;
      42053: inst = 32'hc204ca9;
      42054: inst = 32'h10408000;
      42055: inst = 32'hc404114;
      42056: inst = 32'h8220000;
      42057: inst = 32'hc207e0d;
      42058: inst = 32'h10408000;
      42059: inst = 32'hc404116;
      42060: inst = 32'h8220000;
      42061: inst = 32'hc20d694;
      42062: inst = 32'h10408000;
      42063: inst = 32'hc404117;
      42064: inst = 32'h8220000;
      42065: inst = 32'h10408000;
      42066: inst = 32'hc4047f3;
      42067: inst = 32'h8220000;
      42068: inst = 32'h10408000;
      42069: inst = 32'hc404919;
      42070: inst = 32'h8220000;
      42071: inst = 32'hc20eed7;
      42072: inst = 32'h10408000;
      42073: inst = 32'hc404151;
      42074: inst = 32'h8220000;
      42075: inst = 32'h10408000;
      42076: inst = 32'hc4041b4;
      42077: inst = 32'h8220000;
      42078: inst = 32'h10408000;
      42079: inst = 32'hc404217;
      42080: inst = 32'h8220000;
      42081: inst = 32'h10408000;
      42082: inst = 32'hc404218;
      42083: inst = 32'h8220000;
      42084: inst = 32'h10408000;
      42085: inst = 32'hc404270;
      42086: inst = 32'h8220000;
      42087: inst = 32'h10408000;
      42088: inst = 32'hc404277;
      42089: inst = 32'h8220000;
      42090: inst = 32'h10408000;
      42091: inst = 32'hc4042d0;
      42092: inst = 32'h8220000;
      42093: inst = 32'h10408000;
      42094: inst = 32'hc4042d4;
      42095: inst = 32'h8220000;
      42096: inst = 32'h10408000;
      42097: inst = 32'hc404391;
      42098: inst = 32'h8220000;
      42099: inst = 32'h10408000;
      42100: inst = 32'hc404450;
      42101: inst = 32'h8220000;
      42102: inst = 32'h10408000;
      42103: inst = 32'hc404451;
      42104: inst = 32'h8220000;
      42105: inst = 32'h10408000;
      42106: inst = 32'hc404454;
      42107: inst = 32'h8220000;
      42108: inst = 32'h10408000;
      42109: inst = 32'hc40445b;
      42110: inst = 32'h8220000;
      42111: inst = 32'h10408000;
      42112: inst = 32'hc40451c;
      42113: inst = 32'h8220000;
      42114: inst = 32'h10408000;
      42115: inst = 32'hc4053c8;
      42116: inst = 32'h8220000;
      42117: inst = 32'h10408000;
      42118: inst = 32'hc4053ce;
      42119: inst = 32'h8220000;
      42120: inst = 32'hc20f73a;
      42121: inst = 32'h10408000;
      42122: inst = 32'hc404152;
      42123: inst = 32'h8220000;
      42124: inst = 32'h10408000;
      42125: inst = 32'hc40415b;
      42126: inst = 32'h8220000;
      42127: inst = 32'h10408000;
      42128: inst = 32'hc40415c;
      42129: inst = 32'h8220000;
      42130: inst = 32'h10408000;
      42131: inst = 32'hc40421a;
      42132: inst = 32'h8220000;
      42133: inst = 32'h10408000;
      42134: inst = 32'hc4042d7;
      42135: inst = 32'h8220000;
      42136: inst = 32'h10408000;
      42137: inst = 32'hc4042d8;
      42138: inst = 32'h8220000;
      42139: inst = 32'h10408000;
      42140: inst = 32'hc4042d9;
      42141: inst = 32'h8220000;
      42142: inst = 32'h10408000;
      42143: inst = 32'hc40433b;
      42144: inst = 32'h8220000;
      42145: inst = 32'h10408000;
      42146: inst = 32'hc40439c;
      42147: inst = 32'h8220000;
      42148: inst = 32'h10408000;
      42149: inst = 32'hc4044b3;
      42150: inst = 32'h8220000;
      42151: inst = 32'h10408000;
      42152: inst = 32'hc4044b5;
      42153: inst = 32'h8220000;
      42154: inst = 32'h10408000;
      42155: inst = 32'hc404577;
      42156: inst = 32'h8220000;
      42157: inst = 32'h10408000;
      42158: inst = 32'hc4045d8;
      42159: inst = 32'h8220000;
      42160: inst = 32'h10408000;
      42161: inst = 32'hc4045d9;
      42162: inst = 32'h8220000;
      42163: inst = 32'hc20f75b;
      42164: inst = 32'h10408000;
      42165: inst = 32'hc404153;
      42166: inst = 32'h8220000;
      42167: inst = 32'h10408000;
      42168: inst = 32'hc404157;
      42169: inst = 32'h8220000;
      42170: inst = 32'h10408000;
      42171: inst = 32'hc4041b2;
      42172: inst = 32'h8220000;
      42173: inst = 32'h10408000;
      42174: inst = 32'hc404271;
      42175: inst = 32'h8220000;
      42176: inst = 32'h10408000;
      42177: inst = 32'hc404276;
      42178: inst = 32'h8220000;
      42179: inst = 32'h10408000;
      42180: inst = 32'hc4042dc;
      42181: inst = 32'h8220000;
      42182: inst = 32'h10408000;
      42183: inst = 32'hc404336;
      42184: inst = 32'h8220000;
      42185: inst = 32'h10408000;
      42186: inst = 32'hc404394;
      42187: inst = 32'h8220000;
      42188: inst = 32'h10408000;
      42189: inst = 32'hc4043f0;
      42190: inst = 32'h8220000;
      42191: inst = 32'h10408000;
      42192: inst = 32'hc4043fb;
      42193: inst = 32'h8220000;
      42194: inst = 32'h10408000;
      42195: inst = 32'hc404510;
      42196: inst = 32'h8220000;
      42197: inst = 32'h10408000;
      42198: inst = 32'hc404516;
      42199: inst = 32'h8220000;
      42200: inst = 32'h10408000;
      42201: inst = 32'hc404574;
      42202: inst = 32'h8220000;
      42203: inst = 32'hc20f739;
      42204: inst = 32'h10408000;
      42205: inst = 32'hc404156;
      42206: inst = 32'h8220000;
      42207: inst = 32'h10408000;
      42208: inst = 32'hc4041b6;
      42209: inst = 32'h8220000;
      42210: inst = 32'h10408000;
      42211: inst = 32'hc404213;
      42212: inst = 32'h8220000;
      42213: inst = 32'h10408000;
      42214: inst = 32'hc404399;
      42215: inst = 32'h8220000;
      42216: inst = 32'h10408000;
      42217: inst = 32'hc404517;
      42218: inst = 32'h8220000;
      42219: inst = 32'h10408000;
      42220: inst = 32'hc404576;
      42221: inst = 32'h8220000;
      42222: inst = 32'h10408000;
      42223: inst = 32'hc4045d1;
      42224: inst = 32'h8220000;
      42225: inst = 32'h10408000;
      42226: inst = 32'hc4045dc;
      42227: inst = 32'h8220000;
      42228: inst = 32'hc20ffde;
      42229: inst = 32'h10408000;
      42230: inst = 32'hc404158;
      42231: inst = 32'h8220000;
      42232: inst = 32'h10408000;
      42233: inst = 32'hc4041b9;
      42234: inst = 32'h8220000;
      42235: inst = 32'h10408000;
      42236: inst = 32'hc404392;
      42237: inst = 32'h8220000;
      42238: inst = 32'h10408000;
      42239: inst = 32'hc4043f2;
      42240: inst = 32'h8220000;
      42241: inst = 32'h10408000;
      42242: inst = 32'hc4043f7;
      42243: inst = 32'h8220000;
      42244: inst = 32'h10408000;
      42245: inst = 32'hc4044b9;
      42246: inst = 32'h8220000;
      42247: inst = 32'hc20f75a;
      42248: inst = 32'h10408000;
      42249: inst = 32'hc404159;
      42250: inst = 32'h8220000;
      42251: inst = 32'h10408000;
      42252: inst = 32'hc40415a;
      42253: inst = 32'h8220000;
      42254: inst = 32'h10408000;
      42255: inst = 32'hc404272;
      42256: inst = 32'h8220000;
      42257: inst = 32'h10408000;
      42258: inst = 32'hc404273;
      42259: inst = 32'h8220000;
      42260: inst = 32'h10408000;
      42261: inst = 32'hc404331;
      42262: inst = 32'h8220000;
      42263: inst = 32'h10408000;
      42264: inst = 32'hc4043f3;
      42265: inst = 32'h8220000;
      42266: inst = 32'h10408000;
      42267: inst = 32'hc4043fc;
      42268: inst = 32'h8220000;
      42269: inst = 32'h10408000;
      42270: inst = 32'hc404452;
      42271: inst = 32'h8220000;
      42272: inst = 32'h10408000;
      42273: inst = 32'hc404456;
      42274: inst = 32'h8220000;
      42275: inst = 32'h10408000;
      42276: inst = 32'hc404459;
      42277: inst = 32'h8220000;
      42278: inst = 32'h10408000;
      42279: inst = 32'hc40445a;
      42280: inst = 32'h8220000;
      42281: inst = 32'h10408000;
      42282: inst = 32'hc4044bb;
      42283: inst = 32'h8220000;
      42284: inst = 32'h10408000;
      42285: inst = 32'hc40451a;
      42286: inst = 32'h8220000;
      42287: inst = 32'h10408000;
      42288: inst = 32'hc404570;
      42289: inst = 32'h8220000;
      42290: inst = 32'h10408000;
      42291: inst = 32'hc404573;
      42292: inst = 32'h8220000;
      42293: inst = 32'hc20dbe7;
      42294: inst = 32'h10408000;
      42295: inst = 32'hc404165;
      42296: inst = 32'h8220000;
      42297: inst = 32'hc20f77c;
      42298: inst = 32'h10408000;
      42299: inst = 32'hc404166;
      42300: inst = 32'h8220000;
      42301: inst = 32'h10408000;
      42302: inst = 32'hc4041b8;
      42303: inst = 32'h8220000;
      42304: inst = 32'hc20e3a4;
      42305: inst = 32'h10408000;
      42306: inst = 32'hc40416a;
      42307: inst = 32'h8220000;
      42308: inst = 32'h10408000;
      42309: inst = 32'hc405415;
      42310: inst = 32'h8220000;
      42311: inst = 32'h10408000;
      42312: inst = 32'hc405534;
      42313: inst = 32'h8220000;
      42314: inst = 32'h10408000;
      42315: inst = 32'hc405655;
      42316: inst = 32'h8220000;
      42317: inst = 32'hc20e3c5;
      42318: inst = 32'h10408000;
      42319: inst = 32'hc40416b;
      42320: inst = 32'h8220000;
      42321: inst = 32'h10408000;
      42322: inst = 32'hc40428b;
      42323: inst = 32'h8220000;
      42324: inst = 32'h10408000;
      42325: inst = 32'hc4053b5;
      42326: inst = 32'h8220000;
      42327: inst = 32'h10408000;
      42328: inst = 32'hc405595;
      42329: inst = 32'h8220000;
      42330: inst = 32'h10408000;
      42331: inst = 32'hc4055f5;
      42332: inst = 32'h8220000;
      42333: inst = 32'hc206e0c;
      42334: inst = 32'h10408000;
      42335: inst = 32'hc40416d;
      42336: inst = 32'h8220000;
      42337: inst = 32'hc209e50;
      42338: inst = 32'h10408000;
      42339: inst = 32'hc404176;
      42340: inst = 32'h8220000;
      42341: inst = 32'hc20860e;
      42342: inst = 32'h10408000;
      42343: inst = 32'hc404177;
      42344: inst = 32'h8220000;
      42345: inst = 32'hc20b5f1;
      42346: inst = 32'h10408000;
      42347: inst = 32'hc40417b;
      42348: inst = 32'h8220000;
      42349: inst = 32'hc20ffbd;
      42350: inst = 32'h10408000;
      42351: inst = 32'hc4041b1;
      42352: inst = 32'h8220000;
      42353: inst = 32'h10408000;
      42354: inst = 32'hc404279;
      42355: inst = 32'h8220000;
      42356: inst = 32'h10408000;
      42357: inst = 32'hc404332;
      42358: inst = 32'h8220000;
      42359: inst = 32'h10408000;
      42360: inst = 32'hc404396;
      42361: inst = 32'h8220000;
      42362: inst = 32'h10408000;
      42363: inst = 32'hc404457;
      42364: inst = 32'h8220000;
      42365: inst = 32'h10408000;
      42366: inst = 32'hc40445c;
      42367: inst = 32'h8220000;
      42368: inst = 32'h10408000;
      42369: inst = 32'hc4044bc;
      42370: inst = 32'h8220000;
      42371: inst = 32'hc20f6f8;
      42372: inst = 32'h10408000;
      42373: inst = 32'hc4041b3;
      42374: inst = 32'h8220000;
      42375: inst = 32'h10408000;
      42376: inst = 32'hc404215;
      42377: inst = 32'h8220000;
      42378: inst = 32'h10408000;
      42379: inst = 32'hc40421b;
      42380: inst = 32'h8220000;
      42381: inst = 32'h10408000;
      42382: inst = 32'hc4043f5;
      42383: inst = 32'h8220000;
      42384: inst = 32'h10408000;
      42385: inst = 32'hc4043f8;
      42386: inst = 32'h8220000;
      42387: inst = 32'h10408000;
      42388: inst = 32'hc404572;
      42389: inst = 32'h8220000;
      42390: inst = 32'hc20f719;
      42391: inst = 32'h10408000;
      42392: inst = 32'hc4041ba;
      42393: inst = 32'h8220000;
      42394: inst = 32'h10408000;
      42395: inst = 32'hc4041bb;
      42396: inst = 32'h8220000;
      42397: inst = 32'h10408000;
      42398: inst = 32'hc404335;
      42399: inst = 32'h8220000;
      42400: inst = 32'h10408000;
      42401: inst = 32'hc404337;
      42402: inst = 32'h8220000;
      42403: inst = 32'h10408000;
      42404: inst = 32'hc40433a;
      42405: inst = 32'h8220000;
      42406: inst = 32'h10408000;
      42407: inst = 32'hc404393;
      42408: inst = 32'h8220000;
      42409: inst = 32'h10408000;
      42410: inst = 32'hc4043f4;
      42411: inst = 32'h8220000;
      42412: inst = 32'h10408000;
      42413: inst = 32'hc4044b8;
      42414: inst = 32'h8220000;
      42415: inst = 32'h10408000;
      42416: inst = 32'hc404511;
      42417: inst = 32'h8220000;
      42418: inst = 32'h10408000;
      42419: inst = 32'hc404518;
      42420: inst = 32'h8220000;
      42421: inst = 32'h10408000;
      42422: inst = 32'hc40451b;
      42423: inst = 32'h8220000;
      42424: inst = 32'h10408000;
      42425: inst = 32'hc404575;
      42426: inst = 32'h8220000;
      42427: inst = 32'hc20ffbe;
      42428: inst = 32'h10408000;
      42429: inst = 32'hc4041bc;
      42430: inst = 32'h8220000;
      42431: inst = 32'h10408000;
      42432: inst = 32'hc404275;
      42433: inst = 32'h8220000;
      42434: inst = 32'hc20db85;
      42435: inst = 32'h10408000;
      42436: inst = 32'hc4041c5;
      42437: inst = 32'h8220000;
      42438: inst = 32'h10408000;
      42439: inst = 32'hc404225;
      42440: inst = 32'h8220000;
      42441: inst = 32'h10408000;
      42442: inst = 32'hc404285;
      42443: inst = 32'h8220000;
      42444: inst = 32'h10408000;
      42445: inst = 32'hc4042e5;
      42446: inst = 32'h8220000;
      42447: inst = 32'hc20c44c;
      42448: inst = 32'h10408000;
      42449: inst = 32'hc4041ca;
      42450: inst = 32'h8220000;
      42451: inst = 32'hc20cbe8;
      42452: inst = 32'h10408000;
      42453: inst = 32'hc4041cb;
      42454: inst = 32'h8220000;
      42455: inst = 32'hc20cba5;
      42456: inst = 32'h10408000;
      42457: inst = 32'hc4041cc;
      42458: inst = 32'h8220000;
      42459: inst = 32'h10408000;
      42460: inst = 32'hc40422c;
      42461: inst = 32'h8220000;
      42462: inst = 32'hc20c633;
      42463: inst = 32'h10408000;
      42464: inst = 32'hc4041d0;
      42465: inst = 32'h8220000;
      42466: inst = 32'hc205cca;
      42467: inst = 32'h10408000;
      42468: inst = 32'hc4041d1;
      42469: inst = 32'h8220000;
      42470: inst = 32'hc20e6b6;
      42471: inst = 32'h10408000;
      42472: inst = 32'hc4041d6;
      42473: inst = 32'h8220000;
      42474: inst = 32'h10408000;
      42475: inst = 32'hc40478f;
      42476: inst = 32'h8220000;
      42477: inst = 32'h10408000;
      42478: inst = 32'hc4047eb;
      42479: inst = 32'h8220000;
      42480: inst = 32'h10408000;
      42481: inst = 32'hc4047f2;
      42482: inst = 32'h8220000;
      42483: inst = 32'h10408000;
      42484: inst = 32'hc4048b6;
      42485: inst = 32'h8220000;
      42486: inst = 32'hc2055ca;
      42487: inst = 32'h10408000;
      42488: inst = 32'hc4041d7;
      42489: inst = 32'h8220000;
      42490: inst = 32'hc20de95;
      42491: inst = 32'h10408000;
      42492: inst = 32'hc4041d8;
      42493: inst = 32'h8220000;
      42494: inst = 32'h10408000;
      42495: inst = 32'hc40429b;
      42496: inst = 32'h8220000;
      42497: inst = 32'h10408000;
      42498: inst = 32'hc404792;
      42499: inst = 32'h8220000;
      42500: inst = 32'h10408000;
      42501: inst = 32'hc404798;
      42502: inst = 32'h8220000;
      42503: inst = 32'h10408000;
      42504: inst = 32'hc4047f5;
      42505: inst = 32'h8220000;
      42506: inst = 32'h10408000;
      42507: inst = 32'hc404857;
      42508: inst = 32'h8220000;
      42509: inst = 32'h10408000;
      42510: inst = 32'hc404915;
      42511: inst = 32'h8220000;
      42512: inst = 32'hc2054c9;
      42513: inst = 32'h10408000;
      42514: inst = 32'hc4041db;
      42515: inst = 32'h8220000;
      42516: inst = 32'h10408000;
      42517: inst = 32'hc404230;
      42518: inst = 32'h8220000;
      42519: inst = 32'hc20de75;
      42520: inst = 32'h10408000;
      42521: inst = 32'hc4041dc;
      42522: inst = 32'h8220000;
      42523: inst = 32'hc20f718;
      42524: inst = 32'h10408000;
      42525: inst = 32'hc404210;
      42526: inst = 32'h8220000;
      42527: inst = 32'h10408000;
      42528: inst = 32'hc404278;
      42529: inst = 32'h8220000;
      42530: inst = 32'hc20ff9d;
      42531: inst = 32'h10408000;
      42532: inst = 32'hc404211;
      42533: inst = 32'h8220000;
      42534: inst = 32'h10408000;
      42535: inst = 32'hc404219;
      42536: inst = 32'h8220000;
      42537: inst = 32'h10408000;
      42538: inst = 32'hc4042d6;
      42539: inst = 32'h8220000;
      42540: inst = 32'hc20ff9c;
      42541: inst = 32'h10408000;
      42542: inst = 32'hc404212;
      42543: inst = 32'h8220000;
      42544: inst = 32'h10408000;
      42545: inst = 32'hc404216;
      42546: inst = 32'h8220000;
      42547: inst = 32'h10408000;
      42548: inst = 32'hc40421c;
      42549: inst = 32'h8220000;
      42550: inst = 32'h10408000;
      42551: inst = 32'hc40427b;
      42552: inst = 32'h8220000;
      42553: inst = 32'h10408000;
      42554: inst = 32'hc4042d1;
      42555: inst = 32'h8220000;
      42556: inst = 32'h10408000;
      42557: inst = 32'hc4042d5;
      42558: inst = 32'h8220000;
      42559: inst = 32'h10408000;
      42560: inst = 32'hc40433c;
      42561: inst = 32'h8220000;
      42562: inst = 32'h10408000;
      42563: inst = 32'hc404395;
      42564: inst = 32'h8220000;
      42565: inst = 32'h10408000;
      42566: inst = 32'hc404397;
      42567: inst = 32'h8220000;
      42568: inst = 32'h10408000;
      42569: inst = 32'hc404398;
      42570: inst = 32'h8220000;
      42571: inst = 32'h10408000;
      42572: inst = 32'hc40439a;
      42573: inst = 32'h8220000;
      42574: inst = 32'h10408000;
      42575: inst = 32'hc4043f1;
      42576: inst = 32'h8220000;
      42577: inst = 32'h10408000;
      42578: inst = 32'hc404514;
      42579: inst = 32'h8220000;
      42580: inst = 32'h10408000;
      42581: inst = 32'hc4045d2;
      42582: inst = 32'h8220000;
      42583: inst = 32'hc20a46f;
      42584: inst = 32'h10408000;
      42585: inst = 32'hc40422a;
      42586: inst = 32'h8220000;
      42587: inst = 32'hc20d3c7;
      42588: inst = 32'h10408000;
      42589: inst = 32'hc40422b;
      42590: inst = 32'h8220000;
      42591: inst = 32'h10408000;
      42592: inst = 32'hc405475;
      42593: inst = 32'h8220000;
      42594: inst = 32'hc20ce53;
      42595: inst = 32'h10408000;
      42596: inst = 32'hc40422f;
      42597: inst = 32'h8220000;
      42598: inst = 32'hc207d4d;
      42599: inst = 32'h10408000;
      42600: inst = 32'hc40423b;
      42601: inst = 32'h8220000;
      42602: inst = 32'h10408000;
      42603: inst = 32'hc40423c;
      42604: inst = 32'h8220000;
      42605: inst = 32'hc20ff7c;
      42606: inst = 32'h10408000;
      42607: inst = 32'hc40427c;
      42608: inst = 32'h8220000;
      42609: inst = 32'h10408000;
      42610: inst = 32'hc4042d2;
      42611: inst = 32'h8220000;
      42612: inst = 32'h10408000;
      42613: inst = 32'hc404338;
      42614: inst = 32'h8220000;
      42615: inst = 32'h10408000;
      42616: inst = 32'hc4043f6;
      42617: inst = 32'h8220000;
      42618: inst = 32'h10408000;
      42619: inst = 32'hc4044b4;
      42620: inst = 32'h8220000;
      42621: inst = 32'h10408000;
      42622: inst = 32'hc404571;
      42623: inst = 32'h8220000;
      42624: inst = 32'h10408000;
      42625: inst = 32'hc404578;
      42626: inst = 32'h8220000;
      42627: inst = 32'h10408000;
      42628: inst = 32'hc404579;
      42629: inst = 32'h8220000;
      42630: inst = 32'hc20be12;
      42631: inst = 32'h10408000;
      42632: inst = 32'hc40428f;
      42633: inst = 32'h8220000;
      42634: inst = 32'hc209db0;
      42635: inst = 32'h10408000;
      42636: inst = 32'hc40429c;
      42637: inst = 32'h8220000;
      42638: inst = 32'hc20cb65;
      42639: inst = 32'h10408000;
      42640: inst = 32'hc4043a4;
      42641: inst = 32'h8220000;
      42642: inst = 32'h10408000;
      42643: inst = 32'hc4043ac;
      42644: inst = 32'h8220000;
      42645: inst = 32'hc20cb43;
      42646: inst = 32'h10408000;
      42647: inst = 32'hc4043a5;
      42648: inst = 32'h8220000;
      42649: inst = 32'h10408000;
      42650: inst = 32'hc405355;
      42651: inst = 32'h8220000;
      42652: inst = 32'h10408000;
      42653: inst = 32'hc405712;
      42654: inst = 32'h8220000;
      42655: inst = 32'hc205bce;
      42656: inst = 32'h10408000;
      42657: inst = 32'hc40466b;
      42658: inst = 32'h8220000;
      42659: inst = 32'h10408000;
      42660: inst = 32'hc404670;
      42661: inst = 32'h8220000;
      42662: inst = 32'h10408000;
      42663: inst = 32'hc404674;
      42664: inst = 32'h8220000;
      42665: inst = 32'h10408000;
      42666: inst = 32'hc4046d2;
      42667: inst = 32'h8220000;
      42668: inst = 32'h10408000;
      42669: inst = 32'hc404735;
      42670: inst = 32'h8220000;
      42671: inst = 32'h10408000;
      42672: inst = 32'hc404739;
      42673: inst = 32'h8220000;
      42674: inst = 32'hc205c2c;
      42675: inst = 32'h10408000;
      42676: inst = 32'hc40466c;
      42677: inst = 32'h8220000;
      42678: inst = 32'hc2063ce;
      42679: inst = 32'h10408000;
      42680: inst = 32'hc404671;
      42681: inst = 32'h8220000;
      42682: inst = 32'hc205bed;
      42683: inst = 32'h10408000;
      42684: inst = 32'hc404672;
      42685: inst = 32'h8220000;
      42686: inst = 32'h10408000;
      42687: inst = 32'hc404678;
      42688: inst = 32'h8220000;
      42689: inst = 32'h10408000;
      42690: inst = 32'hc4046d3;
      42691: inst = 32'h8220000;
      42692: inst = 32'h10408000;
      42693: inst = 32'hc4046d8;
      42694: inst = 32'h8220000;
      42695: inst = 32'h10408000;
      42696: inst = 32'hc404733;
      42697: inst = 32'h8220000;
      42698: inst = 32'hc204c8a;
      42699: inst = 32'h10408000;
      42700: inst = 32'hc4046cb;
      42701: inst = 32'h8220000;
      42702: inst = 32'h10408000;
      42703: inst = 32'hc404734;
      42704: inst = 32'h8220000;
      42705: inst = 32'hc20542c;
      42706: inst = 32'h10408000;
      42707: inst = 32'hc4046d4;
      42708: inst = 32'h8220000;
      42709: inst = 32'h10408000;
      42710: inst = 32'hc40472c;
      42711: inst = 32'h8220000;
      42712: inst = 32'hc205c0d;
      42713: inst = 32'h10408000;
      42714: inst = 32'hc4046d9;
      42715: inst = 32'h8220000;
      42716: inst = 32'h10408000;
      42717: inst = 32'hc404731;
      42718: inst = 32'h8220000;
      42719: inst = 32'hc20e6b5;
      42720: inst = 32'h10408000;
      42721: inst = 32'hc40478b;
      42722: inst = 32'h8220000;
      42723: inst = 32'h10408000;
      42724: inst = 32'hc4048b9;
      42725: inst = 32'h8220000;
      42726: inst = 32'hc20ae51;
      42727: inst = 32'h10408000;
      42728: inst = 32'hc40478c;
      42729: inst = 32'h8220000;
      42730: inst = 32'hc20960e;
      42731: inst = 32'h10408000;
      42732: inst = 32'hc40478d;
      42733: inst = 32'h8220000;
      42734: inst = 32'hc20c673;
      42735: inst = 32'h10408000;
      42736: inst = 32'hc40478e;
      42737: inst = 32'h8220000;
      42738: inst = 32'h10408000;
      42739: inst = 32'hc404793;
      42740: inst = 32'h8220000;
      42741: inst = 32'h10408000;
      42742: inst = 32'hc404854;
      42743: inst = 32'h8220000;
      42744: inst = 32'hc20be52;
      42745: inst = 32'h10408000;
      42746: inst = 32'hc404790;
      42747: inst = 32'h8220000;
      42748: inst = 32'h10408000;
      42749: inst = 32'hc404858;
      42750: inst = 32'h8220000;
      42751: inst = 32'h10408000;
      42752: inst = 32'hc404859;
      42753: inst = 32'h8220000;
      42754: inst = 32'hc209e2f;
      42755: inst = 32'h10408000;
      42756: inst = 32'hc404791;
      42757: inst = 32'h8220000;
      42758: inst = 32'h10408000;
      42759: inst = 32'hc404794;
      42760: inst = 32'h8220000;
      42761: inst = 32'hc20ae30;
      42762: inst = 32'h10408000;
      42763: inst = 32'hc4047ec;
      42764: inst = 32'h8220000;
      42765: inst = 32'h10408000;
      42766: inst = 32'hc4047f1;
      42767: inst = 32'h8220000;
      42768: inst = 32'hc20ce73;
      42769: inst = 32'h10408000;
      42770: inst = 32'hc4047ed;
      42771: inst = 32'h8220000;
      42772: inst = 32'h10408000;
      42773: inst = 32'hc4048b4;
      42774: inst = 32'h8220000;
      42775: inst = 32'hc208e0e;
      42776: inst = 32'h10408000;
      42777: inst = 32'hc4047f0;
      42778: inst = 32'h8220000;
      42779: inst = 32'h10408000;
      42780: inst = 32'hc404855;
      42781: inst = 32'h8220000;
      42782: inst = 32'hc2085ed;
      42783: inst = 32'h10408000;
      42784: inst = 32'hc4047f4;
      42785: inst = 32'h8220000;
      42786: inst = 32'h10408000;
      42787: inst = 32'hc4048b8;
      42788: inst = 32'h8220000;
      42789: inst = 32'hc20b651;
      42790: inst = 32'h10408000;
      42791: inst = 32'hc4047f8;
      42792: inst = 32'h8220000;
      42793: inst = 32'h10408000;
      42794: inst = 32'hc404914;
      42795: inst = 32'h8220000;
      42796: inst = 32'hc20c672;
      42797: inst = 32'h10408000;
      42798: inst = 32'hc4047f9;
      42799: inst = 32'h8220000;
      42800: inst = 32'h10408000;
      42801: inst = 32'hc404856;
      42802: inst = 32'h8220000;
      42803: inst = 32'h10408000;
      42804: inst = 32'hc4048b7;
      42805: inst = 32'h8220000;
      42806: inst = 32'hc209e0f;
      42807: inst = 32'h10408000;
      42808: inst = 32'hc4048b5;
      42809: inst = 32'h8220000;
      42810: inst = 32'h10408000;
      42811: inst = 32'hc404918;
      42812: inst = 32'h8220000;
      42813: inst = 32'hc20de94;
      42814: inst = 32'h10408000;
      42815: inst = 32'hc404917;
      42816: inst = 32'h8220000;
      42817: inst = 32'hc20c2e2;
      42818: inst = 32'h10408000;
      42819: inst = 32'hc405352;
      42820: inst = 32'h8220000;
      42821: inst = 32'hc20cb23;
      42822: inst = 32'h10408000;
      42823: inst = 32'hc405353;
      42824: inst = 32'h8220000;
      42825: inst = 32'h10408000;
      42826: inst = 32'hc405356;
      42827: inst = 32'h8220000;
      42828: inst = 32'h10408000;
      42829: inst = 32'hc405357;
      42830: inst = 32'h8220000;
      42831: inst = 32'h10408000;
      42832: inst = 32'hc405358;
      42833: inst = 32'h8220000;
      42834: inst = 32'h10408000;
      42835: inst = 32'hc405359;
      42836: inst = 32'h8220000;
      42837: inst = 32'h10408000;
      42838: inst = 32'hc40535a;
      42839: inst = 32'h8220000;
      42840: inst = 32'h10408000;
      42841: inst = 32'hc405592;
      42842: inst = 32'h8220000;
      42843: inst = 32'h10408000;
      42844: inst = 32'hc4055f2;
      42845: inst = 32'h8220000;
      42846: inst = 32'h10408000;
      42847: inst = 32'hc405652;
      42848: inst = 32'h8220000;
      42849: inst = 32'h10408000;
      42850: inst = 32'hc4056b2;
      42851: inst = 32'h8220000;
      42852: inst = 32'hc20c323;
      42853: inst = 32'h10408000;
      42854: inst = 32'hc40535b;
      42855: inst = 32'h8220000;
      42856: inst = 32'h10408000;
      42857: inst = 32'hc4057d2;
      42858: inst = 32'h8220000;
      42859: inst = 32'hc20e407;
      42860: inst = 32'h10408000;
      42861: inst = 32'hc4053b3;
      42862: inst = 32'h8220000;
      42863: inst = 32'hc207d9a;
      42864: inst = 32'h10408000;
      42865: inst = 32'hc4053b6;
      42866: inst = 32'h8220000;
      42867: inst = 32'hc2065fe;
      42868: inst = 32'h10408000;
      42869: inst = 32'hc4053b7;
      42870: inst = 32'h8220000;
      42871: inst = 32'hc2065fd;
      42872: inst = 32'h10408000;
      42873: inst = 32'hc4053b8;
      42874: inst = 32'h8220000;
      42875: inst = 32'h10408000;
      42876: inst = 32'hc4053b9;
      42877: inst = 32'h8220000;
      42878: inst = 32'hc20661e;
      42879: inst = 32'h10408000;
      42880: inst = 32'hc4053ba;
      42881: inst = 32'h8220000;
      42882: inst = 32'hc20bb86;
      42883: inst = 32'h10408000;
      42884: inst = 32'hc4053bb;
      42885: inst = 32'h8220000;
      42886: inst = 32'h10408000;
      42887: inst = 32'hc4054db;
      42888: inst = 32'h8220000;
      42889: inst = 32'hc20e6fa;
      42890: inst = 32'h10408000;
      42891: inst = 32'hc4053c9;
      42892: inst = 32'h8220000;
      42893: inst = 32'h10408000;
      42894: inst = 32'hc4053cd;
      42895: inst = 32'h8220000;
      42896: inst = 32'h10408000;
      42897: inst = 32'hc4055a7;
      42898: inst = 32'h8220000;
      42899: inst = 32'hc20e6fb;
      42900: inst = 32'h10408000;
      42901: inst = 32'hc4053ca;
      42902: inst = 32'h8220000;
      42903: inst = 32'h10408000;
      42904: inst = 32'hc4053cc;
      42905: inst = 32'h8220000;
      42906: inst = 32'h10408000;
      42907: inst = 32'hc405487;
      42908: inst = 32'h8220000;
      42909: inst = 32'h10408000;
      42910: inst = 32'hc40548f;
      42911: inst = 32'h8220000;
      42912: inst = 32'h10408000;
      42913: inst = 32'hc405547;
      42914: inst = 32'h8220000;
      42915: inst = 32'h10408000;
      42916: inst = 32'hc40554f;
      42917: inst = 32'h8220000;
      42918: inst = 32'hc20defb;
      42919: inst = 32'h10408000;
      42920: inst = 32'hc4053cb;
      42921: inst = 32'h8220000;
      42922: inst = 32'h10408000;
      42923: inst = 32'hc405428;
      42924: inst = 32'h8220000;
      42925: inst = 32'h10408000;
      42926: inst = 32'hc405429;
      42927: inst = 32'h8220000;
      42928: inst = 32'h10408000;
      42929: inst = 32'hc40542a;
      42930: inst = 32'h8220000;
      42931: inst = 32'h10408000;
      42932: inst = 32'hc40542b;
      42933: inst = 32'h8220000;
      42934: inst = 32'h10408000;
      42935: inst = 32'hc40542c;
      42936: inst = 32'h8220000;
      42937: inst = 32'h10408000;
      42938: inst = 32'hc40542d;
      42939: inst = 32'h8220000;
      42940: inst = 32'h10408000;
      42941: inst = 32'hc40542e;
      42942: inst = 32'h8220000;
      42943: inst = 32'h10408000;
      42944: inst = 32'hc405488;
      42945: inst = 32'h8220000;
      42946: inst = 32'h10408000;
      42947: inst = 32'hc405489;
      42948: inst = 32'h8220000;
      42949: inst = 32'h10408000;
      42950: inst = 32'hc40548a;
      42951: inst = 32'h8220000;
      42952: inst = 32'h10408000;
      42953: inst = 32'hc40548b;
      42954: inst = 32'h8220000;
      42955: inst = 32'h10408000;
      42956: inst = 32'hc40548c;
      42957: inst = 32'h8220000;
      42958: inst = 32'h10408000;
      42959: inst = 32'hc40548d;
      42960: inst = 32'h8220000;
      42961: inst = 32'h10408000;
      42962: inst = 32'hc40548e;
      42963: inst = 32'h8220000;
      42964: inst = 32'h10408000;
      42965: inst = 32'hc4054e7;
      42966: inst = 32'h8220000;
      42967: inst = 32'h10408000;
      42968: inst = 32'hc4054ea;
      42969: inst = 32'h8220000;
      42970: inst = 32'h10408000;
      42971: inst = 32'hc4054ed;
      42972: inst = 32'h8220000;
      42973: inst = 32'h10408000;
      42974: inst = 32'hc4054ee;
      42975: inst = 32'h8220000;
      42976: inst = 32'h10408000;
      42977: inst = 32'hc4054ef;
      42978: inst = 32'h8220000;
      42979: inst = 32'h10408000;
      42980: inst = 32'hc40554a;
      42981: inst = 32'h8220000;
      42982: inst = 32'h10408000;
      42983: inst = 32'hc40554d;
      42984: inst = 32'h8220000;
      42985: inst = 32'h10408000;
      42986: inst = 32'hc40554e;
      42987: inst = 32'h8220000;
      42988: inst = 32'h10408000;
      42989: inst = 32'hc4055a8;
      42990: inst = 32'h8220000;
      42991: inst = 32'h10408000;
      42992: inst = 32'hc4055a9;
      42993: inst = 32'h8220000;
      42994: inst = 32'h10408000;
      42995: inst = 32'hc4055aa;
      42996: inst = 32'h8220000;
      42997: inst = 32'h10408000;
      42998: inst = 32'hc4055ab;
      42999: inst = 32'h8220000;
      43000: inst = 32'h10408000;
      43001: inst = 32'hc4055ac;
      43002: inst = 32'h8220000;
      43003: inst = 32'h10408000;
      43004: inst = 32'hc4055ad;
      43005: inst = 32'h8220000;
      43006: inst = 32'h10408000;
      43007: inst = 32'hc4055ae;
      43008: inst = 32'h8220000;
      43009: inst = 32'h10408000;
      43010: inst = 32'hc405609;
      43011: inst = 32'h8220000;
      43012: inst = 32'h10408000;
      43013: inst = 32'hc40560b;
      43014: inst = 32'h8220000;
      43015: inst = 32'h10408000;
      43016: inst = 32'hc405669;
      43017: inst = 32'h8220000;
      43018: inst = 32'hc20cbc7;
      43019: inst = 32'h10408000;
      43020: inst = 32'hc405412;
      43021: inst = 32'h8220000;
      43022: inst = 32'h10408000;
      43023: inst = 32'hc405472;
      43024: inst = 32'h8220000;
      43025: inst = 32'hc20edb1;
      43026: inst = 32'h10408000;
      43027: inst = 32'hc405413;
      43028: inst = 32'h8220000;
      43029: inst = 32'hc20db43;
      43030: inst = 32'h10408000;
      43031: inst = 32'hc405414;
      43032: inst = 32'h8220000;
      43033: inst = 32'hc207d78;
      43034: inst = 32'h10408000;
      43035: inst = 32'hc405416;
      43036: inst = 32'h8220000;
      43037: inst = 32'hc206dbc;
      43038: inst = 32'h10408000;
      43039: inst = 32'hc405417;
      43040: inst = 32'h8220000;
      43041: inst = 32'h10408000;
      43042: inst = 32'hc405477;
      43043: inst = 32'h8220000;
      43044: inst = 32'hc206dbb;
      43045: inst = 32'h10408000;
      43046: inst = 32'hc405418;
      43047: inst = 32'h8220000;
      43048: inst = 32'h10408000;
      43049: inst = 32'hc405419;
      43050: inst = 32'h8220000;
      43051: inst = 32'h10408000;
      43052: inst = 32'hc405478;
      43053: inst = 32'h8220000;
      43054: inst = 32'h10408000;
      43055: inst = 32'hc405479;
      43056: inst = 32'h8220000;
      43057: inst = 32'hc206ddc;
      43058: inst = 32'h10408000;
      43059: inst = 32'hc40541a;
      43060: inst = 32'h8220000;
      43061: inst = 32'h10408000;
      43062: inst = 32'hc40547a;
      43063: inst = 32'h8220000;
      43064: inst = 32'hc20bb66;
      43065: inst = 32'h10408000;
      43066: inst = 32'hc40541b;
      43067: inst = 32'h8220000;
      43068: inst = 32'h10408000;
      43069: inst = 32'hc40547b;
      43070: inst = 32'h8220000;
      43071: inst = 32'h10408000;
      43072: inst = 32'hc40559b;
      43073: inst = 32'h8220000;
      43074: inst = 32'hc20eed8;
      43075: inst = 32'h10408000;
      43076: inst = 32'hc405427;
      43077: inst = 32'h8220000;
      43078: inst = 32'h10408000;
      43079: inst = 32'hc40542f;
      43080: inst = 32'h8220000;
      43081: inst = 32'hc20edd2;
      43082: inst = 32'h10408000;
      43083: inst = 32'hc405473;
      43084: inst = 32'h8220000;
      43085: inst = 32'hc20db42;
      43086: inst = 32'h10408000;
      43087: inst = 32'hc405474;
      43088: inst = 32'h8220000;
      43089: inst = 32'hc207d79;
      43090: inst = 32'h10408000;
      43091: inst = 32'hc405476;
      43092: inst = 32'h8220000;
      43093: inst = 32'hc20e590;
      43094: inst = 32'h10408000;
      43095: inst = 32'hc4054d3;
      43096: inst = 32'h8220000;
      43097: inst = 32'hc20e363;
      43098: inst = 32'h10408000;
      43099: inst = 32'hc4054d4;
      43100: inst = 32'h8220000;
      43101: inst = 32'hc20d3a6;
      43102: inst = 32'h10408000;
      43103: inst = 32'hc4054d5;
      43104: inst = 32'h8220000;
      43105: inst = 32'hc207dba;
      43106: inst = 32'h10408000;
      43107: inst = 32'hc4054d6;
      43108: inst = 32'h8220000;
      43109: inst = 32'hc2075fd;
      43110: inst = 32'h10408000;
      43111: inst = 32'hc4054d7;
      43112: inst = 32'h8220000;
      43113: inst = 32'h10408000;
      43114: inst = 32'hc4054d8;
      43115: inst = 32'h8220000;
      43116: inst = 32'h10408000;
      43117: inst = 32'hc4054d9;
      43118: inst = 32'h8220000;
      43119: inst = 32'hc206e1e;
      43120: inst = 32'h10408000;
      43121: inst = 32'hc4054da;
      43122: inst = 32'h8220000;
      43123: inst = 32'hc204a69;
      43124: inst = 32'h10408000;
      43125: inst = 32'hc4054e8;
      43126: inst = 32'h8220000;
      43127: inst = 32'h10408000;
      43128: inst = 32'hc4054e9;
      43129: inst = 32'h8220000;
      43130: inst = 32'h10408000;
      43131: inst = 32'hc4054eb;
      43132: inst = 32'h8220000;
      43133: inst = 32'h10408000;
      43134: inst = 32'hc4054ec;
      43135: inst = 32'h8220000;
      43136: inst = 32'h10408000;
      43137: inst = 32'hc405548;
      43138: inst = 32'h8220000;
      43139: inst = 32'h10408000;
      43140: inst = 32'hc405549;
      43141: inst = 32'h8220000;
      43142: inst = 32'h10408000;
      43143: inst = 32'hc40554b;
      43144: inst = 32'h8220000;
      43145: inst = 32'h10408000;
      43146: inst = 32'hc40554c;
      43147: inst = 32'h8220000;
      43148: inst = 32'h10408000;
      43149: inst = 32'hc405608;
      43150: inst = 32'h8220000;
      43151: inst = 32'h10408000;
      43152: inst = 32'hc40560a;
      43153: inst = 32'h8220000;
      43154: inst = 32'h10408000;
      43155: inst = 32'hc40560c;
      43156: inst = 32'h8220000;
      43157: inst = 32'h10408000;
      43158: inst = 32'hc405668;
      43159: inst = 32'h8220000;
      43160: inst = 32'h10408000;
      43161: inst = 32'hc40566a;
      43162: inst = 32'h8220000;
      43163: inst = 32'hc20eba3;
      43164: inst = 32'h10408000;
      43165: inst = 32'hc405535;
      43166: inst = 32'h8220000;
      43167: inst = 32'hc207411;
      43168: inst = 32'h10408000;
      43169: inst = 32'hc405536;
      43170: inst = 32'h8220000;
      43171: inst = 32'hc205bf2;
      43172: inst = 32'h10408000;
      43173: inst = 32'hc405537;
      43174: inst = 32'h8220000;
      43175: inst = 32'h10408000;
      43176: inst = 32'hc40553a;
      43177: inst = 32'h8220000;
      43178: inst = 32'hc205c12;
      43179: inst = 32'h10408000;
      43180: inst = 32'hc405538;
      43181: inst = 32'h8220000;
      43182: inst = 32'h10408000;
      43183: inst = 32'hc405539;
      43184: inst = 32'h8220000;
      43185: inst = 32'h10408000;
      43186: inst = 32'hc4055f9;
      43187: inst = 32'h8220000;
      43188: inst = 32'hc20bb25;
      43189: inst = 32'h10408000;
      43190: inst = 32'hc40553b;
      43191: inst = 32'h8220000;
      43192: inst = 32'h10408000;
      43193: inst = 32'hc4056bb;
      43194: inst = 32'h8220000;
      43195: inst = 32'h10408000;
      43196: inst = 32'hc40571b;
      43197: inst = 32'h8220000;
      43198: inst = 32'h10408000;
      43199: inst = 32'hc40577b;
      43200: inst = 32'h8220000;
      43201: inst = 32'hc20dba4;
      43202: inst = 32'h10408000;
      43203: inst = 32'hc405593;
      43204: inst = 32'h8220000;
      43205: inst = 32'h10408000;
      43206: inst = 32'hc4056b4;
      43207: inst = 32'h8220000;
      43208: inst = 32'hc206288;
      43209: inst = 32'h10408000;
      43210: inst = 32'hc405596;
      43211: inst = 32'h8220000;
      43212: inst = 32'hc205bb1;
      43213: inst = 32'h10408000;
      43214: inst = 32'hc405597;
      43215: inst = 32'h8220000;
      43216: inst = 32'hc2052ec;
      43217: inst = 32'h10408000;
      43218: inst = 32'hc405598;
      43219: inst = 32'h8220000;
      43220: inst = 32'hc20532d;
      43221: inst = 32'h10408000;
      43222: inst = 32'hc405599;
      43223: inst = 32'h8220000;
      43224: inst = 32'hc205390;
      43225: inst = 32'h10408000;
      43226: inst = 32'hc40559a;
      43227: inst = 32'h8220000;
      43228: inst = 32'hc20e6d9;
      43229: inst = 32'h10408000;
      43230: inst = 32'hc4055af;
      43231: inst = 32'h8220000;
      43232: inst = 32'hc2062ea;
      43233: inst = 32'h10408000;
      43234: inst = 32'hc4055f6;
      43235: inst = 32'h8220000;
      43236: inst = 32'hc2064f8;
      43237: inst = 32'h10408000;
      43238: inst = 32'hc4055f7;
      43239: inst = 32'h8220000;
      43240: inst = 32'hc205bd1;
      43241: inst = 32'h10408000;
      43242: inst = 32'hc4055f8;
      43243: inst = 32'h8220000;
      43244: inst = 32'hc2064d6;
      43245: inst = 32'h10408000;
      43246: inst = 32'hc4055fa;
      43247: inst = 32'h8220000;
      43248: inst = 32'hc20bba7;
      43249: inst = 32'h10408000;
      43250: inst = 32'hc4055fb;
      43251: inst = 32'h8220000;
      43252: inst = 32'hc20eeb7;
      43253: inst = 32'h10408000;
      43254: inst = 32'hc405607;
      43255: inst = 32'h8220000;
      43256: inst = 32'hc20d699;
      43257: inst = 32'h10408000;
      43258: inst = 32'hc40560d;
      43259: inst = 32'h8220000;
      43260: inst = 32'hc20b553;
      43261: inst = 32'h10408000;
      43262: inst = 32'hc40560e;
      43263: inst = 32'h8220000;
      43264: inst = 32'hc2083cd;
      43265: inst = 32'h10408000;
      43266: inst = 32'hc40560f;
      43267: inst = 32'h8220000;
      43268: inst = 32'hc20736c;
      43269: inst = 32'h10408000;
      43270: inst = 32'hc405610;
      43271: inst = 32'h8220000;
      43272: inst = 32'hc20a4d0;
      43273: inst = 32'h10408000;
      43274: inst = 32'hc405611;
      43275: inst = 32'h8220000;
      43276: inst = 32'hc20de55;
      43277: inst = 32'h10408000;
      43278: inst = 32'hc405612;
      43279: inst = 32'h8220000;
      43280: inst = 32'hc2062eb;
      43281: inst = 32'h10408000;
      43282: inst = 32'hc405656;
      43283: inst = 32'h8220000;
      43284: inst = 32'hc206496;
      43285: inst = 32'h10408000;
      43286: inst = 32'hc405657;
      43287: inst = 32'h8220000;
      43288: inst = 32'hc205bb0;
      43289: inst = 32'h10408000;
      43290: inst = 32'hc405658;
      43291: inst = 32'h8220000;
      43292: inst = 32'hc2063f2;
      43293: inst = 32'h10408000;
      43294: inst = 32'hc405659;
      43295: inst = 32'h8220000;
      43296: inst = 32'hc206475;
      43297: inst = 32'h10408000;
      43298: inst = 32'hc40565a;
      43299: inst = 32'h8220000;
      43300: inst = 32'hc20bb87;
      43301: inst = 32'h10408000;
      43302: inst = 32'hc40565b;
      43303: inst = 32'h8220000;
      43304: inst = 32'hc209492;
      43305: inst = 32'h10408000;
      43306: inst = 32'hc40566b;
      43307: inst = 32'h8220000;
      43308: inst = 32'hc204228;
      43309: inst = 32'h10408000;
      43310: inst = 32'hc40566c;
      43311: inst = 32'h8220000;
      43312: inst = 32'h10408000;
      43313: inst = 32'hc405760;
      43314: inst = 32'h8220000;
      43315: inst = 32'hc20632c;
      43316: inst = 32'h10408000;
      43317: inst = 32'hc40566d;
      43318: inst = 32'h8220000;
      43319: inst = 32'hc20a4d1;
      43320: inst = 32'h10408000;
      43321: inst = 32'hc40566e;
      43322: inst = 32'h8220000;
      43323: inst = 32'hc20cdf4;
      43324: inst = 32'h10408000;
      43325: inst = 32'hc40566f;
      43326: inst = 32'h8220000;
      43327: inst = 32'hc20c593;
      43328: inst = 32'h10408000;
      43329: inst = 32'hc405670;
      43330: inst = 32'h8220000;
      43331: inst = 32'hc20944f;
      43332: inst = 32'h10408000;
      43333: inst = 32'hc405671;
      43334: inst = 32'h8220000;
      43335: inst = 32'hc20734c;
      43336: inst = 32'h10408000;
      43337: inst = 32'hc405672;
      43338: inst = 32'h8220000;
      43339: inst = 32'hc20a4b0;
      43340: inst = 32'h10408000;
      43341: inst = 32'hc405673;
      43342: inst = 32'h8220000;
      43343: inst = 32'hc20e3e6;
      43344: inst = 32'h10408000;
      43345: inst = 32'hc4056b3;
      43346: inst = 32'h8220000;
      43347: inst = 32'hc209ac5;
      43348: inst = 32'h10408000;
      43349: inst = 32'hc4056b5;
      43350: inst = 32'h8220000;
      43351: inst = 32'hc206350;
      43352: inst = 32'h10408000;
      43353: inst = 32'hc4056ba;
      43354: inst = 32'h8220000;
      43355: inst = 32'h10408000;
      43356: inst = 32'hc40571a;
      43357: inst = 32'h8220000;
      43358: inst = 32'h10408000;
      43359: inst = 32'hc405776;
      43360: inst = 32'h8220000;
      43361: inst = 32'hc2052ac;
      43362: inst = 32'h10408000;
      43363: inst = 32'hc4056ca;
      43364: inst = 32'h8220000;
      43365: inst = 32'h10408000;
      43366: inst = 32'hc4056d0;
      43367: inst = 32'h8220000;
      43368: inst = 32'h10408000;
      43369: inst = 32'hc4057bf;
      43370: inst = 32'h8220000;
      43371: inst = 32'hc204a6a;
      43372: inst = 32'h10408000;
      43373: inst = 32'hc4056cb;
      43374: inst = 32'h8220000;
      43375: inst = 32'h10408000;
      43376: inst = 32'hc4056cc;
      43377: inst = 32'h8220000;
      43378: inst = 32'h10408000;
      43379: inst = 32'hc4056cd;
      43380: inst = 32'h8220000;
      43381: inst = 32'h10408000;
      43382: inst = 32'hc4056ce;
      43383: inst = 32'h8220000;
      43384: inst = 32'h10408000;
      43385: inst = 32'hc4057c0;
      43386: inst = 32'h8220000;
      43387: inst = 32'hc20528b;
      43388: inst = 32'h10408000;
      43389: inst = 32'hc4056cf;
      43390: inst = 32'h8220000;
      43391: inst = 32'hc205acd;
      43392: inst = 32'h10408000;
      43393: inst = 32'hc4056d1;
      43394: inst = 32'h8220000;
      43395: inst = 32'hc205aed;
      43396: inst = 32'h10408000;
      43397: inst = 32'hc4056d2;
      43398: inst = 32'h8220000;
      43399: inst = 32'h10408000;
      43400: inst = 32'hc40575f;
      43401: inst = 32'h8220000;
      43402: inst = 32'hc20632f;
      43403: inst = 32'h10408000;
      43404: inst = 32'hc4056d3;
      43405: inst = 32'h8220000;
      43406: inst = 32'h10408000;
      43407: inst = 32'hc405715;
      43408: inst = 32'h8220000;
      43409: inst = 32'hc20634f;
      43410: inst = 32'h10408000;
      43411: inst = 32'hc4056fe;
      43412: inst = 32'h8220000;
      43413: inst = 32'hc204208;
      43414: inst = 32'h10408000;
      43415: inst = 32'hc4056ff;
      43416: inst = 32'h8220000;
      43417: inst = 32'h10408000;
      43418: inst = 32'hc405700;
      43419: inst = 32'h8220000;
      43420: inst = 32'hc209ae6;
      43421: inst = 32'h10408000;
      43422: inst = 32'hc405714;
      43423: inst = 32'h8220000;
      43424: inst = 32'hc206370;
      43425: inst = 32'h10408000;
      43426: inst = 32'hc405716;
      43427: inst = 32'h8220000;
      43428: inst = 32'h10408000;
      43429: inst = 32'hc405777;
      43430: inst = 32'h8220000;
      43431: inst = 32'h10408000;
      43432: inst = 32'hc405778;
      43433: inst = 32'h8220000;
      43434: inst = 32'h10408000;
      43435: inst = 32'hc405779;
      43436: inst = 32'h8220000;
      43437: inst = 32'hc20c303;
      43438: inst = 32'h10408000;
      43439: inst = 32'hc405772;
      43440: inst = 32'h8220000;
      43441: inst = 32'hc20aaa2;
      43442: inst = 32'h10408000;
      43443: inst = 32'hc405773;
      43444: inst = 32'h8220000;
      43445: inst = 32'hc2072ea;
      43446: inst = 32'h10408000;
      43447: inst = 32'hc405774;
      43448: inst = 32'h8220000;
      43449: inst = 32'hc205b72;
      43450: inst = 32'h10408000;
      43451: inst = 32'hc405775;
      43452: inst = 32'h8220000;
      43453: inst = 32'hc206371;
      43454: inst = 32'h10408000;
      43455: inst = 32'hc40577a;
      43456: inst = 32'h8220000;
      43457: inst = 32'hc20bae3;
      43458: inst = 32'h10408000;
      43459: inst = 32'hc4057d3;
      43460: inst = 32'h8220000;
      43461: inst = 32'hc20bb04;
      43462: inst = 32'h10408000;
      43463: inst = 32'hc4057d4;
      43464: inst = 32'h8220000;
      43465: inst = 32'hc20b325;
      43466: inst = 32'h10408000;
      43467: inst = 32'hc4057d5;
      43468: inst = 32'h8220000;
      43469: inst = 32'h10408000;
      43470: inst = 32'hc4057d6;
      43471: inst = 32'h8220000;
      43472: inst = 32'h10408000;
      43473: inst = 32'hc4057d7;
      43474: inst = 32'h8220000;
      43475: inst = 32'h10408000;
      43476: inst = 32'hc4057d8;
      43477: inst = 32'h8220000;
      43478: inst = 32'h10408000;
      43479: inst = 32'hc4057d9;
      43480: inst = 32'h8220000;
      43481: inst = 32'h10408000;
      43482: inst = 32'hc4057da;
      43483: inst = 32'h8220000;
      43484: inst = 32'hc20c344;
      43485: inst = 32'h10408000;
      43486: inst = 32'hc4057db;
      43487: inst = 32'h8220000;
      43488: inst = 32'h58000000;
      43489: inst = 32'h11800000;
      43490: inst = 32'hd800000;
      43491: inst = 32'h11a00000;
      43492: inst = 32'hda00000;
      43493: inst = 32'h25ad5800;
      43494: inst = 32'h15ca6800;
      43495: inst = 32'h21c00001;
      43496: inst = 32'h59200000;
      43497: inst = 32'h298c0001;
      43498: inst = 32'h13e00000;
      43499: inst = 32'hfe0a9e5;
      43500: inst = 32'h5be00000;
      43501: inst = 32'h11800000;
      43502: inst = 32'hd800000;
      43503: inst = 32'h258c5800;
      43504: inst = 32'h15aa6000;
      43505: inst = 32'h13e00000;
      43506: inst = 32'hfe0a9f8;
      43507: inst = 32'h21a00001;
      43508: inst = 32'h5be00000;
      43509: inst = 32'h13e00000;
      43510: inst = 32'hfe0a9ef;
      43511: inst = 32'h5be00000;
      43512: inst = 32'h2d8c5800;
      43513: inst = 32'h2d8a6000;
      43514: inst = 32'h59200000;
      43515: inst = 32'h11800000;
      43516: inst = 32'hd800000;
      43517: inst = 32'h29ab0000;
      43518: inst = 32'h31ad0001;
      43519: inst = 32'h258c5000;
      43520: inst = 32'h21a00000;
      43521: inst = 32'h59200000;
      43522: inst = 32'h13e00000;
      43523: inst = 32'hfe0a9fe;
      43524: inst = 32'h5be00000;
      43525: inst = 32'h10608000;
      43526: inst = 32'hc600000;
      43527: inst = 32'hc20aaaa;
      43528: inst = 32'h4c210000;
      43529: inst = 32'h8230000;
      43530: inst = 32'h104000fe;
      43531: inst = 32'hc40502a;
      43532: inst = 32'h30420001;
      43533: inst = 32'h13e00000;
      43534: inst = 32'hfe0aa0c;
      43535: inst = 32'h1c400000;
      43536: inst = 32'h5be00000;
      43537: inst = 32'h13e00000;
      43538: inst = 32'hfe0aa08;
      43539: inst = 32'h5be00000;
    endcase
  end
endmodule
