`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: lirc572
// Engineer: lirc572
// 
// Create Date: 
// Design Name: NECPU
// Module Name: InstMem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module instMem (
    input  [31:0]  address,
    output reg [31:0] inst
  );
  always @ (address) begin
    inst = 32'd0;
    case (address)
      0: inst = 32'h10000000;
      1: inst = 32'hc000005;
      2: inst = 32'h13e00000;
      3: inst = 32'hfe00055;
      4: inst = 32'h5be00000;
      5: inst = 32'h13c0007f;
      6: inst = 32'hfc02815;
      7: inst = 32'h33de0001;
      8: inst = 32'h13e00000;
      9: inst = 32'hfe00007;
      10: inst = 32'h1fc00000;
      11: inst = 32'h5be00000;
      12: inst = 32'h10000000;
      13: inst = 32'hc000011;
      14: inst = 32'h13e00000;
      15: inst = 32'hfe048ad;
      16: inst = 32'h5be00000;
      17: inst = 32'h13c0007f;
      18: inst = 32'hfc02815;
      19: inst = 32'h33de0001;
      20: inst = 32'h13e00000;
      21: inst = 32'hfe00013;
      22: inst = 32'h1fc00000;
      23: inst = 32'h5be00000;
      24: inst = 32'h10000000;
      25: inst = 32'hc000000;
      26: inst = 32'h10200000;
      27: inst = 32'hc20001f;
      28: inst = 32'h13e00000;
      29: inst = 32'hfe08960;
      30: inst = 32'h5be00000;
      31: inst = 32'h10000000;
      32: inst = 32'hc000024;
      33: inst = 32'h13e00000;
      34: inst = 32'hfe050fe;
      35: inst = 32'h5be00000;
      36: inst = 32'h13c001fc;
      37: inst = 32'hfc0a055;
      38: inst = 32'h33de0001;
      39: inst = 32'h13e00000;
      40: inst = 32'hfe00026;
      41: inst = 32'h1fc00000;
      42: inst = 32'h5be00000;
      43: inst = 32'h10000000;
      44: inst = 32'hc00002b;
      45: inst = 32'h10200000;
      46: inst = 32'hc200032;
      47: inst = 32'h13e00000;
      48: inst = 32'hfe08960;
      49: inst = 32'h5be00000;
      50: inst = 32'h10200000;
      51: inst = 32'hc20000c;
      52: inst = 32'h10400000;
      53: inst = 32'hc400009;
      54: inst = 32'h10000000;
      55: inst = 32'hc00003b;
      56: inst = 32'h13e00000;
      57: inst = 32'hfe0896a;
      58: inst = 32'h5be00000;
      59: inst = 32'h10200000;
      60: inst = 32'hc200000;
      61: inst = 32'h10000000;
      62: inst = 32'hc000042;
      63: inst = 32'h13e00000;
      64: inst = 32'hfe085ad;
      65: inst = 32'h5be00000;
      66: inst = 32'h13e00000;
      67: inst = 32'hfe00045;
      68: inst = 32'h5be00000;
      69: inst = 32'h10608000;
      70: inst = 32'hc600000;
      71: inst = 32'h10200000;
      72: inst = 32'hc20aaaa;
      73: inst = 32'h4c210000;
      74: inst = 32'h8230000;
      75: inst = 32'h104000fe;
      76: inst = 32'hc40502a;
      77: inst = 32'h30420001;
      78: inst = 32'h13e00000;
      79: inst = 32'hfe0004d;
      80: inst = 32'h1c400000;
      81: inst = 32'h5be00000;
      82: inst = 32'h13e00000;
      83: inst = 32'hfe00049;
      84: inst = 32'h5be00000;
      85: inst = 32'hc20eeb6;
      86: inst = 32'h10408000;
      87: inst = 32'hc403fe0;
      88: inst = 32'h8220000;
      89: inst = 32'h10408000;
      90: inst = 32'hc403fe1;
      91: inst = 32'h8220000;
      92: inst = 32'h10408000;
      93: inst = 32'hc403fe2;
      94: inst = 32'h8220000;
      95: inst = 32'h10408000;
      96: inst = 32'hc403fe3;
      97: inst = 32'h8220000;
      98: inst = 32'h10408000;
      99: inst = 32'hc403fe4;
      100: inst = 32'h8220000;
      101: inst = 32'h10408000;
      102: inst = 32'hc403fe5;
      103: inst = 32'h8220000;
      104: inst = 32'h10408000;
      105: inst = 32'hc403fe6;
      106: inst = 32'h8220000;
      107: inst = 32'h10408000;
      108: inst = 32'hc403fe7;
      109: inst = 32'h8220000;
      110: inst = 32'h10408000;
      111: inst = 32'hc403fe8;
      112: inst = 32'h8220000;
      113: inst = 32'h10408000;
      114: inst = 32'hc403fe9;
      115: inst = 32'h8220000;
      116: inst = 32'h10408000;
      117: inst = 32'hc403fea;
      118: inst = 32'h8220000;
      119: inst = 32'h10408000;
      120: inst = 32'hc403fec;
      121: inst = 32'h8220000;
      122: inst = 32'h10408000;
      123: inst = 32'hc403fed;
      124: inst = 32'h8220000;
      125: inst = 32'h10408000;
      126: inst = 32'hc403fee;
      127: inst = 32'h8220000;
      128: inst = 32'h10408000;
      129: inst = 32'hc403fef;
      130: inst = 32'h8220000;
      131: inst = 32'h10408000;
      132: inst = 32'hc403ff0;
      133: inst = 32'h8220000;
      134: inst = 32'h10408000;
      135: inst = 32'hc403ff1;
      136: inst = 32'h8220000;
      137: inst = 32'h10408000;
      138: inst = 32'hc403ff2;
      139: inst = 32'h8220000;
      140: inst = 32'h10408000;
      141: inst = 32'hc403ff3;
      142: inst = 32'h8220000;
      143: inst = 32'h10408000;
      144: inst = 32'hc403ff4;
      145: inst = 32'h8220000;
      146: inst = 32'h10408000;
      147: inst = 32'hc403ff5;
      148: inst = 32'h8220000;
      149: inst = 32'h10408000;
      150: inst = 32'hc403ff6;
      151: inst = 32'h8220000;
      152: inst = 32'h10408000;
      153: inst = 32'hc403ff7;
      154: inst = 32'h8220000;
      155: inst = 32'h10408000;
      156: inst = 32'hc403ff8;
      157: inst = 32'h8220000;
      158: inst = 32'h10408000;
      159: inst = 32'hc403ff9;
      160: inst = 32'h8220000;
      161: inst = 32'h10408000;
      162: inst = 32'hc403ffa;
      163: inst = 32'h8220000;
      164: inst = 32'h10408000;
      165: inst = 32'hc403ffb;
      166: inst = 32'h8220000;
      167: inst = 32'h10408000;
      168: inst = 32'hc403ffc;
      169: inst = 32'h8220000;
      170: inst = 32'h10408000;
      171: inst = 32'hc403ffd;
      172: inst = 32'h8220000;
      173: inst = 32'h10408000;
      174: inst = 32'hc403ffe;
      175: inst = 32'h8220000;
      176: inst = 32'h10408000;
      177: inst = 32'hc403fff;
      178: inst = 32'h8220000;
      179: inst = 32'h10408000;
      180: inst = 32'hc404000;
      181: inst = 32'h8220000;
      182: inst = 32'h10408000;
      183: inst = 32'hc404001;
      184: inst = 32'h8220000;
      185: inst = 32'h10408000;
      186: inst = 32'hc404002;
      187: inst = 32'h8220000;
      188: inst = 32'h10408000;
      189: inst = 32'hc404003;
      190: inst = 32'h8220000;
      191: inst = 32'h10408000;
      192: inst = 32'hc404004;
      193: inst = 32'h8220000;
      194: inst = 32'h10408000;
      195: inst = 32'hc404005;
      196: inst = 32'h8220000;
      197: inst = 32'h10408000;
      198: inst = 32'hc404006;
      199: inst = 32'h8220000;
      200: inst = 32'h10408000;
      201: inst = 32'hc404007;
      202: inst = 32'h8220000;
      203: inst = 32'h10408000;
      204: inst = 32'hc404008;
      205: inst = 32'h8220000;
      206: inst = 32'h10408000;
      207: inst = 32'hc404009;
      208: inst = 32'h8220000;
      209: inst = 32'h10408000;
      210: inst = 32'hc40400a;
      211: inst = 32'h8220000;
      212: inst = 32'h10408000;
      213: inst = 32'hc40400b;
      214: inst = 32'h8220000;
      215: inst = 32'h10408000;
      216: inst = 32'hc40400c;
      217: inst = 32'h8220000;
      218: inst = 32'h10408000;
      219: inst = 32'hc40400d;
      220: inst = 32'h8220000;
      221: inst = 32'h10408000;
      222: inst = 32'hc40400e;
      223: inst = 32'h8220000;
      224: inst = 32'h10408000;
      225: inst = 32'hc40400f;
      226: inst = 32'h8220000;
      227: inst = 32'h10408000;
      228: inst = 32'hc404010;
      229: inst = 32'h8220000;
      230: inst = 32'h10408000;
      231: inst = 32'hc404011;
      232: inst = 32'h8220000;
      233: inst = 32'h10408000;
      234: inst = 32'hc404012;
      235: inst = 32'h8220000;
      236: inst = 32'h10408000;
      237: inst = 32'hc404013;
      238: inst = 32'h8220000;
      239: inst = 32'h10408000;
      240: inst = 32'hc404014;
      241: inst = 32'h8220000;
      242: inst = 32'h10408000;
      243: inst = 32'hc404015;
      244: inst = 32'h8220000;
      245: inst = 32'h10408000;
      246: inst = 32'hc404016;
      247: inst = 32'h8220000;
      248: inst = 32'h10408000;
      249: inst = 32'hc404017;
      250: inst = 32'h8220000;
      251: inst = 32'h10408000;
      252: inst = 32'hc404018;
      253: inst = 32'h8220000;
      254: inst = 32'h10408000;
      255: inst = 32'hc404019;
      256: inst = 32'h8220000;
      257: inst = 32'h10408000;
      258: inst = 32'hc40401a;
      259: inst = 32'h8220000;
      260: inst = 32'h10408000;
      261: inst = 32'hc40401b;
      262: inst = 32'h8220000;
      263: inst = 32'h10408000;
      264: inst = 32'hc40401c;
      265: inst = 32'h8220000;
      266: inst = 32'h10408000;
      267: inst = 32'hc40401d;
      268: inst = 32'h8220000;
      269: inst = 32'h10408000;
      270: inst = 32'hc40401e;
      271: inst = 32'h8220000;
      272: inst = 32'h10408000;
      273: inst = 32'hc40401f;
      274: inst = 32'h8220000;
      275: inst = 32'h10408000;
      276: inst = 32'hc404020;
      277: inst = 32'h8220000;
      278: inst = 32'h10408000;
      279: inst = 32'hc404021;
      280: inst = 32'h8220000;
      281: inst = 32'h10408000;
      282: inst = 32'hc404022;
      283: inst = 32'h8220000;
      284: inst = 32'h10408000;
      285: inst = 32'hc404023;
      286: inst = 32'h8220000;
      287: inst = 32'h10408000;
      288: inst = 32'hc404024;
      289: inst = 32'h8220000;
      290: inst = 32'h10408000;
      291: inst = 32'hc404025;
      292: inst = 32'h8220000;
      293: inst = 32'h10408000;
      294: inst = 32'hc404026;
      295: inst = 32'h8220000;
      296: inst = 32'h10408000;
      297: inst = 32'hc404027;
      298: inst = 32'h8220000;
      299: inst = 32'h10408000;
      300: inst = 32'hc404028;
      301: inst = 32'h8220000;
      302: inst = 32'h10408000;
      303: inst = 32'hc404029;
      304: inst = 32'h8220000;
      305: inst = 32'h10408000;
      306: inst = 32'hc40402a;
      307: inst = 32'h8220000;
      308: inst = 32'h10408000;
      309: inst = 32'hc40402b;
      310: inst = 32'h8220000;
      311: inst = 32'h10408000;
      312: inst = 32'hc40402c;
      313: inst = 32'h8220000;
      314: inst = 32'h10408000;
      315: inst = 32'hc40402d;
      316: inst = 32'h8220000;
      317: inst = 32'h10408000;
      318: inst = 32'hc40402e;
      319: inst = 32'h8220000;
      320: inst = 32'h10408000;
      321: inst = 32'hc40402f;
      322: inst = 32'h8220000;
      323: inst = 32'h10408000;
      324: inst = 32'hc404030;
      325: inst = 32'h8220000;
      326: inst = 32'h10408000;
      327: inst = 32'hc404031;
      328: inst = 32'h8220000;
      329: inst = 32'h10408000;
      330: inst = 32'hc404032;
      331: inst = 32'h8220000;
      332: inst = 32'h10408000;
      333: inst = 32'hc404033;
      334: inst = 32'h8220000;
      335: inst = 32'h10408000;
      336: inst = 32'hc404034;
      337: inst = 32'h8220000;
      338: inst = 32'h10408000;
      339: inst = 32'hc404035;
      340: inst = 32'h8220000;
      341: inst = 32'h10408000;
      342: inst = 32'hc404036;
      343: inst = 32'h8220000;
      344: inst = 32'h10408000;
      345: inst = 32'hc404037;
      346: inst = 32'h8220000;
      347: inst = 32'h10408000;
      348: inst = 32'hc404038;
      349: inst = 32'h8220000;
      350: inst = 32'h10408000;
      351: inst = 32'hc404039;
      352: inst = 32'h8220000;
      353: inst = 32'h10408000;
      354: inst = 32'hc40403a;
      355: inst = 32'h8220000;
      356: inst = 32'h10408000;
      357: inst = 32'hc40403b;
      358: inst = 32'h8220000;
      359: inst = 32'h10408000;
      360: inst = 32'hc40403c;
      361: inst = 32'h8220000;
      362: inst = 32'h10408000;
      363: inst = 32'hc40403d;
      364: inst = 32'h8220000;
      365: inst = 32'h10408000;
      366: inst = 32'hc40403e;
      367: inst = 32'h8220000;
      368: inst = 32'h10408000;
      369: inst = 32'hc40403f;
      370: inst = 32'h8220000;
      371: inst = 32'h10408000;
      372: inst = 32'hc404040;
      373: inst = 32'h8220000;
      374: inst = 32'h10408000;
      375: inst = 32'hc404041;
      376: inst = 32'h8220000;
      377: inst = 32'h10408000;
      378: inst = 32'hc404042;
      379: inst = 32'h8220000;
      380: inst = 32'h10408000;
      381: inst = 32'hc404043;
      382: inst = 32'h8220000;
      383: inst = 32'h10408000;
      384: inst = 32'hc404044;
      385: inst = 32'h8220000;
      386: inst = 32'h10408000;
      387: inst = 32'hc404045;
      388: inst = 32'h8220000;
      389: inst = 32'h10408000;
      390: inst = 32'hc404046;
      391: inst = 32'h8220000;
      392: inst = 32'h10408000;
      393: inst = 32'hc404047;
      394: inst = 32'h8220000;
      395: inst = 32'h10408000;
      396: inst = 32'hc404048;
      397: inst = 32'h8220000;
      398: inst = 32'h10408000;
      399: inst = 32'hc404049;
      400: inst = 32'h8220000;
      401: inst = 32'h10408000;
      402: inst = 32'hc40404a;
      403: inst = 32'h8220000;
      404: inst = 32'h10408000;
      405: inst = 32'hc40404c;
      406: inst = 32'h8220000;
      407: inst = 32'h10408000;
      408: inst = 32'hc40404d;
      409: inst = 32'h8220000;
      410: inst = 32'h10408000;
      411: inst = 32'hc40404e;
      412: inst = 32'h8220000;
      413: inst = 32'h10408000;
      414: inst = 32'hc40404f;
      415: inst = 32'h8220000;
      416: inst = 32'h10408000;
      417: inst = 32'hc404050;
      418: inst = 32'h8220000;
      419: inst = 32'h10408000;
      420: inst = 32'hc404051;
      421: inst = 32'h8220000;
      422: inst = 32'h10408000;
      423: inst = 32'hc404052;
      424: inst = 32'h8220000;
      425: inst = 32'h10408000;
      426: inst = 32'hc404053;
      427: inst = 32'h8220000;
      428: inst = 32'h10408000;
      429: inst = 32'hc404054;
      430: inst = 32'h8220000;
      431: inst = 32'h10408000;
      432: inst = 32'hc404055;
      433: inst = 32'h8220000;
      434: inst = 32'h10408000;
      435: inst = 32'hc404056;
      436: inst = 32'h8220000;
      437: inst = 32'h10408000;
      438: inst = 32'hc404057;
      439: inst = 32'h8220000;
      440: inst = 32'h10408000;
      441: inst = 32'hc404058;
      442: inst = 32'h8220000;
      443: inst = 32'h10408000;
      444: inst = 32'hc404059;
      445: inst = 32'h8220000;
      446: inst = 32'h10408000;
      447: inst = 32'hc40405a;
      448: inst = 32'h8220000;
      449: inst = 32'h10408000;
      450: inst = 32'hc40405b;
      451: inst = 32'h8220000;
      452: inst = 32'h10408000;
      453: inst = 32'hc40405c;
      454: inst = 32'h8220000;
      455: inst = 32'h10408000;
      456: inst = 32'hc40405d;
      457: inst = 32'h8220000;
      458: inst = 32'h10408000;
      459: inst = 32'hc40405e;
      460: inst = 32'h8220000;
      461: inst = 32'h10408000;
      462: inst = 32'hc40405f;
      463: inst = 32'h8220000;
      464: inst = 32'h10408000;
      465: inst = 32'hc404060;
      466: inst = 32'h8220000;
      467: inst = 32'h10408000;
      468: inst = 32'hc404061;
      469: inst = 32'h8220000;
      470: inst = 32'h10408000;
      471: inst = 32'hc404062;
      472: inst = 32'h8220000;
      473: inst = 32'h10408000;
      474: inst = 32'hc404063;
      475: inst = 32'h8220000;
      476: inst = 32'h10408000;
      477: inst = 32'hc404064;
      478: inst = 32'h8220000;
      479: inst = 32'h10408000;
      480: inst = 32'hc404065;
      481: inst = 32'h8220000;
      482: inst = 32'h10408000;
      483: inst = 32'hc404066;
      484: inst = 32'h8220000;
      485: inst = 32'h10408000;
      486: inst = 32'hc404067;
      487: inst = 32'h8220000;
      488: inst = 32'h10408000;
      489: inst = 32'hc404068;
      490: inst = 32'h8220000;
      491: inst = 32'h10408000;
      492: inst = 32'hc404069;
      493: inst = 32'h8220000;
      494: inst = 32'h10408000;
      495: inst = 32'hc40406a;
      496: inst = 32'h8220000;
      497: inst = 32'h10408000;
      498: inst = 32'hc40406b;
      499: inst = 32'h8220000;
      500: inst = 32'h10408000;
      501: inst = 32'hc40406c;
      502: inst = 32'h8220000;
      503: inst = 32'h10408000;
      504: inst = 32'hc40406d;
      505: inst = 32'h8220000;
      506: inst = 32'h10408000;
      507: inst = 32'hc40406e;
      508: inst = 32'h8220000;
      509: inst = 32'h10408000;
      510: inst = 32'hc40406f;
      511: inst = 32'h8220000;
      512: inst = 32'h10408000;
      513: inst = 32'hc404070;
      514: inst = 32'h8220000;
      515: inst = 32'h10408000;
      516: inst = 32'hc404071;
      517: inst = 32'h8220000;
      518: inst = 32'h10408000;
      519: inst = 32'hc404072;
      520: inst = 32'h8220000;
      521: inst = 32'h10408000;
      522: inst = 32'hc404073;
      523: inst = 32'h8220000;
      524: inst = 32'h10408000;
      525: inst = 32'hc404074;
      526: inst = 32'h8220000;
      527: inst = 32'h10408000;
      528: inst = 32'hc404075;
      529: inst = 32'h8220000;
      530: inst = 32'h10408000;
      531: inst = 32'hc404076;
      532: inst = 32'h8220000;
      533: inst = 32'h10408000;
      534: inst = 32'hc404077;
      535: inst = 32'h8220000;
      536: inst = 32'h10408000;
      537: inst = 32'hc404078;
      538: inst = 32'h8220000;
      539: inst = 32'h10408000;
      540: inst = 32'hc404079;
      541: inst = 32'h8220000;
      542: inst = 32'h10408000;
      543: inst = 32'hc40407a;
      544: inst = 32'h8220000;
      545: inst = 32'h10408000;
      546: inst = 32'hc40407b;
      547: inst = 32'h8220000;
      548: inst = 32'h10408000;
      549: inst = 32'hc40407c;
      550: inst = 32'h8220000;
      551: inst = 32'h10408000;
      552: inst = 32'hc40407d;
      553: inst = 32'h8220000;
      554: inst = 32'h10408000;
      555: inst = 32'hc40407e;
      556: inst = 32'h8220000;
      557: inst = 32'h10408000;
      558: inst = 32'hc40407f;
      559: inst = 32'h8220000;
      560: inst = 32'h10408000;
      561: inst = 32'hc404080;
      562: inst = 32'h8220000;
      563: inst = 32'h10408000;
      564: inst = 32'hc404081;
      565: inst = 32'h8220000;
      566: inst = 32'h10408000;
      567: inst = 32'hc404082;
      568: inst = 32'h8220000;
      569: inst = 32'h10408000;
      570: inst = 32'hc404083;
      571: inst = 32'h8220000;
      572: inst = 32'h10408000;
      573: inst = 32'hc404084;
      574: inst = 32'h8220000;
      575: inst = 32'h10408000;
      576: inst = 32'hc404085;
      577: inst = 32'h8220000;
      578: inst = 32'h10408000;
      579: inst = 32'hc404086;
      580: inst = 32'h8220000;
      581: inst = 32'h10408000;
      582: inst = 32'hc404087;
      583: inst = 32'h8220000;
      584: inst = 32'h10408000;
      585: inst = 32'hc404088;
      586: inst = 32'h8220000;
      587: inst = 32'h10408000;
      588: inst = 32'hc404089;
      589: inst = 32'h8220000;
      590: inst = 32'h10408000;
      591: inst = 32'hc40408a;
      592: inst = 32'h8220000;
      593: inst = 32'h10408000;
      594: inst = 32'hc40408b;
      595: inst = 32'h8220000;
      596: inst = 32'h10408000;
      597: inst = 32'hc40408c;
      598: inst = 32'h8220000;
      599: inst = 32'h10408000;
      600: inst = 32'hc40408d;
      601: inst = 32'h8220000;
      602: inst = 32'h10408000;
      603: inst = 32'hc40408e;
      604: inst = 32'h8220000;
      605: inst = 32'h10408000;
      606: inst = 32'hc40408f;
      607: inst = 32'h8220000;
      608: inst = 32'h10408000;
      609: inst = 32'hc404090;
      610: inst = 32'h8220000;
      611: inst = 32'h10408000;
      612: inst = 32'hc404091;
      613: inst = 32'h8220000;
      614: inst = 32'h10408000;
      615: inst = 32'hc404092;
      616: inst = 32'h8220000;
      617: inst = 32'h10408000;
      618: inst = 32'hc404093;
      619: inst = 32'h8220000;
      620: inst = 32'h10408000;
      621: inst = 32'hc404094;
      622: inst = 32'h8220000;
      623: inst = 32'h10408000;
      624: inst = 32'hc404095;
      625: inst = 32'h8220000;
      626: inst = 32'h10408000;
      627: inst = 32'hc404096;
      628: inst = 32'h8220000;
      629: inst = 32'h10408000;
      630: inst = 32'hc404097;
      631: inst = 32'h8220000;
      632: inst = 32'h10408000;
      633: inst = 32'hc404098;
      634: inst = 32'h8220000;
      635: inst = 32'h10408000;
      636: inst = 32'hc404099;
      637: inst = 32'h8220000;
      638: inst = 32'h10408000;
      639: inst = 32'hc40409a;
      640: inst = 32'h8220000;
      641: inst = 32'h10408000;
      642: inst = 32'hc40409b;
      643: inst = 32'h8220000;
      644: inst = 32'h10408000;
      645: inst = 32'hc40409c;
      646: inst = 32'h8220000;
      647: inst = 32'h10408000;
      648: inst = 32'hc40409d;
      649: inst = 32'h8220000;
      650: inst = 32'h10408000;
      651: inst = 32'hc40409e;
      652: inst = 32'h8220000;
      653: inst = 32'h10408000;
      654: inst = 32'hc40409f;
      655: inst = 32'h8220000;
      656: inst = 32'h10408000;
      657: inst = 32'hc4040a0;
      658: inst = 32'h8220000;
      659: inst = 32'h10408000;
      660: inst = 32'hc4040a1;
      661: inst = 32'h8220000;
      662: inst = 32'h10408000;
      663: inst = 32'hc4040a2;
      664: inst = 32'h8220000;
      665: inst = 32'h10408000;
      666: inst = 32'hc4040a3;
      667: inst = 32'h8220000;
      668: inst = 32'h10408000;
      669: inst = 32'hc4040a4;
      670: inst = 32'h8220000;
      671: inst = 32'h10408000;
      672: inst = 32'hc4040a5;
      673: inst = 32'h8220000;
      674: inst = 32'h10408000;
      675: inst = 32'hc4040a6;
      676: inst = 32'h8220000;
      677: inst = 32'h10408000;
      678: inst = 32'hc4040a7;
      679: inst = 32'h8220000;
      680: inst = 32'h10408000;
      681: inst = 32'hc4040a8;
      682: inst = 32'h8220000;
      683: inst = 32'h10408000;
      684: inst = 32'hc4040a9;
      685: inst = 32'h8220000;
      686: inst = 32'h10408000;
      687: inst = 32'hc4040aa;
      688: inst = 32'h8220000;
      689: inst = 32'h10408000;
      690: inst = 32'hc4040ac;
      691: inst = 32'h8220000;
      692: inst = 32'h10408000;
      693: inst = 32'hc4040ad;
      694: inst = 32'h8220000;
      695: inst = 32'h10408000;
      696: inst = 32'hc4040ae;
      697: inst = 32'h8220000;
      698: inst = 32'h10408000;
      699: inst = 32'hc4040af;
      700: inst = 32'h8220000;
      701: inst = 32'h10408000;
      702: inst = 32'hc4040b0;
      703: inst = 32'h8220000;
      704: inst = 32'h10408000;
      705: inst = 32'hc4040b1;
      706: inst = 32'h8220000;
      707: inst = 32'h10408000;
      708: inst = 32'hc4040b2;
      709: inst = 32'h8220000;
      710: inst = 32'h10408000;
      711: inst = 32'hc4040b3;
      712: inst = 32'h8220000;
      713: inst = 32'h10408000;
      714: inst = 32'hc4040b4;
      715: inst = 32'h8220000;
      716: inst = 32'h10408000;
      717: inst = 32'hc4040b5;
      718: inst = 32'h8220000;
      719: inst = 32'h10408000;
      720: inst = 32'hc4040b6;
      721: inst = 32'h8220000;
      722: inst = 32'h10408000;
      723: inst = 32'hc4040b7;
      724: inst = 32'h8220000;
      725: inst = 32'h10408000;
      726: inst = 32'hc4040b8;
      727: inst = 32'h8220000;
      728: inst = 32'h10408000;
      729: inst = 32'hc4040b9;
      730: inst = 32'h8220000;
      731: inst = 32'h10408000;
      732: inst = 32'hc4040ba;
      733: inst = 32'h8220000;
      734: inst = 32'h10408000;
      735: inst = 32'hc4040bb;
      736: inst = 32'h8220000;
      737: inst = 32'h10408000;
      738: inst = 32'hc4040bc;
      739: inst = 32'h8220000;
      740: inst = 32'h10408000;
      741: inst = 32'hc4040bd;
      742: inst = 32'h8220000;
      743: inst = 32'h10408000;
      744: inst = 32'hc4040be;
      745: inst = 32'h8220000;
      746: inst = 32'h10408000;
      747: inst = 32'hc4040bf;
      748: inst = 32'h8220000;
      749: inst = 32'h10408000;
      750: inst = 32'hc4040c0;
      751: inst = 32'h8220000;
      752: inst = 32'h10408000;
      753: inst = 32'hc4040c1;
      754: inst = 32'h8220000;
      755: inst = 32'h10408000;
      756: inst = 32'hc4040c2;
      757: inst = 32'h8220000;
      758: inst = 32'h10408000;
      759: inst = 32'hc4040c3;
      760: inst = 32'h8220000;
      761: inst = 32'h10408000;
      762: inst = 32'hc4040c4;
      763: inst = 32'h8220000;
      764: inst = 32'h10408000;
      765: inst = 32'hc4040c5;
      766: inst = 32'h8220000;
      767: inst = 32'h10408000;
      768: inst = 32'hc4040c6;
      769: inst = 32'h8220000;
      770: inst = 32'h10408000;
      771: inst = 32'hc4040c7;
      772: inst = 32'h8220000;
      773: inst = 32'h10408000;
      774: inst = 32'hc4040c8;
      775: inst = 32'h8220000;
      776: inst = 32'h10408000;
      777: inst = 32'hc4040c9;
      778: inst = 32'h8220000;
      779: inst = 32'h10408000;
      780: inst = 32'hc4040ca;
      781: inst = 32'h8220000;
      782: inst = 32'h10408000;
      783: inst = 32'hc4040cb;
      784: inst = 32'h8220000;
      785: inst = 32'h10408000;
      786: inst = 32'hc4040cc;
      787: inst = 32'h8220000;
      788: inst = 32'h10408000;
      789: inst = 32'hc4040cd;
      790: inst = 32'h8220000;
      791: inst = 32'h10408000;
      792: inst = 32'hc4040ce;
      793: inst = 32'h8220000;
      794: inst = 32'h10408000;
      795: inst = 32'hc4040cf;
      796: inst = 32'h8220000;
      797: inst = 32'h10408000;
      798: inst = 32'hc4040d0;
      799: inst = 32'h8220000;
      800: inst = 32'h10408000;
      801: inst = 32'hc4040d1;
      802: inst = 32'h8220000;
      803: inst = 32'h10408000;
      804: inst = 32'hc4040d2;
      805: inst = 32'h8220000;
      806: inst = 32'h10408000;
      807: inst = 32'hc4040d3;
      808: inst = 32'h8220000;
      809: inst = 32'h10408000;
      810: inst = 32'hc4040d4;
      811: inst = 32'h8220000;
      812: inst = 32'h10408000;
      813: inst = 32'hc4040d5;
      814: inst = 32'h8220000;
      815: inst = 32'h10408000;
      816: inst = 32'hc4040d6;
      817: inst = 32'h8220000;
      818: inst = 32'h10408000;
      819: inst = 32'hc4040d7;
      820: inst = 32'h8220000;
      821: inst = 32'h10408000;
      822: inst = 32'hc4040d8;
      823: inst = 32'h8220000;
      824: inst = 32'h10408000;
      825: inst = 32'hc4040d9;
      826: inst = 32'h8220000;
      827: inst = 32'h10408000;
      828: inst = 32'hc4040da;
      829: inst = 32'h8220000;
      830: inst = 32'h10408000;
      831: inst = 32'hc4040db;
      832: inst = 32'h8220000;
      833: inst = 32'h10408000;
      834: inst = 32'hc4040dc;
      835: inst = 32'h8220000;
      836: inst = 32'h10408000;
      837: inst = 32'hc4040dd;
      838: inst = 32'h8220000;
      839: inst = 32'h10408000;
      840: inst = 32'hc4040de;
      841: inst = 32'h8220000;
      842: inst = 32'h10408000;
      843: inst = 32'hc4040df;
      844: inst = 32'h8220000;
      845: inst = 32'h10408000;
      846: inst = 32'hc4040e0;
      847: inst = 32'h8220000;
      848: inst = 32'h10408000;
      849: inst = 32'hc4040e1;
      850: inst = 32'h8220000;
      851: inst = 32'h10408000;
      852: inst = 32'hc4040e2;
      853: inst = 32'h8220000;
      854: inst = 32'h10408000;
      855: inst = 32'hc4040e3;
      856: inst = 32'h8220000;
      857: inst = 32'h10408000;
      858: inst = 32'hc4040e4;
      859: inst = 32'h8220000;
      860: inst = 32'h10408000;
      861: inst = 32'hc4040e5;
      862: inst = 32'h8220000;
      863: inst = 32'h10408000;
      864: inst = 32'hc4040e6;
      865: inst = 32'h8220000;
      866: inst = 32'h10408000;
      867: inst = 32'hc4040e7;
      868: inst = 32'h8220000;
      869: inst = 32'h10408000;
      870: inst = 32'hc4040e8;
      871: inst = 32'h8220000;
      872: inst = 32'h10408000;
      873: inst = 32'hc4040e9;
      874: inst = 32'h8220000;
      875: inst = 32'h10408000;
      876: inst = 32'hc4040ea;
      877: inst = 32'h8220000;
      878: inst = 32'h10408000;
      879: inst = 32'hc4040eb;
      880: inst = 32'h8220000;
      881: inst = 32'h10408000;
      882: inst = 32'hc4040ec;
      883: inst = 32'h8220000;
      884: inst = 32'h10408000;
      885: inst = 32'hc4040ed;
      886: inst = 32'h8220000;
      887: inst = 32'h10408000;
      888: inst = 32'hc4040ee;
      889: inst = 32'h8220000;
      890: inst = 32'h10408000;
      891: inst = 32'hc4040ef;
      892: inst = 32'h8220000;
      893: inst = 32'h10408000;
      894: inst = 32'hc4040f0;
      895: inst = 32'h8220000;
      896: inst = 32'h10408000;
      897: inst = 32'hc4040f1;
      898: inst = 32'h8220000;
      899: inst = 32'h10408000;
      900: inst = 32'hc4040f2;
      901: inst = 32'h8220000;
      902: inst = 32'h10408000;
      903: inst = 32'hc4040f3;
      904: inst = 32'h8220000;
      905: inst = 32'h10408000;
      906: inst = 32'hc4040f4;
      907: inst = 32'h8220000;
      908: inst = 32'h10408000;
      909: inst = 32'hc4040f5;
      910: inst = 32'h8220000;
      911: inst = 32'h10408000;
      912: inst = 32'hc4040f6;
      913: inst = 32'h8220000;
      914: inst = 32'h10408000;
      915: inst = 32'hc4040f7;
      916: inst = 32'h8220000;
      917: inst = 32'h10408000;
      918: inst = 32'hc4040f8;
      919: inst = 32'h8220000;
      920: inst = 32'h10408000;
      921: inst = 32'hc4040f9;
      922: inst = 32'h8220000;
      923: inst = 32'h10408000;
      924: inst = 32'hc4040fa;
      925: inst = 32'h8220000;
      926: inst = 32'h10408000;
      927: inst = 32'hc4040fb;
      928: inst = 32'h8220000;
      929: inst = 32'h10408000;
      930: inst = 32'hc4040fc;
      931: inst = 32'h8220000;
      932: inst = 32'h10408000;
      933: inst = 32'hc4040fd;
      934: inst = 32'h8220000;
      935: inst = 32'h10408000;
      936: inst = 32'hc4040fe;
      937: inst = 32'h8220000;
      938: inst = 32'h10408000;
      939: inst = 32'hc4040ff;
      940: inst = 32'h8220000;
      941: inst = 32'h10408000;
      942: inst = 32'hc404100;
      943: inst = 32'h8220000;
      944: inst = 32'h10408000;
      945: inst = 32'hc404101;
      946: inst = 32'h8220000;
      947: inst = 32'h10408000;
      948: inst = 32'hc404102;
      949: inst = 32'h8220000;
      950: inst = 32'h10408000;
      951: inst = 32'hc404103;
      952: inst = 32'h8220000;
      953: inst = 32'h10408000;
      954: inst = 32'hc404104;
      955: inst = 32'h8220000;
      956: inst = 32'h10408000;
      957: inst = 32'hc404105;
      958: inst = 32'h8220000;
      959: inst = 32'h10408000;
      960: inst = 32'hc404106;
      961: inst = 32'h8220000;
      962: inst = 32'h10408000;
      963: inst = 32'hc404107;
      964: inst = 32'h8220000;
      965: inst = 32'h10408000;
      966: inst = 32'hc404108;
      967: inst = 32'h8220000;
      968: inst = 32'h10408000;
      969: inst = 32'hc404109;
      970: inst = 32'h8220000;
      971: inst = 32'h10408000;
      972: inst = 32'hc40410a;
      973: inst = 32'h8220000;
      974: inst = 32'h10408000;
      975: inst = 32'hc40410c;
      976: inst = 32'h8220000;
      977: inst = 32'h10408000;
      978: inst = 32'hc40410d;
      979: inst = 32'h8220000;
      980: inst = 32'h10408000;
      981: inst = 32'hc40410e;
      982: inst = 32'h8220000;
      983: inst = 32'h10408000;
      984: inst = 32'hc40410f;
      985: inst = 32'h8220000;
      986: inst = 32'h10408000;
      987: inst = 32'hc404110;
      988: inst = 32'h8220000;
      989: inst = 32'h10408000;
      990: inst = 32'hc404111;
      991: inst = 32'h8220000;
      992: inst = 32'h10408000;
      993: inst = 32'hc404112;
      994: inst = 32'h8220000;
      995: inst = 32'h10408000;
      996: inst = 32'hc404113;
      997: inst = 32'h8220000;
      998: inst = 32'h10408000;
      999: inst = 32'hc404114;
      1000: inst = 32'h8220000;
      1001: inst = 32'h10408000;
      1002: inst = 32'hc404115;
      1003: inst = 32'h8220000;
      1004: inst = 32'h10408000;
      1005: inst = 32'hc404116;
      1006: inst = 32'h8220000;
      1007: inst = 32'h10408000;
      1008: inst = 32'hc404117;
      1009: inst = 32'h8220000;
      1010: inst = 32'h10408000;
      1011: inst = 32'hc404118;
      1012: inst = 32'h8220000;
      1013: inst = 32'h10408000;
      1014: inst = 32'hc404119;
      1015: inst = 32'h8220000;
      1016: inst = 32'h10408000;
      1017: inst = 32'hc40411a;
      1018: inst = 32'h8220000;
      1019: inst = 32'h10408000;
      1020: inst = 32'hc40411b;
      1021: inst = 32'h8220000;
      1022: inst = 32'h10408000;
      1023: inst = 32'hc40411c;
      1024: inst = 32'h8220000;
      1025: inst = 32'h10408000;
      1026: inst = 32'hc40411d;
      1027: inst = 32'h8220000;
      1028: inst = 32'h10408000;
      1029: inst = 32'hc40411e;
      1030: inst = 32'h8220000;
      1031: inst = 32'h10408000;
      1032: inst = 32'hc40411f;
      1033: inst = 32'h8220000;
      1034: inst = 32'h10408000;
      1035: inst = 32'hc404120;
      1036: inst = 32'h8220000;
      1037: inst = 32'h10408000;
      1038: inst = 32'hc404121;
      1039: inst = 32'h8220000;
      1040: inst = 32'h10408000;
      1041: inst = 32'hc404122;
      1042: inst = 32'h8220000;
      1043: inst = 32'h10408000;
      1044: inst = 32'hc404123;
      1045: inst = 32'h8220000;
      1046: inst = 32'h10408000;
      1047: inst = 32'hc404124;
      1048: inst = 32'h8220000;
      1049: inst = 32'h10408000;
      1050: inst = 32'hc404125;
      1051: inst = 32'h8220000;
      1052: inst = 32'h10408000;
      1053: inst = 32'hc404126;
      1054: inst = 32'h8220000;
      1055: inst = 32'h10408000;
      1056: inst = 32'hc404127;
      1057: inst = 32'h8220000;
      1058: inst = 32'h10408000;
      1059: inst = 32'hc404128;
      1060: inst = 32'h8220000;
      1061: inst = 32'h10408000;
      1062: inst = 32'hc404129;
      1063: inst = 32'h8220000;
      1064: inst = 32'h10408000;
      1065: inst = 32'hc40412a;
      1066: inst = 32'h8220000;
      1067: inst = 32'h10408000;
      1068: inst = 32'hc40412b;
      1069: inst = 32'h8220000;
      1070: inst = 32'h10408000;
      1071: inst = 32'hc40412c;
      1072: inst = 32'h8220000;
      1073: inst = 32'h10408000;
      1074: inst = 32'hc40412d;
      1075: inst = 32'h8220000;
      1076: inst = 32'h10408000;
      1077: inst = 32'hc40412e;
      1078: inst = 32'h8220000;
      1079: inst = 32'h10408000;
      1080: inst = 32'hc40412f;
      1081: inst = 32'h8220000;
      1082: inst = 32'h10408000;
      1083: inst = 32'hc404130;
      1084: inst = 32'h8220000;
      1085: inst = 32'h10408000;
      1086: inst = 32'hc404131;
      1087: inst = 32'h8220000;
      1088: inst = 32'h10408000;
      1089: inst = 32'hc404132;
      1090: inst = 32'h8220000;
      1091: inst = 32'h10408000;
      1092: inst = 32'hc404133;
      1093: inst = 32'h8220000;
      1094: inst = 32'h10408000;
      1095: inst = 32'hc404134;
      1096: inst = 32'h8220000;
      1097: inst = 32'h10408000;
      1098: inst = 32'hc404135;
      1099: inst = 32'h8220000;
      1100: inst = 32'h10408000;
      1101: inst = 32'hc404136;
      1102: inst = 32'h8220000;
      1103: inst = 32'h10408000;
      1104: inst = 32'hc404137;
      1105: inst = 32'h8220000;
      1106: inst = 32'h10408000;
      1107: inst = 32'hc404138;
      1108: inst = 32'h8220000;
      1109: inst = 32'h10408000;
      1110: inst = 32'hc404139;
      1111: inst = 32'h8220000;
      1112: inst = 32'h10408000;
      1113: inst = 32'hc40413a;
      1114: inst = 32'h8220000;
      1115: inst = 32'h10408000;
      1116: inst = 32'hc40413b;
      1117: inst = 32'h8220000;
      1118: inst = 32'h10408000;
      1119: inst = 32'hc40413c;
      1120: inst = 32'h8220000;
      1121: inst = 32'h10408000;
      1122: inst = 32'hc40413d;
      1123: inst = 32'h8220000;
      1124: inst = 32'h10408000;
      1125: inst = 32'hc40413e;
      1126: inst = 32'h8220000;
      1127: inst = 32'h10408000;
      1128: inst = 32'hc40413f;
      1129: inst = 32'h8220000;
      1130: inst = 32'h10408000;
      1131: inst = 32'hc404140;
      1132: inst = 32'h8220000;
      1133: inst = 32'h10408000;
      1134: inst = 32'hc404141;
      1135: inst = 32'h8220000;
      1136: inst = 32'h10408000;
      1137: inst = 32'hc404142;
      1138: inst = 32'h8220000;
      1139: inst = 32'h10408000;
      1140: inst = 32'hc404143;
      1141: inst = 32'h8220000;
      1142: inst = 32'h10408000;
      1143: inst = 32'hc404144;
      1144: inst = 32'h8220000;
      1145: inst = 32'h10408000;
      1146: inst = 32'hc404145;
      1147: inst = 32'h8220000;
      1148: inst = 32'h10408000;
      1149: inst = 32'hc404146;
      1150: inst = 32'h8220000;
      1151: inst = 32'h10408000;
      1152: inst = 32'hc404147;
      1153: inst = 32'h8220000;
      1154: inst = 32'h10408000;
      1155: inst = 32'hc404148;
      1156: inst = 32'h8220000;
      1157: inst = 32'h10408000;
      1158: inst = 32'hc404149;
      1159: inst = 32'h8220000;
      1160: inst = 32'h10408000;
      1161: inst = 32'hc40414a;
      1162: inst = 32'h8220000;
      1163: inst = 32'h10408000;
      1164: inst = 32'hc40414b;
      1165: inst = 32'h8220000;
      1166: inst = 32'h10408000;
      1167: inst = 32'hc40414c;
      1168: inst = 32'h8220000;
      1169: inst = 32'h10408000;
      1170: inst = 32'hc40414d;
      1171: inst = 32'h8220000;
      1172: inst = 32'h10408000;
      1173: inst = 32'hc40414e;
      1174: inst = 32'h8220000;
      1175: inst = 32'h10408000;
      1176: inst = 32'hc40414f;
      1177: inst = 32'h8220000;
      1178: inst = 32'h10408000;
      1179: inst = 32'hc404150;
      1180: inst = 32'h8220000;
      1181: inst = 32'h10408000;
      1182: inst = 32'hc404151;
      1183: inst = 32'h8220000;
      1184: inst = 32'h10408000;
      1185: inst = 32'hc404152;
      1186: inst = 32'h8220000;
      1187: inst = 32'h10408000;
      1188: inst = 32'hc404153;
      1189: inst = 32'h8220000;
      1190: inst = 32'h10408000;
      1191: inst = 32'hc404154;
      1192: inst = 32'h8220000;
      1193: inst = 32'h10408000;
      1194: inst = 32'hc404155;
      1195: inst = 32'h8220000;
      1196: inst = 32'h10408000;
      1197: inst = 32'hc404156;
      1198: inst = 32'h8220000;
      1199: inst = 32'h10408000;
      1200: inst = 32'hc404157;
      1201: inst = 32'h8220000;
      1202: inst = 32'h10408000;
      1203: inst = 32'hc404158;
      1204: inst = 32'h8220000;
      1205: inst = 32'h10408000;
      1206: inst = 32'hc404159;
      1207: inst = 32'h8220000;
      1208: inst = 32'h10408000;
      1209: inst = 32'hc40415a;
      1210: inst = 32'h8220000;
      1211: inst = 32'h10408000;
      1212: inst = 32'hc40415b;
      1213: inst = 32'h8220000;
      1214: inst = 32'h10408000;
      1215: inst = 32'hc40415c;
      1216: inst = 32'h8220000;
      1217: inst = 32'h10408000;
      1218: inst = 32'hc40415d;
      1219: inst = 32'h8220000;
      1220: inst = 32'h10408000;
      1221: inst = 32'hc40415e;
      1222: inst = 32'h8220000;
      1223: inst = 32'h10408000;
      1224: inst = 32'hc40415f;
      1225: inst = 32'h8220000;
      1226: inst = 32'h10408000;
      1227: inst = 32'hc404160;
      1228: inst = 32'h8220000;
      1229: inst = 32'h10408000;
      1230: inst = 32'hc404161;
      1231: inst = 32'h8220000;
      1232: inst = 32'h10408000;
      1233: inst = 32'hc404162;
      1234: inst = 32'h8220000;
      1235: inst = 32'h10408000;
      1236: inst = 32'hc404163;
      1237: inst = 32'h8220000;
      1238: inst = 32'h10408000;
      1239: inst = 32'hc404164;
      1240: inst = 32'h8220000;
      1241: inst = 32'h10408000;
      1242: inst = 32'hc404165;
      1243: inst = 32'h8220000;
      1244: inst = 32'h10408000;
      1245: inst = 32'hc404166;
      1246: inst = 32'h8220000;
      1247: inst = 32'h10408000;
      1248: inst = 32'hc404167;
      1249: inst = 32'h8220000;
      1250: inst = 32'h10408000;
      1251: inst = 32'hc404168;
      1252: inst = 32'h8220000;
      1253: inst = 32'h10408000;
      1254: inst = 32'hc404169;
      1255: inst = 32'h8220000;
      1256: inst = 32'h10408000;
      1257: inst = 32'hc40416a;
      1258: inst = 32'h8220000;
      1259: inst = 32'h10408000;
      1260: inst = 32'hc40416c;
      1261: inst = 32'h8220000;
      1262: inst = 32'h10408000;
      1263: inst = 32'hc40416d;
      1264: inst = 32'h8220000;
      1265: inst = 32'h10408000;
      1266: inst = 32'hc40416e;
      1267: inst = 32'h8220000;
      1268: inst = 32'h10408000;
      1269: inst = 32'hc40416f;
      1270: inst = 32'h8220000;
      1271: inst = 32'h10408000;
      1272: inst = 32'hc404170;
      1273: inst = 32'h8220000;
      1274: inst = 32'h10408000;
      1275: inst = 32'hc404171;
      1276: inst = 32'h8220000;
      1277: inst = 32'h10408000;
      1278: inst = 32'hc404172;
      1279: inst = 32'h8220000;
      1280: inst = 32'h10408000;
      1281: inst = 32'hc404173;
      1282: inst = 32'h8220000;
      1283: inst = 32'h10408000;
      1284: inst = 32'hc404174;
      1285: inst = 32'h8220000;
      1286: inst = 32'h10408000;
      1287: inst = 32'hc404175;
      1288: inst = 32'h8220000;
      1289: inst = 32'h10408000;
      1290: inst = 32'hc404176;
      1291: inst = 32'h8220000;
      1292: inst = 32'h10408000;
      1293: inst = 32'hc404177;
      1294: inst = 32'h8220000;
      1295: inst = 32'h10408000;
      1296: inst = 32'hc404178;
      1297: inst = 32'h8220000;
      1298: inst = 32'h10408000;
      1299: inst = 32'hc404179;
      1300: inst = 32'h8220000;
      1301: inst = 32'h10408000;
      1302: inst = 32'hc40417a;
      1303: inst = 32'h8220000;
      1304: inst = 32'h10408000;
      1305: inst = 32'hc40417b;
      1306: inst = 32'h8220000;
      1307: inst = 32'h10408000;
      1308: inst = 32'hc40417c;
      1309: inst = 32'h8220000;
      1310: inst = 32'h10408000;
      1311: inst = 32'hc40417d;
      1312: inst = 32'h8220000;
      1313: inst = 32'h10408000;
      1314: inst = 32'hc40417e;
      1315: inst = 32'h8220000;
      1316: inst = 32'h10408000;
      1317: inst = 32'hc40417f;
      1318: inst = 32'h8220000;
      1319: inst = 32'h10408000;
      1320: inst = 32'hc404180;
      1321: inst = 32'h8220000;
      1322: inst = 32'h10408000;
      1323: inst = 32'hc404181;
      1324: inst = 32'h8220000;
      1325: inst = 32'h10408000;
      1326: inst = 32'hc404182;
      1327: inst = 32'h8220000;
      1328: inst = 32'h10408000;
      1329: inst = 32'hc404183;
      1330: inst = 32'h8220000;
      1331: inst = 32'h10408000;
      1332: inst = 32'hc404184;
      1333: inst = 32'h8220000;
      1334: inst = 32'h10408000;
      1335: inst = 32'hc404185;
      1336: inst = 32'h8220000;
      1337: inst = 32'h10408000;
      1338: inst = 32'hc404186;
      1339: inst = 32'h8220000;
      1340: inst = 32'h10408000;
      1341: inst = 32'hc404187;
      1342: inst = 32'h8220000;
      1343: inst = 32'h10408000;
      1344: inst = 32'hc404188;
      1345: inst = 32'h8220000;
      1346: inst = 32'h10408000;
      1347: inst = 32'hc404189;
      1348: inst = 32'h8220000;
      1349: inst = 32'h10408000;
      1350: inst = 32'hc40418a;
      1351: inst = 32'h8220000;
      1352: inst = 32'h10408000;
      1353: inst = 32'hc40418b;
      1354: inst = 32'h8220000;
      1355: inst = 32'h10408000;
      1356: inst = 32'hc40418c;
      1357: inst = 32'h8220000;
      1358: inst = 32'h10408000;
      1359: inst = 32'hc40418d;
      1360: inst = 32'h8220000;
      1361: inst = 32'h10408000;
      1362: inst = 32'hc40418e;
      1363: inst = 32'h8220000;
      1364: inst = 32'h10408000;
      1365: inst = 32'hc40418f;
      1366: inst = 32'h8220000;
      1367: inst = 32'h10408000;
      1368: inst = 32'hc404190;
      1369: inst = 32'h8220000;
      1370: inst = 32'h10408000;
      1371: inst = 32'hc404191;
      1372: inst = 32'h8220000;
      1373: inst = 32'h10408000;
      1374: inst = 32'hc404192;
      1375: inst = 32'h8220000;
      1376: inst = 32'h10408000;
      1377: inst = 32'hc404193;
      1378: inst = 32'h8220000;
      1379: inst = 32'h10408000;
      1380: inst = 32'hc404194;
      1381: inst = 32'h8220000;
      1382: inst = 32'h10408000;
      1383: inst = 32'hc404195;
      1384: inst = 32'h8220000;
      1385: inst = 32'h10408000;
      1386: inst = 32'hc404196;
      1387: inst = 32'h8220000;
      1388: inst = 32'h10408000;
      1389: inst = 32'hc404197;
      1390: inst = 32'h8220000;
      1391: inst = 32'h10408000;
      1392: inst = 32'hc404198;
      1393: inst = 32'h8220000;
      1394: inst = 32'h10408000;
      1395: inst = 32'hc404199;
      1396: inst = 32'h8220000;
      1397: inst = 32'h10408000;
      1398: inst = 32'hc40419a;
      1399: inst = 32'h8220000;
      1400: inst = 32'h10408000;
      1401: inst = 32'hc40419b;
      1402: inst = 32'h8220000;
      1403: inst = 32'h10408000;
      1404: inst = 32'hc40419c;
      1405: inst = 32'h8220000;
      1406: inst = 32'h10408000;
      1407: inst = 32'hc40419d;
      1408: inst = 32'h8220000;
      1409: inst = 32'h10408000;
      1410: inst = 32'hc40419e;
      1411: inst = 32'h8220000;
      1412: inst = 32'h10408000;
      1413: inst = 32'hc40419f;
      1414: inst = 32'h8220000;
      1415: inst = 32'h10408000;
      1416: inst = 32'hc4041a0;
      1417: inst = 32'h8220000;
      1418: inst = 32'h10408000;
      1419: inst = 32'hc4041a1;
      1420: inst = 32'h8220000;
      1421: inst = 32'h10408000;
      1422: inst = 32'hc4041a2;
      1423: inst = 32'h8220000;
      1424: inst = 32'h10408000;
      1425: inst = 32'hc4041a3;
      1426: inst = 32'h8220000;
      1427: inst = 32'h10408000;
      1428: inst = 32'hc4041a4;
      1429: inst = 32'h8220000;
      1430: inst = 32'h10408000;
      1431: inst = 32'hc4041a5;
      1432: inst = 32'h8220000;
      1433: inst = 32'h10408000;
      1434: inst = 32'hc4041a6;
      1435: inst = 32'h8220000;
      1436: inst = 32'h10408000;
      1437: inst = 32'hc4041a7;
      1438: inst = 32'h8220000;
      1439: inst = 32'h10408000;
      1440: inst = 32'hc4041a8;
      1441: inst = 32'h8220000;
      1442: inst = 32'h10408000;
      1443: inst = 32'hc4041a9;
      1444: inst = 32'h8220000;
      1445: inst = 32'h10408000;
      1446: inst = 32'hc4041aa;
      1447: inst = 32'h8220000;
      1448: inst = 32'h10408000;
      1449: inst = 32'hc4041ab;
      1450: inst = 32'h8220000;
      1451: inst = 32'h10408000;
      1452: inst = 32'hc4041ac;
      1453: inst = 32'h8220000;
      1454: inst = 32'h10408000;
      1455: inst = 32'hc4041ad;
      1456: inst = 32'h8220000;
      1457: inst = 32'h10408000;
      1458: inst = 32'hc4041ae;
      1459: inst = 32'h8220000;
      1460: inst = 32'h10408000;
      1461: inst = 32'hc4041af;
      1462: inst = 32'h8220000;
      1463: inst = 32'h10408000;
      1464: inst = 32'hc4041b0;
      1465: inst = 32'h8220000;
      1466: inst = 32'h10408000;
      1467: inst = 32'hc4041b1;
      1468: inst = 32'h8220000;
      1469: inst = 32'h10408000;
      1470: inst = 32'hc4041b2;
      1471: inst = 32'h8220000;
      1472: inst = 32'h10408000;
      1473: inst = 32'hc4041b3;
      1474: inst = 32'h8220000;
      1475: inst = 32'h10408000;
      1476: inst = 32'hc4041b4;
      1477: inst = 32'h8220000;
      1478: inst = 32'h10408000;
      1479: inst = 32'hc4041b5;
      1480: inst = 32'h8220000;
      1481: inst = 32'h10408000;
      1482: inst = 32'hc4041b6;
      1483: inst = 32'h8220000;
      1484: inst = 32'h10408000;
      1485: inst = 32'hc4041b7;
      1486: inst = 32'h8220000;
      1487: inst = 32'h10408000;
      1488: inst = 32'hc4041b8;
      1489: inst = 32'h8220000;
      1490: inst = 32'h10408000;
      1491: inst = 32'hc4041b9;
      1492: inst = 32'h8220000;
      1493: inst = 32'h10408000;
      1494: inst = 32'hc4041ba;
      1495: inst = 32'h8220000;
      1496: inst = 32'h10408000;
      1497: inst = 32'hc4041bb;
      1498: inst = 32'h8220000;
      1499: inst = 32'h10408000;
      1500: inst = 32'hc4041bc;
      1501: inst = 32'h8220000;
      1502: inst = 32'h10408000;
      1503: inst = 32'hc4041bd;
      1504: inst = 32'h8220000;
      1505: inst = 32'h10408000;
      1506: inst = 32'hc4041be;
      1507: inst = 32'h8220000;
      1508: inst = 32'h10408000;
      1509: inst = 32'hc4041bf;
      1510: inst = 32'h8220000;
      1511: inst = 32'h10408000;
      1512: inst = 32'hc4041c0;
      1513: inst = 32'h8220000;
      1514: inst = 32'h10408000;
      1515: inst = 32'hc4041c1;
      1516: inst = 32'h8220000;
      1517: inst = 32'h10408000;
      1518: inst = 32'hc4041c2;
      1519: inst = 32'h8220000;
      1520: inst = 32'h10408000;
      1521: inst = 32'hc4041c3;
      1522: inst = 32'h8220000;
      1523: inst = 32'h10408000;
      1524: inst = 32'hc4041c4;
      1525: inst = 32'h8220000;
      1526: inst = 32'h10408000;
      1527: inst = 32'hc4041c5;
      1528: inst = 32'h8220000;
      1529: inst = 32'h10408000;
      1530: inst = 32'hc4041c6;
      1531: inst = 32'h8220000;
      1532: inst = 32'h10408000;
      1533: inst = 32'hc4041c7;
      1534: inst = 32'h8220000;
      1535: inst = 32'h10408000;
      1536: inst = 32'hc4041c8;
      1537: inst = 32'h8220000;
      1538: inst = 32'h10408000;
      1539: inst = 32'hc4041c9;
      1540: inst = 32'h8220000;
      1541: inst = 32'h10408000;
      1542: inst = 32'hc4041ca;
      1543: inst = 32'h8220000;
      1544: inst = 32'h10408000;
      1545: inst = 32'hc4041cc;
      1546: inst = 32'h8220000;
      1547: inst = 32'h10408000;
      1548: inst = 32'hc4041cd;
      1549: inst = 32'h8220000;
      1550: inst = 32'h10408000;
      1551: inst = 32'hc4041ce;
      1552: inst = 32'h8220000;
      1553: inst = 32'h10408000;
      1554: inst = 32'hc4041cf;
      1555: inst = 32'h8220000;
      1556: inst = 32'h10408000;
      1557: inst = 32'hc4041d0;
      1558: inst = 32'h8220000;
      1559: inst = 32'h10408000;
      1560: inst = 32'hc4041d1;
      1561: inst = 32'h8220000;
      1562: inst = 32'h10408000;
      1563: inst = 32'hc4041d2;
      1564: inst = 32'h8220000;
      1565: inst = 32'h10408000;
      1566: inst = 32'hc4041d3;
      1567: inst = 32'h8220000;
      1568: inst = 32'h10408000;
      1569: inst = 32'hc4041d4;
      1570: inst = 32'h8220000;
      1571: inst = 32'h10408000;
      1572: inst = 32'hc4041d5;
      1573: inst = 32'h8220000;
      1574: inst = 32'h10408000;
      1575: inst = 32'hc4041d6;
      1576: inst = 32'h8220000;
      1577: inst = 32'h10408000;
      1578: inst = 32'hc4041d7;
      1579: inst = 32'h8220000;
      1580: inst = 32'h10408000;
      1581: inst = 32'hc4041d8;
      1582: inst = 32'h8220000;
      1583: inst = 32'h10408000;
      1584: inst = 32'hc4041d9;
      1585: inst = 32'h8220000;
      1586: inst = 32'h10408000;
      1587: inst = 32'hc404206;
      1588: inst = 32'h8220000;
      1589: inst = 32'h10408000;
      1590: inst = 32'hc404207;
      1591: inst = 32'h8220000;
      1592: inst = 32'h10408000;
      1593: inst = 32'hc404208;
      1594: inst = 32'h8220000;
      1595: inst = 32'h10408000;
      1596: inst = 32'hc404209;
      1597: inst = 32'h8220000;
      1598: inst = 32'h10408000;
      1599: inst = 32'hc40420a;
      1600: inst = 32'h8220000;
      1601: inst = 32'h10408000;
      1602: inst = 32'hc40420b;
      1603: inst = 32'h8220000;
      1604: inst = 32'h10408000;
      1605: inst = 32'hc40420c;
      1606: inst = 32'h8220000;
      1607: inst = 32'h10408000;
      1608: inst = 32'hc40420d;
      1609: inst = 32'h8220000;
      1610: inst = 32'h10408000;
      1611: inst = 32'hc40420e;
      1612: inst = 32'h8220000;
      1613: inst = 32'h10408000;
      1614: inst = 32'hc40420f;
      1615: inst = 32'h8220000;
      1616: inst = 32'h10408000;
      1617: inst = 32'hc404210;
      1618: inst = 32'h8220000;
      1619: inst = 32'h10408000;
      1620: inst = 32'hc404211;
      1621: inst = 32'h8220000;
      1622: inst = 32'h10408000;
      1623: inst = 32'hc404212;
      1624: inst = 32'h8220000;
      1625: inst = 32'h10408000;
      1626: inst = 32'hc404213;
      1627: inst = 32'h8220000;
      1628: inst = 32'h10408000;
      1629: inst = 32'hc404214;
      1630: inst = 32'h8220000;
      1631: inst = 32'h10408000;
      1632: inst = 32'hc404215;
      1633: inst = 32'h8220000;
      1634: inst = 32'h10408000;
      1635: inst = 32'hc404216;
      1636: inst = 32'h8220000;
      1637: inst = 32'h10408000;
      1638: inst = 32'hc404217;
      1639: inst = 32'h8220000;
      1640: inst = 32'h10408000;
      1641: inst = 32'hc404218;
      1642: inst = 32'h8220000;
      1643: inst = 32'h10408000;
      1644: inst = 32'hc404219;
      1645: inst = 32'h8220000;
      1646: inst = 32'h10408000;
      1647: inst = 32'hc40421a;
      1648: inst = 32'h8220000;
      1649: inst = 32'h10408000;
      1650: inst = 32'hc40421b;
      1651: inst = 32'h8220000;
      1652: inst = 32'h10408000;
      1653: inst = 32'hc40421c;
      1654: inst = 32'h8220000;
      1655: inst = 32'h10408000;
      1656: inst = 32'hc40421d;
      1657: inst = 32'h8220000;
      1658: inst = 32'h10408000;
      1659: inst = 32'hc40421e;
      1660: inst = 32'h8220000;
      1661: inst = 32'h10408000;
      1662: inst = 32'hc40421f;
      1663: inst = 32'h8220000;
      1664: inst = 32'h10408000;
      1665: inst = 32'hc404220;
      1666: inst = 32'h8220000;
      1667: inst = 32'h10408000;
      1668: inst = 32'hc404221;
      1669: inst = 32'h8220000;
      1670: inst = 32'h10408000;
      1671: inst = 32'hc404222;
      1672: inst = 32'h8220000;
      1673: inst = 32'h10408000;
      1674: inst = 32'hc404223;
      1675: inst = 32'h8220000;
      1676: inst = 32'h10408000;
      1677: inst = 32'hc404224;
      1678: inst = 32'h8220000;
      1679: inst = 32'h10408000;
      1680: inst = 32'hc404225;
      1681: inst = 32'h8220000;
      1682: inst = 32'h10408000;
      1683: inst = 32'hc404226;
      1684: inst = 32'h8220000;
      1685: inst = 32'h10408000;
      1686: inst = 32'hc404227;
      1687: inst = 32'h8220000;
      1688: inst = 32'h10408000;
      1689: inst = 32'hc404228;
      1690: inst = 32'h8220000;
      1691: inst = 32'h10408000;
      1692: inst = 32'hc404229;
      1693: inst = 32'h8220000;
      1694: inst = 32'h10408000;
      1695: inst = 32'hc40422a;
      1696: inst = 32'h8220000;
      1697: inst = 32'h10408000;
      1698: inst = 32'hc40422c;
      1699: inst = 32'h8220000;
      1700: inst = 32'h10408000;
      1701: inst = 32'hc40422d;
      1702: inst = 32'h8220000;
      1703: inst = 32'h10408000;
      1704: inst = 32'hc40422e;
      1705: inst = 32'h8220000;
      1706: inst = 32'h10408000;
      1707: inst = 32'hc40422f;
      1708: inst = 32'h8220000;
      1709: inst = 32'h10408000;
      1710: inst = 32'hc404230;
      1711: inst = 32'h8220000;
      1712: inst = 32'h10408000;
      1713: inst = 32'hc404231;
      1714: inst = 32'h8220000;
      1715: inst = 32'h10408000;
      1716: inst = 32'hc404232;
      1717: inst = 32'h8220000;
      1718: inst = 32'h10408000;
      1719: inst = 32'hc404233;
      1720: inst = 32'h8220000;
      1721: inst = 32'h10408000;
      1722: inst = 32'hc404234;
      1723: inst = 32'h8220000;
      1724: inst = 32'h10408000;
      1725: inst = 32'hc404235;
      1726: inst = 32'h8220000;
      1727: inst = 32'h10408000;
      1728: inst = 32'hc404236;
      1729: inst = 32'h8220000;
      1730: inst = 32'h10408000;
      1731: inst = 32'hc404237;
      1732: inst = 32'h8220000;
      1733: inst = 32'h10408000;
      1734: inst = 32'hc404238;
      1735: inst = 32'h8220000;
      1736: inst = 32'h10408000;
      1737: inst = 32'hc404239;
      1738: inst = 32'h8220000;
      1739: inst = 32'h10408000;
      1740: inst = 32'hc40423a;
      1741: inst = 32'h8220000;
      1742: inst = 32'h10408000;
      1743: inst = 32'hc40423b;
      1744: inst = 32'h8220000;
      1745: inst = 32'h10408000;
      1746: inst = 32'hc404264;
      1747: inst = 32'h8220000;
      1748: inst = 32'h10408000;
      1749: inst = 32'hc404265;
      1750: inst = 32'h8220000;
      1751: inst = 32'h10408000;
      1752: inst = 32'hc404266;
      1753: inst = 32'h8220000;
      1754: inst = 32'h10408000;
      1755: inst = 32'hc404267;
      1756: inst = 32'h8220000;
      1757: inst = 32'h10408000;
      1758: inst = 32'hc404268;
      1759: inst = 32'h8220000;
      1760: inst = 32'h10408000;
      1761: inst = 32'hc404269;
      1762: inst = 32'h8220000;
      1763: inst = 32'h10408000;
      1764: inst = 32'hc40426a;
      1765: inst = 32'h8220000;
      1766: inst = 32'h10408000;
      1767: inst = 32'hc40426b;
      1768: inst = 32'h8220000;
      1769: inst = 32'h10408000;
      1770: inst = 32'hc40426c;
      1771: inst = 32'h8220000;
      1772: inst = 32'h10408000;
      1773: inst = 32'hc40426d;
      1774: inst = 32'h8220000;
      1775: inst = 32'h10408000;
      1776: inst = 32'hc40426e;
      1777: inst = 32'h8220000;
      1778: inst = 32'h10408000;
      1779: inst = 32'hc40426f;
      1780: inst = 32'h8220000;
      1781: inst = 32'h10408000;
      1782: inst = 32'hc404270;
      1783: inst = 32'h8220000;
      1784: inst = 32'h10408000;
      1785: inst = 32'hc404271;
      1786: inst = 32'h8220000;
      1787: inst = 32'h10408000;
      1788: inst = 32'hc404272;
      1789: inst = 32'h8220000;
      1790: inst = 32'h10408000;
      1791: inst = 32'hc404273;
      1792: inst = 32'h8220000;
      1793: inst = 32'h10408000;
      1794: inst = 32'hc404274;
      1795: inst = 32'h8220000;
      1796: inst = 32'h10408000;
      1797: inst = 32'hc404275;
      1798: inst = 32'h8220000;
      1799: inst = 32'h10408000;
      1800: inst = 32'hc404276;
      1801: inst = 32'h8220000;
      1802: inst = 32'h10408000;
      1803: inst = 32'hc404277;
      1804: inst = 32'h8220000;
      1805: inst = 32'h10408000;
      1806: inst = 32'hc404278;
      1807: inst = 32'h8220000;
      1808: inst = 32'h10408000;
      1809: inst = 32'hc404279;
      1810: inst = 32'h8220000;
      1811: inst = 32'h10408000;
      1812: inst = 32'hc40427a;
      1813: inst = 32'h8220000;
      1814: inst = 32'h10408000;
      1815: inst = 32'hc40427b;
      1816: inst = 32'h8220000;
      1817: inst = 32'h10408000;
      1818: inst = 32'hc40427c;
      1819: inst = 32'h8220000;
      1820: inst = 32'h10408000;
      1821: inst = 32'hc40427d;
      1822: inst = 32'h8220000;
      1823: inst = 32'h10408000;
      1824: inst = 32'hc40427e;
      1825: inst = 32'h8220000;
      1826: inst = 32'h10408000;
      1827: inst = 32'hc40427f;
      1828: inst = 32'h8220000;
      1829: inst = 32'h10408000;
      1830: inst = 32'hc404280;
      1831: inst = 32'h8220000;
      1832: inst = 32'h10408000;
      1833: inst = 32'hc404281;
      1834: inst = 32'h8220000;
      1835: inst = 32'h10408000;
      1836: inst = 32'hc404282;
      1837: inst = 32'h8220000;
      1838: inst = 32'h10408000;
      1839: inst = 32'hc404283;
      1840: inst = 32'h8220000;
      1841: inst = 32'h10408000;
      1842: inst = 32'hc404284;
      1843: inst = 32'h8220000;
      1844: inst = 32'h10408000;
      1845: inst = 32'hc404285;
      1846: inst = 32'h8220000;
      1847: inst = 32'h10408000;
      1848: inst = 32'hc404286;
      1849: inst = 32'h8220000;
      1850: inst = 32'h10408000;
      1851: inst = 32'hc404287;
      1852: inst = 32'h8220000;
      1853: inst = 32'h10408000;
      1854: inst = 32'hc404288;
      1855: inst = 32'h8220000;
      1856: inst = 32'h10408000;
      1857: inst = 32'hc404289;
      1858: inst = 32'h8220000;
      1859: inst = 32'h10408000;
      1860: inst = 32'hc40428a;
      1861: inst = 32'h8220000;
      1862: inst = 32'h10408000;
      1863: inst = 32'hc40428c;
      1864: inst = 32'h8220000;
      1865: inst = 32'h10408000;
      1866: inst = 32'hc40428d;
      1867: inst = 32'h8220000;
      1868: inst = 32'h10408000;
      1869: inst = 32'hc40428e;
      1870: inst = 32'h8220000;
      1871: inst = 32'h10408000;
      1872: inst = 32'hc40428f;
      1873: inst = 32'h8220000;
      1874: inst = 32'h10408000;
      1875: inst = 32'hc404290;
      1876: inst = 32'h8220000;
      1877: inst = 32'h10408000;
      1878: inst = 32'hc404291;
      1879: inst = 32'h8220000;
      1880: inst = 32'h10408000;
      1881: inst = 32'hc404292;
      1882: inst = 32'h8220000;
      1883: inst = 32'h10408000;
      1884: inst = 32'hc404293;
      1885: inst = 32'h8220000;
      1886: inst = 32'h10408000;
      1887: inst = 32'hc404294;
      1888: inst = 32'h8220000;
      1889: inst = 32'h10408000;
      1890: inst = 32'hc404295;
      1891: inst = 32'h8220000;
      1892: inst = 32'h10408000;
      1893: inst = 32'hc404296;
      1894: inst = 32'h8220000;
      1895: inst = 32'h10408000;
      1896: inst = 32'hc404297;
      1897: inst = 32'h8220000;
      1898: inst = 32'h10408000;
      1899: inst = 32'hc404298;
      1900: inst = 32'h8220000;
      1901: inst = 32'h10408000;
      1902: inst = 32'hc404299;
      1903: inst = 32'h8220000;
      1904: inst = 32'h10408000;
      1905: inst = 32'hc40429a;
      1906: inst = 32'h8220000;
      1907: inst = 32'h10408000;
      1908: inst = 32'hc40429b;
      1909: inst = 32'h8220000;
      1910: inst = 32'h10408000;
      1911: inst = 32'hc4042c4;
      1912: inst = 32'h8220000;
      1913: inst = 32'h10408000;
      1914: inst = 32'hc4042c5;
      1915: inst = 32'h8220000;
      1916: inst = 32'h10408000;
      1917: inst = 32'hc4042c6;
      1918: inst = 32'h8220000;
      1919: inst = 32'h10408000;
      1920: inst = 32'hc4042c7;
      1921: inst = 32'h8220000;
      1922: inst = 32'h10408000;
      1923: inst = 32'hc4042c8;
      1924: inst = 32'h8220000;
      1925: inst = 32'h10408000;
      1926: inst = 32'hc4042c9;
      1927: inst = 32'h8220000;
      1928: inst = 32'h10408000;
      1929: inst = 32'hc4042ca;
      1930: inst = 32'h8220000;
      1931: inst = 32'h10408000;
      1932: inst = 32'hc4042cb;
      1933: inst = 32'h8220000;
      1934: inst = 32'h10408000;
      1935: inst = 32'hc4042cc;
      1936: inst = 32'h8220000;
      1937: inst = 32'h10408000;
      1938: inst = 32'hc4042cd;
      1939: inst = 32'h8220000;
      1940: inst = 32'h10408000;
      1941: inst = 32'hc4042ce;
      1942: inst = 32'h8220000;
      1943: inst = 32'h10408000;
      1944: inst = 32'hc4042cf;
      1945: inst = 32'h8220000;
      1946: inst = 32'h10408000;
      1947: inst = 32'hc4042d0;
      1948: inst = 32'h8220000;
      1949: inst = 32'h10408000;
      1950: inst = 32'hc4042d1;
      1951: inst = 32'h8220000;
      1952: inst = 32'h10408000;
      1953: inst = 32'hc4042d2;
      1954: inst = 32'h8220000;
      1955: inst = 32'h10408000;
      1956: inst = 32'hc4042d3;
      1957: inst = 32'h8220000;
      1958: inst = 32'h10408000;
      1959: inst = 32'hc4042d4;
      1960: inst = 32'h8220000;
      1961: inst = 32'h10408000;
      1962: inst = 32'hc4042d5;
      1963: inst = 32'h8220000;
      1964: inst = 32'h10408000;
      1965: inst = 32'hc4042d6;
      1966: inst = 32'h8220000;
      1967: inst = 32'h10408000;
      1968: inst = 32'hc4042d7;
      1969: inst = 32'h8220000;
      1970: inst = 32'h10408000;
      1971: inst = 32'hc4042d8;
      1972: inst = 32'h8220000;
      1973: inst = 32'h10408000;
      1974: inst = 32'hc4042d9;
      1975: inst = 32'h8220000;
      1976: inst = 32'h10408000;
      1977: inst = 32'hc4042da;
      1978: inst = 32'h8220000;
      1979: inst = 32'h10408000;
      1980: inst = 32'hc4042db;
      1981: inst = 32'h8220000;
      1982: inst = 32'h10408000;
      1983: inst = 32'hc4042dc;
      1984: inst = 32'h8220000;
      1985: inst = 32'h10408000;
      1986: inst = 32'hc4042dd;
      1987: inst = 32'h8220000;
      1988: inst = 32'h10408000;
      1989: inst = 32'hc4042de;
      1990: inst = 32'h8220000;
      1991: inst = 32'h10408000;
      1992: inst = 32'hc4042df;
      1993: inst = 32'h8220000;
      1994: inst = 32'h10408000;
      1995: inst = 32'hc4042e0;
      1996: inst = 32'h8220000;
      1997: inst = 32'h10408000;
      1998: inst = 32'hc4042e1;
      1999: inst = 32'h8220000;
      2000: inst = 32'h10408000;
      2001: inst = 32'hc4042e2;
      2002: inst = 32'h8220000;
      2003: inst = 32'h10408000;
      2004: inst = 32'hc4042e3;
      2005: inst = 32'h8220000;
      2006: inst = 32'h10408000;
      2007: inst = 32'hc4042e4;
      2008: inst = 32'h8220000;
      2009: inst = 32'h10408000;
      2010: inst = 32'hc4042e5;
      2011: inst = 32'h8220000;
      2012: inst = 32'h10408000;
      2013: inst = 32'hc4042e6;
      2014: inst = 32'h8220000;
      2015: inst = 32'h10408000;
      2016: inst = 32'hc4042e7;
      2017: inst = 32'h8220000;
      2018: inst = 32'h10408000;
      2019: inst = 32'hc4042e8;
      2020: inst = 32'h8220000;
      2021: inst = 32'h10408000;
      2022: inst = 32'hc4042e9;
      2023: inst = 32'h8220000;
      2024: inst = 32'h10408000;
      2025: inst = 32'hc4042ee;
      2026: inst = 32'h8220000;
      2027: inst = 32'h10408000;
      2028: inst = 32'hc4042ef;
      2029: inst = 32'h8220000;
      2030: inst = 32'h10408000;
      2031: inst = 32'hc4042f0;
      2032: inst = 32'h8220000;
      2033: inst = 32'h10408000;
      2034: inst = 32'hc4042f1;
      2035: inst = 32'h8220000;
      2036: inst = 32'h10408000;
      2037: inst = 32'hc4042f2;
      2038: inst = 32'h8220000;
      2039: inst = 32'h10408000;
      2040: inst = 32'hc4042f3;
      2041: inst = 32'h8220000;
      2042: inst = 32'h10408000;
      2043: inst = 32'hc4042f4;
      2044: inst = 32'h8220000;
      2045: inst = 32'h10408000;
      2046: inst = 32'hc4042f5;
      2047: inst = 32'h8220000;
      2048: inst = 32'h10408000;
      2049: inst = 32'hc4042f6;
      2050: inst = 32'h8220000;
      2051: inst = 32'h10408000;
      2052: inst = 32'hc4042f7;
      2053: inst = 32'h8220000;
      2054: inst = 32'h10408000;
      2055: inst = 32'hc4042f8;
      2056: inst = 32'h8220000;
      2057: inst = 32'h10408000;
      2058: inst = 32'hc4042f9;
      2059: inst = 32'h8220000;
      2060: inst = 32'h10408000;
      2061: inst = 32'hc4042fa;
      2062: inst = 32'h8220000;
      2063: inst = 32'h10408000;
      2064: inst = 32'hc4042fb;
      2065: inst = 32'h8220000;
      2066: inst = 32'h10408000;
      2067: inst = 32'hc404324;
      2068: inst = 32'h8220000;
      2069: inst = 32'h10408000;
      2070: inst = 32'hc404325;
      2071: inst = 32'h8220000;
      2072: inst = 32'h10408000;
      2073: inst = 32'hc404326;
      2074: inst = 32'h8220000;
      2075: inst = 32'h10408000;
      2076: inst = 32'hc404327;
      2077: inst = 32'h8220000;
      2078: inst = 32'h10408000;
      2079: inst = 32'hc404328;
      2080: inst = 32'h8220000;
      2081: inst = 32'h10408000;
      2082: inst = 32'hc404329;
      2083: inst = 32'h8220000;
      2084: inst = 32'h10408000;
      2085: inst = 32'hc40432a;
      2086: inst = 32'h8220000;
      2087: inst = 32'h10408000;
      2088: inst = 32'hc40432b;
      2089: inst = 32'h8220000;
      2090: inst = 32'h10408000;
      2091: inst = 32'hc40432c;
      2092: inst = 32'h8220000;
      2093: inst = 32'h10408000;
      2094: inst = 32'hc40432d;
      2095: inst = 32'h8220000;
      2096: inst = 32'h10408000;
      2097: inst = 32'hc40432e;
      2098: inst = 32'h8220000;
      2099: inst = 32'h10408000;
      2100: inst = 32'hc40432f;
      2101: inst = 32'h8220000;
      2102: inst = 32'h10408000;
      2103: inst = 32'hc404330;
      2104: inst = 32'h8220000;
      2105: inst = 32'h10408000;
      2106: inst = 32'hc404331;
      2107: inst = 32'h8220000;
      2108: inst = 32'h10408000;
      2109: inst = 32'hc404332;
      2110: inst = 32'h8220000;
      2111: inst = 32'h10408000;
      2112: inst = 32'hc404333;
      2113: inst = 32'h8220000;
      2114: inst = 32'h10408000;
      2115: inst = 32'hc404334;
      2116: inst = 32'h8220000;
      2117: inst = 32'h10408000;
      2118: inst = 32'hc404335;
      2119: inst = 32'h8220000;
      2120: inst = 32'h10408000;
      2121: inst = 32'hc404336;
      2122: inst = 32'h8220000;
      2123: inst = 32'h10408000;
      2124: inst = 32'hc404337;
      2125: inst = 32'h8220000;
      2126: inst = 32'h10408000;
      2127: inst = 32'hc404338;
      2128: inst = 32'h8220000;
      2129: inst = 32'h10408000;
      2130: inst = 32'hc404339;
      2131: inst = 32'h8220000;
      2132: inst = 32'h10408000;
      2133: inst = 32'hc40433a;
      2134: inst = 32'h8220000;
      2135: inst = 32'h10408000;
      2136: inst = 32'hc40433b;
      2137: inst = 32'h8220000;
      2138: inst = 32'h10408000;
      2139: inst = 32'hc40433c;
      2140: inst = 32'h8220000;
      2141: inst = 32'h10408000;
      2142: inst = 32'hc40433d;
      2143: inst = 32'h8220000;
      2144: inst = 32'h10408000;
      2145: inst = 32'hc40433e;
      2146: inst = 32'h8220000;
      2147: inst = 32'h10408000;
      2148: inst = 32'hc40433f;
      2149: inst = 32'h8220000;
      2150: inst = 32'h10408000;
      2151: inst = 32'hc404340;
      2152: inst = 32'h8220000;
      2153: inst = 32'h10408000;
      2154: inst = 32'hc404341;
      2155: inst = 32'h8220000;
      2156: inst = 32'h10408000;
      2157: inst = 32'hc404342;
      2158: inst = 32'h8220000;
      2159: inst = 32'h10408000;
      2160: inst = 32'hc404343;
      2161: inst = 32'h8220000;
      2162: inst = 32'h10408000;
      2163: inst = 32'hc404344;
      2164: inst = 32'h8220000;
      2165: inst = 32'h10408000;
      2166: inst = 32'hc404345;
      2167: inst = 32'h8220000;
      2168: inst = 32'h10408000;
      2169: inst = 32'hc404346;
      2170: inst = 32'h8220000;
      2171: inst = 32'h10408000;
      2172: inst = 32'hc404347;
      2173: inst = 32'h8220000;
      2174: inst = 32'h10408000;
      2175: inst = 32'hc404348;
      2176: inst = 32'h8220000;
      2177: inst = 32'h10408000;
      2178: inst = 32'hc40434f;
      2179: inst = 32'h8220000;
      2180: inst = 32'h10408000;
      2181: inst = 32'hc404350;
      2182: inst = 32'h8220000;
      2183: inst = 32'h10408000;
      2184: inst = 32'hc404351;
      2185: inst = 32'h8220000;
      2186: inst = 32'h10408000;
      2187: inst = 32'hc404352;
      2188: inst = 32'h8220000;
      2189: inst = 32'h10408000;
      2190: inst = 32'hc404353;
      2191: inst = 32'h8220000;
      2192: inst = 32'h10408000;
      2193: inst = 32'hc404354;
      2194: inst = 32'h8220000;
      2195: inst = 32'h10408000;
      2196: inst = 32'hc404355;
      2197: inst = 32'h8220000;
      2198: inst = 32'h10408000;
      2199: inst = 32'hc404356;
      2200: inst = 32'h8220000;
      2201: inst = 32'h10408000;
      2202: inst = 32'hc404357;
      2203: inst = 32'h8220000;
      2204: inst = 32'h10408000;
      2205: inst = 32'hc404358;
      2206: inst = 32'h8220000;
      2207: inst = 32'h10408000;
      2208: inst = 32'hc404359;
      2209: inst = 32'h8220000;
      2210: inst = 32'h10408000;
      2211: inst = 32'hc40435a;
      2212: inst = 32'h8220000;
      2213: inst = 32'h10408000;
      2214: inst = 32'hc40435b;
      2215: inst = 32'h8220000;
      2216: inst = 32'h10408000;
      2217: inst = 32'hc404384;
      2218: inst = 32'h8220000;
      2219: inst = 32'h10408000;
      2220: inst = 32'hc404385;
      2221: inst = 32'h8220000;
      2222: inst = 32'h10408000;
      2223: inst = 32'hc404386;
      2224: inst = 32'h8220000;
      2225: inst = 32'h10408000;
      2226: inst = 32'hc404387;
      2227: inst = 32'h8220000;
      2228: inst = 32'h10408000;
      2229: inst = 32'hc404388;
      2230: inst = 32'h8220000;
      2231: inst = 32'h10408000;
      2232: inst = 32'hc404389;
      2233: inst = 32'h8220000;
      2234: inst = 32'h10408000;
      2235: inst = 32'hc40438a;
      2236: inst = 32'h8220000;
      2237: inst = 32'h10408000;
      2238: inst = 32'hc40438b;
      2239: inst = 32'h8220000;
      2240: inst = 32'h10408000;
      2241: inst = 32'hc40438c;
      2242: inst = 32'h8220000;
      2243: inst = 32'h10408000;
      2244: inst = 32'hc40438d;
      2245: inst = 32'h8220000;
      2246: inst = 32'h10408000;
      2247: inst = 32'hc40438e;
      2248: inst = 32'h8220000;
      2249: inst = 32'h10408000;
      2250: inst = 32'hc40438f;
      2251: inst = 32'h8220000;
      2252: inst = 32'h10408000;
      2253: inst = 32'hc404390;
      2254: inst = 32'h8220000;
      2255: inst = 32'h10408000;
      2256: inst = 32'hc404391;
      2257: inst = 32'h8220000;
      2258: inst = 32'h10408000;
      2259: inst = 32'hc404392;
      2260: inst = 32'h8220000;
      2261: inst = 32'h10408000;
      2262: inst = 32'hc404393;
      2263: inst = 32'h8220000;
      2264: inst = 32'h10408000;
      2265: inst = 32'hc404394;
      2266: inst = 32'h8220000;
      2267: inst = 32'h10408000;
      2268: inst = 32'hc404395;
      2269: inst = 32'h8220000;
      2270: inst = 32'h10408000;
      2271: inst = 32'hc404396;
      2272: inst = 32'h8220000;
      2273: inst = 32'h10408000;
      2274: inst = 32'hc404397;
      2275: inst = 32'h8220000;
      2276: inst = 32'h10408000;
      2277: inst = 32'hc404398;
      2278: inst = 32'h8220000;
      2279: inst = 32'h10408000;
      2280: inst = 32'hc404399;
      2281: inst = 32'h8220000;
      2282: inst = 32'h10408000;
      2283: inst = 32'hc40439a;
      2284: inst = 32'h8220000;
      2285: inst = 32'h10408000;
      2286: inst = 32'hc40439b;
      2287: inst = 32'h8220000;
      2288: inst = 32'h10408000;
      2289: inst = 32'hc40439c;
      2290: inst = 32'h8220000;
      2291: inst = 32'h10408000;
      2292: inst = 32'hc40439d;
      2293: inst = 32'h8220000;
      2294: inst = 32'h10408000;
      2295: inst = 32'hc40439e;
      2296: inst = 32'h8220000;
      2297: inst = 32'h10408000;
      2298: inst = 32'hc40439f;
      2299: inst = 32'h8220000;
      2300: inst = 32'h10408000;
      2301: inst = 32'hc4043a0;
      2302: inst = 32'h8220000;
      2303: inst = 32'h10408000;
      2304: inst = 32'hc4043a1;
      2305: inst = 32'h8220000;
      2306: inst = 32'h10408000;
      2307: inst = 32'hc4043a2;
      2308: inst = 32'h8220000;
      2309: inst = 32'h10408000;
      2310: inst = 32'hc4043a3;
      2311: inst = 32'h8220000;
      2312: inst = 32'h10408000;
      2313: inst = 32'hc4043a4;
      2314: inst = 32'h8220000;
      2315: inst = 32'h10408000;
      2316: inst = 32'hc4043a5;
      2317: inst = 32'h8220000;
      2318: inst = 32'h10408000;
      2319: inst = 32'hc4043a6;
      2320: inst = 32'h8220000;
      2321: inst = 32'h10408000;
      2322: inst = 32'hc4043b1;
      2323: inst = 32'h8220000;
      2324: inst = 32'h10408000;
      2325: inst = 32'hc4043b2;
      2326: inst = 32'h8220000;
      2327: inst = 32'h10408000;
      2328: inst = 32'hc4043b3;
      2329: inst = 32'h8220000;
      2330: inst = 32'h10408000;
      2331: inst = 32'hc4043b4;
      2332: inst = 32'h8220000;
      2333: inst = 32'h10408000;
      2334: inst = 32'hc4043b5;
      2335: inst = 32'h8220000;
      2336: inst = 32'h10408000;
      2337: inst = 32'hc4043b6;
      2338: inst = 32'h8220000;
      2339: inst = 32'h10408000;
      2340: inst = 32'hc4043b7;
      2341: inst = 32'h8220000;
      2342: inst = 32'h10408000;
      2343: inst = 32'hc4043b8;
      2344: inst = 32'h8220000;
      2345: inst = 32'h10408000;
      2346: inst = 32'hc4043b9;
      2347: inst = 32'h8220000;
      2348: inst = 32'h10408000;
      2349: inst = 32'hc4043ba;
      2350: inst = 32'h8220000;
      2351: inst = 32'h10408000;
      2352: inst = 32'hc4043bb;
      2353: inst = 32'h8220000;
      2354: inst = 32'h10408000;
      2355: inst = 32'hc4043e4;
      2356: inst = 32'h8220000;
      2357: inst = 32'h10408000;
      2358: inst = 32'hc4043e5;
      2359: inst = 32'h8220000;
      2360: inst = 32'h10408000;
      2361: inst = 32'hc4043e6;
      2362: inst = 32'h8220000;
      2363: inst = 32'h10408000;
      2364: inst = 32'hc4043e7;
      2365: inst = 32'h8220000;
      2366: inst = 32'h10408000;
      2367: inst = 32'hc4043e8;
      2368: inst = 32'h8220000;
      2369: inst = 32'h10408000;
      2370: inst = 32'hc4043e9;
      2371: inst = 32'h8220000;
      2372: inst = 32'h10408000;
      2373: inst = 32'hc4043ea;
      2374: inst = 32'h8220000;
      2375: inst = 32'h10408000;
      2376: inst = 32'hc4043eb;
      2377: inst = 32'h8220000;
      2378: inst = 32'h10408000;
      2379: inst = 32'hc4043ec;
      2380: inst = 32'h8220000;
      2381: inst = 32'h10408000;
      2382: inst = 32'hc4043ed;
      2383: inst = 32'h8220000;
      2384: inst = 32'h10408000;
      2385: inst = 32'hc4043ee;
      2386: inst = 32'h8220000;
      2387: inst = 32'h10408000;
      2388: inst = 32'hc4043ef;
      2389: inst = 32'h8220000;
      2390: inst = 32'h10408000;
      2391: inst = 32'hc4043f0;
      2392: inst = 32'h8220000;
      2393: inst = 32'h10408000;
      2394: inst = 32'hc4043f1;
      2395: inst = 32'h8220000;
      2396: inst = 32'h10408000;
      2397: inst = 32'hc4043f2;
      2398: inst = 32'h8220000;
      2399: inst = 32'h10408000;
      2400: inst = 32'hc4043f3;
      2401: inst = 32'h8220000;
      2402: inst = 32'h10408000;
      2403: inst = 32'hc4043f4;
      2404: inst = 32'h8220000;
      2405: inst = 32'h10408000;
      2406: inst = 32'hc4043f5;
      2407: inst = 32'h8220000;
      2408: inst = 32'h10408000;
      2409: inst = 32'hc4043f6;
      2410: inst = 32'h8220000;
      2411: inst = 32'h10408000;
      2412: inst = 32'hc4043f7;
      2413: inst = 32'h8220000;
      2414: inst = 32'h10408000;
      2415: inst = 32'hc4043f8;
      2416: inst = 32'h8220000;
      2417: inst = 32'h10408000;
      2418: inst = 32'hc4043f9;
      2419: inst = 32'h8220000;
      2420: inst = 32'h10408000;
      2421: inst = 32'hc4043fa;
      2422: inst = 32'h8220000;
      2423: inst = 32'h10408000;
      2424: inst = 32'hc4043fb;
      2425: inst = 32'h8220000;
      2426: inst = 32'h10408000;
      2427: inst = 32'hc4043fc;
      2428: inst = 32'h8220000;
      2429: inst = 32'h10408000;
      2430: inst = 32'hc4043fd;
      2431: inst = 32'h8220000;
      2432: inst = 32'h10408000;
      2433: inst = 32'hc4043fe;
      2434: inst = 32'h8220000;
      2435: inst = 32'h10408000;
      2436: inst = 32'hc4043ff;
      2437: inst = 32'h8220000;
      2438: inst = 32'h10408000;
      2439: inst = 32'hc404400;
      2440: inst = 32'h8220000;
      2441: inst = 32'h10408000;
      2442: inst = 32'hc404401;
      2443: inst = 32'h8220000;
      2444: inst = 32'h10408000;
      2445: inst = 32'hc404402;
      2446: inst = 32'h8220000;
      2447: inst = 32'h10408000;
      2448: inst = 32'hc404403;
      2449: inst = 32'h8220000;
      2450: inst = 32'h10408000;
      2451: inst = 32'hc404404;
      2452: inst = 32'h8220000;
      2453: inst = 32'h10408000;
      2454: inst = 32'hc404405;
      2455: inst = 32'h8220000;
      2456: inst = 32'h10408000;
      2457: inst = 32'hc404412;
      2458: inst = 32'h8220000;
      2459: inst = 32'h10408000;
      2460: inst = 32'hc404413;
      2461: inst = 32'h8220000;
      2462: inst = 32'h10408000;
      2463: inst = 32'hc404414;
      2464: inst = 32'h8220000;
      2465: inst = 32'h10408000;
      2466: inst = 32'hc404415;
      2467: inst = 32'h8220000;
      2468: inst = 32'h10408000;
      2469: inst = 32'hc404416;
      2470: inst = 32'h8220000;
      2471: inst = 32'h10408000;
      2472: inst = 32'hc404417;
      2473: inst = 32'h8220000;
      2474: inst = 32'h10408000;
      2475: inst = 32'hc404418;
      2476: inst = 32'h8220000;
      2477: inst = 32'h10408000;
      2478: inst = 32'hc404419;
      2479: inst = 32'h8220000;
      2480: inst = 32'h10408000;
      2481: inst = 32'hc40441a;
      2482: inst = 32'h8220000;
      2483: inst = 32'h10408000;
      2484: inst = 32'hc40441b;
      2485: inst = 32'h8220000;
      2486: inst = 32'h10408000;
      2487: inst = 32'hc404444;
      2488: inst = 32'h8220000;
      2489: inst = 32'h10408000;
      2490: inst = 32'hc404445;
      2491: inst = 32'h8220000;
      2492: inst = 32'h10408000;
      2493: inst = 32'hc404446;
      2494: inst = 32'h8220000;
      2495: inst = 32'h10408000;
      2496: inst = 32'hc404447;
      2497: inst = 32'h8220000;
      2498: inst = 32'h10408000;
      2499: inst = 32'hc404448;
      2500: inst = 32'h8220000;
      2501: inst = 32'h10408000;
      2502: inst = 32'hc404449;
      2503: inst = 32'h8220000;
      2504: inst = 32'h10408000;
      2505: inst = 32'hc40444a;
      2506: inst = 32'h8220000;
      2507: inst = 32'h10408000;
      2508: inst = 32'hc40444b;
      2509: inst = 32'h8220000;
      2510: inst = 32'h10408000;
      2511: inst = 32'hc40444c;
      2512: inst = 32'h8220000;
      2513: inst = 32'h10408000;
      2514: inst = 32'hc40444d;
      2515: inst = 32'h8220000;
      2516: inst = 32'h10408000;
      2517: inst = 32'hc40444e;
      2518: inst = 32'h8220000;
      2519: inst = 32'h10408000;
      2520: inst = 32'hc40444f;
      2521: inst = 32'h8220000;
      2522: inst = 32'h10408000;
      2523: inst = 32'hc404450;
      2524: inst = 32'h8220000;
      2525: inst = 32'h10408000;
      2526: inst = 32'hc404451;
      2527: inst = 32'h8220000;
      2528: inst = 32'h10408000;
      2529: inst = 32'hc404452;
      2530: inst = 32'h8220000;
      2531: inst = 32'h10408000;
      2532: inst = 32'hc404453;
      2533: inst = 32'h8220000;
      2534: inst = 32'h10408000;
      2535: inst = 32'hc404454;
      2536: inst = 32'h8220000;
      2537: inst = 32'h10408000;
      2538: inst = 32'hc404455;
      2539: inst = 32'h8220000;
      2540: inst = 32'h10408000;
      2541: inst = 32'hc404456;
      2542: inst = 32'h8220000;
      2543: inst = 32'h10408000;
      2544: inst = 32'hc404457;
      2545: inst = 32'h8220000;
      2546: inst = 32'h10408000;
      2547: inst = 32'hc404458;
      2548: inst = 32'h8220000;
      2549: inst = 32'h10408000;
      2550: inst = 32'hc404459;
      2551: inst = 32'h8220000;
      2552: inst = 32'h10408000;
      2553: inst = 32'hc40445a;
      2554: inst = 32'h8220000;
      2555: inst = 32'h10408000;
      2556: inst = 32'hc40445b;
      2557: inst = 32'h8220000;
      2558: inst = 32'h10408000;
      2559: inst = 32'hc40445c;
      2560: inst = 32'h8220000;
      2561: inst = 32'h10408000;
      2562: inst = 32'hc40445d;
      2563: inst = 32'h8220000;
      2564: inst = 32'h10408000;
      2565: inst = 32'hc40445e;
      2566: inst = 32'h8220000;
      2567: inst = 32'h10408000;
      2568: inst = 32'hc40445f;
      2569: inst = 32'h8220000;
      2570: inst = 32'h10408000;
      2571: inst = 32'hc404460;
      2572: inst = 32'h8220000;
      2573: inst = 32'h10408000;
      2574: inst = 32'hc404461;
      2575: inst = 32'h8220000;
      2576: inst = 32'h10408000;
      2577: inst = 32'hc404462;
      2578: inst = 32'h8220000;
      2579: inst = 32'h10408000;
      2580: inst = 32'hc404463;
      2581: inst = 32'h8220000;
      2582: inst = 32'h10408000;
      2583: inst = 32'hc404464;
      2584: inst = 32'h8220000;
      2585: inst = 32'h10408000;
      2586: inst = 32'hc404465;
      2587: inst = 32'h8220000;
      2588: inst = 32'h10408000;
      2589: inst = 32'hc404466;
      2590: inst = 32'h8220000;
      2591: inst = 32'h10408000;
      2592: inst = 32'hc404467;
      2593: inst = 32'h8220000;
      2594: inst = 32'h10408000;
      2595: inst = 32'hc404468;
      2596: inst = 32'h8220000;
      2597: inst = 32'h10408000;
      2598: inst = 32'hc404469;
      2599: inst = 32'h8220000;
      2600: inst = 32'h10408000;
      2601: inst = 32'hc40446e;
      2602: inst = 32'h8220000;
      2603: inst = 32'h10408000;
      2604: inst = 32'hc40446f;
      2605: inst = 32'h8220000;
      2606: inst = 32'h10408000;
      2607: inst = 32'hc404470;
      2608: inst = 32'h8220000;
      2609: inst = 32'h10408000;
      2610: inst = 32'hc404471;
      2611: inst = 32'h8220000;
      2612: inst = 32'h10408000;
      2613: inst = 32'hc404472;
      2614: inst = 32'h8220000;
      2615: inst = 32'h10408000;
      2616: inst = 32'hc404473;
      2617: inst = 32'h8220000;
      2618: inst = 32'h10408000;
      2619: inst = 32'hc404474;
      2620: inst = 32'h8220000;
      2621: inst = 32'h10408000;
      2622: inst = 32'hc404475;
      2623: inst = 32'h8220000;
      2624: inst = 32'h10408000;
      2625: inst = 32'hc404476;
      2626: inst = 32'h8220000;
      2627: inst = 32'h10408000;
      2628: inst = 32'hc404477;
      2629: inst = 32'h8220000;
      2630: inst = 32'h10408000;
      2631: inst = 32'hc404478;
      2632: inst = 32'h8220000;
      2633: inst = 32'h10408000;
      2634: inst = 32'hc404479;
      2635: inst = 32'h8220000;
      2636: inst = 32'h10408000;
      2637: inst = 32'hc40447a;
      2638: inst = 32'h8220000;
      2639: inst = 32'h10408000;
      2640: inst = 32'hc40447b;
      2641: inst = 32'h8220000;
      2642: inst = 32'h10408000;
      2643: inst = 32'hc4044a4;
      2644: inst = 32'h8220000;
      2645: inst = 32'h10408000;
      2646: inst = 32'hc4044a5;
      2647: inst = 32'h8220000;
      2648: inst = 32'h10408000;
      2649: inst = 32'hc4044a6;
      2650: inst = 32'h8220000;
      2651: inst = 32'h10408000;
      2652: inst = 32'hc4044a7;
      2653: inst = 32'h8220000;
      2654: inst = 32'h10408000;
      2655: inst = 32'hc4044a8;
      2656: inst = 32'h8220000;
      2657: inst = 32'h10408000;
      2658: inst = 32'hc4044a9;
      2659: inst = 32'h8220000;
      2660: inst = 32'h10408000;
      2661: inst = 32'hc4044aa;
      2662: inst = 32'h8220000;
      2663: inst = 32'h10408000;
      2664: inst = 32'hc4044ab;
      2665: inst = 32'h8220000;
      2666: inst = 32'h10408000;
      2667: inst = 32'hc4044ac;
      2668: inst = 32'h8220000;
      2669: inst = 32'h10408000;
      2670: inst = 32'hc4044ad;
      2671: inst = 32'h8220000;
      2672: inst = 32'h10408000;
      2673: inst = 32'hc4044ae;
      2674: inst = 32'h8220000;
      2675: inst = 32'h10408000;
      2676: inst = 32'hc4044af;
      2677: inst = 32'h8220000;
      2678: inst = 32'h10408000;
      2679: inst = 32'hc4044b0;
      2680: inst = 32'h8220000;
      2681: inst = 32'h10408000;
      2682: inst = 32'hc4044b1;
      2683: inst = 32'h8220000;
      2684: inst = 32'h10408000;
      2685: inst = 32'hc4044b6;
      2686: inst = 32'h8220000;
      2687: inst = 32'h10408000;
      2688: inst = 32'hc4044b7;
      2689: inst = 32'h8220000;
      2690: inst = 32'h10408000;
      2691: inst = 32'hc4044b8;
      2692: inst = 32'h8220000;
      2693: inst = 32'h10408000;
      2694: inst = 32'hc4044b9;
      2695: inst = 32'h8220000;
      2696: inst = 32'h10408000;
      2697: inst = 32'hc4044ba;
      2698: inst = 32'h8220000;
      2699: inst = 32'h10408000;
      2700: inst = 32'hc4044bb;
      2701: inst = 32'h8220000;
      2702: inst = 32'h10408000;
      2703: inst = 32'hc4044bc;
      2704: inst = 32'h8220000;
      2705: inst = 32'h10408000;
      2706: inst = 32'hc4044bd;
      2707: inst = 32'h8220000;
      2708: inst = 32'h10408000;
      2709: inst = 32'hc4044be;
      2710: inst = 32'h8220000;
      2711: inst = 32'h10408000;
      2712: inst = 32'hc4044bf;
      2713: inst = 32'h8220000;
      2714: inst = 32'h10408000;
      2715: inst = 32'hc4044c0;
      2716: inst = 32'h8220000;
      2717: inst = 32'h10408000;
      2718: inst = 32'hc4044c1;
      2719: inst = 32'h8220000;
      2720: inst = 32'h10408000;
      2721: inst = 32'hc4044c2;
      2722: inst = 32'h8220000;
      2723: inst = 32'h10408000;
      2724: inst = 32'hc4044c3;
      2725: inst = 32'h8220000;
      2726: inst = 32'h10408000;
      2727: inst = 32'hc4044c4;
      2728: inst = 32'h8220000;
      2729: inst = 32'h10408000;
      2730: inst = 32'hc4044c5;
      2731: inst = 32'h8220000;
      2732: inst = 32'h10408000;
      2733: inst = 32'hc4044c6;
      2734: inst = 32'h8220000;
      2735: inst = 32'h10408000;
      2736: inst = 32'hc4044c7;
      2737: inst = 32'h8220000;
      2738: inst = 32'h10408000;
      2739: inst = 32'hc4044c8;
      2740: inst = 32'h8220000;
      2741: inst = 32'h10408000;
      2742: inst = 32'hc4044c9;
      2743: inst = 32'h8220000;
      2744: inst = 32'h10408000;
      2745: inst = 32'hc4044ca;
      2746: inst = 32'h8220000;
      2747: inst = 32'h10408000;
      2748: inst = 32'hc4044cd;
      2749: inst = 32'h8220000;
      2750: inst = 32'h10408000;
      2751: inst = 32'hc4044ce;
      2752: inst = 32'h8220000;
      2753: inst = 32'h10408000;
      2754: inst = 32'hc4044cf;
      2755: inst = 32'h8220000;
      2756: inst = 32'h10408000;
      2757: inst = 32'hc4044d0;
      2758: inst = 32'h8220000;
      2759: inst = 32'h10408000;
      2760: inst = 32'hc4044d1;
      2761: inst = 32'h8220000;
      2762: inst = 32'h10408000;
      2763: inst = 32'hc4044d2;
      2764: inst = 32'h8220000;
      2765: inst = 32'h10408000;
      2766: inst = 32'hc4044d3;
      2767: inst = 32'h8220000;
      2768: inst = 32'h10408000;
      2769: inst = 32'hc4044d4;
      2770: inst = 32'h8220000;
      2771: inst = 32'h10408000;
      2772: inst = 32'hc4044d5;
      2773: inst = 32'h8220000;
      2774: inst = 32'h10408000;
      2775: inst = 32'hc4044d6;
      2776: inst = 32'h8220000;
      2777: inst = 32'h10408000;
      2778: inst = 32'hc4044d7;
      2779: inst = 32'h8220000;
      2780: inst = 32'h10408000;
      2781: inst = 32'hc4044d8;
      2782: inst = 32'h8220000;
      2783: inst = 32'h10408000;
      2784: inst = 32'hc4044d9;
      2785: inst = 32'h8220000;
      2786: inst = 32'h10408000;
      2787: inst = 32'hc4044da;
      2788: inst = 32'h8220000;
      2789: inst = 32'h10408000;
      2790: inst = 32'hc4044db;
      2791: inst = 32'h8220000;
      2792: inst = 32'h10408000;
      2793: inst = 32'hc404504;
      2794: inst = 32'h8220000;
      2795: inst = 32'h10408000;
      2796: inst = 32'hc404505;
      2797: inst = 32'h8220000;
      2798: inst = 32'h10408000;
      2799: inst = 32'hc404506;
      2800: inst = 32'h8220000;
      2801: inst = 32'h10408000;
      2802: inst = 32'hc404507;
      2803: inst = 32'h8220000;
      2804: inst = 32'h10408000;
      2805: inst = 32'hc404508;
      2806: inst = 32'h8220000;
      2807: inst = 32'h10408000;
      2808: inst = 32'hc404509;
      2809: inst = 32'h8220000;
      2810: inst = 32'h10408000;
      2811: inst = 32'hc40450a;
      2812: inst = 32'h8220000;
      2813: inst = 32'h10408000;
      2814: inst = 32'hc40450b;
      2815: inst = 32'h8220000;
      2816: inst = 32'h10408000;
      2817: inst = 32'hc40450c;
      2818: inst = 32'h8220000;
      2819: inst = 32'h10408000;
      2820: inst = 32'hc40450d;
      2821: inst = 32'h8220000;
      2822: inst = 32'h10408000;
      2823: inst = 32'hc40450e;
      2824: inst = 32'h8220000;
      2825: inst = 32'h10408000;
      2826: inst = 32'hc40450f;
      2827: inst = 32'h8220000;
      2828: inst = 32'h10408000;
      2829: inst = 32'hc404510;
      2830: inst = 32'h8220000;
      2831: inst = 32'h10408000;
      2832: inst = 32'hc404511;
      2833: inst = 32'h8220000;
      2834: inst = 32'h10408000;
      2835: inst = 32'hc404512;
      2836: inst = 32'h8220000;
      2837: inst = 32'h10408000;
      2838: inst = 32'hc404515;
      2839: inst = 32'h8220000;
      2840: inst = 32'h10408000;
      2841: inst = 32'hc404516;
      2842: inst = 32'h8220000;
      2843: inst = 32'h10408000;
      2844: inst = 32'hc404517;
      2845: inst = 32'h8220000;
      2846: inst = 32'h10408000;
      2847: inst = 32'hc404518;
      2848: inst = 32'h8220000;
      2849: inst = 32'h10408000;
      2850: inst = 32'hc404519;
      2851: inst = 32'h8220000;
      2852: inst = 32'h10408000;
      2853: inst = 32'hc40451a;
      2854: inst = 32'h8220000;
      2855: inst = 32'h10408000;
      2856: inst = 32'hc40451b;
      2857: inst = 32'h8220000;
      2858: inst = 32'h10408000;
      2859: inst = 32'hc40451c;
      2860: inst = 32'h8220000;
      2861: inst = 32'h10408000;
      2862: inst = 32'hc40451d;
      2863: inst = 32'h8220000;
      2864: inst = 32'h10408000;
      2865: inst = 32'hc40451e;
      2866: inst = 32'h8220000;
      2867: inst = 32'h10408000;
      2868: inst = 32'hc40451f;
      2869: inst = 32'h8220000;
      2870: inst = 32'h10408000;
      2871: inst = 32'hc404520;
      2872: inst = 32'h8220000;
      2873: inst = 32'h10408000;
      2874: inst = 32'hc404521;
      2875: inst = 32'h8220000;
      2876: inst = 32'h10408000;
      2877: inst = 32'hc404522;
      2878: inst = 32'h8220000;
      2879: inst = 32'h10408000;
      2880: inst = 32'hc404523;
      2881: inst = 32'h8220000;
      2882: inst = 32'h10408000;
      2883: inst = 32'hc404524;
      2884: inst = 32'h8220000;
      2885: inst = 32'h10408000;
      2886: inst = 32'hc404525;
      2887: inst = 32'h8220000;
      2888: inst = 32'h10408000;
      2889: inst = 32'hc404526;
      2890: inst = 32'h8220000;
      2891: inst = 32'h10408000;
      2892: inst = 32'hc404527;
      2893: inst = 32'h8220000;
      2894: inst = 32'h10408000;
      2895: inst = 32'hc404528;
      2896: inst = 32'h8220000;
      2897: inst = 32'h10408000;
      2898: inst = 32'hc404529;
      2899: inst = 32'h8220000;
      2900: inst = 32'h10408000;
      2901: inst = 32'hc40452a;
      2902: inst = 32'h8220000;
      2903: inst = 32'h10408000;
      2904: inst = 32'hc40452b;
      2905: inst = 32'h8220000;
      2906: inst = 32'h10408000;
      2907: inst = 32'hc40452c;
      2908: inst = 32'h8220000;
      2909: inst = 32'h10408000;
      2910: inst = 32'hc40452d;
      2911: inst = 32'h8220000;
      2912: inst = 32'h10408000;
      2913: inst = 32'hc40452e;
      2914: inst = 32'h8220000;
      2915: inst = 32'h10408000;
      2916: inst = 32'hc40452f;
      2917: inst = 32'h8220000;
      2918: inst = 32'h10408000;
      2919: inst = 32'hc404530;
      2920: inst = 32'h8220000;
      2921: inst = 32'h10408000;
      2922: inst = 32'hc404531;
      2923: inst = 32'h8220000;
      2924: inst = 32'h10408000;
      2925: inst = 32'hc404532;
      2926: inst = 32'h8220000;
      2927: inst = 32'h10408000;
      2928: inst = 32'hc404533;
      2929: inst = 32'h8220000;
      2930: inst = 32'h10408000;
      2931: inst = 32'hc404534;
      2932: inst = 32'h8220000;
      2933: inst = 32'h10408000;
      2934: inst = 32'hc404535;
      2935: inst = 32'h8220000;
      2936: inst = 32'h10408000;
      2937: inst = 32'hc404536;
      2938: inst = 32'h8220000;
      2939: inst = 32'h10408000;
      2940: inst = 32'hc404537;
      2941: inst = 32'h8220000;
      2942: inst = 32'h10408000;
      2943: inst = 32'hc404538;
      2944: inst = 32'h8220000;
      2945: inst = 32'h10408000;
      2946: inst = 32'hc404539;
      2947: inst = 32'h8220000;
      2948: inst = 32'h10408000;
      2949: inst = 32'hc40453a;
      2950: inst = 32'h8220000;
      2951: inst = 32'h10408000;
      2952: inst = 32'hc40453b;
      2953: inst = 32'h8220000;
      2954: inst = 32'h10408000;
      2955: inst = 32'hc404564;
      2956: inst = 32'h8220000;
      2957: inst = 32'h10408000;
      2958: inst = 32'hc404565;
      2959: inst = 32'h8220000;
      2960: inst = 32'h10408000;
      2961: inst = 32'hc404566;
      2962: inst = 32'h8220000;
      2963: inst = 32'h10408000;
      2964: inst = 32'hc404567;
      2965: inst = 32'h8220000;
      2966: inst = 32'h10408000;
      2967: inst = 32'hc404568;
      2968: inst = 32'h8220000;
      2969: inst = 32'h10408000;
      2970: inst = 32'hc404569;
      2971: inst = 32'h8220000;
      2972: inst = 32'h10408000;
      2973: inst = 32'hc40456a;
      2974: inst = 32'h8220000;
      2975: inst = 32'h10408000;
      2976: inst = 32'hc40456b;
      2977: inst = 32'h8220000;
      2978: inst = 32'h10408000;
      2979: inst = 32'hc40456c;
      2980: inst = 32'h8220000;
      2981: inst = 32'h10408000;
      2982: inst = 32'hc40456d;
      2983: inst = 32'h8220000;
      2984: inst = 32'h10408000;
      2985: inst = 32'hc40456e;
      2986: inst = 32'h8220000;
      2987: inst = 32'h10408000;
      2988: inst = 32'hc40456f;
      2989: inst = 32'h8220000;
      2990: inst = 32'h10408000;
      2991: inst = 32'hc404570;
      2992: inst = 32'h8220000;
      2993: inst = 32'h10408000;
      2994: inst = 32'hc404571;
      2995: inst = 32'h8220000;
      2996: inst = 32'h10408000;
      2997: inst = 32'hc404572;
      2998: inst = 32'h8220000;
      2999: inst = 32'h10408000;
      3000: inst = 32'hc404573;
      3001: inst = 32'h8220000;
      3002: inst = 32'h10408000;
      3003: inst = 32'hc404574;
      3004: inst = 32'h8220000;
      3005: inst = 32'h10408000;
      3006: inst = 32'hc404575;
      3007: inst = 32'h8220000;
      3008: inst = 32'h10408000;
      3009: inst = 32'hc404576;
      3010: inst = 32'h8220000;
      3011: inst = 32'h10408000;
      3012: inst = 32'hc404577;
      3013: inst = 32'h8220000;
      3014: inst = 32'h10408000;
      3015: inst = 32'hc404578;
      3016: inst = 32'h8220000;
      3017: inst = 32'h10408000;
      3018: inst = 32'hc404579;
      3019: inst = 32'h8220000;
      3020: inst = 32'h10408000;
      3021: inst = 32'hc40457a;
      3022: inst = 32'h8220000;
      3023: inst = 32'h10408000;
      3024: inst = 32'hc40457b;
      3025: inst = 32'h8220000;
      3026: inst = 32'h10408000;
      3027: inst = 32'hc40457c;
      3028: inst = 32'h8220000;
      3029: inst = 32'h10408000;
      3030: inst = 32'hc40457d;
      3031: inst = 32'h8220000;
      3032: inst = 32'h10408000;
      3033: inst = 32'hc40457e;
      3034: inst = 32'h8220000;
      3035: inst = 32'h10408000;
      3036: inst = 32'hc40457f;
      3037: inst = 32'h8220000;
      3038: inst = 32'h10408000;
      3039: inst = 32'hc404580;
      3040: inst = 32'h8220000;
      3041: inst = 32'h10408000;
      3042: inst = 32'hc404581;
      3043: inst = 32'h8220000;
      3044: inst = 32'h10408000;
      3045: inst = 32'hc404582;
      3046: inst = 32'h8220000;
      3047: inst = 32'h10408000;
      3048: inst = 32'hc404583;
      3049: inst = 32'h8220000;
      3050: inst = 32'h10408000;
      3051: inst = 32'hc404584;
      3052: inst = 32'h8220000;
      3053: inst = 32'h10408000;
      3054: inst = 32'hc404585;
      3055: inst = 32'h8220000;
      3056: inst = 32'h10408000;
      3057: inst = 32'hc404586;
      3058: inst = 32'h8220000;
      3059: inst = 32'h10408000;
      3060: inst = 32'hc404587;
      3061: inst = 32'h8220000;
      3062: inst = 32'h10408000;
      3063: inst = 32'hc404588;
      3064: inst = 32'h8220000;
      3065: inst = 32'h10408000;
      3066: inst = 32'hc404589;
      3067: inst = 32'h8220000;
      3068: inst = 32'h10408000;
      3069: inst = 32'hc40458a;
      3070: inst = 32'h8220000;
      3071: inst = 32'h10408000;
      3072: inst = 32'hc40458b;
      3073: inst = 32'h8220000;
      3074: inst = 32'h10408000;
      3075: inst = 32'hc40458c;
      3076: inst = 32'h8220000;
      3077: inst = 32'h10408000;
      3078: inst = 32'hc40458d;
      3079: inst = 32'h8220000;
      3080: inst = 32'h10408000;
      3081: inst = 32'hc40458e;
      3082: inst = 32'h8220000;
      3083: inst = 32'h10408000;
      3084: inst = 32'hc40458f;
      3085: inst = 32'h8220000;
      3086: inst = 32'h10408000;
      3087: inst = 32'hc404590;
      3088: inst = 32'h8220000;
      3089: inst = 32'h10408000;
      3090: inst = 32'hc404591;
      3091: inst = 32'h8220000;
      3092: inst = 32'h10408000;
      3093: inst = 32'hc404592;
      3094: inst = 32'h8220000;
      3095: inst = 32'h10408000;
      3096: inst = 32'hc404593;
      3097: inst = 32'h8220000;
      3098: inst = 32'h10408000;
      3099: inst = 32'hc404594;
      3100: inst = 32'h8220000;
      3101: inst = 32'h10408000;
      3102: inst = 32'hc404595;
      3103: inst = 32'h8220000;
      3104: inst = 32'h10408000;
      3105: inst = 32'hc404596;
      3106: inst = 32'h8220000;
      3107: inst = 32'h10408000;
      3108: inst = 32'hc404597;
      3109: inst = 32'h8220000;
      3110: inst = 32'h10408000;
      3111: inst = 32'hc404598;
      3112: inst = 32'h8220000;
      3113: inst = 32'h10408000;
      3114: inst = 32'hc404599;
      3115: inst = 32'h8220000;
      3116: inst = 32'h10408000;
      3117: inst = 32'hc40459a;
      3118: inst = 32'h8220000;
      3119: inst = 32'h10408000;
      3120: inst = 32'hc40459b;
      3121: inst = 32'h8220000;
      3122: inst = 32'h10408000;
      3123: inst = 32'hc4045c4;
      3124: inst = 32'h8220000;
      3125: inst = 32'h10408000;
      3126: inst = 32'hc4045c5;
      3127: inst = 32'h8220000;
      3128: inst = 32'h10408000;
      3129: inst = 32'hc4045c6;
      3130: inst = 32'h8220000;
      3131: inst = 32'h10408000;
      3132: inst = 32'hc4045c7;
      3133: inst = 32'h8220000;
      3134: inst = 32'h10408000;
      3135: inst = 32'hc4045c8;
      3136: inst = 32'h8220000;
      3137: inst = 32'h10408000;
      3138: inst = 32'hc4045c9;
      3139: inst = 32'h8220000;
      3140: inst = 32'h10408000;
      3141: inst = 32'hc4045ca;
      3142: inst = 32'h8220000;
      3143: inst = 32'h10408000;
      3144: inst = 32'hc4045cb;
      3145: inst = 32'h8220000;
      3146: inst = 32'h10408000;
      3147: inst = 32'hc4045cc;
      3148: inst = 32'h8220000;
      3149: inst = 32'h10408000;
      3150: inst = 32'hc4045cd;
      3151: inst = 32'h8220000;
      3152: inst = 32'h10408000;
      3153: inst = 32'hc4045ce;
      3154: inst = 32'h8220000;
      3155: inst = 32'h10408000;
      3156: inst = 32'hc4045cf;
      3157: inst = 32'h8220000;
      3158: inst = 32'h10408000;
      3159: inst = 32'hc4045d0;
      3160: inst = 32'h8220000;
      3161: inst = 32'h10408000;
      3162: inst = 32'hc4045d1;
      3163: inst = 32'h8220000;
      3164: inst = 32'h10408000;
      3165: inst = 32'hc4045d2;
      3166: inst = 32'h8220000;
      3167: inst = 32'h10408000;
      3168: inst = 32'hc4045d3;
      3169: inst = 32'h8220000;
      3170: inst = 32'h10408000;
      3171: inst = 32'hc4045d4;
      3172: inst = 32'h8220000;
      3173: inst = 32'h10408000;
      3174: inst = 32'hc4045d5;
      3175: inst = 32'h8220000;
      3176: inst = 32'h10408000;
      3177: inst = 32'hc4045d6;
      3178: inst = 32'h8220000;
      3179: inst = 32'h10408000;
      3180: inst = 32'hc4045d7;
      3181: inst = 32'h8220000;
      3182: inst = 32'h10408000;
      3183: inst = 32'hc4045d8;
      3184: inst = 32'h8220000;
      3185: inst = 32'h10408000;
      3186: inst = 32'hc4045d9;
      3187: inst = 32'h8220000;
      3188: inst = 32'h10408000;
      3189: inst = 32'hc4045da;
      3190: inst = 32'h8220000;
      3191: inst = 32'h10408000;
      3192: inst = 32'hc4045db;
      3193: inst = 32'h8220000;
      3194: inst = 32'h10408000;
      3195: inst = 32'hc4045dc;
      3196: inst = 32'h8220000;
      3197: inst = 32'h10408000;
      3198: inst = 32'hc4045dd;
      3199: inst = 32'h8220000;
      3200: inst = 32'h10408000;
      3201: inst = 32'hc4045de;
      3202: inst = 32'h8220000;
      3203: inst = 32'h10408000;
      3204: inst = 32'hc4045df;
      3205: inst = 32'h8220000;
      3206: inst = 32'h10408000;
      3207: inst = 32'hc4045e0;
      3208: inst = 32'h8220000;
      3209: inst = 32'h10408000;
      3210: inst = 32'hc4045e1;
      3211: inst = 32'h8220000;
      3212: inst = 32'h10408000;
      3213: inst = 32'hc4045e2;
      3214: inst = 32'h8220000;
      3215: inst = 32'h10408000;
      3216: inst = 32'hc4045e3;
      3217: inst = 32'h8220000;
      3218: inst = 32'h10408000;
      3219: inst = 32'hc4045e4;
      3220: inst = 32'h8220000;
      3221: inst = 32'h10408000;
      3222: inst = 32'hc4045e5;
      3223: inst = 32'h8220000;
      3224: inst = 32'h10408000;
      3225: inst = 32'hc4045e6;
      3226: inst = 32'h8220000;
      3227: inst = 32'h10408000;
      3228: inst = 32'hc4045e7;
      3229: inst = 32'h8220000;
      3230: inst = 32'h10408000;
      3231: inst = 32'hc4045e8;
      3232: inst = 32'h8220000;
      3233: inst = 32'h10408000;
      3234: inst = 32'hc4045e9;
      3235: inst = 32'h8220000;
      3236: inst = 32'h10408000;
      3237: inst = 32'hc4045ea;
      3238: inst = 32'h8220000;
      3239: inst = 32'h10408000;
      3240: inst = 32'hc4045eb;
      3241: inst = 32'h8220000;
      3242: inst = 32'h10408000;
      3243: inst = 32'hc4045ec;
      3244: inst = 32'h8220000;
      3245: inst = 32'h10408000;
      3246: inst = 32'hc4045ed;
      3247: inst = 32'h8220000;
      3248: inst = 32'h10408000;
      3249: inst = 32'hc4045ee;
      3250: inst = 32'h8220000;
      3251: inst = 32'h10408000;
      3252: inst = 32'hc4045ef;
      3253: inst = 32'h8220000;
      3254: inst = 32'h10408000;
      3255: inst = 32'hc4045f0;
      3256: inst = 32'h8220000;
      3257: inst = 32'h10408000;
      3258: inst = 32'hc4045f1;
      3259: inst = 32'h8220000;
      3260: inst = 32'h10408000;
      3261: inst = 32'hc4045f2;
      3262: inst = 32'h8220000;
      3263: inst = 32'h10408000;
      3264: inst = 32'hc4045f3;
      3265: inst = 32'h8220000;
      3266: inst = 32'h10408000;
      3267: inst = 32'hc4045f4;
      3268: inst = 32'h8220000;
      3269: inst = 32'h10408000;
      3270: inst = 32'hc4045f5;
      3271: inst = 32'h8220000;
      3272: inst = 32'h10408000;
      3273: inst = 32'hc4045f6;
      3274: inst = 32'h8220000;
      3275: inst = 32'h10408000;
      3276: inst = 32'hc4045f7;
      3277: inst = 32'h8220000;
      3278: inst = 32'h10408000;
      3279: inst = 32'hc4045f8;
      3280: inst = 32'h8220000;
      3281: inst = 32'h10408000;
      3282: inst = 32'hc4045f9;
      3283: inst = 32'h8220000;
      3284: inst = 32'h10408000;
      3285: inst = 32'hc4045fa;
      3286: inst = 32'h8220000;
      3287: inst = 32'h10408000;
      3288: inst = 32'hc4045fb;
      3289: inst = 32'h8220000;
      3290: inst = 32'h10408000;
      3291: inst = 32'hc404624;
      3292: inst = 32'h8220000;
      3293: inst = 32'h10408000;
      3294: inst = 32'hc404625;
      3295: inst = 32'h8220000;
      3296: inst = 32'h10408000;
      3297: inst = 32'hc404626;
      3298: inst = 32'h8220000;
      3299: inst = 32'h10408000;
      3300: inst = 32'hc404627;
      3301: inst = 32'h8220000;
      3302: inst = 32'h10408000;
      3303: inst = 32'hc404628;
      3304: inst = 32'h8220000;
      3305: inst = 32'h10408000;
      3306: inst = 32'hc404629;
      3307: inst = 32'h8220000;
      3308: inst = 32'h10408000;
      3309: inst = 32'hc40462a;
      3310: inst = 32'h8220000;
      3311: inst = 32'h10408000;
      3312: inst = 32'hc40462b;
      3313: inst = 32'h8220000;
      3314: inst = 32'h10408000;
      3315: inst = 32'hc40462c;
      3316: inst = 32'h8220000;
      3317: inst = 32'h10408000;
      3318: inst = 32'hc40462d;
      3319: inst = 32'h8220000;
      3320: inst = 32'h10408000;
      3321: inst = 32'hc40462e;
      3322: inst = 32'h8220000;
      3323: inst = 32'h10408000;
      3324: inst = 32'hc40462f;
      3325: inst = 32'h8220000;
      3326: inst = 32'h10408000;
      3327: inst = 32'hc404630;
      3328: inst = 32'h8220000;
      3329: inst = 32'h10408000;
      3330: inst = 32'hc404631;
      3331: inst = 32'h8220000;
      3332: inst = 32'h10408000;
      3333: inst = 32'hc404632;
      3334: inst = 32'h8220000;
      3335: inst = 32'h10408000;
      3336: inst = 32'hc404633;
      3337: inst = 32'h8220000;
      3338: inst = 32'h10408000;
      3339: inst = 32'hc404634;
      3340: inst = 32'h8220000;
      3341: inst = 32'h10408000;
      3342: inst = 32'hc404635;
      3343: inst = 32'h8220000;
      3344: inst = 32'h10408000;
      3345: inst = 32'hc404636;
      3346: inst = 32'h8220000;
      3347: inst = 32'h10408000;
      3348: inst = 32'hc404637;
      3349: inst = 32'h8220000;
      3350: inst = 32'h10408000;
      3351: inst = 32'hc404638;
      3352: inst = 32'h8220000;
      3353: inst = 32'h10408000;
      3354: inst = 32'hc404639;
      3355: inst = 32'h8220000;
      3356: inst = 32'h10408000;
      3357: inst = 32'hc40463a;
      3358: inst = 32'h8220000;
      3359: inst = 32'h10408000;
      3360: inst = 32'hc40463b;
      3361: inst = 32'h8220000;
      3362: inst = 32'h10408000;
      3363: inst = 32'hc40463c;
      3364: inst = 32'h8220000;
      3365: inst = 32'h10408000;
      3366: inst = 32'hc40463d;
      3367: inst = 32'h8220000;
      3368: inst = 32'h10408000;
      3369: inst = 32'hc40463e;
      3370: inst = 32'h8220000;
      3371: inst = 32'h10408000;
      3372: inst = 32'hc40463f;
      3373: inst = 32'h8220000;
      3374: inst = 32'h10408000;
      3375: inst = 32'hc404640;
      3376: inst = 32'h8220000;
      3377: inst = 32'h10408000;
      3378: inst = 32'hc404641;
      3379: inst = 32'h8220000;
      3380: inst = 32'h10408000;
      3381: inst = 32'hc404642;
      3382: inst = 32'h8220000;
      3383: inst = 32'h10408000;
      3384: inst = 32'hc404643;
      3385: inst = 32'h8220000;
      3386: inst = 32'h10408000;
      3387: inst = 32'hc404644;
      3388: inst = 32'h8220000;
      3389: inst = 32'h10408000;
      3390: inst = 32'hc404645;
      3391: inst = 32'h8220000;
      3392: inst = 32'h10408000;
      3393: inst = 32'hc404646;
      3394: inst = 32'h8220000;
      3395: inst = 32'h10408000;
      3396: inst = 32'hc404647;
      3397: inst = 32'h8220000;
      3398: inst = 32'h10408000;
      3399: inst = 32'hc404648;
      3400: inst = 32'h8220000;
      3401: inst = 32'h10408000;
      3402: inst = 32'hc404649;
      3403: inst = 32'h8220000;
      3404: inst = 32'h10408000;
      3405: inst = 32'hc40464a;
      3406: inst = 32'h8220000;
      3407: inst = 32'h10408000;
      3408: inst = 32'hc40464b;
      3409: inst = 32'h8220000;
      3410: inst = 32'h10408000;
      3411: inst = 32'hc40464c;
      3412: inst = 32'h8220000;
      3413: inst = 32'h10408000;
      3414: inst = 32'hc40464d;
      3415: inst = 32'h8220000;
      3416: inst = 32'h10408000;
      3417: inst = 32'hc40464e;
      3418: inst = 32'h8220000;
      3419: inst = 32'h10408000;
      3420: inst = 32'hc40464f;
      3421: inst = 32'h8220000;
      3422: inst = 32'h10408000;
      3423: inst = 32'hc404650;
      3424: inst = 32'h8220000;
      3425: inst = 32'h10408000;
      3426: inst = 32'hc404651;
      3427: inst = 32'h8220000;
      3428: inst = 32'h10408000;
      3429: inst = 32'hc404652;
      3430: inst = 32'h8220000;
      3431: inst = 32'h10408000;
      3432: inst = 32'hc404653;
      3433: inst = 32'h8220000;
      3434: inst = 32'h10408000;
      3435: inst = 32'hc404654;
      3436: inst = 32'h8220000;
      3437: inst = 32'h10408000;
      3438: inst = 32'hc404655;
      3439: inst = 32'h8220000;
      3440: inst = 32'h10408000;
      3441: inst = 32'hc404656;
      3442: inst = 32'h8220000;
      3443: inst = 32'h10408000;
      3444: inst = 32'hc404657;
      3445: inst = 32'h8220000;
      3446: inst = 32'h10408000;
      3447: inst = 32'hc404658;
      3448: inst = 32'h8220000;
      3449: inst = 32'h10408000;
      3450: inst = 32'hc404659;
      3451: inst = 32'h8220000;
      3452: inst = 32'h10408000;
      3453: inst = 32'hc40465a;
      3454: inst = 32'h8220000;
      3455: inst = 32'h10408000;
      3456: inst = 32'hc40465b;
      3457: inst = 32'h8220000;
      3458: inst = 32'h10408000;
      3459: inst = 32'hc404684;
      3460: inst = 32'h8220000;
      3461: inst = 32'h10408000;
      3462: inst = 32'hc404685;
      3463: inst = 32'h8220000;
      3464: inst = 32'h10408000;
      3465: inst = 32'hc404686;
      3466: inst = 32'h8220000;
      3467: inst = 32'h10408000;
      3468: inst = 32'hc404687;
      3469: inst = 32'h8220000;
      3470: inst = 32'h10408000;
      3471: inst = 32'hc404688;
      3472: inst = 32'h8220000;
      3473: inst = 32'h10408000;
      3474: inst = 32'hc404689;
      3475: inst = 32'h8220000;
      3476: inst = 32'h10408000;
      3477: inst = 32'hc40468a;
      3478: inst = 32'h8220000;
      3479: inst = 32'h10408000;
      3480: inst = 32'hc40468b;
      3481: inst = 32'h8220000;
      3482: inst = 32'h10408000;
      3483: inst = 32'hc40468c;
      3484: inst = 32'h8220000;
      3485: inst = 32'h10408000;
      3486: inst = 32'hc40468d;
      3487: inst = 32'h8220000;
      3488: inst = 32'h10408000;
      3489: inst = 32'hc40468e;
      3490: inst = 32'h8220000;
      3491: inst = 32'h10408000;
      3492: inst = 32'hc40468f;
      3493: inst = 32'h8220000;
      3494: inst = 32'h10408000;
      3495: inst = 32'hc404690;
      3496: inst = 32'h8220000;
      3497: inst = 32'h10408000;
      3498: inst = 32'hc404691;
      3499: inst = 32'h8220000;
      3500: inst = 32'h10408000;
      3501: inst = 32'hc404692;
      3502: inst = 32'h8220000;
      3503: inst = 32'h10408000;
      3504: inst = 32'hc404693;
      3505: inst = 32'h8220000;
      3506: inst = 32'h10408000;
      3507: inst = 32'hc404694;
      3508: inst = 32'h8220000;
      3509: inst = 32'h10408000;
      3510: inst = 32'hc404695;
      3511: inst = 32'h8220000;
      3512: inst = 32'h10408000;
      3513: inst = 32'hc404696;
      3514: inst = 32'h8220000;
      3515: inst = 32'h10408000;
      3516: inst = 32'hc404697;
      3517: inst = 32'h8220000;
      3518: inst = 32'h10408000;
      3519: inst = 32'hc404698;
      3520: inst = 32'h8220000;
      3521: inst = 32'h10408000;
      3522: inst = 32'hc404699;
      3523: inst = 32'h8220000;
      3524: inst = 32'h10408000;
      3525: inst = 32'hc40469a;
      3526: inst = 32'h8220000;
      3527: inst = 32'h10408000;
      3528: inst = 32'hc40469b;
      3529: inst = 32'h8220000;
      3530: inst = 32'h10408000;
      3531: inst = 32'hc40469c;
      3532: inst = 32'h8220000;
      3533: inst = 32'h10408000;
      3534: inst = 32'hc40469d;
      3535: inst = 32'h8220000;
      3536: inst = 32'h10408000;
      3537: inst = 32'hc40469e;
      3538: inst = 32'h8220000;
      3539: inst = 32'h10408000;
      3540: inst = 32'hc40469f;
      3541: inst = 32'h8220000;
      3542: inst = 32'h10408000;
      3543: inst = 32'hc4046a0;
      3544: inst = 32'h8220000;
      3545: inst = 32'h10408000;
      3546: inst = 32'hc4046a1;
      3547: inst = 32'h8220000;
      3548: inst = 32'h10408000;
      3549: inst = 32'hc4046a2;
      3550: inst = 32'h8220000;
      3551: inst = 32'h10408000;
      3552: inst = 32'hc4046a3;
      3553: inst = 32'h8220000;
      3554: inst = 32'h10408000;
      3555: inst = 32'hc4046a4;
      3556: inst = 32'h8220000;
      3557: inst = 32'h10408000;
      3558: inst = 32'hc4046a5;
      3559: inst = 32'h8220000;
      3560: inst = 32'h10408000;
      3561: inst = 32'hc4046a6;
      3562: inst = 32'h8220000;
      3563: inst = 32'h10408000;
      3564: inst = 32'hc4046a7;
      3565: inst = 32'h8220000;
      3566: inst = 32'h10408000;
      3567: inst = 32'hc4046a8;
      3568: inst = 32'h8220000;
      3569: inst = 32'h10408000;
      3570: inst = 32'hc4046a9;
      3571: inst = 32'h8220000;
      3572: inst = 32'h10408000;
      3573: inst = 32'hc4046aa;
      3574: inst = 32'h8220000;
      3575: inst = 32'h10408000;
      3576: inst = 32'hc4046ab;
      3577: inst = 32'h8220000;
      3578: inst = 32'h10408000;
      3579: inst = 32'hc4046ac;
      3580: inst = 32'h8220000;
      3581: inst = 32'h10408000;
      3582: inst = 32'hc4046ad;
      3583: inst = 32'h8220000;
      3584: inst = 32'h10408000;
      3585: inst = 32'hc4046ae;
      3586: inst = 32'h8220000;
      3587: inst = 32'h10408000;
      3588: inst = 32'hc4046af;
      3589: inst = 32'h8220000;
      3590: inst = 32'h10408000;
      3591: inst = 32'hc4046b0;
      3592: inst = 32'h8220000;
      3593: inst = 32'h10408000;
      3594: inst = 32'hc4046b1;
      3595: inst = 32'h8220000;
      3596: inst = 32'h10408000;
      3597: inst = 32'hc4046b2;
      3598: inst = 32'h8220000;
      3599: inst = 32'h10408000;
      3600: inst = 32'hc4046b3;
      3601: inst = 32'h8220000;
      3602: inst = 32'h10408000;
      3603: inst = 32'hc4046b4;
      3604: inst = 32'h8220000;
      3605: inst = 32'h10408000;
      3606: inst = 32'hc4046b5;
      3607: inst = 32'h8220000;
      3608: inst = 32'h10408000;
      3609: inst = 32'hc4046b6;
      3610: inst = 32'h8220000;
      3611: inst = 32'h10408000;
      3612: inst = 32'hc4046b7;
      3613: inst = 32'h8220000;
      3614: inst = 32'h10408000;
      3615: inst = 32'hc4046b8;
      3616: inst = 32'h8220000;
      3617: inst = 32'h10408000;
      3618: inst = 32'hc4046b9;
      3619: inst = 32'h8220000;
      3620: inst = 32'h10408000;
      3621: inst = 32'hc4046ba;
      3622: inst = 32'h8220000;
      3623: inst = 32'h10408000;
      3624: inst = 32'hc4046bb;
      3625: inst = 32'h8220000;
      3626: inst = 32'h10408000;
      3627: inst = 32'hc4046e4;
      3628: inst = 32'h8220000;
      3629: inst = 32'h10408000;
      3630: inst = 32'hc4046e5;
      3631: inst = 32'h8220000;
      3632: inst = 32'h10408000;
      3633: inst = 32'hc4046e6;
      3634: inst = 32'h8220000;
      3635: inst = 32'h10408000;
      3636: inst = 32'hc4046e7;
      3637: inst = 32'h8220000;
      3638: inst = 32'h10408000;
      3639: inst = 32'hc4046e8;
      3640: inst = 32'h8220000;
      3641: inst = 32'h10408000;
      3642: inst = 32'hc4046e9;
      3643: inst = 32'h8220000;
      3644: inst = 32'h10408000;
      3645: inst = 32'hc4046ea;
      3646: inst = 32'h8220000;
      3647: inst = 32'h10408000;
      3648: inst = 32'hc4046eb;
      3649: inst = 32'h8220000;
      3650: inst = 32'h10408000;
      3651: inst = 32'hc4046ec;
      3652: inst = 32'h8220000;
      3653: inst = 32'h10408000;
      3654: inst = 32'hc4046ed;
      3655: inst = 32'h8220000;
      3656: inst = 32'h10408000;
      3657: inst = 32'hc4046ee;
      3658: inst = 32'h8220000;
      3659: inst = 32'h10408000;
      3660: inst = 32'hc404700;
      3661: inst = 32'h8220000;
      3662: inst = 32'h10408000;
      3663: inst = 32'hc404701;
      3664: inst = 32'h8220000;
      3665: inst = 32'h10408000;
      3666: inst = 32'hc404702;
      3667: inst = 32'h8220000;
      3668: inst = 32'h10408000;
      3669: inst = 32'hc404703;
      3670: inst = 32'h8220000;
      3671: inst = 32'h10408000;
      3672: inst = 32'hc404704;
      3673: inst = 32'h8220000;
      3674: inst = 32'h10408000;
      3675: inst = 32'hc404705;
      3676: inst = 32'h8220000;
      3677: inst = 32'h10408000;
      3678: inst = 32'hc404706;
      3679: inst = 32'h8220000;
      3680: inst = 32'h10408000;
      3681: inst = 32'hc404707;
      3682: inst = 32'h8220000;
      3683: inst = 32'h10408000;
      3684: inst = 32'hc404708;
      3685: inst = 32'h8220000;
      3686: inst = 32'h10408000;
      3687: inst = 32'hc404709;
      3688: inst = 32'h8220000;
      3689: inst = 32'h10408000;
      3690: inst = 32'hc40470a;
      3691: inst = 32'h8220000;
      3692: inst = 32'h10408000;
      3693: inst = 32'hc40470b;
      3694: inst = 32'h8220000;
      3695: inst = 32'h10408000;
      3696: inst = 32'hc40470c;
      3697: inst = 32'h8220000;
      3698: inst = 32'h10408000;
      3699: inst = 32'hc40470d;
      3700: inst = 32'h8220000;
      3701: inst = 32'h10408000;
      3702: inst = 32'hc40470e;
      3703: inst = 32'h8220000;
      3704: inst = 32'h10408000;
      3705: inst = 32'hc40470f;
      3706: inst = 32'h8220000;
      3707: inst = 32'h10408000;
      3708: inst = 32'hc404710;
      3709: inst = 32'h8220000;
      3710: inst = 32'h10408000;
      3711: inst = 32'hc404711;
      3712: inst = 32'h8220000;
      3713: inst = 32'h10408000;
      3714: inst = 32'hc404712;
      3715: inst = 32'h8220000;
      3716: inst = 32'h10408000;
      3717: inst = 32'hc404713;
      3718: inst = 32'h8220000;
      3719: inst = 32'h10408000;
      3720: inst = 32'hc404714;
      3721: inst = 32'h8220000;
      3722: inst = 32'h10408000;
      3723: inst = 32'hc404715;
      3724: inst = 32'h8220000;
      3725: inst = 32'h10408000;
      3726: inst = 32'hc404716;
      3727: inst = 32'h8220000;
      3728: inst = 32'h10408000;
      3729: inst = 32'hc404717;
      3730: inst = 32'h8220000;
      3731: inst = 32'h10408000;
      3732: inst = 32'hc404718;
      3733: inst = 32'h8220000;
      3734: inst = 32'h10408000;
      3735: inst = 32'hc404719;
      3736: inst = 32'h8220000;
      3737: inst = 32'h10408000;
      3738: inst = 32'hc40471a;
      3739: inst = 32'h8220000;
      3740: inst = 32'h10408000;
      3741: inst = 32'hc40471b;
      3742: inst = 32'h8220000;
      3743: inst = 32'h10408000;
      3744: inst = 32'hc404744;
      3745: inst = 32'h8220000;
      3746: inst = 32'h10408000;
      3747: inst = 32'hc404745;
      3748: inst = 32'h8220000;
      3749: inst = 32'h10408000;
      3750: inst = 32'hc404746;
      3751: inst = 32'h8220000;
      3752: inst = 32'h10408000;
      3753: inst = 32'hc404747;
      3754: inst = 32'h8220000;
      3755: inst = 32'h10408000;
      3756: inst = 32'hc404748;
      3757: inst = 32'h8220000;
      3758: inst = 32'h10408000;
      3759: inst = 32'hc404749;
      3760: inst = 32'h8220000;
      3761: inst = 32'h10408000;
      3762: inst = 32'hc40474a;
      3763: inst = 32'h8220000;
      3764: inst = 32'h10408000;
      3765: inst = 32'hc40474b;
      3766: inst = 32'h8220000;
      3767: inst = 32'h10408000;
      3768: inst = 32'hc40474c;
      3769: inst = 32'h8220000;
      3770: inst = 32'h10408000;
      3771: inst = 32'hc40474d;
      3772: inst = 32'h8220000;
      3773: inst = 32'h10408000;
      3774: inst = 32'hc40474e;
      3775: inst = 32'h8220000;
      3776: inst = 32'h10408000;
      3777: inst = 32'hc404760;
      3778: inst = 32'h8220000;
      3779: inst = 32'h10408000;
      3780: inst = 32'hc404761;
      3781: inst = 32'h8220000;
      3782: inst = 32'h10408000;
      3783: inst = 32'hc404762;
      3784: inst = 32'h8220000;
      3785: inst = 32'h10408000;
      3786: inst = 32'hc404763;
      3787: inst = 32'h8220000;
      3788: inst = 32'h10408000;
      3789: inst = 32'hc404764;
      3790: inst = 32'h8220000;
      3791: inst = 32'h10408000;
      3792: inst = 32'hc404765;
      3793: inst = 32'h8220000;
      3794: inst = 32'h10408000;
      3795: inst = 32'hc404766;
      3796: inst = 32'h8220000;
      3797: inst = 32'h10408000;
      3798: inst = 32'hc404767;
      3799: inst = 32'h8220000;
      3800: inst = 32'h10408000;
      3801: inst = 32'hc404768;
      3802: inst = 32'h8220000;
      3803: inst = 32'h10408000;
      3804: inst = 32'hc404769;
      3805: inst = 32'h8220000;
      3806: inst = 32'h10408000;
      3807: inst = 32'hc40476a;
      3808: inst = 32'h8220000;
      3809: inst = 32'h10408000;
      3810: inst = 32'hc40476b;
      3811: inst = 32'h8220000;
      3812: inst = 32'h10408000;
      3813: inst = 32'hc40476c;
      3814: inst = 32'h8220000;
      3815: inst = 32'h10408000;
      3816: inst = 32'hc40476d;
      3817: inst = 32'h8220000;
      3818: inst = 32'h10408000;
      3819: inst = 32'hc40476e;
      3820: inst = 32'h8220000;
      3821: inst = 32'h10408000;
      3822: inst = 32'hc40476f;
      3823: inst = 32'h8220000;
      3824: inst = 32'h10408000;
      3825: inst = 32'hc404770;
      3826: inst = 32'h8220000;
      3827: inst = 32'h10408000;
      3828: inst = 32'hc404771;
      3829: inst = 32'h8220000;
      3830: inst = 32'h10408000;
      3831: inst = 32'hc404772;
      3832: inst = 32'h8220000;
      3833: inst = 32'h10408000;
      3834: inst = 32'hc404773;
      3835: inst = 32'h8220000;
      3836: inst = 32'h10408000;
      3837: inst = 32'hc404774;
      3838: inst = 32'h8220000;
      3839: inst = 32'h10408000;
      3840: inst = 32'hc404775;
      3841: inst = 32'h8220000;
      3842: inst = 32'h10408000;
      3843: inst = 32'hc404776;
      3844: inst = 32'h8220000;
      3845: inst = 32'h10408000;
      3846: inst = 32'hc404777;
      3847: inst = 32'h8220000;
      3848: inst = 32'h10408000;
      3849: inst = 32'hc404778;
      3850: inst = 32'h8220000;
      3851: inst = 32'h10408000;
      3852: inst = 32'hc404779;
      3853: inst = 32'h8220000;
      3854: inst = 32'h10408000;
      3855: inst = 32'hc40477a;
      3856: inst = 32'h8220000;
      3857: inst = 32'h10408000;
      3858: inst = 32'hc40477b;
      3859: inst = 32'h8220000;
      3860: inst = 32'h10408000;
      3861: inst = 32'hc4047a4;
      3862: inst = 32'h8220000;
      3863: inst = 32'h10408000;
      3864: inst = 32'hc4047a5;
      3865: inst = 32'h8220000;
      3866: inst = 32'h10408000;
      3867: inst = 32'hc4047a6;
      3868: inst = 32'h8220000;
      3869: inst = 32'h10408000;
      3870: inst = 32'hc4047a7;
      3871: inst = 32'h8220000;
      3872: inst = 32'h10408000;
      3873: inst = 32'hc4047a8;
      3874: inst = 32'h8220000;
      3875: inst = 32'h10408000;
      3876: inst = 32'hc4047a9;
      3877: inst = 32'h8220000;
      3878: inst = 32'h10408000;
      3879: inst = 32'hc4047aa;
      3880: inst = 32'h8220000;
      3881: inst = 32'h10408000;
      3882: inst = 32'hc4047ab;
      3883: inst = 32'h8220000;
      3884: inst = 32'h10408000;
      3885: inst = 32'hc4047ac;
      3886: inst = 32'h8220000;
      3887: inst = 32'h10408000;
      3888: inst = 32'hc4047ad;
      3889: inst = 32'h8220000;
      3890: inst = 32'h10408000;
      3891: inst = 32'hc4047ae;
      3892: inst = 32'h8220000;
      3893: inst = 32'h10408000;
      3894: inst = 32'hc4047c0;
      3895: inst = 32'h8220000;
      3896: inst = 32'h10408000;
      3897: inst = 32'hc4047c1;
      3898: inst = 32'h8220000;
      3899: inst = 32'h10408000;
      3900: inst = 32'hc4047c2;
      3901: inst = 32'h8220000;
      3902: inst = 32'h10408000;
      3903: inst = 32'hc4047c3;
      3904: inst = 32'h8220000;
      3905: inst = 32'h10408000;
      3906: inst = 32'hc4047c4;
      3907: inst = 32'h8220000;
      3908: inst = 32'h10408000;
      3909: inst = 32'hc4047c5;
      3910: inst = 32'h8220000;
      3911: inst = 32'h10408000;
      3912: inst = 32'hc4047c6;
      3913: inst = 32'h8220000;
      3914: inst = 32'h10408000;
      3915: inst = 32'hc4047c7;
      3916: inst = 32'h8220000;
      3917: inst = 32'h10408000;
      3918: inst = 32'hc4047c8;
      3919: inst = 32'h8220000;
      3920: inst = 32'h10408000;
      3921: inst = 32'hc4047c9;
      3922: inst = 32'h8220000;
      3923: inst = 32'h10408000;
      3924: inst = 32'hc4047ca;
      3925: inst = 32'h8220000;
      3926: inst = 32'h10408000;
      3927: inst = 32'hc4047cb;
      3928: inst = 32'h8220000;
      3929: inst = 32'h10408000;
      3930: inst = 32'hc4047cc;
      3931: inst = 32'h8220000;
      3932: inst = 32'h10408000;
      3933: inst = 32'hc4047cd;
      3934: inst = 32'h8220000;
      3935: inst = 32'h10408000;
      3936: inst = 32'hc4047ce;
      3937: inst = 32'h8220000;
      3938: inst = 32'h10408000;
      3939: inst = 32'hc4047cf;
      3940: inst = 32'h8220000;
      3941: inst = 32'h10408000;
      3942: inst = 32'hc4047d0;
      3943: inst = 32'h8220000;
      3944: inst = 32'h10408000;
      3945: inst = 32'hc4047d1;
      3946: inst = 32'h8220000;
      3947: inst = 32'h10408000;
      3948: inst = 32'hc4047d2;
      3949: inst = 32'h8220000;
      3950: inst = 32'h10408000;
      3951: inst = 32'hc4047d3;
      3952: inst = 32'h8220000;
      3953: inst = 32'h10408000;
      3954: inst = 32'hc4047d4;
      3955: inst = 32'h8220000;
      3956: inst = 32'h10408000;
      3957: inst = 32'hc4047d5;
      3958: inst = 32'h8220000;
      3959: inst = 32'h10408000;
      3960: inst = 32'hc4047d6;
      3961: inst = 32'h8220000;
      3962: inst = 32'h10408000;
      3963: inst = 32'hc4047d7;
      3964: inst = 32'h8220000;
      3965: inst = 32'h10408000;
      3966: inst = 32'hc4047d8;
      3967: inst = 32'h8220000;
      3968: inst = 32'h10408000;
      3969: inst = 32'hc4047d9;
      3970: inst = 32'h8220000;
      3971: inst = 32'h10408000;
      3972: inst = 32'hc4047da;
      3973: inst = 32'h8220000;
      3974: inst = 32'h10408000;
      3975: inst = 32'hc4047db;
      3976: inst = 32'h8220000;
      3977: inst = 32'h10408000;
      3978: inst = 32'hc404804;
      3979: inst = 32'h8220000;
      3980: inst = 32'h10408000;
      3981: inst = 32'hc404805;
      3982: inst = 32'h8220000;
      3983: inst = 32'h10408000;
      3984: inst = 32'hc404806;
      3985: inst = 32'h8220000;
      3986: inst = 32'h10408000;
      3987: inst = 32'hc404807;
      3988: inst = 32'h8220000;
      3989: inst = 32'h10408000;
      3990: inst = 32'hc404808;
      3991: inst = 32'h8220000;
      3992: inst = 32'h10408000;
      3993: inst = 32'hc404809;
      3994: inst = 32'h8220000;
      3995: inst = 32'h10408000;
      3996: inst = 32'hc40480a;
      3997: inst = 32'h8220000;
      3998: inst = 32'h10408000;
      3999: inst = 32'hc40480b;
      4000: inst = 32'h8220000;
      4001: inst = 32'h10408000;
      4002: inst = 32'hc40480c;
      4003: inst = 32'h8220000;
      4004: inst = 32'h10408000;
      4005: inst = 32'hc40480d;
      4006: inst = 32'h8220000;
      4007: inst = 32'h10408000;
      4008: inst = 32'hc40480e;
      4009: inst = 32'h8220000;
      4010: inst = 32'h10408000;
      4011: inst = 32'hc404820;
      4012: inst = 32'h8220000;
      4013: inst = 32'h10408000;
      4014: inst = 32'hc404821;
      4015: inst = 32'h8220000;
      4016: inst = 32'h10408000;
      4017: inst = 32'hc404822;
      4018: inst = 32'h8220000;
      4019: inst = 32'h10408000;
      4020: inst = 32'hc404823;
      4021: inst = 32'h8220000;
      4022: inst = 32'h10408000;
      4023: inst = 32'hc404824;
      4024: inst = 32'h8220000;
      4025: inst = 32'h10408000;
      4026: inst = 32'hc404825;
      4027: inst = 32'h8220000;
      4028: inst = 32'h10408000;
      4029: inst = 32'hc404826;
      4030: inst = 32'h8220000;
      4031: inst = 32'h10408000;
      4032: inst = 32'hc404827;
      4033: inst = 32'h8220000;
      4034: inst = 32'h10408000;
      4035: inst = 32'hc404828;
      4036: inst = 32'h8220000;
      4037: inst = 32'h10408000;
      4038: inst = 32'hc404829;
      4039: inst = 32'h8220000;
      4040: inst = 32'h10408000;
      4041: inst = 32'hc40482a;
      4042: inst = 32'h8220000;
      4043: inst = 32'h10408000;
      4044: inst = 32'hc40482b;
      4045: inst = 32'h8220000;
      4046: inst = 32'h10408000;
      4047: inst = 32'hc40482c;
      4048: inst = 32'h8220000;
      4049: inst = 32'h10408000;
      4050: inst = 32'hc40482d;
      4051: inst = 32'h8220000;
      4052: inst = 32'h10408000;
      4053: inst = 32'hc40482e;
      4054: inst = 32'h8220000;
      4055: inst = 32'h10408000;
      4056: inst = 32'hc40482f;
      4057: inst = 32'h8220000;
      4058: inst = 32'h10408000;
      4059: inst = 32'hc404830;
      4060: inst = 32'h8220000;
      4061: inst = 32'h10408000;
      4062: inst = 32'hc404831;
      4063: inst = 32'h8220000;
      4064: inst = 32'h10408000;
      4065: inst = 32'hc404832;
      4066: inst = 32'h8220000;
      4067: inst = 32'h10408000;
      4068: inst = 32'hc404833;
      4069: inst = 32'h8220000;
      4070: inst = 32'h10408000;
      4071: inst = 32'hc404834;
      4072: inst = 32'h8220000;
      4073: inst = 32'h10408000;
      4074: inst = 32'hc404835;
      4075: inst = 32'h8220000;
      4076: inst = 32'h10408000;
      4077: inst = 32'hc404836;
      4078: inst = 32'h8220000;
      4079: inst = 32'h10408000;
      4080: inst = 32'hc404837;
      4081: inst = 32'h8220000;
      4082: inst = 32'h10408000;
      4083: inst = 32'hc404838;
      4084: inst = 32'h8220000;
      4085: inst = 32'h10408000;
      4086: inst = 32'hc404839;
      4087: inst = 32'h8220000;
      4088: inst = 32'h10408000;
      4089: inst = 32'hc40483a;
      4090: inst = 32'h8220000;
      4091: inst = 32'h10408000;
      4092: inst = 32'hc40483b;
      4093: inst = 32'h8220000;
      4094: inst = 32'h10408000;
      4095: inst = 32'hc404864;
      4096: inst = 32'h8220000;
      4097: inst = 32'h10408000;
      4098: inst = 32'hc404865;
      4099: inst = 32'h8220000;
      4100: inst = 32'h10408000;
      4101: inst = 32'hc404866;
      4102: inst = 32'h8220000;
      4103: inst = 32'h10408000;
      4104: inst = 32'hc404867;
      4105: inst = 32'h8220000;
      4106: inst = 32'h10408000;
      4107: inst = 32'hc404868;
      4108: inst = 32'h8220000;
      4109: inst = 32'h10408000;
      4110: inst = 32'hc404869;
      4111: inst = 32'h8220000;
      4112: inst = 32'h10408000;
      4113: inst = 32'hc40486a;
      4114: inst = 32'h8220000;
      4115: inst = 32'h10408000;
      4116: inst = 32'hc40486b;
      4117: inst = 32'h8220000;
      4118: inst = 32'h10408000;
      4119: inst = 32'hc40486c;
      4120: inst = 32'h8220000;
      4121: inst = 32'h10408000;
      4122: inst = 32'hc40486d;
      4123: inst = 32'h8220000;
      4124: inst = 32'h10408000;
      4125: inst = 32'hc40486e;
      4126: inst = 32'h8220000;
      4127: inst = 32'h10408000;
      4128: inst = 32'hc404880;
      4129: inst = 32'h8220000;
      4130: inst = 32'h10408000;
      4131: inst = 32'hc404881;
      4132: inst = 32'h8220000;
      4133: inst = 32'h10408000;
      4134: inst = 32'hc404882;
      4135: inst = 32'h8220000;
      4136: inst = 32'h10408000;
      4137: inst = 32'hc404883;
      4138: inst = 32'h8220000;
      4139: inst = 32'h10408000;
      4140: inst = 32'hc404884;
      4141: inst = 32'h8220000;
      4142: inst = 32'h10408000;
      4143: inst = 32'hc404885;
      4144: inst = 32'h8220000;
      4145: inst = 32'h10408000;
      4146: inst = 32'hc404886;
      4147: inst = 32'h8220000;
      4148: inst = 32'h10408000;
      4149: inst = 32'hc404887;
      4150: inst = 32'h8220000;
      4151: inst = 32'h10408000;
      4152: inst = 32'hc404888;
      4153: inst = 32'h8220000;
      4154: inst = 32'h10408000;
      4155: inst = 32'hc404889;
      4156: inst = 32'h8220000;
      4157: inst = 32'h10408000;
      4158: inst = 32'hc40488a;
      4159: inst = 32'h8220000;
      4160: inst = 32'h10408000;
      4161: inst = 32'hc40488b;
      4162: inst = 32'h8220000;
      4163: inst = 32'h10408000;
      4164: inst = 32'hc40488c;
      4165: inst = 32'h8220000;
      4166: inst = 32'h10408000;
      4167: inst = 32'hc40488d;
      4168: inst = 32'h8220000;
      4169: inst = 32'h10408000;
      4170: inst = 32'hc40488e;
      4171: inst = 32'h8220000;
      4172: inst = 32'h10408000;
      4173: inst = 32'hc40488f;
      4174: inst = 32'h8220000;
      4175: inst = 32'h10408000;
      4176: inst = 32'hc404890;
      4177: inst = 32'h8220000;
      4178: inst = 32'h10408000;
      4179: inst = 32'hc404891;
      4180: inst = 32'h8220000;
      4181: inst = 32'h10408000;
      4182: inst = 32'hc404892;
      4183: inst = 32'h8220000;
      4184: inst = 32'h10408000;
      4185: inst = 32'hc404893;
      4186: inst = 32'h8220000;
      4187: inst = 32'h10408000;
      4188: inst = 32'hc404894;
      4189: inst = 32'h8220000;
      4190: inst = 32'h10408000;
      4191: inst = 32'hc404895;
      4192: inst = 32'h8220000;
      4193: inst = 32'h10408000;
      4194: inst = 32'hc404896;
      4195: inst = 32'h8220000;
      4196: inst = 32'h10408000;
      4197: inst = 32'hc404897;
      4198: inst = 32'h8220000;
      4199: inst = 32'h10408000;
      4200: inst = 32'hc404898;
      4201: inst = 32'h8220000;
      4202: inst = 32'h10408000;
      4203: inst = 32'hc404899;
      4204: inst = 32'h8220000;
      4205: inst = 32'h10408000;
      4206: inst = 32'hc40489a;
      4207: inst = 32'h8220000;
      4208: inst = 32'h10408000;
      4209: inst = 32'hc40489b;
      4210: inst = 32'h8220000;
      4211: inst = 32'h10408000;
      4212: inst = 32'hc4048c4;
      4213: inst = 32'h8220000;
      4214: inst = 32'h10408000;
      4215: inst = 32'hc4048c5;
      4216: inst = 32'h8220000;
      4217: inst = 32'h10408000;
      4218: inst = 32'hc4048c6;
      4219: inst = 32'h8220000;
      4220: inst = 32'h10408000;
      4221: inst = 32'hc4048c7;
      4222: inst = 32'h8220000;
      4223: inst = 32'h10408000;
      4224: inst = 32'hc4048c8;
      4225: inst = 32'h8220000;
      4226: inst = 32'h10408000;
      4227: inst = 32'hc4048c9;
      4228: inst = 32'h8220000;
      4229: inst = 32'h10408000;
      4230: inst = 32'hc4048ca;
      4231: inst = 32'h8220000;
      4232: inst = 32'h10408000;
      4233: inst = 32'hc4048cb;
      4234: inst = 32'h8220000;
      4235: inst = 32'h10408000;
      4236: inst = 32'hc4048cc;
      4237: inst = 32'h8220000;
      4238: inst = 32'h10408000;
      4239: inst = 32'hc4048cd;
      4240: inst = 32'h8220000;
      4241: inst = 32'h10408000;
      4242: inst = 32'hc4048ce;
      4243: inst = 32'h8220000;
      4244: inst = 32'h10408000;
      4245: inst = 32'hc4048e0;
      4246: inst = 32'h8220000;
      4247: inst = 32'h10408000;
      4248: inst = 32'hc4048e1;
      4249: inst = 32'h8220000;
      4250: inst = 32'h10408000;
      4251: inst = 32'hc4048e2;
      4252: inst = 32'h8220000;
      4253: inst = 32'h10408000;
      4254: inst = 32'hc4048e3;
      4255: inst = 32'h8220000;
      4256: inst = 32'h10408000;
      4257: inst = 32'hc4048e4;
      4258: inst = 32'h8220000;
      4259: inst = 32'h10408000;
      4260: inst = 32'hc4048e5;
      4261: inst = 32'h8220000;
      4262: inst = 32'h10408000;
      4263: inst = 32'hc4048e6;
      4264: inst = 32'h8220000;
      4265: inst = 32'h10408000;
      4266: inst = 32'hc4048e7;
      4267: inst = 32'h8220000;
      4268: inst = 32'h10408000;
      4269: inst = 32'hc4048e8;
      4270: inst = 32'h8220000;
      4271: inst = 32'h10408000;
      4272: inst = 32'hc4048e9;
      4273: inst = 32'h8220000;
      4274: inst = 32'h10408000;
      4275: inst = 32'hc4048ea;
      4276: inst = 32'h8220000;
      4277: inst = 32'h10408000;
      4278: inst = 32'hc4048eb;
      4279: inst = 32'h8220000;
      4280: inst = 32'h10408000;
      4281: inst = 32'hc4048ec;
      4282: inst = 32'h8220000;
      4283: inst = 32'h10408000;
      4284: inst = 32'hc4048ed;
      4285: inst = 32'h8220000;
      4286: inst = 32'h10408000;
      4287: inst = 32'hc4048ee;
      4288: inst = 32'h8220000;
      4289: inst = 32'h10408000;
      4290: inst = 32'hc4048ef;
      4291: inst = 32'h8220000;
      4292: inst = 32'h10408000;
      4293: inst = 32'hc4048f0;
      4294: inst = 32'h8220000;
      4295: inst = 32'h10408000;
      4296: inst = 32'hc4048f1;
      4297: inst = 32'h8220000;
      4298: inst = 32'h10408000;
      4299: inst = 32'hc4048f2;
      4300: inst = 32'h8220000;
      4301: inst = 32'h10408000;
      4302: inst = 32'hc4048f3;
      4303: inst = 32'h8220000;
      4304: inst = 32'h10408000;
      4305: inst = 32'hc4048f4;
      4306: inst = 32'h8220000;
      4307: inst = 32'h10408000;
      4308: inst = 32'hc4048f5;
      4309: inst = 32'h8220000;
      4310: inst = 32'h10408000;
      4311: inst = 32'hc4048f6;
      4312: inst = 32'h8220000;
      4313: inst = 32'h10408000;
      4314: inst = 32'hc4048f7;
      4315: inst = 32'h8220000;
      4316: inst = 32'h10408000;
      4317: inst = 32'hc4048f8;
      4318: inst = 32'h8220000;
      4319: inst = 32'h10408000;
      4320: inst = 32'hc4048f9;
      4321: inst = 32'h8220000;
      4322: inst = 32'h10408000;
      4323: inst = 32'hc4048fa;
      4324: inst = 32'h8220000;
      4325: inst = 32'h10408000;
      4326: inst = 32'hc4048fb;
      4327: inst = 32'h8220000;
      4328: inst = 32'h10408000;
      4329: inst = 32'hc404924;
      4330: inst = 32'h8220000;
      4331: inst = 32'h10408000;
      4332: inst = 32'hc404925;
      4333: inst = 32'h8220000;
      4334: inst = 32'h10408000;
      4335: inst = 32'hc404926;
      4336: inst = 32'h8220000;
      4337: inst = 32'h10408000;
      4338: inst = 32'hc404927;
      4339: inst = 32'h8220000;
      4340: inst = 32'h10408000;
      4341: inst = 32'hc404928;
      4342: inst = 32'h8220000;
      4343: inst = 32'h10408000;
      4344: inst = 32'hc404929;
      4345: inst = 32'h8220000;
      4346: inst = 32'h10408000;
      4347: inst = 32'hc40492a;
      4348: inst = 32'h8220000;
      4349: inst = 32'h10408000;
      4350: inst = 32'hc40492b;
      4351: inst = 32'h8220000;
      4352: inst = 32'h10408000;
      4353: inst = 32'hc40492c;
      4354: inst = 32'h8220000;
      4355: inst = 32'h10408000;
      4356: inst = 32'hc40492d;
      4357: inst = 32'h8220000;
      4358: inst = 32'h10408000;
      4359: inst = 32'hc40492e;
      4360: inst = 32'h8220000;
      4361: inst = 32'h10408000;
      4362: inst = 32'hc404940;
      4363: inst = 32'h8220000;
      4364: inst = 32'h10408000;
      4365: inst = 32'hc404941;
      4366: inst = 32'h8220000;
      4367: inst = 32'h10408000;
      4368: inst = 32'hc404942;
      4369: inst = 32'h8220000;
      4370: inst = 32'h10408000;
      4371: inst = 32'hc404943;
      4372: inst = 32'h8220000;
      4373: inst = 32'h10408000;
      4374: inst = 32'hc404944;
      4375: inst = 32'h8220000;
      4376: inst = 32'h10408000;
      4377: inst = 32'hc404945;
      4378: inst = 32'h8220000;
      4379: inst = 32'h10408000;
      4380: inst = 32'hc404946;
      4381: inst = 32'h8220000;
      4382: inst = 32'h10408000;
      4383: inst = 32'hc404947;
      4384: inst = 32'h8220000;
      4385: inst = 32'h10408000;
      4386: inst = 32'hc404948;
      4387: inst = 32'h8220000;
      4388: inst = 32'h10408000;
      4389: inst = 32'hc404949;
      4390: inst = 32'h8220000;
      4391: inst = 32'h10408000;
      4392: inst = 32'hc40494a;
      4393: inst = 32'h8220000;
      4394: inst = 32'h10408000;
      4395: inst = 32'hc40494b;
      4396: inst = 32'h8220000;
      4397: inst = 32'h10408000;
      4398: inst = 32'hc40494c;
      4399: inst = 32'h8220000;
      4400: inst = 32'h10408000;
      4401: inst = 32'hc40494d;
      4402: inst = 32'h8220000;
      4403: inst = 32'h10408000;
      4404: inst = 32'hc40494e;
      4405: inst = 32'h8220000;
      4406: inst = 32'h10408000;
      4407: inst = 32'hc40494f;
      4408: inst = 32'h8220000;
      4409: inst = 32'h10408000;
      4410: inst = 32'hc404950;
      4411: inst = 32'h8220000;
      4412: inst = 32'h10408000;
      4413: inst = 32'hc404951;
      4414: inst = 32'h8220000;
      4415: inst = 32'h10408000;
      4416: inst = 32'hc404952;
      4417: inst = 32'h8220000;
      4418: inst = 32'h10408000;
      4419: inst = 32'hc404953;
      4420: inst = 32'h8220000;
      4421: inst = 32'h10408000;
      4422: inst = 32'hc404954;
      4423: inst = 32'h8220000;
      4424: inst = 32'h10408000;
      4425: inst = 32'hc404955;
      4426: inst = 32'h8220000;
      4427: inst = 32'h10408000;
      4428: inst = 32'hc404956;
      4429: inst = 32'h8220000;
      4430: inst = 32'h10408000;
      4431: inst = 32'hc404957;
      4432: inst = 32'h8220000;
      4433: inst = 32'h10408000;
      4434: inst = 32'hc404958;
      4435: inst = 32'h8220000;
      4436: inst = 32'h10408000;
      4437: inst = 32'hc404959;
      4438: inst = 32'h8220000;
      4439: inst = 32'h10408000;
      4440: inst = 32'hc40495a;
      4441: inst = 32'h8220000;
      4442: inst = 32'h10408000;
      4443: inst = 32'hc40495b;
      4444: inst = 32'h8220000;
      4445: inst = 32'h10408000;
      4446: inst = 32'hc404984;
      4447: inst = 32'h8220000;
      4448: inst = 32'h10408000;
      4449: inst = 32'hc404985;
      4450: inst = 32'h8220000;
      4451: inst = 32'h10408000;
      4452: inst = 32'hc404986;
      4453: inst = 32'h8220000;
      4454: inst = 32'h10408000;
      4455: inst = 32'hc404987;
      4456: inst = 32'h8220000;
      4457: inst = 32'h10408000;
      4458: inst = 32'hc404988;
      4459: inst = 32'h8220000;
      4460: inst = 32'h10408000;
      4461: inst = 32'hc404989;
      4462: inst = 32'h8220000;
      4463: inst = 32'h10408000;
      4464: inst = 32'hc40498a;
      4465: inst = 32'h8220000;
      4466: inst = 32'h10408000;
      4467: inst = 32'hc40498b;
      4468: inst = 32'h8220000;
      4469: inst = 32'h10408000;
      4470: inst = 32'hc40498c;
      4471: inst = 32'h8220000;
      4472: inst = 32'h10408000;
      4473: inst = 32'hc40498d;
      4474: inst = 32'h8220000;
      4475: inst = 32'h10408000;
      4476: inst = 32'hc40498e;
      4477: inst = 32'h8220000;
      4478: inst = 32'h10408000;
      4479: inst = 32'hc4049a0;
      4480: inst = 32'h8220000;
      4481: inst = 32'h10408000;
      4482: inst = 32'hc4049a1;
      4483: inst = 32'h8220000;
      4484: inst = 32'h10408000;
      4485: inst = 32'hc4049a2;
      4486: inst = 32'h8220000;
      4487: inst = 32'h10408000;
      4488: inst = 32'hc4049a3;
      4489: inst = 32'h8220000;
      4490: inst = 32'h10408000;
      4491: inst = 32'hc4049a4;
      4492: inst = 32'h8220000;
      4493: inst = 32'h10408000;
      4494: inst = 32'hc4049a5;
      4495: inst = 32'h8220000;
      4496: inst = 32'h10408000;
      4497: inst = 32'hc4049a6;
      4498: inst = 32'h8220000;
      4499: inst = 32'h10408000;
      4500: inst = 32'hc4049a7;
      4501: inst = 32'h8220000;
      4502: inst = 32'h10408000;
      4503: inst = 32'hc4049a8;
      4504: inst = 32'h8220000;
      4505: inst = 32'h10408000;
      4506: inst = 32'hc4049a9;
      4507: inst = 32'h8220000;
      4508: inst = 32'h10408000;
      4509: inst = 32'hc4049aa;
      4510: inst = 32'h8220000;
      4511: inst = 32'h10408000;
      4512: inst = 32'hc4049ab;
      4513: inst = 32'h8220000;
      4514: inst = 32'h10408000;
      4515: inst = 32'hc4049ac;
      4516: inst = 32'h8220000;
      4517: inst = 32'h10408000;
      4518: inst = 32'hc4049ad;
      4519: inst = 32'h8220000;
      4520: inst = 32'h10408000;
      4521: inst = 32'hc4049ae;
      4522: inst = 32'h8220000;
      4523: inst = 32'h10408000;
      4524: inst = 32'hc4049af;
      4525: inst = 32'h8220000;
      4526: inst = 32'h10408000;
      4527: inst = 32'hc4049b0;
      4528: inst = 32'h8220000;
      4529: inst = 32'h10408000;
      4530: inst = 32'hc4049b1;
      4531: inst = 32'h8220000;
      4532: inst = 32'h10408000;
      4533: inst = 32'hc4049b2;
      4534: inst = 32'h8220000;
      4535: inst = 32'h10408000;
      4536: inst = 32'hc4049b3;
      4537: inst = 32'h8220000;
      4538: inst = 32'h10408000;
      4539: inst = 32'hc4049b4;
      4540: inst = 32'h8220000;
      4541: inst = 32'h10408000;
      4542: inst = 32'hc4049b5;
      4543: inst = 32'h8220000;
      4544: inst = 32'h10408000;
      4545: inst = 32'hc4049b6;
      4546: inst = 32'h8220000;
      4547: inst = 32'h10408000;
      4548: inst = 32'hc4049b7;
      4549: inst = 32'h8220000;
      4550: inst = 32'h10408000;
      4551: inst = 32'hc4049b8;
      4552: inst = 32'h8220000;
      4553: inst = 32'h10408000;
      4554: inst = 32'hc4049b9;
      4555: inst = 32'h8220000;
      4556: inst = 32'h10408000;
      4557: inst = 32'hc4049ba;
      4558: inst = 32'h8220000;
      4559: inst = 32'h10408000;
      4560: inst = 32'hc4049bb;
      4561: inst = 32'h8220000;
      4562: inst = 32'h10408000;
      4563: inst = 32'hc4049e4;
      4564: inst = 32'h8220000;
      4565: inst = 32'h10408000;
      4566: inst = 32'hc4049e5;
      4567: inst = 32'h8220000;
      4568: inst = 32'h10408000;
      4569: inst = 32'hc4049e6;
      4570: inst = 32'h8220000;
      4571: inst = 32'h10408000;
      4572: inst = 32'hc4049e7;
      4573: inst = 32'h8220000;
      4574: inst = 32'h10408000;
      4575: inst = 32'hc4049e8;
      4576: inst = 32'h8220000;
      4577: inst = 32'h10408000;
      4578: inst = 32'hc4049e9;
      4579: inst = 32'h8220000;
      4580: inst = 32'h10408000;
      4581: inst = 32'hc4049ea;
      4582: inst = 32'h8220000;
      4583: inst = 32'h10408000;
      4584: inst = 32'hc4049eb;
      4585: inst = 32'h8220000;
      4586: inst = 32'h10408000;
      4587: inst = 32'hc4049ec;
      4588: inst = 32'h8220000;
      4589: inst = 32'h10408000;
      4590: inst = 32'hc4049ed;
      4591: inst = 32'h8220000;
      4592: inst = 32'h10408000;
      4593: inst = 32'hc4049ee;
      4594: inst = 32'h8220000;
      4595: inst = 32'h10408000;
      4596: inst = 32'hc404a00;
      4597: inst = 32'h8220000;
      4598: inst = 32'h10408000;
      4599: inst = 32'hc404a01;
      4600: inst = 32'h8220000;
      4601: inst = 32'h10408000;
      4602: inst = 32'hc404a02;
      4603: inst = 32'h8220000;
      4604: inst = 32'h10408000;
      4605: inst = 32'hc404a03;
      4606: inst = 32'h8220000;
      4607: inst = 32'h10408000;
      4608: inst = 32'hc404a04;
      4609: inst = 32'h8220000;
      4610: inst = 32'h10408000;
      4611: inst = 32'hc404a05;
      4612: inst = 32'h8220000;
      4613: inst = 32'h10408000;
      4614: inst = 32'hc404a06;
      4615: inst = 32'h8220000;
      4616: inst = 32'h10408000;
      4617: inst = 32'hc404a07;
      4618: inst = 32'h8220000;
      4619: inst = 32'h10408000;
      4620: inst = 32'hc404a0f;
      4621: inst = 32'h8220000;
      4622: inst = 32'h10408000;
      4623: inst = 32'hc404a10;
      4624: inst = 32'h8220000;
      4625: inst = 32'h10408000;
      4626: inst = 32'hc404a11;
      4627: inst = 32'h8220000;
      4628: inst = 32'h10408000;
      4629: inst = 32'hc404a12;
      4630: inst = 32'h8220000;
      4631: inst = 32'h10408000;
      4632: inst = 32'hc404a13;
      4633: inst = 32'h8220000;
      4634: inst = 32'h10408000;
      4635: inst = 32'hc404a14;
      4636: inst = 32'h8220000;
      4637: inst = 32'h10408000;
      4638: inst = 32'hc404a15;
      4639: inst = 32'h8220000;
      4640: inst = 32'h10408000;
      4641: inst = 32'hc404a16;
      4642: inst = 32'h8220000;
      4643: inst = 32'h10408000;
      4644: inst = 32'hc404a17;
      4645: inst = 32'h8220000;
      4646: inst = 32'h10408000;
      4647: inst = 32'hc404a18;
      4648: inst = 32'h8220000;
      4649: inst = 32'h10408000;
      4650: inst = 32'hc404a19;
      4651: inst = 32'h8220000;
      4652: inst = 32'h10408000;
      4653: inst = 32'hc404a1a;
      4654: inst = 32'h8220000;
      4655: inst = 32'h10408000;
      4656: inst = 32'hc404a1b;
      4657: inst = 32'h8220000;
      4658: inst = 32'h10408000;
      4659: inst = 32'hc404a44;
      4660: inst = 32'h8220000;
      4661: inst = 32'h10408000;
      4662: inst = 32'hc404a45;
      4663: inst = 32'h8220000;
      4664: inst = 32'h10408000;
      4665: inst = 32'hc404a46;
      4666: inst = 32'h8220000;
      4667: inst = 32'h10408000;
      4668: inst = 32'hc404a47;
      4669: inst = 32'h8220000;
      4670: inst = 32'h10408000;
      4671: inst = 32'hc404a48;
      4672: inst = 32'h8220000;
      4673: inst = 32'h10408000;
      4674: inst = 32'hc404a49;
      4675: inst = 32'h8220000;
      4676: inst = 32'h10408000;
      4677: inst = 32'hc404a4a;
      4678: inst = 32'h8220000;
      4679: inst = 32'h10408000;
      4680: inst = 32'hc404a4b;
      4681: inst = 32'h8220000;
      4682: inst = 32'h10408000;
      4683: inst = 32'hc404a4c;
      4684: inst = 32'h8220000;
      4685: inst = 32'h10408000;
      4686: inst = 32'hc404a4d;
      4687: inst = 32'h8220000;
      4688: inst = 32'h10408000;
      4689: inst = 32'hc404a4e;
      4690: inst = 32'h8220000;
      4691: inst = 32'h10408000;
      4692: inst = 32'hc404a60;
      4693: inst = 32'h8220000;
      4694: inst = 32'h10408000;
      4695: inst = 32'hc404a61;
      4696: inst = 32'h8220000;
      4697: inst = 32'h10408000;
      4698: inst = 32'hc404a62;
      4699: inst = 32'h8220000;
      4700: inst = 32'h10408000;
      4701: inst = 32'hc404a63;
      4702: inst = 32'h8220000;
      4703: inst = 32'h10408000;
      4704: inst = 32'hc404a64;
      4705: inst = 32'h8220000;
      4706: inst = 32'h10408000;
      4707: inst = 32'hc404a65;
      4708: inst = 32'h8220000;
      4709: inst = 32'h10408000;
      4710: inst = 32'hc404a66;
      4711: inst = 32'h8220000;
      4712: inst = 32'h10408000;
      4713: inst = 32'hc404a70;
      4714: inst = 32'h8220000;
      4715: inst = 32'h10408000;
      4716: inst = 32'hc404a71;
      4717: inst = 32'h8220000;
      4718: inst = 32'h10408000;
      4719: inst = 32'hc404a72;
      4720: inst = 32'h8220000;
      4721: inst = 32'h10408000;
      4722: inst = 32'hc404a73;
      4723: inst = 32'h8220000;
      4724: inst = 32'h10408000;
      4725: inst = 32'hc404a74;
      4726: inst = 32'h8220000;
      4727: inst = 32'h10408000;
      4728: inst = 32'hc404a75;
      4729: inst = 32'h8220000;
      4730: inst = 32'h10408000;
      4731: inst = 32'hc404a76;
      4732: inst = 32'h8220000;
      4733: inst = 32'h10408000;
      4734: inst = 32'hc404a77;
      4735: inst = 32'h8220000;
      4736: inst = 32'h10408000;
      4737: inst = 32'hc404a78;
      4738: inst = 32'h8220000;
      4739: inst = 32'h10408000;
      4740: inst = 32'hc404a79;
      4741: inst = 32'h8220000;
      4742: inst = 32'h10408000;
      4743: inst = 32'hc404a7a;
      4744: inst = 32'h8220000;
      4745: inst = 32'h10408000;
      4746: inst = 32'hc404a7b;
      4747: inst = 32'h8220000;
      4748: inst = 32'h10408000;
      4749: inst = 32'hc404aa4;
      4750: inst = 32'h8220000;
      4751: inst = 32'h10408000;
      4752: inst = 32'hc404aa5;
      4753: inst = 32'h8220000;
      4754: inst = 32'h10408000;
      4755: inst = 32'hc404aa6;
      4756: inst = 32'h8220000;
      4757: inst = 32'h10408000;
      4758: inst = 32'hc404aa7;
      4759: inst = 32'h8220000;
      4760: inst = 32'h10408000;
      4761: inst = 32'hc404aa8;
      4762: inst = 32'h8220000;
      4763: inst = 32'h10408000;
      4764: inst = 32'hc404aa9;
      4765: inst = 32'h8220000;
      4766: inst = 32'h10408000;
      4767: inst = 32'hc404aaa;
      4768: inst = 32'h8220000;
      4769: inst = 32'h10408000;
      4770: inst = 32'hc404aab;
      4771: inst = 32'h8220000;
      4772: inst = 32'h10408000;
      4773: inst = 32'hc404aac;
      4774: inst = 32'h8220000;
      4775: inst = 32'h10408000;
      4776: inst = 32'hc404aad;
      4777: inst = 32'h8220000;
      4778: inst = 32'h10408000;
      4779: inst = 32'hc404aae;
      4780: inst = 32'h8220000;
      4781: inst = 32'h10408000;
      4782: inst = 32'hc404ac0;
      4783: inst = 32'h8220000;
      4784: inst = 32'h10408000;
      4785: inst = 32'hc404ac1;
      4786: inst = 32'h8220000;
      4787: inst = 32'h10408000;
      4788: inst = 32'hc404ac2;
      4789: inst = 32'h8220000;
      4790: inst = 32'h10408000;
      4791: inst = 32'hc404ac3;
      4792: inst = 32'h8220000;
      4793: inst = 32'h10408000;
      4794: inst = 32'hc404ac4;
      4795: inst = 32'h8220000;
      4796: inst = 32'h10408000;
      4797: inst = 32'hc404ac5;
      4798: inst = 32'h8220000;
      4799: inst = 32'h10408000;
      4800: inst = 32'hc404ac6;
      4801: inst = 32'h8220000;
      4802: inst = 32'h10408000;
      4803: inst = 32'hc404ad0;
      4804: inst = 32'h8220000;
      4805: inst = 32'h10408000;
      4806: inst = 32'hc404ad1;
      4807: inst = 32'h8220000;
      4808: inst = 32'h10408000;
      4809: inst = 32'hc404ad2;
      4810: inst = 32'h8220000;
      4811: inst = 32'h10408000;
      4812: inst = 32'hc404ad3;
      4813: inst = 32'h8220000;
      4814: inst = 32'h10408000;
      4815: inst = 32'hc404ad4;
      4816: inst = 32'h8220000;
      4817: inst = 32'h10408000;
      4818: inst = 32'hc404ad5;
      4819: inst = 32'h8220000;
      4820: inst = 32'h10408000;
      4821: inst = 32'hc404ad6;
      4822: inst = 32'h8220000;
      4823: inst = 32'h10408000;
      4824: inst = 32'hc404ad7;
      4825: inst = 32'h8220000;
      4826: inst = 32'h10408000;
      4827: inst = 32'hc404ad8;
      4828: inst = 32'h8220000;
      4829: inst = 32'h10408000;
      4830: inst = 32'hc404ad9;
      4831: inst = 32'h8220000;
      4832: inst = 32'h10408000;
      4833: inst = 32'hc404ada;
      4834: inst = 32'h8220000;
      4835: inst = 32'h10408000;
      4836: inst = 32'hc404adb;
      4837: inst = 32'h8220000;
      4838: inst = 32'h10408000;
      4839: inst = 32'hc404b04;
      4840: inst = 32'h8220000;
      4841: inst = 32'h10408000;
      4842: inst = 32'hc404b05;
      4843: inst = 32'h8220000;
      4844: inst = 32'h10408000;
      4845: inst = 32'hc404b06;
      4846: inst = 32'h8220000;
      4847: inst = 32'h10408000;
      4848: inst = 32'hc404b07;
      4849: inst = 32'h8220000;
      4850: inst = 32'h10408000;
      4851: inst = 32'hc404b08;
      4852: inst = 32'h8220000;
      4853: inst = 32'h10408000;
      4854: inst = 32'hc404b09;
      4855: inst = 32'h8220000;
      4856: inst = 32'h10408000;
      4857: inst = 32'hc404b0a;
      4858: inst = 32'h8220000;
      4859: inst = 32'h10408000;
      4860: inst = 32'hc404b0b;
      4861: inst = 32'h8220000;
      4862: inst = 32'h10408000;
      4863: inst = 32'hc404b0c;
      4864: inst = 32'h8220000;
      4865: inst = 32'h10408000;
      4866: inst = 32'hc404b0d;
      4867: inst = 32'h8220000;
      4868: inst = 32'h10408000;
      4869: inst = 32'hc404b0e;
      4870: inst = 32'h8220000;
      4871: inst = 32'h10408000;
      4872: inst = 32'hc404b20;
      4873: inst = 32'h8220000;
      4874: inst = 32'h10408000;
      4875: inst = 32'hc404b21;
      4876: inst = 32'h8220000;
      4877: inst = 32'h10408000;
      4878: inst = 32'hc404b22;
      4879: inst = 32'h8220000;
      4880: inst = 32'h10408000;
      4881: inst = 32'hc404b23;
      4882: inst = 32'h8220000;
      4883: inst = 32'h10408000;
      4884: inst = 32'hc404b24;
      4885: inst = 32'h8220000;
      4886: inst = 32'h10408000;
      4887: inst = 32'hc404b25;
      4888: inst = 32'h8220000;
      4889: inst = 32'h10408000;
      4890: inst = 32'hc404b26;
      4891: inst = 32'h8220000;
      4892: inst = 32'h10408000;
      4893: inst = 32'hc404b30;
      4894: inst = 32'h8220000;
      4895: inst = 32'h10408000;
      4896: inst = 32'hc404b31;
      4897: inst = 32'h8220000;
      4898: inst = 32'h10408000;
      4899: inst = 32'hc404b32;
      4900: inst = 32'h8220000;
      4901: inst = 32'h10408000;
      4902: inst = 32'hc404b33;
      4903: inst = 32'h8220000;
      4904: inst = 32'h10408000;
      4905: inst = 32'hc404b34;
      4906: inst = 32'h8220000;
      4907: inst = 32'h10408000;
      4908: inst = 32'hc404b35;
      4909: inst = 32'h8220000;
      4910: inst = 32'h10408000;
      4911: inst = 32'hc404b36;
      4912: inst = 32'h8220000;
      4913: inst = 32'h10408000;
      4914: inst = 32'hc404b37;
      4915: inst = 32'h8220000;
      4916: inst = 32'h10408000;
      4917: inst = 32'hc404b38;
      4918: inst = 32'h8220000;
      4919: inst = 32'h10408000;
      4920: inst = 32'hc404b39;
      4921: inst = 32'h8220000;
      4922: inst = 32'h10408000;
      4923: inst = 32'hc404b3a;
      4924: inst = 32'h8220000;
      4925: inst = 32'h10408000;
      4926: inst = 32'hc404b3b;
      4927: inst = 32'h8220000;
      4928: inst = 32'h10408000;
      4929: inst = 32'hc404b64;
      4930: inst = 32'h8220000;
      4931: inst = 32'h10408000;
      4932: inst = 32'hc404b65;
      4933: inst = 32'h8220000;
      4934: inst = 32'h10408000;
      4935: inst = 32'hc404b66;
      4936: inst = 32'h8220000;
      4937: inst = 32'h10408000;
      4938: inst = 32'hc404b67;
      4939: inst = 32'h8220000;
      4940: inst = 32'h10408000;
      4941: inst = 32'hc404b68;
      4942: inst = 32'h8220000;
      4943: inst = 32'h10408000;
      4944: inst = 32'hc404b69;
      4945: inst = 32'h8220000;
      4946: inst = 32'h10408000;
      4947: inst = 32'hc404b6a;
      4948: inst = 32'h8220000;
      4949: inst = 32'h10408000;
      4950: inst = 32'hc404b6b;
      4951: inst = 32'h8220000;
      4952: inst = 32'h10408000;
      4953: inst = 32'hc404b6c;
      4954: inst = 32'h8220000;
      4955: inst = 32'h10408000;
      4956: inst = 32'hc404b6d;
      4957: inst = 32'h8220000;
      4958: inst = 32'h10408000;
      4959: inst = 32'hc404b6e;
      4960: inst = 32'h8220000;
      4961: inst = 32'h10408000;
      4962: inst = 32'hc404b80;
      4963: inst = 32'h8220000;
      4964: inst = 32'h10408000;
      4965: inst = 32'hc404b81;
      4966: inst = 32'h8220000;
      4967: inst = 32'h10408000;
      4968: inst = 32'hc404b82;
      4969: inst = 32'h8220000;
      4970: inst = 32'h10408000;
      4971: inst = 32'hc404b83;
      4972: inst = 32'h8220000;
      4973: inst = 32'h10408000;
      4974: inst = 32'hc404b84;
      4975: inst = 32'h8220000;
      4976: inst = 32'h10408000;
      4977: inst = 32'hc404b85;
      4978: inst = 32'h8220000;
      4979: inst = 32'h10408000;
      4980: inst = 32'hc404b86;
      4981: inst = 32'h8220000;
      4982: inst = 32'h10408000;
      4983: inst = 32'hc404b90;
      4984: inst = 32'h8220000;
      4985: inst = 32'h10408000;
      4986: inst = 32'hc404b91;
      4987: inst = 32'h8220000;
      4988: inst = 32'h10408000;
      4989: inst = 32'hc404b92;
      4990: inst = 32'h8220000;
      4991: inst = 32'h10408000;
      4992: inst = 32'hc404b93;
      4993: inst = 32'h8220000;
      4994: inst = 32'h10408000;
      4995: inst = 32'hc404b94;
      4996: inst = 32'h8220000;
      4997: inst = 32'h10408000;
      4998: inst = 32'hc404b95;
      4999: inst = 32'h8220000;
      5000: inst = 32'h10408000;
      5001: inst = 32'hc404b96;
      5002: inst = 32'h8220000;
      5003: inst = 32'h10408000;
      5004: inst = 32'hc404b97;
      5005: inst = 32'h8220000;
      5006: inst = 32'h10408000;
      5007: inst = 32'hc404b98;
      5008: inst = 32'h8220000;
      5009: inst = 32'h10408000;
      5010: inst = 32'hc404b99;
      5011: inst = 32'h8220000;
      5012: inst = 32'h10408000;
      5013: inst = 32'hc404b9a;
      5014: inst = 32'h8220000;
      5015: inst = 32'h10408000;
      5016: inst = 32'hc404b9b;
      5017: inst = 32'h8220000;
      5018: inst = 32'h10408000;
      5019: inst = 32'hc404bc4;
      5020: inst = 32'h8220000;
      5021: inst = 32'h10408000;
      5022: inst = 32'hc404bc5;
      5023: inst = 32'h8220000;
      5024: inst = 32'h10408000;
      5025: inst = 32'hc404bc6;
      5026: inst = 32'h8220000;
      5027: inst = 32'h10408000;
      5028: inst = 32'hc404bc7;
      5029: inst = 32'h8220000;
      5030: inst = 32'h10408000;
      5031: inst = 32'hc404bc8;
      5032: inst = 32'h8220000;
      5033: inst = 32'h10408000;
      5034: inst = 32'hc404bc9;
      5035: inst = 32'h8220000;
      5036: inst = 32'h10408000;
      5037: inst = 32'hc404bca;
      5038: inst = 32'h8220000;
      5039: inst = 32'h10408000;
      5040: inst = 32'hc404bcb;
      5041: inst = 32'h8220000;
      5042: inst = 32'h10408000;
      5043: inst = 32'hc404bcc;
      5044: inst = 32'h8220000;
      5045: inst = 32'h10408000;
      5046: inst = 32'hc404bcd;
      5047: inst = 32'h8220000;
      5048: inst = 32'h10408000;
      5049: inst = 32'hc404bce;
      5050: inst = 32'h8220000;
      5051: inst = 32'h10408000;
      5052: inst = 32'hc404be0;
      5053: inst = 32'h8220000;
      5054: inst = 32'h10408000;
      5055: inst = 32'hc404be1;
      5056: inst = 32'h8220000;
      5057: inst = 32'h10408000;
      5058: inst = 32'hc404be2;
      5059: inst = 32'h8220000;
      5060: inst = 32'h10408000;
      5061: inst = 32'hc404be3;
      5062: inst = 32'h8220000;
      5063: inst = 32'h10408000;
      5064: inst = 32'hc404be4;
      5065: inst = 32'h8220000;
      5066: inst = 32'h10408000;
      5067: inst = 32'hc404be5;
      5068: inst = 32'h8220000;
      5069: inst = 32'h10408000;
      5070: inst = 32'hc404be6;
      5071: inst = 32'h8220000;
      5072: inst = 32'h10408000;
      5073: inst = 32'hc404bf0;
      5074: inst = 32'h8220000;
      5075: inst = 32'h10408000;
      5076: inst = 32'hc404bf1;
      5077: inst = 32'h8220000;
      5078: inst = 32'h10408000;
      5079: inst = 32'hc404bf2;
      5080: inst = 32'h8220000;
      5081: inst = 32'h10408000;
      5082: inst = 32'hc404bf3;
      5083: inst = 32'h8220000;
      5084: inst = 32'h10408000;
      5085: inst = 32'hc404bf4;
      5086: inst = 32'h8220000;
      5087: inst = 32'h10408000;
      5088: inst = 32'hc404bf5;
      5089: inst = 32'h8220000;
      5090: inst = 32'h10408000;
      5091: inst = 32'hc404bf6;
      5092: inst = 32'h8220000;
      5093: inst = 32'h10408000;
      5094: inst = 32'hc404bf7;
      5095: inst = 32'h8220000;
      5096: inst = 32'h10408000;
      5097: inst = 32'hc404bf8;
      5098: inst = 32'h8220000;
      5099: inst = 32'h10408000;
      5100: inst = 32'hc404bf9;
      5101: inst = 32'h8220000;
      5102: inst = 32'h10408000;
      5103: inst = 32'hc404c26;
      5104: inst = 32'h8220000;
      5105: inst = 32'h10408000;
      5106: inst = 32'hc404c27;
      5107: inst = 32'h8220000;
      5108: inst = 32'h10408000;
      5109: inst = 32'hc404c28;
      5110: inst = 32'h8220000;
      5111: inst = 32'h10408000;
      5112: inst = 32'hc404c29;
      5113: inst = 32'h8220000;
      5114: inst = 32'h10408000;
      5115: inst = 32'hc404c2a;
      5116: inst = 32'h8220000;
      5117: inst = 32'h10408000;
      5118: inst = 32'hc404c2b;
      5119: inst = 32'h8220000;
      5120: inst = 32'h10408000;
      5121: inst = 32'hc404c2c;
      5122: inst = 32'h8220000;
      5123: inst = 32'h10408000;
      5124: inst = 32'hc404c2d;
      5125: inst = 32'h8220000;
      5126: inst = 32'h10408000;
      5127: inst = 32'hc404c2e;
      5128: inst = 32'h8220000;
      5129: inst = 32'h10408000;
      5130: inst = 32'hc404c40;
      5131: inst = 32'h8220000;
      5132: inst = 32'h10408000;
      5133: inst = 32'hc404c41;
      5134: inst = 32'h8220000;
      5135: inst = 32'h10408000;
      5136: inst = 32'hc404c42;
      5137: inst = 32'h8220000;
      5138: inst = 32'h10408000;
      5139: inst = 32'hc404c43;
      5140: inst = 32'h8220000;
      5141: inst = 32'h10408000;
      5142: inst = 32'hc404c44;
      5143: inst = 32'h8220000;
      5144: inst = 32'h10408000;
      5145: inst = 32'hc404c45;
      5146: inst = 32'h8220000;
      5147: inst = 32'h10408000;
      5148: inst = 32'hc404c46;
      5149: inst = 32'h8220000;
      5150: inst = 32'h10408000;
      5151: inst = 32'hc404c4f;
      5152: inst = 32'h8220000;
      5153: inst = 32'h10408000;
      5154: inst = 32'hc404c50;
      5155: inst = 32'h8220000;
      5156: inst = 32'h10408000;
      5157: inst = 32'hc404c51;
      5158: inst = 32'h8220000;
      5159: inst = 32'h10408000;
      5160: inst = 32'hc404c52;
      5161: inst = 32'h8220000;
      5162: inst = 32'h10408000;
      5163: inst = 32'hc404c53;
      5164: inst = 32'h8220000;
      5165: inst = 32'h10408000;
      5166: inst = 32'hc404c54;
      5167: inst = 32'h8220000;
      5168: inst = 32'h10408000;
      5169: inst = 32'hc404c55;
      5170: inst = 32'h8220000;
      5171: inst = 32'h10408000;
      5172: inst = 32'hc404c56;
      5173: inst = 32'h8220000;
      5174: inst = 32'h10408000;
      5175: inst = 32'hc404c57;
      5176: inst = 32'h8220000;
      5177: inst = 32'h10408000;
      5178: inst = 32'hc404c58;
      5179: inst = 32'h8220000;
      5180: inst = 32'h10408000;
      5181: inst = 32'hc404c59;
      5182: inst = 32'h8220000;
      5183: inst = 32'h10408000;
      5184: inst = 32'hc404c5a;
      5185: inst = 32'h8220000;
      5186: inst = 32'h10408000;
      5187: inst = 32'hc404c5b;
      5188: inst = 32'h8220000;
      5189: inst = 32'h10408000;
      5190: inst = 32'hc404c5c;
      5191: inst = 32'h8220000;
      5192: inst = 32'h10408000;
      5193: inst = 32'hc404c5d;
      5194: inst = 32'h8220000;
      5195: inst = 32'h10408000;
      5196: inst = 32'hc404c5e;
      5197: inst = 32'h8220000;
      5198: inst = 32'h10408000;
      5199: inst = 32'hc404c5f;
      5200: inst = 32'h8220000;
      5201: inst = 32'h10408000;
      5202: inst = 32'hc404c60;
      5203: inst = 32'h8220000;
      5204: inst = 32'h10408000;
      5205: inst = 32'hc404c61;
      5206: inst = 32'h8220000;
      5207: inst = 32'h10408000;
      5208: inst = 32'hc404c62;
      5209: inst = 32'h8220000;
      5210: inst = 32'h10408000;
      5211: inst = 32'hc404c63;
      5212: inst = 32'h8220000;
      5213: inst = 32'h10408000;
      5214: inst = 32'hc404c64;
      5215: inst = 32'h8220000;
      5216: inst = 32'h10408000;
      5217: inst = 32'hc404c65;
      5218: inst = 32'h8220000;
      5219: inst = 32'h10408000;
      5220: inst = 32'hc404c66;
      5221: inst = 32'h8220000;
      5222: inst = 32'h10408000;
      5223: inst = 32'hc404c67;
      5224: inst = 32'h8220000;
      5225: inst = 32'h10408000;
      5226: inst = 32'hc404c68;
      5227: inst = 32'h8220000;
      5228: inst = 32'h10408000;
      5229: inst = 32'hc404c69;
      5230: inst = 32'h8220000;
      5231: inst = 32'h10408000;
      5232: inst = 32'hc404c6a;
      5233: inst = 32'h8220000;
      5234: inst = 32'h10408000;
      5235: inst = 32'hc404c6b;
      5236: inst = 32'h8220000;
      5237: inst = 32'h10408000;
      5238: inst = 32'hc404c6c;
      5239: inst = 32'h8220000;
      5240: inst = 32'h10408000;
      5241: inst = 32'hc404c6d;
      5242: inst = 32'h8220000;
      5243: inst = 32'h10408000;
      5244: inst = 32'hc404c6e;
      5245: inst = 32'h8220000;
      5246: inst = 32'h10408000;
      5247: inst = 32'hc404c6f;
      5248: inst = 32'h8220000;
      5249: inst = 32'h10408000;
      5250: inst = 32'hc404c70;
      5251: inst = 32'h8220000;
      5252: inst = 32'h10408000;
      5253: inst = 32'hc404c71;
      5254: inst = 32'h8220000;
      5255: inst = 32'h10408000;
      5256: inst = 32'hc404c72;
      5257: inst = 32'h8220000;
      5258: inst = 32'h10408000;
      5259: inst = 32'hc404c73;
      5260: inst = 32'h8220000;
      5261: inst = 32'h10408000;
      5262: inst = 32'hc404c74;
      5263: inst = 32'h8220000;
      5264: inst = 32'h10408000;
      5265: inst = 32'hc404c75;
      5266: inst = 32'h8220000;
      5267: inst = 32'h10408000;
      5268: inst = 32'hc404c76;
      5269: inst = 32'h8220000;
      5270: inst = 32'h10408000;
      5271: inst = 32'hc404c77;
      5272: inst = 32'h8220000;
      5273: inst = 32'h10408000;
      5274: inst = 32'hc404c78;
      5275: inst = 32'h8220000;
      5276: inst = 32'h10408000;
      5277: inst = 32'hc404c79;
      5278: inst = 32'h8220000;
      5279: inst = 32'h10408000;
      5280: inst = 32'hc404c7a;
      5281: inst = 32'h8220000;
      5282: inst = 32'h10408000;
      5283: inst = 32'hc404c7b;
      5284: inst = 32'h8220000;
      5285: inst = 32'h10408000;
      5286: inst = 32'hc404c7c;
      5287: inst = 32'h8220000;
      5288: inst = 32'h10408000;
      5289: inst = 32'hc404c7d;
      5290: inst = 32'h8220000;
      5291: inst = 32'h10408000;
      5292: inst = 32'hc404c7e;
      5293: inst = 32'h8220000;
      5294: inst = 32'h10408000;
      5295: inst = 32'hc404c7f;
      5296: inst = 32'h8220000;
      5297: inst = 32'h10408000;
      5298: inst = 32'hc404c80;
      5299: inst = 32'h8220000;
      5300: inst = 32'h10408000;
      5301: inst = 32'hc404c81;
      5302: inst = 32'h8220000;
      5303: inst = 32'h10408000;
      5304: inst = 32'hc404c82;
      5305: inst = 32'h8220000;
      5306: inst = 32'h10408000;
      5307: inst = 32'hc404c83;
      5308: inst = 32'h8220000;
      5309: inst = 32'h10408000;
      5310: inst = 32'hc404c84;
      5311: inst = 32'h8220000;
      5312: inst = 32'h10408000;
      5313: inst = 32'hc404c85;
      5314: inst = 32'h8220000;
      5315: inst = 32'h10408000;
      5316: inst = 32'hc404c86;
      5317: inst = 32'h8220000;
      5318: inst = 32'h10408000;
      5319: inst = 32'hc404c87;
      5320: inst = 32'h8220000;
      5321: inst = 32'h10408000;
      5322: inst = 32'hc404c88;
      5323: inst = 32'h8220000;
      5324: inst = 32'h10408000;
      5325: inst = 32'hc404c89;
      5326: inst = 32'h8220000;
      5327: inst = 32'h10408000;
      5328: inst = 32'hc404c8a;
      5329: inst = 32'h8220000;
      5330: inst = 32'h10408000;
      5331: inst = 32'hc404c8b;
      5332: inst = 32'h8220000;
      5333: inst = 32'h10408000;
      5334: inst = 32'hc404c8c;
      5335: inst = 32'h8220000;
      5336: inst = 32'h10408000;
      5337: inst = 32'hc404c8d;
      5338: inst = 32'h8220000;
      5339: inst = 32'h10408000;
      5340: inst = 32'hc404c8e;
      5341: inst = 32'h8220000;
      5342: inst = 32'h10408000;
      5343: inst = 32'hc404ca0;
      5344: inst = 32'h8220000;
      5345: inst = 32'h10408000;
      5346: inst = 32'hc404ca1;
      5347: inst = 32'h8220000;
      5348: inst = 32'h10408000;
      5349: inst = 32'hc404cb7;
      5350: inst = 32'h8220000;
      5351: inst = 32'h10408000;
      5352: inst = 32'hc404cb8;
      5353: inst = 32'h8220000;
      5354: inst = 32'h10408000;
      5355: inst = 32'hc404cb9;
      5356: inst = 32'h8220000;
      5357: inst = 32'h10408000;
      5358: inst = 32'hc404cba;
      5359: inst = 32'h8220000;
      5360: inst = 32'h10408000;
      5361: inst = 32'hc404cbb;
      5362: inst = 32'h8220000;
      5363: inst = 32'h10408000;
      5364: inst = 32'hc404cbc;
      5365: inst = 32'h8220000;
      5366: inst = 32'h10408000;
      5367: inst = 32'hc404cbd;
      5368: inst = 32'h8220000;
      5369: inst = 32'h10408000;
      5370: inst = 32'hc404cbe;
      5371: inst = 32'h8220000;
      5372: inst = 32'h10408000;
      5373: inst = 32'hc404cbf;
      5374: inst = 32'h8220000;
      5375: inst = 32'h10408000;
      5376: inst = 32'hc404cc0;
      5377: inst = 32'h8220000;
      5378: inst = 32'h10408000;
      5379: inst = 32'hc404cc1;
      5380: inst = 32'h8220000;
      5381: inst = 32'h10408000;
      5382: inst = 32'hc404cc2;
      5383: inst = 32'h8220000;
      5384: inst = 32'h10408000;
      5385: inst = 32'hc404cc3;
      5386: inst = 32'h8220000;
      5387: inst = 32'h10408000;
      5388: inst = 32'hc404cc4;
      5389: inst = 32'h8220000;
      5390: inst = 32'h10408000;
      5391: inst = 32'hc404cc5;
      5392: inst = 32'h8220000;
      5393: inst = 32'h10408000;
      5394: inst = 32'hc404cc6;
      5395: inst = 32'h8220000;
      5396: inst = 32'h10408000;
      5397: inst = 32'hc404cc7;
      5398: inst = 32'h8220000;
      5399: inst = 32'h10408000;
      5400: inst = 32'hc404cc8;
      5401: inst = 32'h8220000;
      5402: inst = 32'h10408000;
      5403: inst = 32'hc404cc9;
      5404: inst = 32'h8220000;
      5405: inst = 32'h10408000;
      5406: inst = 32'hc404cca;
      5407: inst = 32'h8220000;
      5408: inst = 32'h10408000;
      5409: inst = 32'hc404ccb;
      5410: inst = 32'h8220000;
      5411: inst = 32'h10408000;
      5412: inst = 32'hc404ccc;
      5413: inst = 32'h8220000;
      5414: inst = 32'h10408000;
      5415: inst = 32'hc404ccd;
      5416: inst = 32'h8220000;
      5417: inst = 32'h10408000;
      5418: inst = 32'hc404cce;
      5419: inst = 32'h8220000;
      5420: inst = 32'h10408000;
      5421: inst = 32'hc404ccf;
      5422: inst = 32'h8220000;
      5423: inst = 32'h10408000;
      5424: inst = 32'hc404cd0;
      5425: inst = 32'h8220000;
      5426: inst = 32'h10408000;
      5427: inst = 32'hc404cd1;
      5428: inst = 32'h8220000;
      5429: inst = 32'h10408000;
      5430: inst = 32'hc404cd2;
      5431: inst = 32'h8220000;
      5432: inst = 32'h10408000;
      5433: inst = 32'hc404cd3;
      5434: inst = 32'h8220000;
      5435: inst = 32'h10408000;
      5436: inst = 32'hc404cd4;
      5437: inst = 32'h8220000;
      5438: inst = 32'h10408000;
      5439: inst = 32'hc404cd5;
      5440: inst = 32'h8220000;
      5441: inst = 32'h10408000;
      5442: inst = 32'hc404cd6;
      5443: inst = 32'h8220000;
      5444: inst = 32'h10408000;
      5445: inst = 32'hc404cd7;
      5446: inst = 32'h8220000;
      5447: inst = 32'h10408000;
      5448: inst = 32'hc404cd8;
      5449: inst = 32'h8220000;
      5450: inst = 32'h10408000;
      5451: inst = 32'hc404cd9;
      5452: inst = 32'h8220000;
      5453: inst = 32'h10408000;
      5454: inst = 32'hc404cda;
      5455: inst = 32'h8220000;
      5456: inst = 32'h10408000;
      5457: inst = 32'hc404cdb;
      5458: inst = 32'h8220000;
      5459: inst = 32'h10408000;
      5460: inst = 32'hc404cdc;
      5461: inst = 32'h8220000;
      5462: inst = 32'h10408000;
      5463: inst = 32'hc404cdd;
      5464: inst = 32'h8220000;
      5465: inst = 32'h10408000;
      5466: inst = 32'hc404cde;
      5467: inst = 32'h8220000;
      5468: inst = 32'h10408000;
      5469: inst = 32'hc404cdf;
      5470: inst = 32'h8220000;
      5471: inst = 32'h10408000;
      5472: inst = 32'hc404ce0;
      5473: inst = 32'h8220000;
      5474: inst = 32'h10408000;
      5475: inst = 32'hc404ce1;
      5476: inst = 32'h8220000;
      5477: inst = 32'h10408000;
      5478: inst = 32'hc404ce2;
      5479: inst = 32'h8220000;
      5480: inst = 32'h10408000;
      5481: inst = 32'hc404ce3;
      5482: inst = 32'h8220000;
      5483: inst = 32'h10408000;
      5484: inst = 32'hc404ce4;
      5485: inst = 32'h8220000;
      5486: inst = 32'h10408000;
      5487: inst = 32'hc404ce5;
      5488: inst = 32'h8220000;
      5489: inst = 32'h10408000;
      5490: inst = 32'hc404ce6;
      5491: inst = 32'h8220000;
      5492: inst = 32'h10408000;
      5493: inst = 32'hc404ce7;
      5494: inst = 32'h8220000;
      5495: inst = 32'h10408000;
      5496: inst = 32'hc404ce8;
      5497: inst = 32'h8220000;
      5498: inst = 32'h10408000;
      5499: inst = 32'hc404ce9;
      5500: inst = 32'h8220000;
      5501: inst = 32'h10408000;
      5502: inst = 32'hc404cea;
      5503: inst = 32'h8220000;
      5504: inst = 32'h10408000;
      5505: inst = 32'hc404ceb;
      5506: inst = 32'h8220000;
      5507: inst = 32'h10408000;
      5508: inst = 32'hc404cec;
      5509: inst = 32'h8220000;
      5510: inst = 32'h10408000;
      5511: inst = 32'hc404ced;
      5512: inst = 32'h8220000;
      5513: inst = 32'h10408000;
      5514: inst = 32'hc404cee;
      5515: inst = 32'h8220000;
      5516: inst = 32'h10408000;
      5517: inst = 32'hc404d17;
      5518: inst = 32'h8220000;
      5519: inst = 32'h10408000;
      5520: inst = 32'hc404d18;
      5521: inst = 32'h8220000;
      5522: inst = 32'h10408000;
      5523: inst = 32'hc404d19;
      5524: inst = 32'h8220000;
      5525: inst = 32'h10408000;
      5526: inst = 32'hc404d1a;
      5527: inst = 32'h8220000;
      5528: inst = 32'h10408000;
      5529: inst = 32'hc404d1b;
      5530: inst = 32'h8220000;
      5531: inst = 32'h10408000;
      5532: inst = 32'hc404d1c;
      5533: inst = 32'h8220000;
      5534: inst = 32'h10408000;
      5535: inst = 32'hc404d1d;
      5536: inst = 32'h8220000;
      5537: inst = 32'h10408000;
      5538: inst = 32'hc404d1e;
      5539: inst = 32'h8220000;
      5540: inst = 32'h10408000;
      5541: inst = 32'hc404d1f;
      5542: inst = 32'h8220000;
      5543: inst = 32'h10408000;
      5544: inst = 32'hc404d20;
      5545: inst = 32'h8220000;
      5546: inst = 32'h10408000;
      5547: inst = 32'hc404d21;
      5548: inst = 32'h8220000;
      5549: inst = 32'h10408000;
      5550: inst = 32'hc404d22;
      5551: inst = 32'h8220000;
      5552: inst = 32'h10408000;
      5553: inst = 32'hc404d23;
      5554: inst = 32'h8220000;
      5555: inst = 32'h10408000;
      5556: inst = 32'hc404d24;
      5557: inst = 32'h8220000;
      5558: inst = 32'h10408000;
      5559: inst = 32'hc404d25;
      5560: inst = 32'h8220000;
      5561: inst = 32'h10408000;
      5562: inst = 32'hc404d26;
      5563: inst = 32'h8220000;
      5564: inst = 32'h10408000;
      5565: inst = 32'hc404d27;
      5566: inst = 32'h8220000;
      5567: inst = 32'h10408000;
      5568: inst = 32'hc404d28;
      5569: inst = 32'h8220000;
      5570: inst = 32'h10408000;
      5571: inst = 32'hc404d29;
      5572: inst = 32'h8220000;
      5573: inst = 32'h10408000;
      5574: inst = 32'hc404d2a;
      5575: inst = 32'h8220000;
      5576: inst = 32'h10408000;
      5577: inst = 32'hc404d2b;
      5578: inst = 32'h8220000;
      5579: inst = 32'h10408000;
      5580: inst = 32'hc404d2c;
      5581: inst = 32'h8220000;
      5582: inst = 32'h10408000;
      5583: inst = 32'hc404d2d;
      5584: inst = 32'h8220000;
      5585: inst = 32'h10408000;
      5586: inst = 32'hc404d2e;
      5587: inst = 32'h8220000;
      5588: inst = 32'h10408000;
      5589: inst = 32'hc404d2f;
      5590: inst = 32'h8220000;
      5591: inst = 32'h10408000;
      5592: inst = 32'hc404d30;
      5593: inst = 32'h8220000;
      5594: inst = 32'h10408000;
      5595: inst = 32'hc404d31;
      5596: inst = 32'h8220000;
      5597: inst = 32'h10408000;
      5598: inst = 32'hc404d32;
      5599: inst = 32'h8220000;
      5600: inst = 32'h10408000;
      5601: inst = 32'hc404d33;
      5602: inst = 32'h8220000;
      5603: inst = 32'h10408000;
      5604: inst = 32'hc404d34;
      5605: inst = 32'h8220000;
      5606: inst = 32'h10408000;
      5607: inst = 32'hc404d35;
      5608: inst = 32'h8220000;
      5609: inst = 32'h10408000;
      5610: inst = 32'hc404d36;
      5611: inst = 32'h8220000;
      5612: inst = 32'h10408000;
      5613: inst = 32'hc404d37;
      5614: inst = 32'h8220000;
      5615: inst = 32'h10408000;
      5616: inst = 32'hc404d38;
      5617: inst = 32'h8220000;
      5618: inst = 32'h10408000;
      5619: inst = 32'hc404d39;
      5620: inst = 32'h8220000;
      5621: inst = 32'h10408000;
      5622: inst = 32'hc404d3a;
      5623: inst = 32'h8220000;
      5624: inst = 32'h10408000;
      5625: inst = 32'hc404d3b;
      5626: inst = 32'h8220000;
      5627: inst = 32'h10408000;
      5628: inst = 32'hc404d3c;
      5629: inst = 32'h8220000;
      5630: inst = 32'h10408000;
      5631: inst = 32'hc404d3d;
      5632: inst = 32'h8220000;
      5633: inst = 32'h10408000;
      5634: inst = 32'hc404d3e;
      5635: inst = 32'h8220000;
      5636: inst = 32'h10408000;
      5637: inst = 32'hc404d3f;
      5638: inst = 32'h8220000;
      5639: inst = 32'h10408000;
      5640: inst = 32'hc404d40;
      5641: inst = 32'h8220000;
      5642: inst = 32'h10408000;
      5643: inst = 32'hc404d41;
      5644: inst = 32'h8220000;
      5645: inst = 32'h10408000;
      5646: inst = 32'hc404d42;
      5647: inst = 32'h8220000;
      5648: inst = 32'h10408000;
      5649: inst = 32'hc404d43;
      5650: inst = 32'h8220000;
      5651: inst = 32'h10408000;
      5652: inst = 32'hc404d44;
      5653: inst = 32'h8220000;
      5654: inst = 32'h10408000;
      5655: inst = 32'hc404d45;
      5656: inst = 32'h8220000;
      5657: inst = 32'h10408000;
      5658: inst = 32'hc404d46;
      5659: inst = 32'h8220000;
      5660: inst = 32'h10408000;
      5661: inst = 32'hc404d47;
      5662: inst = 32'h8220000;
      5663: inst = 32'h10408000;
      5664: inst = 32'hc404d48;
      5665: inst = 32'h8220000;
      5666: inst = 32'h10408000;
      5667: inst = 32'hc404d49;
      5668: inst = 32'h8220000;
      5669: inst = 32'h10408000;
      5670: inst = 32'hc404d4a;
      5671: inst = 32'h8220000;
      5672: inst = 32'h10408000;
      5673: inst = 32'hc404d4b;
      5674: inst = 32'h8220000;
      5675: inst = 32'h10408000;
      5676: inst = 32'hc404d4c;
      5677: inst = 32'h8220000;
      5678: inst = 32'h10408000;
      5679: inst = 32'hc404d4d;
      5680: inst = 32'h8220000;
      5681: inst = 32'h10408000;
      5682: inst = 32'hc404d4e;
      5683: inst = 32'h8220000;
      5684: inst = 32'h10408000;
      5685: inst = 32'hc404d77;
      5686: inst = 32'h8220000;
      5687: inst = 32'h10408000;
      5688: inst = 32'hc404d78;
      5689: inst = 32'h8220000;
      5690: inst = 32'h10408000;
      5691: inst = 32'hc404d79;
      5692: inst = 32'h8220000;
      5693: inst = 32'h10408000;
      5694: inst = 32'hc404d7a;
      5695: inst = 32'h8220000;
      5696: inst = 32'h10408000;
      5697: inst = 32'hc404d7b;
      5698: inst = 32'h8220000;
      5699: inst = 32'h10408000;
      5700: inst = 32'hc404d7c;
      5701: inst = 32'h8220000;
      5702: inst = 32'h10408000;
      5703: inst = 32'hc404d7d;
      5704: inst = 32'h8220000;
      5705: inst = 32'h10408000;
      5706: inst = 32'hc404d7e;
      5707: inst = 32'h8220000;
      5708: inst = 32'h10408000;
      5709: inst = 32'hc404d7f;
      5710: inst = 32'h8220000;
      5711: inst = 32'h10408000;
      5712: inst = 32'hc404d80;
      5713: inst = 32'h8220000;
      5714: inst = 32'h10408000;
      5715: inst = 32'hc404d81;
      5716: inst = 32'h8220000;
      5717: inst = 32'h10408000;
      5718: inst = 32'hc404d82;
      5719: inst = 32'h8220000;
      5720: inst = 32'h10408000;
      5721: inst = 32'hc404d83;
      5722: inst = 32'h8220000;
      5723: inst = 32'h10408000;
      5724: inst = 32'hc404d84;
      5725: inst = 32'h8220000;
      5726: inst = 32'h10408000;
      5727: inst = 32'hc404d85;
      5728: inst = 32'h8220000;
      5729: inst = 32'h10408000;
      5730: inst = 32'hc404d86;
      5731: inst = 32'h8220000;
      5732: inst = 32'h10408000;
      5733: inst = 32'hc404d87;
      5734: inst = 32'h8220000;
      5735: inst = 32'h10408000;
      5736: inst = 32'hc404d88;
      5737: inst = 32'h8220000;
      5738: inst = 32'h10408000;
      5739: inst = 32'hc404d89;
      5740: inst = 32'h8220000;
      5741: inst = 32'h10408000;
      5742: inst = 32'hc404d8a;
      5743: inst = 32'h8220000;
      5744: inst = 32'h10408000;
      5745: inst = 32'hc404d8b;
      5746: inst = 32'h8220000;
      5747: inst = 32'h10408000;
      5748: inst = 32'hc404d8c;
      5749: inst = 32'h8220000;
      5750: inst = 32'h10408000;
      5751: inst = 32'hc404d8d;
      5752: inst = 32'h8220000;
      5753: inst = 32'h10408000;
      5754: inst = 32'hc404d8e;
      5755: inst = 32'h8220000;
      5756: inst = 32'h10408000;
      5757: inst = 32'hc404d8f;
      5758: inst = 32'h8220000;
      5759: inst = 32'h10408000;
      5760: inst = 32'hc404d90;
      5761: inst = 32'h8220000;
      5762: inst = 32'h10408000;
      5763: inst = 32'hc404d91;
      5764: inst = 32'h8220000;
      5765: inst = 32'h10408000;
      5766: inst = 32'hc404d92;
      5767: inst = 32'h8220000;
      5768: inst = 32'h10408000;
      5769: inst = 32'hc404d93;
      5770: inst = 32'h8220000;
      5771: inst = 32'h10408000;
      5772: inst = 32'hc404d94;
      5773: inst = 32'h8220000;
      5774: inst = 32'h10408000;
      5775: inst = 32'hc404d95;
      5776: inst = 32'h8220000;
      5777: inst = 32'h10408000;
      5778: inst = 32'hc404d96;
      5779: inst = 32'h8220000;
      5780: inst = 32'h10408000;
      5781: inst = 32'hc404d97;
      5782: inst = 32'h8220000;
      5783: inst = 32'h10408000;
      5784: inst = 32'hc404d98;
      5785: inst = 32'h8220000;
      5786: inst = 32'h10408000;
      5787: inst = 32'hc404d99;
      5788: inst = 32'h8220000;
      5789: inst = 32'h10408000;
      5790: inst = 32'hc404d9a;
      5791: inst = 32'h8220000;
      5792: inst = 32'h10408000;
      5793: inst = 32'hc404d9b;
      5794: inst = 32'h8220000;
      5795: inst = 32'h10408000;
      5796: inst = 32'hc404d9c;
      5797: inst = 32'h8220000;
      5798: inst = 32'h10408000;
      5799: inst = 32'hc404d9d;
      5800: inst = 32'h8220000;
      5801: inst = 32'h10408000;
      5802: inst = 32'hc404d9e;
      5803: inst = 32'h8220000;
      5804: inst = 32'h10408000;
      5805: inst = 32'hc404d9f;
      5806: inst = 32'h8220000;
      5807: inst = 32'h10408000;
      5808: inst = 32'hc404da0;
      5809: inst = 32'h8220000;
      5810: inst = 32'h10408000;
      5811: inst = 32'hc404da1;
      5812: inst = 32'h8220000;
      5813: inst = 32'h10408000;
      5814: inst = 32'hc404da2;
      5815: inst = 32'h8220000;
      5816: inst = 32'h10408000;
      5817: inst = 32'hc404da3;
      5818: inst = 32'h8220000;
      5819: inst = 32'h10408000;
      5820: inst = 32'hc404da4;
      5821: inst = 32'h8220000;
      5822: inst = 32'h10408000;
      5823: inst = 32'hc404da5;
      5824: inst = 32'h8220000;
      5825: inst = 32'h10408000;
      5826: inst = 32'hc404da6;
      5827: inst = 32'h8220000;
      5828: inst = 32'h10408000;
      5829: inst = 32'hc404da7;
      5830: inst = 32'h8220000;
      5831: inst = 32'h10408000;
      5832: inst = 32'hc404da8;
      5833: inst = 32'h8220000;
      5834: inst = 32'h10408000;
      5835: inst = 32'hc404da9;
      5836: inst = 32'h8220000;
      5837: inst = 32'h10408000;
      5838: inst = 32'hc404daa;
      5839: inst = 32'h8220000;
      5840: inst = 32'h10408000;
      5841: inst = 32'hc404dab;
      5842: inst = 32'h8220000;
      5843: inst = 32'h10408000;
      5844: inst = 32'hc404dac;
      5845: inst = 32'h8220000;
      5846: inst = 32'h10408000;
      5847: inst = 32'hc404dad;
      5848: inst = 32'h8220000;
      5849: inst = 32'h10408000;
      5850: inst = 32'hc404dae;
      5851: inst = 32'h8220000;
      5852: inst = 32'h10408000;
      5853: inst = 32'hc404dd7;
      5854: inst = 32'h8220000;
      5855: inst = 32'h10408000;
      5856: inst = 32'hc404dd8;
      5857: inst = 32'h8220000;
      5858: inst = 32'h10408000;
      5859: inst = 32'hc404dd9;
      5860: inst = 32'h8220000;
      5861: inst = 32'h10408000;
      5862: inst = 32'hc404dda;
      5863: inst = 32'h8220000;
      5864: inst = 32'h10408000;
      5865: inst = 32'hc404ddb;
      5866: inst = 32'h8220000;
      5867: inst = 32'h10408000;
      5868: inst = 32'hc404ddc;
      5869: inst = 32'h8220000;
      5870: inst = 32'h10408000;
      5871: inst = 32'hc404ddd;
      5872: inst = 32'h8220000;
      5873: inst = 32'h10408000;
      5874: inst = 32'hc404dde;
      5875: inst = 32'h8220000;
      5876: inst = 32'h10408000;
      5877: inst = 32'hc404ddf;
      5878: inst = 32'h8220000;
      5879: inst = 32'h10408000;
      5880: inst = 32'hc404de0;
      5881: inst = 32'h8220000;
      5882: inst = 32'h10408000;
      5883: inst = 32'hc404de1;
      5884: inst = 32'h8220000;
      5885: inst = 32'h10408000;
      5886: inst = 32'hc404de2;
      5887: inst = 32'h8220000;
      5888: inst = 32'h10408000;
      5889: inst = 32'hc404de3;
      5890: inst = 32'h8220000;
      5891: inst = 32'h10408000;
      5892: inst = 32'hc404de4;
      5893: inst = 32'h8220000;
      5894: inst = 32'h10408000;
      5895: inst = 32'hc404de5;
      5896: inst = 32'h8220000;
      5897: inst = 32'h10408000;
      5898: inst = 32'hc404de6;
      5899: inst = 32'h8220000;
      5900: inst = 32'h10408000;
      5901: inst = 32'hc404de7;
      5902: inst = 32'h8220000;
      5903: inst = 32'h10408000;
      5904: inst = 32'hc404de8;
      5905: inst = 32'h8220000;
      5906: inst = 32'h10408000;
      5907: inst = 32'hc404de9;
      5908: inst = 32'h8220000;
      5909: inst = 32'h10408000;
      5910: inst = 32'hc404dea;
      5911: inst = 32'h8220000;
      5912: inst = 32'h10408000;
      5913: inst = 32'hc404deb;
      5914: inst = 32'h8220000;
      5915: inst = 32'h10408000;
      5916: inst = 32'hc404dec;
      5917: inst = 32'h8220000;
      5918: inst = 32'h10408000;
      5919: inst = 32'hc404ded;
      5920: inst = 32'h8220000;
      5921: inst = 32'h10408000;
      5922: inst = 32'hc404dee;
      5923: inst = 32'h8220000;
      5924: inst = 32'h10408000;
      5925: inst = 32'hc404def;
      5926: inst = 32'h8220000;
      5927: inst = 32'h10408000;
      5928: inst = 32'hc404df0;
      5929: inst = 32'h8220000;
      5930: inst = 32'h10408000;
      5931: inst = 32'hc404df1;
      5932: inst = 32'h8220000;
      5933: inst = 32'h10408000;
      5934: inst = 32'hc404df2;
      5935: inst = 32'h8220000;
      5936: inst = 32'h10408000;
      5937: inst = 32'hc404df3;
      5938: inst = 32'h8220000;
      5939: inst = 32'h10408000;
      5940: inst = 32'hc404df4;
      5941: inst = 32'h8220000;
      5942: inst = 32'h10408000;
      5943: inst = 32'hc404df5;
      5944: inst = 32'h8220000;
      5945: inst = 32'h10408000;
      5946: inst = 32'hc404df6;
      5947: inst = 32'h8220000;
      5948: inst = 32'h10408000;
      5949: inst = 32'hc404df7;
      5950: inst = 32'h8220000;
      5951: inst = 32'h10408000;
      5952: inst = 32'hc404df8;
      5953: inst = 32'h8220000;
      5954: inst = 32'h10408000;
      5955: inst = 32'hc404df9;
      5956: inst = 32'h8220000;
      5957: inst = 32'h10408000;
      5958: inst = 32'hc404dfa;
      5959: inst = 32'h8220000;
      5960: inst = 32'h10408000;
      5961: inst = 32'hc404dfb;
      5962: inst = 32'h8220000;
      5963: inst = 32'h10408000;
      5964: inst = 32'hc404dfc;
      5965: inst = 32'h8220000;
      5966: inst = 32'h10408000;
      5967: inst = 32'hc404dfd;
      5968: inst = 32'h8220000;
      5969: inst = 32'h10408000;
      5970: inst = 32'hc404dfe;
      5971: inst = 32'h8220000;
      5972: inst = 32'h10408000;
      5973: inst = 32'hc404dff;
      5974: inst = 32'h8220000;
      5975: inst = 32'h10408000;
      5976: inst = 32'hc404e00;
      5977: inst = 32'h8220000;
      5978: inst = 32'h10408000;
      5979: inst = 32'hc404e01;
      5980: inst = 32'h8220000;
      5981: inst = 32'h10408000;
      5982: inst = 32'hc404e02;
      5983: inst = 32'h8220000;
      5984: inst = 32'h10408000;
      5985: inst = 32'hc404e03;
      5986: inst = 32'h8220000;
      5987: inst = 32'h10408000;
      5988: inst = 32'hc404e04;
      5989: inst = 32'h8220000;
      5990: inst = 32'h10408000;
      5991: inst = 32'hc404e05;
      5992: inst = 32'h8220000;
      5993: inst = 32'h10408000;
      5994: inst = 32'hc404e06;
      5995: inst = 32'h8220000;
      5996: inst = 32'h10408000;
      5997: inst = 32'hc404e07;
      5998: inst = 32'h8220000;
      5999: inst = 32'h10408000;
      6000: inst = 32'hc404e08;
      6001: inst = 32'h8220000;
      6002: inst = 32'h10408000;
      6003: inst = 32'hc404e09;
      6004: inst = 32'h8220000;
      6005: inst = 32'h10408000;
      6006: inst = 32'hc404e0a;
      6007: inst = 32'h8220000;
      6008: inst = 32'h10408000;
      6009: inst = 32'hc404e0b;
      6010: inst = 32'h8220000;
      6011: inst = 32'h10408000;
      6012: inst = 32'hc404e0c;
      6013: inst = 32'h8220000;
      6014: inst = 32'h10408000;
      6015: inst = 32'hc404e0d;
      6016: inst = 32'h8220000;
      6017: inst = 32'h10408000;
      6018: inst = 32'hc404e0e;
      6019: inst = 32'h8220000;
      6020: inst = 32'h10408000;
      6021: inst = 32'hc404e37;
      6022: inst = 32'h8220000;
      6023: inst = 32'h10408000;
      6024: inst = 32'hc404e38;
      6025: inst = 32'h8220000;
      6026: inst = 32'h10408000;
      6027: inst = 32'hc404e39;
      6028: inst = 32'h8220000;
      6029: inst = 32'h10408000;
      6030: inst = 32'hc404e3a;
      6031: inst = 32'h8220000;
      6032: inst = 32'h10408000;
      6033: inst = 32'hc404e3b;
      6034: inst = 32'h8220000;
      6035: inst = 32'h10408000;
      6036: inst = 32'hc404e3c;
      6037: inst = 32'h8220000;
      6038: inst = 32'h10408000;
      6039: inst = 32'hc404e3d;
      6040: inst = 32'h8220000;
      6041: inst = 32'h10408000;
      6042: inst = 32'hc404e3e;
      6043: inst = 32'h8220000;
      6044: inst = 32'h10408000;
      6045: inst = 32'hc404e3f;
      6046: inst = 32'h8220000;
      6047: inst = 32'h10408000;
      6048: inst = 32'hc404e40;
      6049: inst = 32'h8220000;
      6050: inst = 32'h10408000;
      6051: inst = 32'hc404e41;
      6052: inst = 32'h8220000;
      6053: inst = 32'h10408000;
      6054: inst = 32'hc404e42;
      6055: inst = 32'h8220000;
      6056: inst = 32'h10408000;
      6057: inst = 32'hc404e43;
      6058: inst = 32'h8220000;
      6059: inst = 32'h10408000;
      6060: inst = 32'hc404e44;
      6061: inst = 32'h8220000;
      6062: inst = 32'h10408000;
      6063: inst = 32'hc404e45;
      6064: inst = 32'h8220000;
      6065: inst = 32'h10408000;
      6066: inst = 32'hc404e46;
      6067: inst = 32'h8220000;
      6068: inst = 32'h10408000;
      6069: inst = 32'hc404e47;
      6070: inst = 32'h8220000;
      6071: inst = 32'h10408000;
      6072: inst = 32'hc404e48;
      6073: inst = 32'h8220000;
      6074: inst = 32'h10408000;
      6075: inst = 32'hc404e49;
      6076: inst = 32'h8220000;
      6077: inst = 32'h10408000;
      6078: inst = 32'hc404e4a;
      6079: inst = 32'h8220000;
      6080: inst = 32'h10408000;
      6081: inst = 32'hc404e4b;
      6082: inst = 32'h8220000;
      6083: inst = 32'h10408000;
      6084: inst = 32'hc404e4c;
      6085: inst = 32'h8220000;
      6086: inst = 32'h10408000;
      6087: inst = 32'hc404e4d;
      6088: inst = 32'h8220000;
      6089: inst = 32'h10408000;
      6090: inst = 32'hc404e4e;
      6091: inst = 32'h8220000;
      6092: inst = 32'h10408000;
      6093: inst = 32'hc404e4f;
      6094: inst = 32'h8220000;
      6095: inst = 32'h10408000;
      6096: inst = 32'hc404e50;
      6097: inst = 32'h8220000;
      6098: inst = 32'h10408000;
      6099: inst = 32'hc404e51;
      6100: inst = 32'h8220000;
      6101: inst = 32'h10408000;
      6102: inst = 32'hc404e52;
      6103: inst = 32'h8220000;
      6104: inst = 32'h10408000;
      6105: inst = 32'hc404e53;
      6106: inst = 32'h8220000;
      6107: inst = 32'h10408000;
      6108: inst = 32'hc404e54;
      6109: inst = 32'h8220000;
      6110: inst = 32'h10408000;
      6111: inst = 32'hc404e55;
      6112: inst = 32'h8220000;
      6113: inst = 32'h10408000;
      6114: inst = 32'hc404e56;
      6115: inst = 32'h8220000;
      6116: inst = 32'h10408000;
      6117: inst = 32'hc404e57;
      6118: inst = 32'h8220000;
      6119: inst = 32'h10408000;
      6120: inst = 32'hc404e58;
      6121: inst = 32'h8220000;
      6122: inst = 32'h10408000;
      6123: inst = 32'hc404e59;
      6124: inst = 32'h8220000;
      6125: inst = 32'h10408000;
      6126: inst = 32'hc404e5a;
      6127: inst = 32'h8220000;
      6128: inst = 32'h10408000;
      6129: inst = 32'hc404e5b;
      6130: inst = 32'h8220000;
      6131: inst = 32'h10408000;
      6132: inst = 32'hc404e5c;
      6133: inst = 32'h8220000;
      6134: inst = 32'h10408000;
      6135: inst = 32'hc404e5d;
      6136: inst = 32'h8220000;
      6137: inst = 32'h10408000;
      6138: inst = 32'hc404e5e;
      6139: inst = 32'h8220000;
      6140: inst = 32'h10408000;
      6141: inst = 32'hc404e5f;
      6142: inst = 32'h8220000;
      6143: inst = 32'h10408000;
      6144: inst = 32'hc404e60;
      6145: inst = 32'h8220000;
      6146: inst = 32'h10408000;
      6147: inst = 32'hc404e61;
      6148: inst = 32'h8220000;
      6149: inst = 32'h10408000;
      6150: inst = 32'hc404e62;
      6151: inst = 32'h8220000;
      6152: inst = 32'h10408000;
      6153: inst = 32'hc404e63;
      6154: inst = 32'h8220000;
      6155: inst = 32'h10408000;
      6156: inst = 32'hc404e64;
      6157: inst = 32'h8220000;
      6158: inst = 32'h10408000;
      6159: inst = 32'hc404e65;
      6160: inst = 32'h8220000;
      6161: inst = 32'h10408000;
      6162: inst = 32'hc404e66;
      6163: inst = 32'h8220000;
      6164: inst = 32'h10408000;
      6165: inst = 32'hc404e67;
      6166: inst = 32'h8220000;
      6167: inst = 32'h10408000;
      6168: inst = 32'hc404e68;
      6169: inst = 32'h8220000;
      6170: inst = 32'h10408000;
      6171: inst = 32'hc404e69;
      6172: inst = 32'h8220000;
      6173: inst = 32'h10408000;
      6174: inst = 32'hc404e6a;
      6175: inst = 32'h8220000;
      6176: inst = 32'h10408000;
      6177: inst = 32'hc404e6b;
      6178: inst = 32'h8220000;
      6179: inst = 32'h10408000;
      6180: inst = 32'hc404e6c;
      6181: inst = 32'h8220000;
      6182: inst = 32'h10408000;
      6183: inst = 32'hc404e6d;
      6184: inst = 32'h8220000;
      6185: inst = 32'h10408000;
      6186: inst = 32'hc404e6e;
      6187: inst = 32'h8220000;
      6188: inst = 32'h10408000;
      6189: inst = 32'hc404e97;
      6190: inst = 32'h8220000;
      6191: inst = 32'h10408000;
      6192: inst = 32'hc404e98;
      6193: inst = 32'h8220000;
      6194: inst = 32'h10408000;
      6195: inst = 32'hc404e99;
      6196: inst = 32'h8220000;
      6197: inst = 32'h10408000;
      6198: inst = 32'hc404e9a;
      6199: inst = 32'h8220000;
      6200: inst = 32'h10408000;
      6201: inst = 32'hc404e9b;
      6202: inst = 32'h8220000;
      6203: inst = 32'h10408000;
      6204: inst = 32'hc404e9c;
      6205: inst = 32'h8220000;
      6206: inst = 32'h10408000;
      6207: inst = 32'hc404e9d;
      6208: inst = 32'h8220000;
      6209: inst = 32'h10408000;
      6210: inst = 32'hc404e9e;
      6211: inst = 32'h8220000;
      6212: inst = 32'h10408000;
      6213: inst = 32'hc404ea8;
      6214: inst = 32'h8220000;
      6215: inst = 32'h10408000;
      6216: inst = 32'hc404ea9;
      6217: inst = 32'h8220000;
      6218: inst = 32'h10408000;
      6219: inst = 32'hc404eaa;
      6220: inst = 32'h8220000;
      6221: inst = 32'h10408000;
      6222: inst = 32'hc404eab;
      6223: inst = 32'h8220000;
      6224: inst = 32'h10408000;
      6225: inst = 32'hc404eac;
      6226: inst = 32'h8220000;
      6227: inst = 32'h10408000;
      6228: inst = 32'hc404ead;
      6229: inst = 32'h8220000;
      6230: inst = 32'h10408000;
      6231: inst = 32'hc404eae;
      6232: inst = 32'h8220000;
      6233: inst = 32'h10408000;
      6234: inst = 32'hc404eaf;
      6235: inst = 32'h8220000;
      6236: inst = 32'h10408000;
      6237: inst = 32'hc404eb0;
      6238: inst = 32'h8220000;
      6239: inst = 32'h10408000;
      6240: inst = 32'hc404eb1;
      6241: inst = 32'h8220000;
      6242: inst = 32'h10408000;
      6243: inst = 32'hc404eb2;
      6244: inst = 32'h8220000;
      6245: inst = 32'h10408000;
      6246: inst = 32'hc404eb3;
      6247: inst = 32'h8220000;
      6248: inst = 32'h10408000;
      6249: inst = 32'hc404eb4;
      6250: inst = 32'h8220000;
      6251: inst = 32'h10408000;
      6252: inst = 32'hc404eb5;
      6253: inst = 32'h8220000;
      6254: inst = 32'h10408000;
      6255: inst = 32'hc404eb6;
      6256: inst = 32'h8220000;
      6257: inst = 32'h10408000;
      6258: inst = 32'hc404eb7;
      6259: inst = 32'h8220000;
      6260: inst = 32'h10408000;
      6261: inst = 32'hc404ec1;
      6262: inst = 32'h8220000;
      6263: inst = 32'h10408000;
      6264: inst = 32'hc404ec2;
      6265: inst = 32'h8220000;
      6266: inst = 32'h10408000;
      6267: inst = 32'hc404ec3;
      6268: inst = 32'h8220000;
      6269: inst = 32'h10408000;
      6270: inst = 32'hc404ec4;
      6271: inst = 32'h8220000;
      6272: inst = 32'h10408000;
      6273: inst = 32'hc404ec5;
      6274: inst = 32'h8220000;
      6275: inst = 32'h10408000;
      6276: inst = 32'hc404ec6;
      6277: inst = 32'h8220000;
      6278: inst = 32'h10408000;
      6279: inst = 32'hc404ec7;
      6280: inst = 32'h8220000;
      6281: inst = 32'h10408000;
      6282: inst = 32'hc404ec8;
      6283: inst = 32'h8220000;
      6284: inst = 32'h10408000;
      6285: inst = 32'hc404ec9;
      6286: inst = 32'h8220000;
      6287: inst = 32'h10408000;
      6288: inst = 32'hc404eca;
      6289: inst = 32'h8220000;
      6290: inst = 32'h10408000;
      6291: inst = 32'hc404ecb;
      6292: inst = 32'h8220000;
      6293: inst = 32'h10408000;
      6294: inst = 32'hc404ecc;
      6295: inst = 32'h8220000;
      6296: inst = 32'h10408000;
      6297: inst = 32'hc404ecd;
      6298: inst = 32'h8220000;
      6299: inst = 32'h10408000;
      6300: inst = 32'hc404ece;
      6301: inst = 32'h8220000;
      6302: inst = 32'h10408000;
      6303: inst = 32'hc404ef7;
      6304: inst = 32'h8220000;
      6305: inst = 32'h10408000;
      6306: inst = 32'hc404ef8;
      6307: inst = 32'h8220000;
      6308: inst = 32'h10408000;
      6309: inst = 32'hc404ef9;
      6310: inst = 32'h8220000;
      6311: inst = 32'h10408000;
      6312: inst = 32'hc404efa;
      6313: inst = 32'h8220000;
      6314: inst = 32'h10408000;
      6315: inst = 32'hc404efb;
      6316: inst = 32'h8220000;
      6317: inst = 32'h10408000;
      6318: inst = 32'hc404efc;
      6319: inst = 32'h8220000;
      6320: inst = 32'h10408000;
      6321: inst = 32'hc404efd;
      6322: inst = 32'h8220000;
      6323: inst = 32'h10408000;
      6324: inst = 32'hc404efe;
      6325: inst = 32'h8220000;
      6326: inst = 32'h10408000;
      6327: inst = 32'hc404f08;
      6328: inst = 32'h8220000;
      6329: inst = 32'h10408000;
      6330: inst = 32'hc404f09;
      6331: inst = 32'h8220000;
      6332: inst = 32'h10408000;
      6333: inst = 32'hc404f0a;
      6334: inst = 32'h8220000;
      6335: inst = 32'h10408000;
      6336: inst = 32'hc404f0b;
      6337: inst = 32'h8220000;
      6338: inst = 32'h10408000;
      6339: inst = 32'hc404f0c;
      6340: inst = 32'h8220000;
      6341: inst = 32'h10408000;
      6342: inst = 32'hc404f0d;
      6343: inst = 32'h8220000;
      6344: inst = 32'h10408000;
      6345: inst = 32'hc404f0e;
      6346: inst = 32'h8220000;
      6347: inst = 32'h10408000;
      6348: inst = 32'hc404f0f;
      6349: inst = 32'h8220000;
      6350: inst = 32'h10408000;
      6351: inst = 32'hc404f10;
      6352: inst = 32'h8220000;
      6353: inst = 32'h10408000;
      6354: inst = 32'hc404f11;
      6355: inst = 32'h8220000;
      6356: inst = 32'h10408000;
      6357: inst = 32'hc404f12;
      6358: inst = 32'h8220000;
      6359: inst = 32'h10408000;
      6360: inst = 32'hc404f13;
      6361: inst = 32'h8220000;
      6362: inst = 32'h10408000;
      6363: inst = 32'hc404f14;
      6364: inst = 32'h8220000;
      6365: inst = 32'h10408000;
      6366: inst = 32'hc404f15;
      6367: inst = 32'h8220000;
      6368: inst = 32'h10408000;
      6369: inst = 32'hc404f16;
      6370: inst = 32'h8220000;
      6371: inst = 32'h10408000;
      6372: inst = 32'hc404f17;
      6373: inst = 32'h8220000;
      6374: inst = 32'h10408000;
      6375: inst = 32'hc404f21;
      6376: inst = 32'h8220000;
      6377: inst = 32'h10408000;
      6378: inst = 32'hc404f22;
      6379: inst = 32'h8220000;
      6380: inst = 32'h10408000;
      6381: inst = 32'hc404f23;
      6382: inst = 32'h8220000;
      6383: inst = 32'h10408000;
      6384: inst = 32'hc404f24;
      6385: inst = 32'h8220000;
      6386: inst = 32'h10408000;
      6387: inst = 32'hc404f25;
      6388: inst = 32'h8220000;
      6389: inst = 32'h10408000;
      6390: inst = 32'hc404f26;
      6391: inst = 32'h8220000;
      6392: inst = 32'h10408000;
      6393: inst = 32'hc404f27;
      6394: inst = 32'h8220000;
      6395: inst = 32'h10408000;
      6396: inst = 32'hc404f28;
      6397: inst = 32'h8220000;
      6398: inst = 32'h10408000;
      6399: inst = 32'hc404f29;
      6400: inst = 32'h8220000;
      6401: inst = 32'h10408000;
      6402: inst = 32'hc404f2a;
      6403: inst = 32'h8220000;
      6404: inst = 32'h10408000;
      6405: inst = 32'hc404f2b;
      6406: inst = 32'h8220000;
      6407: inst = 32'h10408000;
      6408: inst = 32'hc404f2c;
      6409: inst = 32'h8220000;
      6410: inst = 32'h10408000;
      6411: inst = 32'hc404f2d;
      6412: inst = 32'h8220000;
      6413: inst = 32'h10408000;
      6414: inst = 32'hc404f2e;
      6415: inst = 32'h8220000;
      6416: inst = 32'h10408000;
      6417: inst = 32'hc404f57;
      6418: inst = 32'h8220000;
      6419: inst = 32'h10408000;
      6420: inst = 32'hc404f58;
      6421: inst = 32'h8220000;
      6422: inst = 32'h10408000;
      6423: inst = 32'hc404f59;
      6424: inst = 32'h8220000;
      6425: inst = 32'h10408000;
      6426: inst = 32'hc404f5a;
      6427: inst = 32'h8220000;
      6428: inst = 32'h10408000;
      6429: inst = 32'hc404f5b;
      6430: inst = 32'h8220000;
      6431: inst = 32'h10408000;
      6432: inst = 32'hc404f5c;
      6433: inst = 32'h8220000;
      6434: inst = 32'h10408000;
      6435: inst = 32'hc404f5d;
      6436: inst = 32'h8220000;
      6437: inst = 32'h10408000;
      6438: inst = 32'hc404f5e;
      6439: inst = 32'h8220000;
      6440: inst = 32'h10408000;
      6441: inst = 32'hc404f68;
      6442: inst = 32'h8220000;
      6443: inst = 32'h10408000;
      6444: inst = 32'hc404f69;
      6445: inst = 32'h8220000;
      6446: inst = 32'h10408000;
      6447: inst = 32'hc404f6a;
      6448: inst = 32'h8220000;
      6449: inst = 32'h10408000;
      6450: inst = 32'hc404f6b;
      6451: inst = 32'h8220000;
      6452: inst = 32'h10408000;
      6453: inst = 32'hc404f6c;
      6454: inst = 32'h8220000;
      6455: inst = 32'h10408000;
      6456: inst = 32'hc404f6d;
      6457: inst = 32'h8220000;
      6458: inst = 32'h10408000;
      6459: inst = 32'hc404f6e;
      6460: inst = 32'h8220000;
      6461: inst = 32'h10408000;
      6462: inst = 32'hc404f6f;
      6463: inst = 32'h8220000;
      6464: inst = 32'h10408000;
      6465: inst = 32'hc404f70;
      6466: inst = 32'h8220000;
      6467: inst = 32'h10408000;
      6468: inst = 32'hc404f71;
      6469: inst = 32'h8220000;
      6470: inst = 32'h10408000;
      6471: inst = 32'hc404f72;
      6472: inst = 32'h8220000;
      6473: inst = 32'h10408000;
      6474: inst = 32'hc404f73;
      6475: inst = 32'h8220000;
      6476: inst = 32'h10408000;
      6477: inst = 32'hc404f74;
      6478: inst = 32'h8220000;
      6479: inst = 32'h10408000;
      6480: inst = 32'hc404f75;
      6481: inst = 32'h8220000;
      6482: inst = 32'h10408000;
      6483: inst = 32'hc404f76;
      6484: inst = 32'h8220000;
      6485: inst = 32'h10408000;
      6486: inst = 32'hc404f77;
      6487: inst = 32'h8220000;
      6488: inst = 32'h10408000;
      6489: inst = 32'hc404f81;
      6490: inst = 32'h8220000;
      6491: inst = 32'h10408000;
      6492: inst = 32'hc404f82;
      6493: inst = 32'h8220000;
      6494: inst = 32'h10408000;
      6495: inst = 32'hc404f83;
      6496: inst = 32'h8220000;
      6497: inst = 32'h10408000;
      6498: inst = 32'hc404f84;
      6499: inst = 32'h8220000;
      6500: inst = 32'h10408000;
      6501: inst = 32'hc404f85;
      6502: inst = 32'h8220000;
      6503: inst = 32'h10408000;
      6504: inst = 32'hc404f86;
      6505: inst = 32'h8220000;
      6506: inst = 32'h10408000;
      6507: inst = 32'hc404f87;
      6508: inst = 32'h8220000;
      6509: inst = 32'h10408000;
      6510: inst = 32'hc404f88;
      6511: inst = 32'h8220000;
      6512: inst = 32'h10408000;
      6513: inst = 32'hc404f89;
      6514: inst = 32'h8220000;
      6515: inst = 32'h10408000;
      6516: inst = 32'hc404f8a;
      6517: inst = 32'h8220000;
      6518: inst = 32'h10408000;
      6519: inst = 32'hc404f8b;
      6520: inst = 32'h8220000;
      6521: inst = 32'h10408000;
      6522: inst = 32'hc404f8c;
      6523: inst = 32'h8220000;
      6524: inst = 32'h10408000;
      6525: inst = 32'hc404f8d;
      6526: inst = 32'h8220000;
      6527: inst = 32'h10408000;
      6528: inst = 32'hc404f8e;
      6529: inst = 32'h8220000;
      6530: inst = 32'h10408000;
      6531: inst = 32'hc404fb7;
      6532: inst = 32'h8220000;
      6533: inst = 32'h10408000;
      6534: inst = 32'hc404fb8;
      6535: inst = 32'h8220000;
      6536: inst = 32'h10408000;
      6537: inst = 32'hc404fb9;
      6538: inst = 32'h8220000;
      6539: inst = 32'h10408000;
      6540: inst = 32'hc404fba;
      6541: inst = 32'h8220000;
      6542: inst = 32'h10408000;
      6543: inst = 32'hc404fbb;
      6544: inst = 32'h8220000;
      6545: inst = 32'h10408000;
      6546: inst = 32'hc404fbc;
      6547: inst = 32'h8220000;
      6548: inst = 32'h10408000;
      6549: inst = 32'hc404fbd;
      6550: inst = 32'h8220000;
      6551: inst = 32'h10408000;
      6552: inst = 32'hc404fbe;
      6553: inst = 32'h8220000;
      6554: inst = 32'h10408000;
      6555: inst = 32'hc404fc8;
      6556: inst = 32'h8220000;
      6557: inst = 32'h10408000;
      6558: inst = 32'hc404fc9;
      6559: inst = 32'h8220000;
      6560: inst = 32'h10408000;
      6561: inst = 32'hc404fca;
      6562: inst = 32'h8220000;
      6563: inst = 32'h10408000;
      6564: inst = 32'hc404fcb;
      6565: inst = 32'h8220000;
      6566: inst = 32'h10408000;
      6567: inst = 32'hc404fcc;
      6568: inst = 32'h8220000;
      6569: inst = 32'h10408000;
      6570: inst = 32'hc404fcd;
      6571: inst = 32'h8220000;
      6572: inst = 32'h10408000;
      6573: inst = 32'hc404fce;
      6574: inst = 32'h8220000;
      6575: inst = 32'h10408000;
      6576: inst = 32'hc404fcf;
      6577: inst = 32'h8220000;
      6578: inst = 32'h10408000;
      6579: inst = 32'hc404fd0;
      6580: inst = 32'h8220000;
      6581: inst = 32'h10408000;
      6582: inst = 32'hc404fd1;
      6583: inst = 32'h8220000;
      6584: inst = 32'h10408000;
      6585: inst = 32'hc404fd2;
      6586: inst = 32'h8220000;
      6587: inst = 32'h10408000;
      6588: inst = 32'hc404fd3;
      6589: inst = 32'h8220000;
      6590: inst = 32'h10408000;
      6591: inst = 32'hc404fd4;
      6592: inst = 32'h8220000;
      6593: inst = 32'h10408000;
      6594: inst = 32'hc404fd5;
      6595: inst = 32'h8220000;
      6596: inst = 32'h10408000;
      6597: inst = 32'hc404fd6;
      6598: inst = 32'h8220000;
      6599: inst = 32'h10408000;
      6600: inst = 32'hc404fd7;
      6601: inst = 32'h8220000;
      6602: inst = 32'h10408000;
      6603: inst = 32'hc404fe1;
      6604: inst = 32'h8220000;
      6605: inst = 32'h10408000;
      6606: inst = 32'hc404fe2;
      6607: inst = 32'h8220000;
      6608: inst = 32'h10408000;
      6609: inst = 32'hc404fe3;
      6610: inst = 32'h8220000;
      6611: inst = 32'h10408000;
      6612: inst = 32'hc404fe4;
      6613: inst = 32'h8220000;
      6614: inst = 32'h10408000;
      6615: inst = 32'hc404fe5;
      6616: inst = 32'h8220000;
      6617: inst = 32'h10408000;
      6618: inst = 32'hc404fe6;
      6619: inst = 32'h8220000;
      6620: inst = 32'h10408000;
      6621: inst = 32'hc404fe7;
      6622: inst = 32'h8220000;
      6623: inst = 32'h10408000;
      6624: inst = 32'hc404fe8;
      6625: inst = 32'h8220000;
      6626: inst = 32'h10408000;
      6627: inst = 32'hc404fe9;
      6628: inst = 32'h8220000;
      6629: inst = 32'h10408000;
      6630: inst = 32'hc404fea;
      6631: inst = 32'h8220000;
      6632: inst = 32'h10408000;
      6633: inst = 32'hc404feb;
      6634: inst = 32'h8220000;
      6635: inst = 32'h10408000;
      6636: inst = 32'hc404fec;
      6637: inst = 32'h8220000;
      6638: inst = 32'h10408000;
      6639: inst = 32'hc404fed;
      6640: inst = 32'h8220000;
      6641: inst = 32'h10408000;
      6642: inst = 32'hc404fee;
      6643: inst = 32'h8220000;
      6644: inst = 32'h10408000;
      6645: inst = 32'hc405017;
      6646: inst = 32'h8220000;
      6647: inst = 32'h10408000;
      6648: inst = 32'hc405018;
      6649: inst = 32'h8220000;
      6650: inst = 32'h10408000;
      6651: inst = 32'hc405019;
      6652: inst = 32'h8220000;
      6653: inst = 32'h10408000;
      6654: inst = 32'hc40501a;
      6655: inst = 32'h8220000;
      6656: inst = 32'h10408000;
      6657: inst = 32'hc40501b;
      6658: inst = 32'h8220000;
      6659: inst = 32'h10408000;
      6660: inst = 32'hc40501c;
      6661: inst = 32'h8220000;
      6662: inst = 32'h10408000;
      6663: inst = 32'hc40501d;
      6664: inst = 32'h8220000;
      6665: inst = 32'h10408000;
      6666: inst = 32'hc40501e;
      6667: inst = 32'h8220000;
      6668: inst = 32'h10408000;
      6669: inst = 32'hc405028;
      6670: inst = 32'h8220000;
      6671: inst = 32'h10408000;
      6672: inst = 32'hc405029;
      6673: inst = 32'h8220000;
      6674: inst = 32'h10408000;
      6675: inst = 32'hc40502a;
      6676: inst = 32'h8220000;
      6677: inst = 32'h10408000;
      6678: inst = 32'hc40502b;
      6679: inst = 32'h8220000;
      6680: inst = 32'h10408000;
      6681: inst = 32'hc40502c;
      6682: inst = 32'h8220000;
      6683: inst = 32'h10408000;
      6684: inst = 32'hc40502d;
      6685: inst = 32'h8220000;
      6686: inst = 32'h10408000;
      6687: inst = 32'hc40502e;
      6688: inst = 32'h8220000;
      6689: inst = 32'h10408000;
      6690: inst = 32'hc40502f;
      6691: inst = 32'h8220000;
      6692: inst = 32'h10408000;
      6693: inst = 32'hc405030;
      6694: inst = 32'h8220000;
      6695: inst = 32'h10408000;
      6696: inst = 32'hc405031;
      6697: inst = 32'h8220000;
      6698: inst = 32'h10408000;
      6699: inst = 32'hc405032;
      6700: inst = 32'h8220000;
      6701: inst = 32'h10408000;
      6702: inst = 32'hc405033;
      6703: inst = 32'h8220000;
      6704: inst = 32'h10408000;
      6705: inst = 32'hc405034;
      6706: inst = 32'h8220000;
      6707: inst = 32'h10408000;
      6708: inst = 32'hc405035;
      6709: inst = 32'h8220000;
      6710: inst = 32'h10408000;
      6711: inst = 32'hc405036;
      6712: inst = 32'h8220000;
      6713: inst = 32'h10408000;
      6714: inst = 32'hc405037;
      6715: inst = 32'h8220000;
      6716: inst = 32'h10408000;
      6717: inst = 32'hc405041;
      6718: inst = 32'h8220000;
      6719: inst = 32'h10408000;
      6720: inst = 32'hc405042;
      6721: inst = 32'h8220000;
      6722: inst = 32'h10408000;
      6723: inst = 32'hc405043;
      6724: inst = 32'h8220000;
      6725: inst = 32'h10408000;
      6726: inst = 32'hc405044;
      6727: inst = 32'h8220000;
      6728: inst = 32'h10408000;
      6729: inst = 32'hc405045;
      6730: inst = 32'h8220000;
      6731: inst = 32'h10408000;
      6732: inst = 32'hc405046;
      6733: inst = 32'h8220000;
      6734: inst = 32'h10408000;
      6735: inst = 32'hc405047;
      6736: inst = 32'h8220000;
      6737: inst = 32'h10408000;
      6738: inst = 32'hc405048;
      6739: inst = 32'h8220000;
      6740: inst = 32'h10408000;
      6741: inst = 32'hc405049;
      6742: inst = 32'h8220000;
      6743: inst = 32'h10408000;
      6744: inst = 32'hc40504a;
      6745: inst = 32'h8220000;
      6746: inst = 32'h10408000;
      6747: inst = 32'hc40504b;
      6748: inst = 32'h8220000;
      6749: inst = 32'h10408000;
      6750: inst = 32'hc40504c;
      6751: inst = 32'h8220000;
      6752: inst = 32'h10408000;
      6753: inst = 32'hc40504d;
      6754: inst = 32'h8220000;
      6755: inst = 32'h10408000;
      6756: inst = 32'hc40504e;
      6757: inst = 32'h8220000;
      6758: inst = 32'h10408000;
      6759: inst = 32'hc405077;
      6760: inst = 32'h8220000;
      6761: inst = 32'h10408000;
      6762: inst = 32'hc405078;
      6763: inst = 32'h8220000;
      6764: inst = 32'h10408000;
      6765: inst = 32'hc405079;
      6766: inst = 32'h8220000;
      6767: inst = 32'h10408000;
      6768: inst = 32'hc40507a;
      6769: inst = 32'h8220000;
      6770: inst = 32'h10408000;
      6771: inst = 32'hc40507b;
      6772: inst = 32'h8220000;
      6773: inst = 32'h10408000;
      6774: inst = 32'hc40507c;
      6775: inst = 32'h8220000;
      6776: inst = 32'h10408000;
      6777: inst = 32'hc40507d;
      6778: inst = 32'h8220000;
      6779: inst = 32'h10408000;
      6780: inst = 32'hc40507e;
      6781: inst = 32'h8220000;
      6782: inst = 32'h10408000;
      6783: inst = 32'hc405088;
      6784: inst = 32'h8220000;
      6785: inst = 32'h10408000;
      6786: inst = 32'hc405089;
      6787: inst = 32'h8220000;
      6788: inst = 32'h10408000;
      6789: inst = 32'hc40508a;
      6790: inst = 32'h8220000;
      6791: inst = 32'h10408000;
      6792: inst = 32'hc40508b;
      6793: inst = 32'h8220000;
      6794: inst = 32'h10408000;
      6795: inst = 32'hc40508c;
      6796: inst = 32'h8220000;
      6797: inst = 32'h10408000;
      6798: inst = 32'hc40508d;
      6799: inst = 32'h8220000;
      6800: inst = 32'h10408000;
      6801: inst = 32'hc40508e;
      6802: inst = 32'h8220000;
      6803: inst = 32'h10408000;
      6804: inst = 32'hc40508f;
      6805: inst = 32'h8220000;
      6806: inst = 32'h10408000;
      6807: inst = 32'hc405090;
      6808: inst = 32'h8220000;
      6809: inst = 32'h10408000;
      6810: inst = 32'hc405091;
      6811: inst = 32'h8220000;
      6812: inst = 32'h10408000;
      6813: inst = 32'hc405092;
      6814: inst = 32'h8220000;
      6815: inst = 32'h10408000;
      6816: inst = 32'hc405093;
      6817: inst = 32'h8220000;
      6818: inst = 32'h10408000;
      6819: inst = 32'hc405094;
      6820: inst = 32'h8220000;
      6821: inst = 32'h10408000;
      6822: inst = 32'hc405095;
      6823: inst = 32'h8220000;
      6824: inst = 32'h10408000;
      6825: inst = 32'hc405096;
      6826: inst = 32'h8220000;
      6827: inst = 32'h10408000;
      6828: inst = 32'hc405097;
      6829: inst = 32'h8220000;
      6830: inst = 32'h10408000;
      6831: inst = 32'hc4050a1;
      6832: inst = 32'h8220000;
      6833: inst = 32'h10408000;
      6834: inst = 32'hc4050a2;
      6835: inst = 32'h8220000;
      6836: inst = 32'h10408000;
      6837: inst = 32'hc4050a3;
      6838: inst = 32'h8220000;
      6839: inst = 32'h10408000;
      6840: inst = 32'hc4050a4;
      6841: inst = 32'h8220000;
      6842: inst = 32'h10408000;
      6843: inst = 32'hc4050a5;
      6844: inst = 32'h8220000;
      6845: inst = 32'h10408000;
      6846: inst = 32'hc4050a6;
      6847: inst = 32'h8220000;
      6848: inst = 32'h10408000;
      6849: inst = 32'hc4050a7;
      6850: inst = 32'h8220000;
      6851: inst = 32'h10408000;
      6852: inst = 32'hc4050a8;
      6853: inst = 32'h8220000;
      6854: inst = 32'h10408000;
      6855: inst = 32'hc4050a9;
      6856: inst = 32'h8220000;
      6857: inst = 32'h10408000;
      6858: inst = 32'hc4050aa;
      6859: inst = 32'h8220000;
      6860: inst = 32'h10408000;
      6861: inst = 32'hc4050ab;
      6862: inst = 32'h8220000;
      6863: inst = 32'h10408000;
      6864: inst = 32'hc4050ac;
      6865: inst = 32'h8220000;
      6866: inst = 32'h10408000;
      6867: inst = 32'hc4050ad;
      6868: inst = 32'h8220000;
      6869: inst = 32'h10408000;
      6870: inst = 32'hc4050ae;
      6871: inst = 32'h8220000;
      6872: inst = 32'h10408000;
      6873: inst = 32'hc4050d7;
      6874: inst = 32'h8220000;
      6875: inst = 32'h10408000;
      6876: inst = 32'hc4050d8;
      6877: inst = 32'h8220000;
      6878: inst = 32'h10408000;
      6879: inst = 32'hc4050d9;
      6880: inst = 32'h8220000;
      6881: inst = 32'h10408000;
      6882: inst = 32'hc4050da;
      6883: inst = 32'h8220000;
      6884: inst = 32'h10408000;
      6885: inst = 32'hc4050db;
      6886: inst = 32'h8220000;
      6887: inst = 32'h10408000;
      6888: inst = 32'hc4050dc;
      6889: inst = 32'h8220000;
      6890: inst = 32'h10408000;
      6891: inst = 32'hc4050dd;
      6892: inst = 32'h8220000;
      6893: inst = 32'h10408000;
      6894: inst = 32'hc4050de;
      6895: inst = 32'h8220000;
      6896: inst = 32'h10408000;
      6897: inst = 32'hc4050e8;
      6898: inst = 32'h8220000;
      6899: inst = 32'h10408000;
      6900: inst = 32'hc4050e9;
      6901: inst = 32'h8220000;
      6902: inst = 32'h10408000;
      6903: inst = 32'hc4050ea;
      6904: inst = 32'h8220000;
      6905: inst = 32'h10408000;
      6906: inst = 32'hc4050eb;
      6907: inst = 32'h8220000;
      6908: inst = 32'h10408000;
      6909: inst = 32'hc4050ec;
      6910: inst = 32'h8220000;
      6911: inst = 32'h10408000;
      6912: inst = 32'hc4050ed;
      6913: inst = 32'h8220000;
      6914: inst = 32'h10408000;
      6915: inst = 32'hc4050ee;
      6916: inst = 32'h8220000;
      6917: inst = 32'h10408000;
      6918: inst = 32'hc4050ef;
      6919: inst = 32'h8220000;
      6920: inst = 32'h10408000;
      6921: inst = 32'hc4050f0;
      6922: inst = 32'h8220000;
      6923: inst = 32'h10408000;
      6924: inst = 32'hc4050f1;
      6925: inst = 32'h8220000;
      6926: inst = 32'h10408000;
      6927: inst = 32'hc4050f2;
      6928: inst = 32'h8220000;
      6929: inst = 32'h10408000;
      6930: inst = 32'hc4050f3;
      6931: inst = 32'h8220000;
      6932: inst = 32'h10408000;
      6933: inst = 32'hc4050f4;
      6934: inst = 32'h8220000;
      6935: inst = 32'h10408000;
      6936: inst = 32'hc4050f5;
      6937: inst = 32'h8220000;
      6938: inst = 32'h10408000;
      6939: inst = 32'hc4050f6;
      6940: inst = 32'h8220000;
      6941: inst = 32'h10408000;
      6942: inst = 32'hc4050f7;
      6943: inst = 32'h8220000;
      6944: inst = 32'h10408000;
      6945: inst = 32'hc405101;
      6946: inst = 32'h8220000;
      6947: inst = 32'h10408000;
      6948: inst = 32'hc405102;
      6949: inst = 32'h8220000;
      6950: inst = 32'h10408000;
      6951: inst = 32'hc405103;
      6952: inst = 32'h8220000;
      6953: inst = 32'h10408000;
      6954: inst = 32'hc405104;
      6955: inst = 32'h8220000;
      6956: inst = 32'h10408000;
      6957: inst = 32'hc405105;
      6958: inst = 32'h8220000;
      6959: inst = 32'h10408000;
      6960: inst = 32'hc405106;
      6961: inst = 32'h8220000;
      6962: inst = 32'h10408000;
      6963: inst = 32'hc405107;
      6964: inst = 32'h8220000;
      6965: inst = 32'h10408000;
      6966: inst = 32'hc405108;
      6967: inst = 32'h8220000;
      6968: inst = 32'h10408000;
      6969: inst = 32'hc405109;
      6970: inst = 32'h8220000;
      6971: inst = 32'h10408000;
      6972: inst = 32'hc40510a;
      6973: inst = 32'h8220000;
      6974: inst = 32'h10408000;
      6975: inst = 32'hc40510b;
      6976: inst = 32'h8220000;
      6977: inst = 32'h10408000;
      6978: inst = 32'hc40510c;
      6979: inst = 32'h8220000;
      6980: inst = 32'h10408000;
      6981: inst = 32'hc40510d;
      6982: inst = 32'h8220000;
      6983: inst = 32'h10408000;
      6984: inst = 32'hc40510e;
      6985: inst = 32'h8220000;
      6986: inst = 32'h10408000;
      6987: inst = 32'hc405137;
      6988: inst = 32'h8220000;
      6989: inst = 32'h10408000;
      6990: inst = 32'hc405138;
      6991: inst = 32'h8220000;
      6992: inst = 32'h10408000;
      6993: inst = 32'hc405139;
      6994: inst = 32'h8220000;
      6995: inst = 32'h10408000;
      6996: inst = 32'hc40513a;
      6997: inst = 32'h8220000;
      6998: inst = 32'h10408000;
      6999: inst = 32'hc40513b;
      7000: inst = 32'h8220000;
      7001: inst = 32'h10408000;
      7002: inst = 32'hc40513c;
      7003: inst = 32'h8220000;
      7004: inst = 32'h10408000;
      7005: inst = 32'hc40513d;
      7006: inst = 32'h8220000;
      7007: inst = 32'h10408000;
      7008: inst = 32'hc40513e;
      7009: inst = 32'h8220000;
      7010: inst = 32'h10408000;
      7011: inst = 32'hc405148;
      7012: inst = 32'h8220000;
      7013: inst = 32'h10408000;
      7014: inst = 32'hc405149;
      7015: inst = 32'h8220000;
      7016: inst = 32'h10408000;
      7017: inst = 32'hc40514a;
      7018: inst = 32'h8220000;
      7019: inst = 32'h10408000;
      7020: inst = 32'hc40514b;
      7021: inst = 32'h8220000;
      7022: inst = 32'h10408000;
      7023: inst = 32'hc40514c;
      7024: inst = 32'h8220000;
      7025: inst = 32'h10408000;
      7026: inst = 32'hc40514d;
      7027: inst = 32'h8220000;
      7028: inst = 32'h10408000;
      7029: inst = 32'hc40514e;
      7030: inst = 32'h8220000;
      7031: inst = 32'h10408000;
      7032: inst = 32'hc40514f;
      7033: inst = 32'h8220000;
      7034: inst = 32'h10408000;
      7035: inst = 32'hc405150;
      7036: inst = 32'h8220000;
      7037: inst = 32'h10408000;
      7038: inst = 32'hc405151;
      7039: inst = 32'h8220000;
      7040: inst = 32'h10408000;
      7041: inst = 32'hc405152;
      7042: inst = 32'h8220000;
      7043: inst = 32'h10408000;
      7044: inst = 32'hc405153;
      7045: inst = 32'h8220000;
      7046: inst = 32'h10408000;
      7047: inst = 32'hc405154;
      7048: inst = 32'h8220000;
      7049: inst = 32'h10408000;
      7050: inst = 32'hc405155;
      7051: inst = 32'h8220000;
      7052: inst = 32'h10408000;
      7053: inst = 32'hc405156;
      7054: inst = 32'h8220000;
      7055: inst = 32'h10408000;
      7056: inst = 32'hc405157;
      7057: inst = 32'h8220000;
      7058: inst = 32'h10408000;
      7059: inst = 32'hc405161;
      7060: inst = 32'h8220000;
      7061: inst = 32'h10408000;
      7062: inst = 32'hc405162;
      7063: inst = 32'h8220000;
      7064: inst = 32'h10408000;
      7065: inst = 32'hc405163;
      7066: inst = 32'h8220000;
      7067: inst = 32'h10408000;
      7068: inst = 32'hc405164;
      7069: inst = 32'h8220000;
      7070: inst = 32'h10408000;
      7071: inst = 32'hc405165;
      7072: inst = 32'h8220000;
      7073: inst = 32'h10408000;
      7074: inst = 32'hc405166;
      7075: inst = 32'h8220000;
      7076: inst = 32'h10408000;
      7077: inst = 32'hc405167;
      7078: inst = 32'h8220000;
      7079: inst = 32'h10408000;
      7080: inst = 32'hc405168;
      7081: inst = 32'h8220000;
      7082: inst = 32'h10408000;
      7083: inst = 32'hc405169;
      7084: inst = 32'h8220000;
      7085: inst = 32'h10408000;
      7086: inst = 32'hc40516a;
      7087: inst = 32'h8220000;
      7088: inst = 32'h10408000;
      7089: inst = 32'hc40516b;
      7090: inst = 32'h8220000;
      7091: inst = 32'h10408000;
      7092: inst = 32'hc40516c;
      7093: inst = 32'h8220000;
      7094: inst = 32'h10408000;
      7095: inst = 32'hc40516d;
      7096: inst = 32'h8220000;
      7097: inst = 32'h10408000;
      7098: inst = 32'hc40516e;
      7099: inst = 32'h8220000;
      7100: inst = 32'h10408000;
      7101: inst = 32'hc405197;
      7102: inst = 32'h8220000;
      7103: inst = 32'h10408000;
      7104: inst = 32'hc405198;
      7105: inst = 32'h8220000;
      7106: inst = 32'h10408000;
      7107: inst = 32'hc405199;
      7108: inst = 32'h8220000;
      7109: inst = 32'h10408000;
      7110: inst = 32'hc40519a;
      7111: inst = 32'h8220000;
      7112: inst = 32'h10408000;
      7113: inst = 32'hc40519b;
      7114: inst = 32'h8220000;
      7115: inst = 32'h10408000;
      7116: inst = 32'hc40519c;
      7117: inst = 32'h8220000;
      7118: inst = 32'h10408000;
      7119: inst = 32'hc40519d;
      7120: inst = 32'h8220000;
      7121: inst = 32'h10408000;
      7122: inst = 32'hc4051aa;
      7123: inst = 32'h8220000;
      7124: inst = 32'h10408000;
      7125: inst = 32'hc4051ab;
      7126: inst = 32'h8220000;
      7127: inst = 32'h10408000;
      7128: inst = 32'hc4051ac;
      7129: inst = 32'h8220000;
      7130: inst = 32'h10408000;
      7131: inst = 32'hc4051ad;
      7132: inst = 32'h8220000;
      7133: inst = 32'h10408000;
      7134: inst = 32'hc4051ae;
      7135: inst = 32'h8220000;
      7136: inst = 32'h10408000;
      7137: inst = 32'hc4051af;
      7138: inst = 32'h8220000;
      7139: inst = 32'h10408000;
      7140: inst = 32'hc4051b0;
      7141: inst = 32'h8220000;
      7142: inst = 32'h10408000;
      7143: inst = 32'hc4051b1;
      7144: inst = 32'h8220000;
      7145: inst = 32'h10408000;
      7146: inst = 32'hc4051b2;
      7147: inst = 32'h8220000;
      7148: inst = 32'h10408000;
      7149: inst = 32'hc4051b3;
      7150: inst = 32'h8220000;
      7151: inst = 32'h10408000;
      7152: inst = 32'hc4051b4;
      7153: inst = 32'h8220000;
      7154: inst = 32'h10408000;
      7155: inst = 32'hc4051b5;
      7156: inst = 32'h8220000;
      7157: inst = 32'h10408000;
      7158: inst = 32'hc4051c2;
      7159: inst = 32'h8220000;
      7160: inst = 32'h10408000;
      7161: inst = 32'hc4051c3;
      7162: inst = 32'h8220000;
      7163: inst = 32'h10408000;
      7164: inst = 32'hc4051c4;
      7165: inst = 32'h8220000;
      7166: inst = 32'h10408000;
      7167: inst = 32'hc4051c5;
      7168: inst = 32'h8220000;
      7169: inst = 32'h10408000;
      7170: inst = 32'hc4051c6;
      7171: inst = 32'h8220000;
      7172: inst = 32'h10408000;
      7173: inst = 32'hc4051c7;
      7174: inst = 32'h8220000;
      7175: inst = 32'h10408000;
      7176: inst = 32'hc4051c8;
      7177: inst = 32'h8220000;
      7178: inst = 32'h10408000;
      7179: inst = 32'hc4051c9;
      7180: inst = 32'h8220000;
      7181: inst = 32'h10408000;
      7182: inst = 32'hc4051ca;
      7183: inst = 32'h8220000;
      7184: inst = 32'h10408000;
      7185: inst = 32'hc4051cb;
      7186: inst = 32'h8220000;
      7187: inst = 32'h10408000;
      7188: inst = 32'hc4051cc;
      7189: inst = 32'h8220000;
      7190: inst = 32'h10408000;
      7191: inst = 32'hc4051cd;
      7192: inst = 32'h8220000;
      7193: inst = 32'h10408000;
      7194: inst = 32'hc4051ce;
      7195: inst = 32'h8220000;
      7196: inst = 32'h10408000;
      7197: inst = 32'hc4051f7;
      7198: inst = 32'h8220000;
      7199: inst = 32'h10408000;
      7200: inst = 32'hc4051f8;
      7201: inst = 32'h8220000;
      7202: inst = 32'h10408000;
      7203: inst = 32'hc4051f9;
      7204: inst = 32'h8220000;
      7205: inst = 32'h10408000;
      7206: inst = 32'hc4051fa;
      7207: inst = 32'h8220000;
      7208: inst = 32'h10408000;
      7209: inst = 32'hc4051fb;
      7210: inst = 32'h8220000;
      7211: inst = 32'h10408000;
      7212: inst = 32'hc4051fc;
      7213: inst = 32'h8220000;
      7214: inst = 32'h10408000;
      7215: inst = 32'hc40520a;
      7216: inst = 32'h8220000;
      7217: inst = 32'h10408000;
      7218: inst = 32'hc40520b;
      7219: inst = 32'h8220000;
      7220: inst = 32'h10408000;
      7221: inst = 32'hc40520c;
      7222: inst = 32'h8220000;
      7223: inst = 32'h10408000;
      7224: inst = 32'hc40520d;
      7225: inst = 32'h8220000;
      7226: inst = 32'h10408000;
      7227: inst = 32'hc40520e;
      7228: inst = 32'h8220000;
      7229: inst = 32'h10408000;
      7230: inst = 32'hc40520f;
      7231: inst = 32'h8220000;
      7232: inst = 32'h10408000;
      7233: inst = 32'hc405210;
      7234: inst = 32'h8220000;
      7235: inst = 32'h10408000;
      7236: inst = 32'hc405211;
      7237: inst = 32'h8220000;
      7238: inst = 32'h10408000;
      7239: inst = 32'hc405212;
      7240: inst = 32'h8220000;
      7241: inst = 32'h10408000;
      7242: inst = 32'hc405213;
      7243: inst = 32'h8220000;
      7244: inst = 32'h10408000;
      7245: inst = 32'hc405214;
      7246: inst = 32'h8220000;
      7247: inst = 32'h10408000;
      7248: inst = 32'hc405215;
      7249: inst = 32'h8220000;
      7250: inst = 32'h10408000;
      7251: inst = 32'hc405223;
      7252: inst = 32'h8220000;
      7253: inst = 32'h10408000;
      7254: inst = 32'hc405224;
      7255: inst = 32'h8220000;
      7256: inst = 32'h10408000;
      7257: inst = 32'hc405225;
      7258: inst = 32'h8220000;
      7259: inst = 32'h10408000;
      7260: inst = 32'hc405226;
      7261: inst = 32'h8220000;
      7262: inst = 32'h10408000;
      7263: inst = 32'hc405227;
      7264: inst = 32'h8220000;
      7265: inst = 32'h10408000;
      7266: inst = 32'hc405228;
      7267: inst = 32'h8220000;
      7268: inst = 32'h10408000;
      7269: inst = 32'hc405229;
      7270: inst = 32'h8220000;
      7271: inst = 32'h10408000;
      7272: inst = 32'hc40522a;
      7273: inst = 32'h8220000;
      7274: inst = 32'h10408000;
      7275: inst = 32'hc40522b;
      7276: inst = 32'h8220000;
      7277: inst = 32'h10408000;
      7278: inst = 32'hc40522c;
      7279: inst = 32'h8220000;
      7280: inst = 32'h10408000;
      7281: inst = 32'hc40522d;
      7282: inst = 32'h8220000;
      7283: inst = 32'h10408000;
      7284: inst = 32'hc40522e;
      7285: inst = 32'h8220000;
      7286: inst = 32'h10408000;
      7287: inst = 32'hc405257;
      7288: inst = 32'h8220000;
      7289: inst = 32'h10408000;
      7290: inst = 32'hc405258;
      7291: inst = 32'h8220000;
      7292: inst = 32'h10408000;
      7293: inst = 32'hc405259;
      7294: inst = 32'h8220000;
      7295: inst = 32'h10408000;
      7296: inst = 32'hc40525a;
      7297: inst = 32'h8220000;
      7298: inst = 32'h10408000;
      7299: inst = 32'hc40525b;
      7300: inst = 32'h8220000;
      7301: inst = 32'h10408000;
      7302: inst = 32'hc40526a;
      7303: inst = 32'h8220000;
      7304: inst = 32'h10408000;
      7305: inst = 32'hc40526b;
      7306: inst = 32'h8220000;
      7307: inst = 32'h10408000;
      7308: inst = 32'hc40526c;
      7309: inst = 32'h8220000;
      7310: inst = 32'h10408000;
      7311: inst = 32'hc40526d;
      7312: inst = 32'h8220000;
      7313: inst = 32'h10408000;
      7314: inst = 32'hc40526e;
      7315: inst = 32'h8220000;
      7316: inst = 32'h10408000;
      7317: inst = 32'hc40526f;
      7318: inst = 32'h8220000;
      7319: inst = 32'h10408000;
      7320: inst = 32'hc405270;
      7321: inst = 32'h8220000;
      7322: inst = 32'h10408000;
      7323: inst = 32'hc405271;
      7324: inst = 32'h8220000;
      7325: inst = 32'h10408000;
      7326: inst = 32'hc405272;
      7327: inst = 32'h8220000;
      7328: inst = 32'h10408000;
      7329: inst = 32'hc405273;
      7330: inst = 32'h8220000;
      7331: inst = 32'h10408000;
      7332: inst = 32'hc405274;
      7333: inst = 32'h8220000;
      7334: inst = 32'h10408000;
      7335: inst = 32'hc405275;
      7336: inst = 32'h8220000;
      7337: inst = 32'h10408000;
      7338: inst = 32'hc405284;
      7339: inst = 32'h8220000;
      7340: inst = 32'h10408000;
      7341: inst = 32'hc405285;
      7342: inst = 32'h8220000;
      7343: inst = 32'h10408000;
      7344: inst = 32'hc405286;
      7345: inst = 32'h8220000;
      7346: inst = 32'h10408000;
      7347: inst = 32'hc405287;
      7348: inst = 32'h8220000;
      7349: inst = 32'h10408000;
      7350: inst = 32'hc405288;
      7351: inst = 32'h8220000;
      7352: inst = 32'h10408000;
      7353: inst = 32'hc405289;
      7354: inst = 32'h8220000;
      7355: inst = 32'h10408000;
      7356: inst = 32'hc40528a;
      7357: inst = 32'h8220000;
      7358: inst = 32'h10408000;
      7359: inst = 32'hc40528b;
      7360: inst = 32'h8220000;
      7361: inst = 32'h10408000;
      7362: inst = 32'hc40528c;
      7363: inst = 32'h8220000;
      7364: inst = 32'h10408000;
      7365: inst = 32'hc40528d;
      7366: inst = 32'h8220000;
      7367: inst = 32'h10408000;
      7368: inst = 32'hc40528e;
      7369: inst = 32'h8220000;
      7370: inst = 32'h10408000;
      7371: inst = 32'hc4052b7;
      7372: inst = 32'h8220000;
      7373: inst = 32'h10408000;
      7374: inst = 32'hc4052b8;
      7375: inst = 32'h8220000;
      7376: inst = 32'h10408000;
      7377: inst = 32'hc4052b9;
      7378: inst = 32'h8220000;
      7379: inst = 32'h10408000;
      7380: inst = 32'hc4052ba;
      7381: inst = 32'h8220000;
      7382: inst = 32'h10408000;
      7383: inst = 32'hc4052bb;
      7384: inst = 32'h8220000;
      7385: inst = 32'h10408000;
      7386: inst = 32'hc4052ca;
      7387: inst = 32'h8220000;
      7388: inst = 32'h10408000;
      7389: inst = 32'hc4052cb;
      7390: inst = 32'h8220000;
      7391: inst = 32'h10408000;
      7392: inst = 32'hc4052cc;
      7393: inst = 32'h8220000;
      7394: inst = 32'h10408000;
      7395: inst = 32'hc4052cd;
      7396: inst = 32'h8220000;
      7397: inst = 32'h10408000;
      7398: inst = 32'hc4052ce;
      7399: inst = 32'h8220000;
      7400: inst = 32'h10408000;
      7401: inst = 32'hc4052cf;
      7402: inst = 32'h8220000;
      7403: inst = 32'h10408000;
      7404: inst = 32'hc4052d0;
      7405: inst = 32'h8220000;
      7406: inst = 32'h10408000;
      7407: inst = 32'hc4052d1;
      7408: inst = 32'h8220000;
      7409: inst = 32'h10408000;
      7410: inst = 32'hc4052d2;
      7411: inst = 32'h8220000;
      7412: inst = 32'h10408000;
      7413: inst = 32'hc4052d3;
      7414: inst = 32'h8220000;
      7415: inst = 32'h10408000;
      7416: inst = 32'hc4052d4;
      7417: inst = 32'h8220000;
      7418: inst = 32'h10408000;
      7419: inst = 32'hc4052d5;
      7420: inst = 32'h8220000;
      7421: inst = 32'h10408000;
      7422: inst = 32'hc4052e4;
      7423: inst = 32'h8220000;
      7424: inst = 32'h10408000;
      7425: inst = 32'hc4052e5;
      7426: inst = 32'h8220000;
      7427: inst = 32'h10408000;
      7428: inst = 32'hc4052e6;
      7429: inst = 32'h8220000;
      7430: inst = 32'h10408000;
      7431: inst = 32'hc4052e7;
      7432: inst = 32'h8220000;
      7433: inst = 32'h10408000;
      7434: inst = 32'hc4052e8;
      7435: inst = 32'h8220000;
      7436: inst = 32'h10408000;
      7437: inst = 32'hc4052e9;
      7438: inst = 32'h8220000;
      7439: inst = 32'h10408000;
      7440: inst = 32'hc4052ea;
      7441: inst = 32'h8220000;
      7442: inst = 32'h10408000;
      7443: inst = 32'hc4052eb;
      7444: inst = 32'h8220000;
      7445: inst = 32'h10408000;
      7446: inst = 32'hc4052ec;
      7447: inst = 32'h8220000;
      7448: inst = 32'h10408000;
      7449: inst = 32'hc4052ed;
      7450: inst = 32'h8220000;
      7451: inst = 32'h10408000;
      7452: inst = 32'hc4052ee;
      7453: inst = 32'h8220000;
      7454: inst = 32'hc2094b2;
      7455: inst = 32'h10408000;
      7456: inst = 32'hc403feb;
      7457: inst = 32'h8220000;
      7458: inst = 32'h10408000;
      7459: inst = 32'hc40404b;
      7460: inst = 32'h8220000;
      7461: inst = 32'h10408000;
      7462: inst = 32'hc4040ab;
      7463: inst = 32'h8220000;
      7464: inst = 32'h10408000;
      7465: inst = 32'hc40410b;
      7466: inst = 32'h8220000;
      7467: inst = 32'h10408000;
      7468: inst = 32'hc40416b;
      7469: inst = 32'h8220000;
      7470: inst = 32'h10408000;
      7471: inst = 32'hc4041cb;
      7472: inst = 32'h8220000;
      7473: inst = 32'h10408000;
      7474: inst = 32'hc40422b;
      7475: inst = 32'h8220000;
      7476: inst = 32'h10408000;
      7477: inst = 32'hc40428b;
      7478: inst = 32'h8220000;
      7479: inst = 32'hc20b596;
      7480: inst = 32'h10408000;
      7481: inst = 32'hc4041da;
      7482: inst = 32'h8220000;
      7483: inst = 32'h10408000;
      7484: inst = 32'hc4041db;
      7485: inst = 32'h8220000;
      7486: inst = 32'h10408000;
      7487: inst = 32'hc4041dc;
      7488: inst = 32'h8220000;
      7489: inst = 32'h10408000;
      7490: inst = 32'hc4041dd;
      7491: inst = 32'h8220000;
      7492: inst = 32'h10408000;
      7493: inst = 32'hc4041de;
      7494: inst = 32'h8220000;
      7495: inst = 32'h10408000;
      7496: inst = 32'hc4041df;
      7497: inst = 32'h8220000;
      7498: inst = 32'h10408000;
      7499: inst = 32'hc4041e0;
      7500: inst = 32'h8220000;
      7501: inst = 32'h10408000;
      7502: inst = 32'hc4041e1;
      7503: inst = 32'h8220000;
      7504: inst = 32'h10408000;
      7505: inst = 32'hc4041e2;
      7506: inst = 32'h8220000;
      7507: inst = 32'h10408000;
      7508: inst = 32'hc4041e3;
      7509: inst = 32'h8220000;
      7510: inst = 32'h10408000;
      7511: inst = 32'hc4041e4;
      7512: inst = 32'h8220000;
      7513: inst = 32'h10408000;
      7514: inst = 32'hc4041e5;
      7515: inst = 32'h8220000;
      7516: inst = 32'h10408000;
      7517: inst = 32'hc4041e6;
      7518: inst = 32'h8220000;
      7519: inst = 32'h10408000;
      7520: inst = 32'hc4041e7;
      7521: inst = 32'h8220000;
      7522: inst = 32'h10408000;
      7523: inst = 32'hc4041e8;
      7524: inst = 32'h8220000;
      7525: inst = 32'h10408000;
      7526: inst = 32'hc4041e9;
      7527: inst = 32'h8220000;
      7528: inst = 32'h10408000;
      7529: inst = 32'hc4041ea;
      7530: inst = 32'h8220000;
      7531: inst = 32'h10408000;
      7532: inst = 32'hc4041eb;
      7533: inst = 32'h8220000;
      7534: inst = 32'h10408000;
      7535: inst = 32'hc4041ec;
      7536: inst = 32'h8220000;
      7537: inst = 32'h10408000;
      7538: inst = 32'hc4041ed;
      7539: inst = 32'h8220000;
      7540: inst = 32'h10408000;
      7541: inst = 32'hc4041ee;
      7542: inst = 32'h8220000;
      7543: inst = 32'h10408000;
      7544: inst = 32'hc4041ef;
      7545: inst = 32'h8220000;
      7546: inst = 32'h10408000;
      7547: inst = 32'hc4041f0;
      7548: inst = 32'h8220000;
      7549: inst = 32'h10408000;
      7550: inst = 32'hc4041f1;
      7551: inst = 32'h8220000;
      7552: inst = 32'h10408000;
      7553: inst = 32'hc4041f2;
      7554: inst = 32'h8220000;
      7555: inst = 32'h10408000;
      7556: inst = 32'hc4041f3;
      7557: inst = 32'h8220000;
      7558: inst = 32'h10408000;
      7559: inst = 32'hc4041f4;
      7560: inst = 32'h8220000;
      7561: inst = 32'h10408000;
      7562: inst = 32'hc4041f5;
      7563: inst = 32'h8220000;
      7564: inst = 32'h10408000;
      7565: inst = 32'hc4041f6;
      7566: inst = 32'h8220000;
      7567: inst = 32'h10408000;
      7568: inst = 32'hc4041f7;
      7569: inst = 32'h8220000;
      7570: inst = 32'h10408000;
      7571: inst = 32'hc4041f8;
      7572: inst = 32'h8220000;
      7573: inst = 32'h10408000;
      7574: inst = 32'hc4041f9;
      7575: inst = 32'h8220000;
      7576: inst = 32'h10408000;
      7577: inst = 32'hc4041fa;
      7578: inst = 32'h8220000;
      7579: inst = 32'h10408000;
      7580: inst = 32'hc4041fb;
      7581: inst = 32'h8220000;
      7582: inst = 32'h10408000;
      7583: inst = 32'hc4041fc;
      7584: inst = 32'h8220000;
      7585: inst = 32'h10408000;
      7586: inst = 32'hc4041fd;
      7587: inst = 32'h8220000;
      7588: inst = 32'h10408000;
      7589: inst = 32'hc4041fe;
      7590: inst = 32'h8220000;
      7591: inst = 32'h10408000;
      7592: inst = 32'hc4041ff;
      7593: inst = 32'h8220000;
      7594: inst = 32'h10408000;
      7595: inst = 32'hc404200;
      7596: inst = 32'h8220000;
      7597: inst = 32'h10408000;
      7598: inst = 32'hc404201;
      7599: inst = 32'h8220000;
      7600: inst = 32'h10408000;
      7601: inst = 32'hc404202;
      7602: inst = 32'h8220000;
      7603: inst = 32'h10408000;
      7604: inst = 32'hc404203;
      7605: inst = 32'h8220000;
      7606: inst = 32'h10408000;
      7607: inst = 32'hc404204;
      7608: inst = 32'h8220000;
      7609: inst = 32'h10408000;
      7610: inst = 32'hc404205;
      7611: inst = 32'h8220000;
      7612: inst = 32'h10408000;
      7613: inst = 32'hc404bfa;
      7614: inst = 32'h8220000;
      7615: inst = 32'h10408000;
      7616: inst = 32'hc404bfb;
      7617: inst = 32'h8220000;
      7618: inst = 32'h10408000;
      7619: inst = 32'hc404bfc;
      7620: inst = 32'h8220000;
      7621: inst = 32'h10408000;
      7622: inst = 32'hc404bfd;
      7623: inst = 32'h8220000;
      7624: inst = 32'h10408000;
      7625: inst = 32'hc404bfe;
      7626: inst = 32'h8220000;
      7627: inst = 32'h10408000;
      7628: inst = 32'hc404bff;
      7629: inst = 32'h8220000;
      7630: inst = 32'h10408000;
      7631: inst = 32'hc404c00;
      7632: inst = 32'h8220000;
      7633: inst = 32'h10408000;
      7634: inst = 32'hc404c01;
      7635: inst = 32'h8220000;
      7636: inst = 32'h10408000;
      7637: inst = 32'hc404c02;
      7638: inst = 32'h8220000;
      7639: inst = 32'h10408000;
      7640: inst = 32'hc404c03;
      7641: inst = 32'h8220000;
      7642: inst = 32'h10408000;
      7643: inst = 32'hc404c04;
      7644: inst = 32'h8220000;
      7645: inst = 32'h10408000;
      7646: inst = 32'hc404c05;
      7647: inst = 32'h8220000;
      7648: inst = 32'h10408000;
      7649: inst = 32'hc404c06;
      7650: inst = 32'h8220000;
      7651: inst = 32'h10408000;
      7652: inst = 32'hc404c07;
      7653: inst = 32'h8220000;
      7654: inst = 32'h10408000;
      7655: inst = 32'hc404c08;
      7656: inst = 32'h8220000;
      7657: inst = 32'h10408000;
      7658: inst = 32'hc404c09;
      7659: inst = 32'h8220000;
      7660: inst = 32'h10408000;
      7661: inst = 32'hc404c0a;
      7662: inst = 32'h8220000;
      7663: inst = 32'h10408000;
      7664: inst = 32'hc404c0b;
      7665: inst = 32'h8220000;
      7666: inst = 32'h10408000;
      7667: inst = 32'hc404c0c;
      7668: inst = 32'h8220000;
      7669: inst = 32'h10408000;
      7670: inst = 32'hc404c0d;
      7671: inst = 32'h8220000;
      7672: inst = 32'h10408000;
      7673: inst = 32'hc404c0e;
      7674: inst = 32'h8220000;
      7675: inst = 32'h10408000;
      7676: inst = 32'hc404c0f;
      7677: inst = 32'h8220000;
      7678: inst = 32'h10408000;
      7679: inst = 32'hc404c10;
      7680: inst = 32'h8220000;
      7681: inst = 32'h10408000;
      7682: inst = 32'hc404c11;
      7683: inst = 32'h8220000;
      7684: inst = 32'h10408000;
      7685: inst = 32'hc404c12;
      7686: inst = 32'h8220000;
      7687: inst = 32'h10408000;
      7688: inst = 32'hc404c13;
      7689: inst = 32'h8220000;
      7690: inst = 32'h10408000;
      7691: inst = 32'hc404c14;
      7692: inst = 32'h8220000;
      7693: inst = 32'h10408000;
      7694: inst = 32'hc404c15;
      7695: inst = 32'h8220000;
      7696: inst = 32'h10408000;
      7697: inst = 32'hc404c16;
      7698: inst = 32'h8220000;
      7699: inst = 32'h10408000;
      7700: inst = 32'hc404c17;
      7701: inst = 32'h8220000;
      7702: inst = 32'h10408000;
      7703: inst = 32'hc404c18;
      7704: inst = 32'h8220000;
      7705: inst = 32'h10408000;
      7706: inst = 32'hc404c19;
      7707: inst = 32'h8220000;
      7708: inst = 32'h10408000;
      7709: inst = 32'hc404c1a;
      7710: inst = 32'h8220000;
      7711: inst = 32'h10408000;
      7712: inst = 32'hc404c1b;
      7713: inst = 32'h8220000;
      7714: inst = 32'h10408000;
      7715: inst = 32'hc404c1c;
      7716: inst = 32'h8220000;
      7717: inst = 32'h10408000;
      7718: inst = 32'hc404c1d;
      7719: inst = 32'h8220000;
      7720: inst = 32'h10408000;
      7721: inst = 32'hc404c1e;
      7722: inst = 32'h8220000;
      7723: inst = 32'h10408000;
      7724: inst = 32'hc404c1f;
      7725: inst = 32'h8220000;
      7726: inst = 32'h10408000;
      7727: inst = 32'hc404c20;
      7728: inst = 32'h8220000;
      7729: inst = 32'h10408000;
      7730: inst = 32'hc404c21;
      7731: inst = 32'h8220000;
      7732: inst = 32'h10408000;
      7733: inst = 32'hc404c22;
      7734: inst = 32'h8220000;
      7735: inst = 32'h10408000;
      7736: inst = 32'hc404c23;
      7737: inst = 32'h8220000;
      7738: inst = 32'h10408000;
      7739: inst = 32'hc404c24;
      7740: inst = 32'h8220000;
      7741: inst = 32'h10408000;
      7742: inst = 32'hc404c25;
      7743: inst = 32'h8220000;
      7744: inst = 32'hc20ffff;
      7745: inst = 32'h10408000;
      7746: inst = 32'hc40423c;
      7747: inst = 32'h8220000;
      7748: inst = 32'h10408000;
      7749: inst = 32'hc40423d;
      7750: inst = 32'h8220000;
      7751: inst = 32'h10408000;
      7752: inst = 32'hc40423e;
      7753: inst = 32'h8220000;
      7754: inst = 32'h10408000;
      7755: inst = 32'hc40423f;
      7756: inst = 32'h8220000;
      7757: inst = 32'h10408000;
      7758: inst = 32'hc404240;
      7759: inst = 32'h8220000;
      7760: inst = 32'h10408000;
      7761: inst = 32'hc404241;
      7762: inst = 32'h8220000;
      7763: inst = 32'h10408000;
      7764: inst = 32'hc404242;
      7765: inst = 32'h8220000;
      7766: inst = 32'h10408000;
      7767: inst = 32'hc404243;
      7768: inst = 32'h8220000;
      7769: inst = 32'h10408000;
      7770: inst = 32'hc404244;
      7771: inst = 32'h8220000;
      7772: inst = 32'h10408000;
      7773: inst = 32'hc404245;
      7774: inst = 32'h8220000;
      7775: inst = 32'h10408000;
      7776: inst = 32'hc404246;
      7777: inst = 32'h8220000;
      7778: inst = 32'h10408000;
      7779: inst = 32'hc404247;
      7780: inst = 32'h8220000;
      7781: inst = 32'h10408000;
      7782: inst = 32'hc404248;
      7783: inst = 32'h8220000;
      7784: inst = 32'h10408000;
      7785: inst = 32'hc404249;
      7786: inst = 32'h8220000;
      7787: inst = 32'h10408000;
      7788: inst = 32'hc40424a;
      7789: inst = 32'h8220000;
      7790: inst = 32'h10408000;
      7791: inst = 32'hc40424b;
      7792: inst = 32'h8220000;
      7793: inst = 32'h10408000;
      7794: inst = 32'hc40424c;
      7795: inst = 32'h8220000;
      7796: inst = 32'h10408000;
      7797: inst = 32'hc40424d;
      7798: inst = 32'h8220000;
      7799: inst = 32'h10408000;
      7800: inst = 32'hc40424e;
      7801: inst = 32'h8220000;
      7802: inst = 32'h10408000;
      7803: inst = 32'hc40424f;
      7804: inst = 32'h8220000;
      7805: inst = 32'h10408000;
      7806: inst = 32'hc404250;
      7807: inst = 32'h8220000;
      7808: inst = 32'h10408000;
      7809: inst = 32'hc404251;
      7810: inst = 32'h8220000;
      7811: inst = 32'h10408000;
      7812: inst = 32'hc404252;
      7813: inst = 32'h8220000;
      7814: inst = 32'h10408000;
      7815: inst = 32'hc404253;
      7816: inst = 32'h8220000;
      7817: inst = 32'h10408000;
      7818: inst = 32'hc404254;
      7819: inst = 32'h8220000;
      7820: inst = 32'h10408000;
      7821: inst = 32'hc404255;
      7822: inst = 32'h8220000;
      7823: inst = 32'h10408000;
      7824: inst = 32'hc404256;
      7825: inst = 32'h8220000;
      7826: inst = 32'h10408000;
      7827: inst = 32'hc404257;
      7828: inst = 32'h8220000;
      7829: inst = 32'h10408000;
      7830: inst = 32'hc404258;
      7831: inst = 32'h8220000;
      7832: inst = 32'h10408000;
      7833: inst = 32'hc404259;
      7834: inst = 32'h8220000;
      7835: inst = 32'h10408000;
      7836: inst = 32'hc40425a;
      7837: inst = 32'h8220000;
      7838: inst = 32'h10408000;
      7839: inst = 32'hc40425b;
      7840: inst = 32'h8220000;
      7841: inst = 32'h10408000;
      7842: inst = 32'hc40425c;
      7843: inst = 32'h8220000;
      7844: inst = 32'h10408000;
      7845: inst = 32'hc40425d;
      7846: inst = 32'h8220000;
      7847: inst = 32'h10408000;
      7848: inst = 32'hc40425e;
      7849: inst = 32'h8220000;
      7850: inst = 32'h10408000;
      7851: inst = 32'hc40425f;
      7852: inst = 32'h8220000;
      7853: inst = 32'h10408000;
      7854: inst = 32'hc404260;
      7855: inst = 32'h8220000;
      7856: inst = 32'h10408000;
      7857: inst = 32'hc404261;
      7858: inst = 32'h8220000;
      7859: inst = 32'h10408000;
      7860: inst = 32'hc404262;
      7861: inst = 32'h8220000;
      7862: inst = 32'h10408000;
      7863: inst = 32'hc404263;
      7864: inst = 32'h8220000;
      7865: inst = 32'h10408000;
      7866: inst = 32'hc40429c;
      7867: inst = 32'h8220000;
      7868: inst = 32'h10408000;
      7869: inst = 32'hc40429d;
      7870: inst = 32'h8220000;
      7871: inst = 32'h10408000;
      7872: inst = 32'hc40429e;
      7873: inst = 32'h8220000;
      7874: inst = 32'h10408000;
      7875: inst = 32'hc40429f;
      7876: inst = 32'h8220000;
      7877: inst = 32'h10408000;
      7878: inst = 32'hc4042a0;
      7879: inst = 32'h8220000;
      7880: inst = 32'h10408000;
      7881: inst = 32'hc4042a1;
      7882: inst = 32'h8220000;
      7883: inst = 32'h10408000;
      7884: inst = 32'hc4042a2;
      7885: inst = 32'h8220000;
      7886: inst = 32'h10408000;
      7887: inst = 32'hc4042a3;
      7888: inst = 32'h8220000;
      7889: inst = 32'h10408000;
      7890: inst = 32'hc4042a4;
      7891: inst = 32'h8220000;
      7892: inst = 32'h10408000;
      7893: inst = 32'hc4042a5;
      7894: inst = 32'h8220000;
      7895: inst = 32'h10408000;
      7896: inst = 32'hc4042a6;
      7897: inst = 32'h8220000;
      7898: inst = 32'h10408000;
      7899: inst = 32'hc4042a7;
      7900: inst = 32'h8220000;
      7901: inst = 32'h10408000;
      7902: inst = 32'hc4042a8;
      7903: inst = 32'h8220000;
      7904: inst = 32'h10408000;
      7905: inst = 32'hc4042a9;
      7906: inst = 32'h8220000;
      7907: inst = 32'h10408000;
      7908: inst = 32'hc4042aa;
      7909: inst = 32'h8220000;
      7910: inst = 32'h10408000;
      7911: inst = 32'hc4042ab;
      7912: inst = 32'h8220000;
      7913: inst = 32'h10408000;
      7914: inst = 32'hc4042ac;
      7915: inst = 32'h8220000;
      7916: inst = 32'h10408000;
      7917: inst = 32'hc4042ad;
      7918: inst = 32'h8220000;
      7919: inst = 32'h10408000;
      7920: inst = 32'hc4042ae;
      7921: inst = 32'h8220000;
      7922: inst = 32'h10408000;
      7923: inst = 32'hc4042af;
      7924: inst = 32'h8220000;
      7925: inst = 32'h10408000;
      7926: inst = 32'hc4042b0;
      7927: inst = 32'h8220000;
      7928: inst = 32'h10408000;
      7929: inst = 32'hc4042b1;
      7930: inst = 32'h8220000;
      7931: inst = 32'h10408000;
      7932: inst = 32'hc4042b2;
      7933: inst = 32'h8220000;
      7934: inst = 32'h10408000;
      7935: inst = 32'hc4042b3;
      7936: inst = 32'h8220000;
      7937: inst = 32'h10408000;
      7938: inst = 32'hc4042b4;
      7939: inst = 32'h8220000;
      7940: inst = 32'h10408000;
      7941: inst = 32'hc4042b5;
      7942: inst = 32'h8220000;
      7943: inst = 32'h10408000;
      7944: inst = 32'hc4042b6;
      7945: inst = 32'h8220000;
      7946: inst = 32'h10408000;
      7947: inst = 32'hc4042b7;
      7948: inst = 32'h8220000;
      7949: inst = 32'h10408000;
      7950: inst = 32'hc4042b8;
      7951: inst = 32'h8220000;
      7952: inst = 32'h10408000;
      7953: inst = 32'hc4042b9;
      7954: inst = 32'h8220000;
      7955: inst = 32'h10408000;
      7956: inst = 32'hc4042ba;
      7957: inst = 32'h8220000;
      7958: inst = 32'h10408000;
      7959: inst = 32'hc4042bb;
      7960: inst = 32'h8220000;
      7961: inst = 32'h10408000;
      7962: inst = 32'hc4042bc;
      7963: inst = 32'h8220000;
      7964: inst = 32'h10408000;
      7965: inst = 32'hc4042bd;
      7966: inst = 32'h8220000;
      7967: inst = 32'h10408000;
      7968: inst = 32'hc4042be;
      7969: inst = 32'h8220000;
      7970: inst = 32'h10408000;
      7971: inst = 32'hc4042bf;
      7972: inst = 32'h8220000;
      7973: inst = 32'h10408000;
      7974: inst = 32'hc4042c0;
      7975: inst = 32'h8220000;
      7976: inst = 32'h10408000;
      7977: inst = 32'hc4042c1;
      7978: inst = 32'h8220000;
      7979: inst = 32'h10408000;
      7980: inst = 32'hc4042c2;
      7981: inst = 32'h8220000;
      7982: inst = 32'h10408000;
      7983: inst = 32'hc4042c3;
      7984: inst = 32'h8220000;
      7985: inst = 32'h10408000;
      7986: inst = 32'hc4042fc;
      7987: inst = 32'h8220000;
      7988: inst = 32'h10408000;
      7989: inst = 32'hc4042fd;
      7990: inst = 32'h8220000;
      7991: inst = 32'h10408000;
      7992: inst = 32'hc4042fe;
      7993: inst = 32'h8220000;
      7994: inst = 32'h10408000;
      7995: inst = 32'hc4042ff;
      7996: inst = 32'h8220000;
      7997: inst = 32'h10408000;
      7998: inst = 32'hc404300;
      7999: inst = 32'h8220000;
      8000: inst = 32'h10408000;
      8001: inst = 32'hc404301;
      8002: inst = 32'h8220000;
      8003: inst = 32'h10408000;
      8004: inst = 32'hc404302;
      8005: inst = 32'h8220000;
      8006: inst = 32'h10408000;
      8007: inst = 32'hc404303;
      8008: inst = 32'h8220000;
      8009: inst = 32'h10408000;
      8010: inst = 32'hc404304;
      8011: inst = 32'h8220000;
      8012: inst = 32'h10408000;
      8013: inst = 32'hc404305;
      8014: inst = 32'h8220000;
      8015: inst = 32'h10408000;
      8016: inst = 32'hc404306;
      8017: inst = 32'h8220000;
      8018: inst = 32'h10408000;
      8019: inst = 32'hc404307;
      8020: inst = 32'h8220000;
      8021: inst = 32'h10408000;
      8022: inst = 32'hc404308;
      8023: inst = 32'h8220000;
      8024: inst = 32'h10408000;
      8025: inst = 32'hc404309;
      8026: inst = 32'h8220000;
      8027: inst = 32'h10408000;
      8028: inst = 32'hc40430a;
      8029: inst = 32'h8220000;
      8030: inst = 32'h10408000;
      8031: inst = 32'hc40430b;
      8032: inst = 32'h8220000;
      8033: inst = 32'h10408000;
      8034: inst = 32'hc40430c;
      8035: inst = 32'h8220000;
      8036: inst = 32'h10408000;
      8037: inst = 32'hc40430d;
      8038: inst = 32'h8220000;
      8039: inst = 32'h10408000;
      8040: inst = 32'hc40430e;
      8041: inst = 32'h8220000;
      8042: inst = 32'h10408000;
      8043: inst = 32'hc40430f;
      8044: inst = 32'h8220000;
      8045: inst = 32'h10408000;
      8046: inst = 32'hc404310;
      8047: inst = 32'h8220000;
      8048: inst = 32'h10408000;
      8049: inst = 32'hc404311;
      8050: inst = 32'h8220000;
      8051: inst = 32'h10408000;
      8052: inst = 32'hc404312;
      8053: inst = 32'h8220000;
      8054: inst = 32'h10408000;
      8055: inst = 32'hc404313;
      8056: inst = 32'h8220000;
      8057: inst = 32'h10408000;
      8058: inst = 32'hc404314;
      8059: inst = 32'h8220000;
      8060: inst = 32'h10408000;
      8061: inst = 32'hc404315;
      8062: inst = 32'h8220000;
      8063: inst = 32'h10408000;
      8064: inst = 32'hc404316;
      8065: inst = 32'h8220000;
      8066: inst = 32'h10408000;
      8067: inst = 32'hc404317;
      8068: inst = 32'h8220000;
      8069: inst = 32'h10408000;
      8070: inst = 32'hc404318;
      8071: inst = 32'h8220000;
      8072: inst = 32'h10408000;
      8073: inst = 32'hc404319;
      8074: inst = 32'h8220000;
      8075: inst = 32'h10408000;
      8076: inst = 32'hc40431a;
      8077: inst = 32'h8220000;
      8078: inst = 32'h10408000;
      8079: inst = 32'hc40431b;
      8080: inst = 32'h8220000;
      8081: inst = 32'h10408000;
      8082: inst = 32'hc40431c;
      8083: inst = 32'h8220000;
      8084: inst = 32'h10408000;
      8085: inst = 32'hc40431d;
      8086: inst = 32'h8220000;
      8087: inst = 32'h10408000;
      8088: inst = 32'hc40431e;
      8089: inst = 32'h8220000;
      8090: inst = 32'h10408000;
      8091: inst = 32'hc40431f;
      8092: inst = 32'h8220000;
      8093: inst = 32'h10408000;
      8094: inst = 32'hc404320;
      8095: inst = 32'h8220000;
      8096: inst = 32'h10408000;
      8097: inst = 32'hc404321;
      8098: inst = 32'h8220000;
      8099: inst = 32'h10408000;
      8100: inst = 32'hc404322;
      8101: inst = 32'h8220000;
      8102: inst = 32'h10408000;
      8103: inst = 32'hc404323;
      8104: inst = 32'h8220000;
      8105: inst = 32'h10408000;
      8106: inst = 32'hc40435c;
      8107: inst = 32'h8220000;
      8108: inst = 32'h10408000;
      8109: inst = 32'hc40435d;
      8110: inst = 32'h8220000;
      8111: inst = 32'h10408000;
      8112: inst = 32'hc40435e;
      8113: inst = 32'h8220000;
      8114: inst = 32'h10408000;
      8115: inst = 32'hc40435f;
      8116: inst = 32'h8220000;
      8117: inst = 32'h10408000;
      8118: inst = 32'hc404360;
      8119: inst = 32'h8220000;
      8120: inst = 32'h10408000;
      8121: inst = 32'hc404361;
      8122: inst = 32'h8220000;
      8123: inst = 32'h10408000;
      8124: inst = 32'hc404362;
      8125: inst = 32'h8220000;
      8126: inst = 32'h10408000;
      8127: inst = 32'hc404363;
      8128: inst = 32'h8220000;
      8129: inst = 32'h10408000;
      8130: inst = 32'hc404364;
      8131: inst = 32'h8220000;
      8132: inst = 32'h10408000;
      8133: inst = 32'hc404365;
      8134: inst = 32'h8220000;
      8135: inst = 32'h10408000;
      8136: inst = 32'hc404366;
      8137: inst = 32'h8220000;
      8138: inst = 32'h10408000;
      8139: inst = 32'hc404367;
      8140: inst = 32'h8220000;
      8141: inst = 32'h10408000;
      8142: inst = 32'hc404368;
      8143: inst = 32'h8220000;
      8144: inst = 32'h10408000;
      8145: inst = 32'hc404369;
      8146: inst = 32'h8220000;
      8147: inst = 32'h10408000;
      8148: inst = 32'hc40436a;
      8149: inst = 32'h8220000;
      8150: inst = 32'h10408000;
      8151: inst = 32'hc40436b;
      8152: inst = 32'h8220000;
      8153: inst = 32'h10408000;
      8154: inst = 32'hc40436c;
      8155: inst = 32'h8220000;
      8156: inst = 32'h10408000;
      8157: inst = 32'hc40436d;
      8158: inst = 32'h8220000;
      8159: inst = 32'h10408000;
      8160: inst = 32'hc40436e;
      8161: inst = 32'h8220000;
      8162: inst = 32'h10408000;
      8163: inst = 32'hc40436f;
      8164: inst = 32'h8220000;
      8165: inst = 32'h10408000;
      8166: inst = 32'hc404370;
      8167: inst = 32'h8220000;
      8168: inst = 32'h10408000;
      8169: inst = 32'hc404371;
      8170: inst = 32'h8220000;
      8171: inst = 32'h10408000;
      8172: inst = 32'hc404372;
      8173: inst = 32'h8220000;
      8174: inst = 32'h10408000;
      8175: inst = 32'hc404373;
      8176: inst = 32'h8220000;
      8177: inst = 32'h10408000;
      8178: inst = 32'hc404374;
      8179: inst = 32'h8220000;
      8180: inst = 32'h10408000;
      8181: inst = 32'hc404375;
      8182: inst = 32'h8220000;
      8183: inst = 32'h10408000;
      8184: inst = 32'hc404376;
      8185: inst = 32'h8220000;
      8186: inst = 32'h10408000;
      8187: inst = 32'hc404377;
      8188: inst = 32'h8220000;
      8189: inst = 32'h10408000;
      8190: inst = 32'hc404378;
      8191: inst = 32'h8220000;
      8192: inst = 32'h10408000;
      8193: inst = 32'hc404379;
      8194: inst = 32'h8220000;
      8195: inst = 32'h10408000;
      8196: inst = 32'hc40437a;
      8197: inst = 32'h8220000;
      8198: inst = 32'h10408000;
      8199: inst = 32'hc40437b;
      8200: inst = 32'h8220000;
      8201: inst = 32'h10408000;
      8202: inst = 32'hc40437c;
      8203: inst = 32'h8220000;
      8204: inst = 32'h10408000;
      8205: inst = 32'hc40437d;
      8206: inst = 32'h8220000;
      8207: inst = 32'h10408000;
      8208: inst = 32'hc40437e;
      8209: inst = 32'h8220000;
      8210: inst = 32'h10408000;
      8211: inst = 32'hc40437f;
      8212: inst = 32'h8220000;
      8213: inst = 32'h10408000;
      8214: inst = 32'hc404380;
      8215: inst = 32'h8220000;
      8216: inst = 32'h10408000;
      8217: inst = 32'hc404381;
      8218: inst = 32'h8220000;
      8219: inst = 32'h10408000;
      8220: inst = 32'hc404382;
      8221: inst = 32'h8220000;
      8222: inst = 32'h10408000;
      8223: inst = 32'hc404383;
      8224: inst = 32'h8220000;
      8225: inst = 32'h10408000;
      8226: inst = 32'hc4043bc;
      8227: inst = 32'h8220000;
      8228: inst = 32'h10408000;
      8229: inst = 32'hc4043bd;
      8230: inst = 32'h8220000;
      8231: inst = 32'h10408000;
      8232: inst = 32'hc4043be;
      8233: inst = 32'h8220000;
      8234: inst = 32'h10408000;
      8235: inst = 32'hc4043bf;
      8236: inst = 32'h8220000;
      8237: inst = 32'h10408000;
      8238: inst = 32'hc4043c0;
      8239: inst = 32'h8220000;
      8240: inst = 32'h10408000;
      8241: inst = 32'hc4043c1;
      8242: inst = 32'h8220000;
      8243: inst = 32'h10408000;
      8244: inst = 32'hc4043c2;
      8245: inst = 32'h8220000;
      8246: inst = 32'h10408000;
      8247: inst = 32'hc4043c3;
      8248: inst = 32'h8220000;
      8249: inst = 32'h10408000;
      8250: inst = 32'hc4043c4;
      8251: inst = 32'h8220000;
      8252: inst = 32'h10408000;
      8253: inst = 32'hc4043c5;
      8254: inst = 32'h8220000;
      8255: inst = 32'h10408000;
      8256: inst = 32'hc4043c6;
      8257: inst = 32'h8220000;
      8258: inst = 32'h10408000;
      8259: inst = 32'hc4043c7;
      8260: inst = 32'h8220000;
      8261: inst = 32'h10408000;
      8262: inst = 32'hc4043c8;
      8263: inst = 32'h8220000;
      8264: inst = 32'h10408000;
      8265: inst = 32'hc4043c9;
      8266: inst = 32'h8220000;
      8267: inst = 32'h10408000;
      8268: inst = 32'hc4043ca;
      8269: inst = 32'h8220000;
      8270: inst = 32'h10408000;
      8271: inst = 32'hc4043cb;
      8272: inst = 32'h8220000;
      8273: inst = 32'h10408000;
      8274: inst = 32'hc4043cc;
      8275: inst = 32'h8220000;
      8276: inst = 32'h10408000;
      8277: inst = 32'hc4043cd;
      8278: inst = 32'h8220000;
      8279: inst = 32'h10408000;
      8280: inst = 32'hc4043ce;
      8281: inst = 32'h8220000;
      8282: inst = 32'h10408000;
      8283: inst = 32'hc4043cf;
      8284: inst = 32'h8220000;
      8285: inst = 32'h10408000;
      8286: inst = 32'hc4043d0;
      8287: inst = 32'h8220000;
      8288: inst = 32'h10408000;
      8289: inst = 32'hc4043d1;
      8290: inst = 32'h8220000;
      8291: inst = 32'h10408000;
      8292: inst = 32'hc4043d2;
      8293: inst = 32'h8220000;
      8294: inst = 32'h10408000;
      8295: inst = 32'hc4043d3;
      8296: inst = 32'h8220000;
      8297: inst = 32'h10408000;
      8298: inst = 32'hc4043d4;
      8299: inst = 32'h8220000;
      8300: inst = 32'h10408000;
      8301: inst = 32'hc4043d5;
      8302: inst = 32'h8220000;
      8303: inst = 32'h10408000;
      8304: inst = 32'hc4043d6;
      8305: inst = 32'h8220000;
      8306: inst = 32'h10408000;
      8307: inst = 32'hc4043d7;
      8308: inst = 32'h8220000;
      8309: inst = 32'h10408000;
      8310: inst = 32'hc4043d8;
      8311: inst = 32'h8220000;
      8312: inst = 32'h10408000;
      8313: inst = 32'hc4043d9;
      8314: inst = 32'h8220000;
      8315: inst = 32'h10408000;
      8316: inst = 32'hc4043da;
      8317: inst = 32'h8220000;
      8318: inst = 32'h10408000;
      8319: inst = 32'hc4043db;
      8320: inst = 32'h8220000;
      8321: inst = 32'h10408000;
      8322: inst = 32'hc4043dc;
      8323: inst = 32'h8220000;
      8324: inst = 32'h10408000;
      8325: inst = 32'hc4043dd;
      8326: inst = 32'h8220000;
      8327: inst = 32'h10408000;
      8328: inst = 32'hc4043de;
      8329: inst = 32'h8220000;
      8330: inst = 32'h10408000;
      8331: inst = 32'hc4043df;
      8332: inst = 32'h8220000;
      8333: inst = 32'h10408000;
      8334: inst = 32'hc4043e0;
      8335: inst = 32'h8220000;
      8336: inst = 32'h10408000;
      8337: inst = 32'hc4043e1;
      8338: inst = 32'h8220000;
      8339: inst = 32'h10408000;
      8340: inst = 32'hc4043e2;
      8341: inst = 32'h8220000;
      8342: inst = 32'h10408000;
      8343: inst = 32'hc4043e3;
      8344: inst = 32'h8220000;
      8345: inst = 32'h10408000;
      8346: inst = 32'hc40441c;
      8347: inst = 32'h8220000;
      8348: inst = 32'h10408000;
      8349: inst = 32'hc40441d;
      8350: inst = 32'h8220000;
      8351: inst = 32'h10408000;
      8352: inst = 32'hc40441e;
      8353: inst = 32'h8220000;
      8354: inst = 32'h10408000;
      8355: inst = 32'hc40441f;
      8356: inst = 32'h8220000;
      8357: inst = 32'h10408000;
      8358: inst = 32'hc404420;
      8359: inst = 32'h8220000;
      8360: inst = 32'h10408000;
      8361: inst = 32'hc404421;
      8362: inst = 32'h8220000;
      8363: inst = 32'h10408000;
      8364: inst = 32'hc404422;
      8365: inst = 32'h8220000;
      8366: inst = 32'h10408000;
      8367: inst = 32'hc404423;
      8368: inst = 32'h8220000;
      8369: inst = 32'h10408000;
      8370: inst = 32'hc404424;
      8371: inst = 32'h8220000;
      8372: inst = 32'h10408000;
      8373: inst = 32'hc404425;
      8374: inst = 32'h8220000;
      8375: inst = 32'h10408000;
      8376: inst = 32'hc404426;
      8377: inst = 32'h8220000;
      8378: inst = 32'h10408000;
      8379: inst = 32'hc404427;
      8380: inst = 32'h8220000;
      8381: inst = 32'h10408000;
      8382: inst = 32'hc404428;
      8383: inst = 32'h8220000;
      8384: inst = 32'h10408000;
      8385: inst = 32'hc404429;
      8386: inst = 32'h8220000;
      8387: inst = 32'h10408000;
      8388: inst = 32'hc40442a;
      8389: inst = 32'h8220000;
      8390: inst = 32'h10408000;
      8391: inst = 32'hc40442b;
      8392: inst = 32'h8220000;
      8393: inst = 32'h10408000;
      8394: inst = 32'hc40442c;
      8395: inst = 32'h8220000;
      8396: inst = 32'h10408000;
      8397: inst = 32'hc40442d;
      8398: inst = 32'h8220000;
      8399: inst = 32'h10408000;
      8400: inst = 32'hc40442e;
      8401: inst = 32'h8220000;
      8402: inst = 32'h10408000;
      8403: inst = 32'hc40442f;
      8404: inst = 32'h8220000;
      8405: inst = 32'h10408000;
      8406: inst = 32'hc404430;
      8407: inst = 32'h8220000;
      8408: inst = 32'h10408000;
      8409: inst = 32'hc404431;
      8410: inst = 32'h8220000;
      8411: inst = 32'h10408000;
      8412: inst = 32'hc404432;
      8413: inst = 32'h8220000;
      8414: inst = 32'h10408000;
      8415: inst = 32'hc404433;
      8416: inst = 32'h8220000;
      8417: inst = 32'h10408000;
      8418: inst = 32'hc404434;
      8419: inst = 32'h8220000;
      8420: inst = 32'h10408000;
      8421: inst = 32'hc404435;
      8422: inst = 32'h8220000;
      8423: inst = 32'h10408000;
      8424: inst = 32'hc404436;
      8425: inst = 32'h8220000;
      8426: inst = 32'h10408000;
      8427: inst = 32'hc404437;
      8428: inst = 32'h8220000;
      8429: inst = 32'h10408000;
      8430: inst = 32'hc404438;
      8431: inst = 32'h8220000;
      8432: inst = 32'h10408000;
      8433: inst = 32'hc404439;
      8434: inst = 32'h8220000;
      8435: inst = 32'h10408000;
      8436: inst = 32'hc40443a;
      8437: inst = 32'h8220000;
      8438: inst = 32'h10408000;
      8439: inst = 32'hc40443b;
      8440: inst = 32'h8220000;
      8441: inst = 32'h10408000;
      8442: inst = 32'hc40443c;
      8443: inst = 32'h8220000;
      8444: inst = 32'h10408000;
      8445: inst = 32'hc40443d;
      8446: inst = 32'h8220000;
      8447: inst = 32'h10408000;
      8448: inst = 32'hc40443e;
      8449: inst = 32'h8220000;
      8450: inst = 32'h10408000;
      8451: inst = 32'hc40443f;
      8452: inst = 32'h8220000;
      8453: inst = 32'h10408000;
      8454: inst = 32'hc404440;
      8455: inst = 32'h8220000;
      8456: inst = 32'h10408000;
      8457: inst = 32'hc404441;
      8458: inst = 32'h8220000;
      8459: inst = 32'h10408000;
      8460: inst = 32'hc404442;
      8461: inst = 32'h8220000;
      8462: inst = 32'h10408000;
      8463: inst = 32'hc404443;
      8464: inst = 32'h8220000;
      8465: inst = 32'h10408000;
      8466: inst = 32'hc40447c;
      8467: inst = 32'h8220000;
      8468: inst = 32'h10408000;
      8469: inst = 32'hc40447d;
      8470: inst = 32'h8220000;
      8471: inst = 32'h10408000;
      8472: inst = 32'hc40447e;
      8473: inst = 32'h8220000;
      8474: inst = 32'h10408000;
      8475: inst = 32'hc40447f;
      8476: inst = 32'h8220000;
      8477: inst = 32'h10408000;
      8478: inst = 32'hc404480;
      8479: inst = 32'h8220000;
      8480: inst = 32'h10408000;
      8481: inst = 32'hc404481;
      8482: inst = 32'h8220000;
      8483: inst = 32'h10408000;
      8484: inst = 32'hc404482;
      8485: inst = 32'h8220000;
      8486: inst = 32'h10408000;
      8487: inst = 32'hc404483;
      8488: inst = 32'h8220000;
      8489: inst = 32'h10408000;
      8490: inst = 32'hc404484;
      8491: inst = 32'h8220000;
      8492: inst = 32'h10408000;
      8493: inst = 32'hc404485;
      8494: inst = 32'h8220000;
      8495: inst = 32'h10408000;
      8496: inst = 32'hc404486;
      8497: inst = 32'h8220000;
      8498: inst = 32'h10408000;
      8499: inst = 32'hc404487;
      8500: inst = 32'h8220000;
      8501: inst = 32'h10408000;
      8502: inst = 32'hc404488;
      8503: inst = 32'h8220000;
      8504: inst = 32'h10408000;
      8505: inst = 32'hc404489;
      8506: inst = 32'h8220000;
      8507: inst = 32'h10408000;
      8508: inst = 32'hc40448a;
      8509: inst = 32'h8220000;
      8510: inst = 32'h10408000;
      8511: inst = 32'hc40448b;
      8512: inst = 32'h8220000;
      8513: inst = 32'h10408000;
      8514: inst = 32'hc40448c;
      8515: inst = 32'h8220000;
      8516: inst = 32'h10408000;
      8517: inst = 32'hc40448d;
      8518: inst = 32'h8220000;
      8519: inst = 32'h10408000;
      8520: inst = 32'hc40448e;
      8521: inst = 32'h8220000;
      8522: inst = 32'h10408000;
      8523: inst = 32'hc40448f;
      8524: inst = 32'h8220000;
      8525: inst = 32'h10408000;
      8526: inst = 32'hc404490;
      8527: inst = 32'h8220000;
      8528: inst = 32'h10408000;
      8529: inst = 32'hc404491;
      8530: inst = 32'h8220000;
      8531: inst = 32'h10408000;
      8532: inst = 32'hc404492;
      8533: inst = 32'h8220000;
      8534: inst = 32'h10408000;
      8535: inst = 32'hc404493;
      8536: inst = 32'h8220000;
      8537: inst = 32'h10408000;
      8538: inst = 32'hc404494;
      8539: inst = 32'h8220000;
      8540: inst = 32'h10408000;
      8541: inst = 32'hc404495;
      8542: inst = 32'h8220000;
      8543: inst = 32'h10408000;
      8544: inst = 32'hc404496;
      8545: inst = 32'h8220000;
      8546: inst = 32'h10408000;
      8547: inst = 32'hc404497;
      8548: inst = 32'h8220000;
      8549: inst = 32'h10408000;
      8550: inst = 32'hc404498;
      8551: inst = 32'h8220000;
      8552: inst = 32'h10408000;
      8553: inst = 32'hc404499;
      8554: inst = 32'h8220000;
      8555: inst = 32'h10408000;
      8556: inst = 32'hc40449a;
      8557: inst = 32'h8220000;
      8558: inst = 32'h10408000;
      8559: inst = 32'hc40449b;
      8560: inst = 32'h8220000;
      8561: inst = 32'h10408000;
      8562: inst = 32'hc40449c;
      8563: inst = 32'h8220000;
      8564: inst = 32'h10408000;
      8565: inst = 32'hc40449d;
      8566: inst = 32'h8220000;
      8567: inst = 32'h10408000;
      8568: inst = 32'hc40449e;
      8569: inst = 32'h8220000;
      8570: inst = 32'h10408000;
      8571: inst = 32'hc40449f;
      8572: inst = 32'h8220000;
      8573: inst = 32'h10408000;
      8574: inst = 32'hc4044a0;
      8575: inst = 32'h8220000;
      8576: inst = 32'h10408000;
      8577: inst = 32'hc4044a1;
      8578: inst = 32'h8220000;
      8579: inst = 32'h10408000;
      8580: inst = 32'hc4044a2;
      8581: inst = 32'h8220000;
      8582: inst = 32'h10408000;
      8583: inst = 32'hc4044a3;
      8584: inst = 32'h8220000;
      8585: inst = 32'h10408000;
      8586: inst = 32'hc4044dc;
      8587: inst = 32'h8220000;
      8588: inst = 32'h10408000;
      8589: inst = 32'hc4044dd;
      8590: inst = 32'h8220000;
      8591: inst = 32'h10408000;
      8592: inst = 32'hc4044de;
      8593: inst = 32'h8220000;
      8594: inst = 32'h10408000;
      8595: inst = 32'hc4044df;
      8596: inst = 32'h8220000;
      8597: inst = 32'h10408000;
      8598: inst = 32'hc4044e0;
      8599: inst = 32'h8220000;
      8600: inst = 32'h10408000;
      8601: inst = 32'hc4044e1;
      8602: inst = 32'h8220000;
      8603: inst = 32'h10408000;
      8604: inst = 32'hc4044e2;
      8605: inst = 32'h8220000;
      8606: inst = 32'h10408000;
      8607: inst = 32'hc4044e3;
      8608: inst = 32'h8220000;
      8609: inst = 32'h10408000;
      8610: inst = 32'hc4044e4;
      8611: inst = 32'h8220000;
      8612: inst = 32'h10408000;
      8613: inst = 32'hc4044e5;
      8614: inst = 32'h8220000;
      8615: inst = 32'h10408000;
      8616: inst = 32'hc4044e6;
      8617: inst = 32'h8220000;
      8618: inst = 32'h10408000;
      8619: inst = 32'hc4044e7;
      8620: inst = 32'h8220000;
      8621: inst = 32'h10408000;
      8622: inst = 32'hc4044e8;
      8623: inst = 32'h8220000;
      8624: inst = 32'h10408000;
      8625: inst = 32'hc4044e9;
      8626: inst = 32'h8220000;
      8627: inst = 32'h10408000;
      8628: inst = 32'hc4044ea;
      8629: inst = 32'h8220000;
      8630: inst = 32'h10408000;
      8631: inst = 32'hc4044eb;
      8632: inst = 32'h8220000;
      8633: inst = 32'h10408000;
      8634: inst = 32'hc4044ec;
      8635: inst = 32'h8220000;
      8636: inst = 32'h10408000;
      8637: inst = 32'hc4044ed;
      8638: inst = 32'h8220000;
      8639: inst = 32'h10408000;
      8640: inst = 32'hc4044ee;
      8641: inst = 32'h8220000;
      8642: inst = 32'h10408000;
      8643: inst = 32'hc4044ef;
      8644: inst = 32'h8220000;
      8645: inst = 32'h10408000;
      8646: inst = 32'hc4044f0;
      8647: inst = 32'h8220000;
      8648: inst = 32'h10408000;
      8649: inst = 32'hc4044f1;
      8650: inst = 32'h8220000;
      8651: inst = 32'h10408000;
      8652: inst = 32'hc4044f2;
      8653: inst = 32'h8220000;
      8654: inst = 32'h10408000;
      8655: inst = 32'hc4044f3;
      8656: inst = 32'h8220000;
      8657: inst = 32'h10408000;
      8658: inst = 32'hc4044f4;
      8659: inst = 32'h8220000;
      8660: inst = 32'h10408000;
      8661: inst = 32'hc4044f5;
      8662: inst = 32'h8220000;
      8663: inst = 32'h10408000;
      8664: inst = 32'hc4044f6;
      8665: inst = 32'h8220000;
      8666: inst = 32'h10408000;
      8667: inst = 32'hc4044f7;
      8668: inst = 32'h8220000;
      8669: inst = 32'h10408000;
      8670: inst = 32'hc4044f8;
      8671: inst = 32'h8220000;
      8672: inst = 32'h10408000;
      8673: inst = 32'hc4044f9;
      8674: inst = 32'h8220000;
      8675: inst = 32'h10408000;
      8676: inst = 32'hc4044fa;
      8677: inst = 32'h8220000;
      8678: inst = 32'h10408000;
      8679: inst = 32'hc4044fb;
      8680: inst = 32'h8220000;
      8681: inst = 32'h10408000;
      8682: inst = 32'hc4044fc;
      8683: inst = 32'h8220000;
      8684: inst = 32'h10408000;
      8685: inst = 32'hc4044fd;
      8686: inst = 32'h8220000;
      8687: inst = 32'h10408000;
      8688: inst = 32'hc4044fe;
      8689: inst = 32'h8220000;
      8690: inst = 32'h10408000;
      8691: inst = 32'hc4044ff;
      8692: inst = 32'h8220000;
      8693: inst = 32'h10408000;
      8694: inst = 32'hc404500;
      8695: inst = 32'h8220000;
      8696: inst = 32'h10408000;
      8697: inst = 32'hc404501;
      8698: inst = 32'h8220000;
      8699: inst = 32'h10408000;
      8700: inst = 32'hc404502;
      8701: inst = 32'h8220000;
      8702: inst = 32'h10408000;
      8703: inst = 32'hc404503;
      8704: inst = 32'h8220000;
      8705: inst = 32'h10408000;
      8706: inst = 32'hc40453c;
      8707: inst = 32'h8220000;
      8708: inst = 32'h10408000;
      8709: inst = 32'hc40453d;
      8710: inst = 32'h8220000;
      8711: inst = 32'h10408000;
      8712: inst = 32'hc40453e;
      8713: inst = 32'h8220000;
      8714: inst = 32'h10408000;
      8715: inst = 32'hc40453f;
      8716: inst = 32'h8220000;
      8717: inst = 32'h10408000;
      8718: inst = 32'hc404540;
      8719: inst = 32'h8220000;
      8720: inst = 32'h10408000;
      8721: inst = 32'hc404541;
      8722: inst = 32'h8220000;
      8723: inst = 32'h10408000;
      8724: inst = 32'hc404542;
      8725: inst = 32'h8220000;
      8726: inst = 32'h10408000;
      8727: inst = 32'hc404543;
      8728: inst = 32'h8220000;
      8729: inst = 32'h10408000;
      8730: inst = 32'hc404544;
      8731: inst = 32'h8220000;
      8732: inst = 32'h10408000;
      8733: inst = 32'hc404545;
      8734: inst = 32'h8220000;
      8735: inst = 32'h10408000;
      8736: inst = 32'hc404546;
      8737: inst = 32'h8220000;
      8738: inst = 32'h10408000;
      8739: inst = 32'hc404547;
      8740: inst = 32'h8220000;
      8741: inst = 32'h10408000;
      8742: inst = 32'hc404548;
      8743: inst = 32'h8220000;
      8744: inst = 32'h10408000;
      8745: inst = 32'hc404549;
      8746: inst = 32'h8220000;
      8747: inst = 32'h10408000;
      8748: inst = 32'hc40454a;
      8749: inst = 32'h8220000;
      8750: inst = 32'h10408000;
      8751: inst = 32'hc40454b;
      8752: inst = 32'h8220000;
      8753: inst = 32'h10408000;
      8754: inst = 32'hc40454c;
      8755: inst = 32'h8220000;
      8756: inst = 32'h10408000;
      8757: inst = 32'hc40454d;
      8758: inst = 32'h8220000;
      8759: inst = 32'h10408000;
      8760: inst = 32'hc40454e;
      8761: inst = 32'h8220000;
      8762: inst = 32'h10408000;
      8763: inst = 32'hc40454f;
      8764: inst = 32'h8220000;
      8765: inst = 32'h10408000;
      8766: inst = 32'hc404550;
      8767: inst = 32'h8220000;
      8768: inst = 32'h10408000;
      8769: inst = 32'hc404551;
      8770: inst = 32'h8220000;
      8771: inst = 32'h10408000;
      8772: inst = 32'hc404552;
      8773: inst = 32'h8220000;
      8774: inst = 32'h10408000;
      8775: inst = 32'hc404553;
      8776: inst = 32'h8220000;
      8777: inst = 32'h10408000;
      8778: inst = 32'hc404554;
      8779: inst = 32'h8220000;
      8780: inst = 32'h10408000;
      8781: inst = 32'hc404555;
      8782: inst = 32'h8220000;
      8783: inst = 32'h10408000;
      8784: inst = 32'hc404556;
      8785: inst = 32'h8220000;
      8786: inst = 32'h10408000;
      8787: inst = 32'hc404557;
      8788: inst = 32'h8220000;
      8789: inst = 32'h10408000;
      8790: inst = 32'hc404558;
      8791: inst = 32'h8220000;
      8792: inst = 32'h10408000;
      8793: inst = 32'hc404559;
      8794: inst = 32'h8220000;
      8795: inst = 32'h10408000;
      8796: inst = 32'hc40455a;
      8797: inst = 32'h8220000;
      8798: inst = 32'h10408000;
      8799: inst = 32'hc40455b;
      8800: inst = 32'h8220000;
      8801: inst = 32'h10408000;
      8802: inst = 32'hc40455c;
      8803: inst = 32'h8220000;
      8804: inst = 32'h10408000;
      8805: inst = 32'hc40455d;
      8806: inst = 32'h8220000;
      8807: inst = 32'h10408000;
      8808: inst = 32'hc40455e;
      8809: inst = 32'h8220000;
      8810: inst = 32'h10408000;
      8811: inst = 32'hc40455f;
      8812: inst = 32'h8220000;
      8813: inst = 32'h10408000;
      8814: inst = 32'hc404560;
      8815: inst = 32'h8220000;
      8816: inst = 32'h10408000;
      8817: inst = 32'hc404561;
      8818: inst = 32'h8220000;
      8819: inst = 32'h10408000;
      8820: inst = 32'hc404562;
      8821: inst = 32'h8220000;
      8822: inst = 32'h10408000;
      8823: inst = 32'hc404563;
      8824: inst = 32'h8220000;
      8825: inst = 32'h10408000;
      8826: inst = 32'hc40459c;
      8827: inst = 32'h8220000;
      8828: inst = 32'h10408000;
      8829: inst = 32'hc40459d;
      8830: inst = 32'h8220000;
      8831: inst = 32'h10408000;
      8832: inst = 32'hc40459e;
      8833: inst = 32'h8220000;
      8834: inst = 32'h10408000;
      8835: inst = 32'hc40459f;
      8836: inst = 32'h8220000;
      8837: inst = 32'h10408000;
      8838: inst = 32'hc4045a0;
      8839: inst = 32'h8220000;
      8840: inst = 32'h10408000;
      8841: inst = 32'hc4045a1;
      8842: inst = 32'h8220000;
      8843: inst = 32'h10408000;
      8844: inst = 32'hc4045a2;
      8845: inst = 32'h8220000;
      8846: inst = 32'h10408000;
      8847: inst = 32'hc4045a3;
      8848: inst = 32'h8220000;
      8849: inst = 32'h10408000;
      8850: inst = 32'hc4045a4;
      8851: inst = 32'h8220000;
      8852: inst = 32'h10408000;
      8853: inst = 32'hc4045a5;
      8854: inst = 32'h8220000;
      8855: inst = 32'h10408000;
      8856: inst = 32'hc4045a6;
      8857: inst = 32'h8220000;
      8858: inst = 32'h10408000;
      8859: inst = 32'hc4045a7;
      8860: inst = 32'h8220000;
      8861: inst = 32'h10408000;
      8862: inst = 32'hc4045a8;
      8863: inst = 32'h8220000;
      8864: inst = 32'h10408000;
      8865: inst = 32'hc4045a9;
      8866: inst = 32'h8220000;
      8867: inst = 32'h10408000;
      8868: inst = 32'hc4045aa;
      8869: inst = 32'h8220000;
      8870: inst = 32'h10408000;
      8871: inst = 32'hc4045ab;
      8872: inst = 32'h8220000;
      8873: inst = 32'h10408000;
      8874: inst = 32'hc4045ac;
      8875: inst = 32'h8220000;
      8876: inst = 32'h10408000;
      8877: inst = 32'hc4045ad;
      8878: inst = 32'h8220000;
      8879: inst = 32'h10408000;
      8880: inst = 32'hc4045ae;
      8881: inst = 32'h8220000;
      8882: inst = 32'h10408000;
      8883: inst = 32'hc4045af;
      8884: inst = 32'h8220000;
      8885: inst = 32'h10408000;
      8886: inst = 32'hc4045b0;
      8887: inst = 32'h8220000;
      8888: inst = 32'h10408000;
      8889: inst = 32'hc4045b1;
      8890: inst = 32'h8220000;
      8891: inst = 32'h10408000;
      8892: inst = 32'hc4045b2;
      8893: inst = 32'h8220000;
      8894: inst = 32'h10408000;
      8895: inst = 32'hc4045b3;
      8896: inst = 32'h8220000;
      8897: inst = 32'h10408000;
      8898: inst = 32'hc4045b4;
      8899: inst = 32'h8220000;
      8900: inst = 32'h10408000;
      8901: inst = 32'hc4045b5;
      8902: inst = 32'h8220000;
      8903: inst = 32'h10408000;
      8904: inst = 32'hc4045b6;
      8905: inst = 32'h8220000;
      8906: inst = 32'h10408000;
      8907: inst = 32'hc4045b7;
      8908: inst = 32'h8220000;
      8909: inst = 32'h10408000;
      8910: inst = 32'hc4045b8;
      8911: inst = 32'h8220000;
      8912: inst = 32'h10408000;
      8913: inst = 32'hc4045b9;
      8914: inst = 32'h8220000;
      8915: inst = 32'h10408000;
      8916: inst = 32'hc4045ba;
      8917: inst = 32'h8220000;
      8918: inst = 32'h10408000;
      8919: inst = 32'hc4045bb;
      8920: inst = 32'h8220000;
      8921: inst = 32'h10408000;
      8922: inst = 32'hc4045bc;
      8923: inst = 32'h8220000;
      8924: inst = 32'h10408000;
      8925: inst = 32'hc4045bd;
      8926: inst = 32'h8220000;
      8927: inst = 32'h10408000;
      8928: inst = 32'hc4045be;
      8929: inst = 32'h8220000;
      8930: inst = 32'h10408000;
      8931: inst = 32'hc4045bf;
      8932: inst = 32'h8220000;
      8933: inst = 32'h10408000;
      8934: inst = 32'hc4045c0;
      8935: inst = 32'h8220000;
      8936: inst = 32'h10408000;
      8937: inst = 32'hc4045c1;
      8938: inst = 32'h8220000;
      8939: inst = 32'h10408000;
      8940: inst = 32'hc4045c2;
      8941: inst = 32'h8220000;
      8942: inst = 32'h10408000;
      8943: inst = 32'hc4045c3;
      8944: inst = 32'h8220000;
      8945: inst = 32'h10408000;
      8946: inst = 32'hc4045fc;
      8947: inst = 32'h8220000;
      8948: inst = 32'h10408000;
      8949: inst = 32'hc4045fd;
      8950: inst = 32'h8220000;
      8951: inst = 32'h10408000;
      8952: inst = 32'hc4045fe;
      8953: inst = 32'h8220000;
      8954: inst = 32'h10408000;
      8955: inst = 32'hc4045ff;
      8956: inst = 32'h8220000;
      8957: inst = 32'h10408000;
      8958: inst = 32'hc404600;
      8959: inst = 32'h8220000;
      8960: inst = 32'h10408000;
      8961: inst = 32'hc404601;
      8962: inst = 32'h8220000;
      8963: inst = 32'h10408000;
      8964: inst = 32'hc404602;
      8965: inst = 32'h8220000;
      8966: inst = 32'h10408000;
      8967: inst = 32'hc404603;
      8968: inst = 32'h8220000;
      8969: inst = 32'h10408000;
      8970: inst = 32'hc404604;
      8971: inst = 32'h8220000;
      8972: inst = 32'h10408000;
      8973: inst = 32'hc404605;
      8974: inst = 32'h8220000;
      8975: inst = 32'h10408000;
      8976: inst = 32'hc404606;
      8977: inst = 32'h8220000;
      8978: inst = 32'h10408000;
      8979: inst = 32'hc404607;
      8980: inst = 32'h8220000;
      8981: inst = 32'h10408000;
      8982: inst = 32'hc404608;
      8983: inst = 32'h8220000;
      8984: inst = 32'h10408000;
      8985: inst = 32'hc404609;
      8986: inst = 32'h8220000;
      8987: inst = 32'h10408000;
      8988: inst = 32'hc40460a;
      8989: inst = 32'h8220000;
      8990: inst = 32'h10408000;
      8991: inst = 32'hc40460b;
      8992: inst = 32'h8220000;
      8993: inst = 32'h10408000;
      8994: inst = 32'hc40460c;
      8995: inst = 32'h8220000;
      8996: inst = 32'h10408000;
      8997: inst = 32'hc40460d;
      8998: inst = 32'h8220000;
      8999: inst = 32'h10408000;
      9000: inst = 32'hc40460e;
      9001: inst = 32'h8220000;
      9002: inst = 32'h10408000;
      9003: inst = 32'hc40460f;
      9004: inst = 32'h8220000;
      9005: inst = 32'h10408000;
      9006: inst = 32'hc404610;
      9007: inst = 32'h8220000;
      9008: inst = 32'h10408000;
      9009: inst = 32'hc404611;
      9010: inst = 32'h8220000;
      9011: inst = 32'h10408000;
      9012: inst = 32'hc404612;
      9013: inst = 32'h8220000;
      9014: inst = 32'h10408000;
      9015: inst = 32'hc404613;
      9016: inst = 32'h8220000;
      9017: inst = 32'h10408000;
      9018: inst = 32'hc404614;
      9019: inst = 32'h8220000;
      9020: inst = 32'h10408000;
      9021: inst = 32'hc404615;
      9022: inst = 32'h8220000;
      9023: inst = 32'h10408000;
      9024: inst = 32'hc404616;
      9025: inst = 32'h8220000;
      9026: inst = 32'h10408000;
      9027: inst = 32'hc404617;
      9028: inst = 32'h8220000;
      9029: inst = 32'h10408000;
      9030: inst = 32'hc404618;
      9031: inst = 32'h8220000;
      9032: inst = 32'h10408000;
      9033: inst = 32'hc404619;
      9034: inst = 32'h8220000;
      9035: inst = 32'h10408000;
      9036: inst = 32'hc40461a;
      9037: inst = 32'h8220000;
      9038: inst = 32'h10408000;
      9039: inst = 32'hc40461b;
      9040: inst = 32'h8220000;
      9041: inst = 32'h10408000;
      9042: inst = 32'hc40461c;
      9043: inst = 32'h8220000;
      9044: inst = 32'h10408000;
      9045: inst = 32'hc40461d;
      9046: inst = 32'h8220000;
      9047: inst = 32'h10408000;
      9048: inst = 32'hc40461e;
      9049: inst = 32'h8220000;
      9050: inst = 32'h10408000;
      9051: inst = 32'hc40461f;
      9052: inst = 32'h8220000;
      9053: inst = 32'h10408000;
      9054: inst = 32'hc404620;
      9055: inst = 32'h8220000;
      9056: inst = 32'h10408000;
      9057: inst = 32'hc404621;
      9058: inst = 32'h8220000;
      9059: inst = 32'h10408000;
      9060: inst = 32'hc404622;
      9061: inst = 32'h8220000;
      9062: inst = 32'h10408000;
      9063: inst = 32'hc404623;
      9064: inst = 32'h8220000;
      9065: inst = 32'h10408000;
      9066: inst = 32'hc40465c;
      9067: inst = 32'h8220000;
      9068: inst = 32'h10408000;
      9069: inst = 32'hc40465d;
      9070: inst = 32'h8220000;
      9071: inst = 32'h10408000;
      9072: inst = 32'hc40465e;
      9073: inst = 32'h8220000;
      9074: inst = 32'h10408000;
      9075: inst = 32'hc40465f;
      9076: inst = 32'h8220000;
      9077: inst = 32'h10408000;
      9078: inst = 32'hc404660;
      9079: inst = 32'h8220000;
      9080: inst = 32'h10408000;
      9081: inst = 32'hc404661;
      9082: inst = 32'h8220000;
      9083: inst = 32'h10408000;
      9084: inst = 32'hc404662;
      9085: inst = 32'h8220000;
      9086: inst = 32'h10408000;
      9087: inst = 32'hc404663;
      9088: inst = 32'h8220000;
      9089: inst = 32'h10408000;
      9090: inst = 32'hc404664;
      9091: inst = 32'h8220000;
      9092: inst = 32'h10408000;
      9093: inst = 32'hc404665;
      9094: inst = 32'h8220000;
      9095: inst = 32'h10408000;
      9096: inst = 32'hc404666;
      9097: inst = 32'h8220000;
      9098: inst = 32'h10408000;
      9099: inst = 32'hc404667;
      9100: inst = 32'h8220000;
      9101: inst = 32'h10408000;
      9102: inst = 32'hc404668;
      9103: inst = 32'h8220000;
      9104: inst = 32'h10408000;
      9105: inst = 32'hc404669;
      9106: inst = 32'h8220000;
      9107: inst = 32'h10408000;
      9108: inst = 32'hc40466a;
      9109: inst = 32'h8220000;
      9110: inst = 32'h10408000;
      9111: inst = 32'hc40466b;
      9112: inst = 32'h8220000;
      9113: inst = 32'h10408000;
      9114: inst = 32'hc40466c;
      9115: inst = 32'h8220000;
      9116: inst = 32'h10408000;
      9117: inst = 32'hc40466d;
      9118: inst = 32'h8220000;
      9119: inst = 32'h10408000;
      9120: inst = 32'hc40466e;
      9121: inst = 32'h8220000;
      9122: inst = 32'h10408000;
      9123: inst = 32'hc40466f;
      9124: inst = 32'h8220000;
      9125: inst = 32'h10408000;
      9126: inst = 32'hc404670;
      9127: inst = 32'h8220000;
      9128: inst = 32'h10408000;
      9129: inst = 32'hc404671;
      9130: inst = 32'h8220000;
      9131: inst = 32'h10408000;
      9132: inst = 32'hc404672;
      9133: inst = 32'h8220000;
      9134: inst = 32'h10408000;
      9135: inst = 32'hc404673;
      9136: inst = 32'h8220000;
      9137: inst = 32'h10408000;
      9138: inst = 32'hc404674;
      9139: inst = 32'h8220000;
      9140: inst = 32'h10408000;
      9141: inst = 32'hc404675;
      9142: inst = 32'h8220000;
      9143: inst = 32'h10408000;
      9144: inst = 32'hc404676;
      9145: inst = 32'h8220000;
      9146: inst = 32'h10408000;
      9147: inst = 32'hc404677;
      9148: inst = 32'h8220000;
      9149: inst = 32'h10408000;
      9150: inst = 32'hc404678;
      9151: inst = 32'h8220000;
      9152: inst = 32'h10408000;
      9153: inst = 32'hc404679;
      9154: inst = 32'h8220000;
      9155: inst = 32'h10408000;
      9156: inst = 32'hc40467a;
      9157: inst = 32'h8220000;
      9158: inst = 32'h10408000;
      9159: inst = 32'hc40467b;
      9160: inst = 32'h8220000;
      9161: inst = 32'h10408000;
      9162: inst = 32'hc40467c;
      9163: inst = 32'h8220000;
      9164: inst = 32'h10408000;
      9165: inst = 32'hc40467d;
      9166: inst = 32'h8220000;
      9167: inst = 32'h10408000;
      9168: inst = 32'hc40467e;
      9169: inst = 32'h8220000;
      9170: inst = 32'h10408000;
      9171: inst = 32'hc40467f;
      9172: inst = 32'h8220000;
      9173: inst = 32'h10408000;
      9174: inst = 32'hc404680;
      9175: inst = 32'h8220000;
      9176: inst = 32'h10408000;
      9177: inst = 32'hc404681;
      9178: inst = 32'h8220000;
      9179: inst = 32'h10408000;
      9180: inst = 32'hc404682;
      9181: inst = 32'h8220000;
      9182: inst = 32'h10408000;
      9183: inst = 32'hc404683;
      9184: inst = 32'h8220000;
      9185: inst = 32'h10408000;
      9186: inst = 32'hc4046bc;
      9187: inst = 32'h8220000;
      9188: inst = 32'h10408000;
      9189: inst = 32'hc4046bd;
      9190: inst = 32'h8220000;
      9191: inst = 32'h10408000;
      9192: inst = 32'hc4046be;
      9193: inst = 32'h8220000;
      9194: inst = 32'h10408000;
      9195: inst = 32'hc4046bf;
      9196: inst = 32'h8220000;
      9197: inst = 32'h10408000;
      9198: inst = 32'hc4046c0;
      9199: inst = 32'h8220000;
      9200: inst = 32'h10408000;
      9201: inst = 32'hc4046c1;
      9202: inst = 32'h8220000;
      9203: inst = 32'h10408000;
      9204: inst = 32'hc4046c2;
      9205: inst = 32'h8220000;
      9206: inst = 32'h10408000;
      9207: inst = 32'hc4046c3;
      9208: inst = 32'h8220000;
      9209: inst = 32'h10408000;
      9210: inst = 32'hc4046c4;
      9211: inst = 32'h8220000;
      9212: inst = 32'h10408000;
      9213: inst = 32'hc4046c5;
      9214: inst = 32'h8220000;
      9215: inst = 32'h10408000;
      9216: inst = 32'hc4046c6;
      9217: inst = 32'h8220000;
      9218: inst = 32'h10408000;
      9219: inst = 32'hc4046c7;
      9220: inst = 32'h8220000;
      9221: inst = 32'h10408000;
      9222: inst = 32'hc4046c8;
      9223: inst = 32'h8220000;
      9224: inst = 32'h10408000;
      9225: inst = 32'hc4046c9;
      9226: inst = 32'h8220000;
      9227: inst = 32'h10408000;
      9228: inst = 32'hc4046ca;
      9229: inst = 32'h8220000;
      9230: inst = 32'h10408000;
      9231: inst = 32'hc4046cb;
      9232: inst = 32'h8220000;
      9233: inst = 32'h10408000;
      9234: inst = 32'hc4046cc;
      9235: inst = 32'h8220000;
      9236: inst = 32'h10408000;
      9237: inst = 32'hc4046cd;
      9238: inst = 32'h8220000;
      9239: inst = 32'h10408000;
      9240: inst = 32'hc4046ce;
      9241: inst = 32'h8220000;
      9242: inst = 32'h10408000;
      9243: inst = 32'hc4046cf;
      9244: inst = 32'h8220000;
      9245: inst = 32'h10408000;
      9246: inst = 32'hc4046d0;
      9247: inst = 32'h8220000;
      9248: inst = 32'h10408000;
      9249: inst = 32'hc4046d1;
      9250: inst = 32'h8220000;
      9251: inst = 32'h10408000;
      9252: inst = 32'hc4046d2;
      9253: inst = 32'h8220000;
      9254: inst = 32'h10408000;
      9255: inst = 32'hc4046d3;
      9256: inst = 32'h8220000;
      9257: inst = 32'h10408000;
      9258: inst = 32'hc4046d4;
      9259: inst = 32'h8220000;
      9260: inst = 32'h10408000;
      9261: inst = 32'hc4046d5;
      9262: inst = 32'h8220000;
      9263: inst = 32'h10408000;
      9264: inst = 32'hc4046d6;
      9265: inst = 32'h8220000;
      9266: inst = 32'h10408000;
      9267: inst = 32'hc4046d7;
      9268: inst = 32'h8220000;
      9269: inst = 32'h10408000;
      9270: inst = 32'hc4046d8;
      9271: inst = 32'h8220000;
      9272: inst = 32'h10408000;
      9273: inst = 32'hc4046d9;
      9274: inst = 32'h8220000;
      9275: inst = 32'h10408000;
      9276: inst = 32'hc4046da;
      9277: inst = 32'h8220000;
      9278: inst = 32'h10408000;
      9279: inst = 32'hc4046db;
      9280: inst = 32'h8220000;
      9281: inst = 32'h10408000;
      9282: inst = 32'hc4046dc;
      9283: inst = 32'h8220000;
      9284: inst = 32'h10408000;
      9285: inst = 32'hc4046dd;
      9286: inst = 32'h8220000;
      9287: inst = 32'h10408000;
      9288: inst = 32'hc4046de;
      9289: inst = 32'h8220000;
      9290: inst = 32'h10408000;
      9291: inst = 32'hc4046df;
      9292: inst = 32'h8220000;
      9293: inst = 32'h10408000;
      9294: inst = 32'hc4046e0;
      9295: inst = 32'h8220000;
      9296: inst = 32'h10408000;
      9297: inst = 32'hc4046e1;
      9298: inst = 32'h8220000;
      9299: inst = 32'h10408000;
      9300: inst = 32'hc4046e2;
      9301: inst = 32'h8220000;
      9302: inst = 32'h10408000;
      9303: inst = 32'hc4046e3;
      9304: inst = 32'h8220000;
      9305: inst = 32'h10408000;
      9306: inst = 32'hc40471c;
      9307: inst = 32'h8220000;
      9308: inst = 32'h10408000;
      9309: inst = 32'hc40471d;
      9310: inst = 32'h8220000;
      9311: inst = 32'h10408000;
      9312: inst = 32'hc40471e;
      9313: inst = 32'h8220000;
      9314: inst = 32'h10408000;
      9315: inst = 32'hc40471f;
      9316: inst = 32'h8220000;
      9317: inst = 32'h10408000;
      9318: inst = 32'hc404720;
      9319: inst = 32'h8220000;
      9320: inst = 32'h10408000;
      9321: inst = 32'hc404721;
      9322: inst = 32'h8220000;
      9323: inst = 32'h10408000;
      9324: inst = 32'hc404722;
      9325: inst = 32'h8220000;
      9326: inst = 32'h10408000;
      9327: inst = 32'hc404723;
      9328: inst = 32'h8220000;
      9329: inst = 32'h10408000;
      9330: inst = 32'hc404724;
      9331: inst = 32'h8220000;
      9332: inst = 32'h10408000;
      9333: inst = 32'hc404725;
      9334: inst = 32'h8220000;
      9335: inst = 32'h10408000;
      9336: inst = 32'hc404726;
      9337: inst = 32'h8220000;
      9338: inst = 32'h10408000;
      9339: inst = 32'hc404727;
      9340: inst = 32'h8220000;
      9341: inst = 32'h10408000;
      9342: inst = 32'hc404728;
      9343: inst = 32'h8220000;
      9344: inst = 32'h10408000;
      9345: inst = 32'hc404729;
      9346: inst = 32'h8220000;
      9347: inst = 32'h10408000;
      9348: inst = 32'hc40472a;
      9349: inst = 32'h8220000;
      9350: inst = 32'h10408000;
      9351: inst = 32'hc40472b;
      9352: inst = 32'h8220000;
      9353: inst = 32'h10408000;
      9354: inst = 32'hc40472c;
      9355: inst = 32'h8220000;
      9356: inst = 32'h10408000;
      9357: inst = 32'hc40472d;
      9358: inst = 32'h8220000;
      9359: inst = 32'h10408000;
      9360: inst = 32'hc40472e;
      9361: inst = 32'h8220000;
      9362: inst = 32'h10408000;
      9363: inst = 32'hc40472f;
      9364: inst = 32'h8220000;
      9365: inst = 32'h10408000;
      9366: inst = 32'hc404730;
      9367: inst = 32'h8220000;
      9368: inst = 32'h10408000;
      9369: inst = 32'hc404731;
      9370: inst = 32'h8220000;
      9371: inst = 32'h10408000;
      9372: inst = 32'hc404732;
      9373: inst = 32'h8220000;
      9374: inst = 32'h10408000;
      9375: inst = 32'hc404733;
      9376: inst = 32'h8220000;
      9377: inst = 32'h10408000;
      9378: inst = 32'hc404734;
      9379: inst = 32'h8220000;
      9380: inst = 32'h10408000;
      9381: inst = 32'hc404735;
      9382: inst = 32'h8220000;
      9383: inst = 32'h10408000;
      9384: inst = 32'hc404736;
      9385: inst = 32'h8220000;
      9386: inst = 32'h10408000;
      9387: inst = 32'hc404737;
      9388: inst = 32'h8220000;
      9389: inst = 32'h10408000;
      9390: inst = 32'hc404738;
      9391: inst = 32'h8220000;
      9392: inst = 32'h10408000;
      9393: inst = 32'hc404739;
      9394: inst = 32'h8220000;
      9395: inst = 32'h10408000;
      9396: inst = 32'hc40473a;
      9397: inst = 32'h8220000;
      9398: inst = 32'h10408000;
      9399: inst = 32'hc40473b;
      9400: inst = 32'h8220000;
      9401: inst = 32'h10408000;
      9402: inst = 32'hc40473c;
      9403: inst = 32'h8220000;
      9404: inst = 32'h10408000;
      9405: inst = 32'hc40473d;
      9406: inst = 32'h8220000;
      9407: inst = 32'h10408000;
      9408: inst = 32'hc40473e;
      9409: inst = 32'h8220000;
      9410: inst = 32'h10408000;
      9411: inst = 32'hc40473f;
      9412: inst = 32'h8220000;
      9413: inst = 32'h10408000;
      9414: inst = 32'hc404740;
      9415: inst = 32'h8220000;
      9416: inst = 32'h10408000;
      9417: inst = 32'hc404741;
      9418: inst = 32'h8220000;
      9419: inst = 32'h10408000;
      9420: inst = 32'hc404742;
      9421: inst = 32'h8220000;
      9422: inst = 32'h10408000;
      9423: inst = 32'hc404743;
      9424: inst = 32'h8220000;
      9425: inst = 32'h10408000;
      9426: inst = 32'hc40477c;
      9427: inst = 32'h8220000;
      9428: inst = 32'h10408000;
      9429: inst = 32'hc40477d;
      9430: inst = 32'h8220000;
      9431: inst = 32'h10408000;
      9432: inst = 32'hc40477e;
      9433: inst = 32'h8220000;
      9434: inst = 32'h10408000;
      9435: inst = 32'hc40477f;
      9436: inst = 32'h8220000;
      9437: inst = 32'h10408000;
      9438: inst = 32'hc404780;
      9439: inst = 32'h8220000;
      9440: inst = 32'h10408000;
      9441: inst = 32'hc404781;
      9442: inst = 32'h8220000;
      9443: inst = 32'h10408000;
      9444: inst = 32'hc404782;
      9445: inst = 32'h8220000;
      9446: inst = 32'h10408000;
      9447: inst = 32'hc404783;
      9448: inst = 32'h8220000;
      9449: inst = 32'h10408000;
      9450: inst = 32'hc404784;
      9451: inst = 32'h8220000;
      9452: inst = 32'h10408000;
      9453: inst = 32'hc404785;
      9454: inst = 32'h8220000;
      9455: inst = 32'h10408000;
      9456: inst = 32'hc404786;
      9457: inst = 32'h8220000;
      9458: inst = 32'h10408000;
      9459: inst = 32'hc404787;
      9460: inst = 32'h8220000;
      9461: inst = 32'h10408000;
      9462: inst = 32'hc404788;
      9463: inst = 32'h8220000;
      9464: inst = 32'h10408000;
      9465: inst = 32'hc404789;
      9466: inst = 32'h8220000;
      9467: inst = 32'h10408000;
      9468: inst = 32'hc40478a;
      9469: inst = 32'h8220000;
      9470: inst = 32'h10408000;
      9471: inst = 32'hc40478b;
      9472: inst = 32'h8220000;
      9473: inst = 32'h10408000;
      9474: inst = 32'hc40478c;
      9475: inst = 32'h8220000;
      9476: inst = 32'h10408000;
      9477: inst = 32'hc40478d;
      9478: inst = 32'h8220000;
      9479: inst = 32'h10408000;
      9480: inst = 32'hc40478e;
      9481: inst = 32'h8220000;
      9482: inst = 32'h10408000;
      9483: inst = 32'hc40478f;
      9484: inst = 32'h8220000;
      9485: inst = 32'h10408000;
      9486: inst = 32'hc404790;
      9487: inst = 32'h8220000;
      9488: inst = 32'h10408000;
      9489: inst = 32'hc404791;
      9490: inst = 32'h8220000;
      9491: inst = 32'h10408000;
      9492: inst = 32'hc404792;
      9493: inst = 32'h8220000;
      9494: inst = 32'h10408000;
      9495: inst = 32'hc404793;
      9496: inst = 32'h8220000;
      9497: inst = 32'h10408000;
      9498: inst = 32'hc404794;
      9499: inst = 32'h8220000;
      9500: inst = 32'h10408000;
      9501: inst = 32'hc404795;
      9502: inst = 32'h8220000;
      9503: inst = 32'h10408000;
      9504: inst = 32'hc404796;
      9505: inst = 32'h8220000;
      9506: inst = 32'h10408000;
      9507: inst = 32'hc404797;
      9508: inst = 32'h8220000;
      9509: inst = 32'h10408000;
      9510: inst = 32'hc404798;
      9511: inst = 32'h8220000;
      9512: inst = 32'h10408000;
      9513: inst = 32'hc404799;
      9514: inst = 32'h8220000;
      9515: inst = 32'h10408000;
      9516: inst = 32'hc40479a;
      9517: inst = 32'h8220000;
      9518: inst = 32'h10408000;
      9519: inst = 32'hc40479b;
      9520: inst = 32'h8220000;
      9521: inst = 32'h10408000;
      9522: inst = 32'hc40479c;
      9523: inst = 32'h8220000;
      9524: inst = 32'h10408000;
      9525: inst = 32'hc40479d;
      9526: inst = 32'h8220000;
      9527: inst = 32'h10408000;
      9528: inst = 32'hc40479e;
      9529: inst = 32'h8220000;
      9530: inst = 32'h10408000;
      9531: inst = 32'hc40479f;
      9532: inst = 32'h8220000;
      9533: inst = 32'h10408000;
      9534: inst = 32'hc4047a0;
      9535: inst = 32'h8220000;
      9536: inst = 32'h10408000;
      9537: inst = 32'hc4047a1;
      9538: inst = 32'h8220000;
      9539: inst = 32'h10408000;
      9540: inst = 32'hc4047a2;
      9541: inst = 32'h8220000;
      9542: inst = 32'h10408000;
      9543: inst = 32'hc4047a3;
      9544: inst = 32'h8220000;
      9545: inst = 32'h10408000;
      9546: inst = 32'hc4047dc;
      9547: inst = 32'h8220000;
      9548: inst = 32'h10408000;
      9549: inst = 32'hc4047dd;
      9550: inst = 32'h8220000;
      9551: inst = 32'h10408000;
      9552: inst = 32'hc4047de;
      9553: inst = 32'h8220000;
      9554: inst = 32'h10408000;
      9555: inst = 32'hc4047df;
      9556: inst = 32'h8220000;
      9557: inst = 32'h10408000;
      9558: inst = 32'hc4047e0;
      9559: inst = 32'h8220000;
      9560: inst = 32'h10408000;
      9561: inst = 32'hc4047e1;
      9562: inst = 32'h8220000;
      9563: inst = 32'h10408000;
      9564: inst = 32'hc4047e2;
      9565: inst = 32'h8220000;
      9566: inst = 32'h10408000;
      9567: inst = 32'hc4047e3;
      9568: inst = 32'h8220000;
      9569: inst = 32'h10408000;
      9570: inst = 32'hc4047e4;
      9571: inst = 32'h8220000;
      9572: inst = 32'h10408000;
      9573: inst = 32'hc4047e5;
      9574: inst = 32'h8220000;
      9575: inst = 32'h10408000;
      9576: inst = 32'hc4047e6;
      9577: inst = 32'h8220000;
      9578: inst = 32'h10408000;
      9579: inst = 32'hc4047e7;
      9580: inst = 32'h8220000;
      9581: inst = 32'h10408000;
      9582: inst = 32'hc4047e8;
      9583: inst = 32'h8220000;
      9584: inst = 32'h10408000;
      9585: inst = 32'hc4047e9;
      9586: inst = 32'h8220000;
      9587: inst = 32'h10408000;
      9588: inst = 32'hc4047ea;
      9589: inst = 32'h8220000;
      9590: inst = 32'h10408000;
      9591: inst = 32'hc4047eb;
      9592: inst = 32'h8220000;
      9593: inst = 32'h10408000;
      9594: inst = 32'hc4047ec;
      9595: inst = 32'h8220000;
      9596: inst = 32'h10408000;
      9597: inst = 32'hc4047ed;
      9598: inst = 32'h8220000;
      9599: inst = 32'h10408000;
      9600: inst = 32'hc4047ee;
      9601: inst = 32'h8220000;
      9602: inst = 32'h10408000;
      9603: inst = 32'hc4047ef;
      9604: inst = 32'h8220000;
      9605: inst = 32'h10408000;
      9606: inst = 32'hc4047f0;
      9607: inst = 32'h8220000;
      9608: inst = 32'h10408000;
      9609: inst = 32'hc4047f1;
      9610: inst = 32'h8220000;
      9611: inst = 32'h10408000;
      9612: inst = 32'hc4047f2;
      9613: inst = 32'h8220000;
      9614: inst = 32'h10408000;
      9615: inst = 32'hc4047f3;
      9616: inst = 32'h8220000;
      9617: inst = 32'h10408000;
      9618: inst = 32'hc4047f4;
      9619: inst = 32'h8220000;
      9620: inst = 32'h10408000;
      9621: inst = 32'hc4047f5;
      9622: inst = 32'h8220000;
      9623: inst = 32'h10408000;
      9624: inst = 32'hc4047f6;
      9625: inst = 32'h8220000;
      9626: inst = 32'h10408000;
      9627: inst = 32'hc4047f7;
      9628: inst = 32'h8220000;
      9629: inst = 32'h10408000;
      9630: inst = 32'hc4047f8;
      9631: inst = 32'h8220000;
      9632: inst = 32'h10408000;
      9633: inst = 32'hc4047f9;
      9634: inst = 32'h8220000;
      9635: inst = 32'h10408000;
      9636: inst = 32'hc4047fa;
      9637: inst = 32'h8220000;
      9638: inst = 32'h10408000;
      9639: inst = 32'hc4047fb;
      9640: inst = 32'h8220000;
      9641: inst = 32'h10408000;
      9642: inst = 32'hc4047fc;
      9643: inst = 32'h8220000;
      9644: inst = 32'h10408000;
      9645: inst = 32'hc4047fd;
      9646: inst = 32'h8220000;
      9647: inst = 32'h10408000;
      9648: inst = 32'hc4047fe;
      9649: inst = 32'h8220000;
      9650: inst = 32'h10408000;
      9651: inst = 32'hc4047ff;
      9652: inst = 32'h8220000;
      9653: inst = 32'h10408000;
      9654: inst = 32'hc404800;
      9655: inst = 32'h8220000;
      9656: inst = 32'h10408000;
      9657: inst = 32'hc404801;
      9658: inst = 32'h8220000;
      9659: inst = 32'h10408000;
      9660: inst = 32'hc404802;
      9661: inst = 32'h8220000;
      9662: inst = 32'h10408000;
      9663: inst = 32'hc404803;
      9664: inst = 32'h8220000;
      9665: inst = 32'h10408000;
      9666: inst = 32'hc40483c;
      9667: inst = 32'h8220000;
      9668: inst = 32'h10408000;
      9669: inst = 32'hc40483d;
      9670: inst = 32'h8220000;
      9671: inst = 32'h10408000;
      9672: inst = 32'hc40483e;
      9673: inst = 32'h8220000;
      9674: inst = 32'h10408000;
      9675: inst = 32'hc40483f;
      9676: inst = 32'h8220000;
      9677: inst = 32'h10408000;
      9678: inst = 32'hc404840;
      9679: inst = 32'h8220000;
      9680: inst = 32'h10408000;
      9681: inst = 32'hc404841;
      9682: inst = 32'h8220000;
      9683: inst = 32'h10408000;
      9684: inst = 32'hc404842;
      9685: inst = 32'h8220000;
      9686: inst = 32'h10408000;
      9687: inst = 32'hc404843;
      9688: inst = 32'h8220000;
      9689: inst = 32'h10408000;
      9690: inst = 32'hc404844;
      9691: inst = 32'h8220000;
      9692: inst = 32'h10408000;
      9693: inst = 32'hc404845;
      9694: inst = 32'h8220000;
      9695: inst = 32'h10408000;
      9696: inst = 32'hc404846;
      9697: inst = 32'h8220000;
      9698: inst = 32'h10408000;
      9699: inst = 32'hc404847;
      9700: inst = 32'h8220000;
      9701: inst = 32'h10408000;
      9702: inst = 32'hc404848;
      9703: inst = 32'h8220000;
      9704: inst = 32'h10408000;
      9705: inst = 32'hc404849;
      9706: inst = 32'h8220000;
      9707: inst = 32'h10408000;
      9708: inst = 32'hc40484a;
      9709: inst = 32'h8220000;
      9710: inst = 32'h10408000;
      9711: inst = 32'hc40484b;
      9712: inst = 32'h8220000;
      9713: inst = 32'h10408000;
      9714: inst = 32'hc40484c;
      9715: inst = 32'h8220000;
      9716: inst = 32'h10408000;
      9717: inst = 32'hc40484d;
      9718: inst = 32'h8220000;
      9719: inst = 32'h10408000;
      9720: inst = 32'hc40484e;
      9721: inst = 32'h8220000;
      9722: inst = 32'h10408000;
      9723: inst = 32'hc40484f;
      9724: inst = 32'h8220000;
      9725: inst = 32'h10408000;
      9726: inst = 32'hc404850;
      9727: inst = 32'h8220000;
      9728: inst = 32'h10408000;
      9729: inst = 32'hc404851;
      9730: inst = 32'h8220000;
      9731: inst = 32'h10408000;
      9732: inst = 32'hc404852;
      9733: inst = 32'h8220000;
      9734: inst = 32'h10408000;
      9735: inst = 32'hc404853;
      9736: inst = 32'h8220000;
      9737: inst = 32'h10408000;
      9738: inst = 32'hc404854;
      9739: inst = 32'h8220000;
      9740: inst = 32'h10408000;
      9741: inst = 32'hc404855;
      9742: inst = 32'h8220000;
      9743: inst = 32'h10408000;
      9744: inst = 32'hc404856;
      9745: inst = 32'h8220000;
      9746: inst = 32'h10408000;
      9747: inst = 32'hc404857;
      9748: inst = 32'h8220000;
      9749: inst = 32'h10408000;
      9750: inst = 32'hc404858;
      9751: inst = 32'h8220000;
      9752: inst = 32'h10408000;
      9753: inst = 32'hc404859;
      9754: inst = 32'h8220000;
      9755: inst = 32'h10408000;
      9756: inst = 32'hc40485a;
      9757: inst = 32'h8220000;
      9758: inst = 32'h10408000;
      9759: inst = 32'hc40485b;
      9760: inst = 32'h8220000;
      9761: inst = 32'h10408000;
      9762: inst = 32'hc40485c;
      9763: inst = 32'h8220000;
      9764: inst = 32'h10408000;
      9765: inst = 32'hc40485d;
      9766: inst = 32'h8220000;
      9767: inst = 32'h10408000;
      9768: inst = 32'hc40485e;
      9769: inst = 32'h8220000;
      9770: inst = 32'h10408000;
      9771: inst = 32'hc40485f;
      9772: inst = 32'h8220000;
      9773: inst = 32'h10408000;
      9774: inst = 32'hc404860;
      9775: inst = 32'h8220000;
      9776: inst = 32'h10408000;
      9777: inst = 32'hc404861;
      9778: inst = 32'h8220000;
      9779: inst = 32'h10408000;
      9780: inst = 32'hc404862;
      9781: inst = 32'h8220000;
      9782: inst = 32'h10408000;
      9783: inst = 32'hc404863;
      9784: inst = 32'h8220000;
      9785: inst = 32'h10408000;
      9786: inst = 32'hc40489c;
      9787: inst = 32'h8220000;
      9788: inst = 32'h10408000;
      9789: inst = 32'hc40489d;
      9790: inst = 32'h8220000;
      9791: inst = 32'h10408000;
      9792: inst = 32'hc40489e;
      9793: inst = 32'h8220000;
      9794: inst = 32'h10408000;
      9795: inst = 32'hc40489f;
      9796: inst = 32'h8220000;
      9797: inst = 32'h10408000;
      9798: inst = 32'hc4048a0;
      9799: inst = 32'h8220000;
      9800: inst = 32'h10408000;
      9801: inst = 32'hc4048a1;
      9802: inst = 32'h8220000;
      9803: inst = 32'h10408000;
      9804: inst = 32'hc4048a2;
      9805: inst = 32'h8220000;
      9806: inst = 32'h10408000;
      9807: inst = 32'hc4048a3;
      9808: inst = 32'h8220000;
      9809: inst = 32'h10408000;
      9810: inst = 32'hc4048a4;
      9811: inst = 32'h8220000;
      9812: inst = 32'h10408000;
      9813: inst = 32'hc4048a5;
      9814: inst = 32'h8220000;
      9815: inst = 32'h10408000;
      9816: inst = 32'hc4048a6;
      9817: inst = 32'h8220000;
      9818: inst = 32'h10408000;
      9819: inst = 32'hc4048a7;
      9820: inst = 32'h8220000;
      9821: inst = 32'h10408000;
      9822: inst = 32'hc4048a8;
      9823: inst = 32'h8220000;
      9824: inst = 32'h10408000;
      9825: inst = 32'hc4048a9;
      9826: inst = 32'h8220000;
      9827: inst = 32'h10408000;
      9828: inst = 32'hc4048aa;
      9829: inst = 32'h8220000;
      9830: inst = 32'h10408000;
      9831: inst = 32'hc4048ab;
      9832: inst = 32'h8220000;
      9833: inst = 32'h10408000;
      9834: inst = 32'hc4048ac;
      9835: inst = 32'h8220000;
      9836: inst = 32'h10408000;
      9837: inst = 32'hc4048ad;
      9838: inst = 32'h8220000;
      9839: inst = 32'h10408000;
      9840: inst = 32'hc4048ae;
      9841: inst = 32'h8220000;
      9842: inst = 32'h10408000;
      9843: inst = 32'hc4048af;
      9844: inst = 32'h8220000;
      9845: inst = 32'h10408000;
      9846: inst = 32'hc4048b0;
      9847: inst = 32'h8220000;
      9848: inst = 32'h10408000;
      9849: inst = 32'hc4048b1;
      9850: inst = 32'h8220000;
      9851: inst = 32'h10408000;
      9852: inst = 32'hc4048b2;
      9853: inst = 32'h8220000;
      9854: inst = 32'h10408000;
      9855: inst = 32'hc4048b3;
      9856: inst = 32'h8220000;
      9857: inst = 32'h10408000;
      9858: inst = 32'hc4048b4;
      9859: inst = 32'h8220000;
      9860: inst = 32'h10408000;
      9861: inst = 32'hc4048b5;
      9862: inst = 32'h8220000;
      9863: inst = 32'h10408000;
      9864: inst = 32'hc4048b6;
      9865: inst = 32'h8220000;
      9866: inst = 32'h10408000;
      9867: inst = 32'hc4048b7;
      9868: inst = 32'h8220000;
      9869: inst = 32'h10408000;
      9870: inst = 32'hc4048b8;
      9871: inst = 32'h8220000;
      9872: inst = 32'h10408000;
      9873: inst = 32'hc4048b9;
      9874: inst = 32'h8220000;
      9875: inst = 32'h10408000;
      9876: inst = 32'hc4048ba;
      9877: inst = 32'h8220000;
      9878: inst = 32'h10408000;
      9879: inst = 32'hc4048bb;
      9880: inst = 32'h8220000;
      9881: inst = 32'h10408000;
      9882: inst = 32'hc4048bc;
      9883: inst = 32'h8220000;
      9884: inst = 32'h10408000;
      9885: inst = 32'hc4048bd;
      9886: inst = 32'h8220000;
      9887: inst = 32'h10408000;
      9888: inst = 32'hc4048be;
      9889: inst = 32'h8220000;
      9890: inst = 32'h10408000;
      9891: inst = 32'hc4048bf;
      9892: inst = 32'h8220000;
      9893: inst = 32'h10408000;
      9894: inst = 32'hc4048c0;
      9895: inst = 32'h8220000;
      9896: inst = 32'h10408000;
      9897: inst = 32'hc4048c1;
      9898: inst = 32'h8220000;
      9899: inst = 32'h10408000;
      9900: inst = 32'hc4048c2;
      9901: inst = 32'h8220000;
      9902: inst = 32'h10408000;
      9903: inst = 32'hc4048c3;
      9904: inst = 32'h8220000;
      9905: inst = 32'h10408000;
      9906: inst = 32'hc4048fc;
      9907: inst = 32'h8220000;
      9908: inst = 32'h10408000;
      9909: inst = 32'hc4048fd;
      9910: inst = 32'h8220000;
      9911: inst = 32'h10408000;
      9912: inst = 32'hc4048fe;
      9913: inst = 32'h8220000;
      9914: inst = 32'h10408000;
      9915: inst = 32'hc4048ff;
      9916: inst = 32'h8220000;
      9917: inst = 32'h10408000;
      9918: inst = 32'hc404900;
      9919: inst = 32'h8220000;
      9920: inst = 32'h10408000;
      9921: inst = 32'hc404901;
      9922: inst = 32'h8220000;
      9923: inst = 32'h10408000;
      9924: inst = 32'hc404902;
      9925: inst = 32'h8220000;
      9926: inst = 32'h10408000;
      9927: inst = 32'hc404903;
      9928: inst = 32'h8220000;
      9929: inst = 32'h10408000;
      9930: inst = 32'hc404904;
      9931: inst = 32'h8220000;
      9932: inst = 32'h10408000;
      9933: inst = 32'hc404905;
      9934: inst = 32'h8220000;
      9935: inst = 32'h10408000;
      9936: inst = 32'hc404906;
      9937: inst = 32'h8220000;
      9938: inst = 32'h10408000;
      9939: inst = 32'hc404907;
      9940: inst = 32'h8220000;
      9941: inst = 32'h10408000;
      9942: inst = 32'hc404908;
      9943: inst = 32'h8220000;
      9944: inst = 32'h10408000;
      9945: inst = 32'hc404909;
      9946: inst = 32'h8220000;
      9947: inst = 32'h10408000;
      9948: inst = 32'hc40490a;
      9949: inst = 32'h8220000;
      9950: inst = 32'h10408000;
      9951: inst = 32'hc40490b;
      9952: inst = 32'h8220000;
      9953: inst = 32'h10408000;
      9954: inst = 32'hc40490c;
      9955: inst = 32'h8220000;
      9956: inst = 32'h10408000;
      9957: inst = 32'hc40490d;
      9958: inst = 32'h8220000;
      9959: inst = 32'h10408000;
      9960: inst = 32'hc40490e;
      9961: inst = 32'h8220000;
      9962: inst = 32'h10408000;
      9963: inst = 32'hc40490f;
      9964: inst = 32'h8220000;
      9965: inst = 32'h10408000;
      9966: inst = 32'hc404910;
      9967: inst = 32'h8220000;
      9968: inst = 32'h10408000;
      9969: inst = 32'hc404911;
      9970: inst = 32'h8220000;
      9971: inst = 32'h10408000;
      9972: inst = 32'hc404912;
      9973: inst = 32'h8220000;
      9974: inst = 32'h10408000;
      9975: inst = 32'hc404913;
      9976: inst = 32'h8220000;
      9977: inst = 32'h10408000;
      9978: inst = 32'hc404914;
      9979: inst = 32'h8220000;
      9980: inst = 32'h10408000;
      9981: inst = 32'hc404915;
      9982: inst = 32'h8220000;
      9983: inst = 32'h10408000;
      9984: inst = 32'hc404916;
      9985: inst = 32'h8220000;
      9986: inst = 32'h10408000;
      9987: inst = 32'hc404917;
      9988: inst = 32'h8220000;
      9989: inst = 32'h10408000;
      9990: inst = 32'hc404918;
      9991: inst = 32'h8220000;
      9992: inst = 32'h10408000;
      9993: inst = 32'hc404919;
      9994: inst = 32'h8220000;
      9995: inst = 32'h10408000;
      9996: inst = 32'hc40491a;
      9997: inst = 32'h8220000;
      9998: inst = 32'h10408000;
      9999: inst = 32'hc40491b;
      10000: inst = 32'h8220000;
      10001: inst = 32'h10408000;
      10002: inst = 32'hc40491c;
      10003: inst = 32'h8220000;
      10004: inst = 32'h10408000;
      10005: inst = 32'hc40491d;
      10006: inst = 32'h8220000;
      10007: inst = 32'h10408000;
      10008: inst = 32'hc40491e;
      10009: inst = 32'h8220000;
      10010: inst = 32'h10408000;
      10011: inst = 32'hc40491f;
      10012: inst = 32'h8220000;
      10013: inst = 32'h10408000;
      10014: inst = 32'hc404920;
      10015: inst = 32'h8220000;
      10016: inst = 32'h10408000;
      10017: inst = 32'hc404921;
      10018: inst = 32'h8220000;
      10019: inst = 32'h10408000;
      10020: inst = 32'hc404922;
      10021: inst = 32'h8220000;
      10022: inst = 32'h10408000;
      10023: inst = 32'hc404923;
      10024: inst = 32'h8220000;
      10025: inst = 32'h10408000;
      10026: inst = 32'hc40495c;
      10027: inst = 32'h8220000;
      10028: inst = 32'h10408000;
      10029: inst = 32'hc40495d;
      10030: inst = 32'h8220000;
      10031: inst = 32'h10408000;
      10032: inst = 32'hc40495e;
      10033: inst = 32'h8220000;
      10034: inst = 32'h10408000;
      10035: inst = 32'hc40495f;
      10036: inst = 32'h8220000;
      10037: inst = 32'h10408000;
      10038: inst = 32'hc404960;
      10039: inst = 32'h8220000;
      10040: inst = 32'h10408000;
      10041: inst = 32'hc404961;
      10042: inst = 32'h8220000;
      10043: inst = 32'h10408000;
      10044: inst = 32'hc404962;
      10045: inst = 32'h8220000;
      10046: inst = 32'h10408000;
      10047: inst = 32'hc404963;
      10048: inst = 32'h8220000;
      10049: inst = 32'h10408000;
      10050: inst = 32'hc404964;
      10051: inst = 32'h8220000;
      10052: inst = 32'h10408000;
      10053: inst = 32'hc404965;
      10054: inst = 32'h8220000;
      10055: inst = 32'h10408000;
      10056: inst = 32'hc404966;
      10057: inst = 32'h8220000;
      10058: inst = 32'h10408000;
      10059: inst = 32'hc404967;
      10060: inst = 32'h8220000;
      10061: inst = 32'h10408000;
      10062: inst = 32'hc404968;
      10063: inst = 32'h8220000;
      10064: inst = 32'h10408000;
      10065: inst = 32'hc404969;
      10066: inst = 32'h8220000;
      10067: inst = 32'h10408000;
      10068: inst = 32'hc40496a;
      10069: inst = 32'h8220000;
      10070: inst = 32'h10408000;
      10071: inst = 32'hc40496b;
      10072: inst = 32'h8220000;
      10073: inst = 32'h10408000;
      10074: inst = 32'hc40496c;
      10075: inst = 32'h8220000;
      10076: inst = 32'h10408000;
      10077: inst = 32'hc40496d;
      10078: inst = 32'h8220000;
      10079: inst = 32'h10408000;
      10080: inst = 32'hc40496e;
      10081: inst = 32'h8220000;
      10082: inst = 32'h10408000;
      10083: inst = 32'hc40496f;
      10084: inst = 32'h8220000;
      10085: inst = 32'h10408000;
      10086: inst = 32'hc404970;
      10087: inst = 32'h8220000;
      10088: inst = 32'h10408000;
      10089: inst = 32'hc404971;
      10090: inst = 32'h8220000;
      10091: inst = 32'h10408000;
      10092: inst = 32'hc404972;
      10093: inst = 32'h8220000;
      10094: inst = 32'h10408000;
      10095: inst = 32'hc404973;
      10096: inst = 32'h8220000;
      10097: inst = 32'h10408000;
      10098: inst = 32'hc404974;
      10099: inst = 32'h8220000;
      10100: inst = 32'h10408000;
      10101: inst = 32'hc404975;
      10102: inst = 32'h8220000;
      10103: inst = 32'h10408000;
      10104: inst = 32'hc404976;
      10105: inst = 32'h8220000;
      10106: inst = 32'h10408000;
      10107: inst = 32'hc404977;
      10108: inst = 32'h8220000;
      10109: inst = 32'h10408000;
      10110: inst = 32'hc404978;
      10111: inst = 32'h8220000;
      10112: inst = 32'h10408000;
      10113: inst = 32'hc404979;
      10114: inst = 32'h8220000;
      10115: inst = 32'h10408000;
      10116: inst = 32'hc40497a;
      10117: inst = 32'h8220000;
      10118: inst = 32'h10408000;
      10119: inst = 32'hc40497b;
      10120: inst = 32'h8220000;
      10121: inst = 32'h10408000;
      10122: inst = 32'hc40497c;
      10123: inst = 32'h8220000;
      10124: inst = 32'h10408000;
      10125: inst = 32'hc40497d;
      10126: inst = 32'h8220000;
      10127: inst = 32'h10408000;
      10128: inst = 32'hc40497e;
      10129: inst = 32'h8220000;
      10130: inst = 32'h10408000;
      10131: inst = 32'hc40497f;
      10132: inst = 32'h8220000;
      10133: inst = 32'h10408000;
      10134: inst = 32'hc404980;
      10135: inst = 32'h8220000;
      10136: inst = 32'h10408000;
      10137: inst = 32'hc404981;
      10138: inst = 32'h8220000;
      10139: inst = 32'h10408000;
      10140: inst = 32'hc404982;
      10141: inst = 32'h8220000;
      10142: inst = 32'h10408000;
      10143: inst = 32'hc404983;
      10144: inst = 32'h8220000;
      10145: inst = 32'h10408000;
      10146: inst = 32'hc404992;
      10147: inst = 32'h8220000;
      10148: inst = 32'h10408000;
      10149: inst = 32'hc4049bc;
      10150: inst = 32'h8220000;
      10151: inst = 32'h10408000;
      10152: inst = 32'hc4049bd;
      10153: inst = 32'h8220000;
      10154: inst = 32'h10408000;
      10155: inst = 32'hc4049be;
      10156: inst = 32'h8220000;
      10157: inst = 32'h10408000;
      10158: inst = 32'hc4049bf;
      10159: inst = 32'h8220000;
      10160: inst = 32'h10408000;
      10161: inst = 32'hc4049c0;
      10162: inst = 32'h8220000;
      10163: inst = 32'h10408000;
      10164: inst = 32'hc4049c1;
      10165: inst = 32'h8220000;
      10166: inst = 32'h10408000;
      10167: inst = 32'hc4049c2;
      10168: inst = 32'h8220000;
      10169: inst = 32'h10408000;
      10170: inst = 32'hc4049c3;
      10171: inst = 32'h8220000;
      10172: inst = 32'h10408000;
      10173: inst = 32'hc4049c4;
      10174: inst = 32'h8220000;
      10175: inst = 32'h10408000;
      10176: inst = 32'hc4049c5;
      10177: inst = 32'h8220000;
      10178: inst = 32'h10408000;
      10179: inst = 32'hc4049c6;
      10180: inst = 32'h8220000;
      10181: inst = 32'h10408000;
      10182: inst = 32'hc4049c7;
      10183: inst = 32'h8220000;
      10184: inst = 32'h10408000;
      10185: inst = 32'hc4049c8;
      10186: inst = 32'h8220000;
      10187: inst = 32'h10408000;
      10188: inst = 32'hc4049c9;
      10189: inst = 32'h8220000;
      10190: inst = 32'h10408000;
      10191: inst = 32'hc4049ca;
      10192: inst = 32'h8220000;
      10193: inst = 32'h10408000;
      10194: inst = 32'hc4049cb;
      10195: inst = 32'h8220000;
      10196: inst = 32'h10408000;
      10197: inst = 32'hc4049cc;
      10198: inst = 32'h8220000;
      10199: inst = 32'h10408000;
      10200: inst = 32'hc4049cd;
      10201: inst = 32'h8220000;
      10202: inst = 32'h10408000;
      10203: inst = 32'hc4049ce;
      10204: inst = 32'h8220000;
      10205: inst = 32'h10408000;
      10206: inst = 32'hc4049cf;
      10207: inst = 32'h8220000;
      10208: inst = 32'h10408000;
      10209: inst = 32'hc4049d0;
      10210: inst = 32'h8220000;
      10211: inst = 32'h10408000;
      10212: inst = 32'hc4049d1;
      10213: inst = 32'h8220000;
      10214: inst = 32'h10408000;
      10215: inst = 32'hc4049d2;
      10216: inst = 32'h8220000;
      10217: inst = 32'h10408000;
      10218: inst = 32'hc4049d3;
      10219: inst = 32'h8220000;
      10220: inst = 32'h10408000;
      10221: inst = 32'hc4049d4;
      10222: inst = 32'h8220000;
      10223: inst = 32'h10408000;
      10224: inst = 32'hc4049d5;
      10225: inst = 32'h8220000;
      10226: inst = 32'h10408000;
      10227: inst = 32'hc4049d6;
      10228: inst = 32'h8220000;
      10229: inst = 32'h10408000;
      10230: inst = 32'hc4049d7;
      10231: inst = 32'h8220000;
      10232: inst = 32'h10408000;
      10233: inst = 32'hc4049d8;
      10234: inst = 32'h8220000;
      10235: inst = 32'h10408000;
      10236: inst = 32'hc4049d9;
      10237: inst = 32'h8220000;
      10238: inst = 32'h10408000;
      10239: inst = 32'hc4049da;
      10240: inst = 32'h8220000;
      10241: inst = 32'h10408000;
      10242: inst = 32'hc4049db;
      10243: inst = 32'h8220000;
      10244: inst = 32'h10408000;
      10245: inst = 32'hc4049dc;
      10246: inst = 32'h8220000;
      10247: inst = 32'h10408000;
      10248: inst = 32'hc4049dd;
      10249: inst = 32'h8220000;
      10250: inst = 32'h10408000;
      10251: inst = 32'hc4049de;
      10252: inst = 32'h8220000;
      10253: inst = 32'h10408000;
      10254: inst = 32'hc4049df;
      10255: inst = 32'h8220000;
      10256: inst = 32'h10408000;
      10257: inst = 32'hc4049e0;
      10258: inst = 32'h8220000;
      10259: inst = 32'h10408000;
      10260: inst = 32'hc4049e1;
      10261: inst = 32'h8220000;
      10262: inst = 32'h10408000;
      10263: inst = 32'hc4049e2;
      10264: inst = 32'h8220000;
      10265: inst = 32'h10408000;
      10266: inst = 32'hc4049e3;
      10267: inst = 32'h8220000;
      10268: inst = 32'h10408000;
      10269: inst = 32'hc4049f2;
      10270: inst = 32'h8220000;
      10271: inst = 32'h10408000;
      10272: inst = 32'hc404a1c;
      10273: inst = 32'h8220000;
      10274: inst = 32'h10408000;
      10275: inst = 32'hc404a1d;
      10276: inst = 32'h8220000;
      10277: inst = 32'h10408000;
      10278: inst = 32'hc404a1e;
      10279: inst = 32'h8220000;
      10280: inst = 32'h10408000;
      10281: inst = 32'hc404a1f;
      10282: inst = 32'h8220000;
      10283: inst = 32'h10408000;
      10284: inst = 32'hc404a20;
      10285: inst = 32'h8220000;
      10286: inst = 32'h10408000;
      10287: inst = 32'hc404a21;
      10288: inst = 32'h8220000;
      10289: inst = 32'h10408000;
      10290: inst = 32'hc404a22;
      10291: inst = 32'h8220000;
      10292: inst = 32'h10408000;
      10293: inst = 32'hc404a23;
      10294: inst = 32'h8220000;
      10295: inst = 32'h10408000;
      10296: inst = 32'hc404a24;
      10297: inst = 32'h8220000;
      10298: inst = 32'h10408000;
      10299: inst = 32'hc404a25;
      10300: inst = 32'h8220000;
      10301: inst = 32'h10408000;
      10302: inst = 32'hc404a26;
      10303: inst = 32'h8220000;
      10304: inst = 32'h10408000;
      10305: inst = 32'hc404a27;
      10306: inst = 32'h8220000;
      10307: inst = 32'h10408000;
      10308: inst = 32'hc404a28;
      10309: inst = 32'h8220000;
      10310: inst = 32'h10408000;
      10311: inst = 32'hc404a29;
      10312: inst = 32'h8220000;
      10313: inst = 32'h10408000;
      10314: inst = 32'hc404a2a;
      10315: inst = 32'h8220000;
      10316: inst = 32'h10408000;
      10317: inst = 32'hc404a2b;
      10318: inst = 32'h8220000;
      10319: inst = 32'h10408000;
      10320: inst = 32'hc404a2c;
      10321: inst = 32'h8220000;
      10322: inst = 32'h10408000;
      10323: inst = 32'hc404a2d;
      10324: inst = 32'h8220000;
      10325: inst = 32'h10408000;
      10326: inst = 32'hc404a2e;
      10327: inst = 32'h8220000;
      10328: inst = 32'h10408000;
      10329: inst = 32'hc404a2f;
      10330: inst = 32'h8220000;
      10331: inst = 32'h10408000;
      10332: inst = 32'hc404a30;
      10333: inst = 32'h8220000;
      10334: inst = 32'h10408000;
      10335: inst = 32'hc404a31;
      10336: inst = 32'h8220000;
      10337: inst = 32'h10408000;
      10338: inst = 32'hc404a32;
      10339: inst = 32'h8220000;
      10340: inst = 32'h10408000;
      10341: inst = 32'hc404a33;
      10342: inst = 32'h8220000;
      10343: inst = 32'h10408000;
      10344: inst = 32'hc404a34;
      10345: inst = 32'h8220000;
      10346: inst = 32'h10408000;
      10347: inst = 32'hc404a35;
      10348: inst = 32'h8220000;
      10349: inst = 32'h10408000;
      10350: inst = 32'hc404a36;
      10351: inst = 32'h8220000;
      10352: inst = 32'h10408000;
      10353: inst = 32'hc404a37;
      10354: inst = 32'h8220000;
      10355: inst = 32'h10408000;
      10356: inst = 32'hc404a38;
      10357: inst = 32'h8220000;
      10358: inst = 32'h10408000;
      10359: inst = 32'hc404a39;
      10360: inst = 32'h8220000;
      10361: inst = 32'h10408000;
      10362: inst = 32'hc404a3a;
      10363: inst = 32'h8220000;
      10364: inst = 32'h10408000;
      10365: inst = 32'hc404a3b;
      10366: inst = 32'h8220000;
      10367: inst = 32'h10408000;
      10368: inst = 32'hc404a3c;
      10369: inst = 32'h8220000;
      10370: inst = 32'h10408000;
      10371: inst = 32'hc404a3d;
      10372: inst = 32'h8220000;
      10373: inst = 32'h10408000;
      10374: inst = 32'hc404a3e;
      10375: inst = 32'h8220000;
      10376: inst = 32'h10408000;
      10377: inst = 32'hc404a3f;
      10378: inst = 32'h8220000;
      10379: inst = 32'h10408000;
      10380: inst = 32'hc404a40;
      10381: inst = 32'h8220000;
      10382: inst = 32'h10408000;
      10383: inst = 32'hc404a41;
      10384: inst = 32'h8220000;
      10385: inst = 32'h10408000;
      10386: inst = 32'hc404a42;
      10387: inst = 32'h8220000;
      10388: inst = 32'h10408000;
      10389: inst = 32'hc404a43;
      10390: inst = 32'h8220000;
      10391: inst = 32'h10408000;
      10392: inst = 32'hc404a52;
      10393: inst = 32'h8220000;
      10394: inst = 32'h10408000;
      10395: inst = 32'hc404a7c;
      10396: inst = 32'h8220000;
      10397: inst = 32'h10408000;
      10398: inst = 32'hc404a7d;
      10399: inst = 32'h8220000;
      10400: inst = 32'h10408000;
      10401: inst = 32'hc404a7e;
      10402: inst = 32'h8220000;
      10403: inst = 32'h10408000;
      10404: inst = 32'hc404a7f;
      10405: inst = 32'h8220000;
      10406: inst = 32'h10408000;
      10407: inst = 32'hc404a80;
      10408: inst = 32'h8220000;
      10409: inst = 32'h10408000;
      10410: inst = 32'hc404a81;
      10411: inst = 32'h8220000;
      10412: inst = 32'h10408000;
      10413: inst = 32'hc404a82;
      10414: inst = 32'h8220000;
      10415: inst = 32'h10408000;
      10416: inst = 32'hc404a83;
      10417: inst = 32'h8220000;
      10418: inst = 32'h10408000;
      10419: inst = 32'hc404a84;
      10420: inst = 32'h8220000;
      10421: inst = 32'h10408000;
      10422: inst = 32'hc404a85;
      10423: inst = 32'h8220000;
      10424: inst = 32'h10408000;
      10425: inst = 32'hc404a86;
      10426: inst = 32'h8220000;
      10427: inst = 32'h10408000;
      10428: inst = 32'hc404a87;
      10429: inst = 32'h8220000;
      10430: inst = 32'h10408000;
      10431: inst = 32'hc404a88;
      10432: inst = 32'h8220000;
      10433: inst = 32'h10408000;
      10434: inst = 32'hc404a89;
      10435: inst = 32'h8220000;
      10436: inst = 32'h10408000;
      10437: inst = 32'hc404a8a;
      10438: inst = 32'h8220000;
      10439: inst = 32'h10408000;
      10440: inst = 32'hc404a8b;
      10441: inst = 32'h8220000;
      10442: inst = 32'h10408000;
      10443: inst = 32'hc404a8c;
      10444: inst = 32'h8220000;
      10445: inst = 32'h10408000;
      10446: inst = 32'hc404a8d;
      10447: inst = 32'h8220000;
      10448: inst = 32'h10408000;
      10449: inst = 32'hc404a8e;
      10450: inst = 32'h8220000;
      10451: inst = 32'h10408000;
      10452: inst = 32'hc404a8f;
      10453: inst = 32'h8220000;
      10454: inst = 32'h10408000;
      10455: inst = 32'hc404a90;
      10456: inst = 32'h8220000;
      10457: inst = 32'h10408000;
      10458: inst = 32'hc404a91;
      10459: inst = 32'h8220000;
      10460: inst = 32'h10408000;
      10461: inst = 32'hc404a92;
      10462: inst = 32'h8220000;
      10463: inst = 32'h10408000;
      10464: inst = 32'hc404a93;
      10465: inst = 32'h8220000;
      10466: inst = 32'h10408000;
      10467: inst = 32'hc404a94;
      10468: inst = 32'h8220000;
      10469: inst = 32'h10408000;
      10470: inst = 32'hc404a95;
      10471: inst = 32'h8220000;
      10472: inst = 32'h10408000;
      10473: inst = 32'hc404a96;
      10474: inst = 32'h8220000;
      10475: inst = 32'h10408000;
      10476: inst = 32'hc404a97;
      10477: inst = 32'h8220000;
      10478: inst = 32'h10408000;
      10479: inst = 32'hc404a98;
      10480: inst = 32'h8220000;
      10481: inst = 32'h10408000;
      10482: inst = 32'hc404a99;
      10483: inst = 32'h8220000;
      10484: inst = 32'h10408000;
      10485: inst = 32'hc404a9a;
      10486: inst = 32'h8220000;
      10487: inst = 32'h10408000;
      10488: inst = 32'hc404a9b;
      10489: inst = 32'h8220000;
      10490: inst = 32'h10408000;
      10491: inst = 32'hc404a9c;
      10492: inst = 32'h8220000;
      10493: inst = 32'h10408000;
      10494: inst = 32'hc404a9d;
      10495: inst = 32'h8220000;
      10496: inst = 32'h10408000;
      10497: inst = 32'hc404a9e;
      10498: inst = 32'h8220000;
      10499: inst = 32'h10408000;
      10500: inst = 32'hc404a9f;
      10501: inst = 32'h8220000;
      10502: inst = 32'h10408000;
      10503: inst = 32'hc404aa0;
      10504: inst = 32'h8220000;
      10505: inst = 32'h10408000;
      10506: inst = 32'hc404aa1;
      10507: inst = 32'h8220000;
      10508: inst = 32'h10408000;
      10509: inst = 32'hc404aa2;
      10510: inst = 32'h8220000;
      10511: inst = 32'h10408000;
      10512: inst = 32'hc404aa3;
      10513: inst = 32'h8220000;
      10514: inst = 32'h10408000;
      10515: inst = 32'hc404ab4;
      10516: inst = 32'h8220000;
      10517: inst = 32'h10408000;
      10518: inst = 32'hc404adc;
      10519: inst = 32'h8220000;
      10520: inst = 32'h10408000;
      10521: inst = 32'hc404add;
      10522: inst = 32'h8220000;
      10523: inst = 32'h10408000;
      10524: inst = 32'hc404ade;
      10525: inst = 32'h8220000;
      10526: inst = 32'h10408000;
      10527: inst = 32'hc404adf;
      10528: inst = 32'h8220000;
      10529: inst = 32'h10408000;
      10530: inst = 32'hc404ae0;
      10531: inst = 32'h8220000;
      10532: inst = 32'h10408000;
      10533: inst = 32'hc404ae1;
      10534: inst = 32'h8220000;
      10535: inst = 32'h10408000;
      10536: inst = 32'hc404ae2;
      10537: inst = 32'h8220000;
      10538: inst = 32'h10408000;
      10539: inst = 32'hc404ae3;
      10540: inst = 32'h8220000;
      10541: inst = 32'h10408000;
      10542: inst = 32'hc404ae4;
      10543: inst = 32'h8220000;
      10544: inst = 32'h10408000;
      10545: inst = 32'hc404ae5;
      10546: inst = 32'h8220000;
      10547: inst = 32'h10408000;
      10548: inst = 32'hc404ae6;
      10549: inst = 32'h8220000;
      10550: inst = 32'h10408000;
      10551: inst = 32'hc404ae7;
      10552: inst = 32'h8220000;
      10553: inst = 32'h10408000;
      10554: inst = 32'hc404ae8;
      10555: inst = 32'h8220000;
      10556: inst = 32'h10408000;
      10557: inst = 32'hc404ae9;
      10558: inst = 32'h8220000;
      10559: inst = 32'h10408000;
      10560: inst = 32'hc404aea;
      10561: inst = 32'h8220000;
      10562: inst = 32'h10408000;
      10563: inst = 32'hc404aeb;
      10564: inst = 32'h8220000;
      10565: inst = 32'h10408000;
      10566: inst = 32'hc404aec;
      10567: inst = 32'h8220000;
      10568: inst = 32'h10408000;
      10569: inst = 32'hc404aed;
      10570: inst = 32'h8220000;
      10571: inst = 32'h10408000;
      10572: inst = 32'hc404aee;
      10573: inst = 32'h8220000;
      10574: inst = 32'h10408000;
      10575: inst = 32'hc404aef;
      10576: inst = 32'h8220000;
      10577: inst = 32'h10408000;
      10578: inst = 32'hc404af0;
      10579: inst = 32'h8220000;
      10580: inst = 32'h10408000;
      10581: inst = 32'hc404af1;
      10582: inst = 32'h8220000;
      10583: inst = 32'h10408000;
      10584: inst = 32'hc404af2;
      10585: inst = 32'h8220000;
      10586: inst = 32'h10408000;
      10587: inst = 32'hc404af3;
      10588: inst = 32'h8220000;
      10589: inst = 32'h10408000;
      10590: inst = 32'hc404af4;
      10591: inst = 32'h8220000;
      10592: inst = 32'h10408000;
      10593: inst = 32'hc404af5;
      10594: inst = 32'h8220000;
      10595: inst = 32'h10408000;
      10596: inst = 32'hc404af6;
      10597: inst = 32'h8220000;
      10598: inst = 32'h10408000;
      10599: inst = 32'hc404af7;
      10600: inst = 32'h8220000;
      10601: inst = 32'h10408000;
      10602: inst = 32'hc404af8;
      10603: inst = 32'h8220000;
      10604: inst = 32'h10408000;
      10605: inst = 32'hc404af9;
      10606: inst = 32'h8220000;
      10607: inst = 32'h10408000;
      10608: inst = 32'hc404afa;
      10609: inst = 32'h8220000;
      10610: inst = 32'h10408000;
      10611: inst = 32'hc404afb;
      10612: inst = 32'h8220000;
      10613: inst = 32'h10408000;
      10614: inst = 32'hc404afc;
      10615: inst = 32'h8220000;
      10616: inst = 32'h10408000;
      10617: inst = 32'hc404afd;
      10618: inst = 32'h8220000;
      10619: inst = 32'h10408000;
      10620: inst = 32'hc404afe;
      10621: inst = 32'h8220000;
      10622: inst = 32'h10408000;
      10623: inst = 32'hc404aff;
      10624: inst = 32'h8220000;
      10625: inst = 32'h10408000;
      10626: inst = 32'hc404b00;
      10627: inst = 32'h8220000;
      10628: inst = 32'h10408000;
      10629: inst = 32'hc404b01;
      10630: inst = 32'h8220000;
      10631: inst = 32'h10408000;
      10632: inst = 32'hc404b02;
      10633: inst = 32'h8220000;
      10634: inst = 32'h10408000;
      10635: inst = 32'hc404b03;
      10636: inst = 32'h8220000;
      10637: inst = 32'h10408000;
      10638: inst = 32'hc404b14;
      10639: inst = 32'h8220000;
      10640: inst = 32'h10408000;
      10641: inst = 32'hc404b3c;
      10642: inst = 32'h8220000;
      10643: inst = 32'h10408000;
      10644: inst = 32'hc404b3d;
      10645: inst = 32'h8220000;
      10646: inst = 32'h10408000;
      10647: inst = 32'hc404b3e;
      10648: inst = 32'h8220000;
      10649: inst = 32'h10408000;
      10650: inst = 32'hc404b3f;
      10651: inst = 32'h8220000;
      10652: inst = 32'h10408000;
      10653: inst = 32'hc404b40;
      10654: inst = 32'h8220000;
      10655: inst = 32'h10408000;
      10656: inst = 32'hc404b41;
      10657: inst = 32'h8220000;
      10658: inst = 32'h10408000;
      10659: inst = 32'hc404b42;
      10660: inst = 32'h8220000;
      10661: inst = 32'h10408000;
      10662: inst = 32'hc404b43;
      10663: inst = 32'h8220000;
      10664: inst = 32'h10408000;
      10665: inst = 32'hc404b44;
      10666: inst = 32'h8220000;
      10667: inst = 32'h10408000;
      10668: inst = 32'hc404b45;
      10669: inst = 32'h8220000;
      10670: inst = 32'h10408000;
      10671: inst = 32'hc404b46;
      10672: inst = 32'h8220000;
      10673: inst = 32'h10408000;
      10674: inst = 32'hc404b47;
      10675: inst = 32'h8220000;
      10676: inst = 32'h10408000;
      10677: inst = 32'hc404b48;
      10678: inst = 32'h8220000;
      10679: inst = 32'h10408000;
      10680: inst = 32'hc404b49;
      10681: inst = 32'h8220000;
      10682: inst = 32'h10408000;
      10683: inst = 32'hc404b4a;
      10684: inst = 32'h8220000;
      10685: inst = 32'h10408000;
      10686: inst = 32'hc404b4b;
      10687: inst = 32'h8220000;
      10688: inst = 32'h10408000;
      10689: inst = 32'hc404b4c;
      10690: inst = 32'h8220000;
      10691: inst = 32'h10408000;
      10692: inst = 32'hc404b4d;
      10693: inst = 32'h8220000;
      10694: inst = 32'h10408000;
      10695: inst = 32'hc404b4e;
      10696: inst = 32'h8220000;
      10697: inst = 32'h10408000;
      10698: inst = 32'hc404b4f;
      10699: inst = 32'h8220000;
      10700: inst = 32'h10408000;
      10701: inst = 32'hc404b50;
      10702: inst = 32'h8220000;
      10703: inst = 32'h10408000;
      10704: inst = 32'hc404b51;
      10705: inst = 32'h8220000;
      10706: inst = 32'h10408000;
      10707: inst = 32'hc404b52;
      10708: inst = 32'h8220000;
      10709: inst = 32'h10408000;
      10710: inst = 32'hc404b53;
      10711: inst = 32'h8220000;
      10712: inst = 32'h10408000;
      10713: inst = 32'hc404b54;
      10714: inst = 32'h8220000;
      10715: inst = 32'h10408000;
      10716: inst = 32'hc404b55;
      10717: inst = 32'h8220000;
      10718: inst = 32'h10408000;
      10719: inst = 32'hc404b56;
      10720: inst = 32'h8220000;
      10721: inst = 32'h10408000;
      10722: inst = 32'hc404b57;
      10723: inst = 32'h8220000;
      10724: inst = 32'h10408000;
      10725: inst = 32'hc404b58;
      10726: inst = 32'h8220000;
      10727: inst = 32'h10408000;
      10728: inst = 32'hc404b59;
      10729: inst = 32'h8220000;
      10730: inst = 32'h10408000;
      10731: inst = 32'hc404b5a;
      10732: inst = 32'h8220000;
      10733: inst = 32'h10408000;
      10734: inst = 32'hc404b5b;
      10735: inst = 32'h8220000;
      10736: inst = 32'h10408000;
      10737: inst = 32'hc404b5c;
      10738: inst = 32'h8220000;
      10739: inst = 32'h10408000;
      10740: inst = 32'hc404b5d;
      10741: inst = 32'h8220000;
      10742: inst = 32'h10408000;
      10743: inst = 32'hc404b5e;
      10744: inst = 32'h8220000;
      10745: inst = 32'h10408000;
      10746: inst = 32'hc404b5f;
      10747: inst = 32'h8220000;
      10748: inst = 32'h10408000;
      10749: inst = 32'hc404b60;
      10750: inst = 32'h8220000;
      10751: inst = 32'h10408000;
      10752: inst = 32'hc404b61;
      10753: inst = 32'h8220000;
      10754: inst = 32'h10408000;
      10755: inst = 32'hc404b62;
      10756: inst = 32'h8220000;
      10757: inst = 32'h10408000;
      10758: inst = 32'hc404b63;
      10759: inst = 32'h8220000;
      10760: inst = 32'h10408000;
      10761: inst = 32'hc404b9c;
      10762: inst = 32'h8220000;
      10763: inst = 32'h10408000;
      10764: inst = 32'hc404b9d;
      10765: inst = 32'h8220000;
      10766: inst = 32'h10408000;
      10767: inst = 32'hc404b9e;
      10768: inst = 32'h8220000;
      10769: inst = 32'h10408000;
      10770: inst = 32'hc404b9f;
      10771: inst = 32'h8220000;
      10772: inst = 32'h10408000;
      10773: inst = 32'hc404ba0;
      10774: inst = 32'h8220000;
      10775: inst = 32'h10408000;
      10776: inst = 32'hc404ba1;
      10777: inst = 32'h8220000;
      10778: inst = 32'h10408000;
      10779: inst = 32'hc404ba2;
      10780: inst = 32'h8220000;
      10781: inst = 32'h10408000;
      10782: inst = 32'hc404ba3;
      10783: inst = 32'h8220000;
      10784: inst = 32'h10408000;
      10785: inst = 32'hc404ba4;
      10786: inst = 32'h8220000;
      10787: inst = 32'h10408000;
      10788: inst = 32'hc404ba5;
      10789: inst = 32'h8220000;
      10790: inst = 32'h10408000;
      10791: inst = 32'hc404ba6;
      10792: inst = 32'h8220000;
      10793: inst = 32'h10408000;
      10794: inst = 32'hc404ba7;
      10795: inst = 32'h8220000;
      10796: inst = 32'h10408000;
      10797: inst = 32'hc404ba8;
      10798: inst = 32'h8220000;
      10799: inst = 32'h10408000;
      10800: inst = 32'hc404ba9;
      10801: inst = 32'h8220000;
      10802: inst = 32'h10408000;
      10803: inst = 32'hc404baa;
      10804: inst = 32'h8220000;
      10805: inst = 32'h10408000;
      10806: inst = 32'hc404bab;
      10807: inst = 32'h8220000;
      10808: inst = 32'h10408000;
      10809: inst = 32'hc404bac;
      10810: inst = 32'h8220000;
      10811: inst = 32'h10408000;
      10812: inst = 32'hc404bad;
      10813: inst = 32'h8220000;
      10814: inst = 32'h10408000;
      10815: inst = 32'hc404bae;
      10816: inst = 32'h8220000;
      10817: inst = 32'h10408000;
      10818: inst = 32'hc404baf;
      10819: inst = 32'h8220000;
      10820: inst = 32'h10408000;
      10821: inst = 32'hc404bb0;
      10822: inst = 32'h8220000;
      10823: inst = 32'h10408000;
      10824: inst = 32'hc404bb1;
      10825: inst = 32'h8220000;
      10826: inst = 32'h10408000;
      10827: inst = 32'hc404bb2;
      10828: inst = 32'h8220000;
      10829: inst = 32'h10408000;
      10830: inst = 32'hc404bb3;
      10831: inst = 32'h8220000;
      10832: inst = 32'h10408000;
      10833: inst = 32'hc404bb4;
      10834: inst = 32'h8220000;
      10835: inst = 32'h10408000;
      10836: inst = 32'hc404bb5;
      10837: inst = 32'h8220000;
      10838: inst = 32'h10408000;
      10839: inst = 32'hc404bb6;
      10840: inst = 32'h8220000;
      10841: inst = 32'h10408000;
      10842: inst = 32'hc404bb7;
      10843: inst = 32'h8220000;
      10844: inst = 32'h10408000;
      10845: inst = 32'hc404bb8;
      10846: inst = 32'h8220000;
      10847: inst = 32'h10408000;
      10848: inst = 32'hc404bb9;
      10849: inst = 32'h8220000;
      10850: inst = 32'h10408000;
      10851: inst = 32'hc404bba;
      10852: inst = 32'h8220000;
      10853: inst = 32'h10408000;
      10854: inst = 32'hc404bbb;
      10855: inst = 32'h8220000;
      10856: inst = 32'h10408000;
      10857: inst = 32'hc404bbc;
      10858: inst = 32'h8220000;
      10859: inst = 32'h10408000;
      10860: inst = 32'hc404bbd;
      10861: inst = 32'h8220000;
      10862: inst = 32'h10408000;
      10863: inst = 32'hc404bbe;
      10864: inst = 32'h8220000;
      10865: inst = 32'h10408000;
      10866: inst = 32'hc404bbf;
      10867: inst = 32'h8220000;
      10868: inst = 32'h10408000;
      10869: inst = 32'hc404bc0;
      10870: inst = 32'h8220000;
      10871: inst = 32'h10408000;
      10872: inst = 32'hc404bc1;
      10873: inst = 32'h8220000;
      10874: inst = 32'h10408000;
      10875: inst = 32'hc404bc2;
      10876: inst = 32'h8220000;
      10877: inst = 32'h10408000;
      10878: inst = 32'hc404bc3;
      10879: inst = 32'h8220000;
      10880: inst = 32'hc20ee75;
      10881: inst = 32'h10408000;
      10882: inst = 32'hc4042ea;
      10883: inst = 32'h8220000;
      10884: inst = 32'h10408000;
      10885: inst = 32'hc4043a7;
      10886: inst = 32'h8220000;
      10887: inst = 32'hc20d42c;
      10888: inst = 32'h10408000;
      10889: inst = 32'hc4042eb;
      10890: inst = 32'h8220000;
      10891: inst = 32'h10408000;
      10892: inst = 32'hc4042ec;
      10893: inst = 32'h8220000;
      10894: inst = 32'h10408000;
      10895: inst = 32'hc4043a8;
      10896: inst = 32'h8220000;
      10897: inst = 32'hc20ee55;
      10898: inst = 32'h10408000;
      10899: inst = 32'hc4042ed;
      10900: inst = 32'h8220000;
      10901: inst = 32'h10408000;
      10902: inst = 32'hc4043b0;
      10903: inst = 32'h8220000;
      10904: inst = 32'hc20e571;
      10905: inst = 32'h10408000;
      10906: inst = 32'hc404349;
      10907: inst = 32'h8220000;
      10908: inst = 32'h10408000;
      10909: inst = 32'hc40434e;
      10910: inst = 32'h8220000;
      10911: inst = 32'h10408000;
      10912: inst = 32'hc404406;
      10913: inst = 32'h8220000;
      10914: inst = 32'h10408000;
      10915: inst = 32'hc404411;
      10916: inst = 32'h8220000;
      10917: inst = 32'hc20cb28;
      10918: inst = 32'h10408000;
      10919: inst = 32'hc40434a;
      10920: inst = 32'h8220000;
      10921: inst = 32'h10408000;
      10922: inst = 32'hc40434d;
      10923: inst = 32'h8220000;
      10924: inst = 32'h10408000;
      10925: inst = 32'hc404407;
      10926: inst = 32'h8220000;
      10927: inst = 32'h10408000;
      10928: inst = 32'hc404410;
      10929: inst = 32'h8220000;
      10930: inst = 32'hc20cac7;
      10931: inst = 32'h10408000;
      10932: inst = 32'hc40434b;
      10933: inst = 32'h8220000;
      10934: inst = 32'h10408000;
      10935: inst = 32'hc40434c;
      10936: inst = 32'h8220000;
      10937: inst = 32'h10408000;
      10938: inst = 32'hc4043a9;
      10939: inst = 32'h8220000;
      10940: inst = 32'h10408000;
      10941: inst = 32'hc4043aa;
      10942: inst = 32'h8220000;
      10943: inst = 32'h10408000;
      10944: inst = 32'hc4043ab;
      10945: inst = 32'h8220000;
      10946: inst = 32'h10408000;
      10947: inst = 32'hc4043ac;
      10948: inst = 32'h8220000;
      10949: inst = 32'h10408000;
      10950: inst = 32'hc4043ad;
      10951: inst = 32'h8220000;
      10952: inst = 32'h10408000;
      10953: inst = 32'hc4043ae;
      10954: inst = 32'h8220000;
      10955: inst = 32'h10408000;
      10956: inst = 32'hc404408;
      10957: inst = 32'h8220000;
      10958: inst = 32'h10408000;
      10959: inst = 32'hc404409;
      10960: inst = 32'h8220000;
      10961: inst = 32'h10408000;
      10962: inst = 32'hc40440a;
      10963: inst = 32'h8220000;
      10964: inst = 32'h10408000;
      10965: inst = 32'hc40440b;
      10966: inst = 32'h8220000;
      10967: inst = 32'h10408000;
      10968: inst = 32'hc40440c;
      10969: inst = 32'h8220000;
      10970: inst = 32'h10408000;
      10971: inst = 32'hc40440d;
      10972: inst = 32'h8220000;
      10973: inst = 32'h10408000;
      10974: inst = 32'hc40440e;
      10975: inst = 32'h8220000;
      10976: inst = 32'h10408000;
      10977: inst = 32'hc40440f;
      10978: inst = 32'h8220000;
      10979: inst = 32'hc20d40c;
      10980: inst = 32'h10408000;
      10981: inst = 32'hc4043af;
      10982: inst = 32'h8220000;
      10983: inst = 32'hc20ee8e;
      10984: inst = 32'h10408000;
      10985: inst = 32'hc40446a;
      10986: inst = 32'h8220000;
      10987: inst = 32'h10408000;
      10988: inst = 32'hc4044b5;
      10989: inst = 32'h8220000;
      10990: inst = 32'hc20ee48;
      10991: inst = 32'h10408000;
      10992: inst = 32'hc40446b;
      10993: inst = 32'h8220000;
      10994: inst = 32'h10408000;
      10995: inst = 32'hc40446c;
      10996: inst = 32'h8220000;
      10997: inst = 32'h10408000;
      10998: inst = 32'hc4044b3;
      10999: inst = 32'h8220000;
      11000: inst = 32'h10408000;
      11001: inst = 32'hc4044b4;
      11002: inst = 32'h8220000;
      11003: inst = 32'hc20ee90;
      11004: inst = 32'h10408000;
      11005: inst = 32'hc40446d;
      11006: inst = 32'h8220000;
      11007: inst = 32'h10408000;
      11008: inst = 32'hc4044b2;
      11009: inst = 32'h8220000;
      11010: inst = 32'hc20eeb5;
      11011: inst = 32'h10408000;
      11012: inst = 32'hc4044cb;
      11013: inst = 32'h8220000;
      11014: inst = 32'h10408000;
      11015: inst = 32'hc4044cc;
      11016: inst = 32'h8220000;
      11017: inst = 32'h10408000;
      11018: inst = 32'hc404513;
      11019: inst = 32'h8220000;
      11020: inst = 32'h10408000;
      11021: inst = 32'hc404514;
      11022: inst = 32'h8220000;
      11023: inst = 32'hc20c2e2;
      11024: inst = 32'h10408000;
      11025: inst = 32'hc4046ef;
      11026: inst = 32'h8220000;
      11027: inst = 32'h10408000;
      11028: inst = 32'hc4046f0;
      11029: inst = 32'h8220000;
      11030: inst = 32'h10408000;
      11031: inst = 32'hc4046f1;
      11032: inst = 32'h8220000;
      11033: inst = 32'h10408000;
      11034: inst = 32'hc4046f2;
      11035: inst = 32'h8220000;
      11036: inst = 32'h10408000;
      11037: inst = 32'hc4046f3;
      11038: inst = 32'h8220000;
      11039: inst = 32'h10408000;
      11040: inst = 32'hc4046f4;
      11041: inst = 32'h8220000;
      11042: inst = 32'h10408000;
      11043: inst = 32'hc4046f5;
      11044: inst = 32'h8220000;
      11045: inst = 32'h10408000;
      11046: inst = 32'hc4046f6;
      11047: inst = 32'h8220000;
      11048: inst = 32'h10408000;
      11049: inst = 32'hc4046f7;
      11050: inst = 32'h8220000;
      11051: inst = 32'h10408000;
      11052: inst = 32'hc4046f8;
      11053: inst = 32'h8220000;
      11054: inst = 32'h10408000;
      11055: inst = 32'hc4046f9;
      11056: inst = 32'h8220000;
      11057: inst = 32'h10408000;
      11058: inst = 32'hc4046fa;
      11059: inst = 32'h8220000;
      11060: inst = 32'h10408000;
      11061: inst = 32'hc4046fb;
      11062: inst = 32'h8220000;
      11063: inst = 32'h10408000;
      11064: inst = 32'hc4046fc;
      11065: inst = 32'h8220000;
      11066: inst = 32'h10408000;
      11067: inst = 32'hc4046fd;
      11068: inst = 32'h8220000;
      11069: inst = 32'h10408000;
      11070: inst = 32'hc4046fe;
      11071: inst = 32'h8220000;
      11072: inst = 32'h10408000;
      11073: inst = 32'hc4046ff;
      11074: inst = 32'h8220000;
      11075: inst = 32'h10408000;
      11076: inst = 32'hc40474f;
      11077: inst = 32'h8220000;
      11078: inst = 32'h10408000;
      11079: inst = 32'hc40475f;
      11080: inst = 32'h8220000;
      11081: inst = 32'h10408000;
      11082: inst = 32'hc4047af;
      11083: inst = 32'h8220000;
      11084: inst = 32'h10408000;
      11085: inst = 32'hc4047bf;
      11086: inst = 32'h8220000;
      11087: inst = 32'h10408000;
      11088: inst = 32'hc40480f;
      11089: inst = 32'h8220000;
      11090: inst = 32'h10408000;
      11091: inst = 32'hc40481f;
      11092: inst = 32'h8220000;
      11093: inst = 32'h10408000;
      11094: inst = 32'hc40486f;
      11095: inst = 32'h8220000;
      11096: inst = 32'h10408000;
      11097: inst = 32'hc40487f;
      11098: inst = 32'h8220000;
      11099: inst = 32'h10408000;
      11100: inst = 32'hc4048cf;
      11101: inst = 32'h8220000;
      11102: inst = 32'h10408000;
      11103: inst = 32'hc4048df;
      11104: inst = 32'h8220000;
      11105: inst = 32'h10408000;
      11106: inst = 32'hc40492f;
      11107: inst = 32'h8220000;
      11108: inst = 32'h10408000;
      11109: inst = 32'hc40493f;
      11110: inst = 32'h8220000;
      11111: inst = 32'h10408000;
      11112: inst = 32'hc40498f;
      11113: inst = 32'h8220000;
      11114: inst = 32'h10408000;
      11115: inst = 32'hc40499f;
      11116: inst = 32'h8220000;
      11117: inst = 32'h10408000;
      11118: inst = 32'hc4049ef;
      11119: inst = 32'h8220000;
      11120: inst = 32'h10408000;
      11121: inst = 32'hc4049ff;
      11122: inst = 32'h8220000;
      11123: inst = 32'h10408000;
      11124: inst = 32'hc404a4f;
      11125: inst = 32'h8220000;
      11126: inst = 32'h10408000;
      11127: inst = 32'hc404a5f;
      11128: inst = 32'h8220000;
      11129: inst = 32'h10408000;
      11130: inst = 32'hc404aaf;
      11131: inst = 32'h8220000;
      11132: inst = 32'h10408000;
      11133: inst = 32'hc404abf;
      11134: inst = 32'h8220000;
      11135: inst = 32'h10408000;
      11136: inst = 32'hc404b0f;
      11137: inst = 32'h8220000;
      11138: inst = 32'h10408000;
      11139: inst = 32'hc404b1f;
      11140: inst = 32'h8220000;
      11141: inst = 32'h10408000;
      11142: inst = 32'hc404b6f;
      11143: inst = 32'h8220000;
      11144: inst = 32'h10408000;
      11145: inst = 32'hc404b7f;
      11146: inst = 32'h8220000;
      11147: inst = 32'h10408000;
      11148: inst = 32'hc404bcf;
      11149: inst = 32'h8220000;
      11150: inst = 32'h10408000;
      11151: inst = 32'hc404bdf;
      11152: inst = 32'h8220000;
      11153: inst = 32'h10408000;
      11154: inst = 32'hc404c2f;
      11155: inst = 32'h8220000;
      11156: inst = 32'h10408000;
      11157: inst = 32'hc404c3f;
      11158: inst = 32'h8220000;
      11159: inst = 32'h10408000;
      11160: inst = 32'hc404c8f;
      11161: inst = 32'h8220000;
      11162: inst = 32'h10408000;
      11163: inst = 32'hc404c9f;
      11164: inst = 32'h8220000;
      11165: inst = 32'h10408000;
      11166: inst = 32'hc404cef;
      11167: inst = 32'h8220000;
      11168: inst = 32'h10408000;
      11169: inst = 32'hc404cff;
      11170: inst = 32'h8220000;
      11171: inst = 32'h10408000;
      11172: inst = 32'hc404d4f;
      11173: inst = 32'h8220000;
      11174: inst = 32'h10408000;
      11175: inst = 32'hc404d5f;
      11176: inst = 32'h8220000;
      11177: inst = 32'h10408000;
      11178: inst = 32'hc404daf;
      11179: inst = 32'h8220000;
      11180: inst = 32'h10408000;
      11181: inst = 32'hc404dbf;
      11182: inst = 32'h8220000;
      11183: inst = 32'h10408000;
      11184: inst = 32'hc404e0f;
      11185: inst = 32'h8220000;
      11186: inst = 32'h10408000;
      11187: inst = 32'hc404e1f;
      11188: inst = 32'h8220000;
      11189: inst = 32'h10408000;
      11190: inst = 32'hc404e6f;
      11191: inst = 32'h8220000;
      11192: inst = 32'h10408000;
      11193: inst = 32'hc404e7f;
      11194: inst = 32'h8220000;
      11195: inst = 32'h10408000;
      11196: inst = 32'hc404ecf;
      11197: inst = 32'h8220000;
      11198: inst = 32'h10408000;
      11199: inst = 32'hc404edf;
      11200: inst = 32'h8220000;
      11201: inst = 32'h10408000;
      11202: inst = 32'hc404f2f;
      11203: inst = 32'h8220000;
      11204: inst = 32'h10408000;
      11205: inst = 32'hc404f3f;
      11206: inst = 32'h8220000;
      11207: inst = 32'h10408000;
      11208: inst = 32'hc404f8f;
      11209: inst = 32'h8220000;
      11210: inst = 32'h10408000;
      11211: inst = 32'hc404f9f;
      11212: inst = 32'h8220000;
      11213: inst = 32'h10408000;
      11214: inst = 32'hc404fef;
      11215: inst = 32'h8220000;
      11216: inst = 32'h10408000;
      11217: inst = 32'hc404fff;
      11218: inst = 32'h8220000;
      11219: inst = 32'h10408000;
      11220: inst = 32'hc40504f;
      11221: inst = 32'h8220000;
      11222: inst = 32'h10408000;
      11223: inst = 32'hc40505f;
      11224: inst = 32'h8220000;
      11225: inst = 32'h10408000;
      11226: inst = 32'hc4050af;
      11227: inst = 32'h8220000;
      11228: inst = 32'h10408000;
      11229: inst = 32'hc4050bf;
      11230: inst = 32'h8220000;
      11231: inst = 32'h10408000;
      11232: inst = 32'hc40510f;
      11233: inst = 32'h8220000;
      11234: inst = 32'h10408000;
      11235: inst = 32'hc40511f;
      11236: inst = 32'h8220000;
      11237: inst = 32'h10408000;
      11238: inst = 32'hc40516f;
      11239: inst = 32'h8220000;
      11240: inst = 32'h10408000;
      11241: inst = 32'hc40517f;
      11242: inst = 32'h8220000;
      11243: inst = 32'h10408000;
      11244: inst = 32'hc4051cf;
      11245: inst = 32'h8220000;
      11246: inst = 32'h10408000;
      11247: inst = 32'hc4051df;
      11248: inst = 32'h8220000;
      11249: inst = 32'h10408000;
      11250: inst = 32'hc40522f;
      11251: inst = 32'h8220000;
      11252: inst = 32'h10408000;
      11253: inst = 32'hc40523f;
      11254: inst = 32'h8220000;
      11255: inst = 32'h10408000;
      11256: inst = 32'hc40528f;
      11257: inst = 32'h8220000;
      11258: inst = 32'h10408000;
      11259: inst = 32'hc40529f;
      11260: inst = 32'h8220000;
      11261: inst = 32'h10408000;
      11262: inst = 32'hc4052ef;
      11263: inst = 32'h8220000;
      11264: inst = 32'h10408000;
      11265: inst = 32'hc4052f0;
      11266: inst = 32'h8220000;
      11267: inst = 32'h10408000;
      11268: inst = 32'hc4052f1;
      11269: inst = 32'h8220000;
      11270: inst = 32'h10408000;
      11271: inst = 32'hc4052f2;
      11272: inst = 32'h8220000;
      11273: inst = 32'h10408000;
      11274: inst = 32'hc4052f3;
      11275: inst = 32'h8220000;
      11276: inst = 32'h10408000;
      11277: inst = 32'hc4052f4;
      11278: inst = 32'h8220000;
      11279: inst = 32'h10408000;
      11280: inst = 32'hc4052f5;
      11281: inst = 32'h8220000;
      11282: inst = 32'h10408000;
      11283: inst = 32'hc4052f6;
      11284: inst = 32'h8220000;
      11285: inst = 32'h10408000;
      11286: inst = 32'hc4052f7;
      11287: inst = 32'h8220000;
      11288: inst = 32'h10408000;
      11289: inst = 32'hc4052f8;
      11290: inst = 32'h8220000;
      11291: inst = 32'h10408000;
      11292: inst = 32'hc4052f9;
      11293: inst = 32'h8220000;
      11294: inst = 32'h10408000;
      11295: inst = 32'hc4052fa;
      11296: inst = 32'h8220000;
      11297: inst = 32'h10408000;
      11298: inst = 32'hc4052fb;
      11299: inst = 32'h8220000;
      11300: inst = 32'h10408000;
      11301: inst = 32'hc4052fc;
      11302: inst = 32'h8220000;
      11303: inst = 32'h10408000;
      11304: inst = 32'hc4052fd;
      11305: inst = 32'h8220000;
      11306: inst = 32'h10408000;
      11307: inst = 32'hc4052fe;
      11308: inst = 32'h8220000;
      11309: inst = 32'h10408000;
      11310: inst = 32'hc4052ff;
      11311: inst = 32'h8220000;
      11312: inst = 32'hc20dbc5;
      11313: inst = 32'h10408000;
      11314: inst = 32'hc404750;
      11315: inst = 32'h8220000;
      11316: inst = 32'h10408000;
      11317: inst = 32'hc404751;
      11318: inst = 32'h8220000;
      11319: inst = 32'h10408000;
      11320: inst = 32'hc404752;
      11321: inst = 32'h8220000;
      11322: inst = 32'h10408000;
      11323: inst = 32'hc404753;
      11324: inst = 32'h8220000;
      11325: inst = 32'h10408000;
      11326: inst = 32'hc404754;
      11327: inst = 32'h8220000;
      11328: inst = 32'h10408000;
      11329: inst = 32'hc404755;
      11330: inst = 32'h8220000;
      11331: inst = 32'h10408000;
      11332: inst = 32'hc404756;
      11333: inst = 32'h8220000;
      11334: inst = 32'h10408000;
      11335: inst = 32'hc404757;
      11336: inst = 32'h8220000;
      11337: inst = 32'h10408000;
      11338: inst = 32'hc404758;
      11339: inst = 32'h8220000;
      11340: inst = 32'h10408000;
      11341: inst = 32'hc404759;
      11342: inst = 32'h8220000;
      11343: inst = 32'h10408000;
      11344: inst = 32'hc40475a;
      11345: inst = 32'h8220000;
      11346: inst = 32'h10408000;
      11347: inst = 32'hc40475b;
      11348: inst = 32'h8220000;
      11349: inst = 32'h10408000;
      11350: inst = 32'hc40475c;
      11351: inst = 32'h8220000;
      11352: inst = 32'h10408000;
      11353: inst = 32'hc40475d;
      11354: inst = 32'h8220000;
      11355: inst = 32'h10408000;
      11356: inst = 32'hc40475e;
      11357: inst = 32'h8220000;
      11358: inst = 32'h10408000;
      11359: inst = 32'hc4047b0;
      11360: inst = 32'h8220000;
      11361: inst = 32'h10408000;
      11362: inst = 32'hc4047b1;
      11363: inst = 32'h8220000;
      11364: inst = 32'h10408000;
      11365: inst = 32'hc4047b2;
      11366: inst = 32'h8220000;
      11367: inst = 32'h10408000;
      11368: inst = 32'hc4047b3;
      11369: inst = 32'h8220000;
      11370: inst = 32'h10408000;
      11371: inst = 32'hc4047b4;
      11372: inst = 32'h8220000;
      11373: inst = 32'h10408000;
      11374: inst = 32'hc4047b5;
      11375: inst = 32'h8220000;
      11376: inst = 32'h10408000;
      11377: inst = 32'hc4047b6;
      11378: inst = 32'h8220000;
      11379: inst = 32'h10408000;
      11380: inst = 32'hc4047b7;
      11381: inst = 32'h8220000;
      11382: inst = 32'h10408000;
      11383: inst = 32'hc4047b8;
      11384: inst = 32'h8220000;
      11385: inst = 32'h10408000;
      11386: inst = 32'hc4047b9;
      11387: inst = 32'h8220000;
      11388: inst = 32'h10408000;
      11389: inst = 32'hc4047ba;
      11390: inst = 32'h8220000;
      11391: inst = 32'h10408000;
      11392: inst = 32'hc4047bb;
      11393: inst = 32'h8220000;
      11394: inst = 32'h10408000;
      11395: inst = 32'hc4047bc;
      11396: inst = 32'h8220000;
      11397: inst = 32'h10408000;
      11398: inst = 32'hc4047bd;
      11399: inst = 32'h8220000;
      11400: inst = 32'h10408000;
      11401: inst = 32'hc4047be;
      11402: inst = 32'h8220000;
      11403: inst = 32'h10408000;
      11404: inst = 32'hc404810;
      11405: inst = 32'h8220000;
      11406: inst = 32'h10408000;
      11407: inst = 32'hc404811;
      11408: inst = 32'h8220000;
      11409: inst = 32'h10408000;
      11410: inst = 32'hc404812;
      11411: inst = 32'h8220000;
      11412: inst = 32'h10408000;
      11413: inst = 32'hc404813;
      11414: inst = 32'h8220000;
      11415: inst = 32'h10408000;
      11416: inst = 32'hc404814;
      11417: inst = 32'h8220000;
      11418: inst = 32'h10408000;
      11419: inst = 32'hc404815;
      11420: inst = 32'h8220000;
      11421: inst = 32'h10408000;
      11422: inst = 32'hc404816;
      11423: inst = 32'h8220000;
      11424: inst = 32'h10408000;
      11425: inst = 32'hc404817;
      11426: inst = 32'h8220000;
      11427: inst = 32'h10408000;
      11428: inst = 32'hc404818;
      11429: inst = 32'h8220000;
      11430: inst = 32'h10408000;
      11431: inst = 32'hc404819;
      11432: inst = 32'h8220000;
      11433: inst = 32'h10408000;
      11434: inst = 32'hc40481a;
      11435: inst = 32'h8220000;
      11436: inst = 32'h10408000;
      11437: inst = 32'hc40481b;
      11438: inst = 32'h8220000;
      11439: inst = 32'h10408000;
      11440: inst = 32'hc40481c;
      11441: inst = 32'h8220000;
      11442: inst = 32'h10408000;
      11443: inst = 32'hc40481d;
      11444: inst = 32'h8220000;
      11445: inst = 32'h10408000;
      11446: inst = 32'hc40481e;
      11447: inst = 32'h8220000;
      11448: inst = 32'h10408000;
      11449: inst = 32'hc404870;
      11450: inst = 32'h8220000;
      11451: inst = 32'h10408000;
      11452: inst = 32'hc404871;
      11453: inst = 32'h8220000;
      11454: inst = 32'h10408000;
      11455: inst = 32'hc404872;
      11456: inst = 32'h8220000;
      11457: inst = 32'h10408000;
      11458: inst = 32'hc404873;
      11459: inst = 32'h8220000;
      11460: inst = 32'h10408000;
      11461: inst = 32'hc404874;
      11462: inst = 32'h8220000;
      11463: inst = 32'h10408000;
      11464: inst = 32'hc404875;
      11465: inst = 32'h8220000;
      11466: inst = 32'h10408000;
      11467: inst = 32'hc404876;
      11468: inst = 32'h8220000;
      11469: inst = 32'h10408000;
      11470: inst = 32'hc404877;
      11471: inst = 32'h8220000;
      11472: inst = 32'h10408000;
      11473: inst = 32'hc404878;
      11474: inst = 32'h8220000;
      11475: inst = 32'h10408000;
      11476: inst = 32'hc404879;
      11477: inst = 32'h8220000;
      11478: inst = 32'h10408000;
      11479: inst = 32'hc40487a;
      11480: inst = 32'h8220000;
      11481: inst = 32'h10408000;
      11482: inst = 32'hc40487b;
      11483: inst = 32'h8220000;
      11484: inst = 32'h10408000;
      11485: inst = 32'hc40487c;
      11486: inst = 32'h8220000;
      11487: inst = 32'h10408000;
      11488: inst = 32'hc40487d;
      11489: inst = 32'h8220000;
      11490: inst = 32'h10408000;
      11491: inst = 32'hc40487e;
      11492: inst = 32'h8220000;
      11493: inst = 32'h10408000;
      11494: inst = 32'hc4048d0;
      11495: inst = 32'h8220000;
      11496: inst = 32'h10408000;
      11497: inst = 32'hc4048d1;
      11498: inst = 32'h8220000;
      11499: inst = 32'h10408000;
      11500: inst = 32'hc4048d2;
      11501: inst = 32'h8220000;
      11502: inst = 32'h10408000;
      11503: inst = 32'hc4048d3;
      11504: inst = 32'h8220000;
      11505: inst = 32'h10408000;
      11506: inst = 32'hc4048d4;
      11507: inst = 32'h8220000;
      11508: inst = 32'h10408000;
      11509: inst = 32'hc4048d5;
      11510: inst = 32'h8220000;
      11511: inst = 32'h10408000;
      11512: inst = 32'hc4048d6;
      11513: inst = 32'h8220000;
      11514: inst = 32'h10408000;
      11515: inst = 32'hc4048d7;
      11516: inst = 32'h8220000;
      11517: inst = 32'h10408000;
      11518: inst = 32'hc4048d8;
      11519: inst = 32'h8220000;
      11520: inst = 32'h10408000;
      11521: inst = 32'hc4048d9;
      11522: inst = 32'h8220000;
      11523: inst = 32'h10408000;
      11524: inst = 32'hc4048da;
      11525: inst = 32'h8220000;
      11526: inst = 32'h10408000;
      11527: inst = 32'hc4048db;
      11528: inst = 32'h8220000;
      11529: inst = 32'h10408000;
      11530: inst = 32'hc4048dc;
      11531: inst = 32'h8220000;
      11532: inst = 32'h10408000;
      11533: inst = 32'hc4048dd;
      11534: inst = 32'h8220000;
      11535: inst = 32'h10408000;
      11536: inst = 32'hc4048de;
      11537: inst = 32'h8220000;
      11538: inst = 32'h10408000;
      11539: inst = 32'hc404930;
      11540: inst = 32'h8220000;
      11541: inst = 32'h10408000;
      11542: inst = 32'hc404931;
      11543: inst = 32'h8220000;
      11544: inst = 32'h10408000;
      11545: inst = 32'hc404936;
      11546: inst = 32'h8220000;
      11547: inst = 32'h10408000;
      11548: inst = 32'hc404937;
      11549: inst = 32'h8220000;
      11550: inst = 32'h10408000;
      11551: inst = 32'hc404938;
      11552: inst = 32'h8220000;
      11553: inst = 32'h10408000;
      11554: inst = 32'hc404939;
      11555: inst = 32'h8220000;
      11556: inst = 32'h10408000;
      11557: inst = 32'hc40493a;
      11558: inst = 32'h8220000;
      11559: inst = 32'h10408000;
      11560: inst = 32'hc40493b;
      11561: inst = 32'h8220000;
      11562: inst = 32'h10408000;
      11563: inst = 32'hc40493c;
      11564: inst = 32'h8220000;
      11565: inst = 32'h10408000;
      11566: inst = 32'hc40493d;
      11567: inst = 32'h8220000;
      11568: inst = 32'h10408000;
      11569: inst = 32'hc40493e;
      11570: inst = 32'h8220000;
      11571: inst = 32'h10408000;
      11572: inst = 32'hc404990;
      11573: inst = 32'h8220000;
      11574: inst = 32'h10408000;
      11575: inst = 32'hc404991;
      11576: inst = 32'h8220000;
      11577: inst = 32'h10408000;
      11578: inst = 32'hc404996;
      11579: inst = 32'h8220000;
      11580: inst = 32'h10408000;
      11581: inst = 32'hc404997;
      11582: inst = 32'h8220000;
      11583: inst = 32'h10408000;
      11584: inst = 32'hc404998;
      11585: inst = 32'h8220000;
      11586: inst = 32'h10408000;
      11587: inst = 32'hc404999;
      11588: inst = 32'h8220000;
      11589: inst = 32'h10408000;
      11590: inst = 32'hc40499a;
      11591: inst = 32'h8220000;
      11592: inst = 32'h10408000;
      11593: inst = 32'hc40499b;
      11594: inst = 32'h8220000;
      11595: inst = 32'h10408000;
      11596: inst = 32'hc40499c;
      11597: inst = 32'h8220000;
      11598: inst = 32'h10408000;
      11599: inst = 32'hc40499d;
      11600: inst = 32'h8220000;
      11601: inst = 32'h10408000;
      11602: inst = 32'hc40499e;
      11603: inst = 32'h8220000;
      11604: inst = 32'h10408000;
      11605: inst = 32'hc4049f0;
      11606: inst = 32'h8220000;
      11607: inst = 32'h10408000;
      11608: inst = 32'hc4049f1;
      11609: inst = 32'h8220000;
      11610: inst = 32'h10408000;
      11611: inst = 32'hc4049f6;
      11612: inst = 32'h8220000;
      11613: inst = 32'h10408000;
      11614: inst = 32'hc4049f7;
      11615: inst = 32'h8220000;
      11616: inst = 32'h10408000;
      11617: inst = 32'hc4049f8;
      11618: inst = 32'h8220000;
      11619: inst = 32'h10408000;
      11620: inst = 32'hc4049f9;
      11621: inst = 32'h8220000;
      11622: inst = 32'h10408000;
      11623: inst = 32'hc4049fa;
      11624: inst = 32'h8220000;
      11625: inst = 32'h10408000;
      11626: inst = 32'hc4049fb;
      11627: inst = 32'h8220000;
      11628: inst = 32'h10408000;
      11629: inst = 32'hc4049fc;
      11630: inst = 32'h8220000;
      11631: inst = 32'h10408000;
      11632: inst = 32'hc4049fd;
      11633: inst = 32'h8220000;
      11634: inst = 32'h10408000;
      11635: inst = 32'hc4049fe;
      11636: inst = 32'h8220000;
      11637: inst = 32'h10408000;
      11638: inst = 32'hc404a50;
      11639: inst = 32'h8220000;
      11640: inst = 32'h10408000;
      11641: inst = 32'hc404a51;
      11642: inst = 32'h8220000;
      11643: inst = 32'h10408000;
      11644: inst = 32'hc404a56;
      11645: inst = 32'h8220000;
      11646: inst = 32'h10408000;
      11647: inst = 32'hc404a57;
      11648: inst = 32'h8220000;
      11649: inst = 32'h10408000;
      11650: inst = 32'hc404a58;
      11651: inst = 32'h8220000;
      11652: inst = 32'h10408000;
      11653: inst = 32'hc404a59;
      11654: inst = 32'h8220000;
      11655: inst = 32'h10408000;
      11656: inst = 32'hc404a5a;
      11657: inst = 32'h8220000;
      11658: inst = 32'h10408000;
      11659: inst = 32'hc404a5b;
      11660: inst = 32'h8220000;
      11661: inst = 32'h10408000;
      11662: inst = 32'hc404a5c;
      11663: inst = 32'h8220000;
      11664: inst = 32'h10408000;
      11665: inst = 32'hc404a5d;
      11666: inst = 32'h8220000;
      11667: inst = 32'h10408000;
      11668: inst = 32'hc404a5e;
      11669: inst = 32'h8220000;
      11670: inst = 32'h10408000;
      11671: inst = 32'hc404ab0;
      11672: inst = 32'h8220000;
      11673: inst = 32'h10408000;
      11674: inst = 32'hc404ab1;
      11675: inst = 32'h8220000;
      11676: inst = 32'h10408000;
      11677: inst = 32'hc404ab6;
      11678: inst = 32'h8220000;
      11679: inst = 32'h10408000;
      11680: inst = 32'hc404ab7;
      11681: inst = 32'h8220000;
      11682: inst = 32'h10408000;
      11683: inst = 32'hc404ab8;
      11684: inst = 32'h8220000;
      11685: inst = 32'h10408000;
      11686: inst = 32'hc404ab9;
      11687: inst = 32'h8220000;
      11688: inst = 32'h10408000;
      11689: inst = 32'hc404aba;
      11690: inst = 32'h8220000;
      11691: inst = 32'h10408000;
      11692: inst = 32'hc404abb;
      11693: inst = 32'h8220000;
      11694: inst = 32'h10408000;
      11695: inst = 32'hc404abc;
      11696: inst = 32'h8220000;
      11697: inst = 32'h10408000;
      11698: inst = 32'hc404abd;
      11699: inst = 32'h8220000;
      11700: inst = 32'h10408000;
      11701: inst = 32'hc404abe;
      11702: inst = 32'h8220000;
      11703: inst = 32'h10408000;
      11704: inst = 32'hc404b10;
      11705: inst = 32'h8220000;
      11706: inst = 32'h10408000;
      11707: inst = 32'hc404b11;
      11708: inst = 32'h8220000;
      11709: inst = 32'h10408000;
      11710: inst = 32'hc404b16;
      11711: inst = 32'h8220000;
      11712: inst = 32'h10408000;
      11713: inst = 32'hc404b17;
      11714: inst = 32'h8220000;
      11715: inst = 32'h10408000;
      11716: inst = 32'hc404b18;
      11717: inst = 32'h8220000;
      11718: inst = 32'h10408000;
      11719: inst = 32'hc404b19;
      11720: inst = 32'h8220000;
      11721: inst = 32'h10408000;
      11722: inst = 32'hc404b1a;
      11723: inst = 32'h8220000;
      11724: inst = 32'h10408000;
      11725: inst = 32'hc404b1b;
      11726: inst = 32'h8220000;
      11727: inst = 32'h10408000;
      11728: inst = 32'hc404b1c;
      11729: inst = 32'h8220000;
      11730: inst = 32'h10408000;
      11731: inst = 32'hc404b1d;
      11732: inst = 32'h8220000;
      11733: inst = 32'h10408000;
      11734: inst = 32'hc404b1e;
      11735: inst = 32'h8220000;
      11736: inst = 32'h10408000;
      11737: inst = 32'hc404b70;
      11738: inst = 32'h8220000;
      11739: inst = 32'h10408000;
      11740: inst = 32'hc404b71;
      11741: inst = 32'h8220000;
      11742: inst = 32'h10408000;
      11743: inst = 32'hc404b76;
      11744: inst = 32'h8220000;
      11745: inst = 32'h10408000;
      11746: inst = 32'hc404b77;
      11747: inst = 32'h8220000;
      11748: inst = 32'h10408000;
      11749: inst = 32'hc404b78;
      11750: inst = 32'h8220000;
      11751: inst = 32'h10408000;
      11752: inst = 32'hc404b79;
      11753: inst = 32'h8220000;
      11754: inst = 32'h10408000;
      11755: inst = 32'hc404b7a;
      11756: inst = 32'h8220000;
      11757: inst = 32'h10408000;
      11758: inst = 32'hc404b7b;
      11759: inst = 32'h8220000;
      11760: inst = 32'h10408000;
      11761: inst = 32'hc404b7c;
      11762: inst = 32'h8220000;
      11763: inst = 32'h10408000;
      11764: inst = 32'hc404b7d;
      11765: inst = 32'h8220000;
      11766: inst = 32'h10408000;
      11767: inst = 32'hc404b7e;
      11768: inst = 32'h8220000;
      11769: inst = 32'h10408000;
      11770: inst = 32'hc404bd0;
      11771: inst = 32'h8220000;
      11772: inst = 32'h10408000;
      11773: inst = 32'hc404bd1;
      11774: inst = 32'h8220000;
      11775: inst = 32'h10408000;
      11776: inst = 32'hc404bd2;
      11777: inst = 32'h8220000;
      11778: inst = 32'h10408000;
      11779: inst = 32'hc404bd3;
      11780: inst = 32'h8220000;
      11781: inst = 32'h10408000;
      11782: inst = 32'hc404bd4;
      11783: inst = 32'h8220000;
      11784: inst = 32'h10408000;
      11785: inst = 32'hc404bd5;
      11786: inst = 32'h8220000;
      11787: inst = 32'h10408000;
      11788: inst = 32'hc404bd6;
      11789: inst = 32'h8220000;
      11790: inst = 32'h10408000;
      11791: inst = 32'hc404bd7;
      11792: inst = 32'h8220000;
      11793: inst = 32'h10408000;
      11794: inst = 32'hc404bd8;
      11795: inst = 32'h8220000;
      11796: inst = 32'h10408000;
      11797: inst = 32'hc404bd9;
      11798: inst = 32'h8220000;
      11799: inst = 32'h10408000;
      11800: inst = 32'hc404bda;
      11801: inst = 32'h8220000;
      11802: inst = 32'h10408000;
      11803: inst = 32'hc404bdb;
      11804: inst = 32'h8220000;
      11805: inst = 32'h10408000;
      11806: inst = 32'hc404bdc;
      11807: inst = 32'h8220000;
      11808: inst = 32'h10408000;
      11809: inst = 32'hc404bdd;
      11810: inst = 32'h8220000;
      11811: inst = 32'h10408000;
      11812: inst = 32'hc404bde;
      11813: inst = 32'h8220000;
      11814: inst = 32'h10408000;
      11815: inst = 32'hc404c30;
      11816: inst = 32'h8220000;
      11817: inst = 32'h10408000;
      11818: inst = 32'hc404c31;
      11819: inst = 32'h8220000;
      11820: inst = 32'h10408000;
      11821: inst = 32'hc404c32;
      11822: inst = 32'h8220000;
      11823: inst = 32'h10408000;
      11824: inst = 32'hc404c33;
      11825: inst = 32'h8220000;
      11826: inst = 32'h10408000;
      11827: inst = 32'hc404c34;
      11828: inst = 32'h8220000;
      11829: inst = 32'h10408000;
      11830: inst = 32'hc404c35;
      11831: inst = 32'h8220000;
      11832: inst = 32'h10408000;
      11833: inst = 32'hc404c36;
      11834: inst = 32'h8220000;
      11835: inst = 32'h10408000;
      11836: inst = 32'hc404c37;
      11837: inst = 32'h8220000;
      11838: inst = 32'h10408000;
      11839: inst = 32'hc404c38;
      11840: inst = 32'h8220000;
      11841: inst = 32'h10408000;
      11842: inst = 32'hc404c39;
      11843: inst = 32'h8220000;
      11844: inst = 32'h10408000;
      11845: inst = 32'hc404c3a;
      11846: inst = 32'h8220000;
      11847: inst = 32'h10408000;
      11848: inst = 32'hc404c3b;
      11849: inst = 32'h8220000;
      11850: inst = 32'h10408000;
      11851: inst = 32'hc404c3c;
      11852: inst = 32'h8220000;
      11853: inst = 32'h10408000;
      11854: inst = 32'hc404c3d;
      11855: inst = 32'h8220000;
      11856: inst = 32'h10408000;
      11857: inst = 32'hc404c3e;
      11858: inst = 32'h8220000;
      11859: inst = 32'h10408000;
      11860: inst = 32'hc404c90;
      11861: inst = 32'h8220000;
      11862: inst = 32'h10408000;
      11863: inst = 32'hc404c91;
      11864: inst = 32'h8220000;
      11865: inst = 32'h10408000;
      11866: inst = 32'hc404c92;
      11867: inst = 32'h8220000;
      11868: inst = 32'h10408000;
      11869: inst = 32'hc404c93;
      11870: inst = 32'h8220000;
      11871: inst = 32'h10408000;
      11872: inst = 32'hc404c94;
      11873: inst = 32'h8220000;
      11874: inst = 32'h10408000;
      11875: inst = 32'hc404c95;
      11876: inst = 32'h8220000;
      11877: inst = 32'h10408000;
      11878: inst = 32'hc404c96;
      11879: inst = 32'h8220000;
      11880: inst = 32'h10408000;
      11881: inst = 32'hc404c97;
      11882: inst = 32'h8220000;
      11883: inst = 32'h10408000;
      11884: inst = 32'hc404c98;
      11885: inst = 32'h8220000;
      11886: inst = 32'h10408000;
      11887: inst = 32'hc404c99;
      11888: inst = 32'h8220000;
      11889: inst = 32'h10408000;
      11890: inst = 32'hc404c9a;
      11891: inst = 32'h8220000;
      11892: inst = 32'h10408000;
      11893: inst = 32'hc404c9b;
      11894: inst = 32'h8220000;
      11895: inst = 32'h10408000;
      11896: inst = 32'hc404c9c;
      11897: inst = 32'h8220000;
      11898: inst = 32'h10408000;
      11899: inst = 32'hc404c9d;
      11900: inst = 32'h8220000;
      11901: inst = 32'h10408000;
      11902: inst = 32'hc404c9e;
      11903: inst = 32'h8220000;
      11904: inst = 32'h10408000;
      11905: inst = 32'hc404cf0;
      11906: inst = 32'h8220000;
      11907: inst = 32'h10408000;
      11908: inst = 32'hc404cf1;
      11909: inst = 32'h8220000;
      11910: inst = 32'h10408000;
      11911: inst = 32'hc404cf2;
      11912: inst = 32'h8220000;
      11913: inst = 32'h10408000;
      11914: inst = 32'hc404cf3;
      11915: inst = 32'h8220000;
      11916: inst = 32'h10408000;
      11917: inst = 32'hc404cf4;
      11918: inst = 32'h8220000;
      11919: inst = 32'h10408000;
      11920: inst = 32'hc404cf5;
      11921: inst = 32'h8220000;
      11922: inst = 32'h10408000;
      11923: inst = 32'hc404cf6;
      11924: inst = 32'h8220000;
      11925: inst = 32'h10408000;
      11926: inst = 32'hc404cf7;
      11927: inst = 32'h8220000;
      11928: inst = 32'h10408000;
      11929: inst = 32'hc404cf8;
      11930: inst = 32'h8220000;
      11931: inst = 32'h10408000;
      11932: inst = 32'hc404cf9;
      11933: inst = 32'h8220000;
      11934: inst = 32'h10408000;
      11935: inst = 32'hc404cfa;
      11936: inst = 32'h8220000;
      11937: inst = 32'h10408000;
      11938: inst = 32'hc404cfe;
      11939: inst = 32'h8220000;
      11940: inst = 32'h10408000;
      11941: inst = 32'hc404d50;
      11942: inst = 32'h8220000;
      11943: inst = 32'h10408000;
      11944: inst = 32'hc404d51;
      11945: inst = 32'h8220000;
      11946: inst = 32'h10408000;
      11947: inst = 32'hc404d52;
      11948: inst = 32'h8220000;
      11949: inst = 32'h10408000;
      11950: inst = 32'hc404d53;
      11951: inst = 32'h8220000;
      11952: inst = 32'h10408000;
      11953: inst = 32'hc404d54;
      11954: inst = 32'h8220000;
      11955: inst = 32'h10408000;
      11956: inst = 32'hc404d55;
      11957: inst = 32'h8220000;
      11958: inst = 32'h10408000;
      11959: inst = 32'hc404d56;
      11960: inst = 32'h8220000;
      11961: inst = 32'h10408000;
      11962: inst = 32'hc404d57;
      11963: inst = 32'h8220000;
      11964: inst = 32'h10408000;
      11965: inst = 32'hc404d58;
      11966: inst = 32'h8220000;
      11967: inst = 32'h10408000;
      11968: inst = 32'hc404d59;
      11969: inst = 32'h8220000;
      11970: inst = 32'h10408000;
      11971: inst = 32'hc404d5a;
      11972: inst = 32'h8220000;
      11973: inst = 32'h10408000;
      11974: inst = 32'hc404d5c;
      11975: inst = 32'h8220000;
      11976: inst = 32'h10408000;
      11977: inst = 32'hc404d5d;
      11978: inst = 32'h8220000;
      11979: inst = 32'h10408000;
      11980: inst = 32'hc404d5e;
      11981: inst = 32'h8220000;
      11982: inst = 32'h10408000;
      11983: inst = 32'hc404db0;
      11984: inst = 32'h8220000;
      11985: inst = 32'h10408000;
      11986: inst = 32'hc404db1;
      11987: inst = 32'h8220000;
      11988: inst = 32'h10408000;
      11989: inst = 32'hc404db2;
      11990: inst = 32'h8220000;
      11991: inst = 32'h10408000;
      11992: inst = 32'hc404db3;
      11993: inst = 32'h8220000;
      11994: inst = 32'h10408000;
      11995: inst = 32'hc404db4;
      11996: inst = 32'h8220000;
      11997: inst = 32'h10408000;
      11998: inst = 32'hc404db5;
      11999: inst = 32'h8220000;
      12000: inst = 32'h10408000;
      12001: inst = 32'hc404db6;
      12002: inst = 32'h8220000;
      12003: inst = 32'h10408000;
      12004: inst = 32'hc404db7;
      12005: inst = 32'h8220000;
      12006: inst = 32'h10408000;
      12007: inst = 32'hc404db8;
      12008: inst = 32'h8220000;
      12009: inst = 32'h10408000;
      12010: inst = 32'hc404db9;
      12011: inst = 32'h8220000;
      12012: inst = 32'h10408000;
      12013: inst = 32'hc404dba;
      12014: inst = 32'h8220000;
      12015: inst = 32'h10408000;
      12016: inst = 32'hc404dbb;
      12017: inst = 32'h8220000;
      12018: inst = 32'h10408000;
      12019: inst = 32'hc404dbc;
      12020: inst = 32'h8220000;
      12021: inst = 32'h10408000;
      12022: inst = 32'hc404dbd;
      12023: inst = 32'h8220000;
      12024: inst = 32'h10408000;
      12025: inst = 32'hc404dbe;
      12026: inst = 32'h8220000;
      12027: inst = 32'h10408000;
      12028: inst = 32'hc404e10;
      12029: inst = 32'h8220000;
      12030: inst = 32'h10408000;
      12031: inst = 32'hc404e11;
      12032: inst = 32'h8220000;
      12033: inst = 32'h10408000;
      12034: inst = 32'hc404e12;
      12035: inst = 32'h8220000;
      12036: inst = 32'h10408000;
      12037: inst = 32'hc404e13;
      12038: inst = 32'h8220000;
      12039: inst = 32'h10408000;
      12040: inst = 32'hc404e14;
      12041: inst = 32'h8220000;
      12042: inst = 32'h10408000;
      12043: inst = 32'hc404e15;
      12044: inst = 32'h8220000;
      12045: inst = 32'h10408000;
      12046: inst = 32'hc404e16;
      12047: inst = 32'h8220000;
      12048: inst = 32'h10408000;
      12049: inst = 32'hc404e17;
      12050: inst = 32'h8220000;
      12051: inst = 32'h10408000;
      12052: inst = 32'hc404e18;
      12053: inst = 32'h8220000;
      12054: inst = 32'h10408000;
      12055: inst = 32'hc404e19;
      12056: inst = 32'h8220000;
      12057: inst = 32'h10408000;
      12058: inst = 32'hc404e1a;
      12059: inst = 32'h8220000;
      12060: inst = 32'h10408000;
      12061: inst = 32'hc404e1b;
      12062: inst = 32'h8220000;
      12063: inst = 32'h10408000;
      12064: inst = 32'hc404e1c;
      12065: inst = 32'h8220000;
      12066: inst = 32'h10408000;
      12067: inst = 32'hc404e1d;
      12068: inst = 32'h8220000;
      12069: inst = 32'h10408000;
      12070: inst = 32'hc404e1e;
      12071: inst = 32'h8220000;
      12072: inst = 32'h10408000;
      12073: inst = 32'hc404e70;
      12074: inst = 32'h8220000;
      12075: inst = 32'h10408000;
      12076: inst = 32'hc404e71;
      12077: inst = 32'h8220000;
      12078: inst = 32'h10408000;
      12079: inst = 32'hc404e72;
      12080: inst = 32'h8220000;
      12081: inst = 32'h10408000;
      12082: inst = 32'hc404e73;
      12083: inst = 32'h8220000;
      12084: inst = 32'h10408000;
      12085: inst = 32'hc404e74;
      12086: inst = 32'h8220000;
      12087: inst = 32'h10408000;
      12088: inst = 32'hc404e75;
      12089: inst = 32'h8220000;
      12090: inst = 32'h10408000;
      12091: inst = 32'hc404e76;
      12092: inst = 32'h8220000;
      12093: inst = 32'h10408000;
      12094: inst = 32'hc404e77;
      12095: inst = 32'h8220000;
      12096: inst = 32'h10408000;
      12097: inst = 32'hc404e78;
      12098: inst = 32'h8220000;
      12099: inst = 32'h10408000;
      12100: inst = 32'hc404e79;
      12101: inst = 32'h8220000;
      12102: inst = 32'h10408000;
      12103: inst = 32'hc404e7a;
      12104: inst = 32'h8220000;
      12105: inst = 32'h10408000;
      12106: inst = 32'hc404e7b;
      12107: inst = 32'h8220000;
      12108: inst = 32'h10408000;
      12109: inst = 32'hc404e7c;
      12110: inst = 32'h8220000;
      12111: inst = 32'h10408000;
      12112: inst = 32'hc404e7d;
      12113: inst = 32'h8220000;
      12114: inst = 32'h10408000;
      12115: inst = 32'hc404e7e;
      12116: inst = 32'h8220000;
      12117: inst = 32'h10408000;
      12118: inst = 32'hc404ed0;
      12119: inst = 32'h8220000;
      12120: inst = 32'h10408000;
      12121: inst = 32'hc404ed1;
      12122: inst = 32'h8220000;
      12123: inst = 32'h10408000;
      12124: inst = 32'hc404ed2;
      12125: inst = 32'h8220000;
      12126: inst = 32'h10408000;
      12127: inst = 32'hc404ed3;
      12128: inst = 32'h8220000;
      12129: inst = 32'h10408000;
      12130: inst = 32'hc404ed4;
      12131: inst = 32'h8220000;
      12132: inst = 32'h10408000;
      12133: inst = 32'hc404ed5;
      12134: inst = 32'h8220000;
      12135: inst = 32'h10408000;
      12136: inst = 32'hc404ed6;
      12137: inst = 32'h8220000;
      12138: inst = 32'h10408000;
      12139: inst = 32'hc404ed7;
      12140: inst = 32'h8220000;
      12141: inst = 32'h10408000;
      12142: inst = 32'hc404ed8;
      12143: inst = 32'h8220000;
      12144: inst = 32'h10408000;
      12145: inst = 32'hc404ed9;
      12146: inst = 32'h8220000;
      12147: inst = 32'h10408000;
      12148: inst = 32'hc404eda;
      12149: inst = 32'h8220000;
      12150: inst = 32'h10408000;
      12151: inst = 32'hc404edb;
      12152: inst = 32'h8220000;
      12153: inst = 32'h10408000;
      12154: inst = 32'hc404edc;
      12155: inst = 32'h8220000;
      12156: inst = 32'h10408000;
      12157: inst = 32'hc404edd;
      12158: inst = 32'h8220000;
      12159: inst = 32'h10408000;
      12160: inst = 32'hc404ede;
      12161: inst = 32'h8220000;
      12162: inst = 32'h10408000;
      12163: inst = 32'hc404f30;
      12164: inst = 32'h8220000;
      12165: inst = 32'h10408000;
      12166: inst = 32'hc404f31;
      12167: inst = 32'h8220000;
      12168: inst = 32'h10408000;
      12169: inst = 32'hc404f32;
      12170: inst = 32'h8220000;
      12171: inst = 32'h10408000;
      12172: inst = 32'hc404f33;
      12173: inst = 32'h8220000;
      12174: inst = 32'h10408000;
      12175: inst = 32'hc404f34;
      12176: inst = 32'h8220000;
      12177: inst = 32'h10408000;
      12178: inst = 32'hc404f35;
      12179: inst = 32'h8220000;
      12180: inst = 32'h10408000;
      12181: inst = 32'hc404f36;
      12182: inst = 32'h8220000;
      12183: inst = 32'h10408000;
      12184: inst = 32'hc404f37;
      12185: inst = 32'h8220000;
      12186: inst = 32'h10408000;
      12187: inst = 32'hc404f38;
      12188: inst = 32'h8220000;
      12189: inst = 32'h10408000;
      12190: inst = 32'hc404f39;
      12191: inst = 32'h8220000;
      12192: inst = 32'h10408000;
      12193: inst = 32'hc404f3a;
      12194: inst = 32'h8220000;
      12195: inst = 32'h10408000;
      12196: inst = 32'hc404f3b;
      12197: inst = 32'h8220000;
      12198: inst = 32'h10408000;
      12199: inst = 32'hc404f3c;
      12200: inst = 32'h8220000;
      12201: inst = 32'h10408000;
      12202: inst = 32'hc404f3d;
      12203: inst = 32'h8220000;
      12204: inst = 32'h10408000;
      12205: inst = 32'hc404f3e;
      12206: inst = 32'h8220000;
      12207: inst = 32'h10408000;
      12208: inst = 32'hc404f90;
      12209: inst = 32'h8220000;
      12210: inst = 32'h10408000;
      12211: inst = 32'hc404f91;
      12212: inst = 32'h8220000;
      12213: inst = 32'h10408000;
      12214: inst = 32'hc404f92;
      12215: inst = 32'h8220000;
      12216: inst = 32'h10408000;
      12217: inst = 32'hc404f93;
      12218: inst = 32'h8220000;
      12219: inst = 32'h10408000;
      12220: inst = 32'hc404f94;
      12221: inst = 32'h8220000;
      12222: inst = 32'h10408000;
      12223: inst = 32'hc404f95;
      12224: inst = 32'h8220000;
      12225: inst = 32'h10408000;
      12226: inst = 32'hc404f96;
      12227: inst = 32'h8220000;
      12228: inst = 32'h10408000;
      12229: inst = 32'hc404f97;
      12230: inst = 32'h8220000;
      12231: inst = 32'h10408000;
      12232: inst = 32'hc404f98;
      12233: inst = 32'h8220000;
      12234: inst = 32'h10408000;
      12235: inst = 32'hc404f99;
      12236: inst = 32'h8220000;
      12237: inst = 32'h10408000;
      12238: inst = 32'hc404f9a;
      12239: inst = 32'h8220000;
      12240: inst = 32'h10408000;
      12241: inst = 32'hc404f9b;
      12242: inst = 32'h8220000;
      12243: inst = 32'h10408000;
      12244: inst = 32'hc404f9c;
      12245: inst = 32'h8220000;
      12246: inst = 32'h10408000;
      12247: inst = 32'hc404f9d;
      12248: inst = 32'h8220000;
      12249: inst = 32'h10408000;
      12250: inst = 32'hc404f9e;
      12251: inst = 32'h8220000;
      12252: inst = 32'h10408000;
      12253: inst = 32'hc404ff0;
      12254: inst = 32'h8220000;
      12255: inst = 32'h10408000;
      12256: inst = 32'hc404ff1;
      12257: inst = 32'h8220000;
      12258: inst = 32'h10408000;
      12259: inst = 32'hc404ff2;
      12260: inst = 32'h8220000;
      12261: inst = 32'h10408000;
      12262: inst = 32'hc404ff3;
      12263: inst = 32'h8220000;
      12264: inst = 32'h10408000;
      12265: inst = 32'hc404ff4;
      12266: inst = 32'h8220000;
      12267: inst = 32'h10408000;
      12268: inst = 32'hc404ff5;
      12269: inst = 32'h8220000;
      12270: inst = 32'h10408000;
      12271: inst = 32'hc404ff6;
      12272: inst = 32'h8220000;
      12273: inst = 32'h10408000;
      12274: inst = 32'hc404ff7;
      12275: inst = 32'h8220000;
      12276: inst = 32'h10408000;
      12277: inst = 32'hc404ff8;
      12278: inst = 32'h8220000;
      12279: inst = 32'h10408000;
      12280: inst = 32'hc404ff9;
      12281: inst = 32'h8220000;
      12282: inst = 32'h10408000;
      12283: inst = 32'hc404ffa;
      12284: inst = 32'h8220000;
      12285: inst = 32'h10408000;
      12286: inst = 32'hc404ffb;
      12287: inst = 32'h8220000;
      12288: inst = 32'h10408000;
      12289: inst = 32'hc404ffc;
      12290: inst = 32'h8220000;
      12291: inst = 32'h10408000;
      12292: inst = 32'hc404ffd;
      12293: inst = 32'h8220000;
      12294: inst = 32'h10408000;
      12295: inst = 32'hc404ffe;
      12296: inst = 32'h8220000;
      12297: inst = 32'h10408000;
      12298: inst = 32'hc405050;
      12299: inst = 32'h8220000;
      12300: inst = 32'h10408000;
      12301: inst = 32'hc405051;
      12302: inst = 32'h8220000;
      12303: inst = 32'h10408000;
      12304: inst = 32'hc405052;
      12305: inst = 32'h8220000;
      12306: inst = 32'h10408000;
      12307: inst = 32'hc405053;
      12308: inst = 32'h8220000;
      12309: inst = 32'h10408000;
      12310: inst = 32'hc405054;
      12311: inst = 32'h8220000;
      12312: inst = 32'h10408000;
      12313: inst = 32'hc405055;
      12314: inst = 32'h8220000;
      12315: inst = 32'h10408000;
      12316: inst = 32'hc405056;
      12317: inst = 32'h8220000;
      12318: inst = 32'h10408000;
      12319: inst = 32'hc405057;
      12320: inst = 32'h8220000;
      12321: inst = 32'h10408000;
      12322: inst = 32'hc405058;
      12323: inst = 32'h8220000;
      12324: inst = 32'h10408000;
      12325: inst = 32'hc405059;
      12326: inst = 32'h8220000;
      12327: inst = 32'h10408000;
      12328: inst = 32'hc40505a;
      12329: inst = 32'h8220000;
      12330: inst = 32'h10408000;
      12331: inst = 32'hc40505b;
      12332: inst = 32'h8220000;
      12333: inst = 32'h10408000;
      12334: inst = 32'hc40505c;
      12335: inst = 32'h8220000;
      12336: inst = 32'h10408000;
      12337: inst = 32'hc40505d;
      12338: inst = 32'h8220000;
      12339: inst = 32'h10408000;
      12340: inst = 32'hc40505e;
      12341: inst = 32'h8220000;
      12342: inst = 32'h10408000;
      12343: inst = 32'hc4050b0;
      12344: inst = 32'h8220000;
      12345: inst = 32'h10408000;
      12346: inst = 32'hc4050b1;
      12347: inst = 32'h8220000;
      12348: inst = 32'h10408000;
      12349: inst = 32'hc4050b2;
      12350: inst = 32'h8220000;
      12351: inst = 32'h10408000;
      12352: inst = 32'hc4050b3;
      12353: inst = 32'h8220000;
      12354: inst = 32'h10408000;
      12355: inst = 32'hc4050b4;
      12356: inst = 32'h8220000;
      12357: inst = 32'h10408000;
      12358: inst = 32'hc4050b5;
      12359: inst = 32'h8220000;
      12360: inst = 32'h10408000;
      12361: inst = 32'hc4050b6;
      12362: inst = 32'h8220000;
      12363: inst = 32'h10408000;
      12364: inst = 32'hc4050b7;
      12365: inst = 32'h8220000;
      12366: inst = 32'h10408000;
      12367: inst = 32'hc4050b8;
      12368: inst = 32'h8220000;
      12369: inst = 32'h10408000;
      12370: inst = 32'hc4050b9;
      12371: inst = 32'h8220000;
      12372: inst = 32'h10408000;
      12373: inst = 32'hc4050ba;
      12374: inst = 32'h8220000;
      12375: inst = 32'h10408000;
      12376: inst = 32'hc4050bb;
      12377: inst = 32'h8220000;
      12378: inst = 32'h10408000;
      12379: inst = 32'hc4050bc;
      12380: inst = 32'h8220000;
      12381: inst = 32'h10408000;
      12382: inst = 32'hc4050bd;
      12383: inst = 32'h8220000;
      12384: inst = 32'h10408000;
      12385: inst = 32'hc4050be;
      12386: inst = 32'h8220000;
      12387: inst = 32'h10408000;
      12388: inst = 32'hc405110;
      12389: inst = 32'h8220000;
      12390: inst = 32'h10408000;
      12391: inst = 32'hc405111;
      12392: inst = 32'h8220000;
      12393: inst = 32'h10408000;
      12394: inst = 32'hc405112;
      12395: inst = 32'h8220000;
      12396: inst = 32'h10408000;
      12397: inst = 32'hc405113;
      12398: inst = 32'h8220000;
      12399: inst = 32'h10408000;
      12400: inst = 32'hc405114;
      12401: inst = 32'h8220000;
      12402: inst = 32'h10408000;
      12403: inst = 32'hc405115;
      12404: inst = 32'h8220000;
      12405: inst = 32'h10408000;
      12406: inst = 32'hc405116;
      12407: inst = 32'h8220000;
      12408: inst = 32'h10408000;
      12409: inst = 32'hc405117;
      12410: inst = 32'h8220000;
      12411: inst = 32'h10408000;
      12412: inst = 32'hc405118;
      12413: inst = 32'h8220000;
      12414: inst = 32'h10408000;
      12415: inst = 32'hc405119;
      12416: inst = 32'h8220000;
      12417: inst = 32'h10408000;
      12418: inst = 32'hc40511a;
      12419: inst = 32'h8220000;
      12420: inst = 32'h10408000;
      12421: inst = 32'hc40511b;
      12422: inst = 32'h8220000;
      12423: inst = 32'h10408000;
      12424: inst = 32'hc40511c;
      12425: inst = 32'h8220000;
      12426: inst = 32'h10408000;
      12427: inst = 32'hc40511d;
      12428: inst = 32'h8220000;
      12429: inst = 32'h10408000;
      12430: inst = 32'hc40511e;
      12431: inst = 32'h8220000;
      12432: inst = 32'h10408000;
      12433: inst = 32'hc405170;
      12434: inst = 32'h8220000;
      12435: inst = 32'h10408000;
      12436: inst = 32'hc405171;
      12437: inst = 32'h8220000;
      12438: inst = 32'h10408000;
      12439: inst = 32'hc405172;
      12440: inst = 32'h8220000;
      12441: inst = 32'h10408000;
      12442: inst = 32'hc405173;
      12443: inst = 32'h8220000;
      12444: inst = 32'h10408000;
      12445: inst = 32'hc405174;
      12446: inst = 32'h8220000;
      12447: inst = 32'h10408000;
      12448: inst = 32'hc405175;
      12449: inst = 32'h8220000;
      12450: inst = 32'h10408000;
      12451: inst = 32'hc405176;
      12452: inst = 32'h8220000;
      12453: inst = 32'h10408000;
      12454: inst = 32'hc405177;
      12455: inst = 32'h8220000;
      12456: inst = 32'h10408000;
      12457: inst = 32'hc405178;
      12458: inst = 32'h8220000;
      12459: inst = 32'h10408000;
      12460: inst = 32'hc405179;
      12461: inst = 32'h8220000;
      12462: inst = 32'h10408000;
      12463: inst = 32'hc40517a;
      12464: inst = 32'h8220000;
      12465: inst = 32'h10408000;
      12466: inst = 32'hc40517b;
      12467: inst = 32'h8220000;
      12468: inst = 32'h10408000;
      12469: inst = 32'hc40517c;
      12470: inst = 32'h8220000;
      12471: inst = 32'h10408000;
      12472: inst = 32'hc40517d;
      12473: inst = 32'h8220000;
      12474: inst = 32'h10408000;
      12475: inst = 32'hc40517e;
      12476: inst = 32'h8220000;
      12477: inst = 32'h10408000;
      12478: inst = 32'hc4051d0;
      12479: inst = 32'h8220000;
      12480: inst = 32'h10408000;
      12481: inst = 32'hc4051d1;
      12482: inst = 32'h8220000;
      12483: inst = 32'h10408000;
      12484: inst = 32'hc4051d2;
      12485: inst = 32'h8220000;
      12486: inst = 32'h10408000;
      12487: inst = 32'hc4051d3;
      12488: inst = 32'h8220000;
      12489: inst = 32'h10408000;
      12490: inst = 32'hc4051d4;
      12491: inst = 32'h8220000;
      12492: inst = 32'h10408000;
      12493: inst = 32'hc4051d5;
      12494: inst = 32'h8220000;
      12495: inst = 32'h10408000;
      12496: inst = 32'hc4051d6;
      12497: inst = 32'h8220000;
      12498: inst = 32'h10408000;
      12499: inst = 32'hc4051d7;
      12500: inst = 32'h8220000;
      12501: inst = 32'h10408000;
      12502: inst = 32'hc4051d8;
      12503: inst = 32'h8220000;
      12504: inst = 32'h10408000;
      12505: inst = 32'hc4051d9;
      12506: inst = 32'h8220000;
      12507: inst = 32'h10408000;
      12508: inst = 32'hc4051da;
      12509: inst = 32'h8220000;
      12510: inst = 32'h10408000;
      12511: inst = 32'hc4051db;
      12512: inst = 32'h8220000;
      12513: inst = 32'h10408000;
      12514: inst = 32'hc4051dc;
      12515: inst = 32'h8220000;
      12516: inst = 32'h10408000;
      12517: inst = 32'hc4051dd;
      12518: inst = 32'h8220000;
      12519: inst = 32'h10408000;
      12520: inst = 32'hc4051de;
      12521: inst = 32'h8220000;
      12522: inst = 32'h10408000;
      12523: inst = 32'hc405230;
      12524: inst = 32'h8220000;
      12525: inst = 32'h10408000;
      12526: inst = 32'hc405231;
      12527: inst = 32'h8220000;
      12528: inst = 32'h10408000;
      12529: inst = 32'hc405232;
      12530: inst = 32'h8220000;
      12531: inst = 32'h10408000;
      12532: inst = 32'hc405233;
      12533: inst = 32'h8220000;
      12534: inst = 32'h10408000;
      12535: inst = 32'hc405234;
      12536: inst = 32'h8220000;
      12537: inst = 32'h10408000;
      12538: inst = 32'hc405235;
      12539: inst = 32'h8220000;
      12540: inst = 32'h10408000;
      12541: inst = 32'hc405236;
      12542: inst = 32'h8220000;
      12543: inst = 32'h10408000;
      12544: inst = 32'hc405237;
      12545: inst = 32'h8220000;
      12546: inst = 32'h10408000;
      12547: inst = 32'hc405238;
      12548: inst = 32'h8220000;
      12549: inst = 32'h10408000;
      12550: inst = 32'hc405239;
      12551: inst = 32'h8220000;
      12552: inst = 32'h10408000;
      12553: inst = 32'hc40523a;
      12554: inst = 32'h8220000;
      12555: inst = 32'h10408000;
      12556: inst = 32'hc40523b;
      12557: inst = 32'h8220000;
      12558: inst = 32'h10408000;
      12559: inst = 32'hc40523c;
      12560: inst = 32'h8220000;
      12561: inst = 32'h10408000;
      12562: inst = 32'hc40523d;
      12563: inst = 32'h8220000;
      12564: inst = 32'h10408000;
      12565: inst = 32'hc40523e;
      12566: inst = 32'h8220000;
      12567: inst = 32'h10408000;
      12568: inst = 32'hc405290;
      12569: inst = 32'h8220000;
      12570: inst = 32'h10408000;
      12571: inst = 32'hc405291;
      12572: inst = 32'h8220000;
      12573: inst = 32'h10408000;
      12574: inst = 32'hc405292;
      12575: inst = 32'h8220000;
      12576: inst = 32'h10408000;
      12577: inst = 32'hc405293;
      12578: inst = 32'h8220000;
      12579: inst = 32'h10408000;
      12580: inst = 32'hc405294;
      12581: inst = 32'h8220000;
      12582: inst = 32'h10408000;
      12583: inst = 32'hc405295;
      12584: inst = 32'h8220000;
      12585: inst = 32'h10408000;
      12586: inst = 32'hc405296;
      12587: inst = 32'h8220000;
      12588: inst = 32'h10408000;
      12589: inst = 32'hc405297;
      12590: inst = 32'h8220000;
      12591: inst = 32'h10408000;
      12592: inst = 32'hc405298;
      12593: inst = 32'h8220000;
      12594: inst = 32'h10408000;
      12595: inst = 32'hc405299;
      12596: inst = 32'h8220000;
      12597: inst = 32'h10408000;
      12598: inst = 32'hc40529a;
      12599: inst = 32'h8220000;
      12600: inst = 32'h10408000;
      12601: inst = 32'hc40529b;
      12602: inst = 32'h8220000;
      12603: inst = 32'h10408000;
      12604: inst = 32'hc40529c;
      12605: inst = 32'h8220000;
      12606: inst = 32'h10408000;
      12607: inst = 32'hc40529d;
      12608: inst = 32'h8220000;
      12609: inst = 32'h10408000;
      12610: inst = 32'hc40529e;
      12611: inst = 32'h8220000;
      12612: inst = 32'hc20ef7c;
      12613: inst = 32'h10408000;
      12614: inst = 32'hc404932;
      12615: inst = 32'h8220000;
      12616: inst = 32'h10408000;
      12617: inst = 32'hc404933;
      12618: inst = 32'h8220000;
      12619: inst = 32'h10408000;
      12620: inst = 32'hc404934;
      12621: inst = 32'h8220000;
      12622: inst = 32'h10408000;
      12623: inst = 32'hc404935;
      12624: inst = 32'h8220000;
      12625: inst = 32'h10408000;
      12626: inst = 32'hc404993;
      12627: inst = 32'h8220000;
      12628: inst = 32'h10408000;
      12629: inst = 32'hc404994;
      12630: inst = 32'h8220000;
      12631: inst = 32'h10408000;
      12632: inst = 32'hc404995;
      12633: inst = 32'h8220000;
      12634: inst = 32'h10408000;
      12635: inst = 32'hc4049f3;
      12636: inst = 32'h8220000;
      12637: inst = 32'h10408000;
      12638: inst = 32'hc4049f4;
      12639: inst = 32'h8220000;
      12640: inst = 32'h10408000;
      12641: inst = 32'hc4049f5;
      12642: inst = 32'h8220000;
      12643: inst = 32'h10408000;
      12644: inst = 32'hc404a53;
      12645: inst = 32'h8220000;
      12646: inst = 32'h10408000;
      12647: inst = 32'hc404a54;
      12648: inst = 32'h8220000;
      12649: inst = 32'h10408000;
      12650: inst = 32'hc404a55;
      12651: inst = 32'h8220000;
      12652: inst = 32'h10408000;
      12653: inst = 32'hc404ab2;
      12654: inst = 32'h8220000;
      12655: inst = 32'h10408000;
      12656: inst = 32'hc404ab3;
      12657: inst = 32'h8220000;
      12658: inst = 32'h10408000;
      12659: inst = 32'hc404ab5;
      12660: inst = 32'h8220000;
      12661: inst = 32'h10408000;
      12662: inst = 32'hc404b12;
      12663: inst = 32'h8220000;
      12664: inst = 32'h10408000;
      12665: inst = 32'hc404b13;
      12666: inst = 32'h8220000;
      12667: inst = 32'h10408000;
      12668: inst = 32'hc404b15;
      12669: inst = 32'h8220000;
      12670: inst = 32'h10408000;
      12671: inst = 32'hc404b72;
      12672: inst = 32'h8220000;
      12673: inst = 32'h10408000;
      12674: inst = 32'hc404b73;
      12675: inst = 32'h8220000;
      12676: inst = 32'h10408000;
      12677: inst = 32'hc404b74;
      12678: inst = 32'h8220000;
      12679: inst = 32'h10408000;
      12680: inst = 32'hc404b75;
      12681: inst = 32'h8220000;
      12682: inst = 32'hc20eed7;
      12683: inst = 32'h10408000;
      12684: inst = 32'hc404a08;
      12685: inst = 32'h8220000;
      12686: inst = 32'h10408000;
      12687: inst = 32'hc404a0e;
      12688: inst = 32'h8220000;
      12689: inst = 32'hc20e6fa;
      12690: inst = 32'h10408000;
      12691: inst = 32'hc404a09;
      12692: inst = 32'h8220000;
      12693: inst = 32'h10408000;
      12694: inst = 32'hc404a0d;
      12695: inst = 32'h8220000;
      12696: inst = 32'h10408000;
      12697: inst = 32'hc404be7;
      12698: inst = 32'h8220000;
      12699: inst = 32'hc20e6fb;
      12700: inst = 32'h10408000;
      12701: inst = 32'hc404a0a;
      12702: inst = 32'h8220000;
      12703: inst = 32'h10408000;
      12704: inst = 32'hc404a0c;
      12705: inst = 32'h8220000;
      12706: inst = 32'h10408000;
      12707: inst = 32'hc404ac7;
      12708: inst = 32'h8220000;
      12709: inst = 32'h10408000;
      12710: inst = 32'hc404acf;
      12711: inst = 32'h8220000;
      12712: inst = 32'h10408000;
      12713: inst = 32'hc404b87;
      12714: inst = 32'h8220000;
      12715: inst = 32'h10408000;
      12716: inst = 32'hc404b8f;
      12717: inst = 32'h8220000;
      12718: inst = 32'h10408000;
      12719: inst = 32'hc404c4d;
      12720: inst = 32'h8220000;
      12721: inst = 32'hc20defb;
      12722: inst = 32'h10408000;
      12723: inst = 32'hc404a0b;
      12724: inst = 32'h8220000;
      12725: inst = 32'h10408000;
      12726: inst = 32'hc404a68;
      12727: inst = 32'h8220000;
      12728: inst = 32'h10408000;
      12729: inst = 32'hc404a69;
      12730: inst = 32'h8220000;
      12731: inst = 32'h10408000;
      12732: inst = 32'hc404a6a;
      12733: inst = 32'h8220000;
      12734: inst = 32'h10408000;
      12735: inst = 32'hc404a6b;
      12736: inst = 32'h8220000;
      12737: inst = 32'h10408000;
      12738: inst = 32'hc404a6c;
      12739: inst = 32'h8220000;
      12740: inst = 32'h10408000;
      12741: inst = 32'hc404a6d;
      12742: inst = 32'h8220000;
      12743: inst = 32'h10408000;
      12744: inst = 32'hc404a6e;
      12745: inst = 32'h8220000;
      12746: inst = 32'h10408000;
      12747: inst = 32'hc404ac8;
      12748: inst = 32'h8220000;
      12749: inst = 32'h10408000;
      12750: inst = 32'hc404ac9;
      12751: inst = 32'h8220000;
      12752: inst = 32'h10408000;
      12753: inst = 32'hc404aca;
      12754: inst = 32'h8220000;
      12755: inst = 32'h10408000;
      12756: inst = 32'hc404acb;
      12757: inst = 32'h8220000;
      12758: inst = 32'h10408000;
      12759: inst = 32'hc404acc;
      12760: inst = 32'h8220000;
      12761: inst = 32'h10408000;
      12762: inst = 32'hc404acd;
      12763: inst = 32'h8220000;
      12764: inst = 32'h10408000;
      12765: inst = 32'hc404ace;
      12766: inst = 32'h8220000;
      12767: inst = 32'h10408000;
      12768: inst = 32'hc404b27;
      12769: inst = 32'h8220000;
      12770: inst = 32'h10408000;
      12771: inst = 32'hc404b2a;
      12772: inst = 32'h8220000;
      12773: inst = 32'h10408000;
      12774: inst = 32'hc404b2d;
      12775: inst = 32'h8220000;
      12776: inst = 32'h10408000;
      12777: inst = 32'hc404b2e;
      12778: inst = 32'h8220000;
      12779: inst = 32'h10408000;
      12780: inst = 32'hc404b2f;
      12781: inst = 32'h8220000;
      12782: inst = 32'h10408000;
      12783: inst = 32'hc404b8a;
      12784: inst = 32'h8220000;
      12785: inst = 32'h10408000;
      12786: inst = 32'hc404b8d;
      12787: inst = 32'h8220000;
      12788: inst = 32'h10408000;
      12789: inst = 32'hc404b8e;
      12790: inst = 32'h8220000;
      12791: inst = 32'h10408000;
      12792: inst = 32'hc404be8;
      12793: inst = 32'h8220000;
      12794: inst = 32'h10408000;
      12795: inst = 32'hc404be9;
      12796: inst = 32'h8220000;
      12797: inst = 32'h10408000;
      12798: inst = 32'hc404bea;
      12799: inst = 32'h8220000;
      12800: inst = 32'h10408000;
      12801: inst = 32'hc404beb;
      12802: inst = 32'h8220000;
      12803: inst = 32'h10408000;
      12804: inst = 32'hc404bec;
      12805: inst = 32'h8220000;
      12806: inst = 32'h10408000;
      12807: inst = 32'hc404bed;
      12808: inst = 32'h8220000;
      12809: inst = 32'h10408000;
      12810: inst = 32'hc404bee;
      12811: inst = 32'h8220000;
      12812: inst = 32'h10408000;
      12813: inst = 32'hc404c49;
      12814: inst = 32'h8220000;
      12815: inst = 32'h10408000;
      12816: inst = 32'hc404c4b;
      12817: inst = 32'h8220000;
      12818: inst = 32'h10408000;
      12819: inst = 32'hc404ca9;
      12820: inst = 32'h8220000;
      12821: inst = 32'h10408000;
      12822: inst = 32'hc404cab;
      12823: inst = 32'h8220000;
      12824: inst = 32'hc20eed8;
      12825: inst = 32'h10408000;
      12826: inst = 32'hc404a67;
      12827: inst = 32'h8220000;
      12828: inst = 32'h10408000;
      12829: inst = 32'hc404a6f;
      12830: inst = 32'h8220000;
      12831: inst = 32'hc204a69;
      12832: inst = 32'h10408000;
      12833: inst = 32'hc404b28;
      12834: inst = 32'h8220000;
      12835: inst = 32'h10408000;
      12836: inst = 32'hc404b29;
      12837: inst = 32'h8220000;
      12838: inst = 32'h10408000;
      12839: inst = 32'hc404b2b;
      12840: inst = 32'h8220000;
      12841: inst = 32'h10408000;
      12842: inst = 32'hc404b2c;
      12843: inst = 32'h8220000;
      12844: inst = 32'h10408000;
      12845: inst = 32'hc404b88;
      12846: inst = 32'h8220000;
      12847: inst = 32'h10408000;
      12848: inst = 32'hc404b89;
      12849: inst = 32'h8220000;
      12850: inst = 32'h10408000;
      12851: inst = 32'hc404b8b;
      12852: inst = 32'h8220000;
      12853: inst = 32'h10408000;
      12854: inst = 32'hc404b8c;
      12855: inst = 32'h8220000;
      12856: inst = 32'h10408000;
      12857: inst = 32'hc404c48;
      12858: inst = 32'h8220000;
      12859: inst = 32'h10408000;
      12860: inst = 32'hc404c4a;
      12861: inst = 32'h8220000;
      12862: inst = 32'h10408000;
      12863: inst = 32'hc404c4c;
      12864: inst = 32'h8220000;
      12865: inst = 32'h10408000;
      12866: inst = 32'hc404ca8;
      12867: inst = 32'h8220000;
      12868: inst = 32'h10408000;
      12869: inst = 32'hc404caa;
      12870: inst = 32'h8220000;
      12871: inst = 32'h10408000;
      12872: inst = 32'hc404cac;
      12873: inst = 32'h8220000;
      12874: inst = 32'h10408000;
      12875: inst = 32'hc405085;
      12876: inst = 32'h8220000;
      12877: inst = 32'h10408000;
      12878: inst = 32'hc40509a;
      12879: inst = 32'h8220000;
      12880: inst = 32'h10408000;
      12881: inst = 32'hc4050e4;
      12882: inst = 32'h8220000;
      12883: inst = 32'h10408000;
      12884: inst = 32'hc4050e5;
      12885: inst = 32'h8220000;
      12886: inst = 32'h10408000;
      12887: inst = 32'hc4050fa;
      12888: inst = 32'h8220000;
      12889: inst = 32'h10408000;
      12890: inst = 32'hc4050fb;
      12891: inst = 32'h8220000;
      12892: inst = 32'h10408000;
      12893: inst = 32'hc405143;
      12894: inst = 32'h8220000;
      12895: inst = 32'h10408000;
      12896: inst = 32'hc405144;
      12897: inst = 32'h8220000;
      12898: inst = 32'h10408000;
      12899: inst = 32'hc405145;
      12900: inst = 32'h8220000;
      12901: inst = 32'h10408000;
      12902: inst = 32'hc40515a;
      12903: inst = 32'h8220000;
      12904: inst = 32'h10408000;
      12905: inst = 32'hc40515b;
      12906: inst = 32'h8220000;
      12907: inst = 32'h10408000;
      12908: inst = 32'hc40515c;
      12909: inst = 32'h8220000;
      12910: inst = 32'h10408000;
      12911: inst = 32'hc4051a2;
      12912: inst = 32'h8220000;
      12913: inst = 32'h10408000;
      12914: inst = 32'hc4051a3;
      12915: inst = 32'h8220000;
      12916: inst = 32'h10408000;
      12917: inst = 32'hc4051a4;
      12918: inst = 32'h8220000;
      12919: inst = 32'h10408000;
      12920: inst = 32'hc4051a5;
      12921: inst = 32'h8220000;
      12922: inst = 32'h10408000;
      12923: inst = 32'hc4051ba;
      12924: inst = 32'h8220000;
      12925: inst = 32'h10408000;
      12926: inst = 32'hc4051bb;
      12927: inst = 32'h8220000;
      12928: inst = 32'h10408000;
      12929: inst = 32'hc4051bc;
      12930: inst = 32'h8220000;
      12931: inst = 32'h10408000;
      12932: inst = 32'hc4051bd;
      12933: inst = 32'h8220000;
      12934: inst = 32'h10408000;
      12935: inst = 32'hc405202;
      12936: inst = 32'h8220000;
      12937: inst = 32'h10408000;
      12938: inst = 32'hc405203;
      12939: inst = 32'h8220000;
      12940: inst = 32'h10408000;
      12941: inst = 32'hc405204;
      12942: inst = 32'h8220000;
      12943: inst = 32'h10408000;
      12944: inst = 32'hc405205;
      12945: inst = 32'h8220000;
      12946: inst = 32'h10408000;
      12947: inst = 32'hc40521a;
      12948: inst = 32'h8220000;
      12949: inst = 32'h10408000;
      12950: inst = 32'hc40521b;
      12951: inst = 32'h8220000;
      12952: inst = 32'h10408000;
      12953: inst = 32'hc40521c;
      12954: inst = 32'h8220000;
      12955: inst = 32'h10408000;
      12956: inst = 32'hc40521d;
      12957: inst = 32'h8220000;
      12958: inst = 32'h10408000;
      12959: inst = 32'hc405262;
      12960: inst = 32'h8220000;
      12961: inst = 32'h10408000;
      12962: inst = 32'hc405263;
      12963: inst = 32'h8220000;
      12964: inst = 32'h10408000;
      12965: inst = 32'hc405264;
      12966: inst = 32'h8220000;
      12967: inst = 32'h10408000;
      12968: inst = 32'hc405265;
      12969: inst = 32'h8220000;
      12970: inst = 32'h10408000;
      12971: inst = 32'hc40527a;
      12972: inst = 32'h8220000;
      12973: inst = 32'h10408000;
      12974: inst = 32'hc40527b;
      12975: inst = 32'h8220000;
      12976: inst = 32'h10408000;
      12977: inst = 32'hc40527c;
      12978: inst = 32'h8220000;
      12979: inst = 32'h10408000;
      12980: inst = 32'hc40527d;
      12981: inst = 32'h8220000;
      12982: inst = 32'h10408000;
      12983: inst = 32'hc4052c2;
      12984: inst = 32'h8220000;
      12985: inst = 32'h10408000;
      12986: inst = 32'hc4052c3;
      12987: inst = 32'h8220000;
      12988: inst = 32'h10408000;
      12989: inst = 32'hc4052c4;
      12990: inst = 32'h8220000;
      12991: inst = 32'h10408000;
      12992: inst = 32'hc4052db;
      12993: inst = 32'h8220000;
      12994: inst = 32'h10408000;
      12995: inst = 32'hc4052dc;
      12996: inst = 32'h8220000;
      12997: inst = 32'h10408000;
      12998: inst = 32'hc4052dd;
      12999: inst = 32'h8220000;
      13000: inst = 32'h10408000;
      13001: inst = 32'hc405322;
      13002: inst = 32'h8220000;
      13003: inst = 32'h10408000;
      13004: inst = 32'hc405323;
      13005: inst = 32'h8220000;
      13006: inst = 32'h10408000;
      13007: inst = 32'hc405324;
      13008: inst = 32'h8220000;
      13009: inst = 32'h10408000;
      13010: inst = 32'hc40533b;
      13011: inst = 32'h8220000;
      13012: inst = 32'h10408000;
      13013: inst = 32'hc40533c;
      13014: inst = 32'h8220000;
      13015: inst = 32'h10408000;
      13016: inst = 32'hc40533d;
      13017: inst = 32'h8220000;
      13018: inst = 32'h10408000;
      13019: inst = 32'hc40537f;
      13020: inst = 32'h8220000;
      13021: inst = 32'h10408000;
      13022: inst = 32'hc405382;
      13023: inst = 32'h8220000;
      13024: inst = 32'h10408000;
      13025: inst = 32'hc405383;
      13026: inst = 32'h8220000;
      13027: inst = 32'h10408000;
      13028: inst = 32'hc405384;
      13029: inst = 32'h8220000;
      13030: inst = 32'h10408000;
      13031: inst = 32'hc40539b;
      13032: inst = 32'h8220000;
      13033: inst = 32'h10408000;
      13034: inst = 32'hc40539c;
      13035: inst = 32'h8220000;
      13036: inst = 32'h10408000;
      13037: inst = 32'hc40539d;
      13038: inst = 32'h8220000;
      13039: inst = 32'h10408000;
      13040: inst = 32'hc4053a0;
      13041: inst = 32'h8220000;
      13042: inst = 32'h10408000;
      13043: inst = 32'hc4053de;
      13044: inst = 32'h8220000;
      13045: inst = 32'h10408000;
      13046: inst = 32'hc4053df;
      13047: inst = 32'h8220000;
      13048: inst = 32'h10408000;
      13049: inst = 32'hc4053e2;
      13050: inst = 32'h8220000;
      13051: inst = 32'h10408000;
      13052: inst = 32'hc4053e3;
      13053: inst = 32'h8220000;
      13054: inst = 32'h10408000;
      13055: inst = 32'hc4053fc;
      13056: inst = 32'h8220000;
      13057: inst = 32'h10408000;
      13058: inst = 32'hc4053fd;
      13059: inst = 32'h8220000;
      13060: inst = 32'h10408000;
      13061: inst = 32'hc405400;
      13062: inst = 32'h8220000;
      13063: inst = 32'h10408000;
      13064: inst = 32'hc405401;
      13065: inst = 32'h8220000;
      13066: inst = 32'h10408000;
      13067: inst = 32'hc40543d;
      13068: inst = 32'h8220000;
      13069: inst = 32'h10408000;
      13070: inst = 32'hc40543e;
      13071: inst = 32'h8220000;
      13072: inst = 32'h10408000;
      13073: inst = 32'hc40543f;
      13074: inst = 32'h8220000;
      13075: inst = 32'h10408000;
      13076: inst = 32'hc405442;
      13077: inst = 32'h8220000;
      13078: inst = 32'h10408000;
      13079: inst = 32'hc405443;
      13080: inst = 32'h8220000;
      13081: inst = 32'h10408000;
      13082: inst = 32'hc40545c;
      13083: inst = 32'h8220000;
      13084: inst = 32'h10408000;
      13085: inst = 32'hc40545d;
      13086: inst = 32'h8220000;
      13087: inst = 32'h10408000;
      13088: inst = 32'hc405460;
      13089: inst = 32'h8220000;
      13090: inst = 32'h10408000;
      13091: inst = 32'hc405461;
      13092: inst = 32'h8220000;
      13093: inst = 32'h10408000;
      13094: inst = 32'hc405462;
      13095: inst = 32'h8220000;
      13096: inst = 32'h10408000;
      13097: inst = 32'hc40549d;
      13098: inst = 32'h8220000;
      13099: inst = 32'h10408000;
      13100: inst = 32'hc40549e;
      13101: inst = 32'h8220000;
      13102: inst = 32'h10408000;
      13103: inst = 32'hc4054a0;
      13104: inst = 32'h8220000;
      13105: inst = 32'h10408000;
      13106: inst = 32'hc4054a1;
      13107: inst = 32'h8220000;
      13108: inst = 32'h10408000;
      13109: inst = 32'hc4054a2;
      13110: inst = 32'h8220000;
      13111: inst = 32'h10408000;
      13112: inst = 32'hc4054a3;
      13113: inst = 32'h8220000;
      13114: inst = 32'h10408000;
      13115: inst = 32'hc4054bc;
      13116: inst = 32'h8220000;
      13117: inst = 32'h10408000;
      13118: inst = 32'hc4054bd;
      13119: inst = 32'h8220000;
      13120: inst = 32'h10408000;
      13121: inst = 32'hc4054be;
      13122: inst = 32'h8220000;
      13123: inst = 32'h10408000;
      13124: inst = 32'hc4054bf;
      13125: inst = 32'h8220000;
      13126: inst = 32'h10408000;
      13127: inst = 32'hc4054c1;
      13128: inst = 32'h8220000;
      13129: inst = 32'h10408000;
      13130: inst = 32'hc4054c2;
      13131: inst = 32'h8220000;
      13132: inst = 32'h10408000;
      13133: inst = 32'hc4054fc;
      13134: inst = 32'h8220000;
      13135: inst = 32'h10408000;
      13136: inst = 32'hc4054fd;
      13137: inst = 32'h8220000;
      13138: inst = 32'h10408000;
      13139: inst = 32'hc4054fe;
      13140: inst = 32'h8220000;
      13141: inst = 32'h10408000;
      13142: inst = 32'hc405502;
      13143: inst = 32'h8220000;
      13144: inst = 32'h10408000;
      13145: inst = 32'hc40551d;
      13146: inst = 32'h8220000;
      13147: inst = 32'h10408000;
      13148: inst = 32'hc405521;
      13149: inst = 32'h8220000;
      13150: inst = 32'h10408000;
      13151: inst = 32'hc405522;
      13152: inst = 32'h8220000;
      13153: inst = 32'h10408000;
      13154: inst = 32'hc405523;
      13155: inst = 32'h8220000;
      13156: inst = 32'h10408000;
      13157: inst = 32'hc40555b;
      13158: inst = 32'h8220000;
      13159: inst = 32'h10408000;
      13160: inst = 32'hc40555c;
      13161: inst = 32'h8220000;
      13162: inst = 32'h10408000;
      13163: inst = 32'hc40555d;
      13164: inst = 32'h8220000;
      13165: inst = 32'h10408000;
      13166: inst = 32'hc405562;
      13167: inst = 32'h8220000;
      13168: inst = 32'h10408000;
      13169: inst = 32'hc40557d;
      13170: inst = 32'h8220000;
      13171: inst = 32'h10408000;
      13172: inst = 32'hc405582;
      13173: inst = 32'h8220000;
      13174: inst = 32'h10408000;
      13175: inst = 32'hc405583;
      13176: inst = 32'h8220000;
      13177: inst = 32'h10408000;
      13178: inst = 32'hc405584;
      13179: inst = 32'h8220000;
      13180: inst = 32'h10408000;
      13181: inst = 32'hc4055ba;
      13182: inst = 32'h8220000;
      13183: inst = 32'h10408000;
      13184: inst = 32'hc4055bb;
      13185: inst = 32'h8220000;
      13186: inst = 32'h10408000;
      13187: inst = 32'hc4055bc;
      13188: inst = 32'h8220000;
      13189: inst = 32'h10408000;
      13190: inst = 32'hc4055bd;
      13191: inst = 32'h8220000;
      13192: inst = 32'h10408000;
      13193: inst = 32'hc4055c2;
      13194: inst = 32'h8220000;
      13195: inst = 32'h10408000;
      13196: inst = 32'hc4055dd;
      13197: inst = 32'h8220000;
      13198: inst = 32'h10408000;
      13199: inst = 32'hc4055e2;
      13200: inst = 32'h8220000;
      13201: inst = 32'h10408000;
      13202: inst = 32'hc4055e3;
      13203: inst = 32'h8220000;
      13204: inst = 32'h10408000;
      13205: inst = 32'hc4055e4;
      13206: inst = 32'h8220000;
      13207: inst = 32'h10408000;
      13208: inst = 32'hc4055e5;
      13209: inst = 32'h8220000;
      13210: inst = 32'h10408000;
      13211: inst = 32'hc40561a;
      13212: inst = 32'h8220000;
      13213: inst = 32'h10408000;
      13214: inst = 32'hc40561b;
      13215: inst = 32'h8220000;
      13216: inst = 32'h10408000;
      13217: inst = 32'hc40561c;
      13218: inst = 32'h8220000;
      13219: inst = 32'h10408000;
      13220: inst = 32'hc40561d;
      13221: inst = 32'h8220000;
      13222: inst = 32'h10408000;
      13223: inst = 32'hc405642;
      13224: inst = 32'h8220000;
      13225: inst = 32'h10408000;
      13226: inst = 32'hc405643;
      13227: inst = 32'h8220000;
      13228: inst = 32'h10408000;
      13229: inst = 32'hc405644;
      13230: inst = 32'h8220000;
      13231: inst = 32'h10408000;
      13232: inst = 32'hc405645;
      13233: inst = 32'h8220000;
      13234: inst = 32'h10408000;
      13235: inst = 32'hc405679;
      13236: inst = 32'h8220000;
      13237: inst = 32'h10408000;
      13238: inst = 32'hc40567a;
      13239: inst = 32'h8220000;
      13240: inst = 32'h10408000;
      13241: inst = 32'hc40567b;
      13242: inst = 32'h8220000;
      13243: inst = 32'h10408000;
      13244: inst = 32'hc40567c;
      13245: inst = 32'h8220000;
      13246: inst = 32'h10408000;
      13247: inst = 32'hc4056a3;
      13248: inst = 32'h8220000;
      13249: inst = 32'h10408000;
      13250: inst = 32'hc4056a4;
      13251: inst = 32'h8220000;
      13252: inst = 32'h10408000;
      13253: inst = 32'hc4056a5;
      13254: inst = 32'h8220000;
      13255: inst = 32'h10408000;
      13256: inst = 32'hc4056a6;
      13257: inst = 32'h8220000;
      13258: inst = 32'hc20e6d9;
      13259: inst = 32'h10408000;
      13260: inst = 32'hc404bef;
      13261: inst = 32'h8220000;
      13262: inst = 32'h10408000;
      13263: inst = 32'hc404c4e;
      13264: inst = 32'h8220000;
      13265: inst = 32'hc20eeb7;
      13266: inst = 32'h10408000;
      13267: inst = 32'hc404c47;
      13268: inst = 32'h8220000;
      13269: inst = 32'hc20d615;
      13270: inst = 32'h10408000;
      13271: inst = 32'hc404ca2;
      13272: inst = 32'h8220000;
      13273: inst = 32'h10408000;
      13274: inst = 32'hc404d00;
      13275: inst = 32'h8220000;
      13276: inst = 32'hc209c91;
      13277: inst = 32'h10408000;
      13278: inst = 32'hc404ca3;
      13279: inst = 32'h8220000;
      13280: inst = 32'h10408000;
      13281: inst = 32'hc404d01;
      13282: inst = 32'h8220000;
      13283: inst = 32'hc207bf0;
      13284: inst = 32'h10408000;
      13285: inst = 32'hc404ca4;
      13286: inst = 32'h8220000;
      13287: inst = 32'h10408000;
      13288: inst = 32'hc404ca5;
      13289: inst = 32'h8220000;
      13290: inst = 32'h10408000;
      13291: inst = 32'hc404ca6;
      13292: inst = 32'h8220000;
      13293: inst = 32'h10408000;
      13294: inst = 32'hc404ca7;
      13295: inst = 32'h8220000;
      13296: inst = 32'h10408000;
      13297: inst = 32'hc404d02;
      13298: inst = 32'h8220000;
      13299: inst = 32'h10408000;
      13300: inst = 32'hc404d03;
      13301: inst = 32'h8220000;
      13302: inst = 32'h10408000;
      13303: inst = 32'hc404d04;
      13304: inst = 32'h8220000;
      13305: inst = 32'h10408000;
      13306: inst = 32'hc404d05;
      13307: inst = 32'h8220000;
      13308: inst = 32'h10408000;
      13309: inst = 32'hc404d06;
      13310: inst = 32'h8220000;
      13311: inst = 32'h10408000;
      13312: inst = 32'hc404d07;
      13313: inst = 32'h8220000;
      13314: inst = 32'h10408000;
      13315: inst = 32'hc404d08;
      13316: inst = 32'h8220000;
      13317: inst = 32'h10408000;
      13318: inst = 32'hc404d09;
      13319: inst = 32'h8220000;
      13320: inst = 32'h10408000;
      13321: inst = 32'hc404d0a;
      13322: inst = 32'h8220000;
      13323: inst = 32'h10408000;
      13324: inst = 32'hc404d0b;
      13325: inst = 32'h8220000;
      13326: inst = 32'h10408000;
      13327: inst = 32'hc404d0c;
      13328: inst = 32'h8220000;
      13329: inst = 32'h10408000;
      13330: inst = 32'hc404d0d;
      13331: inst = 32'h8220000;
      13332: inst = 32'h10408000;
      13333: inst = 32'hc404d0e;
      13334: inst = 32'h8220000;
      13335: inst = 32'h10408000;
      13336: inst = 32'hc404d0f;
      13337: inst = 32'h8220000;
      13338: inst = 32'h10408000;
      13339: inst = 32'hc404d10;
      13340: inst = 32'h8220000;
      13341: inst = 32'h10408000;
      13342: inst = 32'hc404d11;
      13343: inst = 32'h8220000;
      13344: inst = 32'h10408000;
      13345: inst = 32'hc404d12;
      13346: inst = 32'h8220000;
      13347: inst = 32'h10408000;
      13348: inst = 32'hc404d13;
      13349: inst = 32'h8220000;
      13350: inst = 32'h10408000;
      13351: inst = 32'hc404d14;
      13352: inst = 32'h8220000;
      13353: inst = 32'h10408000;
      13354: inst = 32'hc4055c3;
      13355: inst = 32'h8220000;
      13356: inst = 32'h10408000;
      13357: inst = 32'hc4055dc;
      13358: inst = 32'h8220000;
      13359: inst = 32'hc20ad55;
      13360: inst = 32'h10408000;
      13361: inst = 32'hc404cad;
      13362: inst = 32'h8220000;
      13363: inst = 32'hc208410;
      13364: inst = 32'h10408000;
      13365: inst = 32'hc404cae;
      13366: inst = 32'h8220000;
      13367: inst = 32'h10408000;
      13368: inst = 32'hc404caf;
      13369: inst = 32'h8220000;
      13370: inst = 32'h10408000;
      13371: inst = 32'hc404cb0;
      13372: inst = 32'h8220000;
      13373: inst = 32'h10408000;
      13374: inst = 32'hc404cb1;
      13375: inst = 32'h8220000;
      13376: inst = 32'h10408000;
      13377: inst = 32'hc404cb2;
      13378: inst = 32'h8220000;
      13379: inst = 32'h10408000;
      13380: inst = 32'hc404cb3;
      13381: inst = 32'h8220000;
      13382: inst = 32'h10408000;
      13383: inst = 32'hc404cb4;
      13384: inst = 32'h8220000;
      13385: inst = 32'h10408000;
      13386: inst = 32'hc404cb5;
      13387: inst = 32'h8220000;
      13388: inst = 32'h10408000;
      13389: inst = 32'hc40537d;
      13390: inst = 32'h8220000;
      13391: inst = 32'h10408000;
      13392: inst = 32'hc405385;
      13393: inst = 32'h8220000;
      13394: inst = 32'h10408000;
      13395: inst = 32'hc40539a;
      13396: inst = 32'h8220000;
      13397: inst = 32'h10408000;
      13398: inst = 32'hc4053a2;
      13399: inst = 32'h8220000;
      13400: inst = 32'h10408000;
      13401: inst = 32'hc4054a4;
      13402: inst = 32'h8220000;
      13403: inst = 32'h10408000;
      13404: inst = 32'hc4054bb;
      13405: inst = 32'h8220000;
      13406: inst = 32'h10408000;
      13407: inst = 32'hc405741;
      13408: inst = 32'h8220000;
      13409: inst = 32'h10408000;
      13410: inst = 32'hc40575e;
      13411: inst = 32'h8220000;
      13412: inst = 32'hc209470;
      13413: inst = 32'h10408000;
      13414: inst = 32'hc404cb6;
      13415: inst = 32'h8220000;
      13416: inst = 32'h10408000;
      13417: inst = 32'hc404d15;
      13418: inst = 32'h8220000;
      13419: inst = 32'hc20a534;
      13420: inst = 32'h10408000;
      13421: inst = 32'hc404cfb;
      13422: inst = 32'h8220000;
      13423: inst = 32'hc208c51;
      13424: inst = 32'h10408000;
      13425: inst = 32'hc404cfc;
      13426: inst = 32'h8220000;
      13427: inst = 32'h10408000;
      13428: inst = 32'hc404cfd;
      13429: inst = 32'h8220000;
      13430: inst = 32'h10408000;
      13431: inst = 32'hc4053da;
      13432: inst = 32'h8220000;
      13433: inst = 32'h10408000;
      13434: inst = 32'hc4053dc;
      13435: inst = 32'h8220000;
      13436: inst = 32'h10408000;
      13437: inst = 32'hc405403;
      13438: inst = 32'h8220000;
      13439: inst = 32'h10408000;
      13440: inst = 32'hc405405;
      13441: inst = 32'h8220000;
      13442: inst = 32'h10408000;
      13443: inst = 32'hc4054fa;
      13444: inst = 32'h8220000;
      13445: inst = 32'h10408000;
      13446: inst = 32'hc405525;
      13447: inst = 32'h8220000;
      13448: inst = 32'h10408000;
      13449: inst = 32'hc405557;
      13450: inst = 32'h8220000;
      13451: inst = 32'h10408000;
      13452: inst = 32'hc40555f;
      13453: inst = 32'h8220000;
      13454: inst = 32'h10408000;
      13455: inst = 32'hc405580;
      13456: inst = 32'h8220000;
      13457: inst = 32'h10408000;
      13458: inst = 32'hc405588;
      13459: inst = 32'h8220000;
      13460: inst = 32'h10408000;
      13461: inst = 32'hc405618;
      13462: inst = 32'h8220000;
      13463: inst = 32'h10408000;
      13464: inst = 32'hc405627;
      13465: inst = 32'h8220000;
      13466: inst = 32'h10408000;
      13467: inst = 32'hc405638;
      13468: inst = 32'h8220000;
      13469: inst = 32'h10408000;
      13470: inst = 32'hc405647;
      13471: inst = 32'h8220000;
      13472: inst = 32'h10408000;
      13473: inst = 32'hc40570b;
      13474: inst = 32'h8220000;
      13475: inst = 32'hc206b6d;
      13476: inst = 32'h10408000;
      13477: inst = 32'hc404d16;
      13478: inst = 32'h8220000;
      13479: inst = 32'h10408000;
      13480: inst = 32'hc404d75;
      13481: inst = 32'h8220000;
      13482: inst = 32'h10408000;
      13483: inst = 32'hc404d76;
      13484: inst = 32'h8220000;
      13485: inst = 32'h10408000;
      13486: inst = 32'hc404dd5;
      13487: inst = 32'h8220000;
      13488: inst = 32'h10408000;
      13489: inst = 32'hc404dd6;
      13490: inst = 32'h8220000;
      13491: inst = 32'h10408000;
      13492: inst = 32'hc404e35;
      13493: inst = 32'h8220000;
      13494: inst = 32'h10408000;
      13495: inst = 32'hc404e36;
      13496: inst = 32'h8220000;
      13497: inst = 32'h10408000;
      13498: inst = 32'hc404e95;
      13499: inst = 32'h8220000;
      13500: inst = 32'h10408000;
      13501: inst = 32'hc404e96;
      13502: inst = 32'h8220000;
      13503: inst = 32'h10408000;
      13504: inst = 32'hc404ef5;
      13505: inst = 32'h8220000;
      13506: inst = 32'h10408000;
      13507: inst = 32'hc404ef6;
      13508: inst = 32'h8220000;
      13509: inst = 32'h10408000;
      13510: inst = 32'hc404f55;
      13511: inst = 32'h8220000;
      13512: inst = 32'h10408000;
      13513: inst = 32'hc404f56;
      13514: inst = 32'h8220000;
      13515: inst = 32'h10408000;
      13516: inst = 32'hc404fb5;
      13517: inst = 32'h8220000;
      13518: inst = 32'h10408000;
      13519: inst = 32'hc404fb6;
      13520: inst = 32'h8220000;
      13521: inst = 32'h10408000;
      13522: inst = 32'hc405015;
      13523: inst = 32'h8220000;
      13524: inst = 32'h10408000;
      13525: inst = 32'hc405016;
      13526: inst = 32'h8220000;
      13527: inst = 32'h10408000;
      13528: inst = 32'hc405075;
      13529: inst = 32'h8220000;
      13530: inst = 32'h10408000;
      13531: inst = 32'hc405076;
      13532: inst = 32'h8220000;
      13533: inst = 32'h10408000;
      13534: inst = 32'hc4050d5;
      13535: inst = 32'h8220000;
      13536: inst = 32'h10408000;
      13537: inst = 32'hc4050d6;
      13538: inst = 32'h8220000;
      13539: inst = 32'h10408000;
      13540: inst = 32'hc405135;
      13541: inst = 32'h8220000;
      13542: inst = 32'h10408000;
      13543: inst = 32'hc405136;
      13544: inst = 32'h8220000;
      13545: inst = 32'h10408000;
      13546: inst = 32'hc405195;
      13547: inst = 32'h8220000;
      13548: inst = 32'h10408000;
      13549: inst = 32'hc405196;
      13550: inst = 32'h8220000;
      13551: inst = 32'h10408000;
      13552: inst = 32'hc4051f5;
      13553: inst = 32'h8220000;
      13554: inst = 32'h10408000;
      13555: inst = 32'hc4051f6;
      13556: inst = 32'h8220000;
      13557: inst = 32'h10408000;
      13558: inst = 32'hc405255;
      13559: inst = 32'h8220000;
      13560: inst = 32'h10408000;
      13561: inst = 32'hc405256;
      13562: inst = 32'h8220000;
      13563: inst = 32'h10408000;
      13564: inst = 32'hc4052b5;
      13565: inst = 32'h8220000;
      13566: inst = 32'h10408000;
      13567: inst = 32'hc4052b6;
      13568: inst = 32'h8220000;
      13569: inst = 32'h10408000;
      13570: inst = 32'hc405325;
      13571: inst = 32'h8220000;
      13572: inst = 32'h10408000;
      13573: inst = 32'hc40533a;
      13574: inst = 32'h8220000;
      13575: inst = 32'hc20c638;
      13576: inst = 32'h10408000;
      13577: inst = 32'hc404d5b;
      13578: inst = 32'h8220000;
      13579: inst = 32'hc208c71;
      13580: inst = 32'h10408000;
      13581: inst = 32'hc404d60;
      13582: inst = 32'h8220000;
      13583: inst = 32'h10408000;
      13584: inst = 32'hc404d61;
      13585: inst = 32'h8220000;
      13586: inst = 32'h10408000;
      13587: inst = 32'hc404d62;
      13588: inst = 32'h8220000;
      13589: inst = 32'h10408000;
      13590: inst = 32'hc404d63;
      13591: inst = 32'h8220000;
      13592: inst = 32'h10408000;
      13593: inst = 32'hc404d64;
      13594: inst = 32'h8220000;
      13595: inst = 32'h10408000;
      13596: inst = 32'hc404d65;
      13597: inst = 32'h8220000;
      13598: inst = 32'h10408000;
      13599: inst = 32'hc404d66;
      13600: inst = 32'h8220000;
      13601: inst = 32'h10408000;
      13602: inst = 32'hc404d67;
      13603: inst = 32'h8220000;
      13604: inst = 32'h10408000;
      13605: inst = 32'hc404d68;
      13606: inst = 32'h8220000;
      13607: inst = 32'h10408000;
      13608: inst = 32'hc404d69;
      13609: inst = 32'h8220000;
      13610: inst = 32'h10408000;
      13611: inst = 32'hc404d6a;
      13612: inst = 32'h8220000;
      13613: inst = 32'h10408000;
      13614: inst = 32'hc404d6b;
      13615: inst = 32'h8220000;
      13616: inst = 32'h10408000;
      13617: inst = 32'hc404d6c;
      13618: inst = 32'h8220000;
      13619: inst = 32'h10408000;
      13620: inst = 32'hc404d6d;
      13621: inst = 32'h8220000;
      13622: inst = 32'h10408000;
      13623: inst = 32'hc404d6e;
      13624: inst = 32'h8220000;
      13625: inst = 32'h10408000;
      13626: inst = 32'hc404d6f;
      13627: inst = 32'h8220000;
      13628: inst = 32'h10408000;
      13629: inst = 32'hc404d70;
      13630: inst = 32'h8220000;
      13631: inst = 32'h10408000;
      13632: inst = 32'hc404d71;
      13633: inst = 32'h8220000;
      13634: inst = 32'h10408000;
      13635: inst = 32'hc404d72;
      13636: inst = 32'h8220000;
      13637: inst = 32'h10408000;
      13638: inst = 32'hc404d73;
      13639: inst = 32'h8220000;
      13640: inst = 32'h10408000;
      13641: inst = 32'hc404d74;
      13642: inst = 32'h8220000;
      13643: inst = 32'h10408000;
      13644: inst = 32'hc404dc0;
      13645: inst = 32'h8220000;
      13646: inst = 32'h10408000;
      13647: inst = 32'hc404dca;
      13648: inst = 32'h8220000;
      13649: inst = 32'h10408000;
      13650: inst = 32'hc404dd4;
      13651: inst = 32'h8220000;
      13652: inst = 32'h10408000;
      13653: inst = 32'hc404e20;
      13654: inst = 32'h8220000;
      13655: inst = 32'h10408000;
      13656: inst = 32'hc404e2a;
      13657: inst = 32'h8220000;
      13658: inst = 32'h10408000;
      13659: inst = 32'hc404e34;
      13660: inst = 32'h8220000;
      13661: inst = 32'h10408000;
      13662: inst = 32'hc404e80;
      13663: inst = 32'h8220000;
      13664: inst = 32'h10408000;
      13665: inst = 32'hc404e8a;
      13666: inst = 32'h8220000;
      13667: inst = 32'h10408000;
      13668: inst = 32'hc404e94;
      13669: inst = 32'h8220000;
      13670: inst = 32'h10408000;
      13671: inst = 32'hc404ee0;
      13672: inst = 32'h8220000;
      13673: inst = 32'h10408000;
      13674: inst = 32'hc404eea;
      13675: inst = 32'h8220000;
      13676: inst = 32'h10408000;
      13677: inst = 32'hc404ef4;
      13678: inst = 32'h8220000;
      13679: inst = 32'h10408000;
      13680: inst = 32'hc404f40;
      13681: inst = 32'h8220000;
      13682: inst = 32'h10408000;
      13683: inst = 32'hc404f4a;
      13684: inst = 32'h8220000;
      13685: inst = 32'h10408000;
      13686: inst = 32'hc404f54;
      13687: inst = 32'h8220000;
      13688: inst = 32'h10408000;
      13689: inst = 32'hc404fa0;
      13690: inst = 32'h8220000;
      13691: inst = 32'h10408000;
      13692: inst = 32'hc404faa;
      13693: inst = 32'h8220000;
      13694: inst = 32'h10408000;
      13695: inst = 32'hc404fb4;
      13696: inst = 32'h8220000;
      13697: inst = 32'h10408000;
      13698: inst = 32'hc405000;
      13699: inst = 32'h8220000;
      13700: inst = 32'h10408000;
      13701: inst = 32'hc40500a;
      13702: inst = 32'h8220000;
      13703: inst = 32'h10408000;
      13704: inst = 32'hc405014;
      13705: inst = 32'h8220000;
      13706: inst = 32'h10408000;
      13707: inst = 32'hc405060;
      13708: inst = 32'h8220000;
      13709: inst = 32'h10408000;
      13710: inst = 32'hc40506a;
      13711: inst = 32'h8220000;
      13712: inst = 32'h10408000;
      13713: inst = 32'hc405074;
      13714: inst = 32'h8220000;
      13715: inst = 32'h10408000;
      13716: inst = 32'hc4050c0;
      13717: inst = 32'h8220000;
      13718: inst = 32'h10408000;
      13719: inst = 32'hc4050ca;
      13720: inst = 32'h8220000;
      13721: inst = 32'h10408000;
      13722: inst = 32'hc4050d4;
      13723: inst = 32'h8220000;
      13724: inst = 32'h10408000;
      13725: inst = 32'hc405120;
      13726: inst = 32'h8220000;
      13727: inst = 32'h10408000;
      13728: inst = 32'hc40512a;
      13729: inst = 32'h8220000;
      13730: inst = 32'h10408000;
      13731: inst = 32'hc405134;
      13732: inst = 32'h8220000;
      13733: inst = 32'h10408000;
      13734: inst = 32'hc405180;
      13735: inst = 32'h8220000;
      13736: inst = 32'h10408000;
      13737: inst = 32'hc40518a;
      13738: inst = 32'h8220000;
      13739: inst = 32'h10408000;
      13740: inst = 32'hc405194;
      13741: inst = 32'h8220000;
      13742: inst = 32'h10408000;
      13743: inst = 32'hc4051a8;
      13744: inst = 32'h8220000;
      13745: inst = 32'h10408000;
      13746: inst = 32'hc4051a9;
      13747: inst = 32'h8220000;
      13748: inst = 32'h10408000;
      13749: inst = 32'hc4051b7;
      13750: inst = 32'h8220000;
      13751: inst = 32'h10408000;
      13752: inst = 32'hc4051e0;
      13753: inst = 32'h8220000;
      13754: inst = 32'h10408000;
      13755: inst = 32'hc4051ea;
      13756: inst = 32'h8220000;
      13757: inst = 32'h10408000;
      13758: inst = 32'hc4051f4;
      13759: inst = 32'h8220000;
      13760: inst = 32'h10408000;
      13761: inst = 32'hc405208;
      13762: inst = 32'h8220000;
      13763: inst = 32'h10408000;
      13764: inst = 32'hc405217;
      13765: inst = 32'h8220000;
      13766: inst = 32'h10408000;
      13767: inst = 32'hc405240;
      13768: inst = 32'h8220000;
      13769: inst = 32'h10408000;
      13770: inst = 32'hc40524a;
      13771: inst = 32'h8220000;
      13772: inst = 32'h10408000;
      13773: inst = 32'hc405254;
      13774: inst = 32'h8220000;
      13775: inst = 32'h10408000;
      13776: inst = 32'hc40525e;
      13777: inst = 32'h8220000;
      13778: inst = 32'h10408000;
      13779: inst = 32'hc405268;
      13780: inst = 32'h8220000;
      13781: inst = 32'h10408000;
      13782: inst = 32'hc405277;
      13783: inst = 32'h8220000;
      13784: inst = 32'h10408000;
      13785: inst = 32'hc405281;
      13786: inst = 32'h8220000;
      13787: inst = 32'h10408000;
      13788: inst = 32'hc4052a0;
      13789: inst = 32'h8220000;
      13790: inst = 32'h10408000;
      13791: inst = 32'hc4052a1;
      13792: inst = 32'h8220000;
      13793: inst = 32'h10408000;
      13794: inst = 32'hc4052a2;
      13795: inst = 32'h8220000;
      13796: inst = 32'h10408000;
      13797: inst = 32'hc4052a3;
      13798: inst = 32'h8220000;
      13799: inst = 32'h10408000;
      13800: inst = 32'hc4052a4;
      13801: inst = 32'h8220000;
      13802: inst = 32'h10408000;
      13803: inst = 32'hc4052a5;
      13804: inst = 32'h8220000;
      13805: inst = 32'h10408000;
      13806: inst = 32'hc4052a6;
      13807: inst = 32'h8220000;
      13808: inst = 32'h10408000;
      13809: inst = 32'hc4052a7;
      13810: inst = 32'h8220000;
      13811: inst = 32'h10408000;
      13812: inst = 32'hc4052a8;
      13813: inst = 32'h8220000;
      13814: inst = 32'h10408000;
      13815: inst = 32'hc4052a9;
      13816: inst = 32'h8220000;
      13817: inst = 32'h10408000;
      13818: inst = 32'hc4052aa;
      13819: inst = 32'h8220000;
      13820: inst = 32'h10408000;
      13821: inst = 32'hc4052ab;
      13822: inst = 32'h8220000;
      13823: inst = 32'h10408000;
      13824: inst = 32'hc4052ac;
      13825: inst = 32'h8220000;
      13826: inst = 32'h10408000;
      13827: inst = 32'hc4052ad;
      13828: inst = 32'h8220000;
      13829: inst = 32'h10408000;
      13830: inst = 32'hc4052ae;
      13831: inst = 32'h8220000;
      13832: inst = 32'h10408000;
      13833: inst = 32'hc4052af;
      13834: inst = 32'h8220000;
      13835: inst = 32'h10408000;
      13836: inst = 32'hc4052b0;
      13837: inst = 32'h8220000;
      13838: inst = 32'h10408000;
      13839: inst = 32'hc4052b1;
      13840: inst = 32'h8220000;
      13841: inst = 32'h10408000;
      13842: inst = 32'hc4052b2;
      13843: inst = 32'h8220000;
      13844: inst = 32'h10408000;
      13845: inst = 32'hc4052b3;
      13846: inst = 32'h8220000;
      13847: inst = 32'h10408000;
      13848: inst = 32'hc4052b4;
      13849: inst = 32'h8220000;
      13850: inst = 32'h10408000;
      13851: inst = 32'hc4052bd;
      13852: inst = 32'h8220000;
      13853: inst = 32'h10408000;
      13854: inst = 32'hc4052be;
      13855: inst = 32'h8220000;
      13856: inst = 32'h10408000;
      13857: inst = 32'hc4052c8;
      13858: inst = 32'h8220000;
      13859: inst = 32'h10408000;
      13860: inst = 32'hc4052d7;
      13861: inst = 32'h8220000;
      13862: inst = 32'h10408000;
      13863: inst = 32'hc4052e1;
      13864: inst = 32'h8220000;
      13865: inst = 32'h10408000;
      13866: inst = 32'hc4052e2;
      13867: inst = 32'h8220000;
      13868: inst = 32'h10408000;
      13869: inst = 32'hc40531c;
      13870: inst = 32'h8220000;
      13871: inst = 32'h10408000;
      13872: inst = 32'hc40531d;
      13873: inst = 32'h8220000;
      13874: inst = 32'h10408000;
      13875: inst = 32'hc40531e;
      13876: inst = 32'h8220000;
      13877: inst = 32'h10408000;
      13878: inst = 32'hc40531f;
      13879: inst = 32'h8220000;
      13880: inst = 32'h10408000;
      13881: inst = 32'hc405320;
      13882: inst = 32'h8220000;
      13883: inst = 32'h10408000;
      13884: inst = 32'hc405326;
      13885: inst = 32'h8220000;
      13886: inst = 32'h10408000;
      13887: inst = 32'hc405327;
      13888: inst = 32'h8220000;
      13889: inst = 32'h10408000;
      13890: inst = 32'hc405328;
      13891: inst = 32'h8220000;
      13892: inst = 32'h10408000;
      13893: inst = 32'hc405337;
      13894: inst = 32'h8220000;
      13895: inst = 32'h10408000;
      13896: inst = 32'hc405338;
      13897: inst = 32'h8220000;
      13898: inst = 32'h10408000;
      13899: inst = 32'hc405339;
      13900: inst = 32'h8220000;
      13901: inst = 32'h10408000;
      13902: inst = 32'hc40533f;
      13903: inst = 32'h8220000;
      13904: inst = 32'h10408000;
      13905: inst = 32'hc405340;
      13906: inst = 32'h8220000;
      13907: inst = 32'h10408000;
      13908: inst = 32'hc405341;
      13909: inst = 32'h8220000;
      13910: inst = 32'h10408000;
      13911: inst = 32'hc405342;
      13912: inst = 32'h8220000;
      13913: inst = 32'h10408000;
      13914: inst = 32'hc405343;
      13915: inst = 32'h8220000;
      13916: inst = 32'h10408000;
      13917: inst = 32'hc40537b;
      13918: inst = 32'h8220000;
      13919: inst = 32'h10408000;
      13920: inst = 32'hc40537c;
      13921: inst = 32'h8220000;
      13922: inst = 32'h10408000;
      13923: inst = 32'hc405386;
      13924: inst = 32'h8220000;
      13925: inst = 32'h10408000;
      13926: inst = 32'hc405387;
      13927: inst = 32'h8220000;
      13928: inst = 32'h10408000;
      13929: inst = 32'hc405388;
      13930: inst = 32'h8220000;
      13931: inst = 32'h10408000;
      13932: inst = 32'hc405397;
      13933: inst = 32'h8220000;
      13934: inst = 32'h10408000;
      13935: inst = 32'hc405398;
      13936: inst = 32'h8220000;
      13937: inst = 32'h10408000;
      13938: inst = 32'hc405399;
      13939: inst = 32'h8220000;
      13940: inst = 32'h10408000;
      13941: inst = 32'hc4053a3;
      13942: inst = 32'h8220000;
      13943: inst = 32'h10408000;
      13944: inst = 32'hc4053a4;
      13945: inst = 32'h8220000;
      13946: inst = 32'h10408000;
      13947: inst = 32'hc4053db;
      13948: inst = 32'h8220000;
      13949: inst = 32'h10408000;
      13950: inst = 32'hc4053e5;
      13951: inst = 32'h8220000;
      13952: inst = 32'h10408000;
      13953: inst = 32'hc4053e6;
      13954: inst = 32'h8220000;
      13955: inst = 32'h10408000;
      13956: inst = 32'hc4053e7;
      13957: inst = 32'h8220000;
      13958: inst = 32'h10408000;
      13959: inst = 32'hc4053f8;
      13960: inst = 32'h8220000;
      13961: inst = 32'h10408000;
      13962: inst = 32'hc4053f9;
      13963: inst = 32'h8220000;
      13964: inst = 32'h10408000;
      13965: inst = 32'hc4053fa;
      13966: inst = 32'h8220000;
      13967: inst = 32'h10408000;
      13968: inst = 32'hc405404;
      13969: inst = 32'h8220000;
      13970: inst = 32'h10408000;
      13971: inst = 32'hc40543a;
      13972: inst = 32'h8220000;
      13973: inst = 32'h10408000;
      13974: inst = 32'hc40543b;
      13975: inst = 32'h8220000;
      13976: inst = 32'h10408000;
      13977: inst = 32'hc405445;
      13978: inst = 32'h8220000;
      13979: inst = 32'h10408000;
      13980: inst = 32'hc405446;
      13981: inst = 32'h8220000;
      13982: inst = 32'h10408000;
      13983: inst = 32'hc405447;
      13984: inst = 32'h8220000;
      13985: inst = 32'h10408000;
      13986: inst = 32'hc405458;
      13987: inst = 32'h8220000;
      13988: inst = 32'h10408000;
      13989: inst = 32'hc405459;
      13990: inst = 32'h8220000;
      13991: inst = 32'h10408000;
      13992: inst = 32'hc40545a;
      13993: inst = 32'h8220000;
      13994: inst = 32'h10408000;
      13995: inst = 32'hc405464;
      13996: inst = 32'h8220000;
      13997: inst = 32'h10408000;
      13998: inst = 32'hc405465;
      13999: inst = 32'h8220000;
      14000: inst = 32'h10408000;
      14001: inst = 32'hc405499;
      14002: inst = 32'h8220000;
      14003: inst = 32'h10408000;
      14004: inst = 32'hc40549a;
      14005: inst = 32'h8220000;
      14006: inst = 32'h10408000;
      14007: inst = 32'hc4054a5;
      14008: inst = 32'h8220000;
      14009: inst = 32'h10408000;
      14010: inst = 32'hc4054a6;
      14011: inst = 32'h8220000;
      14012: inst = 32'h10408000;
      14013: inst = 32'hc4054a7;
      14014: inst = 32'h8220000;
      14015: inst = 32'h10408000;
      14016: inst = 32'hc4054b8;
      14017: inst = 32'h8220000;
      14018: inst = 32'h10408000;
      14019: inst = 32'hc4054b9;
      14020: inst = 32'h8220000;
      14021: inst = 32'h10408000;
      14022: inst = 32'hc4054ba;
      14023: inst = 32'h8220000;
      14024: inst = 32'h10408000;
      14025: inst = 32'hc4054c5;
      14026: inst = 32'h8220000;
      14027: inst = 32'h10408000;
      14028: inst = 32'hc4054c6;
      14029: inst = 32'h8220000;
      14030: inst = 32'h10408000;
      14031: inst = 32'hc4054f8;
      14032: inst = 32'h8220000;
      14033: inst = 32'h10408000;
      14034: inst = 32'hc4054f9;
      14035: inst = 32'h8220000;
      14036: inst = 32'h10408000;
      14037: inst = 32'hc405500;
      14038: inst = 32'h8220000;
      14039: inst = 32'h10408000;
      14040: inst = 32'hc405504;
      14041: inst = 32'h8220000;
      14042: inst = 32'h10408000;
      14043: inst = 32'hc405505;
      14044: inst = 32'h8220000;
      14045: inst = 32'h10408000;
      14046: inst = 32'hc405506;
      14047: inst = 32'h8220000;
      14048: inst = 32'h10408000;
      14049: inst = 32'hc405507;
      14050: inst = 32'h8220000;
      14051: inst = 32'h10408000;
      14052: inst = 32'hc405518;
      14053: inst = 32'h8220000;
      14054: inst = 32'h10408000;
      14055: inst = 32'hc405519;
      14056: inst = 32'h8220000;
      14057: inst = 32'h10408000;
      14058: inst = 32'hc40551a;
      14059: inst = 32'h8220000;
      14060: inst = 32'h10408000;
      14061: inst = 32'hc40551b;
      14062: inst = 32'h8220000;
      14063: inst = 32'h10408000;
      14064: inst = 32'hc40551f;
      14065: inst = 32'h8220000;
      14066: inst = 32'h10408000;
      14067: inst = 32'hc405526;
      14068: inst = 32'h8220000;
      14069: inst = 32'h10408000;
      14070: inst = 32'hc405527;
      14071: inst = 32'h8220000;
      14072: inst = 32'h10408000;
      14073: inst = 32'hc405558;
      14074: inst = 32'h8220000;
      14075: inst = 32'h10408000;
      14076: inst = 32'hc405559;
      14077: inst = 32'h8220000;
      14078: inst = 32'h10408000;
      14079: inst = 32'hc405560;
      14080: inst = 32'h8220000;
      14081: inst = 32'h10408000;
      14082: inst = 32'hc405564;
      14083: inst = 32'h8220000;
      14084: inst = 32'h10408000;
      14085: inst = 32'hc405565;
      14086: inst = 32'h8220000;
      14087: inst = 32'h10408000;
      14088: inst = 32'hc405566;
      14089: inst = 32'h8220000;
      14090: inst = 32'h10408000;
      14091: inst = 32'hc405567;
      14092: inst = 32'h8220000;
      14093: inst = 32'h10408000;
      14094: inst = 32'hc405578;
      14095: inst = 32'h8220000;
      14096: inst = 32'h10408000;
      14097: inst = 32'hc405579;
      14098: inst = 32'h8220000;
      14099: inst = 32'h10408000;
      14100: inst = 32'hc40557a;
      14101: inst = 32'h8220000;
      14102: inst = 32'h10408000;
      14103: inst = 32'hc40557b;
      14104: inst = 32'h8220000;
      14105: inst = 32'h10408000;
      14106: inst = 32'hc40557f;
      14107: inst = 32'h8220000;
      14108: inst = 32'h10408000;
      14109: inst = 32'hc405586;
      14110: inst = 32'h8220000;
      14111: inst = 32'h10408000;
      14112: inst = 32'hc405587;
      14113: inst = 32'h8220000;
      14114: inst = 32'h10408000;
      14115: inst = 32'hc4055b7;
      14116: inst = 32'h8220000;
      14117: inst = 32'h10408000;
      14118: inst = 32'hc4055b8;
      14119: inst = 32'h8220000;
      14120: inst = 32'h10408000;
      14121: inst = 32'hc4055bf;
      14122: inst = 32'h8220000;
      14123: inst = 32'h10408000;
      14124: inst = 32'hc4055c0;
      14125: inst = 32'h8220000;
      14126: inst = 32'h10408000;
      14127: inst = 32'hc4055c4;
      14128: inst = 32'h8220000;
      14129: inst = 32'h10408000;
      14130: inst = 32'hc4055c5;
      14131: inst = 32'h8220000;
      14132: inst = 32'h10408000;
      14133: inst = 32'hc4055c6;
      14134: inst = 32'h8220000;
      14135: inst = 32'h10408000;
      14136: inst = 32'hc4055c7;
      14137: inst = 32'h8220000;
      14138: inst = 32'h10408000;
      14139: inst = 32'hc4055d8;
      14140: inst = 32'h8220000;
      14141: inst = 32'h10408000;
      14142: inst = 32'hc4055d9;
      14143: inst = 32'h8220000;
      14144: inst = 32'h10408000;
      14145: inst = 32'hc4055da;
      14146: inst = 32'h8220000;
      14147: inst = 32'h10408000;
      14148: inst = 32'hc4055db;
      14149: inst = 32'h8220000;
      14150: inst = 32'h10408000;
      14151: inst = 32'hc4055df;
      14152: inst = 32'h8220000;
      14153: inst = 32'h10408000;
      14154: inst = 32'hc4055e0;
      14155: inst = 32'h8220000;
      14156: inst = 32'h10408000;
      14157: inst = 32'hc4055e7;
      14158: inst = 32'h8220000;
      14159: inst = 32'h10408000;
      14160: inst = 32'hc4055e8;
      14161: inst = 32'h8220000;
      14162: inst = 32'h10408000;
      14163: inst = 32'hc405616;
      14164: inst = 32'h8220000;
      14165: inst = 32'h10408000;
      14166: inst = 32'hc405617;
      14167: inst = 32'h8220000;
      14168: inst = 32'h10408000;
      14169: inst = 32'hc40561f;
      14170: inst = 32'h8220000;
      14171: inst = 32'h10408000;
      14172: inst = 32'hc405620;
      14173: inst = 32'h8220000;
      14174: inst = 32'h10408000;
      14175: inst = 32'hc405623;
      14176: inst = 32'h8220000;
      14177: inst = 32'h10408000;
      14178: inst = 32'hc405624;
      14179: inst = 32'h8220000;
      14180: inst = 32'h10408000;
      14181: inst = 32'hc405625;
      14182: inst = 32'h8220000;
      14183: inst = 32'h10408000;
      14184: inst = 32'hc405626;
      14185: inst = 32'h8220000;
      14186: inst = 32'h10408000;
      14187: inst = 32'hc405639;
      14188: inst = 32'h8220000;
      14189: inst = 32'h10408000;
      14190: inst = 32'hc40563a;
      14191: inst = 32'h8220000;
      14192: inst = 32'h10408000;
      14193: inst = 32'hc40563b;
      14194: inst = 32'h8220000;
      14195: inst = 32'h10408000;
      14196: inst = 32'hc40563c;
      14197: inst = 32'h8220000;
      14198: inst = 32'h10408000;
      14199: inst = 32'hc40563f;
      14200: inst = 32'h8220000;
      14201: inst = 32'h10408000;
      14202: inst = 32'hc405640;
      14203: inst = 32'h8220000;
      14204: inst = 32'h10408000;
      14205: inst = 32'hc405648;
      14206: inst = 32'h8220000;
      14207: inst = 32'h10408000;
      14208: inst = 32'hc405649;
      14209: inst = 32'h8220000;
      14210: inst = 32'h10408000;
      14211: inst = 32'hc405675;
      14212: inst = 32'h8220000;
      14213: inst = 32'h10408000;
      14214: inst = 32'hc405676;
      14215: inst = 32'h8220000;
      14216: inst = 32'h10408000;
      14217: inst = 32'hc405677;
      14218: inst = 32'h8220000;
      14219: inst = 32'h10408000;
      14220: inst = 32'hc40567e;
      14221: inst = 32'h8220000;
      14222: inst = 32'h10408000;
      14223: inst = 32'hc40567f;
      14224: inst = 32'h8220000;
      14225: inst = 32'h10408000;
      14226: inst = 32'hc405680;
      14227: inst = 32'h8220000;
      14228: inst = 32'h10408000;
      14229: inst = 32'hc405683;
      14230: inst = 32'h8220000;
      14231: inst = 32'h10408000;
      14232: inst = 32'hc405684;
      14233: inst = 32'h8220000;
      14234: inst = 32'h10408000;
      14235: inst = 32'hc405685;
      14236: inst = 32'h8220000;
      14237: inst = 32'h10408000;
      14238: inst = 32'hc405686;
      14239: inst = 32'h8220000;
      14240: inst = 32'h10408000;
      14241: inst = 32'hc405699;
      14242: inst = 32'h8220000;
      14243: inst = 32'h10408000;
      14244: inst = 32'hc40569a;
      14245: inst = 32'h8220000;
      14246: inst = 32'h10408000;
      14247: inst = 32'hc40569b;
      14248: inst = 32'h8220000;
      14249: inst = 32'h10408000;
      14250: inst = 32'hc40569c;
      14251: inst = 32'h8220000;
      14252: inst = 32'h10408000;
      14253: inst = 32'hc40569f;
      14254: inst = 32'h8220000;
      14255: inst = 32'h10408000;
      14256: inst = 32'hc4056a0;
      14257: inst = 32'h8220000;
      14258: inst = 32'h10408000;
      14259: inst = 32'hc4056a1;
      14260: inst = 32'h8220000;
      14261: inst = 32'h10408000;
      14262: inst = 32'hc4056a8;
      14263: inst = 32'h8220000;
      14264: inst = 32'h10408000;
      14265: inst = 32'hc4056a9;
      14266: inst = 32'h8220000;
      14267: inst = 32'h10408000;
      14268: inst = 32'hc4056aa;
      14269: inst = 32'h8220000;
      14270: inst = 32'h10408000;
      14271: inst = 32'hc4056d4;
      14272: inst = 32'h8220000;
      14273: inst = 32'h10408000;
      14274: inst = 32'hc4056d5;
      14275: inst = 32'h8220000;
      14276: inst = 32'h10408000;
      14277: inst = 32'hc4056d6;
      14278: inst = 32'h8220000;
      14279: inst = 32'h10408000;
      14280: inst = 32'hc4056d7;
      14281: inst = 32'h8220000;
      14282: inst = 32'h10408000;
      14283: inst = 32'hc4056d8;
      14284: inst = 32'h8220000;
      14285: inst = 32'h10408000;
      14286: inst = 32'hc4056d9;
      14287: inst = 32'h8220000;
      14288: inst = 32'h10408000;
      14289: inst = 32'hc4056da;
      14290: inst = 32'h8220000;
      14291: inst = 32'h10408000;
      14292: inst = 32'hc4056db;
      14293: inst = 32'h8220000;
      14294: inst = 32'h10408000;
      14295: inst = 32'hc4056dc;
      14296: inst = 32'h8220000;
      14297: inst = 32'h10408000;
      14298: inst = 32'hc4056dd;
      14299: inst = 32'h8220000;
      14300: inst = 32'h10408000;
      14301: inst = 32'hc4056de;
      14302: inst = 32'h8220000;
      14303: inst = 32'h10408000;
      14304: inst = 32'hc4056df;
      14305: inst = 32'h8220000;
      14306: inst = 32'h10408000;
      14307: inst = 32'hc4056e0;
      14308: inst = 32'h8220000;
      14309: inst = 32'h10408000;
      14310: inst = 32'hc4056e3;
      14311: inst = 32'h8220000;
      14312: inst = 32'h10408000;
      14313: inst = 32'hc4056e4;
      14314: inst = 32'h8220000;
      14315: inst = 32'h10408000;
      14316: inst = 32'hc4056e5;
      14317: inst = 32'h8220000;
      14318: inst = 32'h10408000;
      14319: inst = 32'hc4056e6;
      14320: inst = 32'h8220000;
      14321: inst = 32'h10408000;
      14322: inst = 32'hc4056f9;
      14323: inst = 32'h8220000;
      14324: inst = 32'h10408000;
      14325: inst = 32'hc4056fa;
      14326: inst = 32'h8220000;
      14327: inst = 32'h10408000;
      14328: inst = 32'hc4056fb;
      14329: inst = 32'h8220000;
      14330: inst = 32'h10408000;
      14331: inst = 32'hc4056fc;
      14332: inst = 32'h8220000;
      14333: inst = 32'h10408000;
      14334: inst = 32'hc4056ff;
      14335: inst = 32'h8220000;
      14336: inst = 32'h10408000;
      14337: inst = 32'hc405700;
      14338: inst = 32'h8220000;
      14339: inst = 32'h10408000;
      14340: inst = 32'hc405701;
      14341: inst = 32'h8220000;
      14342: inst = 32'h10408000;
      14343: inst = 32'hc405702;
      14344: inst = 32'h8220000;
      14345: inst = 32'h10408000;
      14346: inst = 32'hc405703;
      14347: inst = 32'h8220000;
      14348: inst = 32'h10408000;
      14349: inst = 32'hc405704;
      14350: inst = 32'h8220000;
      14351: inst = 32'h10408000;
      14352: inst = 32'hc405705;
      14353: inst = 32'h8220000;
      14354: inst = 32'h10408000;
      14355: inst = 32'hc405706;
      14356: inst = 32'h8220000;
      14357: inst = 32'h10408000;
      14358: inst = 32'hc405707;
      14359: inst = 32'h8220000;
      14360: inst = 32'h10408000;
      14361: inst = 32'hc405708;
      14362: inst = 32'h8220000;
      14363: inst = 32'h10408000;
      14364: inst = 32'hc405709;
      14365: inst = 32'h8220000;
      14366: inst = 32'h10408000;
      14367: inst = 32'hc40570a;
      14368: inst = 32'h8220000;
      14369: inst = 32'h10408000;
      14370: inst = 32'hc405734;
      14371: inst = 32'h8220000;
      14372: inst = 32'h10408000;
      14373: inst = 32'hc405735;
      14374: inst = 32'h8220000;
      14375: inst = 32'h10408000;
      14376: inst = 32'hc405736;
      14377: inst = 32'h8220000;
      14378: inst = 32'h10408000;
      14379: inst = 32'hc405737;
      14380: inst = 32'h8220000;
      14381: inst = 32'h10408000;
      14382: inst = 32'hc405738;
      14383: inst = 32'h8220000;
      14384: inst = 32'h10408000;
      14385: inst = 32'hc405739;
      14386: inst = 32'h8220000;
      14387: inst = 32'h10408000;
      14388: inst = 32'hc40573a;
      14389: inst = 32'h8220000;
      14390: inst = 32'h10408000;
      14391: inst = 32'hc40573b;
      14392: inst = 32'h8220000;
      14393: inst = 32'h10408000;
      14394: inst = 32'hc40573c;
      14395: inst = 32'h8220000;
      14396: inst = 32'h10408000;
      14397: inst = 32'hc40573d;
      14398: inst = 32'h8220000;
      14399: inst = 32'h10408000;
      14400: inst = 32'hc40573e;
      14401: inst = 32'h8220000;
      14402: inst = 32'h10408000;
      14403: inst = 32'hc40573f;
      14404: inst = 32'h8220000;
      14405: inst = 32'h10408000;
      14406: inst = 32'hc405740;
      14407: inst = 32'h8220000;
      14408: inst = 32'h10408000;
      14409: inst = 32'hc405742;
      14410: inst = 32'h8220000;
      14411: inst = 32'h10408000;
      14412: inst = 32'hc405743;
      14413: inst = 32'h8220000;
      14414: inst = 32'h10408000;
      14415: inst = 32'hc405744;
      14416: inst = 32'h8220000;
      14417: inst = 32'h10408000;
      14418: inst = 32'hc405745;
      14419: inst = 32'h8220000;
      14420: inst = 32'h10408000;
      14421: inst = 32'hc405746;
      14422: inst = 32'h8220000;
      14423: inst = 32'h10408000;
      14424: inst = 32'hc405759;
      14425: inst = 32'h8220000;
      14426: inst = 32'h10408000;
      14427: inst = 32'hc40575a;
      14428: inst = 32'h8220000;
      14429: inst = 32'h10408000;
      14430: inst = 32'hc40575b;
      14431: inst = 32'h8220000;
      14432: inst = 32'h10408000;
      14433: inst = 32'hc40575c;
      14434: inst = 32'h8220000;
      14435: inst = 32'h10408000;
      14436: inst = 32'hc40575d;
      14437: inst = 32'h8220000;
      14438: inst = 32'h10408000;
      14439: inst = 32'hc40575f;
      14440: inst = 32'h8220000;
      14441: inst = 32'h10408000;
      14442: inst = 32'hc405760;
      14443: inst = 32'h8220000;
      14444: inst = 32'h10408000;
      14445: inst = 32'hc405761;
      14446: inst = 32'h8220000;
      14447: inst = 32'h10408000;
      14448: inst = 32'hc405762;
      14449: inst = 32'h8220000;
      14450: inst = 32'h10408000;
      14451: inst = 32'hc405763;
      14452: inst = 32'h8220000;
      14453: inst = 32'h10408000;
      14454: inst = 32'hc405764;
      14455: inst = 32'h8220000;
      14456: inst = 32'h10408000;
      14457: inst = 32'hc405765;
      14458: inst = 32'h8220000;
      14459: inst = 32'h10408000;
      14460: inst = 32'hc405766;
      14461: inst = 32'h8220000;
      14462: inst = 32'h10408000;
      14463: inst = 32'hc405767;
      14464: inst = 32'h8220000;
      14465: inst = 32'h10408000;
      14466: inst = 32'hc405768;
      14467: inst = 32'h8220000;
      14468: inst = 32'h10408000;
      14469: inst = 32'hc405769;
      14470: inst = 32'h8220000;
      14471: inst = 32'h10408000;
      14472: inst = 32'hc40576a;
      14473: inst = 32'h8220000;
      14474: inst = 32'h10408000;
      14475: inst = 32'hc40576b;
      14476: inst = 32'h8220000;
      14477: inst = 32'h10408000;
      14478: inst = 32'hc405793;
      14479: inst = 32'h8220000;
      14480: inst = 32'h10408000;
      14481: inst = 32'hc405794;
      14482: inst = 32'h8220000;
      14483: inst = 32'h10408000;
      14484: inst = 32'hc405795;
      14485: inst = 32'h8220000;
      14486: inst = 32'h10408000;
      14487: inst = 32'hc405796;
      14488: inst = 32'h8220000;
      14489: inst = 32'h10408000;
      14490: inst = 32'hc405797;
      14491: inst = 32'h8220000;
      14492: inst = 32'h10408000;
      14493: inst = 32'hc405798;
      14494: inst = 32'h8220000;
      14495: inst = 32'h10408000;
      14496: inst = 32'hc405799;
      14497: inst = 32'h8220000;
      14498: inst = 32'h10408000;
      14499: inst = 32'hc40579a;
      14500: inst = 32'h8220000;
      14501: inst = 32'h10408000;
      14502: inst = 32'hc40579b;
      14503: inst = 32'h8220000;
      14504: inst = 32'h10408000;
      14505: inst = 32'hc40579c;
      14506: inst = 32'h8220000;
      14507: inst = 32'h10408000;
      14508: inst = 32'hc40579d;
      14509: inst = 32'h8220000;
      14510: inst = 32'h10408000;
      14511: inst = 32'hc40579e;
      14512: inst = 32'h8220000;
      14513: inst = 32'h10408000;
      14514: inst = 32'hc40579f;
      14515: inst = 32'h8220000;
      14516: inst = 32'h10408000;
      14517: inst = 32'hc4057a0;
      14518: inst = 32'h8220000;
      14519: inst = 32'h10408000;
      14520: inst = 32'hc4057a1;
      14521: inst = 32'h8220000;
      14522: inst = 32'h10408000;
      14523: inst = 32'hc4057a2;
      14524: inst = 32'h8220000;
      14525: inst = 32'h10408000;
      14526: inst = 32'hc4057a3;
      14527: inst = 32'h8220000;
      14528: inst = 32'h10408000;
      14529: inst = 32'hc4057a4;
      14530: inst = 32'h8220000;
      14531: inst = 32'h10408000;
      14532: inst = 32'hc4057a5;
      14533: inst = 32'h8220000;
      14534: inst = 32'h10408000;
      14535: inst = 32'hc4057a6;
      14536: inst = 32'h8220000;
      14537: inst = 32'h10408000;
      14538: inst = 32'hc4057b9;
      14539: inst = 32'h8220000;
      14540: inst = 32'h10408000;
      14541: inst = 32'hc4057ba;
      14542: inst = 32'h8220000;
      14543: inst = 32'h10408000;
      14544: inst = 32'hc4057bb;
      14545: inst = 32'h8220000;
      14546: inst = 32'h10408000;
      14547: inst = 32'hc4057bc;
      14548: inst = 32'h8220000;
      14549: inst = 32'h10408000;
      14550: inst = 32'hc4057bd;
      14551: inst = 32'h8220000;
      14552: inst = 32'h10408000;
      14553: inst = 32'hc4057be;
      14554: inst = 32'h8220000;
      14555: inst = 32'h10408000;
      14556: inst = 32'hc4057bf;
      14557: inst = 32'h8220000;
      14558: inst = 32'h10408000;
      14559: inst = 32'hc4057c0;
      14560: inst = 32'h8220000;
      14561: inst = 32'h10408000;
      14562: inst = 32'hc4057c1;
      14563: inst = 32'h8220000;
      14564: inst = 32'h10408000;
      14565: inst = 32'hc4057c2;
      14566: inst = 32'h8220000;
      14567: inst = 32'h10408000;
      14568: inst = 32'hc4057c3;
      14569: inst = 32'h8220000;
      14570: inst = 32'h10408000;
      14571: inst = 32'hc4057c4;
      14572: inst = 32'h8220000;
      14573: inst = 32'h10408000;
      14574: inst = 32'hc4057c5;
      14575: inst = 32'h8220000;
      14576: inst = 32'h10408000;
      14577: inst = 32'hc4057c6;
      14578: inst = 32'h8220000;
      14579: inst = 32'h10408000;
      14580: inst = 32'hc4057c7;
      14581: inst = 32'h8220000;
      14582: inst = 32'h10408000;
      14583: inst = 32'hc4057c8;
      14584: inst = 32'h8220000;
      14585: inst = 32'h10408000;
      14586: inst = 32'hc4057c9;
      14587: inst = 32'h8220000;
      14588: inst = 32'h10408000;
      14589: inst = 32'hc4057ca;
      14590: inst = 32'h8220000;
      14591: inst = 32'h10408000;
      14592: inst = 32'hc4057cb;
      14593: inst = 32'h8220000;
      14594: inst = 32'h10408000;
      14595: inst = 32'hc4057cc;
      14596: inst = 32'h8220000;
      14597: inst = 32'hc20bdd7;
      14598: inst = 32'h10408000;
      14599: inst = 32'hc404dc1;
      14600: inst = 32'h8220000;
      14601: inst = 32'h10408000;
      14602: inst = 32'hc404dc2;
      14603: inst = 32'h8220000;
      14604: inst = 32'h10408000;
      14605: inst = 32'hc404dc3;
      14606: inst = 32'h8220000;
      14607: inst = 32'h10408000;
      14608: inst = 32'hc404dc4;
      14609: inst = 32'h8220000;
      14610: inst = 32'h10408000;
      14611: inst = 32'hc404dc5;
      14612: inst = 32'h8220000;
      14613: inst = 32'h10408000;
      14614: inst = 32'hc404dc6;
      14615: inst = 32'h8220000;
      14616: inst = 32'h10408000;
      14617: inst = 32'hc404dc7;
      14618: inst = 32'h8220000;
      14619: inst = 32'h10408000;
      14620: inst = 32'hc404dc8;
      14621: inst = 32'h8220000;
      14622: inst = 32'h10408000;
      14623: inst = 32'hc404dc9;
      14624: inst = 32'h8220000;
      14625: inst = 32'h10408000;
      14626: inst = 32'hc404dcb;
      14627: inst = 32'h8220000;
      14628: inst = 32'h10408000;
      14629: inst = 32'hc404dcc;
      14630: inst = 32'h8220000;
      14631: inst = 32'h10408000;
      14632: inst = 32'hc404dcd;
      14633: inst = 32'h8220000;
      14634: inst = 32'h10408000;
      14635: inst = 32'hc404dce;
      14636: inst = 32'h8220000;
      14637: inst = 32'h10408000;
      14638: inst = 32'hc404dcf;
      14639: inst = 32'h8220000;
      14640: inst = 32'h10408000;
      14641: inst = 32'hc404dd0;
      14642: inst = 32'h8220000;
      14643: inst = 32'h10408000;
      14644: inst = 32'hc404dd1;
      14645: inst = 32'h8220000;
      14646: inst = 32'h10408000;
      14647: inst = 32'hc404dd2;
      14648: inst = 32'h8220000;
      14649: inst = 32'h10408000;
      14650: inst = 32'hc404dd3;
      14651: inst = 32'h8220000;
      14652: inst = 32'h10408000;
      14653: inst = 32'hc404e21;
      14654: inst = 32'h8220000;
      14655: inst = 32'h10408000;
      14656: inst = 32'hc404e22;
      14657: inst = 32'h8220000;
      14658: inst = 32'h10408000;
      14659: inst = 32'hc404e23;
      14660: inst = 32'h8220000;
      14661: inst = 32'h10408000;
      14662: inst = 32'hc404e24;
      14663: inst = 32'h8220000;
      14664: inst = 32'h10408000;
      14665: inst = 32'hc404e25;
      14666: inst = 32'h8220000;
      14667: inst = 32'h10408000;
      14668: inst = 32'hc404e26;
      14669: inst = 32'h8220000;
      14670: inst = 32'h10408000;
      14671: inst = 32'hc404e27;
      14672: inst = 32'h8220000;
      14673: inst = 32'h10408000;
      14674: inst = 32'hc404e28;
      14675: inst = 32'h8220000;
      14676: inst = 32'h10408000;
      14677: inst = 32'hc404e29;
      14678: inst = 32'h8220000;
      14679: inst = 32'h10408000;
      14680: inst = 32'hc404e2b;
      14681: inst = 32'h8220000;
      14682: inst = 32'h10408000;
      14683: inst = 32'hc404e2c;
      14684: inst = 32'h8220000;
      14685: inst = 32'h10408000;
      14686: inst = 32'hc404e2d;
      14687: inst = 32'h8220000;
      14688: inst = 32'h10408000;
      14689: inst = 32'hc404e2e;
      14690: inst = 32'h8220000;
      14691: inst = 32'h10408000;
      14692: inst = 32'hc404e2f;
      14693: inst = 32'h8220000;
      14694: inst = 32'h10408000;
      14695: inst = 32'hc404e30;
      14696: inst = 32'h8220000;
      14697: inst = 32'h10408000;
      14698: inst = 32'hc404e31;
      14699: inst = 32'h8220000;
      14700: inst = 32'h10408000;
      14701: inst = 32'hc404e32;
      14702: inst = 32'h8220000;
      14703: inst = 32'h10408000;
      14704: inst = 32'hc404e33;
      14705: inst = 32'h8220000;
      14706: inst = 32'h10408000;
      14707: inst = 32'hc404e81;
      14708: inst = 32'h8220000;
      14709: inst = 32'h10408000;
      14710: inst = 32'hc404e82;
      14711: inst = 32'h8220000;
      14712: inst = 32'h10408000;
      14713: inst = 32'hc404e83;
      14714: inst = 32'h8220000;
      14715: inst = 32'h10408000;
      14716: inst = 32'hc404e84;
      14717: inst = 32'h8220000;
      14718: inst = 32'h10408000;
      14719: inst = 32'hc404e85;
      14720: inst = 32'h8220000;
      14721: inst = 32'h10408000;
      14722: inst = 32'hc404e86;
      14723: inst = 32'h8220000;
      14724: inst = 32'h10408000;
      14725: inst = 32'hc404e87;
      14726: inst = 32'h8220000;
      14727: inst = 32'h10408000;
      14728: inst = 32'hc404e88;
      14729: inst = 32'h8220000;
      14730: inst = 32'h10408000;
      14731: inst = 32'hc404e89;
      14732: inst = 32'h8220000;
      14733: inst = 32'h10408000;
      14734: inst = 32'hc404e8b;
      14735: inst = 32'h8220000;
      14736: inst = 32'h10408000;
      14737: inst = 32'hc404e8c;
      14738: inst = 32'h8220000;
      14739: inst = 32'h10408000;
      14740: inst = 32'hc404e8d;
      14741: inst = 32'h8220000;
      14742: inst = 32'h10408000;
      14743: inst = 32'hc404e8e;
      14744: inst = 32'h8220000;
      14745: inst = 32'h10408000;
      14746: inst = 32'hc404e8f;
      14747: inst = 32'h8220000;
      14748: inst = 32'h10408000;
      14749: inst = 32'hc404e90;
      14750: inst = 32'h8220000;
      14751: inst = 32'h10408000;
      14752: inst = 32'hc404e91;
      14753: inst = 32'h8220000;
      14754: inst = 32'h10408000;
      14755: inst = 32'hc404e92;
      14756: inst = 32'h8220000;
      14757: inst = 32'h10408000;
      14758: inst = 32'hc404e93;
      14759: inst = 32'h8220000;
      14760: inst = 32'h10408000;
      14761: inst = 32'hc404ee1;
      14762: inst = 32'h8220000;
      14763: inst = 32'h10408000;
      14764: inst = 32'hc404ee2;
      14765: inst = 32'h8220000;
      14766: inst = 32'h10408000;
      14767: inst = 32'hc404ee3;
      14768: inst = 32'h8220000;
      14769: inst = 32'h10408000;
      14770: inst = 32'hc404ee4;
      14771: inst = 32'h8220000;
      14772: inst = 32'h10408000;
      14773: inst = 32'hc404ee5;
      14774: inst = 32'h8220000;
      14775: inst = 32'h10408000;
      14776: inst = 32'hc404ee6;
      14777: inst = 32'h8220000;
      14778: inst = 32'h10408000;
      14779: inst = 32'hc404ee7;
      14780: inst = 32'h8220000;
      14781: inst = 32'h10408000;
      14782: inst = 32'hc404ee8;
      14783: inst = 32'h8220000;
      14784: inst = 32'h10408000;
      14785: inst = 32'hc404ee9;
      14786: inst = 32'h8220000;
      14787: inst = 32'h10408000;
      14788: inst = 32'hc404eeb;
      14789: inst = 32'h8220000;
      14790: inst = 32'h10408000;
      14791: inst = 32'hc404eec;
      14792: inst = 32'h8220000;
      14793: inst = 32'h10408000;
      14794: inst = 32'hc404eed;
      14795: inst = 32'h8220000;
      14796: inst = 32'h10408000;
      14797: inst = 32'hc404eee;
      14798: inst = 32'h8220000;
      14799: inst = 32'h10408000;
      14800: inst = 32'hc404eef;
      14801: inst = 32'h8220000;
      14802: inst = 32'h10408000;
      14803: inst = 32'hc404ef0;
      14804: inst = 32'h8220000;
      14805: inst = 32'h10408000;
      14806: inst = 32'hc404ef1;
      14807: inst = 32'h8220000;
      14808: inst = 32'h10408000;
      14809: inst = 32'hc404ef2;
      14810: inst = 32'h8220000;
      14811: inst = 32'h10408000;
      14812: inst = 32'hc404ef3;
      14813: inst = 32'h8220000;
      14814: inst = 32'h10408000;
      14815: inst = 32'hc404f41;
      14816: inst = 32'h8220000;
      14817: inst = 32'h10408000;
      14818: inst = 32'hc404f42;
      14819: inst = 32'h8220000;
      14820: inst = 32'h10408000;
      14821: inst = 32'hc404f43;
      14822: inst = 32'h8220000;
      14823: inst = 32'h10408000;
      14824: inst = 32'hc404f44;
      14825: inst = 32'h8220000;
      14826: inst = 32'h10408000;
      14827: inst = 32'hc404f45;
      14828: inst = 32'h8220000;
      14829: inst = 32'h10408000;
      14830: inst = 32'hc404f46;
      14831: inst = 32'h8220000;
      14832: inst = 32'h10408000;
      14833: inst = 32'hc404f47;
      14834: inst = 32'h8220000;
      14835: inst = 32'h10408000;
      14836: inst = 32'hc404f48;
      14837: inst = 32'h8220000;
      14838: inst = 32'h10408000;
      14839: inst = 32'hc404f49;
      14840: inst = 32'h8220000;
      14841: inst = 32'h10408000;
      14842: inst = 32'hc404f4b;
      14843: inst = 32'h8220000;
      14844: inst = 32'h10408000;
      14845: inst = 32'hc404f4c;
      14846: inst = 32'h8220000;
      14847: inst = 32'h10408000;
      14848: inst = 32'hc404f4d;
      14849: inst = 32'h8220000;
      14850: inst = 32'h10408000;
      14851: inst = 32'hc404f4e;
      14852: inst = 32'h8220000;
      14853: inst = 32'h10408000;
      14854: inst = 32'hc404f4f;
      14855: inst = 32'h8220000;
      14856: inst = 32'h10408000;
      14857: inst = 32'hc404f50;
      14858: inst = 32'h8220000;
      14859: inst = 32'h10408000;
      14860: inst = 32'hc404f51;
      14861: inst = 32'h8220000;
      14862: inst = 32'h10408000;
      14863: inst = 32'hc404f52;
      14864: inst = 32'h8220000;
      14865: inst = 32'h10408000;
      14866: inst = 32'hc404f53;
      14867: inst = 32'h8220000;
      14868: inst = 32'h10408000;
      14869: inst = 32'hc404fa1;
      14870: inst = 32'h8220000;
      14871: inst = 32'h10408000;
      14872: inst = 32'hc404fa2;
      14873: inst = 32'h8220000;
      14874: inst = 32'h10408000;
      14875: inst = 32'hc404fa3;
      14876: inst = 32'h8220000;
      14877: inst = 32'h10408000;
      14878: inst = 32'hc404fa4;
      14879: inst = 32'h8220000;
      14880: inst = 32'h10408000;
      14881: inst = 32'hc404fa5;
      14882: inst = 32'h8220000;
      14883: inst = 32'h10408000;
      14884: inst = 32'hc404fa6;
      14885: inst = 32'h8220000;
      14886: inst = 32'h10408000;
      14887: inst = 32'hc404fa7;
      14888: inst = 32'h8220000;
      14889: inst = 32'h10408000;
      14890: inst = 32'hc404fa9;
      14891: inst = 32'h8220000;
      14892: inst = 32'h10408000;
      14893: inst = 32'hc404fab;
      14894: inst = 32'h8220000;
      14895: inst = 32'h10408000;
      14896: inst = 32'hc404fad;
      14897: inst = 32'h8220000;
      14898: inst = 32'h10408000;
      14899: inst = 32'hc404fae;
      14900: inst = 32'h8220000;
      14901: inst = 32'h10408000;
      14902: inst = 32'hc404faf;
      14903: inst = 32'h8220000;
      14904: inst = 32'h10408000;
      14905: inst = 32'hc404fb0;
      14906: inst = 32'h8220000;
      14907: inst = 32'h10408000;
      14908: inst = 32'hc404fb1;
      14909: inst = 32'h8220000;
      14910: inst = 32'h10408000;
      14911: inst = 32'hc404fb2;
      14912: inst = 32'h8220000;
      14913: inst = 32'h10408000;
      14914: inst = 32'hc404fb3;
      14915: inst = 32'h8220000;
      14916: inst = 32'h10408000;
      14917: inst = 32'hc405001;
      14918: inst = 32'h8220000;
      14919: inst = 32'h10408000;
      14920: inst = 32'hc405002;
      14921: inst = 32'h8220000;
      14922: inst = 32'h10408000;
      14923: inst = 32'hc405003;
      14924: inst = 32'h8220000;
      14925: inst = 32'h10408000;
      14926: inst = 32'hc405004;
      14927: inst = 32'h8220000;
      14928: inst = 32'h10408000;
      14929: inst = 32'hc405005;
      14930: inst = 32'h8220000;
      14931: inst = 32'h10408000;
      14932: inst = 32'hc405006;
      14933: inst = 32'h8220000;
      14934: inst = 32'h10408000;
      14935: inst = 32'hc405007;
      14936: inst = 32'h8220000;
      14937: inst = 32'h10408000;
      14938: inst = 32'hc405009;
      14939: inst = 32'h8220000;
      14940: inst = 32'h10408000;
      14941: inst = 32'hc40500b;
      14942: inst = 32'h8220000;
      14943: inst = 32'h10408000;
      14944: inst = 32'hc40500d;
      14945: inst = 32'h8220000;
      14946: inst = 32'h10408000;
      14947: inst = 32'hc40500e;
      14948: inst = 32'h8220000;
      14949: inst = 32'h10408000;
      14950: inst = 32'hc40500f;
      14951: inst = 32'h8220000;
      14952: inst = 32'h10408000;
      14953: inst = 32'hc405010;
      14954: inst = 32'h8220000;
      14955: inst = 32'h10408000;
      14956: inst = 32'hc405011;
      14957: inst = 32'h8220000;
      14958: inst = 32'h10408000;
      14959: inst = 32'hc405012;
      14960: inst = 32'h8220000;
      14961: inst = 32'h10408000;
      14962: inst = 32'hc405013;
      14963: inst = 32'h8220000;
      14964: inst = 32'h10408000;
      14965: inst = 32'hc405061;
      14966: inst = 32'h8220000;
      14967: inst = 32'h10408000;
      14968: inst = 32'hc405062;
      14969: inst = 32'h8220000;
      14970: inst = 32'h10408000;
      14971: inst = 32'hc405063;
      14972: inst = 32'h8220000;
      14973: inst = 32'h10408000;
      14974: inst = 32'hc405064;
      14975: inst = 32'h8220000;
      14976: inst = 32'h10408000;
      14977: inst = 32'hc405065;
      14978: inst = 32'h8220000;
      14979: inst = 32'h10408000;
      14980: inst = 32'hc405066;
      14981: inst = 32'h8220000;
      14982: inst = 32'h10408000;
      14983: inst = 32'hc405067;
      14984: inst = 32'h8220000;
      14985: inst = 32'h10408000;
      14986: inst = 32'hc405068;
      14987: inst = 32'h8220000;
      14988: inst = 32'h10408000;
      14989: inst = 32'hc405069;
      14990: inst = 32'h8220000;
      14991: inst = 32'h10408000;
      14992: inst = 32'hc40506b;
      14993: inst = 32'h8220000;
      14994: inst = 32'h10408000;
      14995: inst = 32'hc40506c;
      14996: inst = 32'h8220000;
      14997: inst = 32'h10408000;
      14998: inst = 32'hc40506d;
      14999: inst = 32'h8220000;
      15000: inst = 32'h10408000;
      15001: inst = 32'hc40506e;
      15002: inst = 32'h8220000;
      15003: inst = 32'h10408000;
      15004: inst = 32'hc40506f;
      15005: inst = 32'h8220000;
      15006: inst = 32'h10408000;
      15007: inst = 32'hc405070;
      15008: inst = 32'h8220000;
      15009: inst = 32'h10408000;
      15010: inst = 32'hc405071;
      15011: inst = 32'h8220000;
      15012: inst = 32'h10408000;
      15013: inst = 32'hc405072;
      15014: inst = 32'h8220000;
      15015: inst = 32'h10408000;
      15016: inst = 32'hc405073;
      15017: inst = 32'h8220000;
      15018: inst = 32'h10408000;
      15019: inst = 32'hc4050c1;
      15020: inst = 32'h8220000;
      15021: inst = 32'h10408000;
      15022: inst = 32'hc4050c2;
      15023: inst = 32'h8220000;
      15024: inst = 32'h10408000;
      15025: inst = 32'hc4050c3;
      15026: inst = 32'h8220000;
      15027: inst = 32'h10408000;
      15028: inst = 32'hc4050c4;
      15029: inst = 32'h8220000;
      15030: inst = 32'h10408000;
      15031: inst = 32'hc4050c5;
      15032: inst = 32'h8220000;
      15033: inst = 32'h10408000;
      15034: inst = 32'hc4050c6;
      15035: inst = 32'h8220000;
      15036: inst = 32'h10408000;
      15037: inst = 32'hc4050c7;
      15038: inst = 32'h8220000;
      15039: inst = 32'h10408000;
      15040: inst = 32'hc4050c8;
      15041: inst = 32'h8220000;
      15042: inst = 32'h10408000;
      15043: inst = 32'hc4050c9;
      15044: inst = 32'h8220000;
      15045: inst = 32'h10408000;
      15046: inst = 32'hc4050cb;
      15047: inst = 32'h8220000;
      15048: inst = 32'h10408000;
      15049: inst = 32'hc4050cc;
      15050: inst = 32'h8220000;
      15051: inst = 32'h10408000;
      15052: inst = 32'hc4050cd;
      15053: inst = 32'h8220000;
      15054: inst = 32'h10408000;
      15055: inst = 32'hc4050ce;
      15056: inst = 32'h8220000;
      15057: inst = 32'h10408000;
      15058: inst = 32'hc4050cf;
      15059: inst = 32'h8220000;
      15060: inst = 32'h10408000;
      15061: inst = 32'hc4050d0;
      15062: inst = 32'h8220000;
      15063: inst = 32'h10408000;
      15064: inst = 32'hc4050d1;
      15065: inst = 32'h8220000;
      15066: inst = 32'h10408000;
      15067: inst = 32'hc4050d2;
      15068: inst = 32'h8220000;
      15069: inst = 32'h10408000;
      15070: inst = 32'hc4050d3;
      15071: inst = 32'h8220000;
      15072: inst = 32'h10408000;
      15073: inst = 32'hc405121;
      15074: inst = 32'h8220000;
      15075: inst = 32'h10408000;
      15076: inst = 32'hc405122;
      15077: inst = 32'h8220000;
      15078: inst = 32'h10408000;
      15079: inst = 32'hc405123;
      15080: inst = 32'h8220000;
      15081: inst = 32'h10408000;
      15082: inst = 32'hc405124;
      15083: inst = 32'h8220000;
      15084: inst = 32'h10408000;
      15085: inst = 32'hc405125;
      15086: inst = 32'h8220000;
      15087: inst = 32'h10408000;
      15088: inst = 32'hc405126;
      15089: inst = 32'h8220000;
      15090: inst = 32'h10408000;
      15091: inst = 32'hc405127;
      15092: inst = 32'h8220000;
      15093: inst = 32'h10408000;
      15094: inst = 32'hc405128;
      15095: inst = 32'h8220000;
      15096: inst = 32'h10408000;
      15097: inst = 32'hc405129;
      15098: inst = 32'h8220000;
      15099: inst = 32'h10408000;
      15100: inst = 32'hc40512b;
      15101: inst = 32'h8220000;
      15102: inst = 32'h10408000;
      15103: inst = 32'hc40512c;
      15104: inst = 32'h8220000;
      15105: inst = 32'h10408000;
      15106: inst = 32'hc40512d;
      15107: inst = 32'h8220000;
      15108: inst = 32'h10408000;
      15109: inst = 32'hc40512e;
      15110: inst = 32'h8220000;
      15111: inst = 32'h10408000;
      15112: inst = 32'hc40512f;
      15113: inst = 32'h8220000;
      15114: inst = 32'h10408000;
      15115: inst = 32'hc405130;
      15116: inst = 32'h8220000;
      15117: inst = 32'h10408000;
      15118: inst = 32'hc405131;
      15119: inst = 32'h8220000;
      15120: inst = 32'h10408000;
      15121: inst = 32'hc405132;
      15122: inst = 32'h8220000;
      15123: inst = 32'h10408000;
      15124: inst = 32'hc405133;
      15125: inst = 32'h8220000;
      15126: inst = 32'h10408000;
      15127: inst = 32'hc405181;
      15128: inst = 32'h8220000;
      15129: inst = 32'h10408000;
      15130: inst = 32'hc405182;
      15131: inst = 32'h8220000;
      15132: inst = 32'h10408000;
      15133: inst = 32'hc405183;
      15134: inst = 32'h8220000;
      15135: inst = 32'h10408000;
      15136: inst = 32'hc405184;
      15137: inst = 32'h8220000;
      15138: inst = 32'h10408000;
      15139: inst = 32'hc405185;
      15140: inst = 32'h8220000;
      15141: inst = 32'h10408000;
      15142: inst = 32'hc405186;
      15143: inst = 32'h8220000;
      15144: inst = 32'h10408000;
      15145: inst = 32'hc405187;
      15146: inst = 32'h8220000;
      15147: inst = 32'h10408000;
      15148: inst = 32'hc405188;
      15149: inst = 32'h8220000;
      15150: inst = 32'h10408000;
      15151: inst = 32'hc405189;
      15152: inst = 32'h8220000;
      15153: inst = 32'h10408000;
      15154: inst = 32'hc40518b;
      15155: inst = 32'h8220000;
      15156: inst = 32'h10408000;
      15157: inst = 32'hc40518c;
      15158: inst = 32'h8220000;
      15159: inst = 32'h10408000;
      15160: inst = 32'hc40518d;
      15161: inst = 32'h8220000;
      15162: inst = 32'h10408000;
      15163: inst = 32'hc40518e;
      15164: inst = 32'h8220000;
      15165: inst = 32'h10408000;
      15166: inst = 32'hc40518f;
      15167: inst = 32'h8220000;
      15168: inst = 32'h10408000;
      15169: inst = 32'hc405190;
      15170: inst = 32'h8220000;
      15171: inst = 32'h10408000;
      15172: inst = 32'hc405191;
      15173: inst = 32'h8220000;
      15174: inst = 32'h10408000;
      15175: inst = 32'hc405192;
      15176: inst = 32'h8220000;
      15177: inst = 32'h10408000;
      15178: inst = 32'hc405193;
      15179: inst = 32'h8220000;
      15180: inst = 32'h10408000;
      15181: inst = 32'hc4051e1;
      15182: inst = 32'h8220000;
      15183: inst = 32'h10408000;
      15184: inst = 32'hc4051e2;
      15185: inst = 32'h8220000;
      15186: inst = 32'h10408000;
      15187: inst = 32'hc4051e3;
      15188: inst = 32'h8220000;
      15189: inst = 32'h10408000;
      15190: inst = 32'hc4051e4;
      15191: inst = 32'h8220000;
      15192: inst = 32'h10408000;
      15193: inst = 32'hc4051e5;
      15194: inst = 32'h8220000;
      15195: inst = 32'h10408000;
      15196: inst = 32'hc4051e6;
      15197: inst = 32'h8220000;
      15198: inst = 32'h10408000;
      15199: inst = 32'hc4051e7;
      15200: inst = 32'h8220000;
      15201: inst = 32'h10408000;
      15202: inst = 32'hc4051e8;
      15203: inst = 32'h8220000;
      15204: inst = 32'h10408000;
      15205: inst = 32'hc4051e9;
      15206: inst = 32'h8220000;
      15207: inst = 32'h10408000;
      15208: inst = 32'hc4051eb;
      15209: inst = 32'h8220000;
      15210: inst = 32'h10408000;
      15211: inst = 32'hc4051ec;
      15212: inst = 32'h8220000;
      15213: inst = 32'h10408000;
      15214: inst = 32'hc4051ed;
      15215: inst = 32'h8220000;
      15216: inst = 32'h10408000;
      15217: inst = 32'hc4051ee;
      15218: inst = 32'h8220000;
      15219: inst = 32'h10408000;
      15220: inst = 32'hc4051ef;
      15221: inst = 32'h8220000;
      15222: inst = 32'h10408000;
      15223: inst = 32'hc4051f0;
      15224: inst = 32'h8220000;
      15225: inst = 32'h10408000;
      15226: inst = 32'hc4051f1;
      15227: inst = 32'h8220000;
      15228: inst = 32'h10408000;
      15229: inst = 32'hc4051f2;
      15230: inst = 32'h8220000;
      15231: inst = 32'h10408000;
      15232: inst = 32'hc4051f3;
      15233: inst = 32'h8220000;
      15234: inst = 32'h10408000;
      15235: inst = 32'hc405241;
      15236: inst = 32'h8220000;
      15237: inst = 32'h10408000;
      15238: inst = 32'hc405242;
      15239: inst = 32'h8220000;
      15240: inst = 32'h10408000;
      15241: inst = 32'hc405243;
      15242: inst = 32'h8220000;
      15243: inst = 32'h10408000;
      15244: inst = 32'hc405244;
      15245: inst = 32'h8220000;
      15246: inst = 32'h10408000;
      15247: inst = 32'hc405245;
      15248: inst = 32'h8220000;
      15249: inst = 32'h10408000;
      15250: inst = 32'hc405246;
      15251: inst = 32'h8220000;
      15252: inst = 32'h10408000;
      15253: inst = 32'hc405247;
      15254: inst = 32'h8220000;
      15255: inst = 32'h10408000;
      15256: inst = 32'hc405248;
      15257: inst = 32'h8220000;
      15258: inst = 32'h10408000;
      15259: inst = 32'hc405249;
      15260: inst = 32'h8220000;
      15261: inst = 32'h10408000;
      15262: inst = 32'hc40524b;
      15263: inst = 32'h8220000;
      15264: inst = 32'h10408000;
      15265: inst = 32'hc40524c;
      15266: inst = 32'h8220000;
      15267: inst = 32'h10408000;
      15268: inst = 32'hc40524d;
      15269: inst = 32'h8220000;
      15270: inst = 32'h10408000;
      15271: inst = 32'hc40524e;
      15272: inst = 32'h8220000;
      15273: inst = 32'h10408000;
      15274: inst = 32'hc40524f;
      15275: inst = 32'h8220000;
      15276: inst = 32'h10408000;
      15277: inst = 32'hc405250;
      15278: inst = 32'h8220000;
      15279: inst = 32'h10408000;
      15280: inst = 32'hc405251;
      15281: inst = 32'h8220000;
      15282: inst = 32'h10408000;
      15283: inst = 32'hc405252;
      15284: inst = 32'h8220000;
      15285: inst = 32'h10408000;
      15286: inst = 32'hc405253;
      15287: inst = 32'h8220000;
      15288: inst = 32'hc20bd73;
      15289: inst = 32'h10408000;
      15290: inst = 32'hc404e9f;
      15291: inst = 32'h8220000;
      15292: inst = 32'h10408000;
      15293: inst = 32'hc404ec0;
      15294: inst = 32'h8220000;
      15295: inst = 32'hc205aed;
      15296: inst = 32'h10408000;
      15297: inst = 32'hc404ea0;
      15298: inst = 32'h8220000;
      15299: inst = 32'h10408000;
      15300: inst = 32'hc404ea1;
      15301: inst = 32'h8220000;
      15302: inst = 32'h10408000;
      15303: inst = 32'hc404ea2;
      15304: inst = 32'h8220000;
      15305: inst = 32'h10408000;
      15306: inst = 32'hc404ea3;
      15307: inst = 32'h8220000;
      15308: inst = 32'h10408000;
      15309: inst = 32'hc404ea4;
      15310: inst = 32'h8220000;
      15311: inst = 32'h10408000;
      15312: inst = 32'hc404ebb;
      15313: inst = 32'h8220000;
      15314: inst = 32'h10408000;
      15315: inst = 32'hc404ebc;
      15316: inst = 32'h8220000;
      15317: inst = 32'h10408000;
      15318: inst = 32'hc404ebd;
      15319: inst = 32'h8220000;
      15320: inst = 32'h10408000;
      15321: inst = 32'hc404ebe;
      15322: inst = 32'h8220000;
      15323: inst = 32'h10408000;
      15324: inst = 32'hc404ebf;
      15325: inst = 32'h8220000;
      15326: inst = 32'h10408000;
      15327: inst = 32'hc404f00;
      15328: inst = 32'h8220000;
      15329: inst = 32'h10408000;
      15330: inst = 32'hc404f01;
      15331: inst = 32'h8220000;
      15332: inst = 32'h10408000;
      15333: inst = 32'hc404f02;
      15334: inst = 32'h8220000;
      15335: inst = 32'h10408000;
      15336: inst = 32'hc404f03;
      15337: inst = 32'h8220000;
      15338: inst = 32'h10408000;
      15339: inst = 32'hc404f04;
      15340: inst = 32'h8220000;
      15341: inst = 32'h10408000;
      15342: inst = 32'hc404f05;
      15343: inst = 32'h8220000;
      15344: inst = 32'h10408000;
      15345: inst = 32'hc404f1a;
      15346: inst = 32'h8220000;
      15347: inst = 32'h10408000;
      15348: inst = 32'hc404f1b;
      15349: inst = 32'h8220000;
      15350: inst = 32'h10408000;
      15351: inst = 32'hc404f1c;
      15352: inst = 32'h8220000;
      15353: inst = 32'h10408000;
      15354: inst = 32'hc404f1d;
      15355: inst = 32'h8220000;
      15356: inst = 32'h10408000;
      15357: inst = 32'hc404f1e;
      15358: inst = 32'h8220000;
      15359: inst = 32'h10408000;
      15360: inst = 32'hc404f1f;
      15361: inst = 32'h8220000;
      15362: inst = 32'h10408000;
      15363: inst = 32'hc404f60;
      15364: inst = 32'h8220000;
      15365: inst = 32'h10408000;
      15366: inst = 32'hc404f61;
      15367: inst = 32'h8220000;
      15368: inst = 32'h10408000;
      15369: inst = 32'hc404f62;
      15370: inst = 32'h8220000;
      15371: inst = 32'h10408000;
      15372: inst = 32'hc404f63;
      15373: inst = 32'h8220000;
      15374: inst = 32'h10408000;
      15375: inst = 32'hc404f64;
      15376: inst = 32'h8220000;
      15377: inst = 32'h10408000;
      15378: inst = 32'hc404f65;
      15379: inst = 32'h8220000;
      15380: inst = 32'h10408000;
      15381: inst = 32'hc404f66;
      15382: inst = 32'h8220000;
      15383: inst = 32'h10408000;
      15384: inst = 32'hc404f67;
      15385: inst = 32'h8220000;
      15386: inst = 32'h10408000;
      15387: inst = 32'hc404f78;
      15388: inst = 32'h8220000;
      15389: inst = 32'h10408000;
      15390: inst = 32'hc404f79;
      15391: inst = 32'h8220000;
      15392: inst = 32'h10408000;
      15393: inst = 32'hc404f7a;
      15394: inst = 32'h8220000;
      15395: inst = 32'h10408000;
      15396: inst = 32'hc404f7b;
      15397: inst = 32'h8220000;
      15398: inst = 32'h10408000;
      15399: inst = 32'hc404f7c;
      15400: inst = 32'h8220000;
      15401: inst = 32'h10408000;
      15402: inst = 32'hc404f7d;
      15403: inst = 32'h8220000;
      15404: inst = 32'h10408000;
      15405: inst = 32'hc404f7e;
      15406: inst = 32'h8220000;
      15407: inst = 32'h10408000;
      15408: inst = 32'hc404f7f;
      15409: inst = 32'h8220000;
      15410: inst = 32'h10408000;
      15411: inst = 32'hc404fc0;
      15412: inst = 32'h8220000;
      15413: inst = 32'h10408000;
      15414: inst = 32'hc404fc1;
      15415: inst = 32'h8220000;
      15416: inst = 32'h10408000;
      15417: inst = 32'hc404fc2;
      15418: inst = 32'h8220000;
      15419: inst = 32'h10408000;
      15420: inst = 32'hc404fc3;
      15421: inst = 32'h8220000;
      15422: inst = 32'h10408000;
      15423: inst = 32'hc404fc4;
      15424: inst = 32'h8220000;
      15425: inst = 32'h10408000;
      15426: inst = 32'hc404fc6;
      15427: inst = 32'h8220000;
      15428: inst = 32'h10408000;
      15429: inst = 32'hc404fc7;
      15430: inst = 32'h8220000;
      15431: inst = 32'h10408000;
      15432: inst = 32'hc404fd8;
      15433: inst = 32'h8220000;
      15434: inst = 32'h10408000;
      15435: inst = 32'hc404fd9;
      15436: inst = 32'h8220000;
      15437: inst = 32'h10408000;
      15438: inst = 32'hc404fdb;
      15439: inst = 32'h8220000;
      15440: inst = 32'h10408000;
      15441: inst = 32'hc404fdc;
      15442: inst = 32'h8220000;
      15443: inst = 32'h10408000;
      15444: inst = 32'hc404fdd;
      15445: inst = 32'h8220000;
      15446: inst = 32'h10408000;
      15447: inst = 32'hc404fde;
      15448: inst = 32'h8220000;
      15449: inst = 32'h10408000;
      15450: inst = 32'hc404fdf;
      15451: inst = 32'h8220000;
      15452: inst = 32'h10408000;
      15453: inst = 32'hc405020;
      15454: inst = 32'h8220000;
      15455: inst = 32'h10408000;
      15456: inst = 32'hc405021;
      15457: inst = 32'h8220000;
      15458: inst = 32'h10408000;
      15459: inst = 32'hc405022;
      15460: inst = 32'h8220000;
      15461: inst = 32'h10408000;
      15462: inst = 32'hc405023;
      15463: inst = 32'h8220000;
      15464: inst = 32'h10408000;
      15465: inst = 32'hc405026;
      15466: inst = 32'h8220000;
      15467: inst = 32'h10408000;
      15468: inst = 32'hc405027;
      15469: inst = 32'h8220000;
      15470: inst = 32'h10408000;
      15471: inst = 32'hc405038;
      15472: inst = 32'h8220000;
      15473: inst = 32'h10408000;
      15474: inst = 32'hc405039;
      15475: inst = 32'h8220000;
      15476: inst = 32'h10408000;
      15477: inst = 32'hc40503c;
      15478: inst = 32'h8220000;
      15479: inst = 32'h10408000;
      15480: inst = 32'hc40503d;
      15481: inst = 32'h8220000;
      15482: inst = 32'h10408000;
      15483: inst = 32'hc40503e;
      15484: inst = 32'h8220000;
      15485: inst = 32'h10408000;
      15486: inst = 32'hc40503f;
      15487: inst = 32'h8220000;
      15488: inst = 32'h10408000;
      15489: inst = 32'hc40507f;
      15490: inst = 32'h8220000;
      15491: inst = 32'h10408000;
      15492: inst = 32'hc405080;
      15493: inst = 32'h8220000;
      15494: inst = 32'h10408000;
      15495: inst = 32'hc405081;
      15496: inst = 32'h8220000;
      15497: inst = 32'h10408000;
      15498: inst = 32'hc405082;
      15499: inst = 32'h8220000;
      15500: inst = 32'h10408000;
      15501: inst = 32'hc405086;
      15502: inst = 32'h8220000;
      15503: inst = 32'h10408000;
      15504: inst = 32'hc405087;
      15505: inst = 32'h8220000;
      15506: inst = 32'h10408000;
      15507: inst = 32'hc405098;
      15508: inst = 32'h8220000;
      15509: inst = 32'h10408000;
      15510: inst = 32'hc405099;
      15511: inst = 32'h8220000;
      15512: inst = 32'h10408000;
      15513: inst = 32'hc40509d;
      15514: inst = 32'h8220000;
      15515: inst = 32'h10408000;
      15516: inst = 32'hc40509e;
      15517: inst = 32'h8220000;
      15518: inst = 32'h10408000;
      15519: inst = 32'hc40509f;
      15520: inst = 32'h8220000;
      15521: inst = 32'h10408000;
      15522: inst = 32'hc4050a0;
      15523: inst = 32'h8220000;
      15524: inst = 32'h10408000;
      15525: inst = 32'hc4050df;
      15526: inst = 32'h8220000;
      15527: inst = 32'h10408000;
      15528: inst = 32'hc4050e0;
      15529: inst = 32'h8220000;
      15530: inst = 32'h10408000;
      15531: inst = 32'hc4050e1;
      15532: inst = 32'h8220000;
      15533: inst = 32'h10408000;
      15534: inst = 32'hc4050e2;
      15535: inst = 32'h8220000;
      15536: inst = 32'h10408000;
      15537: inst = 32'hc4050e6;
      15538: inst = 32'h8220000;
      15539: inst = 32'h10408000;
      15540: inst = 32'hc4050e7;
      15541: inst = 32'h8220000;
      15542: inst = 32'h10408000;
      15543: inst = 32'hc4050f8;
      15544: inst = 32'h8220000;
      15545: inst = 32'h10408000;
      15546: inst = 32'hc4050f9;
      15547: inst = 32'h8220000;
      15548: inst = 32'h10408000;
      15549: inst = 32'hc4050fd;
      15550: inst = 32'h8220000;
      15551: inst = 32'h10408000;
      15552: inst = 32'hc4050fe;
      15553: inst = 32'h8220000;
      15554: inst = 32'h10408000;
      15555: inst = 32'hc4050ff;
      15556: inst = 32'h8220000;
      15557: inst = 32'h10408000;
      15558: inst = 32'hc405100;
      15559: inst = 32'h8220000;
      15560: inst = 32'h10408000;
      15561: inst = 32'hc40513f;
      15562: inst = 32'h8220000;
      15563: inst = 32'h10408000;
      15564: inst = 32'hc405140;
      15565: inst = 32'h8220000;
      15566: inst = 32'h10408000;
      15567: inst = 32'hc405141;
      15568: inst = 32'h8220000;
      15569: inst = 32'h10408000;
      15570: inst = 32'hc405146;
      15571: inst = 32'h8220000;
      15572: inst = 32'h10408000;
      15573: inst = 32'hc405147;
      15574: inst = 32'h8220000;
      15575: inst = 32'h10408000;
      15576: inst = 32'hc405158;
      15577: inst = 32'h8220000;
      15578: inst = 32'h10408000;
      15579: inst = 32'hc405159;
      15580: inst = 32'h8220000;
      15581: inst = 32'h10408000;
      15582: inst = 32'hc40515e;
      15583: inst = 32'h8220000;
      15584: inst = 32'h10408000;
      15585: inst = 32'hc40515f;
      15586: inst = 32'h8220000;
      15587: inst = 32'h10408000;
      15588: inst = 32'hc405160;
      15589: inst = 32'h8220000;
      15590: inst = 32'h10408000;
      15591: inst = 32'hc40519f;
      15592: inst = 32'h8220000;
      15593: inst = 32'h10408000;
      15594: inst = 32'hc4051a0;
      15595: inst = 32'h8220000;
      15596: inst = 32'h10408000;
      15597: inst = 32'hc4051a6;
      15598: inst = 32'h8220000;
      15599: inst = 32'h10408000;
      15600: inst = 32'hc4051a7;
      15601: inst = 32'h8220000;
      15602: inst = 32'h10408000;
      15603: inst = 32'hc4051b8;
      15604: inst = 32'h8220000;
      15605: inst = 32'h10408000;
      15606: inst = 32'hc4051b9;
      15607: inst = 32'h8220000;
      15608: inst = 32'h10408000;
      15609: inst = 32'hc4051bf;
      15610: inst = 32'h8220000;
      15611: inst = 32'h10408000;
      15612: inst = 32'hc4051c0;
      15613: inst = 32'h8220000;
      15614: inst = 32'h10408000;
      15615: inst = 32'hc4051ff;
      15616: inst = 32'h8220000;
      15617: inst = 32'h10408000;
      15618: inst = 32'hc405200;
      15619: inst = 32'h8220000;
      15620: inst = 32'h10408000;
      15621: inst = 32'hc405206;
      15622: inst = 32'h8220000;
      15623: inst = 32'h10408000;
      15624: inst = 32'hc405207;
      15625: inst = 32'h8220000;
      15626: inst = 32'h10408000;
      15627: inst = 32'hc405218;
      15628: inst = 32'h8220000;
      15629: inst = 32'h10408000;
      15630: inst = 32'hc405219;
      15631: inst = 32'h8220000;
      15632: inst = 32'h10408000;
      15633: inst = 32'hc40521f;
      15634: inst = 32'h8220000;
      15635: inst = 32'h10408000;
      15636: inst = 32'hc405220;
      15637: inst = 32'h8220000;
      15638: inst = 32'h10408000;
      15639: inst = 32'hc40525f;
      15640: inst = 32'h8220000;
      15641: inst = 32'h10408000;
      15642: inst = 32'hc405260;
      15643: inst = 32'h8220000;
      15644: inst = 32'h10408000;
      15645: inst = 32'hc405266;
      15646: inst = 32'h8220000;
      15647: inst = 32'h10408000;
      15648: inst = 32'hc405267;
      15649: inst = 32'h8220000;
      15650: inst = 32'h10408000;
      15651: inst = 32'hc405278;
      15652: inst = 32'h8220000;
      15653: inst = 32'h10408000;
      15654: inst = 32'hc405279;
      15655: inst = 32'h8220000;
      15656: inst = 32'h10408000;
      15657: inst = 32'hc40527f;
      15658: inst = 32'h8220000;
      15659: inst = 32'h10408000;
      15660: inst = 32'hc405280;
      15661: inst = 32'h8220000;
      15662: inst = 32'h10408000;
      15663: inst = 32'hc4052bf;
      15664: inst = 32'h8220000;
      15665: inst = 32'h10408000;
      15666: inst = 32'hc4052c0;
      15667: inst = 32'h8220000;
      15668: inst = 32'h10408000;
      15669: inst = 32'hc4052c6;
      15670: inst = 32'h8220000;
      15671: inst = 32'h10408000;
      15672: inst = 32'hc4052c7;
      15673: inst = 32'h8220000;
      15674: inst = 32'h10408000;
      15675: inst = 32'hc4052d8;
      15676: inst = 32'h8220000;
      15677: inst = 32'h10408000;
      15678: inst = 32'hc4052d9;
      15679: inst = 32'h8220000;
      15680: inst = 32'h10408000;
      15681: inst = 32'hc4052df;
      15682: inst = 32'h8220000;
      15683: inst = 32'h10408000;
      15684: inst = 32'hc4052e0;
      15685: inst = 32'h8220000;
      15686: inst = 32'hc207bae;
      15687: inst = 32'h10408000;
      15688: inst = 32'hc404ea5;
      15689: inst = 32'h8220000;
      15690: inst = 32'h10408000;
      15691: inst = 32'hc404eba;
      15692: inst = 32'h8220000;
      15693: inst = 32'hc20c5b4;
      15694: inst = 32'h10408000;
      15695: inst = 32'hc404ea6;
      15696: inst = 32'h8220000;
      15697: inst = 32'h10408000;
      15698: inst = 32'hc404eb9;
      15699: inst = 32'h8220000;
      15700: inst = 32'hc20d5f4;
      15701: inst = 32'h10408000;
      15702: inst = 32'hc404ea7;
      15703: inst = 32'h8220000;
      15704: inst = 32'h10408000;
      15705: inst = 32'hc404eb8;
      15706: inst = 32'h8220000;
      15707: inst = 32'hc20a4b1;
      15708: inst = 32'h10408000;
      15709: inst = 32'hc404eff;
      15710: inst = 32'h8220000;
      15711: inst = 32'h10408000;
      15712: inst = 32'hc404f20;
      15713: inst = 32'h8220000;
      15714: inst = 32'h10408000;
      15715: inst = 32'hc404fbf;
      15716: inst = 32'h8220000;
      15717: inst = 32'h10408000;
      15718: inst = 32'hc404fe0;
      15719: inst = 32'h8220000;
      15720: inst = 32'hc2062ed;
      15721: inst = 32'h10408000;
      15722: inst = 32'hc404f06;
      15723: inst = 32'h8220000;
      15724: inst = 32'h10408000;
      15725: inst = 32'hc404f19;
      15726: inst = 32'h8220000;
      15727: inst = 32'hc209450;
      15728: inst = 32'h10408000;
      15729: inst = 32'hc404f07;
      15730: inst = 32'h8220000;
      15731: inst = 32'h10408000;
      15732: inst = 32'hc404f18;
      15733: inst = 32'h8220000;
      15734: inst = 32'h10408000;
      15735: inst = 32'hc405209;
      15736: inst = 32'h8220000;
      15737: inst = 32'h10408000;
      15738: inst = 32'hc405216;
      15739: inst = 32'h8220000;
      15740: inst = 32'hc20a4d1;
      15741: inst = 32'h10408000;
      15742: inst = 32'hc404f5f;
      15743: inst = 32'h8220000;
      15744: inst = 32'h10408000;
      15745: inst = 32'hc404f80;
      15746: inst = 32'h8220000;
      15747: inst = 32'hc204a49;
      15748: inst = 32'h10408000;
      15749: inst = 32'hc404fa8;
      15750: inst = 32'h8220000;
      15751: inst = 32'h10408000;
      15752: inst = 32'hc404fac;
      15753: inst = 32'h8220000;
      15754: inst = 32'h10408000;
      15755: inst = 32'hc405008;
      15756: inst = 32'h8220000;
      15757: inst = 32'h10408000;
      15758: inst = 32'hc40500c;
      15759: inst = 32'h8220000;
      15760: inst = 32'hc205acb;
      15761: inst = 32'h10408000;
      15762: inst = 32'hc404fc5;
      15763: inst = 32'h8220000;
      15764: inst = 32'h10408000;
      15765: inst = 32'hc404fda;
      15766: inst = 32'h8220000;
      15767: inst = 32'h10408000;
      15768: inst = 32'hc405336;
      15769: inst = 32'h8220000;
      15770: inst = 32'h10408000;
      15771: inst = 32'hc405380;
      15772: inst = 32'h8220000;
      15773: inst = 32'h10408000;
      15774: inst = 32'hc40539f;
      15775: inst = 32'h8220000;
      15776: inst = 32'h10408000;
      15777: inst = 32'hc4053dd;
      15778: inst = 32'h8220000;
      15779: inst = 32'h10408000;
      15780: inst = 32'hc405402;
      15781: inst = 32'h8220000;
      15782: inst = 32'hc20630d;
      15783: inst = 32'h10408000;
      15784: inst = 32'hc40501f;
      15785: inst = 32'h8220000;
      15786: inst = 32'h10408000;
      15787: inst = 32'hc405040;
      15788: inst = 32'h8220000;
      15789: inst = 32'hc205aec;
      15790: inst = 32'h10408000;
      15791: inst = 32'hc405024;
      15792: inst = 32'h8220000;
      15793: inst = 32'h10408000;
      15794: inst = 32'hc40503b;
      15795: inst = 32'h8220000;
      15796: inst = 32'h10408000;
      15797: inst = 32'hc405083;
      15798: inst = 32'h8220000;
      15799: inst = 32'h10408000;
      15800: inst = 32'hc40509c;
      15801: inst = 32'h8220000;
      15802: inst = 32'h10408000;
      15803: inst = 32'hc4051a1;
      15804: inst = 32'h8220000;
      15805: inst = 32'h10408000;
      15806: inst = 32'hc4051be;
      15807: inst = 32'h8220000;
      15808: inst = 32'h10408000;
      15809: inst = 32'hc405329;
      15810: inst = 32'h8220000;
      15811: inst = 32'h10408000;
      15812: inst = 32'hc405568;
      15813: inst = 32'h8220000;
      15814: inst = 32'h10408000;
      15815: inst = 32'hc405577;
      15816: inst = 32'h8220000;
      15817: inst = 32'h10408000;
      15818: inst = 32'hc4057a7;
      15819: inst = 32'h8220000;
      15820: inst = 32'h10408000;
      15821: inst = 32'hc4057b8;
      15822: inst = 32'h8220000;
      15823: inst = 32'hc205269;
      15824: inst = 32'h10408000;
      15825: inst = 32'hc405025;
      15826: inst = 32'h8220000;
      15827: inst = 32'h10408000;
      15828: inst = 32'hc40503a;
      15829: inst = 32'h8220000;
      15830: inst = 32'h10408000;
      15831: inst = 32'hc40537e;
      15832: inst = 32'h8220000;
      15833: inst = 32'h10408000;
      15834: inst = 32'hc4053a1;
      15835: inst = 32'h8220000;
      15836: inst = 32'h10408000;
      15837: inst = 32'hc40549c;
      15838: inst = 32'h8220000;
      15839: inst = 32'h10408000;
      15840: inst = 32'hc4054c3;
      15841: inst = 32'h8220000;
      15842: inst = 32'hc20528a;
      15843: inst = 32'h10408000;
      15844: inst = 32'hc405084;
      15845: inst = 32'h8220000;
      15846: inst = 32'h10408000;
      15847: inst = 32'hc40509b;
      15848: inst = 32'h8220000;
      15849: inst = 32'h10408000;
      15850: inst = 32'hc4050e3;
      15851: inst = 32'h8220000;
      15852: inst = 32'h10408000;
      15853: inst = 32'hc4050fc;
      15854: inst = 32'h8220000;
      15855: inst = 32'h10408000;
      15856: inst = 32'hc4052c5;
      15857: inst = 32'h8220000;
      15858: inst = 32'h10408000;
      15859: inst = 32'hc4052da;
      15860: inst = 32'h8220000;
      15861: inst = 32'h10408000;
      15862: inst = 32'hc4053e9;
      15863: inst = 32'h8220000;
      15864: inst = 32'h10408000;
      15865: inst = 32'hc4053f6;
      15866: inst = 32'h8220000;
      15867: inst = 32'h10408000;
      15868: inst = 32'hc405449;
      15869: inst = 32'h8220000;
      15870: inst = 32'h10408000;
      15871: inst = 32'hc405456;
      15872: inst = 32'h8220000;
      15873: inst = 32'h10408000;
      15874: inst = 32'hc4054a9;
      15875: inst = 32'h8220000;
      15876: inst = 32'h10408000;
      15877: inst = 32'hc4054b6;
      15878: inst = 32'h8220000;
      15879: inst = 32'h10408000;
      15880: inst = 32'hc405509;
      15881: inst = 32'h8220000;
      15882: inst = 32'h10408000;
      15883: inst = 32'hc405516;
      15884: inst = 32'h8220000;
      15885: inst = 32'h10408000;
      15886: inst = 32'hc40555e;
      15887: inst = 32'h8220000;
      15888: inst = 32'h10408000;
      15889: inst = 32'hc405569;
      15890: inst = 32'h8220000;
      15891: inst = 32'h10408000;
      15892: inst = 32'hc405576;
      15893: inst = 32'h8220000;
      15894: inst = 32'h10408000;
      15895: inst = 32'hc405581;
      15896: inst = 32'h8220000;
      15897: inst = 32'h10408000;
      15898: inst = 32'hc4055c9;
      15899: inst = 32'h8220000;
      15900: inst = 32'h10408000;
      15901: inst = 32'hc4055d6;
      15902: inst = 32'h8220000;
      15903: inst = 32'h10408000;
      15904: inst = 32'hc405628;
      15905: inst = 32'h8220000;
      15906: inst = 32'h10408000;
      15907: inst = 32'hc405629;
      15908: inst = 32'h8220000;
      15909: inst = 32'h10408000;
      15910: inst = 32'hc405636;
      15911: inst = 32'h8220000;
      15912: inst = 32'h10408000;
      15913: inst = 32'hc405637;
      15914: inst = 32'h8220000;
      15915: inst = 32'h10408000;
      15916: inst = 32'hc40567d;
      15917: inst = 32'h8220000;
      15918: inst = 32'h10408000;
      15919: inst = 32'hc405688;
      15920: inst = 32'h8220000;
      15921: inst = 32'h10408000;
      15922: inst = 32'hc405689;
      15923: inst = 32'h8220000;
      15924: inst = 32'h10408000;
      15925: inst = 32'hc405696;
      15926: inst = 32'h8220000;
      15927: inst = 32'h10408000;
      15928: inst = 32'hc405697;
      15929: inst = 32'h8220000;
      15930: inst = 32'h10408000;
      15931: inst = 32'hc4056a2;
      15932: inst = 32'h8220000;
      15933: inst = 32'h10408000;
      15934: inst = 32'hc4056e8;
      15935: inst = 32'h8220000;
      15936: inst = 32'h10408000;
      15937: inst = 32'hc4056e9;
      15938: inst = 32'h8220000;
      15939: inst = 32'h10408000;
      15940: inst = 32'hc4056f6;
      15941: inst = 32'h8220000;
      15942: inst = 32'h10408000;
      15943: inst = 32'hc4056f7;
      15944: inst = 32'h8220000;
      15945: inst = 32'h10408000;
      15946: inst = 32'hc405748;
      15947: inst = 32'h8220000;
      15948: inst = 32'h10408000;
      15949: inst = 32'hc405749;
      15950: inst = 32'h8220000;
      15951: inst = 32'h10408000;
      15952: inst = 32'hc405756;
      15953: inst = 32'h8220000;
      15954: inst = 32'h10408000;
      15955: inst = 32'hc405757;
      15956: inst = 32'h8220000;
      15957: inst = 32'h10408000;
      15958: inst = 32'hc4057a8;
      15959: inst = 32'h8220000;
      15960: inst = 32'h10408000;
      15961: inst = 32'hc4057a9;
      15962: inst = 32'h8220000;
      15963: inst = 32'h10408000;
      15964: inst = 32'hc4057b6;
      15965: inst = 32'h8220000;
      15966: inst = 32'h10408000;
      15967: inst = 32'hc4057b7;
      15968: inst = 32'h8220000;
      15969: inst = 32'hc205aab;
      15970: inst = 32'h10408000;
      15971: inst = 32'hc405142;
      15972: inst = 32'h8220000;
      15973: inst = 32'h10408000;
      15974: inst = 32'hc40515d;
      15975: inst = 32'h8220000;
      15976: inst = 32'hc20cdd4;
      15977: inst = 32'h10408000;
      15978: inst = 32'hc40519e;
      15979: inst = 32'h8220000;
      15980: inst = 32'h10408000;
      15981: inst = 32'hc4051c1;
      15982: inst = 32'h8220000;
      15983: inst = 32'hc209471;
      15984: inst = 32'h10408000;
      15985: inst = 32'hc4051b6;
      15986: inst = 32'h8220000;
      15987: inst = 32'hc20de55;
      15988: inst = 32'h10408000;
      15989: inst = 32'hc4051fd;
      15990: inst = 32'h8220000;
      15991: inst = 32'h10408000;
      15992: inst = 32'hc405222;
      15993: inst = 32'h8220000;
      15994: inst = 32'hc209492;
      15995: inst = 32'h10408000;
      15996: inst = 32'hc4051fe;
      15997: inst = 32'h8220000;
      15998: inst = 32'h10408000;
      15999: inst = 32'hc405221;
      16000: inst = 32'h8220000;
      16001: inst = 32'hc205acc;
      16002: inst = 32'h10408000;
      16003: inst = 32'hc405201;
      16004: inst = 32'h8220000;
      16005: inst = 32'h10408000;
      16006: inst = 32'hc40521e;
      16007: inst = 32'h8220000;
      16008: inst = 32'h10408000;
      16009: inst = 32'hc405261;
      16010: inst = 32'h8220000;
      16011: inst = 32'h10408000;
      16012: inst = 32'hc40527e;
      16013: inst = 32'h8220000;
      16014: inst = 32'h10408000;
      16015: inst = 32'hc4052c1;
      16016: inst = 32'h8220000;
      16017: inst = 32'h10408000;
      16018: inst = 32'hc4052de;
      16019: inst = 32'h8220000;
      16020: inst = 32'hc20e696;
      16021: inst = 32'h10408000;
      16022: inst = 32'hc40525c;
      16023: inst = 32'h8220000;
      16024: inst = 32'h10408000;
      16025: inst = 32'hc405283;
      16026: inst = 32'h8220000;
      16027: inst = 32'hc209cb2;
      16028: inst = 32'h10408000;
      16029: inst = 32'hc40525d;
      16030: inst = 32'h8220000;
      16031: inst = 32'h10408000;
      16032: inst = 32'hc405282;
      16033: inst = 32'h8220000;
      16034: inst = 32'hc208c2f;
      16035: inst = 32'h10408000;
      16036: inst = 32'hc405269;
      16037: inst = 32'h8220000;
      16038: inst = 32'h10408000;
      16039: inst = 32'hc405276;
      16040: inst = 32'h8220000;
      16041: inst = 32'hc20ad33;
      16042: inst = 32'h10408000;
      16043: inst = 32'hc4052bc;
      16044: inst = 32'h8220000;
      16045: inst = 32'h10408000;
      16046: inst = 32'hc4052e3;
      16047: inst = 32'h8220000;
      16048: inst = 32'hc2083ee;
      16049: inst = 32'h10408000;
      16050: inst = 32'hc4052c9;
      16051: inst = 32'h8220000;
      16052: inst = 32'h10408000;
      16053: inst = 32'hc4052d6;
      16054: inst = 32'h8220000;
      16055: inst = 32'hc206b50;
      16056: inst = 32'h10408000;
      16057: inst = 32'hc405300;
      16058: inst = 32'h8220000;
      16059: inst = 32'h10408000;
      16060: inst = 32'hc405301;
      16061: inst = 32'h8220000;
      16062: inst = 32'h10408000;
      16063: inst = 32'hc405302;
      16064: inst = 32'h8220000;
      16065: inst = 32'h10408000;
      16066: inst = 32'hc405303;
      16067: inst = 32'h8220000;
      16068: inst = 32'h10408000;
      16069: inst = 32'hc405304;
      16070: inst = 32'h8220000;
      16071: inst = 32'h10408000;
      16072: inst = 32'hc405305;
      16073: inst = 32'h8220000;
      16074: inst = 32'h10408000;
      16075: inst = 32'hc405306;
      16076: inst = 32'h8220000;
      16077: inst = 32'h10408000;
      16078: inst = 32'hc405307;
      16079: inst = 32'h8220000;
      16080: inst = 32'h10408000;
      16081: inst = 32'hc405308;
      16082: inst = 32'h8220000;
      16083: inst = 32'h10408000;
      16084: inst = 32'hc405309;
      16085: inst = 32'h8220000;
      16086: inst = 32'h10408000;
      16087: inst = 32'hc40530a;
      16088: inst = 32'h8220000;
      16089: inst = 32'h10408000;
      16090: inst = 32'hc40530b;
      16091: inst = 32'h8220000;
      16092: inst = 32'h10408000;
      16093: inst = 32'hc40530c;
      16094: inst = 32'h8220000;
      16095: inst = 32'h10408000;
      16096: inst = 32'hc40530d;
      16097: inst = 32'h8220000;
      16098: inst = 32'h10408000;
      16099: inst = 32'hc40530e;
      16100: inst = 32'h8220000;
      16101: inst = 32'h10408000;
      16102: inst = 32'hc40530f;
      16103: inst = 32'h8220000;
      16104: inst = 32'h10408000;
      16105: inst = 32'hc405310;
      16106: inst = 32'h8220000;
      16107: inst = 32'h10408000;
      16108: inst = 32'hc405311;
      16109: inst = 32'h8220000;
      16110: inst = 32'h10408000;
      16111: inst = 32'hc405312;
      16112: inst = 32'h8220000;
      16113: inst = 32'h10408000;
      16114: inst = 32'hc405313;
      16115: inst = 32'h8220000;
      16116: inst = 32'h10408000;
      16117: inst = 32'hc405314;
      16118: inst = 32'h8220000;
      16119: inst = 32'h10408000;
      16120: inst = 32'hc405315;
      16121: inst = 32'h8220000;
      16122: inst = 32'h10408000;
      16123: inst = 32'hc405316;
      16124: inst = 32'h8220000;
      16125: inst = 32'h10408000;
      16126: inst = 32'hc405317;
      16127: inst = 32'h8220000;
      16128: inst = 32'h10408000;
      16129: inst = 32'hc405318;
      16130: inst = 32'h8220000;
      16131: inst = 32'h10408000;
      16132: inst = 32'hc405319;
      16133: inst = 32'h8220000;
      16134: inst = 32'h10408000;
      16135: inst = 32'hc40531a;
      16136: inst = 32'h8220000;
      16137: inst = 32'h10408000;
      16138: inst = 32'hc40532a;
      16139: inst = 32'h8220000;
      16140: inst = 32'h10408000;
      16141: inst = 32'hc40532b;
      16142: inst = 32'h8220000;
      16143: inst = 32'h10408000;
      16144: inst = 32'hc40532c;
      16145: inst = 32'h8220000;
      16146: inst = 32'h10408000;
      16147: inst = 32'hc40532d;
      16148: inst = 32'h8220000;
      16149: inst = 32'h10408000;
      16150: inst = 32'hc40532e;
      16151: inst = 32'h8220000;
      16152: inst = 32'h10408000;
      16153: inst = 32'hc40532f;
      16154: inst = 32'h8220000;
      16155: inst = 32'h10408000;
      16156: inst = 32'hc405330;
      16157: inst = 32'h8220000;
      16158: inst = 32'h10408000;
      16159: inst = 32'hc405331;
      16160: inst = 32'h8220000;
      16161: inst = 32'h10408000;
      16162: inst = 32'hc405332;
      16163: inst = 32'h8220000;
      16164: inst = 32'h10408000;
      16165: inst = 32'hc405333;
      16166: inst = 32'h8220000;
      16167: inst = 32'h10408000;
      16168: inst = 32'hc405334;
      16169: inst = 32'h8220000;
      16170: inst = 32'h10408000;
      16171: inst = 32'hc405335;
      16172: inst = 32'h8220000;
      16173: inst = 32'h10408000;
      16174: inst = 32'hc405345;
      16175: inst = 32'h8220000;
      16176: inst = 32'h10408000;
      16177: inst = 32'hc405346;
      16178: inst = 32'h8220000;
      16179: inst = 32'h10408000;
      16180: inst = 32'hc405347;
      16181: inst = 32'h8220000;
      16182: inst = 32'h10408000;
      16183: inst = 32'hc405348;
      16184: inst = 32'h8220000;
      16185: inst = 32'h10408000;
      16186: inst = 32'hc405349;
      16187: inst = 32'h8220000;
      16188: inst = 32'h10408000;
      16189: inst = 32'hc40534a;
      16190: inst = 32'h8220000;
      16191: inst = 32'h10408000;
      16192: inst = 32'hc40534b;
      16193: inst = 32'h8220000;
      16194: inst = 32'h10408000;
      16195: inst = 32'hc40534c;
      16196: inst = 32'h8220000;
      16197: inst = 32'h10408000;
      16198: inst = 32'hc40534d;
      16199: inst = 32'h8220000;
      16200: inst = 32'h10408000;
      16201: inst = 32'hc40534e;
      16202: inst = 32'h8220000;
      16203: inst = 32'h10408000;
      16204: inst = 32'hc40534f;
      16205: inst = 32'h8220000;
      16206: inst = 32'h10408000;
      16207: inst = 32'hc405350;
      16208: inst = 32'h8220000;
      16209: inst = 32'h10408000;
      16210: inst = 32'hc405351;
      16211: inst = 32'h8220000;
      16212: inst = 32'h10408000;
      16213: inst = 32'hc405352;
      16214: inst = 32'h8220000;
      16215: inst = 32'h10408000;
      16216: inst = 32'hc405353;
      16217: inst = 32'h8220000;
      16218: inst = 32'h10408000;
      16219: inst = 32'hc405354;
      16220: inst = 32'h8220000;
      16221: inst = 32'h10408000;
      16222: inst = 32'hc405355;
      16223: inst = 32'h8220000;
      16224: inst = 32'h10408000;
      16225: inst = 32'hc405356;
      16226: inst = 32'h8220000;
      16227: inst = 32'h10408000;
      16228: inst = 32'hc405357;
      16229: inst = 32'h8220000;
      16230: inst = 32'h10408000;
      16231: inst = 32'hc405358;
      16232: inst = 32'h8220000;
      16233: inst = 32'h10408000;
      16234: inst = 32'hc405359;
      16235: inst = 32'h8220000;
      16236: inst = 32'h10408000;
      16237: inst = 32'hc40535a;
      16238: inst = 32'h8220000;
      16239: inst = 32'h10408000;
      16240: inst = 32'hc40535b;
      16241: inst = 32'h8220000;
      16242: inst = 32'h10408000;
      16243: inst = 32'hc40535c;
      16244: inst = 32'h8220000;
      16245: inst = 32'h10408000;
      16246: inst = 32'hc40535d;
      16247: inst = 32'h8220000;
      16248: inst = 32'h10408000;
      16249: inst = 32'hc40535e;
      16250: inst = 32'h8220000;
      16251: inst = 32'h10408000;
      16252: inst = 32'hc40535f;
      16253: inst = 32'h8220000;
      16254: inst = 32'h10408000;
      16255: inst = 32'hc405360;
      16256: inst = 32'h8220000;
      16257: inst = 32'h10408000;
      16258: inst = 32'hc405361;
      16259: inst = 32'h8220000;
      16260: inst = 32'h10408000;
      16261: inst = 32'hc405362;
      16262: inst = 32'h8220000;
      16263: inst = 32'h10408000;
      16264: inst = 32'hc405363;
      16265: inst = 32'h8220000;
      16266: inst = 32'h10408000;
      16267: inst = 32'hc405364;
      16268: inst = 32'h8220000;
      16269: inst = 32'h10408000;
      16270: inst = 32'hc405365;
      16271: inst = 32'h8220000;
      16272: inst = 32'h10408000;
      16273: inst = 32'hc405366;
      16274: inst = 32'h8220000;
      16275: inst = 32'h10408000;
      16276: inst = 32'hc405367;
      16277: inst = 32'h8220000;
      16278: inst = 32'h10408000;
      16279: inst = 32'hc405368;
      16280: inst = 32'h8220000;
      16281: inst = 32'h10408000;
      16282: inst = 32'hc405369;
      16283: inst = 32'h8220000;
      16284: inst = 32'h10408000;
      16285: inst = 32'hc40536a;
      16286: inst = 32'h8220000;
      16287: inst = 32'h10408000;
      16288: inst = 32'hc40536b;
      16289: inst = 32'h8220000;
      16290: inst = 32'h10408000;
      16291: inst = 32'hc40536c;
      16292: inst = 32'h8220000;
      16293: inst = 32'h10408000;
      16294: inst = 32'hc40536d;
      16295: inst = 32'h8220000;
      16296: inst = 32'h10408000;
      16297: inst = 32'hc40536e;
      16298: inst = 32'h8220000;
      16299: inst = 32'h10408000;
      16300: inst = 32'hc40536f;
      16301: inst = 32'h8220000;
      16302: inst = 32'h10408000;
      16303: inst = 32'hc405370;
      16304: inst = 32'h8220000;
      16305: inst = 32'h10408000;
      16306: inst = 32'hc405371;
      16307: inst = 32'h8220000;
      16308: inst = 32'h10408000;
      16309: inst = 32'hc405372;
      16310: inst = 32'h8220000;
      16311: inst = 32'h10408000;
      16312: inst = 32'hc405373;
      16313: inst = 32'h8220000;
      16314: inst = 32'h10408000;
      16315: inst = 32'hc405374;
      16316: inst = 32'h8220000;
      16317: inst = 32'h10408000;
      16318: inst = 32'hc405375;
      16319: inst = 32'h8220000;
      16320: inst = 32'h10408000;
      16321: inst = 32'hc405376;
      16322: inst = 32'h8220000;
      16323: inst = 32'h10408000;
      16324: inst = 32'hc405377;
      16325: inst = 32'h8220000;
      16326: inst = 32'h10408000;
      16327: inst = 32'hc405378;
      16328: inst = 32'h8220000;
      16329: inst = 32'h10408000;
      16330: inst = 32'hc405379;
      16331: inst = 32'h8220000;
      16332: inst = 32'h10408000;
      16333: inst = 32'hc40538a;
      16334: inst = 32'h8220000;
      16335: inst = 32'h10408000;
      16336: inst = 32'hc40538b;
      16337: inst = 32'h8220000;
      16338: inst = 32'h10408000;
      16339: inst = 32'hc40538c;
      16340: inst = 32'h8220000;
      16341: inst = 32'h10408000;
      16342: inst = 32'hc40538d;
      16343: inst = 32'h8220000;
      16344: inst = 32'h10408000;
      16345: inst = 32'hc40538e;
      16346: inst = 32'h8220000;
      16347: inst = 32'h10408000;
      16348: inst = 32'hc40538f;
      16349: inst = 32'h8220000;
      16350: inst = 32'h10408000;
      16351: inst = 32'hc405390;
      16352: inst = 32'h8220000;
      16353: inst = 32'h10408000;
      16354: inst = 32'hc405391;
      16355: inst = 32'h8220000;
      16356: inst = 32'h10408000;
      16357: inst = 32'hc405392;
      16358: inst = 32'h8220000;
      16359: inst = 32'h10408000;
      16360: inst = 32'hc405393;
      16361: inst = 32'h8220000;
      16362: inst = 32'h10408000;
      16363: inst = 32'hc405394;
      16364: inst = 32'h8220000;
      16365: inst = 32'h10408000;
      16366: inst = 32'hc405395;
      16367: inst = 32'h8220000;
      16368: inst = 32'h10408000;
      16369: inst = 32'hc4053a6;
      16370: inst = 32'h8220000;
      16371: inst = 32'h10408000;
      16372: inst = 32'hc4053a7;
      16373: inst = 32'h8220000;
      16374: inst = 32'h10408000;
      16375: inst = 32'hc4053a8;
      16376: inst = 32'h8220000;
      16377: inst = 32'h10408000;
      16378: inst = 32'hc4053a9;
      16379: inst = 32'h8220000;
      16380: inst = 32'h10408000;
      16381: inst = 32'hc4053aa;
      16382: inst = 32'h8220000;
      16383: inst = 32'h10408000;
      16384: inst = 32'hc4053ab;
      16385: inst = 32'h8220000;
      16386: inst = 32'h10408000;
      16387: inst = 32'hc4053ac;
      16388: inst = 32'h8220000;
      16389: inst = 32'h10408000;
      16390: inst = 32'hc4053ad;
      16391: inst = 32'h8220000;
      16392: inst = 32'h10408000;
      16393: inst = 32'hc4053ae;
      16394: inst = 32'h8220000;
      16395: inst = 32'h10408000;
      16396: inst = 32'hc4053af;
      16397: inst = 32'h8220000;
      16398: inst = 32'h10408000;
      16399: inst = 32'hc4053b0;
      16400: inst = 32'h8220000;
      16401: inst = 32'h10408000;
      16402: inst = 32'hc4053b1;
      16403: inst = 32'h8220000;
      16404: inst = 32'h10408000;
      16405: inst = 32'hc4053b2;
      16406: inst = 32'h8220000;
      16407: inst = 32'h10408000;
      16408: inst = 32'hc4053b3;
      16409: inst = 32'h8220000;
      16410: inst = 32'h10408000;
      16411: inst = 32'hc4053b4;
      16412: inst = 32'h8220000;
      16413: inst = 32'h10408000;
      16414: inst = 32'hc4053b5;
      16415: inst = 32'h8220000;
      16416: inst = 32'h10408000;
      16417: inst = 32'hc4053b6;
      16418: inst = 32'h8220000;
      16419: inst = 32'h10408000;
      16420: inst = 32'hc4053b7;
      16421: inst = 32'h8220000;
      16422: inst = 32'h10408000;
      16423: inst = 32'hc4053b8;
      16424: inst = 32'h8220000;
      16425: inst = 32'h10408000;
      16426: inst = 32'hc4053b9;
      16427: inst = 32'h8220000;
      16428: inst = 32'h10408000;
      16429: inst = 32'hc4053ba;
      16430: inst = 32'h8220000;
      16431: inst = 32'h10408000;
      16432: inst = 32'hc4053bb;
      16433: inst = 32'h8220000;
      16434: inst = 32'h10408000;
      16435: inst = 32'hc4053bc;
      16436: inst = 32'h8220000;
      16437: inst = 32'h10408000;
      16438: inst = 32'hc4053bd;
      16439: inst = 32'h8220000;
      16440: inst = 32'h10408000;
      16441: inst = 32'hc4053be;
      16442: inst = 32'h8220000;
      16443: inst = 32'h10408000;
      16444: inst = 32'hc4053bf;
      16445: inst = 32'h8220000;
      16446: inst = 32'h10408000;
      16447: inst = 32'hc4053c0;
      16448: inst = 32'h8220000;
      16449: inst = 32'h10408000;
      16450: inst = 32'hc4053c1;
      16451: inst = 32'h8220000;
      16452: inst = 32'h10408000;
      16453: inst = 32'hc4053c2;
      16454: inst = 32'h8220000;
      16455: inst = 32'h10408000;
      16456: inst = 32'hc4053c3;
      16457: inst = 32'h8220000;
      16458: inst = 32'h10408000;
      16459: inst = 32'hc4053c4;
      16460: inst = 32'h8220000;
      16461: inst = 32'h10408000;
      16462: inst = 32'hc4053c5;
      16463: inst = 32'h8220000;
      16464: inst = 32'h10408000;
      16465: inst = 32'hc4053c6;
      16466: inst = 32'h8220000;
      16467: inst = 32'h10408000;
      16468: inst = 32'hc4053c7;
      16469: inst = 32'h8220000;
      16470: inst = 32'h10408000;
      16471: inst = 32'hc4053c8;
      16472: inst = 32'h8220000;
      16473: inst = 32'h10408000;
      16474: inst = 32'hc4053c9;
      16475: inst = 32'h8220000;
      16476: inst = 32'h10408000;
      16477: inst = 32'hc4053ca;
      16478: inst = 32'h8220000;
      16479: inst = 32'h10408000;
      16480: inst = 32'hc4053cb;
      16481: inst = 32'h8220000;
      16482: inst = 32'h10408000;
      16483: inst = 32'hc4053cc;
      16484: inst = 32'h8220000;
      16485: inst = 32'h10408000;
      16486: inst = 32'hc4053cd;
      16487: inst = 32'h8220000;
      16488: inst = 32'h10408000;
      16489: inst = 32'hc4053ce;
      16490: inst = 32'h8220000;
      16491: inst = 32'h10408000;
      16492: inst = 32'hc4053cf;
      16493: inst = 32'h8220000;
      16494: inst = 32'h10408000;
      16495: inst = 32'hc4053d0;
      16496: inst = 32'h8220000;
      16497: inst = 32'h10408000;
      16498: inst = 32'hc4053d1;
      16499: inst = 32'h8220000;
      16500: inst = 32'h10408000;
      16501: inst = 32'hc4053d2;
      16502: inst = 32'h8220000;
      16503: inst = 32'h10408000;
      16504: inst = 32'hc4053d3;
      16505: inst = 32'h8220000;
      16506: inst = 32'h10408000;
      16507: inst = 32'hc4053d4;
      16508: inst = 32'h8220000;
      16509: inst = 32'h10408000;
      16510: inst = 32'hc4053d5;
      16511: inst = 32'h8220000;
      16512: inst = 32'h10408000;
      16513: inst = 32'hc4053d6;
      16514: inst = 32'h8220000;
      16515: inst = 32'h10408000;
      16516: inst = 32'hc4053d7;
      16517: inst = 32'h8220000;
      16518: inst = 32'h10408000;
      16519: inst = 32'hc4053d8;
      16520: inst = 32'h8220000;
      16521: inst = 32'h10408000;
      16522: inst = 32'hc4053ea;
      16523: inst = 32'h8220000;
      16524: inst = 32'h10408000;
      16525: inst = 32'hc4053eb;
      16526: inst = 32'h8220000;
      16527: inst = 32'h10408000;
      16528: inst = 32'hc4053ec;
      16529: inst = 32'h8220000;
      16530: inst = 32'h10408000;
      16531: inst = 32'hc4053ed;
      16532: inst = 32'h8220000;
      16533: inst = 32'h10408000;
      16534: inst = 32'hc4053ee;
      16535: inst = 32'h8220000;
      16536: inst = 32'h10408000;
      16537: inst = 32'hc4053ef;
      16538: inst = 32'h8220000;
      16539: inst = 32'h10408000;
      16540: inst = 32'hc4053f0;
      16541: inst = 32'h8220000;
      16542: inst = 32'h10408000;
      16543: inst = 32'hc4053f1;
      16544: inst = 32'h8220000;
      16545: inst = 32'h10408000;
      16546: inst = 32'hc4053f2;
      16547: inst = 32'h8220000;
      16548: inst = 32'h10408000;
      16549: inst = 32'hc4053f3;
      16550: inst = 32'h8220000;
      16551: inst = 32'h10408000;
      16552: inst = 32'hc4053f4;
      16553: inst = 32'h8220000;
      16554: inst = 32'h10408000;
      16555: inst = 32'hc4053f5;
      16556: inst = 32'h8220000;
      16557: inst = 32'h10408000;
      16558: inst = 32'hc405407;
      16559: inst = 32'h8220000;
      16560: inst = 32'h10408000;
      16561: inst = 32'hc405408;
      16562: inst = 32'h8220000;
      16563: inst = 32'h10408000;
      16564: inst = 32'hc405409;
      16565: inst = 32'h8220000;
      16566: inst = 32'h10408000;
      16567: inst = 32'hc40540a;
      16568: inst = 32'h8220000;
      16569: inst = 32'h10408000;
      16570: inst = 32'hc40540b;
      16571: inst = 32'h8220000;
      16572: inst = 32'h10408000;
      16573: inst = 32'hc40540c;
      16574: inst = 32'h8220000;
      16575: inst = 32'h10408000;
      16576: inst = 32'hc40540d;
      16577: inst = 32'h8220000;
      16578: inst = 32'h10408000;
      16579: inst = 32'hc40540e;
      16580: inst = 32'h8220000;
      16581: inst = 32'h10408000;
      16582: inst = 32'hc40540f;
      16583: inst = 32'h8220000;
      16584: inst = 32'h10408000;
      16585: inst = 32'hc405410;
      16586: inst = 32'h8220000;
      16587: inst = 32'h10408000;
      16588: inst = 32'hc405411;
      16589: inst = 32'h8220000;
      16590: inst = 32'h10408000;
      16591: inst = 32'hc405412;
      16592: inst = 32'h8220000;
      16593: inst = 32'h10408000;
      16594: inst = 32'hc405413;
      16595: inst = 32'h8220000;
      16596: inst = 32'h10408000;
      16597: inst = 32'hc405414;
      16598: inst = 32'h8220000;
      16599: inst = 32'h10408000;
      16600: inst = 32'hc405415;
      16601: inst = 32'h8220000;
      16602: inst = 32'h10408000;
      16603: inst = 32'hc405416;
      16604: inst = 32'h8220000;
      16605: inst = 32'h10408000;
      16606: inst = 32'hc405417;
      16607: inst = 32'h8220000;
      16608: inst = 32'h10408000;
      16609: inst = 32'hc405418;
      16610: inst = 32'h8220000;
      16611: inst = 32'h10408000;
      16612: inst = 32'hc405419;
      16613: inst = 32'h8220000;
      16614: inst = 32'h10408000;
      16615: inst = 32'hc40541a;
      16616: inst = 32'h8220000;
      16617: inst = 32'h10408000;
      16618: inst = 32'hc40541b;
      16619: inst = 32'h8220000;
      16620: inst = 32'h10408000;
      16621: inst = 32'hc40541c;
      16622: inst = 32'h8220000;
      16623: inst = 32'h10408000;
      16624: inst = 32'hc40541d;
      16625: inst = 32'h8220000;
      16626: inst = 32'h10408000;
      16627: inst = 32'hc40541e;
      16628: inst = 32'h8220000;
      16629: inst = 32'h10408000;
      16630: inst = 32'hc40541f;
      16631: inst = 32'h8220000;
      16632: inst = 32'h10408000;
      16633: inst = 32'hc405420;
      16634: inst = 32'h8220000;
      16635: inst = 32'h10408000;
      16636: inst = 32'hc405421;
      16637: inst = 32'h8220000;
      16638: inst = 32'h10408000;
      16639: inst = 32'hc405422;
      16640: inst = 32'h8220000;
      16641: inst = 32'h10408000;
      16642: inst = 32'hc405423;
      16643: inst = 32'h8220000;
      16644: inst = 32'h10408000;
      16645: inst = 32'hc405424;
      16646: inst = 32'h8220000;
      16647: inst = 32'h10408000;
      16648: inst = 32'hc405425;
      16649: inst = 32'h8220000;
      16650: inst = 32'h10408000;
      16651: inst = 32'hc405426;
      16652: inst = 32'h8220000;
      16653: inst = 32'h10408000;
      16654: inst = 32'hc405427;
      16655: inst = 32'h8220000;
      16656: inst = 32'h10408000;
      16657: inst = 32'hc405428;
      16658: inst = 32'h8220000;
      16659: inst = 32'h10408000;
      16660: inst = 32'hc405429;
      16661: inst = 32'h8220000;
      16662: inst = 32'h10408000;
      16663: inst = 32'hc40542a;
      16664: inst = 32'h8220000;
      16665: inst = 32'h10408000;
      16666: inst = 32'hc40542b;
      16667: inst = 32'h8220000;
      16668: inst = 32'h10408000;
      16669: inst = 32'hc40542c;
      16670: inst = 32'h8220000;
      16671: inst = 32'h10408000;
      16672: inst = 32'hc40542d;
      16673: inst = 32'h8220000;
      16674: inst = 32'h10408000;
      16675: inst = 32'hc40542e;
      16676: inst = 32'h8220000;
      16677: inst = 32'h10408000;
      16678: inst = 32'hc40542f;
      16679: inst = 32'h8220000;
      16680: inst = 32'h10408000;
      16681: inst = 32'hc405430;
      16682: inst = 32'h8220000;
      16683: inst = 32'h10408000;
      16684: inst = 32'hc405431;
      16685: inst = 32'h8220000;
      16686: inst = 32'h10408000;
      16687: inst = 32'hc405432;
      16688: inst = 32'h8220000;
      16689: inst = 32'h10408000;
      16690: inst = 32'hc405433;
      16691: inst = 32'h8220000;
      16692: inst = 32'h10408000;
      16693: inst = 32'hc405434;
      16694: inst = 32'h8220000;
      16695: inst = 32'h10408000;
      16696: inst = 32'hc405435;
      16697: inst = 32'h8220000;
      16698: inst = 32'h10408000;
      16699: inst = 32'hc405436;
      16700: inst = 32'h8220000;
      16701: inst = 32'h10408000;
      16702: inst = 32'hc405437;
      16703: inst = 32'h8220000;
      16704: inst = 32'h10408000;
      16705: inst = 32'hc405438;
      16706: inst = 32'h8220000;
      16707: inst = 32'h10408000;
      16708: inst = 32'hc40544a;
      16709: inst = 32'h8220000;
      16710: inst = 32'h10408000;
      16711: inst = 32'hc40544b;
      16712: inst = 32'h8220000;
      16713: inst = 32'h10408000;
      16714: inst = 32'hc40544c;
      16715: inst = 32'h8220000;
      16716: inst = 32'h10408000;
      16717: inst = 32'hc40544d;
      16718: inst = 32'h8220000;
      16719: inst = 32'h10408000;
      16720: inst = 32'hc40544e;
      16721: inst = 32'h8220000;
      16722: inst = 32'h10408000;
      16723: inst = 32'hc40544f;
      16724: inst = 32'h8220000;
      16725: inst = 32'h10408000;
      16726: inst = 32'hc405450;
      16727: inst = 32'h8220000;
      16728: inst = 32'h10408000;
      16729: inst = 32'hc405451;
      16730: inst = 32'h8220000;
      16731: inst = 32'h10408000;
      16732: inst = 32'hc405452;
      16733: inst = 32'h8220000;
      16734: inst = 32'h10408000;
      16735: inst = 32'hc405453;
      16736: inst = 32'h8220000;
      16737: inst = 32'h10408000;
      16738: inst = 32'hc405454;
      16739: inst = 32'h8220000;
      16740: inst = 32'h10408000;
      16741: inst = 32'hc405455;
      16742: inst = 32'h8220000;
      16743: inst = 32'h10408000;
      16744: inst = 32'hc405467;
      16745: inst = 32'h8220000;
      16746: inst = 32'h10408000;
      16747: inst = 32'hc405468;
      16748: inst = 32'h8220000;
      16749: inst = 32'h10408000;
      16750: inst = 32'hc405469;
      16751: inst = 32'h8220000;
      16752: inst = 32'h10408000;
      16753: inst = 32'hc40546a;
      16754: inst = 32'h8220000;
      16755: inst = 32'h10408000;
      16756: inst = 32'hc40546b;
      16757: inst = 32'h8220000;
      16758: inst = 32'h10408000;
      16759: inst = 32'hc40546c;
      16760: inst = 32'h8220000;
      16761: inst = 32'h10408000;
      16762: inst = 32'hc40546d;
      16763: inst = 32'h8220000;
      16764: inst = 32'h10408000;
      16765: inst = 32'hc40546e;
      16766: inst = 32'h8220000;
      16767: inst = 32'h10408000;
      16768: inst = 32'hc40546f;
      16769: inst = 32'h8220000;
      16770: inst = 32'h10408000;
      16771: inst = 32'hc405470;
      16772: inst = 32'h8220000;
      16773: inst = 32'h10408000;
      16774: inst = 32'hc405471;
      16775: inst = 32'h8220000;
      16776: inst = 32'h10408000;
      16777: inst = 32'hc405472;
      16778: inst = 32'h8220000;
      16779: inst = 32'h10408000;
      16780: inst = 32'hc405473;
      16781: inst = 32'h8220000;
      16782: inst = 32'h10408000;
      16783: inst = 32'hc405474;
      16784: inst = 32'h8220000;
      16785: inst = 32'h10408000;
      16786: inst = 32'hc405475;
      16787: inst = 32'h8220000;
      16788: inst = 32'h10408000;
      16789: inst = 32'hc405476;
      16790: inst = 32'h8220000;
      16791: inst = 32'h10408000;
      16792: inst = 32'hc405477;
      16793: inst = 32'h8220000;
      16794: inst = 32'h10408000;
      16795: inst = 32'hc405478;
      16796: inst = 32'h8220000;
      16797: inst = 32'h10408000;
      16798: inst = 32'hc405479;
      16799: inst = 32'h8220000;
      16800: inst = 32'h10408000;
      16801: inst = 32'hc40547a;
      16802: inst = 32'h8220000;
      16803: inst = 32'h10408000;
      16804: inst = 32'hc40547b;
      16805: inst = 32'h8220000;
      16806: inst = 32'h10408000;
      16807: inst = 32'hc40547c;
      16808: inst = 32'h8220000;
      16809: inst = 32'h10408000;
      16810: inst = 32'hc40547d;
      16811: inst = 32'h8220000;
      16812: inst = 32'h10408000;
      16813: inst = 32'hc40547e;
      16814: inst = 32'h8220000;
      16815: inst = 32'h10408000;
      16816: inst = 32'hc40547f;
      16817: inst = 32'h8220000;
      16818: inst = 32'h10408000;
      16819: inst = 32'hc405480;
      16820: inst = 32'h8220000;
      16821: inst = 32'h10408000;
      16822: inst = 32'hc405481;
      16823: inst = 32'h8220000;
      16824: inst = 32'h10408000;
      16825: inst = 32'hc405482;
      16826: inst = 32'h8220000;
      16827: inst = 32'h10408000;
      16828: inst = 32'hc405483;
      16829: inst = 32'h8220000;
      16830: inst = 32'h10408000;
      16831: inst = 32'hc405484;
      16832: inst = 32'h8220000;
      16833: inst = 32'h10408000;
      16834: inst = 32'hc405485;
      16835: inst = 32'h8220000;
      16836: inst = 32'h10408000;
      16837: inst = 32'hc405486;
      16838: inst = 32'h8220000;
      16839: inst = 32'h10408000;
      16840: inst = 32'hc405487;
      16841: inst = 32'h8220000;
      16842: inst = 32'h10408000;
      16843: inst = 32'hc405488;
      16844: inst = 32'h8220000;
      16845: inst = 32'h10408000;
      16846: inst = 32'hc405489;
      16847: inst = 32'h8220000;
      16848: inst = 32'h10408000;
      16849: inst = 32'hc40548a;
      16850: inst = 32'h8220000;
      16851: inst = 32'h10408000;
      16852: inst = 32'hc40548b;
      16853: inst = 32'h8220000;
      16854: inst = 32'h10408000;
      16855: inst = 32'hc40548c;
      16856: inst = 32'h8220000;
      16857: inst = 32'h10408000;
      16858: inst = 32'hc40548d;
      16859: inst = 32'h8220000;
      16860: inst = 32'h10408000;
      16861: inst = 32'hc40548e;
      16862: inst = 32'h8220000;
      16863: inst = 32'h10408000;
      16864: inst = 32'hc40548f;
      16865: inst = 32'h8220000;
      16866: inst = 32'h10408000;
      16867: inst = 32'hc405490;
      16868: inst = 32'h8220000;
      16869: inst = 32'h10408000;
      16870: inst = 32'hc405491;
      16871: inst = 32'h8220000;
      16872: inst = 32'h10408000;
      16873: inst = 32'hc405492;
      16874: inst = 32'h8220000;
      16875: inst = 32'h10408000;
      16876: inst = 32'hc405493;
      16877: inst = 32'h8220000;
      16878: inst = 32'h10408000;
      16879: inst = 32'hc405494;
      16880: inst = 32'h8220000;
      16881: inst = 32'h10408000;
      16882: inst = 32'hc405495;
      16883: inst = 32'h8220000;
      16884: inst = 32'h10408000;
      16885: inst = 32'hc405496;
      16886: inst = 32'h8220000;
      16887: inst = 32'h10408000;
      16888: inst = 32'hc405497;
      16889: inst = 32'h8220000;
      16890: inst = 32'h10408000;
      16891: inst = 32'hc4054aa;
      16892: inst = 32'h8220000;
      16893: inst = 32'h10408000;
      16894: inst = 32'hc4054ab;
      16895: inst = 32'h8220000;
      16896: inst = 32'h10408000;
      16897: inst = 32'hc4054ac;
      16898: inst = 32'h8220000;
      16899: inst = 32'h10408000;
      16900: inst = 32'hc4054ad;
      16901: inst = 32'h8220000;
      16902: inst = 32'h10408000;
      16903: inst = 32'hc4054ae;
      16904: inst = 32'h8220000;
      16905: inst = 32'h10408000;
      16906: inst = 32'hc4054af;
      16907: inst = 32'h8220000;
      16908: inst = 32'h10408000;
      16909: inst = 32'hc4054b0;
      16910: inst = 32'h8220000;
      16911: inst = 32'h10408000;
      16912: inst = 32'hc4054b1;
      16913: inst = 32'h8220000;
      16914: inst = 32'h10408000;
      16915: inst = 32'hc4054b2;
      16916: inst = 32'h8220000;
      16917: inst = 32'h10408000;
      16918: inst = 32'hc4054b3;
      16919: inst = 32'h8220000;
      16920: inst = 32'h10408000;
      16921: inst = 32'hc4054b4;
      16922: inst = 32'h8220000;
      16923: inst = 32'h10408000;
      16924: inst = 32'hc4054b5;
      16925: inst = 32'h8220000;
      16926: inst = 32'h10408000;
      16927: inst = 32'hc4054c8;
      16928: inst = 32'h8220000;
      16929: inst = 32'h10408000;
      16930: inst = 32'hc4054c9;
      16931: inst = 32'h8220000;
      16932: inst = 32'h10408000;
      16933: inst = 32'hc4054ca;
      16934: inst = 32'h8220000;
      16935: inst = 32'h10408000;
      16936: inst = 32'hc4054cb;
      16937: inst = 32'h8220000;
      16938: inst = 32'h10408000;
      16939: inst = 32'hc4054cc;
      16940: inst = 32'h8220000;
      16941: inst = 32'h10408000;
      16942: inst = 32'hc4054cd;
      16943: inst = 32'h8220000;
      16944: inst = 32'h10408000;
      16945: inst = 32'hc4054ce;
      16946: inst = 32'h8220000;
      16947: inst = 32'h10408000;
      16948: inst = 32'hc4054cf;
      16949: inst = 32'h8220000;
      16950: inst = 32'h10408000;
      16951: inst = 32'hc4054d0;
      16952: inst = 32'h8220000;
      16953: inst = 32'h10408000;
      16954: inst = 32'hc4054d1;
      16955: inst = 32'h8220000;
      16956: inst = 32'h10408000;
      16957: inst = 32'hc4054d2;
      16958: inst = 32'h8220000;
      16959: inst = 32'h10408000;
      16960: inst = 32'hc4054d3;
      16961: inst = 32'h8220000;
      16962: inst = 32'h10408000;
      16963: inst = 32'hc4054d4;
      16964: inst = 32'h8220000;
      16965: inst = 32'h10408000;
      16966: inst = 32'hc4054d5;
      16967: inst = 32'h8220000;
      16968: inst = 32'h10408000;
      16969: inst = 32'hc4054d6;
      16970: inst = 32'h8220000;
      16971: inst = 32'h10408000;
      16972: inst = 32'hc4054d7;
      16973: inst = 32'h8220000;
      16974: inst = 32'h10408000;
      16975: inst = 32'hc4054d8;
      16976: inst = 32'h8220000;
      16977: inst = 32'h10408000;
      16978: inst = 32'hc4054d9;
      16979: inst = 32'h8220000;
      16980: inst = 32'h10408000;
      16981: inst = 32'hc4054da;
      16982: inst = 32'h8220000;
      16983: inst = 32'h10408000;
      16984: inst = 32'hc4054db;
      16985: inst = 32'h8220000;
      16986: inst = 32'h10408000;
      16987: inst = 32'hc4054dc;
      16988: inst = 32'h8220000;
      16989: inst = 32'h10408000;
      16990: inst = 32'hc4054dd;
      16991: inst = 32'h8220000;
      16992: inst = 32'h10408000;
      16993: inst = 32'hc4054de;
      16994: inst = 32'h8220000;
      16995: inst = 32'h10408000;
      16996: inst = 32'hc4054df;
      16997: inst = 32'h8220000;
      16998: inst = 32'h10408000;
      16999: inst = 32'hc4054e0;
      17000: inst = 32'h8220000;
      17001: inst = 32'h10408000;
      17002: inst = 32'hc4054e1;
      17003: inst = 32'h8220000;
      17004: inst = 32'h10408000;
      17005: inst = 32'hc4054e2;
      17006: inst = 32'h8220000;
      17007: inst = 32'h10408000;
      17008: inst = 32'hc4054e3;
      17009: inst = 32'h8220000;
      17010: inst = 32'h10408000;
      17011: inst = 32'hc4054e4;
      17012: inst = 32'h8220000;
      17013: inst = 32'h10408000;
      17014: inst = 32'hc4054e5;
      17015: inst = 32'h8220000;
      17016: inst = 32'h10408000;
      17017: inst = 32'hc4054e6;
      17018: inst = 32'h8220000;
      17019: inst = 32'h10408000;
      17020: inst = 32'hc4054e7;
      17021: inst = 32'h8220000;
      17022: inst = 32'h10408000;
      17023: inst = 32'hc4054e8;
      17024: inst = 32'h8220000;
      17025: inst = 32'h10408000;
      17026: inst = 32'hc4054e9;
      17027: inst = 32'h8220000;
      17028: inst = 32'h10408000;
      17029: inst = 32'hc4054ea;
      17030: inst = 32'h8220000;
      17031: inst = 32'h10408000;
      17032: inst = 32'hc4054eb;
      17033: inst = 32'h8220000;
      17034: inst = 32'h10408000;
      17035: inst = 32'hc4054ec;
      17036: inst = 32'h8220000;
      17037: inst = 32'h10408000;
      17038: inst = 32'hc4054ed;
      17039: inst = 32'h8220000;
      17040: inst = 32'h10408000;
      17041: inst = 32'hc4054ee;
      17042: inst = 32'h8220000;
      17043: inst = 32'h10408000;
      17044: inst = 32'hc4054ef;
      17045: inst = 32'h8220000;
      17046: inst = 32'h10408000;
      17047: inst = 32'hc4054f0;
      17048: inst = 32'h8220000;
      17049: inst = 32'h10408000;
      17050: inst = 32'hc4054f1;
      17051: inst = 32'h8220000;
      17052: inst = 32'h10408000;
      17053: inst = 32'hc4054f2;
      17054: inst = 32'h8220000;
      17055: inst = 32'h10408000;
      17056: inst = 32'hc4054f3;
      17057: inst = 32'h8220000;
      17058: inst = 32'h10408000;
      17059: inst = 32'hc4054f4;
      17060: inst = 32'h8220000;
      17061: inst = 32'h10408000;
      17062: inst = 32'hc4054f5;
      17063: inst = 32'h8220000;
      17064: inst = 32'h10408000;
      17065: inst = 32'hc4054f6;
      17066: inst = 32'h8220000;
      17067: inst = 32'h10408000;
      17068: inst = 32'hc40550a;
      17069: inst = 32'h8220000;
      17070: inst = 32'h10408000;
      17071: inst = 32'hc40550b;
      17072: inst = 32'h8220000;
      17073: inst = 32'h10408000;
      17074: inst = 32'hc40550c;
      17075: inst = 32'h8220000;
      17076: inst = 32'h10408000;
      17077: inst = 32'hc40550d;
      17078: inst = 32'h8220000;
      17079: inst = 32'h10408000;
      17080: inst = 32'hc40550e;
      17081: inst = 32'h8220000;
      17082: inst = 32'h10408000;
      17083: inst = 32'hc40550f;
      17084: inst = 32'h8220000;
      17085: inst = 32'h10408000;
      17086: inst = 32'hc405510;
      17087: inst = 32'h8220000;
      17088: inst = 32'h10408000;
      17089: inst = 32'hc405511;
      17090: inst = 32'h8220000;
      17091: inst = 32'h10408000;
      17092: inst = 32'hc405512;
      17093: inst = 32'h8220000;
      17094: inst = 32'h10408000;
      17095: inst = 32'hc405513;
      17096: inst = 32'h8220000;
      17097: inst = 32'h10408000;
      17098: inst = 32'hc405514;
      17099: inst = 32'h8220000;
      17100: inst = 32'h10408000;
      17101: inst = 32'hc405515;
      17102: inst = 32'h8220000;
      17103: inst = 32'h10408000;
      17104: inst = 32'hc405529;
      17105: inst = 32'h8220000;
      17106: inst = 32'h10408000;
      17107: inst = 32'hc40552a;
      17108: inst = 32'h8220000;
      17109: inst = 32'h10408000;
      17110: inst = 32'hc40552b;
      17111: inst = 32'h8220000;
      17112: inst = 32'h10408000;
      17113: inst = 32'hc40552c;
      17114: inst = 32'h8220000;
      17115: inst = 32'h10408000;
      17116: inst = 32'hc40552d;
      17117: inst = 32'h8220000;
      17118: inst = 32'h10408000;
      17119: inst = 32'hc40552e;
      17120: inst = 32'h8220000;
      17121: inst = 32'h10408000;
      17122: inst = 32'hc40552f;
      17123: inst = 32'h8220000;
      17124: inst = 32'h10408000;
      17125: inst = 32'hc405530;
      17126: inst = 32'h8220000;
      17127: inst = 32'h10408000;
      17128: inst = 32'hc405531;
      17129: inst = 32'h8220000;
      17130: inst = 32'h10408000;
      17131: inst = 32'hc405532;
      17132: inst = 32'h8220000;
      17133: inst = 32'h10408000;
      17134: inst = 32'hc405533;
      17135: inst = 32'h8220000;
      17136: inst = 32'h10408000;
      17137: inst = 32'hc405534;
      17138: inst = 32'h8220000;
      17139: inst = 32'h10408000;
      17140: inst = 32'hc405535;
      17141: inst = 32'h8220000;
      17142: inst = 32'h10408000;
      17143: inst = 32'hc405536;
      17144: inst = 32'h8220000;
      17145: inst = 32'h10408000;
      17146: inst = 32'hc405537;
      17147: inst = 32'h8220000;
      17148: inst = 32'h10408000;
      17149: inst = 32'hc405538;
      17150: inst = 32'h8220000;
      17151: inst = 32'h10408000;
      17152: inst = 32'hc405539;
      17153: inst = 32'h8220000;
      17154: inst = 32'h10408000;
      17155: inst = 32'hc40553a;
      17156: inst = 32'h8220000;
      17157: inst = 32'h10408000;
      17158: inst = 32'hc40553b;
      17159: inst = 32'h8220000;
      17160: inst = 32'h10408000;
      17161: inst = 32'hc40553c;
      17162: inst = 32'h8220000;
      17163: inst = 32'h10408000;
      17164: inst = 32'hc40553d;
      17165: inst = 32'h8220000;
      17166: inst = 32'h10408000;
      17167: inst = 32'hc40553e;
      17168: inst = 32'h8220000;
      17169: inst = 32'h10408000;
      17170: inst = 32'hc40553f;
      17171: inst = 32'h8220000;
      17172: inst = 32'h10408000;
      17173: inst = 32'hc405540;
      17174: inst = 32'h8220000;
      17175: inst = 32'h10408000;
      17176: inst = 32'hc405541;
      17177: inst = 32'h8220000;
      17178: inst = 32'h10408000;
      17179: inst = 32'hc405542;
      17180: inst = 32'h8220000;
      17181: inst = 32'h10408000;
      17182: inst = 32'hc405543;
      17183: inst = 32'h8220000;
      17184: inst = 32'h10408000;
      17185: inst = 32'hc405544;
      17186: inst = 32'h8220000;
      17187: inst = 32'h10408000;
      17188: inst = 32'hc405545;
      17189: inst = 32'h8220000;
      17190: inst = 32'h10408000;
      17191: inst = 32'hc405546;
      17192: inst = 32'h8220000;
      17193: inst = 32'h10408000;
      17194: inst = 32'hc405547;
      17195: inst = 32'h8220000;
      17196: inst = 32'h10408000;
      17197: inst = 32'hc405548;
      17198: inst = 32'h8220000;
      17199: inst = 32'h10408000;
      17200: inst = 32'hc405549;
      17201: inst = 32'h8220000;
      17202: inst = 32'h10408000;
      17203: inst = 32'hc40554a;
      17204: inst = 32'h8220000;
      17205: inst = 32'h10408000;
      17206: inst = 32'hc40554b;
      17207: inst = 32'h8220000;
      17208: inst = 32'h10408000;
      17209: inst = 32'hc40554c;
      17210: inst = 32'h8220000;
      17211: inst = 32'h10408000;
      17212: inst = 32'hc40554d;
      17213: inst = 32'h8220000;
      17214: inst = 32'h10408000;
      17215: inst = 32'hc40554e;
      17216: inst = 32'h8220000;
      17217: inst = 32'h10408000;
      17218: inst = 32'hc40554f;
      17219: inst = 32'h8220000;
      17220: inst = 32'h10408000;
      17221: inst = 32'hc405550;
      17222: inst = 32'h8220000;
      17223: inst = 32'h10408000;
      17224: inst = 32'hc405551;
      17225: inst = 32'h8220000;
      17226: inst = 32'h10408000;
      17227: inst = 32'hc405552;
      17228: inst = 32'h8220000;
      17229: inst = 32'h10408000;
      17230: inst = 32'hc405553;
      17231: inst = 32'h8220000;
      17232: inst = 32'h10408000;
      17233: inst = 32'hc405554;
      17234: inst = 32'h8220000;
      17235: inst = 32'h10408000;
      17236: inst = 32'hc405555;
      17237: inst = 32'h8220000;
      17238: inst = 32'h10408000;
      17239: inst = 32'hc40556a;
      17240: inst = 32'h8220000;
      17241: inst = 32'h10408000;
      17242: inst = 32'hc40556b;
      17243: inst = 32'h8220000;
      17244: inst = 32'h10408000;
      17245: inst = 32'hc40556c;
      17246: inst = 32'h8220000;
      17247: inst = 32'h10408000;
      17248: inst = 32'hc40556d;
      17249: inst = 32'h8220000;
      17250: inst = 32'h10408000;
      17251: inst = 32'hc40556e;
      17252: inst = 32'h8220000;
      17253: inst = 32'h10408000;
      17254: inst = 32'hc40556f;
      17255: inst = 32'h8220000;
      17256: inst = 32'h10408000;
      17257: inst = 32'hc405570;
      17258: inst = 32'h8220000;
      17259: inst = 32'h10408000;
      17260: inst = 32'hc405571;
      17261: inst = 32'h8220000;
      17262: inst = 32'h10408000;
      17263: inst = 32'hc405572;
      17264: inst = 32'h8220000;
      17265: inst = 32'h10408000;
      17266: inst = 32'hc405573;
      17267: inst = 32'h8220000;
      17268: inst = 32'h10408000;
      17269: inst = 32'hc405574;
      17270: inst = 32'h8220000;
      17271: inst = 32'h10408000;
      17272: inst = 32'hc405575;
      17273: inst = 32'h8220000;
      17274: inst = 32'h10408000;
      17275: inst = 32'hc40558a;
      17276: inst = 32'h8220000;
      17277: inst = 32'h10408000;
      17278: inst = 32'hc40558b;
      17279: inst = 32'h8220000;
      17280: inst = 32'h10408000;
      17281: inst = 32'hc40558c;
      17282: inst = 32'h8220000;
      17283: inst = 32'h10408000;
      17284: inst = 32'hc40558d;
      17285: inst = 32'h8220000;
      17286: inst = 32'h10408000;
      17287: inst = 32'hc40558e;
      17288: inst = 32'h8220000;
      17289: inst = 32'h10408000;
      17290: inst = 32'hc40558f;
      17291: inst = 32'h8220000;
      17292: inst = 32'h10408000;
      17293: inst = 32'hc405590;
      17294: inst = 32'h8220000;
      17295: inst = 32'h10408000;
      17296: inst = 32'hc405591;
      17297: inst = 32'h8220000;
      17298: inst = 32'h10408000;
      17299: inst = 32'hc405592;
      17300: inst = 32'h8220000;
      17301: inst = 32'h10408000;
      17302: inst = 32'hc405593;
      17303: inst = 32'h8220000;
      17304: inst = 32'h10408000;
      17305: inst = 32'hc405594;
      17306: inst = 32'h8220000;
      17307: inst = 32'h10408000;
      17308: inst = 32'hc405595;
      17309: inst = 32'h8220000;
      17310: inst = 32'h10408000;
      17311: inst = 32'hc405596;
      17312: inst = 32'h8220000;
      17313: inst = 32'h10408000;
      17314: inst = 32'hc405597;
      17315: inst = 32'h8220000;
      17316: inst = 32'h10408000;
      17317: inst = 32'hc405598;
      17318: inst = 32'h8220000;
      17319: inst = 32'h10408000;
      17320: inst = 32'hc405599;
      17321: inst = 32'h8220000;
      17322: inst = 32'h10408000;
      17323: inst = 32'hc40559a;
      17324: inst = 32'h8220000;
      17325: inst = 32'h10408000;
      17326: inst = 32'hc40559b;
      17327: inst = 32'h8220000;
      17328: inst = 32'h10408000;
      17329: inst = 32'hc40559c;
      17330: inst = 32'h8220000;
      17331: inst = 32'h10408000;
      17332: inst = 32'hc40559d;
      17333: inst = 32'h8220000;
      17334: inst = 32'h10408000;
      17335: inst = 32'hc40559e;
      17336: inst = 32'h8220000;
      17337: inst = 32'h10408000;
      17338: inst = 32'hc40559f;
      17339: inst = 32'h8220000;
      17340: inst = 32'h10408000;
      17341: inst = 32'hc4055a0;
      17342: inst = 32'h8220000;
      17343: inst = 32'h10408000;
      17344: inst = 32'hc4055a1;
      17345: inst = 32'h8220000;
      17346: inst = 32'h10408000;
      17347: inst = 32'hc4055a2;
      17348: inst = 32'h8220000;
      17349: inst = 32'h10408000;
      17350: inst = 32'hc4055a3;
      17351: inst = 32'h8220000;
      17352: inst = 32'h10408000;
      17353: inst = 32'hc4055a4;
      17354: inst = 32'h8220000;
      17355: inst = 32'h10408000;
      17356: inst = 32'hc4055a5;
      17357: inst = 32'h8220000;
      17358: inst = 32'h10408000;
      17359: inst = 32'hc4055a6;
      17360: inst = 32'h8220000;
      17361: inst = 32'h10408000;
      17362: inst = 32'hc4055a7;
      17363: inst = 32'h8220000;
      17364: inst = 32'h10408000;
      17365: inst = 32'hc4055a8;
      17366: inst = 32'h8220000;
      17367: inst = 32'h10408000;
      17368: inst = 32'hc4055a9;
      17369: inst = 32'h8220000;
      17370: inst = 32'h10408000;
      17371: inst = 32'hc4055aa;
      17372: inst = 32'h8220000;
      17373: inst = 32'h10408000;
      17374: inst = 32'hc4055ab;
      17375: inst = 32'h8220000;
      17376: inst = 32'h10408000;
      17377: inst = 32'hc4055ac;
      17378: inst = 32'h8220000;
      17379: inst = 32'h10408000;
      17380: inst = 32'hc4055ad;
      17381: inst = 32'h8220000;
      17382: inst = 32'h10408000;
      17383: inst = 32'hc4055ae;
      17384: inst = 32'h8220000;
      17385: inst = 32'h10408000;
      17386: inst = 32'hc4055af;
      17387: inst = 32'h8220000;
      17388: inst = 32'h10408000;
      17389: inst = 32'hc4055b0;
      17390: inst = 32'h8220000;
      17391: inst = 32'h10408000;
      17392: inst = 32'hc4055b1;
      17393: inst = 32'h8220000;
      17394: inst = 32'h10408000;
      17395: inst = 32'hc4055b2;
      17396: inst = 32'h8220000;
      17397: inst = 32'h10408000;
      17398: inst = 32'hc4055b3;
      17399: inst = 32'h8220000;
      17400: inst = 32'h10408000;
      17401: inst = 32'hc4055b4;
      17402: inst = 32'h8220000;
      17403: inst = 32'h10408000;
      17404: inst = 32'hc4055ca;
      17405: inst = 32'h8220000;
      17406: inst = 32'h10408000;
      17407: inst = 32'hc4055cb;
      17408: inst = 32'h8220000;
      17409: inst = 32'h10408000;
      17410: inst = 32'hc4055cc;
      17411: inst = 32'h8220000;
      17412: inst = 32'h10408000;
      17413: inst = 32'hc4055cd;
      17414: inst = 32'h8220000;
      17415: inst = 32'h10408000;
      17416: inst = 32'hc4055ce;
      17417: inst = 32'h8220000;
      17418: inst = 32'h10408000;
      17419: inst = 32'hc4055cf;
      17420: inst = 32'h8220000;
      17421: inst = 32'h10408000;
      17422: inst = 32'hc4055d0;
      17423: inst = 32'h8220000;
      17424: inst = 32'h10408000;
      17425: inst = 32'hc4055d1;
      17426: inst = 32'h8220000;
      17427: inst = 32'h10408000;
      17428: inst = 32'hc4055d2;
      17429: inst = 32'h8220000;
      17430: inst = 32'h10408000;
      17431: inst = 32'hc4055d3;
      17432: inst = 32'h8220000;
      17433: inst = 32'h10408000;
      17434: inst = 32'hc4055d4;
      17435: inst = 32'h8220000;
      17436: inst = 32'h10408000;
      17437: inst = 32'hc4055d5;
      17438: inst = 32'h8220000;
      17439: inst = 32'h10408000;
      17440: inst = 32'hc4055eb;
      17441: inst = 32'h8220000;
      17442: inst = 32'h10408000;
      17443: inst = 32'hc4055ec;
      17444: inst = 32'h8220000;
      17445: inst = 32'h10408000;
      17446: inst = 32'hc4055ed;
      17447: inst = 32'h8220000;
      17448: inst = 32'h10408000;
      17449: inst = 32'hc4055ee;
      17450: inst = 32'h8220000;
      17451: inst = 32'h10408000;
      17452: inst = 32'hc4055ef;
      17453: inst = 32'h8220000;
      17454: inst = 32'h10408000;
      17455: inst = 32'hc4055f0;
      17456: inst = 32'h8220000;
      17457: inst = 32'h10408000;
      17458: inst = 32'hc4055f1;
      17459: inst = 32'h8220000;
      17460: inst = 32'h10408000;
      17461: inst = 32'hc4055f2;
      17462: inst = 32'h8220000;
      17463: inst = 32'h10408000;
      17464: inst = 32'hc4055f3;
      17465: inst = 32'h8220000;
      17466: inst = 32'h10408000;
      17467: inst = 32'hc4055f4;
      17468: inst = 32'h8220000;
      17469: inst = 32'h10408000;
      17470: inst = 32'hc4055f5;
      17471: inst = 32'h8220000;
      17472: inst = 32'h10408000;
      17473: inst = 32'hc4055f6;
      17474: inst = 32'h8220000;
      17475: inst = 32'h10408000;
      17476: inst = 32'hc4055f7;
      17477: inst = 32'h8220000;
      17478: inst = 32'h10408000;
      17479: inst = 32'hc4055f8;
      17480: inst = 32'h8220000;
      17481: inst = 32'h10408000;
      17482: inst = 32'hc4055f9;
      17483: inst = 32'h8220000;
      17484: inst = 32'h10408000;
      17485: inst = 32'hc4055fa;
      17486: inst = 32'h8220000;
      17487: inst = 32'h10408000;
      17488: inst = 32'hc4055fb;
      17489: inst = 32'h8220000;
      17490: inst = 32'h10408000;
      17491: inst = 32'hc4055fc;
      17492: inst = 32'h8220000;
      17493: inst = 32'h10408000;
      17494: inst = 32'hc4055fd;
      17495: inst = 32'h8220000;
      17496: inst = 32'h10408000;
      17497: inst = 32'hc4055fe;
      17498: inst = 32'h8220000;
      17499: inst = 32'h10408000;
      17500: inst = 32'hc4055ff;
      17501: inst = 32'h8220000;
      17502: inst = 32'h10408000;
      17503: inst = 32'hc405600;
      17504: inst = 32'h8220000;
      17505: inst = 32'h10408000;
      17506: inst = 32'hc405601;
      17507: inst = 32'h8220000;
      17508: inst = 32'h10408000;
      17509: inst = 32'hc405602;
      17510: inst = 32'h8220000;
      17511: inst = 32'h10408000;
      17512: inst = 32'hc405603;
      17513: inst = 32'h8220000;
      17514: inst = 32'h10408000;
      17515: inst = 32'hc405604;
      17516: inst = 32'h8220000;
      17517: inst = 32'h10408000;
      17518: inst = 32'hc405605;
      17519: inst = 32'h8220000;
      17520: inst = 32'h10408000;
      17521: inst = 32'hc405606;
      17522: inst = 32'h8220000;
      17523: inst = 32'h10408000;
      17524: inst = 32'hc405607;
      17525: inst = 32'h8220000;
      17526: inst = 32'h10408000;
      17527: inst = 32'hc405608;
      17528: inst = 32'h8220000;
      17529: inst = 32'h10408000;
      17530: inst = 32'hc405609;
      17531: inst = 32'h8220000;
      17532: inst = 32'h10408000;
      17533: inst = 32'hc40560a;
      17534: inst = 32'h8220000;
      17535: inst = 32'h10408000;
      17536: inst = 32'hc40560b;
      17537: inst = 32'h8220000;
      17538: inst = 32'h10408000;
      17539: inst = 32'hc40560c;
      17540: inst = 32'h8220000;
      17541: inst = 32'h10408000;
      17542: inst = 32'hc40560d;
      17543: inst = 32'h8220000;
      17544: inst = 32'h10408000;
      17545: inst = 32'hc40560e;
      17546: inst = 32'h8220000;
      17547: inst = 32'h10408000;
      17548: inst = 32'hc40560f;
      17549: inst = 32'h8220000;
      17550: inst = 32'h10408000;
      17551: inst = 32'hc405610;
      17552: inst = 32'h8220000;
      17553: inst = 32'h10408000;
      17554: inst = 32'hc405611;
      17555: inst = 32'h8220000;
      17556: inst = 32'h10408000;
      17557: inst = 32'hc405612;
      17558: inst = 32'h8220000;
      17559: inst = 32'h10408000;
      17560: inst = 32'hc405613;
      17561: inst = 32'h8220000;
      17562: inst = 32'h10408000;
      17563: inst = 32'hc405614;
      17564: inst = 32'h8220000;
      17565: inst = 32'h10408000;
      17566: inst = 32'hc40562a;
      17567: inst = 32'h8220000;
      17568: inst = 32'h10408000;
      17569: inst = 32'hc40562b;
      17570: inst = 32'h8220000;
      17571: inst = 32'h10408000;
      17572: inst = 32'hc40562c;
      17573: inst = 32'h8220000;
      17574: inst = 32'h10408000;
      17575: inst = 32'hc40562d;
      17576: inst = 32'h8220000;
      17577: inst = 32'h10408000;
      17578: inst = 32'hc40562e;
      17579: inst = 32'h8220000;
      17580: inst = 32'h10408000;
      17581: inst = 32'hc40562f;
      17582: inst = 32'h8220000;
      17583: inst = 32'h10408000;
      17584: inst = 32'hc405630;
      17585: inst = 32'h8220000;
      17586: inst = 32'h10408000;
      17587: inst = 32'hc405631;
      17588: inst = 32'h8220000;
      17589: inst = 32'h10408000;
      17590: inst = 32'hc405632;
      17591: inst = 32'h8220000;
      17592: inst = 32'h10408000;
      17593: inst = 32'hc405633;
      17594: inst = 32'h8220000;
      17595: inst = 32'h10408000;
      17596: inst = 32'hc405634;
      17597: inst = 32'h8220000;
      17598: inst = 32'h10408000;
      17599: inst = 32'hc405635;
      17600: inst = 32'h8220000;
      17601: inst = 32'h10408000;
      17602: inst = 32'hc40564b;
      17603: inst = 32'h8220000;
      17604: inst = 32'h10408000;
      17605: inst = 32'hc40564c;
      17606: inst = 32'h8220000;
      17607: inst = 32'h10408000;
      17608: inst = 32'hc40564d;
      17609: inst = 32'h8220000;
      17610: inst = 32'h10408000;
      17611: inst = 32'hc40564e;
      17612: inst = 32'h8220000;
      17613: inst = 32'h10408000;
      17614: inst = 32'hc40564f;
      17615: inst = 32'h8220000;
      17616: inst = 32'h10408000;
      17617: inst = 32'hc405650;
      17618: inst = 32'h8220000;
      17619: inst = 32'h10408000;
      17620: inst = 32'hc405651;
      17621: inst = 32'h8220000;
      17622: inst = 32'h10408000;
      17623: inst = 32'hc405652;
      17624: inst = 32'h8220000;
      17625: inst = 32'h10408000;
      17626: inst = 32'hc405653;
      17627: inst = 32'h8220000;
      17628: inst = 32'h10408000;
      17629: inst = 32'hc405654;
      17630: inst = 32'h8220000;
      17631: inst = 32'h10408000;
      17632: inst = 32'hc405655;
      17633: inst = 32'h8220000;
      17634: inst = 32'h10408000;
      17635: inst = 32'hc405656;
      17636: inst = 32'h8220000;
      17637: inst = 32'h10408000;
      17638: inst = 32'hc405657;
      17639: inst = 32'h8220000;
      17640: inst = 32'h10408000;
      17641: inst = 32'hc405658;
      17642: inst = 32'h8220000;
      17643: inst = 32'h10408000;
      17644: inst = 32'hc405659;
      17645: inst = 32'h8220000;
      17646: inst = 32'h10408000;
      17647: inst = 32'hc40565a;
      17648: inst = 32'h8220000;
      17649: inst = 32'h10408000;
      17650: inst = 32'hc40565b;
      17651: inst = 32'h8220000;
      17652: inst = 32'h10408000;
      17653: inst = 32'hc40565c;
      17654: inst = 32'h8220000;
      17655: inst = 32'h10408000;
      17656: inst = 32'hc40565d;
      17657: inst = 32'h8220000;
      17658: inst = 32'h10408000;
      17659: inst = 32'hc40565e;
      17660: inst = 32'h8220000;
      17661: inst = 32'h10408000;
      17662: inst = 32'hc40565f;
      17663: inst = 32'h8220000;
      17664: inst = 32'h10408000;
      17665: inst = 32'hc405660;
      17666: inst = 32'h8220000;
      17667: inst = 32'h10408000;
      17668: inst = 32'hc405661;
      17669: inst = 32'h8220000;
      17670: inst = 32'h10408000;
      17671: inst = 32'hc405662;
      17672: inst = 32'h8220000;
      17673: inst = 32'h10408000;
      17674: inst = 32'hc405663;
      17675: inst = 32'h8220000;
      17676: inst = 32'h10408000;
      17677: inst = 32'hc405664;
      17678: inst = 32'h8220000;
      17679: inst = 32'h10408000;
      17680: inst = 32'hc405665;
      17681: inst = 32'h8220000;
      17682: inst = 32'h10408000;
      17683: inst = 32'hc405666;
      17684: inst = 32'h8220000;
      17685: inst = 32'h10408000;
      17686: inst = 32'hc405667;
      17687: inst = 32'h8220000;
      17688: inst = 32'h10408000;
      17689: inst = 32'hc405668;
      17690: inst = 32'h8220000;
      17691: inst = 32'h10408000;
      17692: inst = 32'hc405669;
      17693: inst = 32'h8220000;
      17694: inst = 32'h10408000;
      17695: inst = 32'hc40566a;
      17696: inst = 32'h8220000;
      17697: inst = 32'h10408000;
      17698: inst = 32'hc40566b;
      17699: inst = 32'h8220000;
      17700: inst = 32'h10408000;
      17701: inst = 32'hc40566c;
      17702: inst = 32'h8220000;
      17703: inst = 32'h10408000;
      17704: inst = 32'hc40566d;
      17705: inst = 32'h8220000;
      17706: inst = 32'h10408000;
      17707: inst = 32'hc40566e;
      17708: inst = 32'h8220000;
      17709: inst = 32'h10408000;
      17710: inst = 32'hc40566f;
      17711: inst = 32'h8220000;
      17712: inst = 32'h10408000;
      17713: inst = 32'hc405670;
      17714: inst = 32'h8220000;
      17715: inst = 32'h10408000;
      17716: inst = 32'hc405671;
      17717: inst = 32'h8220000;
      17718: inst = 32'h10408000;
      17719: inst = 32'hc405672;
      17720: inst = 32'h8220000;
      17721: inst = 32'h10408000;
      17722: inst = 32'hc405673;
      17723: inst = 32'h8220000;
      17724: inst = 32'h10408000;
      17725: inst = 32'hc40568a;
      17726: inst = 32'h8220000;
      17727: inst = 32'h10408000;
      17728: inst = 32'hc40568b;
      17729: inst = 32'h8220000;
      17730: inst = 32'h10408000;
      17731: inst = 32'hc40568c;
      17732: inst = 32'h8220000;
      17733: inst = 32'h10408000;
      17734: inst = 32'hc40568d;
      17735: inst = 32'h8220000;
      17736: inst = 32'h10408000;
      17737: inst = 32'hc40568e;
      17738: inst = 32'h8220000;
      17739: inst = 32'h10408000;
      17740: inst = 32'hc40568f;
      17741: inst = 32'h8220000;
      17742: inst = 32'h10408000;
      17743: inst = 32'hc405690;
      17744: inst = 32'h8220000;
      17745: inst = 32'h10408000;
      17746: inst = 32'hc405691;
      17747: inst = 32'h8220000;
      17748: inst = 32'h10408000;
      17749: inst = 32'hc405692;
      17750: inst = 32'h8220000;
      17751: inst = 32'h10408000;
      17752: inst = 32'hc405693;
      17753: inst = 32'h8220000;
      17754: inst = 32'h10408000;
      17755: inst = 32'hc405694;
      17756: inst = 32'h8220000;
      17757: inst = 32'h10408000;
      17758: inst = 32'hc405695;
      17759: inst = 32'h8220000;
      17760: inst = 32'h10408000;
      17761: inst = 32'hc4056ac;
      17762: inst = 32'h8220000;
      17763: inst = 32'h10408000;
      17764: inst = 32'hc4056ad;
      17765: inst = 32'h8220000;
      17766: inst = 32'h10408000;
      17767: inst = 32'hc4056ae;
      17768: inst = 32'h8220000;
      17769: inst = 32'h10408000;
      17770: inst = 32'hc4056af;
      17771: inst = 32'h8220000;
      17772: inst = 32'h10408000;
      17773: inst = 32'hc4056b0;
      17774: inst = 32'h8220000;
      17775: inst = 32'h10408000;
      17776: inst = 32'hc4056b1;
      17777: inst = 32'h8220000;
      17778: inst = 32'h10408000;
      17779: inst = 32'hc4056b2;
      17780: inst = 32'h8220000;
      17781: inst = 32'h10408000;
      17782: inst = 32'hc4056b3;
      17783: inst = 32'h8220000;
      17784: inst = 32'h10408000;
      17785: inst = 32'hc4056b4;
      17786: inst = 32'h8220000;
      17787: inst = 32'h10408000;
      17788: inst = 32'hc4056b5;
      17789: inst = 32'h8220000;
      17790: inst = 32'h10408000;
      17791: inst = 32'hc4056b6;
      17792: inst = 32'h8220000;
      17793: inst = 32'h10408000;
      17794: inst = 32'hc4056b7;
      17795: inst = 32'h8220000;
      17796: inst = 32'h10408000;
      17797: inst = 32'hc4056b8;
      17798: inst = 32'h8220000;
      17799: inst = 32'h10408000;
      17800: inst = 32'hc4056b9;
      17801: inst = 32'h8220000;
      17802: inst = 32'h10408000;
      17803: inst = 32'hc4056ba;
      17804: inst = 32'h8220000;
      17805: inst = 32'h10408000;
      17806: inst = 32'hc4056bb;
      17807: inst = 32'h8220000;
      17808: inst = 32'h10408000;
      17809: inst = 32'hc4056bc;
      17810: inst = 32'h8220000;
      17811: inst = 32'h10408000;
      17812: inst = 32'hc4056bd;
      17813: inst = 32'h8220000;
      17814: inst = 32'h10408000;
      17815: inst = 32'hc4056be;
      17816: inst = 32'h8220000;
      17817: inst = 32'h10408000;
      17818: inst = 32'hc4056bf;
      17819: inst = 32'h8220000;
      17820: inst = 32'h10408000;
      17821: inst = 32'hc4056c0;
      17822: inst = 32'h8220000;
      17823: inst = 32'h10408000;
      17824: inst = 32'hc4056c1;
      17825: inst = 32'h8220000;
      17826: inst = 32'h10408000;
      17827: inst = 32'hc4056c2;
      17828: inst = 32'h8220000;
      17829: inst = 32'h10408000;
      17830: inst = 32'hc4056c3;
      17831: inst = 32'h8220000;
      17832: inst = 32'h10408000;
      17833: inst = 32'hc4056c4;
      17834: inst = 32'h8220000;
      17835: inst = 32'h10408000;
      17836: inst = 32'hc4056c5;
      17837: inst = 32'h8220000;
      17838: inst = 32'h10408000;
      17839: inst = 32'hc4056c6;
      17840: inst = 32'h8220000;
      17841: inst = 32'h10408000;
      17842: inst = 32'hc4056c7;
      17843: inst = 32'h8220000;
      17844: inst = 32'h10408000;
      17845: inst = 32'hc4056c8;
      17846: inst = 32'h8220000;
      17847: inst = 32'h10408000;
      17848: inst = 32'hc4056c9;
      17849: inst = 32'h8220000;
      17850: inst = 32'h10408000;
      17851: inst = 32'hc4056ca;
      17852: inst = 32'h8220000;
      17853: inst = 32'h10408000;
      17854: inst = 32'hc4056cb;
      17855: inst = 32'h8220000;
      17856: inst = 32'h10408000;
      17857: inst = 32'hc4056cc;
      17858: inst = 32'h8220000;
      17859: inst = 32'h10408000;
      17860: inst = 32'hc4056cd;
      17861: inst = 32'h8220000;
      17862: inst = 32'h10408000;
      17863: inst = 32'hc4056ce;
      17864: inst = 32'h8220000;
      17865: inst = 32'h10408000;
      17866: inst = 32'hc4056cf;
      17867: inst = 32'h8220000;
      17868: inst = 32'h10408000;
      17869: inst = 32'hc4056d0;
      17870: inst = 32'h8220000;
      17871: inst = 32'h10408000;
      17872: inst = 32'hc4056d1;
      17873: inst = 32'h8220000;
      17874: inst = 32'h10408000;
      17875: inst = 32'hc4056d2;
      17876: inst = 32'h8220000;
      17877: inst = 32'h10408000;
      17878: inst = 32'hc4056ea;
      17879: inst = 32'h8220000;
      17880: inst = 32'h10408000;
      17881: inst = 32'hc4056eb;
      17882: inst = 32'h8220000;
      17883: inst = 32'h10408000;
      17884: inst = 32'hc4056ec;
      17885: inst = 32'h8220000;
      17886: inst = 32'h10408000;
      17887: inst = 32'hc4056ed;
      17888: inst = 32'h8220000;
      17889: inst = 32'h10408000;
      17890: inst = 32'hc4056ee;
      17891: inst = 32'h8220000;
      17892: inst = 32'h10408000;
      17893: inst = 32'hc4056ef;
      17894: inst = 32'h8220000;
      17895: inst = 32'h10408000;
      17896: inst = 32'hc4056f0;
      17897: inst = 32'h8220000;
      17898: inst = 32'h10408000;
      17899: inst = 32'hc4056f1;
      17900: inst = 32'h8220000;
      17901: inst = 32'h10408000;
      17902: inst = 32'hc4056f2;
      17903: inst = 32'h8220000;
      17904: inst = 32'h10408000;
      17905: inst = 32'hc4056f3;
      17906: inst = 32'h8220000;
      17907: inst = 32'h10408000;
      17908: inst = 32'hc4056f4;
      17909: inst = 32'h8220000;
      17910: inst = 32'h10408000;
      17911: inst = 32'hc4056f5;
      17912: inst = 32'h8220000;
      17913: inst = 32'h10408000;
      17914: inst = 32'hc40570d;
      17915: inst = 32'h8220000;
      17916: inst = 32'h10408000;
      17917: inst = 32'hc40570e;
      17918: inst = 32'h8220000;
      17919: inst = 32'h10408000;
      17920: inst = 32'hc40570f;
      17921: inst = 32'h8220000;
      17922: inst = 32'h10408000;
      17923: inst = 32'hc405710;
      17924: inst = 32'h8220000;
      17925: inst = 32'h10408000;
      17926: inst = 32'hc405711;
      17927: inst = 32'h8220000;
      17928: inst = 32'h10408000;
      17929: inst = 32'hc405712;
      17930: inst = 32'h8220000;
      17931: inst = 32'h10408000;
      17932: inst = 32'hc405713;
      17933: inst = 32'h8220000;
      17934: inst = 32'h10408000;
      17935: inst = 32'hc405714;
      17936: inst = 32'h8220000;
      17937: inst = 32'h10408000;
      17938: inst = 32'hc405715;
      17939: inst = 32'h8220000;
      17940: inst = 32'h10408000;
      17941: inst = 32'hc405716;
      17942: inst = 32'h8220000;
      17943: inst = 32'h10408000;
      17944: inst = 32'hc405717;
      17945: inst = 32'h8220000;
      17946: inst = 32'h10408000;
      17947: inst = 32'hc405718;
      17948: inst = 32'h8220000;
      17949: inst = 32'h10408000;
      17950: inst = 32'hc405719;
      17951: inst = 32'h8220000;
      17952: inst = 32'h10408000;
      17953: inst = 32'hc40571a;
      17954: inst = 32'h8220000;
      17955: inst = 32'h10408000;
      17956: inst = 32'hc40571b;
      17957: inst = 32'h8220000;
      17958: inst = 32'h10408000;
      17959: inst = 32'hc40571c;
      17960: inst = 32'h8220000;
      17961: inst = 32'h10408000;
      17962: inst = 32'hc40571d;
      17963: inst = 32'h8220000;
      17964: inst = 32'h10408000;
      17965: inst = 32'hc40571e;
      17966: inst = 32'h8220000;
      17967: inst = 32'h10408000;
      17968: inst = 32'hc40571f;
      17969: inst = 32'h8220000;
      17970: inst = 32'h10408000;
      17971: inst = 32'hc405720;
      17972: inst = 32'h8220000;
      17973: inst = 32'h10408000;
      17974: inst = 32'hc405721;
      17975: inst = 32'h8220000;
      17976: inst = 32'h10408000;
      17977: inst = 32'hc405722;
      17978: inst = 32'h8220000;
      17979: inst = 32'h10408000;
      17980: inst = 32'hc405723;
      17981: inst = 32'h8220000;
      17982: inst = 32'h10408000;
      17983: inst = 32'hc405724;
      17984: inst = 32'h8220000;
      17985: inst = 32'h10408000;
      17986: inst = 32'hc405725;
      17987: inst = 32'h8220000;
      17988: inst = 32'h10408000;
      17989: inst = 32'hc405726;
      17990: inst = 32'h8220000;
      17991: inst = 32'h10408000;
      17992: inst = 32'hc405727;
      17993: inst = 32'h8220000;
      17994: inst = 32'h10408000;
      17995: inst = 32'hc405728;
      17996: inst = 32'h8220000;
      17997: inst = 32'h10408000;
      17998: inst = 32'hc405729;
      17999: inst = 32'h8220000;
      18000: inst = 32'h10408000;
      18001: inst = 32'hc40572a;
      18002: inst = 32'h8220000;
      18003: inst = 32'h10408000;
      18004: inst = 32'hc40572b;
      18005: inst = 32'h8220000;
      18006: inst = 32'h10408000;
      18007: inst = 32'hc40572c;
      18008: inst = 32'h8220000;
      18009: inst = 32'h10408000;
      18010: inst = 32'hc40572d;
      18011: inst = 32'h8220000;
      18012: inst = 32'h10408000;
      18013: inst = 32'hc40572e;
      18014: inst = 32'h8220000;
      18015: inst = 32'h10408000;
      18016: inst = 32'hc40572f;
      18017: inst = 32'h8220000;
      18018: inst = 32'h10408000;
      18019: inst = 32'hc405730;
      18020: inst = 32'h8220000;
      18021: inst = 32'h10408000;
      18022: inst = 32'hc405731;
      18023: inst = 32'h8220000;
      18024: inst = 32'h10408000;
      18025: inst = 32'hc40574a;
      18026: inst = 32'h8220000;
      18027: inst = 32'h10408000;
      18028: inst = 32'hc40574b;
      18029: inst = 32'h8220000;
      18030: inst = 32'h10408000;
      18031: inst = 32'hc40574c;
      18032: inst = 32'h8220000;
      18033: inst = 32'h10408000;
      18034: inst = 32'hc40574d;
      18035: inst = 32'h8220000;
      18036: inst = 32'h10408000;
      18037: inst = 32'hc40574e;
      18038: inst = 32'h8220000;
      18039: inst = 32'h10408000;
      18040: inst = 32'hc40574f;
      18041: inst = 32'h8220000;
      18042: inst = 32'h10408000;
      18043: inst = 32'hc405750;
      18044: inst = 32'h8220000;
      18045: inst = 32'h10408000;
      18046: inst = 32'hc405751;
      18047: inst = 32'h8220000;
      18048: inst = 32'h10408000;
      18049: inst = 32'hc405752;
      18050: inst = 32'h8220000;
      18051: inst = 32'h10408000;
      18052: inst = 32'hc405753;
      18053: inst = 32'h8220000;
      18054: inst = 32'h10408000;
      18055: inst = 32'hc405754;
      18056: inst = 32'h8220000;
      18057: inst = 32'h10408000;
      18058: inst = 32'hc405755;
      18059: inst = 32'h8220000;
      18060: inst = 32'h10408000;
      18061: inst = 32'hc40576e;
      18062: inst = 32'h8220000;
      18063: inst = 32'h10408000;
      18064: inst = 32'hc40576f;
      18065: inst = 32'h8220000;
      18066: inst = 32'h10408000;
      18067: inst = 32'hc405770;
      18068: inst = 32'h8220000;
      18069: inst = 32'h10408000;
      18070: inst = 32'hc405771;
      18071: inst = 32'h8220000;
      18072: inst = 32'h10408000;
      18073: inst = 32'hc405772;
      18074: inst = 32'h8220000;
      18075: inst = 32'h10408000;
      18076: inst = 32'hc405773;
      18077: inst = 32'h8220000;
      18078: inst = 32'h10408000;
      18079: inst = 32'hc405774;
      18080: inst = 32'h8220000;
      18081: inst = 32'h10408000;
      18082: inst = 32'hc405775;
      18083: inst = 32'h8220000;
      18084: inst = 32'h10408000;
      18085: inst = 32'hc405776;
      18086: inst = 32'h8220000;
      18087: inst = 32'h10408000;
      18088: inst = 32'hc405777;
      18089: inst = 32'h8220000;
      18090: inst = 32'h10408000;
      18091: inst = 32'hc405778;
      18092: inst = 32'h8220000;
      18093: inst = 32'h10408000;
      18094: inst = 32'hc405779;
      18095: inst = 32'h8220000;
      18096: inst = 32'h10408000;
      18097: inst = 32'hc40577a;
      18098: inst = 32'h8220000;
      18099: inst = 32'h10408000;
      18100: inst = 32'hc40577b;
      18101: inst = 32'h8220000;
      18102: inst = 32'h10408000;
      18103: inst = 32'hc40577c;
      18104: inst = 32'h8220000;
      18105: inst = 32'h10408000;
      18106: inst = 32'hc40577d;
      18107: inst = 32'h8220000;
      18108: inst = 32'h10408000;
      18109: inst = 32'hc40577e;
      18110: inst = 32'h8220000;
      18111: inst = 32'h10408000;
      18112: inst = 32'hc40577f;
      18113: inst = 32'h8220000;
      18114: inst = 32'h10408000;
      18115: inst = 32'hc405780;
      18116: inst = 32'h8220000;
      18117: inst = 32'h10408000;
      18118: inst = 32'hc405781;
      18119: inst = 32'h8220000;
      18120: inst = 32'h10408000;
      18121: inst = 32'hc405782;
      18122: inst = 32'h8220000;
      18123: inst = 32'h10408000;
      18124: inst = 32'hc405783;
      18125: inst = 32'h8220000;
      18126: inst = 32'h10408000;
      18127: inst = 32'hc405784;
      18128: inst = 32'h8220000;
      18129: inst = 32'h10408000;
      18130: inst = 32'hc405785;
      18131: inst = 32'h8220000;
      18132: inst = 32'h10408000;
      18133: inst = 32'hc405786;
      18134: inst = 32'h8220000;
      18135: inst = 32'h10408000;
      18136: inst = 32'hc405787;
      18137: inst = 32'h8220000;
      18138: inst = 32'h10408000;
      18139: inst = 32'hc405788;
      18140: inst = 32'h8220000;
      18141: inst = 32'h10408000;
      18142: inst = 32'hc405789;
      18143: inst = 32'h8220000;
      18144: inst = 32'h10408000;
      18145: inst = 32'hc40578a;
      18146: inst = 32'h8220000;
      18147: inst = 32'h10408000;
      18148: inst = 32'hc40578b;
      18149: inst = 32'h8220000;
      18150: inst = 32'h10408000;
      18151: inst = 32'hc40578c;
      18152: inst = 32'h8220000;
      18153: inst = 32'h10408000;
      18154: inst = 32'hc40578d;
      18155: inst = 32'h8220000;
      18156: inst = 32'h10408000;
      18157: inst = 32'hc40578e;
      18158: inst = 32'h8220000;
      18159: inst = 32'h10408000;
      18160: inst = 32'hc40578f;
      18161: inst = 32'h8220000;
      18162: inst = 32'h10408000;
      18163: inst = 32'hc405790;
      18164: inst = 32'h8220000;
      18165: inst = 32'h10408000;
      18166: inst = 32'hc405791;
      18167: inst = 32'h8220000;
      18168: inst = 32'h10408000;
      18169: inst = 32'hc4057aa;
      18170: inst = 32'h8220000;
      18171: inst = 32'h10408000;
      18172: inst = 32'hc4057ab;
      18173: inst = 32'h8220000;
      18174: inst = 32'h10408000;
      18175: inst = 32'hc4057ac;
      18176: inst = 32'h8220000;
      18177: inst = 32'h10408000;
      18178: inst = 32'hc4057ad;
      18179: inst = 32'h8220000;
      18180: inst = 32'h10408000;
      18181: inst = 32'hc4057ae;
      18182: inst = 32'h8220000;
      18183: inst = 32'h10408000;
      18184: inst = 32'hc4057af;
      18185: inst = 32'h8220000;
      18186: inst = 32'h10408000;
      18187: inst = 32'hc4057b0;
      18188: inst = 32'h8220000;
      18189: inst = 32'h10408000;
      18190: inst = 32'hc4057b1;
      18191: inst = 32'h8220000;
      18192: inst = 32'h10408000;
      18193: inst = 32'hc4057b2;
      18194: inst = 32'h8220000;
      18195: inst = 32'h10408000;
      18196: inst = 32'hc4057b3;
      18197: inst = 32'h8220000;
      18198: inst = 32'h10408000;
      18199: inst = 32'hc4057b4;
      18200: inst = 32'h8220000;
      18201: inst = 32'h10408000;
      18202: inst = 32'hc4057b5;
      18203: inst = 32'h8220000;
      18204: inst = 32'h10408000;
      18205: inst = 32'hc4057ce;
      18206: inst = 32'h8220000;
      18207: inst = 32'h10408000;
      18208: inst = 32'hc4057cf;
      18209: inst = 32'h8220000;
      18210: inst = 32'h10408000;
      18211: inst = 32'hc4057d0;
      18212: inst = 32'h8220000;
      18213: inst = 32'h10408000;
      18214: inst = 32'hc4057d1;
      18215: inst = 32'h8220000;
      18216: inst = 32'h10408000;
      18217: inst = 32'hc4057d2;
      18218: inst = 32'h8220000;
      18219: inst = 32'h10408000;
      18220: inst = 32'hc4057d3;
      18221: inst = 32'h8220000;
      18222: inst = 32'h10408000;
      18223: inst = 32'hc4057d4;
      18224: inst = 32'h8220000;
      18225: inst = 32'h10408000;
      18226: inst = 32'hc4057d5;
      18227: inst = 32'h8220000;
      18228: inst = 32'h10408000;
      18229: inst = 32'hc4057d6;
      18230: inst = 32'h8220000;
      18231: inst = 32'h10408000;
      18232: inst = 32'hc4057d7;
      18233: inst = 32'h8220000;
      18234: inst = 32'h10408000;
      18235: inst = 32'hc4057d8;
      18236: inst = 32'h8220000;
      18237: inst = 32'h10408000;
      18238: inst = 32'hc4057d9;
      18239: inst = 32'h8220000;
      18240: inst = 32'h10408000;
      18241: inst = 32'hc4057da;
      18242: inst = 32'h8220000;
      18243: inst = 32'h10408000;
      18244: inst = 32'hc4057db;
      18245: inst = 32'h8220000;
      18246: inst = 32'h10408000;
      18247: inst = 32'hc4057dc;
      18248: inst = 32'h8220000;
      18249: inst = 32'h10408000;
      18250: inst = 32'hc4057dd;
      18251: inst = 32'h8220000;
      18252: inst = 32'h10408000;
      18253: inst = 32'hc4057de;
      18254: inst = 32'h8220000;
      18255: inst = 32'h10408000;
      18256: inst = 32'hc4057df;
      18257: inst = 32'h8220000;
      18258: inst = 32'hc207bd0;
      18259: inst = 32'h10408000;
      18260: inst = 32'hc40531b;
      18261: inst = 32'h8220000;
      18262: inst = 32'h10408000;
      18263: inst = 32'hc405344;
      18264: inst = 32'h8220000;
      18265: inst = 32'hc207bcf;
      18266: inst = 32'h10408000;
      18267: inst = 32'hc405321;
      18268: inst = 32'h8220000;
      18269: inst = 32'h10408000;
      18270: inst = 32'hc40533e;
      18271: inst = 32'h8220000;
      18272: inst = 32'h10408000;
      18273: inst = 32'hc405381;
      18274: inst = 32'h8220000;
      18275: inst = 32'h10408000;
      18276: inst = 32'hc40539e;
      18277: inst = 32'h8220000;
      18278: inst = 32'h10408000;
      18279: inst = 32'hc4053e1;
      18280: inst = 32'h8220000;
      18281: inst = 32'h10408000;
      18282: inst = 32'hc4053fe;
      18283: inst = 32'h8220000;
      18284: inst = 32'h10408000;
      18285: inst = 32'hc405441;
      18286: inst = 32'h8220000;
      18287: inst = 32'h10408000;
      18288: inst = 32'hc405448;
      18289: inst = 32'h8220000;
      18290: inst = 32'h10408000;
      18291: inst = 32'hc405457;
      18292: inst = 32'h8220000;
      18293: inst = 32'h10408000;
      18294: inst = 32'hc40545e;
      18295: inst = 32'h8220000;
      18296: inst = 32'h10408000;
      18297: inst = 32'hc405501;
      18298: inst = 32'h8220000;
      18299: inst = 32'h10408000;
      18300: inst = 32'hc40551e;
      18301: inst = 32'h8220000;
      18302: inst = 32'h10408000;
      18303: inst = 32'hc405561;
      18304: inst = 32'h8220000;
      18305: inst = 32'h10408000;
      18306: inst = 32'hc40557e;
      18307: inst = 32'h8220000;
      18308: inst = 32'h10408000;
      18309: inst = 32'hc4055b9;
      18310: inst = 32'h8220000;
      18311: inst = 32'h10408000;
      18312: inst = 32'hc4055c1;
      18313: inst = 32'h8220000;
      18314: inst = 32'h10408000;
      18315: inst = 32'hc4055de;
      18316: inst = 32'h8220000;
      18317: inst = 32'h10408000;
      18318: inst = 32'hc4055e6;
      18319: inst = 32'h8220000;
      18320: inst = 32'h10408000;
      18321: inst = 32'hc40561e;
      18322: inst = 32'h8220000;
      18323: inst = 32'h10408000;
      18324: inst = 32'hc405621;
      18325: inst = 32'h8220000;
      18326: inst = 32'h10408000;
      18327: inst = 32'hc40563e;
      18328: inst = 32'h8220000;
      18329: inst = 32'h10408000;
      18330: inst = 32'hc405641;
      18331: inst = 32'h8220000;
      18332: inst = 32'h10408000;
      18333: inst = 32'hc405681;
      18334: inst = 32'h8220000;
      18335: inst = 32'h10408000;
      18336: inst = 32'hc405698;
      18337: inst = 32'h8220000;
      18338: inst = 32'h10408000;
      18339: inst = 32'hc40569e;
      18340: inst = 32'h8220000;
      18341: inst = 32'h10408000;
      18342: inst = 32'hc4056e1;
      18343: inst = 32'h8220000;
      18344: inst = 32'h10408000;
      18345: inst = 32'hc4056fe;
      18346: inst = 32'h8220000;
      18347: inst = 32'hc207390;
      18348: inst = 32'h10408000;
      18349: inst = 32'hc40537a;
      18350: inst = 32'h8220000;
      18351: inst = 32'h10408000;
      18352: inst = 32'hc4053a5;
      18353: inst = 32'h8220000;
      18354: inst = 32'hc2052aa;
      18355: inst = 32'h10408000;
      18356: inst = 32'hc405389;
      18357: inst = 32'h8220000;
      18358: inst = 32'h10408000;
      18359: inst = 32'hc405396;
      18360: inst = 32'h8220000;
      18361: inst = 32'h10408000;
      18362: inst = 32'hc4054fb;
      18363: inst = 32'h8220000;
      18364: inst = 32'h10408000;
      18365: inst = 32'hc405503;
      18366: inst = 32'h8220000;
      18367: inst = 32'h10408000;
      18368: inst = 32'hc40551c;
      18369: inst = 32'h8220000;
      18370: inst = 32'h10408000;
      18371: inst = 32'hc405524;
      18372: inst = 32'h8220000;
      18373: inst = 32'h10408000;
      18374: inst = 32'hc4055c8;
      18375: inst = 32'h8220000;
      18376: inst = 32'h10408000;
      18377: inst = 32'hc4055d7;
      18378: inst = 32'h8220000;
      18379: inst = 32'h10408000;
      18380: inst = 32'hc405619;
      18381: inst = 32'h8220000;
      18382: inst = 32'h10408000;
      18383: inst = 32'hc405622;
      18384: inst = 32'h8220000;
      18385: inst = 32'h10408000;
      18386: inst = 32'hc40563d;
      18387: inst = 32'h8220000;
      18388: inst = 32'h10408000;
      18389: inst = 32'hc405646;
      18390: inst = 32'h8220000;
      18391: inst = 32'hc206b70;
      18392: inst = 32'h10408000;
      18393: inst = 32'hc4053d9;
      18394: inst = 32'h8220000;
      18395: inst = 32'h10408000;
      18396: inst = 32'hc405406;
      18397: inst = 32'h8220000;
      18398: inst = 32'h10408000;
      18399: inst = 32'hc405556;
      18400: inst = 32'h8220000;
      18401: inst = 32'h10408000;
      18402: inst = 32'hc405589;
      18403: inst = 32'h8220000;
      18404: inst = 32'h10408000;
      18405: inst = 32'hc4055b5;
      18406: inst = 32'h8220000;
      18407: inst = 32'h10408000;
      18408: inst = 32'hc4055ea;
      18409: inst = 32'h8220000;
      18410: inst = 32'h10408000;
      18411: inst = 32'hc405732;
      18412: inst = 32'h8220000;
      18413: inst = 32'h10408000;
      18414: inst = 32'hc40576d;
      18415: inst = 32'h8220000;
      18416: inst = 32'hc20736e;
      18417: inst = 32'h10408000;
      18418: inst = 32'hc4053e0;
      18419: inst = 32'h8220000;
      18420: inst = 32'h10408000;
      18421: inst = 32'hc4053ff;
      18422: inst = 32'h8220000;
      18423: inst = 32'hc205aaa;
      18424: inst = 32'h10408000;
      18425: inst = 32'hc4053e4;
      18426: inst = 32'h8220000;
      18427: inst = 32'h10408000;
      18428: inst = 32'hc4053fb;
      18429: inst = 32'h8220000;
      18430: inst = 32'hc208431;
      18431: inst = 32'h10408000;
      18432: inst = 32'hc4053e8;
      18433: inst = 32'h8220000;
      18434: inst = 32'h10408000;
      18435: inst = 32'hc4053f7;
      18436: inst = 32'h8220000;
      18437: inst = 32'h10408000;
      18438: inst = 32'hc405439;
      18439: inst = 32'h8220000;
      18440: inst = 32'h10408000;
      18441: inst = 32'hc405466;
      18442: inst = 32'h8220000;
      18443: inst = 32'h10408000;
      18444: inst = 32'hc4055b6;
      18445: inst = 32'h8220000;
      18446: inst = 32'h10408000;
      18447: inst = 32'hc4055e9;
      18448: inst = 32'h8220000;
      18449: inst = 32'h10408000;
      18450: inst = 32'hc405733;
      18451: inst = 32'h8220000;
      18452: inst = 32'h10408000;
      18453: inst = 32'hc40576c;
      18454: inst = 32'h8220000;
      18455: inst = 32'hc206b4d;
      18456: inst = 32'h10408000;
      18457: inst = 32'hc40543c;
      18458: inst = 32'h8220000;
      18459: inst = 32'h10408000;
      18460: inst = 32'hc405444;
      18461: inst = 32'h8220000;
      18462: inst = 32'h10408000;
      18463: inst = 32'hc40545b;
      18464: inst = 32'h8220000;
      18465: inst = 32'h10408000;
      18466: inst = 32'hc405463;
      18467: inst = 32'h8220000;
      18468: inst = 32'h10408000;
      18469: inst = 32'hc405563;
      18470: inst = 32'h8220000;
      18471: inst = 32'h10408000;
      18472: inst = 32'hc40557c;
      18473: inst = 32'h8220000;
      18474: inst = 32'h10408000;
      18475: inst = 32'hc405682;
      18476: inst = 32'h8220000;
      18477: inst = 32'h10408000;
      18478: inst = 32'hc40569d;
      18479: inst = 32'h8220000;
      18480: inst = 32'hc208430;
      18481: inst = 32'h10408000;
      18482: inst = 32'hc405440;
      18483: inst = 32'h8220000;
      18484: inst = 32'h10408000;
      18485: inst = 32'hc40545f;
      18486: inst = 32'h8220000;
      18487: inst = 32'hc207bf1;
      18488: inst = 32'h10408000;
      18489: inst = 32'hc405498;
      18490: inst = 32'h8220000;
      18491: inst = 32'h10408000;
      18492: inst = 32'hc4054c7;
      18493: inst = 32'h8220000;
      18494: inst = 32'h10408000;
      18495: inst = 32'hc405615;
      18496: inst = 32'h8220000;
      18497: inst = 32'h10408000;
      18498: inst = 32'hc40564a;
      18499: inst = 32'h8220000;
      18500: inst = 32'hc207bef;
      18501: inst = 32'h10408000;
      18502: inst = 32'hc40549b;
      18503: inst = 32'h8220000;
      18504: inst = 32'h10408000;
      18505: inst = 32'hc4054c4;
      18506: inst = 32'h8220000;
      18507: inst = 32'h10408000;
      18508: inst = 32'hc405687;
      18509: inst = 32'h8220000;
      18510: inst = 32'h10408000;
      18511: inst = 32'hc4056e2;
      18512: inst = 32'h8220000;
      18513: inst = 32'h10408000;
      18514: inst = 32'hc4056fd;
      18515: inst = 32'h8220000;
      18516: inst = 32'hc205aeb;
      18517: inst = 32'h10408000;
      18518: inst = 32'hc40549f;
      18519: inst = 32'h8220000;
      18520: inst = 32'h10408000;
      18521: inst = 32'hc4054c0;
      18522: inst = 32'h8220000;
      18523: inst = 32'hc206b6e;
      18524: inst = 32'h10408000;
      18525: inst = 32'hc4054a8;
      18526: inst = 32'h8220000;
      18527: inst = 32'h10408000;
      18528: inst = 32'hc4054b7;
      18529: inst = 32'h8220000;
      18530: inst = 32'h10408000;
      18531: inst = 32'hc4056e7;
      18532: inst = 32'h8220000;
      18533: inst = 32'h10408000;
      18534: inst = 32'hc4056f8;
      18535: inst = 32'h8220000;
      18536: inst = 32'hc2073b0;
      18537: inst = 32'h10408000;
      18538: inst = 32'hc4054f7;
      18539: inst = 32'h8220000;
      18540: inst = 32'h10408000;
      18541: inst = 32'hc405528;
      18542: inst = 32'h8220000;
      18543: inst = 32'h10408000;
      18544: inst = 32'hc405674;
      18545: inst = 32'h8220000;
      18546: inst = 32'h10408000;
      18547: inst = 32'hc4056ab;
      18548: inst = 32'h8220000;
      18549: inst = 32'hc2073ae;
      18550: inst = 32'h10408000;
      18551: inst = 32'hc4054ff;
      18552: inst = 32'h8220000;
      18553: inst = 32'h10408000;
      18554: inst = 32'hc405520;
      18555: inst = 32'h8220000;
      18556: inst = 32'hc20632d;
      18557: inst = 32'h10408000;
      18558: inst = 32'hc405508;
      18559: inst = 32'h8220000;
      18560: inst = 32'h10408000;
      18561: inst = 32'hc405517;
      18562: inst = 32'h8220000;
      18563: inst = 32'h10408000;
      18564: inst = 32'hc405747;
      18565: inst = 32'h8220000;
      18566: inst = 32'h10408000;
      18567: inst = 32'hc405758;
      18568: inst = 32'h8220000;
      18569: inst = 32'hc206b2d;
      18570: inst = 32'h10408000;
      18571: inst = 32'hc40555a;
      18572: inst = 32'h8220000;
      18573: inst = 32'h10408000;
      18574: inst = 32'hc405585;
      18575: inst = 32'h8220000;
      18576: inst = 32'hc20630c;
      18577: inst = 32'h10408000;
      18578: inst = 32'hc4055be;
      18579: inst = 32'h8220000;
      18580: inst = 32'h10408000;
      18581: inst = 32'hc4055e1;
      18582: inst = 32'h8220000;
      18583: inst = 32'h10408000;
      18584: inst = 32'hc405678;
      18585: inst = 32'h8220000;
      18586: inst = 32'hc20632c;
      18587: inst = 32'h10408000;
      18588: inst = 32'hc4056a7;
      18589: inst = 32'h8220000;
      18590: inst = 32'hc206b90;
      18591: inst = 32'h10408000;
      18592: inst = 32'hc4056d3;
      18593: inst = 32'h8220000;
      18594: inst = 32'h10408000;
      18595: inst = 32'hc40570c;
      18596: inst = 32'h8220000;
      18597: inst = 32'hc207c11;
      18598: inst = 32'h10408000;
      18599: inst = 32'hc405792;
      18600: inst = 32'h8220000;
      18601: inst = 32'h10408000;
      18602: inst = 32'hc4057cd;
      18603: inst = 32'h8220000;
      18604: inst = 32'h58000000;
      18605: inst = 32'hc20ea25;
      18606: inst = 32'h10408000;
      18607: inst = 32'hc40464d;
      18608: inst = 32'h8220000;
      18609: inst = 32'h10408000;
      18610: inst = 32'hc40464e;
      18611: inst = 32'h8220000;
      18612: inst = 32'h10408000;
      18613: inst = 32'hc40464f;
      18614: inst = 32'h8220000;
      18615: inst = 32'h10408000;
      18616: inst = 32'hc404650;
      18617: inst = 32'h8220000;
      18618: inst = 32'h10408000;
      18619: inst = 32'hc404651;
      18620: inst = 32'h8220000;
      18621: inst = 32'h10408000;
      18622: inst = 32'hc404652;
      18623: inst = 32'h8220000;
      18624: inst = 32'h10408000;
      18625: inst = 32'hc404653;
      18626: inst = 32'h8220000;
      18627: inst = 32'h10408000;
      18628: inst = 32'hc404654;
      18629: inst = 32'h8220000;
      18630: inst = 32'h10408000;
      18631: inst = 32'hc404655;
      18632: inst = 32'h8220000;
      18633: inst = 32'h10408000;
      18634: inst = 32'hc404659;
      18635: inst = 32'h8220000;
      18636: inst = 32'h10408000;
      18637: inst = 32'hc40465a;
      18638: inst = 32'h8220000;
      18639: inst = 32'h10408000;
      18640: inst = 32'hc40465b;
      18641: inst = 32'h8220000;
      18642: inst = 32'h10408000;
      18643: inst = 32'hc40465c;
      18644: inst = 32'h8220000;
      18645: inst = 32'h10408000;
      18646: inst = 32'hc40465d;
      18647: inst = 32'h8220000;
      18648: inst = 32'h10408000;
      18649: inst = 32'hc40465e;
      18650: inst = 32'h8220000;
      18651: inst = 32'h10408000;
      18652: inst = 32'hc40465f;
      18653: inst = 32'h8220000;
      18654: inst = 32'h10408000;
      18655: inst = 32'hc404660;
      18656: inst = 32'h8220000;
      18657: inst = 32'h10408000;
      18658: inst = 32'hc404661;
      18659: inst = 32'h8220000;
      18660: inst = 32'h10408000;
      18661: inst = 32'hc404663;
      18662: inst = 32'h8220000;
      18663: inst = 32'h10408000;
      18664: inst = 32'hc404664;
      18665: inst = 32'h8220000;
      18666: inst = 32'h10408000;
      18667: inst = 32'hc404665;
      18668: inst = 32'h8220000;
      18669: inst = 32'h10408000;
      18670: inst = 32'hc404666;
      18671: inst = 32'h8220000;
      18672: inst = 32'h10408000;
      18673: inst = 32'hc404667;
      18674: inst = 32'h8220000;
      18675: inst = 32'h10408000;
      18676: inst = 32'hc404668;
      18677: inst = 32'h8220000;
      18678: inst = 32'h10408000;
      18679: inst = 32'hc404669;
      18680: inst = 32'h8220000;
      18681: inst = 32'h10408000;
      18682: inst = 32'hc40466a;
      18683: inst = 32'h8220000;
      18684: inst = 32'h10408000;
      18685: inst = 32'hc40466b;
      18686: inst = 32'h8220000;
      18687: inst = 32'h10408000;
      18688: inst = 32'hc404671;
      18689: inst = 32'h8220000;
      18690: inst = 32'h10408000;
      18691: inst = 32'hc404672;
      18692: inst = 32'h8220000;
      18693: inst = 32'h10408000;
      18694: inst = 32'hc404673;
      18695: inst = 32'h8220000;
      18696: inst = 32'h10408000;
      18697: inst = 32'hc404674;
      18698: inst = 32'h8220000;
      18699: inst = 32'h10408000;
      18700: inst = 32'hc404675;
      18701: inst = 32'h8220000;
      18702: inst = 32'h10408000;
      18703: inst = 32'hc404676;
      18704: inst = 32'h8220000;
      18705: inst = 32'h10408000;
      18706: inst = 32'hc404677;
      18707: inst = 32'h8220000;
      18708: inst = 32'h10408000;
      18709: inst = 32'hc404678;
      18710: inst = 32'h8220000;
      18711: inst = 32'h10408000;
      18712: inst = 32'hc404679;
      18713: inst = 32'h8220000;
      18714: inst = 32'h10408000;
      18715: inst = 32'hc40467c;
      18716: inst = 32'h8220000;
      18717: inst = 32'h10408000;
      18718: inst = 32'hc40467d;
      18719: inst = 32'h8220000;
      18720: inst = 32'h10408000;
      18721: inst = 32'hc40467e;
      18722: inst = 32'h8220000;
      18723: inst = 32'h10408000;
      18724: inst = 32'hc40467f;
      18725: inst = 32'h8220000;
      18726: inst = 32'h10408000;
      18727: inst = 32'hc404680;
      18728: inst = 32'h8220000;
      18729: inst = 32'h10408000;
      18730: inst = 32'hc404681;
      18731: inst = 32'h8220000;
      18732: inst = 32'h10408000;
      18733: inst = 32'hc404682;
      18734: inst = 32'h8220000;
      18735: inst = 32'h10408000;
      18736: inst = 32'hc404683;
      18737: inst = 32'h8220000;
      18738: inst = 32'h10408000;
      18739: inst = 32'hc404684;
      18740: inst = 32'h8220000;
      18741: inst = 32'h10408000;
      18742: inst = 32'hc404685;
      18743: inst = 32'h8220000;
      18744: inst = 32'h10408000;
      18745: inst = 32'hc40468b;
      18746: inst = 32'h8220000;
      18747: inst = 32'h10408000;
      18748: inst = 32'hc40468c;
      18749: inst = 32'h8220000;
      18750: inst = 32'h10408000;
      18751: inst = 32'hc40468d;
      18752: inst = 32'h8220000;
      18753: inst = 32'h10408000;
      18754: inst = 32'hc40468e;
      18755: inst = 32'h8220000;
      18756: inst = 32'h10408000;
      18757: inst = 32'hc40468f;
      18758: inst = 32'h8220000;
      18759: inst = 32'h10408000;
      18760: inst = 32'hc404690;
      18761: inst = 32'h8220000;
      18762: inst = 32'h10408000;
      18763: inst = 32'hc404691;
      18764: inst = 32'h8220000;
      18765: inst = 32'h10408000;
      18766: inst = 32'hc404692;
      18767: inst = 32'h8220000;
      18768: inst = 32'h10408000;
      18769: inst = 32'hc404693;
      18770: inst = 32'h8220000;
      18771: inst = 32'h10408000;
      18772: inst = 32'hc4046ac;
      18773: inst = 32'h8220000;
      18774: inst = 32'h10408000;
      18775: inst = 32'hc4046ad;
      18776: inst = 32'h8220000;
      18777: inst = 32'h10408000;
      18778: inst = 32'hc4046ae;
      18779: inst = 32'h8220000;
      18780: inst = 32'h10408000;
      18781: inst = 32'hc4046af;
      18782: inst = 32'h8220000;
      18783: inst = 32'h10408000;
      18784: inst = 32'hc4046b0;
      18785: inst = 32'h8220000;
      18786: inst = 32'h10408000;
      18787: inst = 32'hc4046b1;
      18788: inst = 32'h8220000;
      18789: inst = 32'h10408000;
      18790: inst = 32'hc4046b2;
      18791: inst = 32'h8220000;
      18792: inst = 32'h10408000;
      18793: inst = 32'hc4046b3;
      18794: inst = 32'h8220000;
      18795: inst = 32'h10408000;
      18796: inst = 32'hc4046b4;
      18797: inst = 32'h8220000;
      18798: inst = 32'h10408000;
      18799: inst = 32'hc4046b5;
      18800: inst = 32'h8220000;
      18801: inst = 32'h10408000;
      18802: inst = 32'hc4046b8;
      18803: inst = 32'h8220000;
      18804: inst = 32'h10408000;
      18805: inst = 32'hc4046b9;
      18806: inst = 32'h8220000;
      18807: inst = 32'h10408000;
      18808: inst = 32'hc4046ba;
      18809: inst = 32'h8220000;
      18810: inst = 32'h10408000;
      18811: inst = 32'hc4046bb;
      18812: inst = 32'h8220000;
      18813: inst = 32'h10408000;
      18814: inst = 32'hc4046bc;
      18815: inst = 32'h8220000;
      18816: inst = 32'h10408000;
      18817: inst = 32'hc4046bd;
      18818: inst = 32'h8220000;
      18819: inst = 32'h10408000;
      18820: inst = 32'hc4046be;
      18821: inst = 32'h8220000;
      18822: inst = 32'h10408000;
      18823: inst = 32'hc4046bf;
      18824: inst = 32'h8220000;
      18825: inst = 32'h10408000;
      18826: inst = 32'hc4046c0;
      18827: inst = 32'h8220000;
      18828: inst = 32'h10408000;
      18829: inst = 32'hc4046c1;
      18830: inst = 32'h8220000;
      18831: inst = 32'h10408000;
      18832: inst = 32'hc4046c3;
      18833: inst = 32'h8220000;
      18834: inst = 32'h10408000;
      18835: inst = 32'hc4046c4;
      18836: inst = 32'h8220000;
      18837: inst = 32'h10408000;
      18838: inst = 32'hc4046c5;
      18839: inst = 32'h8220000;
      18840: inst = 32'h10408000;
      18841: inst = 32'hc4046c6;
      18842: inst = 32'h8220000;
      18843: inst = 32'h10408000;
      18844: inst = 32'hc4046c7;
      18845: inst = 32'h8220000;
      18846: inst = 32'h10408000;
      18847: inst = 32'hc4046c8;
      18848: inst = 32'h8220000;
      18849: inst = 32'h10408000;
      18850: inst = 32'hc4046c9;
      18851: inst = 32'h8220000;
      18852: inst = 32'h10408000;
      18853: inst = 32'hc4046ca;
      18854: inst = 32'h8220000;
      18855: inst = 32'h10408000;
      18856: inst = 32'hc4046cb;
      18857: inst = 32'h8220000;
      18858: inst = 32'h10408000;
      18859: inst = 32'hc4046d0;
      18860: inst = 32'h8220000;
      18861: inst = 32'h10408000;
      18862: inst = 32'hc4046d1;
      18863: inst = 32'h8220000;
      18864: inst = 32'h10408000;
      18865: inst = 32'hc4046d2;
      18866: inst = 32'h8220000;
      18867: inst = 32'h10408000;
      18868: inst = 32'hc4046d3;
      18869: inst = 32'h8220000;
      18870: inst = 32'h10408000;
      18871: inst = 32'hc4046d4;
      18872: inst = 32'h8220000;
      18873: inst = 32'h10408000;
      18874: inst = 32'hc4046d5;
      18875: inst = 32'h8220000;
      18876: inst = 32'h10408000;
      18877: inst = 32'hc4046d6;
      18878: inst = 32'h8220000;
      18879: inst = 32'h10408000;
      18880: inst = 32'hc4046d7;
      18881: inst = 32'h8220000;
      18882: inst = 32'h10408000;
      18883: inst = 32'hc4046d8;
      18884: inst = 32'h8220000;
      18885: inst = 32'h10408000;
      18886: inst = 32'hc4046da;
      18887: inst = 32'h8220000;
      18888: inst = 32'h10408000;
      18889: inst = 32'hc4046dc;
      18890: inst = 32'h8220000;
      18891: inst = 32'h10408000;
      18892: inst = 32'hc4046dd;
      18893: inst = 32'h8220000;
      18894: inst = 32'h10408000;
      18895: inst = 32'hc4046de;
      18896: inst = 32'h8220000;
      18897: inst = 32'h10408000;
      18898: inst = 32'hc4046df;
      18899: inst = 32'h8220000;
      18900: inst = 32'h10408000;
      18901: inst = 32'hc4046e0;
      18902: inst = 32'h8220000;
      18903: inst = 32'h10408000;
      18904: inst = 32'hc4046e1;
      18905: inst = 32'h8220000;
      18906: inst = 32'h10408000;
      18907: inst = 32'hc4046e2;
      18908: inst = 32'h8220000;
      18909: inst = 32'h10408000;
      18910: inst = 32'hc4046e3;
      18911: inst = 32'h8220000;
      18912: inst = 32'h10408000;
      18913: inst = 32'hc4046e4;
      18914: inst = 32'h8220000;
      18915: inst = 32'h10408000;
      18916: inst = 32'hc4046e5;
      18917: inst = 32'h8220000;
      18918: inst = 32'h10408000;
      18919: inst = 32'hc4046ea;
      18920: inst = 32'h8220000;
      18921: inst = 32'h10408000;
      18922: inst = 32'hc4046eb;
      18923: inst = 32'h8220000;
      18924: inst = 32'h10408000;
      18925: inst = 32'hc4046ec;
      18926: inst = 32'h8220000;
      18927: inst = 32'h10408000;
      18928: inst = 32'hc4046ed;
      18929: inst = 32'h8220000;
      18930: inst = 32'h10408000;
      18931: inst = 32'hc4046ee;
      18932: inst = 32'h8220000;
      18933: inst = 32'h10408000;
      18934: inst = 32'hc4046ef;
      18935: inst = 32'h8220000;
      18936: inst = 32'h10408000;
      18937: inst = 32'hc4046f0;
      18938: inst = 32'h8220000;
      18939: inst = 32'h10408000;
      18940: inst = 32'hc4046f1;
      18941: inst = 32'h8220000;
      18942: inst = 32'h10408000;
      18943: inst = 32'hc4046f2;
      18944: inst = 32'h8220000;
      18945: inst = 32'h10408000;
      18946: inst = 32'hc4046f3;
      18947: inst = 32'h8220000;
      18948: inst = 32'h10408000;
      18949: inst = 32'hc40470b;
      18950: inst = 32'h8220000;
      18951: inst = 32'h10408000;
      18952: inst = 32'hc40470c;
      18953: inst = 32'h8220000;
      18954: inst = 32'h10408000;
      18955: inst = 32'hc40470d;
      18956: inst = 32'h8220000;
      18957: inst = 32'h10408000;
      18958: inst = 32'hc404717;
      18959: inst = 32'h8220000;
      18960: inst = 32'h10408000;
      18961: inst = 32'hc404718;
      18962: inst = 32'h8220000;
      18963: inst = 32'h10408000;
      18964: inst = 32'hc404719;
      18965: inst = 32'h8220000;
      18966: inst = 32'h10408000;
      18967: inst = 32'hc404728;
      18968: inst = 32'h8220000;
      18969: inst = 32'h10408000;
      18970: inst = 32'hc404729;
      18971: inst = 32'h8220000;
      18972: inst = 32'h10408000;
      18973: inst = 32'hc40472a;
      18974: inst = 32'h8220000;
      18975: inst = 32'h10408000;
      18976: inst = 32'hc40472b;
      18977: inst = 32'h8220000;
      18978: inst = 32'h10408000;
      18979: inst = 32'hc404730;
      18980: inst = 32'h8220000;
      18981: inst = 32'h10408000;
      18982: inst = 32'hc404731;
      18983: inst = 32'h8220000;
      18984: inst = 32'h10408000;
      18985: inst = 32'hc404735;
      18986: inst = 32'h8220000;
      18987: inst = 32'h10408000;
      18988: inst = 32'hc404736;
      18989: inst = 32'h8220000;
      18990: inst = 32'h10408000;
      18991: inst = 32'hc404737;
      18992: inst = 32'h8220000;
      18993: inst = 32'h10408000;
      18994: inst = 32'hc404739;
      18995: inst = 32'h8220000;
      18996: inst = 32'h10408000;
      18997: inst = 32'hc40473a;
      18998: inst = 32'h8220000;
      18999: inst = 32'h10408000;
      19000: inst = 32'hc404742;
      19001: inst = 32'h8220000;
      19002: inst = 32'h10408000;
      19003: inst = 32'hc404743;
      19004: inst = 32'h8220000;
      19005: inst = 32'h10408000;
      19006: inst = 32'hc404744;
      19007: inst = 32'h8220000;
      19008: inst = 32'h10408000;
      19009: inst = 32'hc404745;
      19010: inst = 32'h8220000;
      19011: inst = 32'h10408000;
      19012: inst = 32'hc404749;
      19013: inst = 32'h8220000;
      19014: inst = 32'h10408000;
      19015: inst = 32'hc40474a;
      19016: inst = 32'h8220000;
      19017: inst = 32'h10408000;
      19018: inst = 32'hc40474b;
      19019: inst = 32'h8220000;
      19020: inst = 32'h10408000;
      19021: inst = 32'hc40476b;
      19022: inst = 32'h8220000;
      19023: inst = 32'h10408000;
      19024: inst = 32'hc40476c;
      19025: inst = 32'h8220000;
      19026: inst = 32'h10408000;
      19027: inst = 32'hc404777;
      19028: inst = 32'h8220000;
      19029: inst = 32'h10408000;
      19030: inst = 32'hc404778;
      19031: inst = 32'h8220000;
      19032: inst = 32'h10408000;
      19033: inst = 32'hc404788;
      19034: inst = 32'h8220000;
      19035: inst = 32'h10408000;
      19036: inst = 32'hc404789;
      19037: inst = 32'h8220000;
      19038: inst = 32'h10408000;
      19039: inst = 32'hc40478a;
      19040: inst = 32'h8220000;
      19041: inst = 32'h10408000;
      19042: inst = 32'hc404790;
      19043: inst = 32'h8220000;
      19044: inst = 32'h10408000;
      19045: inst = 32'hc404791;
      19046: inst = 32'h8220000;
      19047: inst = 32'h10408000;
      19048: inst = 32'hc404795;
      19049: inst = 32'h8220000;
      19050: inst = 32'h10408000;
      19051: inst = 32'hc404799;
      19052: inst = 32'h8220000;
      19053: inst = 32'h10408000;
      19054: inst = 32'hc40479a;
      19055: inst = 32'h8220000;
      19056: inst = 32'h10408000;
      19057: inst = 32'hc4047a2;
      19058: inst = 32'h8220000;
      19059: inst = 32'h10408000;
      19060: inst = 32'hc4047a3;
      19061: inst = 32'h8220000;
      19062: inst = 32'h10408000;
      19063: inst = 32'hc4047a4;
      19064: inst = 32'h8220000;
      19065: inst = 32'h10408000;
      19066: inst = 32'hc4047a9;
      19067: inst = 32'h8220000;
      19068: inst = 32'h10408000;
      19069: inst = 32'hc4047aa;
      19070: inst = 32'h8220000;
      19071: inst = 32'h10408000;
      19072: inst = 32'hc4047cb;
      19073: inst = 32'h8220000;
      19074: inst = 32'h10408000;
      19075: inst = 32'hc4047cc;
      19076: inst = 32'h8220000;
      19077: inst = 32'h10408000;
      19078: inst = 32'hc4047ce;
      19079: inst = 32'h8220000;
      19080: inst = 32'h10408000;
      19081: inst = 32'hc4047cf;
      19082: inst = 32'h8220000;
      19083: inst = 32'h10408000;
      19084: inst = 32'hc4047d0;
      19085: inst = 32'h8220000;
      19086: inst = 32'h10408000;
      19087: inst = 32'hc4047d1;
      19088: inst = 32'h8220000;
      19089: inst = 32'h10408000;
      19090: inst = 32'hc4047d2;
      19091: inst = 32'h8220000;
      19092: inst = 32'h10408000;
      19093: inst = 32'hc4047d7;
      19094: inst = 32'h8220000;
      19095: inst = 32'h10408000;
      19096: inst = 32'hc4047d8;
      19097: inst = 32'h8220000;
      19098: inst = 32'h10408000;
      19099: inst = 32'hc4047da;
      19100: inst = 32'h8220000;
      19101: inst = 32'h10408000;
      19102: inst = 32'hc4047db;
      19103: inst = 32'h8220000;
      19104: inst = 32'h10408000;
      19105: inst = 32'hc4047dc;
      19106: inst = 32'h8220000;
      19107: inst = 32'h10408000;
      19108: inst = 32'hc4047dd;
      19109: inst = 32'h8220000;
      19110: inst = 32'h10408000;
      19111: inst = 32'hc4047de;
      19112: inst = 32'h8220000;
      19113: inst = 32'h10408000;
      19114: inst = 32'hc4047e7;
      19115: inst = 32'h8220000;
      19116: inst = 32'h10408000;
      19117: inst = 32'hc4047e8;
      19118: inst = 32'h8220000;
      19119: inst = 32'h10408000;
      19120: inst = 32'hc4047e9;
      19121: inst = 32'h8220000;
      19122: inst = 32'h10408000;
      19123: inst = 32'hc4047f0;
      19124: inst = 32'h8220000;
      19125: inst = 32'h10408000;
      19126: inst = 32'hc4047f1;
      19127: inst = 32'h8220000;
      19128: inst = 32'h10408000;
      19129: inst = 32'hc4047f9;
      19130: inst = 32'h8220000;
      19131: inst = 32'h10408000;
      19132: inst = 32'hc4047fa;
      19133: inst = 32'h8220000;
      19134: inst = 32'h10408000;
      19135: inst = 32'hc404800;
      19136: inst = 32'h8220000;
      19137: inst = 32'h10408000;
      19138: inst = 32'hc404801;
      19139: inst = 32'h8220000;
      19140: inst = 32'h10408000;
      19141: inst = 32'hc404802;
      19142: inst = 32'h8220000;
      19143: inst = 32'h10408000;
      19144: inst = 32'hc404803;
      19145: inst = 32'h8220000;
      19146: inst = 32'h10408000;
      19147: inst = 32'hc404809;
      19148: inst = 32'h8220000;
      19149: inst = 32'h10408000;
      19150: inst = 32'hc40480a;
      19151: inst = 32'h8220000;
      19152: inst = 32'h10408000;
      19153: inst = 32'hc40480c;
      19154: inst = 32'h8220000;
      19155: inst = 32'h10408000;
      19156: inst = 32'hc40480d;
      19157: inst = 32'h8220000;
      19158: inst = 32'h10408000;
      19159: inst = 32'hc40480e;
      19160: inst = 32'h8220000;
      19161: inst = 32'h10408000;
      19162: inst = 32'hc40480f;
      19163: inst = 32'h8220000;
      19164: inst = 32'h10408000;
      19165: inst = 32'hc404810;
      19166: inst = 32'h8220000;
      19167: inst = 32'h10408000;
      19168: inst = 32'hc404811;
      19169: inst = 32'h8220000;
      19170: inst = 32'h10408000;
      19171: inst = 32'hc40482b;
      19172: inst = 32'h8220000;
      19173: inst = 32'h10408000;
      19174: inst = 32'hc40482c;
      19175: inst = 32'h8220000;
      19176: inst = 32'h10408000;
      19177: inst = 32'hc40482e;
      19178: inst = 32'h8220000;
      19179: inst = 32'h10408000;
      19180: inst = 32'hc40482f;
      19181: inst = 32'h8220000;
      19182: inst = 32'h10408000;
      19183: inst = 32'hc404830;
      19184: inst = 32'h8220000;
      19185: inst = 32'h10408000;
      19186: inst = 32'hc404831;
      19187: inst = 32'h8220000;
      19188: inst = 32'h10408000;
      19189: inst = 32'hc404832;
      19190: inst = 32'h8220000;
      19191: inst = 32'h10408000;
      19192: inst = 32'hc404837;
      19193: inst = 32'h8220000;
      19194: inst = 32'h10408000;
      19195: inst = 32'hc404838;
      19196: inst = 32'h8220000;
      19197: inst = 32'h10408000;
      19198: inst = 32'hc40483a;
      19199: inst = 32'h8220000;
      19200: inst = 32'h10408000;
      19201: inst = 32'hc40483b;
      19202: inst = 32'h8220000;
      19203: inst = 32'h10408000;
      19204: inst = 32'hc40483c;
      19205: inst = 32'h8220000;
      19206: inst = 32'h10408000;
      19207: inst = 32'hc40483d;
      19208: inst = 32'h8220000;
      19209: inst = 32'h10408000;
      19210: inst = 32'hc40483e;
      19211: inst = 32'h8220000;
      19212: inst = 32'h10408000;
      19213: inst = 32'hc404846;
      19214: inst = 32'h8220000;
      19215: inst = 32'h10408000;
      19216: inst = 32'hc404847;
      19217: inst = 32'h8220000;
      19218: inst = 32'h10408000;
      19219: inst = 32'hc404848;
      19220: inst = 32'h8220000;
      19221: inst = 32'h10408000;
      19222: inst = 32'hc404850;
      19223: inst = 32'h8220000;
      19224: inst = 32'h10408000;
      19225: inst = 32'hc404851;
      19226: inst = 32'h8220000;
      19227: inst = 32'h10408000;
      19228: inst = 32'hc404859;
      19229: inst = 32'h8220000;
      19230: inst = 32'h10408000;
      19231: inst = 32'hc40485a;
      19232: inst = 32'h8220000;
      19233: inst = 32'h10408000;
      19234: inst = 32'hc40485f;
      19235: inst = 32'h8220000;
      19236: inst = 32'h10408000;
      19237: inst = 32'hc404860;
      19238: inst = 32'h8220000;
      19239: inst = 32'h10408000;
      19240: inst = 32'hc404861;
      19241: inst = 32'h8220000;
      19242: inst = 32'h10408000;
      19243: inst = 32'hc404862;
      19244: inst = 32'h8220000;
      19245: inst = 32'h10408000;
      19246: inst = 32'hc404869;
      19247: inst = 32'h8220000;
      19248: inst = 32'h10408000;
      19249: inst = 32'hc40486a;
      19250: inst = 32'h8220000;
      19251: inst = 32'h10408000;
      19252: inst = 32'hc40486c;
      19253: inst = 32'h8220000;
      19254: inst = 32'h10408000;
      19255: inst = 32'hc40486d;
      19256: inst = 32'h8220000;
      19257: inst = 32'h10408000;
      19258: inst = 32'hc40486e;
      19259: inst = 32'h8220000;
      19260: inst = 32'h10408000;
      19261: inst = 32'hc40486f;
      19262: inst = 32'h8220000;
      19263: inst = 32'h10408000;
      19264: inst = 32'hc404870;
      19265: inst = 32'h8220000;
      19266: inst = 32'h10408000;
      19267: inst = 32'hc404871;
      19268: inst = 32'h8220000;
      19269: inst = 32'h10408000;
      19270: inst = 32'hc404872;
      19271: inst = 32'h8220000;
      19272: inst = 32'h10408000;
      19273: inst = 32'hc40488b;
      19274: inst = 32'h8220000;
      19275: inst = 32'h10408000;
      19276: inst = 32'hc40488c;
      19277: inst = 32'h8220000;
      19278: inst = 32'h10408000;
      19279: inst = 32'hc404897;
      19280: inst = 32'h8220000;
      19281: inst = 32'h10408000;
      19282: inst = 32'hc404898;
      19283: inst = 32'h8220000;
      19284: inst = 32'h10408000;
      19285: inst = 32'hc4048a6;
      19286: inst = 32'h8220000;
      19287: inst = 32'h10408000;
      19288: inst = 32'hc4048b0;
      19289: inst = 32'h8220000;
      19290: inst = 32'h10408000;
      19291: inst = 32'hc4048b1;
      19292: inst = 32'h8220000;
      19293: inst = 32'h10408000;
      19294: inst = 32'hc4048b4;
      19295: inst = 32'h8220000;
      19296: inst = 32'h10408000;
      19297: inst = 32'hc4048b5;
      19298: inst = 32'h8220000;
      19299: inst = 32'h10408000;
      19300: inst = 32'hc4048b9;
      19301: inst = 32'h8220000;
      19302: inst = 32'h10408000;
      19303: inst = 32'hc4048ba;
      19304: inst = 32'h8220000;
      19305: inst = 32'h10408000;
      19306: inst = 32'hc4048bf;
      19307: inst = 32'h8220000;
      19308: inst = 32'h10408000;
      19309: inst = 32'hc4048c9;
      19310: inst = 32'h8220000;
      19311: inst = 32'h10408000;
      19312: inst = 32'hc4048ca;
      19313: inst = 32'h8220000;
      19314: inst = 32'h10408000;
      19315: inst = 32'hc4048d1;
      19316: inst = 32'h8220000;
      19317: inst = 32'h10408000;
      19318: inst = 32'hc4048d2;
      19319: inst = 32'h8220000;
      19320: inst = 32'h10408000;
      19321: inst = 32'hc4048d3;
      19322: inst = 32'h8220000;
      19323: inst = 32'h10408000;
      19324: inst = 32'hc4048eb;
      19325: inst = 32'h8220000;
      19326: inst = 32'h10408000;
      19327: inst = 32'hc4048ec;
      19328: inst = 32'h8220000;
      19329: inst = 32'h10408000;
      19330: inst = 32'hc4048ed;
      19331: inst = 32'h8220000;
      19332: inst = 32'h10408000;
      19333: inst = 32'hc4048ee;
      19334: inst = 32'h8220000;
      19335: inst = 32'h10408000;
      19336: inst = 32'hc4048ef;
      19337: inst = 32'h8220000;
      19338: inst = 32'h10408000;
      19339: inst = 32'hc4048f0;
      19340: inst = 32'h8220000;
      19341: inst = 32'h10408000;
      19342: inst = 32'hc4048f1;
      19343: inst = 32'h8220000;
      19344: inst = 32'h10408000;
      19345: inst = 32'hc4048f2;
      19346: inst = 32'h8220000;
      19347: inst = 32'h10408000;
      19348: inst = 32'hc4048f3;
      19349: inst = 32'h8220000;
      19350: inst = 32'h10408000;
      19351: inst = 32'hc4048f4;
      19352: inst = 32'h8220000;
      19353: inst = 32'h10408000;
      19354: inst = 32'hc4048f5;
      19355: inst = 32'h8220000;
      19356: inst = 32'h10408000;
      19357: inst = 32'hc4048f7;
      19358: inst = 32'h8220000;
      19359: inst = 32'h10408000;
      19360: inst = 32'hc4048f8;
      19361: inst = 32'h8220000;
      19362: inst = 32'h10408000;
      19363: inst = 32'hc4048f9;
      19364: inst = 32'h8220000;
      19365: inst = 32'h10408000;
      19366: inst = 32'hc4048fa;
      19367: inst = 32'h8220000;
      19368: inst = 32'h10408000;
      19369: inst = 32'hc4048fb;
      19370: inst = 32'h8220000;
      19371: inst = 32'h10408000;
      19372: inst = 32'hc4048fc;
      19373: inst = 32'h8220000;
      19374: inst = 32'h10408000;
      19375: inst = 32'hc4048fd;
      19376: inst = 32'h8220000;
      19377: inst = 32'h10408000;
      19378: inst = 32'hc4048fe;
      19379: inst = 32'h8220000;
      19380: inst = 32'h10408000;
      19381: inst = 32'hc4048ff;
      19382: inst = 32'h8220000;
      19383: inst = 32'h10408000;
      19384: inst = 32'hc404900;
      19385: inst = 32'h8220000;
      19386: inst = 32'h10408000;
      19387: inst = 32'hc404901;
      19388: inst = 32'h8220000;
      19389: inst = 32'h10408000;
      19390: inst = 32'hc404904;
      19391: inst = 32'h8220000;
      19392: inst = 32'h10408000;
      19393: inst = 32'hc404905;
      19394: inst = 32'h8220000;
      19395: inst = 32'h10408000;
      19396: inst = 32'hc404906;
      19397: inst = 32'h8220000;
      19398: inst = 32'h10408000;
      19399: inst = 32'hc404907;
      19400: inst = 32'h8220000;
      19401: inst = 32'h10408000;
      19402: inst = 32'hc404908;
      19403: inst = 32'h8220000;
      19404: inst = 32'h10408000;
      19405: inst = 32'hc404909;
      19406: inst = 32'h8220000;
      19407: inst = 32'h10408000;
      19408: inst = 32'hc40490a;
      19409: inst = 32'h8220000;
      19410: inst = 32'h10408000;
      19411: inst = 32'hc40490b;
      19412: inst = 32'h8220000;
      19413: inst = 32'h10408000;
      19414: inst = 32'hc40490c;
      19415: inst = 32'h8220000;
      19416: inst = 32'h10408000;
      19417: inst = 32'hc40490d;
      19418: inst = 32'h8220000;
      19419: inst = 32'h10408000;
      19420: inst = 32'hc404910;
      19421: inst = 32'h8220000;
      19422: inst = 32'h10408000;
      19423: inst = 32'hc404911;
      19424: inst = 32'h8220000;
      19425: inst = 32'h10408000;
      19426: inst = 32'hc404912;
      19427: inst = 32'h8220000;
      19428: inst = 32'h10408000;
      19429: inst = 32'hc404913;
      19430: inst = 32'h8220000;
      19431: inst = 32'h10408000;
      19432: inst = 32'hc404914;
      19433: inst = 32'h8220000;
      19434: inst = 32'h10408000;
      19435: inst = 32'hc404915;
      19436: inst = 32'h8220000;
      19437: inst = 32'h10408000;
      19438: inst = 32'hc404916;
      19439: inst = 32'h8220000;
      19440: inst = 32'h10408000;
      19441: inst = 32'hc404917;
      19442: inst = 32'h8220000;
      19443: inst = 32'h10408000;
      19444: inst = 32'hc404918;
      19445: inst = 32'h8220000;
      19446: inst = 32'h10408000;
      19447: inst = 32'hc404919;
      19448: inst = 32'h8220000;
      19449: inst = 32'h10408000;
      19450: inst = 32'hc40491a;
      19451: inst = 32'h8220000;
      19452: inst = 32'h10408000;
      19453: inst = 32'hc40491e;
      19454: inst = 32'h8220000;
      19455: inst = 32'h10408000;
      19456: inst = 32'hc40491f;
      19457: inst = 32'h8220000;
      19458: inst = 32'h10408000;
      19459: inst = 32'hc404920;
      19460: inst = 32'h8220000;
      19461: inst = 32'h10408000;
      19462: inst = 32'hc404921;
      19463: inst = 32'h8220000;
      19464: inst = 32'h10408000;
      19465: inst = 32'hc404922;
      19466: inst = 32'h8220000;
      19467: inst = 32'h10408000;
      19468: inst = 32'hc404923;
      19469: inst = 32'h8220000;
      19470: inst = 32'h10408000;
      19471: inst = 32'hc404924;
      19472: inst = 32'h8220000;
      19473: inst = 32'h10408000;
      19474: inst = 32'hc404925;
      19475: inst = 32'h8220000;
      19476: inst = 32'h10408000;
      19477: inst = 32'hc404926;
      19478: inst = 32'h8220000;
      19479: inst = 32'h10408000;
      19480: inst = 32'hc404927;
      19481: inst = 32'h8220000;
      19482: inst = 32'h10408000;
      19483: inst = 32'hc404929;
      19484: inst = 32'h8220000;
      19485: inst = 32'h10408000;
      19486: inst = 32'hc40492a;
      19487: inst = 32'h8220000;
      19488: inst = 32'h10408000;
      19489: inst = 32'hc40492b;
      19490: inst = 32'h8220000;
      19491: inst = 32'h10408000;
      19492: inst = 32'hc40492c;
      19493: inst = 32'h8220000;
      19494: inst = 32'h10408000;
      19495: inst = 32'hc40492d;
      19496: inst = 32'h8220000;
      19497: inst = 32'h10408000;
      19498: inst = 32'hc40492e;
      19499: inst = 32'h8220000;
      19500: inst = 32'h10408000;
      19501: inst = 32'hc40492f;
      19502: inst = 32'h8220000;
      19503: inst = 32'h10408000;
      19504: inst = 32'hc404930;
      19505: inst = 32'h8220000;
      19506: inst = 32'h10408000;
      19507: inst = 32'hc404931;
      19508: inst = 32'h8220000;
      19509: inst = 32'h10408000;
      19510: inst = 32'hc404932;
      19511: inst = 32'h8220000;
      19512: inst = 32'h10408000;
      19513: inst = 32'hc404933;
      19514: inst = 32'h8220000;
      19515: inst = 32'h10408000;
      19516: inst = 32'hc40494b;
      19517: inst = 32'h8220000;
      19518: inst = 32'h10408000;
      19519: inst = 32'hc40494c;
      19520: inst = 32'h8220000;
      19521: inst = 32'h10408000;
      19522: inst = 32'hc40494d;
      19523: inst = 32'h8220000;
      19524: inst = 32'h10408000;
      19525: inst = 32'hc40494e;
      19526: inst = 32'h8220000;
      19527: inst = 32'h10408000;
      19528: inst = 32'hc40494f;
      19529: inst = 32'h8220000;
      19530: inst = 32'h10408000;
      19531: inst = 32'hc404950;
      19532: inst = 32'h8220000;
      19533: inst = 32'h10408000;
      19534: inst = 32'hc404951;
      19535: inst = 32'h8220000;
      19536: inst = 32'h10408000;
      19537: inst = 32'hc404952;
      19538: inst = 32'h8220000;
      19539: inst = 32'h10408000;
      19540: inst = 32'hc404953;
      19541: inst = 32'h8220000;
      19542: inst = 32'h10408000;
      19543: inst = 32'hc404954;
      19544: inst = 32'h8220000;
      19545: inst = 32'h10408000;
      19546: inst = 32'hc404957;
      19547: inst = 32'h8220000;
      19548: inst = 32'h10408000;
      19549: inst = 32'hc404958;
      19550: inst = 32'h8220000;
      19551: inst = 32'h10408000;
      19552: inst = 32'hc404959;
      19553: inst = 32'h8220000;
      19554: inst = 32'h10408000;
      19555: inst = 32'hc40495a;
      19556: inst = 32'h8220000;
      19557: inst = 32'h10408000;
      19558: inst = 32'hc40495b;
      19559: inst = 32'h8220000;
      19560: inst = 32'h10408000;
      19561: inst = 32'hc40495c;
      19562: inst = 32'h8220000;
      19563: inst = 32'h10408000;
      19564: inst = 32'hc40495d;
      19565: inst = 32'h8220000;
      19566: inst = 32'h10408000;
      19567: inst = 32'hc40495e;
      19568: inst = 32'h8220000;
      19569: inst = 32'h10408000;
      19570: inst = 32'hc40495f;
      19571: inst = 32'h8220000;
      19572: inst = 32'h10408000;
      19573: inst = 32'hc404960;
      19574: inst = 32'h8220000;
      19575: inst = 32'h10408000;
      19576: inst = 32'hc404961;
      19577: inst = 32'h8220000;
      19578: inst = 32'h10408000;
      19579: inst = 32'hc404963;
      19580: inst = 32'h8220000;
      19581: inst = 32'h10408000;
      19582: inst = 32'hc404964;
      19583: inst = 32'h8220000;
      19584: inst = 32'h10408000;
      19585: inst = 32'hc404965;
      19586: inst = 32'h8220000;
      19587: inst = 32'h10408000;
      19588: inst = 32'hc404966;
      19589: inst = 32'h8220000;
      19590: inst = 32'h10408000;
      19591: inst = 32'hc404967;
      19592: inst = 32'h8220000;
      19593: inst = 32'h10408000;
      19594: inst = 32'hc404968;
      19595: inst = 32'h8220000;
      19596: inst = 32'h10408000;
      19597: inst = 32'hc404969;
      19598: inst = 32'h8220000;
      19599: inst = 32'h10408000;
      19600: inst = 32'hc40496a;
      19601: inst = 32'h8220000;
      19602: inst = 32'h10408000;
      19603: inst = 32'hc40496b;
      19604: inst = 32'h8220000;
      19605: inst = 32'h10408000;
      19606: inst = 32'hc40496c;
      19607: inst = 32'h8220000;
      19608: inst = 32'h10408000;
      19609: inst = 32'hc40496d;
      19610: inst = 32'h8220000;
      19611: inst = 32'h10408000;
      19612: inst = 32'hc404970;
      19613: inst = 32'h8220000;
      19614: inst = 32'h10408000;
      19615: inst = 32'hc404971;
      19616: inst = 32'h8220000;
      19617: inst = 32'h10408000;
      19618: inst = 32'hc404972;
      19619: inst = 32'h8220000;
      19620: inst = 32'h10408000;
      19621: inst = 32'hc404973;
      19622: inst = 32'h8220000;
      19623: inst = 32'h10408000;
      19624: inst = 32'hc404974;
      19625: inst = 32'h8220000;
      19626: inst = 32'h10408000;
      19627: inst = 32'hc404975;
      19628: inst = 32'h8220000;
      19629: inst = 32'h10408000;
      19630: inst = 32'hc404976;
      19631: inst = 32'h8220000;
      19632: inst = 32'h10408000;
      19633: inst = 32'hc404977;
      19634: inst = 32'h8220000;
      19635: inst = 32'h10408000;
      19636: inst = 32'hc404978;
      19637: inst = 32'h8220000;
      19638: inst = 32'h10408000;
      19639: inst = 32'hc404979;
      19640: inst = 32'h8220000;
      19641: inst = 32'h10408000;
      19642: inst = 32'hc40497d;
      19643: inst = 32'h8220000;
      19644: inst = 32'h10408000;
      19645: inst = 32'hc40497e;
      19646: inst = 32'h8220000;
      19647: inst = 32'h10408000;
      19648: inst = 32'hc40497f;
      19649: inst = 32'h8220000;
      19650: inst = 32'h10408000;
      19651: inst = 32'hc404980;
      19652: inst = 32'h8220000;
      19653: inst = 32'h10408000;
      19654: inst = 32'hc404981;
      19655: inst = 32'h8220000;
      19656: inst = 32'h10408000;
      19657: inst = 32'hc404982;
      19658: inst = 32'h8220000;
      19659: inst = 32'h10408000;
      19660: inst = 32'hc404983;
      19661: inst = 32'h8220000;
      19662: inst = 32'h10408000;
      19663: inst = 32'hc404984;
      19664: inst = 32'h8220000;
      19665: inst = 32'h10408000;
      19666: inst = 32'hc404985;
      19667: inst = 32'h8220000;
      19668: inst = 32'h10408000;
      19669: inst = 32'hc404986;
      19670: inst = 32'h8220000;
      19671: inst = 32'h10408000;
      19672: inst = 32'hc404987;
      19673: inst = 32'h8220000;
      19674: inst = 32'h10408000;
      19675: inst = 32'hc404989;
      19676: inst = 32'h8220000;
      19677: inst = 32'h10408000;
      19678: inst = 32'hc40498a;
      19679: inst = 32'h8220000;
      19680: inst = 32'h10408000;
      19681: inst = 32'hc40498b;
      19682: inst = 32'h8220000;
      19683: inst = 32'h10408000;
      19684: inst = 32'hc40498c;
      19685: inst = 32'h8220000;
      19686: inst = 32'h10408000;
      19687: inst = 32'hc40498d;
      19688: inst = 32'h8220000;
      19689: inst = 32'h10408000;
      19690: inst = 32'hc40498e;
      19691: inst = 32'h8220000;
      19692: inst = 32'h10408000;
      19693: inst = 32'hc40498f;
      19694: inst = 32'h8220000;
      19695: inst = 32'h10408000;
      19696: inst = 32'hc404990;
      19697: inst = 32'h8220000;
      19698: inst = 32'h10408000;
      19699: inst = 32'hc404991;
      19700: inst = 32'h8220000;
      19701: inst = 32'h10408000;
      19702: inst = 32'hc404992;
      19703: inst = 32'h8220000;
      19704: inst = 32'h10408000;
      19705: inst = 32'hc404993;
      19706: inst = 32'h8220000;
      19707: inst = 32'h10408000;
      19708: inst = 32'hc404dcd;
      19709: inst = 32'h8220000;
      19710: inst = 32'h10408000;
      19711: inst = 32'hc404dce;
      19712: inst = 32'h8220000;
      19713: inst = 32'h10408000;
      19714: inst = 32'hc404dcf;
      19715: inst = 32'h8220000;
      19716: inst = 32'h10408000;
      19717: inst = 32'hc404dd0;
      19718: inst = 32'h8220000;
      19719: inst = 32'h10408000;
      19720: inst = 32'hc404dd1;
      19721: inst = 32'h8220000;
      19722: inst = 32'h10408000;
      19723: inst = 32'hc404dd2;
      19724: inst = 32'h8220000;
      19725: inst = 32'h10408000;
      19726: inst = 32'hc404dd3;
      19727: inst = 32'h8220000;
      19728: inst = 32'h10408000;
      19729: inst = 32'hc404dd4;
      19730: inst = 32'h8220000;
      19731: inst = 32'h10408000;
      19732: inst = 32'hc404dd5;
      19733: inst = 32'h8220000;
      19734: inst = 32'h10408000;
      19735: inst = 32'hc404dd7;
      19736: inst = 32'h8220000;
      19737: inst = 32'h10408000;
      19738: inst = 32'hc404dd8;
      19739: inst = 32'h8220000;
      19740: inst = 32'h10408000;
      19741: inst = 32'hc404dd9;
      19742: inst = 32'h8220000;
      19743: inst = 32'h10408000;
      19744: inst = 32'hc404dda;
      19745: inst = 32'h8220000;
      19746: inst = 32'h10408000;
      19747: inst = 32'hc404ddb;
      19748: inst = 32'h8220000;
      19749: inst = 32'h10408000;
      19750: inst = 32'hc404ddc;
      19751: inst = 32'h8220000;
      19752: inst = 32'h10408000;
      19753: inst = 32'hc404ddd;
      19754: inst = 32'h8220000;
      19755: inst = 32'h10408000;
      19756: inst = 32'hc404dde;
      19757: inst = 32'h8220000;
      19758: inst = 32'h10408000;
      19759: inst = 32'hc404ddf;
      19760: inst = 32'h8220000;
      19761: inst = 32'h10408000;
      19762: inst = 32'hc404de0;
      19763: inst = 32'h8220000;
      19764: inst = 32'h10408000;
      19765: inst = 32'hc404de1;
      19766: inst = 32'h8220000;
      19767: inst = 32'h10408000;
      19768: inst = 32'hc404de2;
      19769: inst = 32'h8220000;
      19770: inst = 32'h10408000;
      19771: inst = 32'hc404de4;
      19772: inst = 32'h8220000;
      19773: inst = 32'h10408000;
      19774: inst = 32'hc404de5;
      19775: inst = 32'h8220000;
      19776: inst = 32'h10408000;
      19777: inst = 32'hc404de6;
      19778: inst = 32'h8220000;
      19779: inst = 32'h10408000;
      19780: inst = 32'hc404de7;
      19781: inst = 32'h8220000;
      19782: inst = 32'h10408000;
      19783: inst = 32'hc404de8;
      19784: inst = 32'h8220000;
      19785: inst = 32'h10408000;
      19786: inst = 32'hc404de9;
      19787: inst = 32'h8220000;
      19788: inst = 32'h10408000;
      19789: inst = 32'hc404dea;
      19790: inst = 32'h8220000;
      19791: inst = 32'h10408000;
      19792: inst = 32'hc404deb;
      19793: inst = 32'h8220000;
      19794: inst = 32'h10408000;
      19795: inst = 32'hc404dec;
      19796: inst = 32'h8220000;
      19797: inst = 32'h10408000;
      19798: inst = 32'hc404ded;
      19799: inst = 32'h8220000;
      19800: inst = 32'h10408000;
      19801: inst = 32'hc404df0;
      19802: inst = 32'h8220000;
      19803: inst = 32'h10408000;
      19804: inst = 32'hc404df1;
      19805: inst = 32'h8220000;
      19806: inst = 32'h10408000;
      19807: inst = 32'hc404df2;
      19808: inst = 32'h8220000;
      19809: inst = 32'h10408000;
      19810: inst = 32'hc404dfc;
      19811: inst = 32'h8220000;
      19812: inst = 32'h10408000;
      19813: inst = 32'hc404dfd;
      19814: inst = 32'h8220000;
      19815: inst = 32'h10408000;
      19816: inst = 32'hc404dfe;
      19817: inst = 32'h8220000;
      19818: inst = 32'h10408000;
      19819: inst = 32'hc404dff;
      19820: inst = 32'h8220000;
      19821: inst = 32'h10408000;
      19822: inst = 32'hc404e00;
      19823: inst = 32'h8220000;
      19824: inst = 32'h10408000;
      19825: inst = 32'hc404e01;
      19826: inst = 32'h8220000;
      19827: inst = 32'h10408000;
      19828: inst = 32'hc404e02;
      19829: inst = 32'h8220000;
      19830: inst = 32'h10408000;
      19831: inst = 32'hc404e03;
      19832: inst = 32'h8220000;
      19833: inst = 32'h10408000;
      19834: inst = 32'hc404e04;
      19835: inst = 32'h8220000;
      19836: inst = 32'h10408000;
      19837: inst = 32'hc404e05;
      19838: inst = 32'h8220000;
      19839: inst = 32'h10408000;
      19840: inst = 32'hc404e06;
      19841: inst = 32'h8220000;
      19842: inst = 32'h10408000;
      19843: inst = 32'hc404e07;
      19844: inst = 32'h8220000;
      19845: inst = 32'h10408000;
      19846: inst = 32'hc404e0b;
      19847: inst = 32'h8220000;
      19848: inst = 32'h10408000;
      19849: inst = 32'hc404e0c;
      19850: inst = 32'h8220000;
      19851: inst = 32'h10408000;
      19852: inst = 32'hc404e0d;
      19853: inst = 32'h8220000;
      19854: inst = 32'h10408000;
      19855: inst = 32'hc404e0e;
      19856: inst = 32'h8220000;
      19857: inst = 32'h10408000;
      19858: inst = 32'hc404e0f;
      19859: inst = 32'h8220000;
      19860: inst = 32'h10408000;
      19861: inst = 32'hc404e10;
      19862: inst = 32'h8220000;
      19863: inst = 32'h10408000;
      19864: inst = 32'hc404e11;
      19865: inst = 32'h8220000;
      19866: inst = 32'h10408000;
      19867: inst = 32'hc404e12;
      19868: inst = 32'h8220000;
      19869: inst = 32'h10408000;
      19870: inst = 32'hc404e13;
      19871: inst = 32'h8220000;
      19872: inst = 32'h10408000;
      19873: inst = 32'hc404e2c;
      19874: inst = 32'h8220000;
      19875: inst = 32'h10408000;
      19876: inst = 32'hc404e2d;
      19877: inst = 32'h8220000;
      19878: inst = 32'h10408000;
      19879: inst = 32'hc404e2e;
      19880: inst = 32'h8220000;
      19881: inst = 32'h10408000;
      19882: inst = 32'hc404e2f;
      19883: inst = 32'h8220000;
      19884: inst = 32'h10408000;
      19885: inst = 32'hc404e30;
      19886: inst = 32'h8220000;
      19887: inst = 32'h10408000;
      19888: inst = 32'hc404e31;
      19889: inst = 32'h8220000;
      19890: inst = 32'h10408000;
      19891: inst = 32'hc404e32;
      19892: inst = 32'h8220000;
      19893: inst = 32'h10408000;
      19894: inst = 32'hc404e33;
      19895: inst = 32'h8220000;
      19896: inst = 32'h10408000;
      19897: inst = 32'hc404e34;
      19898: inst = 32'h8220000;
      19899: inst = 32'h10408000;
      19900: inst = 32'hc404e35;
      19901: inst = 32'h8220000;
      19902: inst = 32'h10408000;
      19903: inst = 32'hc404e38;
      19904: inst = 32'h8220000;
      19905: inst = 32'h10408000;
      19906: inst = 32'hc404e39;
      19907: inst = 32'h8220000;
      19908: inst = 32'h10408000;
      19909: inst = 32'hc404e3a;
      19910: inst = 32'h8220000;
      19911: inst = 32'h10408000;
      19912: inst = 32'hc404e3b;
      19913: inst = 32'h8220000;
      19914: inst = 32'h10408000;
      19915: inst = 32'hc404e3c;
      19916: inst = 32'h8220000;
      19917: inst = 32'h10408000;
      19918: inst = 32'hc404e3d;
      19919: inst = 32'h8220000;
      19920: inst = 32'h10408000;
      19921: inst = 32'hc404e3e;
      19922: inst = 32'h8220000;
      19923: inst = 32'h10408000;
      19924: inst = 32'hc404e3f;
      19925: inst = 32'h8220000;
      19926: inst = 32'h10408000;
      19927: inst = 32'hc404e40;
      19928: inst = 32'h8220000;
      19929: inst = 32'h10408000;
      19930: inst = 32'hc404e41;
      19931: inst = 32'h8220000;
      19932: inst = 32'h10408000;
      19933: inst = 32'hc404e42;
      19934: inst = 32'h8220000;
      19935: inst = 32'h10408000;
      19936: inst = 32'hc404e44;
      19937: inst = 32'h8220000;
      19938: inst = 32'h10408000;
      19939: inst = 32'hc404e45;
      19940: inst = 32'h8220000;
      19941: inst = 32'h10408000;
      19942: inst = 32'hc404e46;
      19943: inst = 32'h8220000;
      19944: inst = 32'h10408000;
      19945: inst = 32'hc404e47;
      19946: inst = 32'h8220000;
      19947: inst = 32'h10408000;
      19948: inst = 32'hc404e48;
      19949: inst = 32'h8220000;
      19950: inst = 32'h10408000;
      19951: inst = 32'hc404e49;
      19952: inst = 32'h8220000;
      19953: inst = 32'h10408000;
      19954: inst = 32'hc404e4a;
      19955: inst = 32'h8220000;
      19956: inst = 32'h10408000;
      19957: inst = 32'hc404e4b;
      19958: inst = 32'h8220000;
      19959: inst = 32'h10408000;
      19960: inst = 32'hc404e4c;
      19961: inst = 32'h8220000;
      19962: inst = 32'h10408000;
      19963: inst = 32'hc404e4d;
      19964: inst = 32'h8220000;
      19965: inst = 32'h10408000;
      19966: inst = 32'hc404e50;
      19967: inst = 32'h8220000;
      19968: inst = 32'h10408000;
      19969: inst = 32'hc404e51;
      19970: inst = 32'h8220000;
      19971: inst = 32'h10408000;
      19972: inst = 32'hc404e52;
      19973: inst = 32'h8220000;
      19974: inst = 32'h10408000;
      19975: inst = 32'hc404e53;
      19976: inst = 32'h8220000;
      19977: inst = 32'h10408000;
      19978: inst = 32'hc404e5c;
      19979: inst = 32'h8220000;
      19980: inst = 32'h10408000;
      19981: inst = 32'hc404e5d;
      19982: inst = 32'h8220000;
      19983: inst = 32'h10408000;
      19984: inst = 32'hc404e5e;
      19985: inst = 32'h8220000;
      19986: inst = 32'h10408000;
      19987: inst = 32'hc404e5f;
      19988: inst = 32'h8220000;
      19989: inst = 32'h10408000;
      19990: inst = 32'hc404e60;
      19991: inst = 32'h8220000;
      19992: inst = 32'h10408000;
      19993: inst = 32'hc404e61;
      19994: inst = 32'h8220000;
      19995: inst = 32'h10408000;
      19996: inst = 32'hc404e62;
      19997: inst = 32'h8220000;
      19998: inst = 32'h10408000;
      19999: inst = 32'hc404e63;
      20000: inst = 32'h8220000;
      20001: inst = 32'h10408000;
      20002: inst = 32'hc404e64;
      20003: inst = 32'h8220000;
      20004: inst = 32'h10408000;
      20005: inst = 32'hc404e65;
      20006: inst = 32'h8220000;
      20007: inst = 32'h10408000;
      20008: inst = 32'hc404e66;
      20009: inst = 32'h8220000;
      20010: inst = 32'h10408000;
      20011: inst = 32'hc404e6a;
      20012: inst = 32'h8220000;
      20013: inst = 32'h10408000;
      20014: inst = 32'hc404e6b;
      20015: inst = 32'h8220000;
      20016: inst = 32'h10408000;
      20017: inst = 32'hc404e6c;
      20018: inst = 32'h8220000;
      20019: inst = 32'h10408000;
      20020: inst = 32'hc404e6d;
      20021: inst = 32'h8220000;
      20022: inst = 32'h10408000;
      20023: inst = 32'hc404e6e;
      20024: inst = 32'h8220000;
      20025: inst = 32'h10408000;
      20026: inst = 32'hc404e6f;
      20027: inst = 32'h8220000;
      20028: inst = 32'h10408000;
      20029: inst = 32'hc404e70;
      20030: inst = 32'h8220000;
      20031: inst = 32'h10408000;
      20032: inst = 32'hc404e71;
      20033: inst = 32'h8220000;
      20034: inst = 32'h10408000;
      20035: inst = 32'hc404e72;
      20036: inst = 32'h8220000;
      20037: inst = 32'h10408000;
      20038: inst = 32'hc404e73;
      20039: inst = 32'h8220000;
      20040: inst = 32'h10408000;
      20041: inst = 32'hc404e8b;
      20042: inst = 32'h8220000;
      20043: inst = 32'h10408000;
      20044: inst = 32'hc404e8c;
      20045: inst = 32'h8220000;
      20046: inst = 32'h10408000;
      20047: inst = 32'hc404e8d;
      20048: inst = 32'h8220000;
      20049: inst = 32'h10408000;
      20050: inst = 32'hc404e99;
      20051: inst = 32'h8220000;
      20052: inst = 32'h10408000;
      20053: inst = 32'hc404e9a;
      20054: inst = 32'h8220000;
      20055: inst = 32'h10408000;
      20056: inst = 32'hc404e9b;
      20057: inst = 32'h8220000;
      20058: inst = 32'h10408000;
      20059: inst = 32'hc404e9c;
      20060: inst = 32'h8220000;
      20061: inst = 32'h10408000;
      20062: inst = 32'hc404ea4;
      20063: inst = 32'h8220000;
      20064: inst = 32'h10408000;
      20065: inst = 32'hc404ea5;
      20066: inst = 32'h8220000;
      20067: inst = 32'h10408000;
      20068: inst = 32'hc404eac;
      20069: inst = 32'h8220000;
      20070: inst = 32'h10408000;
      20071: inst = 32'hc404ead;
      20072: inst = 32'h8220000;
      20073: inst = 32'h10408000;
      20074: inst = 32'hc404eb0;
      20075: inst = 32'h8220000;
      20076: inst = 32'h10408000;
      20077: inst = 32'hc404eb1;
      20078: inst = 32'h8220000;
      20079: inst = 32'h10408000;
      20080: inst = 32'hc404eb2;
      20081: inst = 32'h8220000;
      20082: inst = 32'h10408000;
      20083: inst = 32'hc404eb3;
      20084: inst = 32'h8220000;
      20085: inst = 32'h10408000;
      20086: inst = 32'hc404eb4;
      20087: inst = 32'h8220000;
      20088: inst = 32'h10408000;
      20089: inst = 32'hc404ebc;
      20090: inst = 32'h8220000;
      20091: inst = 32'h10408000;
      20092: inst = 32'hc404ebd;
      20093: inst = 32'h8220000;
      20094: inst = 32'h10408000;
      20095: inst = 32'hc404ec2;
      20096: inst = 32'h8220000;
      20097: inst = 32'h10408000;
      20098: inst = 32'hc404ec3;
      20099: inst = 32'h8220000;
      20100: inst = 32'h10408000;
      20101: inst = 32'hc404ec4;
      20102: inst = 32'h8220000;
      20103: inst = 32'h10408000;
      20104: inst = 32'hc404ec5;
      20105: inst = 32'h8220000;
      20106: inst = 32'h10408000;
      20107: inst = 32'hc404ec9;
      20108: inst = 32'h8220000;
      20109: inst = 32'h10408000;
      20110: inst = 32'hc404eca;
      20111: inst = 32'h8220000;
      20112: inst = 32'h10408000;
      20113: inst = 32'hc404eeb;
      20114: inst = 32'h8220000;
      20115: inst = 32'h10408000;
      20116: inst = 32'hc404eec;
      20117: inst = 32'h8220000;
      20118: inst = 32'h10408000;
      20119: inst = 32'hc404efa;
      20120: inst = 32'h8220000;
      20121: inst = 32'h10408000;
      20122: inst = 32'hc404efb;
      20123: inst = 32'h8220000;
      20124: inst = 32'h10408000;
      20125: inst = 32'hc404efc;
      20126: inst = 32'h8220000;
      20127: inst = 32'h10408000;
      20128: inst = 32'hc404f04;
      20129: inst = 32'h8220000;
      20130: inst = 32'h10408000;
      20131: inst = 32'hc404f05;
      20132: inst = 32'h8220000;
      20133: inst = 32'h10408000;
      20134: inst = 32'hc404f0c;
      20135: inst = 32'h8220000;
      20136: inst = 32'h10408000;
      20137: inst = 32'hc404f0d;
      20138: inst = 32'h8220000;
      20139: inst = 32'h10408000;
      20140: inst = 32'hc404f10;
      20141: inst = 32'h8220000;
      20142: inst = 32'h10408000;
      20143: inst = 32'hc404f12;
      20144: inst = 32'h8220000;
      20145: inst = 32'h10408000;
      20146: inst = 32'hc404f13;
      20147: inst = 32'h8220000;
      20148: inst = 32'h10408000;
      20149: inst = 32'hc404f14;
      20150: inst = 32'h8220000;
      20151: inst = 32'h10408000;
      20152: inst = 32'hc404f15;
      20153: inst = 32'h8220000;
      20154: inst = 32'h10408000;
      20155: inst = 32'hc404f1c;
      20156: inst = 32'h8220000;
      20157: inst = 32'h10408000;
      20158: inst = 32'hc404f1d;
      20159: inst = 32'h8220000;
      20160: inst = 32'h10408000;
      20161: inst = 32'hc404f22;
      20162: inst = 32'h8220000;
      20163: inst = 32'h10408000;
      20164: inst = 32'hc404f23;
      20165: inst = 32'h8220000;
      20166: inst = 32'h10408000;
      20167: inst = 32'hc404f24;
      20168: inst = 32'h8220000;
      20169: inst = 32'h10408000;
      20170: inst = 32'hc404f29;
      20171: inst = 32'h8220000;
      20172: inst = 32'h10408000;
      20173: inst = 32'hc404f2a;
      20174: inst = 32'h8220000;
      20175: inst = 32'h10408000;
      20176: inst = 32'hc404f4b;
      20177: inst = 32'h8220000;
      20178: inst = 32'h10408000;
      20179: inst = 32'hc404f4c;
      20180: inst = 32'h8220000;
      20181: inst = 32'h10408000;
      20182: inst = 32'hc404f4e;
      20183: inst = 32'h8220000;
      20184: inst = 32'h10408000;
      20185: inst = 32'hc404f4f;
      20186: inst = 32'h8220000;
      20187: inst = 32'h10408000;
      20188: inst = 32'hc404f50;
      20189: inst = 32'h8220000;
      20190: inst = 32'h10408000;
      20191: inst = 32'hc404f51;
      20192: inst = 32'h8220000;
      20193: inst = 32'h10408000;
      20194: inst = 32'hc404f52;
      20195: inst = 32'h8220000;
      20196: inst = 32'h10408000;
      20197: inst = 32'hc404f5b;
      20198: inst = 32'h8220000;
      20199: inst = 32'h10408000;
      20200: inst = 32'hc404f5c;
      20201: inst = 32'h8220000;
      20202: inst = 32'h10408000;
      20203: inst = 32'hc404f5d;
      20204: inst = 32'h8220000;
      20205: inst = 32'h10408000;
      20206: inst = 32'hc404f64;
      20207: inst = 32'h8220000;
      20208: inst = 32'h10408000;
      20209: inst = 32'hc404f65;
      20210: inst = 32'h8220000;
      20211: inst = 32'h10408000;
      20212: inst = 32'hc404f6c;
      20213: inst = 32'h8220000;
      20214: inst = 32'h10408000;
      20215: inst = 32'hc404f70;
      20216: inst = 32'h8220000;
      20217: inst = 32'h10408000;
      20218: inst = 32'hc404f71;
      20219: inst = 32'h8220000;
      20220: inst = 32'h10408000;
      20221: inst = 32'hc404f72;
      20222: inst = 32'h8220000;
      20223: inst = 32'h10408000;
      20224: inst = 32'hc404f73;
      20225: inst = 32'h8220000;
      20226: inst = 32'h10408000;
      20227: inst = 32'hc404f74;
      20228: inst = 32'h8220000;
      20229: inst = 32'h10408000;
      20230: inst = 32'hc404f75;
      20231: inst = 32'h8220000;
      20232: inst = 32'h10408000;
      20233: inst = 32'hc404f76;
      20234: inst = 32'h8220000;
      20235: inst = 32'h10408000;
      20236: inst = 32'hc404f7c;
      20237: inst = 32'h8220000;
      20238: inst = 32'h10408000;
      20239: inst = 32'hc404f7d;
      20240: inst = 32'h8220000;
      20241: inst = 32'h10408000;
      20242: inst = 32'hc404f7f;
      20243: inst = 32'h8220000;
      20244: inst = 32'h10408000;
      20245: inst = 32'hc404f80;
      20246: inst = 32'h8220000;
      20247: inst = 32'h10408000;
      20248: inst = 32'hc404f81;
      20249: inst = 32'h8220000;
      20250: inst = 32'h10408000;
      20251: inst = 32'hc404f82;
      20252: inst = 32'h8220000;
      20253: inst = 32'h10408000;
      20254: inst = 32'hc404f83;
      20255: inst = 32'h8220000;
      20256: inst = 32'h10408000;
      20257: inst = 32'hc404f89;
      20258: inst = 32'h8220000;
      20259: inst = 32'h10408000;
      20260: inst = 32'hc404f8a;
      20261: inst = 32'h8220000;
      20262: inst = 32'h10408000;
      20263: inst = 32'hc404f8c;
      20264: inst = 32'h8220000;
      20265: inst = 32'h10408000;
      20266: inst = 32'hc404f8d;
      20267: inst = 32'h8220000;
      20268: inst = 32'h10408000;
      20269: inst = 32'hc404f8e;
      20270: inst = 32'h8220000;
      20271: inst = 32'h10408000;
      20272: inst = 32'hc404f8f;
      20273: inst = 32'h8220000;
      20274: inst = 32'h10408000;
      20275: inst = 32'hc404f90;
      20276: inst = 32'h8220000;
      20277: inst = 32'h10408000;
      20278: inst = 32'hc404fab;
      20279: inst = 32'h8220000;
      20280: inst = 32'h10408000;
      20281: inst = 32'hc404fac;
      20282: inst = 32'h8220000;
      20283: inst = 32'h10408000;
      20284: inst = 32'hc404fae;
      20285: inst = 32'h8220000;
      20286: inst = 32'h10408000;
      20287: inst = 32'hc404faf;
      20288: inst = 32'h8220000;
      20289: inst = 32'h10408000;
      20290: inst = 32'hc404fb0;
      20291: inst = 32'h8220000;
      20292: inst = 32'h10408000;
      20293: inst = 32'hc404fb1;
      20294: inst = 32'h8220000;
      20295: inst = 32'h10408000;
      20296: inst = 32'hc404fb2;
      20297: inst = 32'h8220000;
      20298: inst = 32'h10408000;
      20299: inst = 32'hc404fbc;
      20300: inst = 32'h8220000;
      20301: inst = 32'h10408000;
      20302: inst = 32'hc404fbd;
      20303: inst = 32'h8220000;
      20304: inst = 32'h10408000;
      20305: inst = 32'hc404fbe;
      20306: inst = 32'h8220000;
      20307: inst = 32'h10408000;
      20308: inst = 32'hc404fc4;
      20309: inst = 32'h8220000;
      20310: inst = 32'h10408000;
      20311: inst = 32'hc404fc5;
      20312: inst = 32'h8220000;
      20313: inst = 32'h10408000;
      20314: inst = 32'hc404fd0;
      20315: inst = 32'h8220000;
      20316: inst = 32'h10408000;
      20317: inst = 32'hc404fd1;
      20318: inst = 32'h8220000;
      20319: inst = 32'h10408000;
      20320: inst = 32'hc404fd2;
      20321: inst = 32'h8220000;
      20322: inst = 32'h10408000;
      20323: inst = 32'hc404fd4;
      20324: inst = 32'h8220000;
      20325: inst = 32'h10408000;
      20326: inst = 32'hc404fd5;
      20327: inst = 32'h8220000;
      20328: inst = 32'h10408000;
      20329: inst = 32'hc404fd6;
      20330: inst = 32'h8220000;
      20331: inst = 32'h10408000;
      20332: inst = 32'hc404fd7;
      20333: inst = 32'h8220000;
      20334: inst = 32'h10408000;
      20335: inst = 32'hc404fdc;
      20336: inst = 32'h8220000;
      20337: inst = 32'h10408000;
      20338: inst = 32'hc404fdd;
      20339: inst = 32'h8220000;
      20340: inst = 32'h10408000;
      20341: inst = 32'hc404fdf;
      20342: inst = 32'h8220000;
      20343: inst = 32'h10408000;
      20344: inst = 32'hc404fe0;
      20345: inst = 32'h8220000;
      20346: inst = 32'h10408000;
      20347: inst = 32'hc404fe1;
      20348: inst = 32'h8220000;
      20349: inst = 32'h10408000;
      20350: inst = 32'hc404fe2;
      20351: inst = 32'h8220000;
      20352: inst = 32'h10408000;
      20353: inst = 32'hc404fe9;
      20354: inst = 32'h8220000;
      20355: inst = 32'h10408000;
      20356: inst = 32'hc404fea;
      20357: inst = 32'h8220000;
      20358: inst = 32'h10408000;
      20359: inst = 32'hc404fec;
      20360: inst = 32'h8220000;
      20361: inst = 32'h10408000;
      20362: inst = 32'hc404fed;
      20363: inst = 32'h8220000;
      20364: inst = 32'h10408000;
      20365: inst = 32'hc404fee;
      20366: inst = 32'h8220000;
      20367: inst = 32'h10408000;
      20368: inst = 32'hc404fef;
      20369: inst = 32'h8220000;
      20370: inst = 32'h10408000;
      20371: inst = 32'hc404ff0;
      20372: inst = 32'h8220000;
      20373: inst = 32'h10408000;
      20374: inst = 32'hc40500b;
      20375: inst = 32'h8220000;
      20376: inst = 32'h10408000;
      20377: inst = 32'hc40500c;
      20378: inst = 32'h8220000;
      20379: inst = 32'h10408000;
      20380: inst = 32'hc40501d;
      20381: inst = 32'h8220000;
      20382: inst = 32'h10408000;
      20383: inst = 32'hc40501e;
      20384: inst = 32'h8220000;
      20385: inst = 32'h10408000;
      20386: inst = 32'hc40501f;
      20387: inst = 32'h8220000;
      20388: inst = 32'h10408000;
      20389: inst = 32'hc405024;
      20390: inst = 32'h8220000;
      20391: inst = 32'h10408000;
      20392: inst = 32'hc405025;
      20393: inst = 32'h8220000;
      20394: inst = 32'h10408000;
      20395: inst = 32'hc405030;
      20396: inst = 32'h8220000;
      20397: inst = 32'h10408000;
      20398: inst = 32'hc405031;
      20399: inst = 32'h8220000;
      20400: inst = 32'h10408000;
      20401: inst = 32'hc405032;
      20402: inst = 32'h8220000;
      20403: inst = 32'h10408000;
      20404: inst = 32'hc405033;
      20405: inst = 32'h8220000;
      20406: inst = 32'h10408000;
      20407: inst = 32'hc405034;
      20408: inst = 32'h8220000;
      20409: inst = 32'h10408000;
      20410: inst = 32'hc405035;
      20411: inst = 32'h8220000;
      20412: inst = 32'h10408000;
      20413: inst = 32'hc405036;
      20414: inst = 32'h8220000;
      20415: inst = 32'h10408000;
      20416: inst = 32'hc405037;
      20417: inst = 32'h8220000;
      20418: inst = 32'h10408000;
      20419: inst = 32'hc405038;
      20420: inst = 32'h8220000;
      20421: inst = 32'h10408000;
      20422: inst = 32'hc40503c;
      20423: inst = 32'h8220000;
      20424: inst = 32'h10408000;
      20425: inst = 32'hc40503d;
      20426: inst = 32'h8220000;
      20427: inst = 32'h10408000;
      20428: inst = 32'hc405049;
      20429: inst = 32'h8220000;
      20430: inst = 32'h10408000;
      20431: inst = 32'hc40504a;
      20432: inst = 32'h8220000;
      20433: inst = 32'h10408000;
      20434: inst = 32'hc40506b;
      20435: inst = 32'h8220000;
      20436: inst = 32'h10408000;
      20437: inst = 32'hc40506c;
      20438: inst = 32'h8220000;
      20439: inst = 32'h10408000;
      20440: inst = 32'hc40506d;
      20441: inst = 32'h8220000;
      20442: inst = 32'h10408000;
      20443: inst = 32'hc40506e;
      20444: inst = 32'h8220000;
      20445: inst = 32'h10408000;
      20446: inst = 32'hc40506f;
      20447: inst = 32'h8220000;
      20448: inst = 32'h10408000;
      20449: inst = 32'hc405070;
      20450: inst = 32'h8220000;
      20451: inst = 32'h10408000;
      20452: inst = 32'hc405071;
      20453: inst = 32'h8220000;
      20454: inst = 32'h10408000;
      20455: inst = 32'hc405072;
      20456: inst = 32'h8220000;
      20457: inst = 32'h10408000;
      20458: inst = 32'hc405073;
      20459: inst = 32'h8220000;
      20460: inst = 32'h10408000;
      20461: inst = 32'hc405074;
      20462: inst = 32'h8220000;
      20463: inst = 32'h10408000;
      20464: inst = 32'hc405075;
      20465: inst = 32'h8220000;
      20466: inst = 32'h10408000;
      20467: inst = 32'hc405077;
      20468: inst = 32'h8220000;
      20469: inst = 32'h10408000;
      20470: inst = 32'hc405078;
      20471: inst = 32'h8220000;
      20472: inst = 32'h10408000;
      20473: inst = 32'hc405079;
      20474: inst = 32'h8220000;
      20475: inst = 32'h10408000;
      20476: inst = 32'hc40507a;
      20477: inst = 32'h8220000;
      20478: inst = 32'h10408000;
      20479: inst = 32'hc40507b;
      20480: inst = 32'h8220000;
      20481: inst = 32'h10408000;
      20482: inst = 32'hc40507c;
      20483: inst = 32'h8220000;
      20484: inst = 32'h10408000;
      20485: inst = 32'hc40507d;
      20486: inst = 32'h8220000;
      20487: inst = 32'h10408000;
      20488: inst = 32'hc40507e;
      20489: inst = 32'h8220000;
      20490: inst = 32'h10408000;
      20491: inst = 32'hc40507f;
      20492: inst = 32'h8220000;
      20493: inst = 32'h10408000;
      20494: inst = 32'hc405080;
      20495: inst = 32'h8220000;
      20496: inst = 32'h10408000;
      20497: inst = 32'hc405084;
      20498: inst = 32'h8220000;
      20499: inst = 32'h10408000;
      20500: inst = 32'hc405085;
      20501: inst = 32'h8220000;
      20502: inst = 32'h10408000;
      20503: inst = 32'hc405086;
      20504: inst = 32'h8220000;
      20505: inst = 32'h10408000;
      20506: inst = 32'hc405087;
      20507: inst = 32'h8220000;
      20508: inst = 32'h10408000;
      20509: inst = 32'hc405088;
      20510: inst = 32'h8220000;
      20511: inst = 32'h10408000;
      20512: inst = 32'hc405089;
      20513: inst = 32'h8220000;
      20514: inst = 32'h10408000;
      20515: inst = 32'hc40508a;
      20516: inst = 32'h8220000;
      20517: inst = 32'h10408000;
      20518: inst = 32'hc40508b;
      20519: inst = 32'h8220000;
      20520: inst = 32'h10408000;
      20521: inst = 32'hc40508c;
      20522: inst = 32'h8220000;
      20523: inst = 32'h10408000;
      20524: inst = 32'hc40508d;
      20525: inst = 32'h8220000;
      20526: inst = 32'h10408000;
      20527: inst = 32'hc405090;
      20528: inst = 32'h8220000;
      20529: inst = 32'h10408000;
      20530: inst = 32'hc405091;
      20531: inst = 32'h8220000;
      20532: inst = 32'h10408000;
      20533: inst = 32'hc405096;
      20534: inst = 32'h8220000;
      20535: inst = 32'h10408000;
      20536: inst = 32'hc405097;
      20537: inst = 32'h8220000;
      20538: inst = 32'h10408000;
      20539: inst = 32'hc405098;
      20540: inst = 32'h8220000;
      20541: inst = 32'h10408000;
      20542: inst = 32'hc405099;
      20543: inst = 32'h8220000;
      20544: inst = 32'h10408000;
      20545: inst = 32'hc40509c;
      20546: inst = 32'h8220000;
      20547: inst = 32'h10408000;
      20548: inst = 32'hc40509d;
      20549: inst = 32'h8220000;
      20550: inst = 32'h10408000;
      20551: inst = 32'hc4050a9;
      20552: inst = 32'h8220000;
      20553: inst = 32'h10408000;
      20554: inst = 32'hc4050aa;
      20555: inst = 32'h8220000;
      20556: inst = 32'h10408000;
      20557: inst = 32'hc4050ab;
      20558: inst = 32'h8220000;
      20559: inst = 32'h10408000;
      20560: inst = 32'hc4050ac;
      20561: inst = 32'h8220000;
      20562: inst = 32'h10408000;
      20563: inst = 32'hc4050ad;
      20564: inst = 32'h8220000;
      20565: inst = 32'h10408000;
      20566: inst = 32'hc4050ae;
      20567: inst = 32'h8220000;
      20568: inst = 32'h10408000;
      20569: inst = 32'hc4050af;
      20570: inst = 32'h8220000;
      20571: inst = 32'h10408000;
      20572: inst = 32'hc4050b0;
      20573: inst = 32'h8220000;
      20574: inst = 32'h10408000;
      20575: inst = 32'hc4050b1;
      20576: inst = 32'h8220000;
      20577: inst = 32'h10408000;
      20578: inst = 32'hc4050b2;
      20579: inst = 32'h8220000;
      20580: inst = 32'h10408000;
      20581: inst = 32'hc4050b3;
      20582: inst = 32'h8220000;
      20583: inst = 32'h10408000;
      20584: inst = 32'hc4050cb;
      20585: inst = 32'h8220000;
      20586: inst = 32'h10408000;
      20587: inst = 32'hc4050cc;
      20588: inst = 32'h8220000;
      20589: inst = 32'h10408000;
      20590: inst = 32'hc4050cd;
      20591: inst = 32'h8220000;
      20592: inst = 32'h10408000;
      20593: inst = 32'hc4050ce;
      20594: inst = 32'h8220000;
      20595: inst = 32'h10408000;
      20596: inst = 32'hc4050cf;
      20597: inst = 32'h8220000;
      20598: inst = 32'h10408000;
      20599: inst = 32'hc4050d0;
      20600: inst = 32'h8220000;
      20601: inst = 32'h10408000;
      20602: inst = 32'hc4050d1;
      20603: inst = 32'h8220000;
      20604: inst = 32'h10408000;
      20605: inst = 32'hc4050d2;
      20606: inst = 32'h8220000;
      20607: inst = 32'h10408000;
      20608: inst = 32'hc4050d3;
      20609: inst = 32'h8220000;
      20610: inst = 32'h10408000;
      20611: inst = 32'hc4050d4;
      20612: inst = 32'h8220000;
      20613: inst = 32'h10408000;
      20614: inst = 32'hc4050d7;
      20615: inst = 32'h8220000;
      20616: inst = 32'h10408000;
      20617: inst = 32'hc4050d8;
      20618: inst = 32'h8220000;
      20619: inst = 32'h10408000;
      20620: inst = 32'hc4050d9;
      20621: inst = 32'h8220000;
      20622: inst = 32'h10408000;
      20623: inst = 32'hc4050da;
      20624: inst = 32'h8220000;
      20625: inst = 32'h10408000;
      20626: inst = 32'hc4050db;
      20627: inst = 32'h8220000;
      20628: inst = 32'h10408000;
      20629: inst = 32'hc4050dc;
      20630: inst = 32'h8220000;
      20631: inst = 32'h10408000;
      20632: inst = 32'hc4050dd;
      20633: inst = 32'h8220000;
      20634: inst = 32'h10408000;
      20635: inst = 32'hc4050de;
      20636: inst = 32'h8220000;
      20637: inst = 32'h10408000;
      20638: inst = 32'hc4050df;
      20639: inst = 32'h8220000;
      20640: inst = 32'h10408000;
      20641: inst = 32'hc4050e0;
      20642: inst = 32'h8220000;
      20643: inst = 32'h10408000;
      20644: inst = 32'hc4050e1;
      20645: inst = 32'h8220000;
      20646: inst = 32'h10408000;
      20647: inst = 32'hc4050e5;
      20648: inst = 32'h8220000;
      20649: inst = 32'h10408000;
      20650: inst = 32'hc4050e6;
      20651: inst = 32'h8220000;
      20652: inst = 32'h10408000;
      20653: inst = 32'hc4050e7;
      20654: inst = 32'h8220000;
      20655: inst = 32'h10408000;
      20656: inst = 32'hc4050e8;
      20657: inst = 32'h8220000;
      20658: inst = 32'h10408000;
      20659: inst = 32'hc4050e9;
      20660: inst = 32'h8220000;
      20661: inst = 32'h10408000;
      20662: inst = 32'hc4050ea;
      20663: inst = 32'h8220000;
      20664: inst = 32'h10408000;
      20665: inst = 32'hc4050eb;
      20666: inst = 32'h8220000;
      20667: inst = 32'h10408000;
      20668: inst = 32'hc4050ec;
      20669: inst = 32'h8220000;
      20670: inst = 32'h10408000;
      20671: inst = 32'hc4050ed;
      20672: inst = 32'h8220000;
      20673: inst = 32'h10408000;
      20674: inst = 32'hc4050f0;
      20675: inst = 32'h8220000;
      20676: inst = 32'h10408000;
      20677: inst = 32'hc4050f1;
      20678: inst = 32'h8220000;
      20679: inst = 32'h10408000;
      20680: inst = 32'hc4050f6;
      20681: inst = 32'h8220000;
      20682: inst = 32'h10408000;
      20683: inst = 32'hc4050f7;
      20684: inst = 32'h8220000;
      20685: inst = 32'h10408000;
      20686: inst = 32'hc4050f8;
      20687: inst = 32'h8220000;
      20688: inst = 32'h10408000;
      20689: inst = 32'hc4050f9;
      20690: inst = 32'h8220000;
      20691: inst = 32'h10408000;
      20692: inst = 32'hc4050fa;
      20693: inst = 32'h8220000;
      20694: inst = 32'h10408000;
      20695: inst = 32'hc4050fc;
      20696: inst = 32'h8220000;
      20697: inst = 32'h10408000;
      20698: inst = 32'hc4050fd;
      20699: inst = 32'h8220000;
      20700: inst = 32'h10408000;
      20701: inst = 32'hc405109;
      20702: inst = 32'h8220000;
      20703: inst = 32'h10408000;
      20704: inst = 32'hc40510a;
      20705: inst = 32'h8220000;
      20706: inst = 32'h10408000;
      20707: inst = 32'hc40510b;
      20708: inst = 32'h8220000;
      20709: inst = 32'h10408000;
      20710: inst = 32'hc40510c;
      20711: inst = 32'h8220000;
      20712: inst = 32'h10408000;
      20713: inst = 32'hc40510d;
      20714: inst = 32'h8220000;
      20715: inst = 32'h10408000;
      20716: inst = 32'hc40510e;
      20717: inst = 32'h8220000;
      20718: inst = 32'h10408000;
      20719: inst = 32'hc40510f;
      20720: inst = 32'h8220000;
      20721: inst = 32'h10408000;
      20722: inst = 32'hc405110;
      20723: inst = 32'h8220000;
      20724: inst = 32'h10408000;
      20725: inst = 32'hc405111;
      20726: inst = 32'h8220000;
      20727: inst = 32'h10408000;
      20728: inst = 32'hc405112;
      20729: inst = 32'h8220000;
      20730: inst = 32'h10408000;
      20731: inst = 32'hc405113;
      20732: inst = 32'h8220000;
      20733: inst = 32'h58000000;
      20734: inst = 32'hc20529c;
      20735: inst = 32'h10408000;
      20736: inst = 32'hc404224;
      20737: inst = 32'h8220000;
      20738: inst = 32'h10408000;
      20739: inst = 32'hc404225;
      20740: inst = 32'h8220000;
      20741: inst = 32'h10408000;
      20742: inst = 32'hc404226;
      20743: inst = 32'h8220000;
      20744: inst = 32'h10408000;
      20745: inst = 32'hc404227;
      20746: inst = 32'h8220000;
      20747: inst = 32'h10408000;
      20748: inst = 32'hc404228;
      20749: inst = 32'h8220000;
      20750: inst = 32'h10408000;
      20751: inst = 32'hc404229;
      20752: inst = 32'h8220000;
      20753: inst = 32'h10408000;
      20754: inst = 32'hc40422a;
      20755: inst = 32'h8220000;
      20756: inst = 32'h10408000;
      20757: inst = 32'hc40422b;
      20758: inst = 32'h8220000;
      20759: inst = 32'h10408000;
      20760: inst = 32'hc40422c;
      20761: inst = 32'h8220000;
      20762: inst = 32'h10408000;
      20763: inst = 32'hc40422d;
      20764: inst = 32'h8220000;
      20765: inst = 32'h10408000;
      20766: inst = 32'hc40422e;
      20767: inst = 32'h8220000;
      20768: inst = 32'h10408000;
      20769: inst = 32'hc40422f;
      20770: inst = 32'h8220000;
      20771: inst = 32'h10408000;
      20772: inst = 32'hc404230;
      20773: inst = 32'h8220000;
      20774: inst = 32'h10408000;
      20775: inst = 32'hc404231;
      20776: inst = 32'h8220000;
      20777: inst = 32'h10408000;
      20778: inst = 32'hc404232;
      20779: inst = 32'h8220000;
      20780: inst = 32'h10408000;
      20781: inst = 32'hc404233;
      20782: inst = 32'h8220000;
      20783: inst = 32'h10408000;
      20784: inst = 32'hc404234;
      20785: inst = 32'h8220000;
      20786: inst = 32'h10408000;
      20787: inst = 32'hc404235;
      20788: inst = 32'h8220000;
      20789: inst = 32'h10408000;
      20790: inst = 32'hc404236;
      20791: inst = 32'h8220000;
      20792: inst = 32'h10408000;
      20793: inst = 32'hc404237;
      20794: inst = 32'h8220000;
      20795: inst = 32'h10408000;
      20796: inst = 32'hc404238;
      20797: inst = 32'h8220000;
      20798: inst = 32'h10408000;
      20799: inst = 32'hc404239;
      20800: inst = 32'h8220000;
      20801: inst = 32'h10408000;
      20802: inst = 32'hc40423a;
      20803: inst = 32'h8220000;
      20804: inst = 32'h10408000;
      20805: inst = 32'hc40423b;
      20806: inst = 32'h8220000;
      20807: inst = 32'h10408000;
      20808: inst = 32'hc40423c;
      20809: inst = 32'h8220000;
      20810: inst = 32'h10408000;
      20811: inst = 32'hc40423d;
      20812: inst = 32'h8220000;
      20813: inst = 32'h10408000;
      20814: inst = 32'hc40423e;
      20815: inst = 32'h8220000;
      20816: inst = 32'h10408000;
      20817: inst = 32'hc40423f;
      20818: inst = 32'h8220000;
      20819: inst = 32'h10408000;
      20820: inst = 32'hc404240;
      20821: inst = 32'h8220000;
      20822: inst = 32'h10408000;
      20823: inst = 32'hc404241;
      20824: inst = 32'h8220000;
      20825: inst = 32'h10408000;
      20826: inst = 32'hc404242;
      20827: inst = 32'h8220000;
      20828: inst = 32'h10408000;
      20829: inst = 32'hc404243;
      20830: inst = 32'h8220000;
      20831: inst = 32'h10408000;
      20832: inst = 32'hc404244;
      20833: inst = 32'h8220000;
      20834: inst = 32'h10408000;
      20835: inst = 32'hc404245;
      20836: inst = 32'h8220000;
      20837: inst = 32'h10408000;
      20838: inst = 32'hc404246;
      20839: inst = 32'h8220000;
      20840: inst = 32'h10408000;
      20841: inst = 32'hc404247;
      20842: inst = 32'h8220000;
      20843: inst = 32'h10408000;
      20844: inst = 32'hc404248;
      20845: inst = 32'h8220000;
      20846: inst = 32'h10408000;
      20847: inst = 32'hc404249;
      20848: inst = 32'h8220000;
      20849: inst = 32'h10408000;
      20850: inst = 32'hc40424a;
      20851: inst = 32'h8220000;
      20852: inst = 32'h10408000;
      20853: inst = 32'hc40424b;
      20854: inst = 32'h8220000;
      20855: inst = 32'h10408000;
      20856: inst = 32'hc40424c;
      20857: inst = 32'h8220000;
      20858: inst = 32'h10408000;
      20859: inst = 32'hc40424d;
      20860: inst = 32'h8220000;
      20861: inst = 32'h10408000;
      20862: inst = 32'hc40424e;
      20863: inst = 32'h8220000;
      20864: inst = 32'h10408000;
      20865: inst = 32'hc40424f;
      20866: inst = 32'h8220000;
      20867: inst = 32'h10408000;
      20868: inst = 32'hc404250;
      20869: inst = 32'h8220000;
      20870: inst = 32'h10408000;
      20871: inst = 32'hc404251;
      20872: inst = 32'h8220000;
      20873: inst = 32'h10408000;
      20874: inst = 32'hc404252;
      20875: inst = 32'h8220000;
      20876: inst = 32'h10408000;
      20877: inst = 32'hc404253;
      20878: inst = 32'h8220000;
      20879: inst = 32'h10408000;
      20880: inst = 32'hc404254;
      20881: inst = 32'h8220000;
      20882: inst = 32'h10408000;
      20883: inst = 32'hc404255;
      20884: inst = 32'h8220000;
      20885: inst = 32'h10408000;
      20886: inst = 32'hc404256;
      20887: inst = 32'h8220000;
      20888: inst = 32'h10408000;
      20889: inst = 32'hc404257;
      20890: inst = 32'h8220000;
      20891: inst = 32'h10408000;
      20892: inst = 32'hc404258;
      20893: inst = 32'h8220000;
      20894: inst = 32'h10408000;
      20895: inst = 32'hc404259;
      20896: inst = 32'h8220000;
      20897: inst = 32'h10408000;
      20898: inst = 32'hc40425a;
      20899: inst = 32'h8220000;
      20900: inst = 32'h10408000;
      20901: inst = 32'hc40425b;
      20902: inst = 32'h8220000;
      20903: inst = 32'h10408000;
      20904: inst = 32'hc40425c;
      20905: inst = 32'h8220000;
      20906: inst = 32'h10408000;
      20907: inst = 32'hc40425d;
      20908: inst = 32'h8220000;
      20909: inst = 32'h10408000;
      20910: inst = 32'hc40425e;
      20911: inst = 32'h8220000;
      20912: inst = 32'h10408000;
      20913: inst = 32'hc40425f;
      20914: inst = 32'h8220000;
      20915: inst = 32'h10408000;
      20916: inst = 32'hc404260;
      20917: inst = 32'h8220000;
      20918: inst = 32'h10408000;
      20919: inst = 32'hc404261;
      20920: inst = 32'h8220000;
      20921: inst = 32'h10408000;
      20922: inst = 32'hc404262;
      20923: inst = 32'h8220000;
      20924: inst = 32'h10408000;
      20925: inst = 32'hc404263;
      20926: inst = 32'h8220000;
      20927: inst = 32'h10408000;
      20928: inst = 32'hc404264;
      20929: inst = 32'h8220000;
      20930: inst = 32'h10408000;
      20931: inst = 32'hc404265;
      20932: inst = 32'h8220000;
      20933: inst = 32'h10408000;
      20934: inst = 32'hc404266;
      20935: inst = 32'h8220000;
      20936: inst = 32'h10408000;
      20937: inst = 32'hc404267;
      20938: inst = 32'h8220000;
      20939: inst = 32'h10408000;
      20940: inst = 32'hc404268;
      20941: inst = 32'h8220000;
      20942: inst = 32'h10408000;
      20943: inst = 32'hc404269;
      20944: inst = 32'h8220000;
      20945: inst = 32'h10408000;
      20946: inst = 32'hc40426a;
      20947: inst = 32'h8220000;
      20948: inst = 32'h10408000;
      20949: inst = 32'hc40426b;
      20950: inst = 32'h8220000;
      20951: inst = 32'h10408000;
      20952: inst = 32'hc40426c;
      20953: inst = 32'h8220000;
      20954: inst = 32'h10408000;
      20955: inst = 32'hc40426d;
      20956: inst = 32'h8220000;
      20957: inst = 32'h10408000;
      20958: inst = 32'hc40426e;
      20959: inst = 32'h8220000;
      20960: inst = 32'h10408000;
      20961: inst = 32'hc40426f;
      20962: inst = 32'h8220000;
      20963: inst = 32'h10408000;
      20964: inst = 32'hc404270;
      20965: inst = 32'h8220000;
      20966: inst = 32'h10408000;
      20967: inst = 32'hc404271;
      20968: inst = 32'h8220000;
      20969: inst = 32'h10408000;
      20970: inst = 32'hc404272;
      20971: inst = 32'h8220000;
      20972: inst = 32'h10408000;
      20973: inst = 32'hc404273;
      20974: inst = 32'h8220000;
      20975: inst = 32'h10408000;
      20976: inst = 32'hc404274;
      20977: inst = 32'h8220000;
      20978: inst = 32'h10408000;
      20979: inst = 32'hc404275;
      20980: inst = 32'h8220000;
      20981: inst = 32'h10408000;
      20982: inst = 32'hc404276;
      20983: inst = 32'h8220000;
      20984: inst = 32'h10408000;
      20985: inst = 32'hc404277;
      20986: inst = 32'h8220000;
      20987: inst = 32'h10408000;
      20988: inst = 32'hc404278;
      20989: inst = 32'h8220000;
      20990: inst = 32'h10408000;
      20991: inst = 32'hc404279;
      20992: inst = 32'h8220000;
      20993: inst = 32'h10408000;
      20994: inst = 32'hc40427a;
      20995: inst = 32'h8220000;
      20996: inst = 32'h10408000;
      20997: inst = 32'hc40427b;
      20998: inst = 32'h8220000;
      20999: inst = 32'h10408000;
      21000: inst = 32'hc404284;
      21001: inst = 32'h8220000;
      21002: inst = 32'h10408000;
      21003: inst = 32'hc404285;
      21004: inst = 32'h8220000;
      21005: inst = 32'h10408000;
      21006: inst = 32'hc404286;
      21007: inst = 32'h8220000;
      21008: inst = 32'h10408000;
      21009: inst = 32'hc404287;
      21010: inst = 32'h8220000;
      21011: inst = 32'h10408000;
      21012: inst = 32'hc404288;
      21013: inst = 32'h8220000;
      21014: inst = 32'h10408000;
      21015: inst = 32'hc404289;
      21016: inst = 32'h8220000;
      21017: inst = 32'h10408000;
      21018: inst = 32'hc40428a;
      21019: inst = 32'h8220000;
      21020: inst = 32'h10408000;
      21021: inst = 32'hc40428b;
      21022: inst = 32'h8220000;
      21023: inst = 32'h10408000;
      21024: inst = 32'hc40428c;
      21025: inst = 32'h8220000;
      21026: inst = 32'h10408000;
      21027: inst = 32'hc40428d;
      21028: inst = 32'h8220000;
      21029: inst = 32'h10408000;
      21030: inst = 32'hc40428e;
      21031: inst = 32'h8220000;
      21032: inst = 32'h10408000;
      21033: inst = 32'hc40428f;
      21034: inst = 32'h8220000;
      21035: inst = 32'h10408000;
      21036: inst = 32'hc404290;
      21037: inst = 32'h8220000;
      21038: inst = 32'h10408000;
      21039: inst = 32'hc404291;
      21040: inst = 32'h8220000;
      21041: inst = 32'h10408000;
      21042: inst = 32'hc404292;
      21043: inst = 32'h8220000;
      21044: inst = 32'h10408000;
      21045: inst = 32'hc404293;
      21046: inst = 32'h8220000;
      21047: inst = 32'h10408000;
      21048: inst = 32'hc404294;
      21049: inst = 32'h8220000;
      21050: inst = 32'h10408000;
      21051: inst = 32'hc404295;
      21052: inst = 32'h8220000;
      21053: inst = 32'h10408000;
      21054: inst = 32'hc404296;
      21055: inst = 32'h8220000;
      21056: inst = 32'h10408000;
      21057: inst = 32'hc404297;
      21058: inst = 32'h8220000;
      21059: inst = 32'h10408000;
      21060: inst = 32'hc404298;
      21061: inst = 32'h8220000;
      21062: inst = 32'h10408000;
      21063: inst = 32'hc404299;
      21064: inst = 32'h8220000;
      21065: inst = 32'h10408000;
      21066: inst = 32'hc40429a;
      21067: inst = 32'h8220000;
      21068: inst = 32'h10408000;
      21069: inst = 32'hc40429b;
      21070: inst = 32'h8220000;
      21071: inst = 32'h10408000;
      21072: inst = 32'hc40429c;
      21073: inst = 32'h8220000;
      21074: inst = 32'h10408000;
      21075: inst = 32'hc40429d;
      21076: inst = 32'h8220000;
      21077: inst = 32'h10408000;
      21078: inst = 32'hc40429e;
      21079: inst = 32'h8220000;
      21080: inst = 32'h10408000;
      21081: inst = 32'hc40429f;
      21082: inst = 32'h8220000;
      21083: inst = 32'h10408000;
      21084: inst = 32'hc4042a0;
      21085: inst = 32'h8220000;
      21086: inst = 32'h10408000;
      21087: inst = 32'hc4042a1;
      21088: inst = 32'h8220000;
      21089: inst = 32'h10408000;
      21090: inst = 32'hc4042a2;
      21091: inst = 32'h8220000;
      21092: inst = 32'h10408000;
      21093: inst = 32'hc4042a3;
      21094: inst = 32'h8220000;
      21095: inst = 32'h10408000;
      21096: inst = 32'hc4042a4;
      21097: inst = 32'h8220000;
      21098: inst = 32'h10408000;
      21099: inst = 32'hc4042a5;
      21100: inst = 32'h8220000;
      21101: inst = 32'h10408000;
      21102: inst = 32'hc4042a6;
      21103: inst = 32'h8220000;
      21104: inst = 32'h10408000;
      21105: inst = 32'hc4042a7;
      21106: inst = 32'h8220000;
      21107: inst = 32'h10408000;
      21108: inst = 32'hc4042a8;
      21109: inst = 32'h8220000;
      21110: inst = 32'h10408000;
      21111: inst = 32'hc4042a9;
      21112: inst = 32'h8220000;
      21113: inst = 32'h10408000;
      21114: inst = 32'hc4042aa;
      21115: inst = 32'h8220000;
      21116: inst = 32'h10408000;
      21117: inst = 32'hc4042ab;
      21118: inst = 32'h8220000;
      21119: inst = 32'h10408000;
      21120: inst = 32'hc4042ac;
      21121: inst = 32'h8220000;
      21122: inst = 32'h10408000;
      21123: inst = 32'hc4042ad;
      21124: inst = 32'h8220000;
      21125: inst = 32'h10408000;
      21126: inst = 32'hc4042ae;
      21127: inst = 32'h8220000;
      21128: inst = 32'h10408000;
      21129: inst = 32'hc4042af;
      21130: inst = 32'h8220000;
      21131: inst = 32'h10408000;
      21132: inst = 32'hc4042b0;
      21133: inst = 32'h8220000;
      21134: inst = 32'h10408000;
      21135: inst = 32'hc4042b1;
      21136: inst = 32'h8220000;
      21137: inst = 32'h10408000;
      21138: inst = 32'hc4042b2;
      21139: inst = 32'h8220000;
      21140: inst = 32'h10408000;
      21141: inst = 32'hc4042b3;
      21142: inst = 32'h8220000;
      21143: inst = 32'h10408000;
      21144: inst = 32'hc4042b4;
      21145: inst = 32'h8220000;
      21146: inst = 32'h10408000;
      21147: inst = 32'hc4042b5;
      21148: inst = 32'h8220000;
      21149: inst = 32'h10408000;
      21150: inst = 32'hc4042b6;
      21151: inst = 32'h8220000;
      21152: inst = 32'h10408000;
      21153: inst = 32'hc4042b7;
      21154: inst = 32'h8220000;
      21155: inst = 32'h10408000;
      21156: inst = 32'hc4042b8;
      21157: inst = 32'h8220000;
      21158: inst = 32'h10408000;
      21159: inst = 32'hc4042b9;
      21160: inst = 32'h8220000;
      21161: inst = 32'h10408000;
      21162: inst = 32'hc4042ba;
      21163: inst = 32'h8220000;
      21164: inst = 32'h10408000;
      21165: inst = 32'hc4042bb;
      21166: inst = 32'h8220000;
      21167: inst = 32'h10408000;
      21168: inst = 32'hc4042bc;
      21169: inst = 32'h8220000;
      21170: inst = 32'h10408000;
      21171: inst = 32'hc4042bd;
      21172: inst = 32'h8220000;
      21173: inst = 32'h10408000;
      21174: inst = 32'hc4042be;
      21175: inst = 32'h8220000;
      21176: inst = 32'h10408000;
      21177: inst = 32'hc4042bf;
      21178: inst = 32'h8220000;
      21179: inst = 32'h10408000;
      21180: inst = 32'hc4042c0;
      21181: inst = 32'h8220000;
      21182: inst = 32'h10408000;
      21183: inst = 32'hc4042c1;
      21184: inst = 32'h8220000;
      21185: inst = 32'h10408000;
      21186: inst = 32'hc4042c2;
      21187: inst = 32'h8220000;
      21188: inst = 32'h10408000;
      21189: inst = 32'hc4042c3;
      21190: inst = 32'h8220000;
      21191: inst = 32'h10408000;
      21192: inst = 32'hc4042c4;
      21193: inst = 32'h8220000;
      21194: inst = 32'h10408000;
      21195: inst = 32'hc4042c5;
      21196: inst = 32'h8220000;
      21197: inst = 32'h10408000;
      21198: inst = 32'hc4042c6;
      21199: inst = 32'h8220000;
      21200: inst = 32'h10408000;
      21201: inst = 32'hc4042c7;
      21202: inst = 32'h8220000;
      21203: inst = 32'h10408000;
      21204: inst = 32'hc4042c8;
      21205: inst = 32'h8220000;
      21206: inst = 32'h10408000;
      21207: inst = 32'hc4042c9;
      21208: inst = 32'h8220000;
      21209: inst = 32'h10408000;
      21210: inst = 32'hc4042ca;
      21211: inst = 32'h8220000;
      21212: inst = 32'h10408000;
      21213: inst = 32'hc4042cb;
      21214: inst = 32'h8220000;
      21215: inst = 32'h10408000;
      21216: inst = 32'hc4042cc;
      21217: inst = 32'h8220000;
      21218: inst = 32'h10408000;
      21219: inst = 32'hc4042cd;
      21220: inst = 32'h8220000;
      21221: inst = 32'h10408000;
      21222: inst = 32'hc4042ce;
      21223: inst = 32'h8220000;
      21224: inst = 32'h10408000;
      21225: inst = 32'hc4042cf;
      21226: inst = 32'h8220000;
      21227: inst = 32'h10408000;
      21228: inst = 32'hc4042d0;
      21229: inst = 32'h8220000;
      21230: inst = 32'h10408000;
      21231: inst = 32'hc4042d1;
      21232: inst = 32'h8220000;
      21233: inst = 32'h10408000;
      21234: inst = 32'hc4042d2;
      21235: inst = 32'h8220000;
      21236: inst = 32'h10408000;
      21237: inst = 32'hc4042d3;
      21238: inst = 32'h8220000;
      21239: inst = 32'h10408000;
      21240: inst = 32'hc4042d4;
      21241: inst = 32'h8220000;
      21242: inst = 32'h10408000;
      21243: inst = 32'hc4042d5;
      21244: inst = 32'h8220000;
      21245: inst = 32'h10408000;
      21246: inst = 32'hc4042d6;
      21247: inst = 32'h8220000;
      21248: inst = 32'h10408000;
      21249: inst = 32'hc4042d7;
      21250: inst = 32'h8220000;
      21251: inst = 32'h10408000;
      21252: inst = 32'hc4042d8;
      21253: inst = 32'h8220000;
      21254: inst = 32'h10408000;
      21255: inst = 32'hc4042d9;
      21256: inst = 32'h8220000;
      21257: inst = 32'h10408000;
      21258: inst = 32'hc4042da;
      21259: inst = 32'h8220000;
      21260: inst = 32'h10408000;
      21261: inst = 32'hc4042db;
      21262: inst = 32'h8220000;
      21263: inst = 32'h10408000;
      21264: inst = 32'hc4042e4;
      21265: inst = 32'h8220000;
      21266: inst = 32'h10408000;
      21267: inst = 32'hc4042e5;
      21268: inst = 32'h8220000;
      21269: inst = 32'h10408000;
      21270: inst = 32'hc4042e6;
      21271: inst = 32'h8220000;
      21272: inst = 32'h10408000;
      21273: inst = 32'hc404339;
      21274: inst = 32'h8220000;
      21275: inst = 32'h10408000;
      21276: inst = 32'hc40433a;
      21277: inst = 32'h8220000;
      21278: inst = 32'h10408000;
      21279: inst = 32'hc40433b;
      21280: inst = 32'h8220000;
      21281: inst = 32'h10408000;
      21282: inst = 32'hc404344;
      21283: inst = 32'h8220000;
      21284: inst = 32'h10408000;
      21285: inst = 32'hc404345;
      21286: inst = 32'h8220000;
      21287: inst = 32'h10408000;
      21288: inst = 32'hc40439a;
      21289: inst = 32'h8220000;
      21290: inst = 32'h10408000;
      21291: inst = 32'hc40439b;
      21292: inst = 32'h8220000;
      21293: inst = 32'h10408000;
      21294: inst = 32'hc4043a4;
      21295: inst = 32'h8220000;
      21296: inst = 32'h10408000;
      21297: inst = 32'hc4043a5;
      21298: inst = 32'h8220000;
      21299: inst = 32'h10408000;
      21300: inst = 32'hc4043fa;
      21301: inst = 32'h8220000;
      21302: inst = 32'h10408000;
      21303: inst = 32'hc4043fb;
      21304: inst = 32'h8220000;
      21305: inst = 32'h10408000;
      21306: inst = 32'hc404404;
      21307: inst = 32'h8220000;
      21308: inst = 32'h10408000;
      21309: inst = 32'hc404405;
      21310: inst = 32'h8220000;
      21311: inst = 32'h10408000;
      21312: inst = 32'hc40445a;
      21313: inst = 32'h8220000;
      21314: inst = 32'h10408000;
      21315: inst = 32'hc40445b;
      21316: inst = 32'h8220000;
      21317: inst = 32'h10408000;
      21318: inst = 32'hc404464;
      21319: inst = 32'h8220000;
      21320: inst = 32'h10408000;
      21321: inst = 32'hc404465;
      21322: inst = 32'h8220000;
      21323: inst = 32'h10408000;
      21324: inst = 32'hc4044ba;
      21325: inst = 32'h8220000;
      21326: inst = 32'h10408000;
      21327: inst = 32'hc4044bb;
      21328: inst = 32'h8220000;
      21329: inst = 32'h10408000;
      21330: inst = 32'hc4044c4;
      21331: inst = 32'h8220000;
      21332: inst = 32'h10408000;
      21333: inst = 32'hc4044c5;
      21334: inst = 32'h8220000;
      21335: inst = 32'h10408000;
      21336: inst = 32'hc40451a;
      21337: inst = 32'h8220000;
      21338: inst = 32'h10408000;
      21339: inst = 32'hc40451b;
      21340: inst = 32'h8220000;
      21341: inst = 32'h10408000;
      21342: inst = 32'hc404524;
      21343: inst = 32'h8220000;
      21344: inst = 32'h10408000;
      21345: inst = 32'hc404525;
      21346: inst = 32'h8220000;
      21347: inst = 32'h10408000;
      21348: inst = 32'hc40457a;
      21349: inst = 32'h8220000;
      21350: inst = 32'h10408000;
      21351: inst = 32'hc40457b;
      21352: inst = 32'h8220000;
      21353: inst = 32'h10408000;
      21354: inst = 32'hc404584;
      21355: inst = 32'h8220000;
      21356: inst = 32'h10408000;
      21357: inst = 32'hc404585;
      21358: inst = 32'h8220000;
      21359: inst = 32'h10408000;
      21360: inst = 32'hc4045da;
      21361: inst = 32'h8220000;
      21362: inst = 32'h10408000;
      21363: inst = 32'hc4045db;
      21364: inst = 32'h8220000;
      21365: inst = 32'h10408000;
      21366: inst = 32'hc4045e4;
      21367: inst = 32'h8220000;
      21368: inst = 32'h10408000;
      21369: inst = 32'hc4045e5;
      21370: inst = 32'h8220000;
      21371: inst = 32'h10408000;
      21372: inst = 32'hc40463a;
      21373: inst = 32'h8220000;
      21374: inst = 32'h10408000;
      21375: inst = 32'hc40463b;
      21376: inst = 32'h8220000;
      21377: inst = 32'h10408000;
      21378: inst = 32'hc404644;
      21379: inst = 32'h8220000;
      21380: inst = 32'h10408000;
      21381: inst = 32'hc404645;
      21382: inst = 32'h8220000;
      21383: inst = 32'h10408000;
      21384: inst = 32'hc40469a;
      21385: inst = 32'h8220000;
      21386: inst = 32'h10408000;
      21387: inst = 32'hc40469b;
      21388: inst = 32'h8220000;
      21389: inst = 32'h10408000;
      21390: inst = 32'hc4046a4;
      21391: inst = 32'h8220000;
      21392: inst = 32'h10408000;
      21393: inst = 32'hc4046a5;
      21394: inst = 32'h8220000;
      21395: inst = 32'h10408000;
      21396: inst = 32'hc4046fa;
      21397: inst = 32'h8220000;
      21398: inst = 32'h10408000;
      21399: inst = 32'hc4046fb;
      21400: inst = 32'h8220000;
      21401: inst = 32'h10408000;
      21402: inst = 32'hc404704;
      21403: inst = 32'h8220000;
      21404: inst = 32'h10408000;
      21405: inst = 32'hc404705;
      21406: inst = 32'h8220000;
      21407: inst = 32'h10408000;
      21408: inst = 32'hc40475a;
      21409: inst = 32'h8220000;
      21410: inst = 32'h10408000;
      21411: inst = 32'hc40475b;
      21412: inst = 32'h8220000;
      21413: inst = 32'h10408000;
      21414: inst = 32'hc404764;
      21415: inst = 32'h8220000;
      21416: inst = 32'h10408000;
      21417: inst = 32'hc404765;
      21418: inst = 32'h8220000;
      21419: inst = 32'h10408000;
      21420: inst = 32'hc4047ba;
      21421: inst = 32'h8220000;
      21422: inst = 32'h10408000;
      21423: inst = 32'hc4047bb;
      21424: inst = 32'h8220000;
      21425: inst = 32'h10408000;
      21426: inst = 32'hc4047c4;
      21427: inst = 32'h8220000;
      21428: inst = 32'h10408000;
      21429: inst = 32'hc4047c5;
      21430: inst = 32'h8220000;
      21431: inst = 32'h10408000;
      21432: inst = 32'hc40481a;
      21433: inst = 32'h8220000;
      21434: inst = 32'h10408000;
      21435: inst = 32'hc40481b;
      21436: inst = 32'h8220000;
      21437: inst = 32'h10408000;
      21438: inst = 32'hc404824;
      21439: inst = 32'h8220000;
      21440: inst = 32'h10408000;
      21441: inst = 32'hc404825;
      21442: inst = 32'h8220000;
      21443: inst = 32'h10408000;
      21444: inst = 32'hc40487a;
      21445: inst = 32'h8220000;
      21446: inst = 32'h10408000;
      21447: inst = 32'hc40487b;
      21448: inst = 32'h8220000;
      21449: inst = 32'h10408000;
      21450: inst = 32'hc404884;
      21451: inst = 32'h8220000;
      21452: inst = 32'h10408000;
      21453: inst = 32'hc404885;
      21454: inst = 32'h8220000;
      21455: inst = 32'h10408000;
      21456: inst = 32'hc4048da;
      21457: inst = 32'h8220000;
      21458: inst = 32'h10408000;
      21459: inst = 32'hc4048db;
      21460: inst = 32'h8220000;
      21461: inst = 32'h10408000;
      21462: inst = 32'hc4048e4;
      21463: inst = 32'h8220000;
      21464: inst = 32'h10408000;
      21465: inst = 32'hc4048e5;
      21466: inst = 32'h8220000;
      21467: inst = 32'h10408000;
      21468: inst = 32'hc40493a;
      21469: inst = 32'h8220000;
      21470: inst = 32'h10408000;
      21471: inst = 32'hc40493b;
      21472: inst = 32'h8220000;
      21473: inst = 32'h10408000;
      21474: inst = 32'hc404944;
      21475: inst = 32'h8220000;
      21476: inst = 32'h10408000;
      21477: inst = 32'hc404945;
      21478: inst = 32'h8220000;
      21479: inst = 32'h10408000;
      21480: inst = 32'hc40499a;
      21481: inst = 32'h8220000;
      21482: inst = 32'h10408000;
      21483: inst = 32'hc40499b;
      21484: inst = 32'h8220000;
      21485: inst = 32'h10408000;
      21486: inst = 32'hc4049a4;
      21487: inst = 32'h8220000;
      21488: inst = 32'h10408000;
      21489: inst = 32'hc4049a5;
      21490: inst = 32'h8220000;
      21491: inst = 32'h10408000;
      21492: inst = 32'hc4049fa;
      21493: inst = 32'h8220000;
      21494: inst = 32'h10408000;
      21495: inst = 32'hc4049fb;
      21496: inst = 32'h8220000;
      21497: inst = 32'h10408000;
      21498: inst = 32'hc404a04;
      21499: inst = 32'h8220000;
      21500: inst = 32'h10408000;
      21501: inst = 32'hc404a05;
      21502: inst = 32'h8220000;
      21503: inst = 32'h10408000;
      21504: inst = 32'hc404a5a;
      21505: inst = 32'h8220000;
      21506: inst = 32'h10408000;
      21507: inst = 32'hc404a5b;
      21508: inst = 32'h8220000;
      21509: inst = 32'h10408000;
      21510: inst = 32'hc404a64;
      21511: inst = 32'h8220000;
      21512: inst = 32'h10408000;
      21513: inst = 32'hc404a65;
      21514: inst = 32'h8220000;
      21515: inst = 32'h10408000;
      21516: inst = 32'hc404aba;
      21517: inst = 32'h8220000;
      21518: inst = 32'h10408000;
      21519: inst = 32'hc404abb;
      21520: inst = 32'h8220000;
      21521: inst = 32'h10408000;
      21522: inst = 32'hc404ac4;
      21523: inst = 32'h8220000;
      21524: inst = 32'h10408000;
      21525: inst = 32'hc404ac5;
      21526: inst = 32'h8220000;
      21527: inst = 32'h10408000;
      21528: inst = 32'hc404b1a;
      21529: inst = 32'h8220000;
      21530: inst = 32'h10408000;
      21531: inst = 32'hc404b1b;
      21532: inst = 32'h8220000;
      21533: inst = 32'h10408000;
      21534: inst = 32'hc404b24;
      21535: inst = 32'h8220000;
      21536: inst = 32'h10408000;
      21537: inst = 32'hc404b25;
      21538: inst = 32'h8220000;
      21539: inst = 32'h10408000;
      21540: inst = 32'hc404b7a;
      21541: inst = 32'h8220000;
      21542: inst = 32'h10408000;
      21543: inst = 32'hc404b7b;
      21544: inst = 32'h8220000;
      21545: inst = 32'h10408000;
      21546: inst = 32'hc404b84;
      21547: inst = 32'h8220000;
      21548: inst = 32'h10408000;
      21549: inst = 32'hc404b85;
      21550: inst = 32'h8220000;
      21551: inst = 32'h10408000;
      21552: inst = 32'hc404bda;
      21553: inst = 32'h8220000;
      21554: inst = 32'h10408000;
      21555: inst = 32'hc404bdb;
      21556: inst = 32'h8220000;
      21557: inst = 32'h10408000;
      21558: inst = 32'hc404be4;
      21559: inst = 32'h8220000;
      21560: inst = 32'h10408000;
      21561: inst = 32'hc404be5;
      21562: inst = 32'h8220000;
      21563: inst = 32'h10408000;
      21564: inst = 32'hc404c3a;
      21565: inst = 32'h8220000;
      21566: inst = 32'h10408000;
      21567: inst = 32'hc404c3b;
      21568: inst = 32'h8220000;
      21569: inst = 32'h10408000;
      21570: inst = 32'hc404c44;
      21571: inst = 32'h8220000;
      21572: inst = 32'h10408000;
      21573: inst = 32'hc404c45;
      21574: inst = 32'h8220000;
      21575: inst = 32'h10408000;
      21576: inst = 32'hc404c9a;
      21577: inst = 32'h8220000;
      21578: inst = 32'h10408000;
      21579: inst = 32'hc404c9b;
      21580: inst = 32'h8220000;
      21581: inst = 32'h10408000;
      21582: inst = 32'hc404ca4;
      21583: inst = 32'h8220000;
      21584: inst = 32'h10408000;
      21585: inst = 32'hc404ca5;
      21586: inst = 32'h8220000;
      21587: inst = 32'h10408000;
      21588: inst = 32'hc404cfa;
      21589: inst = 32'h8220000;
      21590: inst = 32'h10408000;
      21591: inst = 32'hc404cfb;
      21592: inst = 32'h8220000;
      21593: inst = 32'h10408000;
      21594: inst = 32'hc404d04;
      21595: inst = 32'h8220000;
      21596: inst = 32'h10408000;
      21597: inst = 32'hc404d05;
      21598: inst = 32'h8220000;
      21599: inst = 32'h10408000;
      21600: inst = 32'hc404d5a;
      21601: inst = 32'h8220000;
      21602: inst = 32'h10408000;
      21603: inst = 32'hc404d5b;
      21604: inst = 32'h8220000;
      21605: inst = 32'h10408000;
      21606: inst = 32'hc404d64;
      21607: inst = 32'h8220000;
      21608: inst = 32'h10408000;
      21609: inst = 32'hc404d65;
      21610: inst = 32'h8220000;
      21611: inst = 32'h10408000;
      21612: inst = 32'hc404dba;
      21613: inst = 32'h8220000;
      21614: inst = 32'h10408000;
      21615: inst = 32'hc404dbb;
      21616: inst = 32'h8220000;
      21617: inst = 32'h10408000;
      21618: inst = 32'hc404dc4;
      21619: inst = 32'h8220000;
      21620: inst = 32'h10408000;
      21621: inst = 32'hc404dc5;
      21622: inst = 32'h8220000;
      21623: inst = 32'h10408000;
      21624: inst = 32'hc404e1a;
      21625: inst = 32'h8220000;
      21626: inst = 32'h10408000;
      21627: inst = 32'hc404e1b;
      21628: inst = 32'h8220000;
      21629: inst = 32'h10408000;
      21630: inst = 32'hc404e24;
      21631: inst = 32'h8220000;
      21632: inst = 32'h10408000;
      21633: inst = 32'hc404e25;
      21634: inst = 32'h8220000;
      21635: inst = 32'h10408000;
      21636: inst = 32'hc404e7a;
      21637: inst = 32'h8220000;
      21638: inst = 32'h10408000;
      21639: inst = 32'hc404e7b;
      21640: inst = 32'h8220000;
      21641: inst = 32'h10408000;
      21642: inst = 32'hc404e84;
      21643: inst = 32'h8220000;
      21644: inst = 32'h10408000;
      21645: inst = 32'hc404e85;
      21646: inst = 32'h8220000;
      21647: inst = 32'h10408000;
      21648: inst = 32'hc404eda;
      21649: inst = 32'h8220000;
      21650: inst = 32'h10408000;
      21651: inst = 32'hc404edb;
      21652: inst = 32'h8220000;
      21653: inst = 32'h10408000;
      21654: inst = 32'hc404ee4;
      21655: inst = 32'h8220000;
      21656: inst = 32'h10408000;
      21657: inst = 32'hc404ee5;
      21658: inst = 32'h8220000;
      21659: inst = 32'h10408000;
      21660: inst = 32'hc404f3a;
      21661: inst = 32'h8220000;
      21662: inst = 32'h10408000;
      21663: inst = 32'hc404f3b;
      21664: inst = 32'h8220000;
      21665: inst = 32'h10408000;
      21666: inst = 32'hc404f44;
      21667: inst = 32'h8220000;
      21668: inst = 32'h10408000;
      21669: inst = 32'hc404f45;
      21670: inst = 32'h8220000;
      21671: inst = 32'h10408000;
      21672: inst = 32'hc404f9a;
      21673: inst = 32'h8220000;
      21674: inst = 32'h10408000;
      21675: inst = 32'hc404f9b;
      21676: inst = 32'h8220000;
      21677: inst = 32'h10408000;
      21678: inst = 32'hc404fa4;
      21679: inst = 32'h8220000;
      21680: inst = 32'h10408000;
      21681: inst = 32'hc404fa5;
      21682: inst = 32'h8220000;
      21683: inst = 32'h10408000;
      21684: inst = 32'hc404ffa;
      21685: inst = 32'h8220000;
      21686: inst = 32'h10408000;
      21687: inst = 32'hc404ffb;
      21688: inst = 32'h8220000;
      21689: inst = 32'h10408000;
      21690: inst = 32'hc405004;
      21691: inst = 32'h8220000;
      21692: inst = 32'h10408000;
      21693: inst = 32'hc405005;
      21694: inst = 32'h8220000;
      21695: inst = 32'h10408000;
      21696: inst = 32'hc40505a;
      21697: inst = 32'h8220000;
      21698: inst = 32'h10408000;
      21699: inst = 32'hc40505b;
      21700: inst = 32'h8220000;
      21701: inst = 32'h10408000;
      21702: inst = 32'hc405064;
      21703: inst = 32'h8220000;
      21704: inst = 32'h10408000;
      21705: inst = 32'hc405065;
      21706: inst = 32'h8220000;
      21707: inst = 32'h10408000;
      21708: inst = 32'hc4050ba;
      21709: inst = 32'h8220000;
      21710: inst = 32'h10408000;
      21711: inst = 32'hc4050bb;
      21712: inst = 32'h8220000;
      21713: inst = 32'h10408000;
      21714: inst = 32'hc4050c4;
      21715: inst = 32'h8220000;
      21716: inst = 32'h10408000;
      21717: inst = 32'hc4050c5;
      21718: inst = 32'h8220000;
      21719: inst = 32'h10408000;
      21720: inst = 32'hc40511a;
      21721: inst = 32'h8220000;
      21722: inst = 32'h10408000;
      21723: inst = 32'hc40511b;
      21724: inst = 32'h8220000;
      21725: inst = 32'h10408000;
      21726: inst = 32'hc405124;
      21727: inst = 32'h8220000;
      21728: inst = 32'h10408000;
      21729: inst = 32'hc405125;
      21730: inst = 32'h8220000;
      21731: inst = 32'h10408000;
      21732: inst = 32'hc40517a;
      21733: inst = 32'h8220000;
      21734: inst = 32'h10408000;
      21735: inst = 32'hc40517b;
      21736: inst = 32'h8220000;
      21737: inst = 32'h10408000;
      21738: inst = 32'hc405184;
      21739: inst = 32'h8220000;
      21740: inst = 32'h10408000;
      21741: inst = 32'hc405185;
      21742: inst = 32'h8220000;
      21743: inst = 32'h10408000;
      21744: inst = 32'hc4051da;
      21745: inst = 32'h8220000;
      21746: inst = 32'h10408000;
      21747: inst = 32'hc4051db;
      21748: inst = 32'h8220000;
      21749: inst = 32'h10408000;
      21750: inst = 32'hc4051e4;
      21751: inst = 32'h8220000;
      21752: inst = 32'h10408000;
      21753: inst = 32'hc4051e5;
      21754: inst = 32'h8220000;
      21755: inst = 32'h10408000;
      21756: inst = 32'hc40523a;
      21757: inst = 32'h8220000;
      21758: inst = 32'h10408000;
      21759: inst = 32'hc40523b;
      21760: inst = 32'h8220000;
      21761: inst = 32'h10408000;
      21762: inst = 32'hc405244;
      21763: inst = 32'h8220000;
      21764: inst = 32'h10408000;
      21765: inst = 32'hc405245;
      21766: inst = 32'h8220000;
      21767: inst = 32'h10408000;
      21768: inst = 32'hc40529a;
      21769: inst = 32'h8220000;
      21770: inst = 32'h10408000;
      21771: inst = 32'hc40529b;
      21772: inst = 32'h8220000;
      21773: inst = 32'h10408000;
      21774: inst = 32'hc4052a4;
      21775: inst = 32'h8220000;
      21776: inst = 32'h10408000;
      21777: inst = 32'hc4052a5;
      21778: inst = 32'h8220000;
      21779: inst = 32'h10408000;
      21780: inst = 32'hc4052fa;
      21781: inst = 32'h8220000;
      21782: inst = 32'h10408000;
      21783: inst = 32'hc4052fb;
      21784: inst = 32'h8220000;
      21785: inst = 32'h10408000;
      21786: inst = 32'hc405304;
      21787: inst = 32'h8220000;
      21788: inst = 32'h10408000;
      21789: inst = 32'hc405305;
      21790: inst = 32'h8220000;
      21791: inst = 32'h10408000;
      21792: inst = 32'hc40535a;
      21793: inst = 32'h8220000;
      21794: inst = 32'h10408000;
      21795: inst = 32'hc40535b;
      21796: inst = 32'h8220000;
      21797: inst = 32'h10408000;
      21798: inst = 32'hc405364;
      21799: inst = 32'h8220000;
      21800: inst = 32'h10408000;
      21801: inst = 32'hc405365;
      21802: inst = 32'h8220000;
      21803: inst = 32'h10408000;
      21804: inst = 32'hc4053ba;
      21805: inst = 32'h8220000;
      21806: inst = 32'h10408000;
      21807: inst = 32'hc4053bb;
      21808: inst = 32'h8220000;
      21809: inst = 32'h10408000;
      21810: inst = 32'hc4053c4;
      21811: inst = 32'h8220000;
      21812: inst = 32'h10408000;
      21813: inst = 32'hc4053c5;
      21814: inst = 32'h8220000;
      21815: inst = 32'h10408000;
      21816: inst = 32'hc40541a;
      21817: inst = 32'h8220000;
      21818: inst = 32'h10408000;
      21819: inst = 32'hc40541b;
      21820: inst = 32'h8220000;
      21821: inst = 32'h10408000;
      21822: inst = 32'hc405424;
      21823: inst = 32'h8220000;
      21824: inst = 32'h10408000;
      21825: inst = 32'hc405425;
      21826: inst = 32'h8220000;
      21827: inst = 32'h10408000;
      21828: inst = 32'hc405426;
      21829: inst = 32'h8220000;
      21830: inst = 32'h10408000;
      21831: inst = 32'hc405479;
      21832: inst = 32'h8220000;
      21833: inst = 32'h10408000;
      21834: inst = 32'hc40547a;
      21835: inst = 32'h8220000;
      21836: inst = 32'h10408000;
      21837: inst = 32'hc40547b;
      21838: inst = 32'h8220000;
      21839: inst = 32'h10408000;
      21840: inst = 32'hc405484;
      21841: inst = 32'h8220000;
      21842: inst = 32'h10408000;
      21843: inst = 32'hc405485;
      21844: inst = 32'h8220000;
      21845: inst = 32'h10408000;
      21846: inst = 32'hc405486;
      21847: inst = 32'h8220000;
      21848: inst = 32'h10408000;
      21849: inst = 32'hc405487;
      21850: inst = 32'h8220000;
      21851: inst = 32'h10408000;
      21852: inst = 32'hc405488;
      21853: inst = 32'h8220000;
      21854: inst = 32'h10408000;
      21855: inst = 32'hc405489;
      21856: inst = 32'h8220000;
      21857: inst = 32'h10408000;
      21858: inst = 32'hc40548a;
      21859: inst = 32'h8220000;
      21860: inst = 32'h10408000;
      21861: inst = 32'hc40548b;
      21862: inst = 32'h8220000;
      21863: inst = 32'h10408000;
      21864: inst = 32'hc40548c;
      21865: inst = 32'h8220000;
      21866: inst = 32'h10408000;
      21867: inst = 32'hc40548d;
      21868: inst = 32'h8220000;
      21869: inst = 32'h10408000;
      21870: inst = 32'hc40548e;
      21871: inst = 32'h8220000;
      21872: inst = 32'h10408000;
      21873: inst = 32'hc40548f;
      21874: inst = 32'h8220000;
      21875: inst = 32'h10408000;
      21876: inst = 32'hc405490;
      21877: inst = 32'h8220000;
      21878: inst = 32'h10408000;
      21879: inst = 32'hc405491;
      21880: inst = 32'h8220000;
      21881: inst = 32'h10408000;
      21882: inst = 32'hc405492;
      21883: inst = 32'h8220000;
      21884: inst = 32'h10408000;
      21885: inst = 32'hc405493;
      21886: inst = 32'h8220000;
      21887: inst = 32'h10408000;
      21888: inst = 32'hc405494;
      21889: inst = 32'h8220000;
      21890: inst = 32'h10408000;
      21891: inst = 32'hc405495;
      21892: inst = 32'h8220000;
      21893: inst = 32'h10408000;
      21894: inst = 32'hc405496;
      21895: inst = 32'h8220000;
      21896: inst = 32'h10408000;
      21897: inst = 32'hc405497;
      21898: inst = 32'h8220000;
      21899: inst = 32'h10408000;
      21900: inst = 32'hc405498;
      21901: inst = 32'h8220000;
      21902: inst = 32'h10408000;
      21903: inst = 32'hc405499;
      21904: inst = 32'h8220000;
      21905: inst = 32'h10408000;
      21906: inst = 32'hc40549a;
      21907: inst = 32'h8220000;
      21908: inst = 32'h10408000;
      21909: inst = 32'hc40549b;
      21910: inst = 32'h8220000;
      21911: inst = 32'h10408000;
      21912: inst = 32'hc40549c;
      21913: inst = 32'h8220000;
      21914: inst = 32'h10408000;
      21915: inst = 32'hc40549d;
      21916: inst = 32'h8220000;
      21917: inst = 32'h10408000;
      21918: inst = 32'hc40549e;
      21919: inst = 32'h8220000;
      21920: inst = 32'h10408000;
      21921: inst = 32'hc40549f;
      21922: inst = 32'h8220000;
      21923: inst = 32'h10408000;
      21924: inst = 32'hc4054a0;
      21925: inst = 32'h8220000;
      21926: inst = 32'h10408000;
      21927: inst = 32'hc4054a1;
      21928: inst = 32'h8220000;
      21929: inst = 32'h10408000;
      21930: inst = 32'hc4054a2;
      21931: inst = 32'h8220000;
      21932: inst = 32'h10408000;
      21933: inst = 32'hc4054a3;
      21934: inst = 32'h8220000;
      21935: inst = 32'h10408000;
      21936: inst = 32'hc4054a4;
      21937: inst = 32'h8220000;
      21938: inst = 32'h10408000;
      21939: inst = 32'hc4054a5;
      21940: inst = 32'h8220000;
      21941: inst = 32'h10408000;
      21942: inst = 32'hc4054a6;
      21943: inst = 32'h8220000;
      21944: inst = 32'h10408000;
      21945: inst = 32'hc4054a7;
      21946: inst = 32'h8220000;
      21947: inst = 32'h10408000;
      21948: inst = 32'hc4054a8;
      21949: inst = 32'h8220000;
      21950: inst = 32'h10408000;
      21951: inst = 32'hc4054a9;
      21952: inst = 32'h8220000;
      21953: inst = 32'h10408000;
      21954: inst = 32'hc4054aa;
      21955: inst = 32'h8220000;
      21956: inst = 32'h10408000;
      21957: inst = 32'hc4054ab;
      21958: inst = 32'h8220000;
      21959: inst = 32'h10408000;
      21960: inst = 32'hc4054ac;
      21961: inst = 32'h8220000;
      21962: inst = 32'h10408000;
      21963: inst = 32'hc4054ad;
      21964: inst = 32'h8220000;
      21965: inst = 32'h10408000;
      21966: inst = 32'hc4054ae;
      21967: inst = 32'h8220000;
      21968: inst = 32'h10408000;
      21969: inst = 32'hc4054af;
      21970: inst = 32'h8220000;
      21971: inst = 32'h10408000;
      21972: inst = 32'hc4054b0;
      21973: inst = 32'h8220000;
      21974: inst = 32'h10408000;
      21975: inst = 32'hc4054b1;
      21976: inst = 32'h8220000;
      21977: inst = 32'h10408000;
      21978: inst = 32'hc4054b2;
      21979: inst = 32'h8220000;
      21980: inst = 32'h10408000;
      21981: inst = 32'hc4054b3;
      21982: inst = 32'h8220000;
      21983: inst = 32'h10408000;
      21984: inst = 32'hc4054b4;
      21985: inst = 32'h8220000;
      21986: inst = 32'h10408000;
      21987: inst = 32'hc4054b5;
      21988: inst = 32'h8220000;
      21989: inst = 32'h10408000;
      21990: inst = 32'hc4054b6;
      21991: inst = 32'h8220000;
      21992: inst = 32'h10408000;
      21993: inst = 32'hc4054b7;
      21994: inst = 32'h8220000;
      21995: inst = 32'h10408000;
      21996: inst = 32'hc4054b8;
      21997: inst = 32'h8220000;
      21998: inst = 32'h10408000;
      21999: inst = 32'hc4054b9;
      22000: inst = 32'h8220000;
      22001: inst = 32'h10408000;
      22002: inst = 32'hc4054ba;
      22003: inst = 32'h8220000;
      22004: inst = 32'h10408000;
      22005: inst = 32'hc4054bb;
      22006: inst = 32'h8220000;
      22007: inst = 32'h10408000;
      22008: inst = 32'hc4054bc;
      22009: inst = 32'h8220000;
      22010: inst = 32'h10408000;
      22011: inst = 32'hc4054bd;
      22012: inst = 32'h8220000;
      22013: inst = 32'h10408000;
      22014: inst = 32'hc4054be;
      22015: inst = 32'h8220000;
      22016: inst = 32'h10408000;
      22017: inst = 32'hc4054bf;
      22018: inst = 32'h8220000;
      22019: inst = 32'h10408000;
      22020: inst = 32'hc4054c0;
      22021: inst = 32'h8220000;
      22022: inst = 32'h10408000;
      22023: inst = 32'hc4054c1;
      22024: inst = 32'h8220000;
      22025: inst = 32'h10408000;
      22026: inst = 32'hc4054c2;
      22027: inst = 32'h8220000;
      22028: inst = 32'h10408000;
      22029: inst = 32'hc4054c3;
      22030: inst = 32'h8220000;
      22031: inst = 32'h10408000;
      22032: inst = 32'hc4054c4;
      22033: inst = 32'h8220000;
      22034: inst = 32'h10408000;
      22035: inst = 32'hc4054c5;
      22036: inst = 32'h8220000;
      22037: inst = 32'h10408000;
      22038: inst = 32'hc4054c6;
      22039: inst = 32'h8220000;
      22040: inst = 32'h10408000;
      22041: inst = 32'hc4054c7;
      22042: inst = 32'h8220000;
      22043: inst = 32'h10408000;
      22044: inst = 32'hc4054c8;
      22045: inst = 32'h8220000;
      22046: inst = 32'h10408000;
      22047: inst = 32'hc4054c9;
      22048: inst = 32'h8220000;
      22049: inst = 32'h10408000;
      22050: inst = 32'hc4054ca;
      22051: inst = 32'h8220000;
      22052: inst = 32'h10408000;
      22053: inst = 32'hc4054cb;
      22054: inst = 32'h8220000;
      22055: inst = 32'h10408000;
      22056: inst = 32'hc4054cc;
      22057: inst = 32'h8220000;
      22058: inst = 32'h10408000;
      22059: inst = 32'hc4054cd;
      22060: inst = 32'h8220000;
      22061: inst = 32'h10408000;
      22062: inst = 32'hc4054ce;
      22063: inst = 32'h8220000;
      22064: inst = 32'h10408000;
      22065: inst = 32'hc4054cf;
      22066: inst = 32'h8220000;
      22067: inst = 32'h10408000;
      22068: inst = 32'hc4054d0;
      22069: inst = 32'h8220000;
      22070: inst = 32'h10408000;
      22071: inst = 32'hc4054d1;
      22072: inst = 32'h8220000;
      22073: inst = 32'h10408000;
      22074: inst = 32'hc4054d2;
      22075: inst = 32'h8220000;
      22076: inst = 32'h10408000;
      22077: inst = 32'hc4054d3;
      22078: inst = 32'h8220000;
      22079: inst = 32'h10408000;
      22080: inst = 32'hc4054d4;
      22081: inst = 32'h8220000;
      22082: inst = 32'h10408000;
      22083: inst = 32'hc4054d5;
      22084: inst = 32'h8220000;
      22085: inst = 32'h10408000;
      22086: inst = 32'hc4054d6;
      22087: inst = 32'h8220000;
      22088: inst = 32'h10408000;
      22089: inst = 32'hc4054d7;
      22090: inst = 32'h8220000;
      22091: inst = 32'h10408000;
      22092: inst = 32'hc4054d8;
      22093: inst = 32'h8220000;
      22094: inst = 32'h10408000;
      22095: inst = 32'hc4054d9;
      22096: inst = 32'h8220000;
      22097: inst = 32'h10408000;
      22098: inst = 32'hc4054da;
      22099: inst = 32'h8220000;
      22100: inst = 32'h10408000;
      22101: inst = 32'hc4054db;
      22102: inst = 32'h8220000;
      22103: inst = 32'h10408000;
      22104: inst = 32'hc4054e4;
      22105: inst = 32'h8220000;
      22106: inst = 32'h10408000;
      22107: inst = 32'hc4054e5;
      22108: inst = 32'h8220000;
      22109: inst = 32'h10408000;
      22110: inst = 32'hc4054e6;
      22111: inst = 32'h8220000;
      22112: inst = 32'h10408000;
      22113: inst = 32'hc4054e7;
      22114: inst = 32'h8220000;
      22115: inst = 32'h10408000;
      22116: inst = 32'hc4054e8;
      22117: inst = 32'h8220000;
      22118: inst = 32'h10408000;
      22119: inst = 32'hc4054e9;
      22120: inst = 32'h8220000;
      22121: inst = 32'h10408000;
      22122: inst = 32'hc4054ea;
      22123: inst = 32'h8220000;
      22124: inst = 32'h10408000;
      22125: inst = 32'hc4054eb;
      22126: inst = 32'h8220000;
      22127: inst = 32'h10408000;
      22128: inst = 32'hc4054ec;
      22129: inst = 32'h8220000;
      22130: inst = 32'h10408000;
      22131: inst = 32'hc4054ed;
      22132: inst = 32'h8220000;
      22133: inst = 32'h10408000;
      22134: inst = 32'hc4054ee;
      22135: inst = 32'h8220000;
      22136: inst = 32'h10408000;
      22137: inst = 32'hc4054ef;
      22138: inst = 32'h8220000;
      22139: inst = 32'h10408000;
      22140: inst = 32'hc4054f0;
      22141: inst = 32'h8220000;
      22142: inst = 32'h10408000;
      22143: inst = 32'hc4054f1;
      22144: inst = 32'h8220000;
      22145: inst = 32'h10408000;
      22146: inst = 32'hc4054f2;
      22147: inst = 32'h8220000;
      22148: inst = 32'h10408000;
      22149: inst = 32'hc4054f3;
      22150: inst = 32'h8220000;
      22151: inst = 32'h10408000;
      22152: inst = 32'hc4054f4;
      22153: inst = 32'h8220000;
      22154: inst = 32'h10408000;
      22155: inst = 32'hc4054f5;
      22156: inst = 32'h8220000;
      22157: inst = 32'h10408000;
      22158: inst = 32'hc4054f6;
      22159: inst = 32'h8220000;
      22160: inst = 32'h10408000;
      22161: inst = 32'hc4054f7;
      22162: inst = 32'h8220000;
      22163: inst = 32'h10408000;
      22164: inst = 32'hc4054f8;
      22165: inst = 32'h8220000;
      22166: inst = 32'h10408000;
      22167: inst = 32'hc4054f9;
      22168: inst = 32'h8220000;
      22169: inst = 32'h10408000;
      22170: inst = 32'hc4054fa;
      22171: inst = 32'h8220000;
      22172: inst = 32'h10408000;
      22173: inst = 32'hc4054fb;
      22174: inst = 32'h8220000;
      22175: inst = 32'h10408000;
      22176: inst = 32'hc4054fc;
      22177: inst = 32'h8220000;
      22178: inst = 32'h10408000;
      22179: inst = 32'hc4054fd;
      22180: inst = 32'h8220000;
      22181: inst = 32'h10408000;
      22182: inst = 32'hc4054fe;
      22183: inst = 32'h8220000;
      22184: inst = 32'h10408000;
      22185: inst = 32'hc4054ff;
      22186: inst = 32'h8220000;
      22187: inst = 32'h10408000;
      22188: inst = 32'hc405500;
      22189: inst = 32'h8220000;
      22190: inst = 32'h10408000;
      22191: inst = 32'hc405501;
      22192: inst = 32'h8220000;
      22193: inst = 32'h10408000;
      22194: inst = 32'hc405502;
      22195: inst = 32'h8220000;
      22196: inst = 32'h10408000;
      22197: inst = 32'hc405503;
      22198: inst = 32'h8220000;
      22199: inst = 32'h10408000;
      22200: inst = 32'hc405504;
      22201: inst = 32'h8220000;
      22202: inst = 32'h10408000;
      22203: inst = 32'hc405505;
      22204: inst = 32'h8220000;
      22205: inst = 32'h10408000;
      22206: inst = 32'hc405506;
      22207: inst = 32'h8220000;
      22208: inst = 32'h10408000;
      22209: inst = 32'hc405507;
      22210: inst = 32'h8220000;
      22211: inst = 32'h10408000;
      22212: inst = 32'hc405508;
      22213: inst = 32'h8220000;
      22214: inst = 32'h10408000;
      22215: inst = 32'hc405509;
      22216: inst = 32'h8220000;
      22217: inst = 32'h10408000;
      22218: inst = 32'hc40550a;
      22219: inst = 32'h8220000;
      22220: inst = 32'h10408000;
      22221: inst = 32'hc40550b;
      22222: inst = 32'h8220000;
      22223: inst = 32'h10408000;
      22224: inst = 32'hc40550c;
      22225: inst = 32'h8220000;
      22226: inst = 32'h10408000;
      22227: inst = 32'hc40550d;
      22228: inst = 32'h8220000;
      22229: inst = 32'h10408000;
      22230: inst = 32'hc40550e;
      22231: inst = 32'h8220000;
      22232: inst = 32'h10408000;
      22233: inst = 32'hc40550f;
      22234: inst = 32'h8220000;
      22235: inst = 32'h10408000;
      22236: inst = 32'hc405510;
      22237: inst = 32'h8220000;
      22238: inst = 32'h10408000;
      22239: inst = 32'hc405511;
      22240: inst = 32'h8220000;
      22241: inst = 32'h10408000;
      22242: inst = 32'hc405512;
      22243: inst = 32'h8220000;
      22244: inst = 32'h10408000;
      22245: inst = 32'hc405513;
      22246: inst = 32'h8220000;
      22247: inst = 32'h10408000;
      22248: inst = 32'hc405514;
      22249: inst = 32'h8220000;
      22250: inst = 32'h10408000;
      22251: inst = 32'hc405515;
      22252: inst = 32'h8220000;
      22253: inst = 32'h10408000;
      22254: inst = 32'hc405516;
      22255: inst = 32'h8220000;
      22256: inst = 32'h10408000;
      22257: inst = 32'hc405517;
      22258: inst = 32'h8220000;
      22259: inst = 32'h10408000;
      22260: inst = 32'hc405518;
      22261: inst = 32'h8220000;
      22262: inst = 32'h10408000;
      22263: inst = 32'hc405519;
      22264: inst = 32'h8220000;
      22265: inst = 32'h10408000;
      22266: inst = 32'hc40551a;
      22267: inst = 32'h8220000;
      22268: inst = 32'h10408000;
      22269: inst = 32'hc40551b;
      22270: inst = 32'h8220000;
      22271: inst = 32'h10408000;
      22272: inst = 32'hc40551c;
      22273: inst = 32'h8220000;
      22274: inst = 32'h10408000;
      22275: inst = 32'hc40551d;
      22276: inst = 32'h8220000;
      22277: inst = 32'h10408000;
      22278: inst = 32'hc40551e;
      22279: inst = 32'h8220000;
      22280: inst = 32'h10408000;
      22281: inst = 32'hc40551f;
      22282: inst = 32'h8220000;
      22283: inst = 32'h10408000;
      22284: inst = 32'hc405520;
      22285: inst = 32'h8220000;
      22286: inst = 32'h10408000;
      22287: inst = 32'hc405521;
      22288: inst = 32'h8220000;
      22289: inst = 32'h10408000;
      22290: inst = 32'hc405522;
      22291: inst = 32'h8220000;
      22292: inst = 32'h10408000;
      22293: inst = 32'hc405523;
      22294: inst = 32'h8220000;
      22295: inst = 32'h10408000;
      22296: inst = 32'hc405524;
      22297: inst = 32'h8220000;
      22298: inst = 32'h10408000;
      22299: inst = 32'hc405525;
      22300: inst = 32'h8220000;
      22301: inst = 32'h10408000;
      22302: inst = 32'hc405526;
      22303: inst = 32'h8220000;
      22304: inst = 32'h10408000;
      22305: inst = 32'hc405527;
      22306: inst = 32'h8220000;
      22307: inst = 32'h10408000;
      22308: inst = 32'hc405528;
      22309: inst = 32'h8220000;
      22310: inst = 32'h10408000;
      22311: inst = 32'hc405529;
      22312: inst = 32'h8220000;
      22313: inst = 32'h10408000;
      22314: inst = 32'hc40552a;
      22315: inst = 32'h8220000;
      22316: inst = 32'h10408000;
      22317: inst = 32'hc40552b;
      22318: inst = 32'h8220000;
      22319: inst = 32'h10408000;
      22320: inst = 32'hc40552c;
      22321: inst = 32'h8220000;
      22322: inst = 32'h10408000;
      22323: inst = 32'hc40552d;
      22324: inst = 32'h8220000;
      22325: inst = 32'h10408000;
      22326: inst = 32'hc40552e;
      22327: inst = 32'h8220000;
      22328: inst = 32'h10408000;
      22329: inst = 32'hc40552f;
      22330: inst = 32'h8220000;
      22331: inst = 32'h10408000;
      22332: inst = 32'hc405530;
      22333: inst = 32'h8220000;
      22334: inst = 32'h10408000;
      22335: inst = 32'hc405531;
      22336: inst = 32'h8220000;
      22337: inst = 32'h10408000;
      22338: inst = 32'hc405532;
      22339: inst = 32'h8220000;
      22340: inst = 32'h10408000;
      22341: inst = 32'hc405533;
      22342: inst = 32'h8220000;
      22343: inst = 32'h10408000;
      22344: inst = 32'hc405534;
      22345: inst = 32'h8220000;
      22346: inst = 32'h10408000;
      22347: inst = 32'hc405535;
      22348: inst = 32'h8220000;
      22349: inst = 32'h10408000;
      22350: inst = 32'hc405536;
      22351: inst = 32'h8220000;
      22352: inst = 32'h10408000;
      22353: inst = 32'hc405537;
      22354: inst = 32'h8220000;
      22355: inst = 32'h10408000;
      22356: inst = 32'hc405538;
      22357: inst = 32'h8220000;
      22358: inst = 32'h10408000;
      22359: inst = 32'hc405539;
      22360: inst = 32'h8220000;
      22361: inst = 32'h10408000;
      22362: inst = 32'hc40553a;
      22363: inst = 32'h8220000;
      22364: inst = 32'h10408000;
      22365: inst = 32'hc40553b;
      22366: inst = 32'h8220000;
      22367: inst = 32'hc204a7a;
      22368: inst = 32'h10408000;
      22369: inst = 32'hc4042e7;
      22370: inst = 32'h8220000;
      22371: inst = 32'h10408000;
      22372: inst = 32'hc404338;
      22373: inst = 32'h8220000;
      22374: inst = 32'h10408000;
      22375: inst = 32'hc404346;
      22376: inst = 32'h8220000;
      22377: inst = 32'h10408000;
      22378: inst = 32'hc404399;
      22379: inst = 32'h8220000;
      22380: inst = 32'h10408000;
      22381: inst = 32'hc4053c6;
      22382: inst = 32'h8220000;
      22383: inst = 32'h10408000;
      22384: inst = 32'hc405419;
      22385: inst = 32'h8220000;
      22386: inst = 32'h10408000;
      22387: inst = 32'hc405427;
      22388: inst = 32'h8220000;
      22389: inst = 32'h10408000;
      22390: inst = 32'hc405478;
      22391: inst = 32'h8220000;
      22392: inst = 32'hc2031b0;
      22393: inst = 32'h10408000;
      22394: inst = 32'hc4042e8;
      22395: inst = 32'h8220000;
      22396: inst = 32'h10408000;
      22397: inst = 32'hc404337;
      22398: inst = 32'h8220000;
      22399: inst = 32'h10408000;
      22400: inst = 32'hc4043a6;
      22401: inst = 32'h8220000;
      22402: inst = 32'h10408000;
      22403: inst = 32'hc4043f9;
      22404: inst = 32'h8220000;
      22405: inst = 32'h10408000;
      22406: inst = 32'hc405366;
      22407: inst = 32'h8220000;
      22408: inst = 32'h10408000;
      22409: inst = 32'hc4053b9;
      22410: inst = 32'h8220000;
      22411: inst = 32'h10408000;
      22412: inst = 32'hc405428;
      22413: inst = 32'h8220000;
      22414: inst = 32'h10408000;
      22415: inst = 32'hc405477;
      22416: inst = 32'h8220000;
      22417: inst = 32'hc20296d;
      22418: inst = 32'h10408000;
      22419: inst = 32'hc4042e9;
      22420: inst = 32'h8220000;
      22421: inst = 32'h10408000;
      22422: inst = 32'hc4042ea;
      22423: inst = 32'h8220000;
      22424: inst = 32'h10408000;
      22425: inst = 32'hc4042eb;
      22426: inst = 32'h8220000;
      22427: inst = 32'h10408000;
      22428: inst = 32'hc4042ec;
      22429: inst = 32'h8220000;
      22430: inst = 32'h10408000;
      22431: inst = 32'hc4042ed;
      22432: inst = 32'h8220000;
      22433: inst = 32'h10408000;
      22434: inst = 32'hc4042ee;
      22435: inst = 32'h8220000;
      22436: inst = 32'h10408000;
      22437: inst = 32'hc4042ef;
      22438: inst = 32'h8220000;
      22439: inst = 32'h10408000;
      22440: inst = 32'hc4042f0;
      22441: inst = 32'h8220000;
      22442: inst = 32'h10408000;
      22443: inst = 32'hc4042f1;
      22444: inst = 32'h8220000;
      22445: inst = 32'h10408000;
      22446: inst = 32'hc4042f2;
      22447: inst = 32'h8220000;
      22448: inst = 32'h10408000;
      22449: inst = 32'hc4042f3;
      22450: inst = 32'h8220000;
      22451: inst = 32'h10408000;
      22452: inst = 32'hc4042f4;
      22453: inst = 32'h8220000;
      22454: inst = 32'h10408000;
      22455: inst = 32'hc4042f5;
      22456: inst = 32'h8220000;
      22457: inst = 32'h10408000;
      22458: inst = 32'hc4042f6;
      22459: inst = 32'h8220000;
      22460: inst = 32'h10408000;
      22461: inst = 32'hc4042f7;
      22462: inst = 32'h8220000;
      22463: inst = 32'h10408000;
      22464: inst = 32'hc4042f8;
      22465: inst = 32'h8220000;
      22466: inst = 32'h10408000;
      22467: inst = 32'hc4042f9;
      22468: inst = 32'h8220000;
      22469: inst = 32'h10408000;
      22470: inst = 32'hc4042fa;
      22471: inst = 32'h8220000;
      22472: inst = 32'h10408000;
      22473: inst = 32'hc4042fb;
      22474: inst = 32'h8220000;
      22475: inst = 32'h10408000;
      22476: inst = 32'hc4042fc;
      22477: inst = 32'h8220000;
      22478: inst = 32'h10408000;
      22479: inst = 32'hc4042fd;
      22480: inst = 32'h8220000;
      22481: inst = 32'h10408000;
      22482: inst = 32'hc4042fe;
      22483: inst = 32'h8220000;
      22484: inst = 32'h10408000;
      22485: inst = 32'hc4042ff;
      22486: inst = 32'h8220000;
      22487: inst = 32'h10408000;
      22488: inst = 32'hc404300;
      22489: inst = 32'h8220000;
      22490: inst = 32'h10408000;
      22491: inst = 32'hc404301;
      22492: inst = 32'h8220000;
      22493: inst = 32'h10408000;
      22494: inst = 32'hc404302;
      22495: inst = 32'h8220000;
      22496: inst = 32'h10408000;
      22497: inst = 32'hc404303;
      22498: inst = 32'h8220000;
      22499: inst = 32'h10408000;
      22500: inst = 32'hc404304;
      22501: inst = 32'h8220000;
      22502: inst = 32'h10408000;
      22503: inst = 32'hc404305;
      22504: inst = 32'h8220000;
      22505: inst = 32'h10408000;
      22506: inst = 32'hc404306;
      22507: inst = 32'h8220000;
      22508: inst = 32'h10408000;
      22509: inst = 32'hc404307;
      22510: inst = 32'h8220000;
      22511: inst = 32'h10408000;
      22512: inst = 32'hc404308;
      22513: inst = 32'h8220000;
      22514: inst = 32'h10408000;
      22515: inst = 32'hc404309;
      22516: inst = 32'h8220000;
      22517: inst = 32'h10408000;
      22518: inst = 32'hc40430a;
      22519: inst = 32'h8220000;
      22520: inst = 32'h10408000;
      22521: inst = 32'hc40430b;
      22522: inst = 32'h8220000;
      22523: inst = 32'h10408000;
      22524: inst = 32'hc40430c;
      22525: inst = 32'h8220000;
      22526: inst = 32'h10408000;
      22527: inst = 32'hc40430d;
      22528: inst = 32'h8220000;
      22529: inst = 32'h10408000;
      22530: inst = 32'hc40430e;
      22531: inst = 32'h8220000;
      22532: inst = 32'h10408000;
      22533: inst = 32'hc40430f;
      22534: inst = 32'h8220000;
      22535: inst = 32'h10408000;
      22536: inst = 32'hc404310;
      22537: inst = 32'h8220000;
      22538: inst = 32'h10408000;
      22539: inst = 32'hc404311;
      22540: inst = 32'h8220000;
      22541: inst = 32'h10408000;
      22542: inst = 32'hc404312;
      22543: inst = 32'h8220000;
      22544: inst = 32'h10408000;
      22545: inst = 32'hc404313;
      22546: inst = 32'h8220000;
      22547: inst = 32'h10408000;
      22548: inst = 32'hc404314;
      22549: inst = 32'h8220000;
      22550: inst = 32'h10408000;
      22551: inst = 32'hc404315;
      22552: inst = 32'h8220000;
      22553: inst = 32'h10408000;
      22554: inst = 32'hc404316;
      22555: inst = 32'h8220000;
      22556: inst = 32'h10408000;
      22557: inst = 32'hc404317;
      22558: inst = 32'h8220000;
      22559: inst = 32'h10408000;
      22560: inst = 32'hc404318;
      22561: inst = 32'h8220000;
      22562: inst = 32'h10408000;
      22563: inst = 32'hc404319;
      22564: inst = 32'h8220000;
      22565: inst = 32'h10408000;
      22566: inst = 32'hc40431a;
      22567: inst = 32'h8220000;
      22568: inst = 32'h10408000;
      22569: inst = 32'hc40431b;
      22570: inst = 32'h8220000;
      22571: inst = 32'h10408000;
      22572: inst = 32'hc40431c;
      22573: inst = 32'h8220000;
      22574: inst = 32'h10408000;
      22575: inst = 32'hc40431d;
      22576: inst = 32'h8220000;
      22577: inst = 32'h10408000;
      22578: inst = 32'hc40431e;
      22579: inst = 32'h8220000;
      22580: inst = 32'h10408000;
      22581: inst = 32'hc40431f;
      22582: inst = 32'h8220000;
      22583: inst = 32'h10408000;
      22584: inst = 32'hc404320;
      22585: inst = 32'h8220000;
      22586: inst = 32'h10408000;
      22587: inst = 32'hc404321;
      22588: inst = 32'h8220000;
      22589: inst = 32'h10408000;
      22590: inst = 32'hc404322;
      22591: inst = 32'h8220000;
      22592: inst = 32'h10408000;
      22593: inst = 32'hc404323;
      22594: inst = 32'h8220000;
      22595: inst = 32'h10408000;
      22596: inst = 32'hc404324;
      22597: inst = 32'h8220000;
      22598: inst = 32'h10408000;
      22599: inst = 32'hc404325;
      22600: inst = 32'h8220000;
      22601: inst = 32'h10408000;
      22602: inst = 32'hc404326;
      22603: inst = 32'h8220000;
      22604: inst = 32'h10408000;
      22605: inst = 32'hc404327;
      22606: inst = 32'h8220000;
      22607: inst = 32'h10408000;
      22608: inst = 32'hc404328;
      22609: inst = 32'h8220000;
      22610: inst = 32'h10408000;
      22611: inst = 32'hc404329;
      22612: inst = 32'h8220000;
      22613: inst = 32'h10408000;
      22614: inst = 32'hc40432a;
      22615: inst = 32'h8220000;
      22616: inst = 32'h10408000;
      22617: inst = 32'hc40432b;
      22618: inst = 32'h8220000;
      22619: inst = 32'h10408000;
      22620: inst = 32'hc40432c;
      22621: inst = 32'h8220000;
      22622: inst = 32'h10408000;
      22623: inst = 32'hc40432d;
      22624: inst = 32'h8220000;
      22625: inst = 32'h10408000;
      22626: inst = 32'hc40432e;
      22627: inst = 32'h8220000;
      22628: inst = 32'h10408000;
      22629: inst = 32'hc40432f;
      22630: inst = 32'h8220000;
      22631: inst = 32'h10408000;
      22632: inst = 32'hc404330;
      22633: inst = 32'h8220000;
      22634: inst = 32'h10408000;
      22635: inst = 32'hc404331;
      22636: inst = 32'h8220000;
      22637: inst = 32'h10408000;
      22638: inst = 32'hc404332;
      22639: inst = 32'h8220000;
      22640: inst = 32'h10408000;
      22641: inst = 32'hc404333;
      22642: inst = 32'h8220000;
      22643: inst = 32'h10408000;
      22644: inst = 32'hc404334;
      22645: inst = 32'h8220000;
      22646: inst = 32'h10408000;
      22647: inst = 32'hc404335;
      22648: inst = 32'h8220000;
      22649: inst = 32'h10408000;
      22650: inst = 32'hc404336;
      22651: inst = 32'h8220000;
      22652: inst = 32'h10408000;
      22653: inst = 32'hc405429;
      22654: inst = 32'h8220000;
      22655: inst = 32'h10408000;
      22656: inst = 32'hc40542a;
      22657: inst = 32'h8220000;
      22658: inst = 32'h10408000;
      22659: inst = 32'hc40542b;
      22660: inst = 32'h8220000;
      22661: inst = 32'h10408000;
      22662: inst = 32'hc40542c;
      22663: inst = 32'h8220000;
      22664: inst = 32'h10408000;
      22665: inst = 32'hc40542d;
      22666: inst = 32'h8220000;
      22667: inst = 32'h10408000;
      22668: inst = 32'hc40542e;
      22669: inst = 32'h8220000;
      22670: inst = 32'h10408000;
      22671: inst = 32'hc40542f;
      22672: inst = 32'h8220000;
      22673: inst = 32'h10408000;
      22674: inst = 32'hc405430;
      22675: inst = 32'h8220000;
      22676: inst = 32'h10408000;
      22677: inst = 32'hc405431;
      22678: inst = 32'h8220000;
      22679: inst = 32'h10408000;
      22680: inst = 32'hc405432;
      22681: inst = 32'h8220000;
      22682: inst = 32'h10408000;
      22683: inst = 32'hc405433;
      22684: inst = 32'h8220000;
      22685: inst = 32'h10408000;
      22686: inst = 32'hc405434;
      22687: inst = 32'h8220000;
      22688: inst = 32'h10408000;
      22689: inst = 32'hc405435;
      22690: inst = 32'h8220000;
      22691: inst = 32'h10408000;
      22692: inst = 32'hc405436;
      22693: inst = 32'h8220000;
      22694: inst = 32'h10408000;
      22695: inst = 32'hc405437;
      22696: inst = 32'h8220000;
      22697: inst = 32'h10408000;
      22698: inst = 32'hc405438;
      22699: inst = 32'h8220000;
      22700: inst = 32'h10408000;
      22701: inst = 32'hc405439;
      22702: inst = 32'h8220000;
      22703: inst = 32'h10408000;
      22704: inst = 32'hc40543a;
      22705: inst = 32'h8220000;
      22706: inst = 32'h10408000;
      22707: inst = 32'hc40543b;
      22708: inst = 32'h8220000;
      22709: inst = 32'h10408000;
      22710: inst = 32'hc40543c;
      22711: inst = 32'h8220000;
      22712: inst = 32'h10408000;
      22713: inst = 32'hc40543d;
      22714: inst = 32'h8220000;
      22715: inst = 32'h10408000;
      22716: inst = 32'hc40543e;
      22717: inst = 32'h8220000;
      22718: inst = 32'h10408000;
      22719: inst = 32'hc40543f;
      22720: inst = 32'h8220000;
      22721: inst = 32'h10408000;
      22722: inst = 32'hc405440;
      22723: inst = 32'h8220000;
      22724: inst = 32'h10408000;
      22725: inst = 32'hc405441;
      22726: inst = 32'h8220000;
      22727: inst = 32'h10408000;
      22728: inst = 32'hc405442;
      22729: inst = 32'h8220000;
      22730: inst = 32'h10408000;
      22731: inst = 32'hc405443;
      22732: inst = 32'h8220000;
      22733: inst = 32'h10408000;
      22734: inst = 32'hc405444;
      22735: inst = 32'h8220000;
      22736: inst = 32'h10408000;
      22737: inst = 32'hc405445;
      22738: inst = 32'h8220000;
      22739: inst = 32'h10408000;
      22740: inst = 32'hc405446;
      22741: inst = 32'h8220000;
      22742: inst = 32'h10408000;
      22743: inst = 32'hc405447;
      22744: inst = 32'h8220000;
      22745: inst = 32'h10408000;
      22746: inst = 32'hc405448;
      22747: inst = 32'h8220000;
      22748: inst = 32'h10408000;
      22749: inst = 32'hc405449;
      22750: inst = 32'h8220000;
      22751: inst = 32'h10408000;
      22752: inst = 32'hc40544a;
      22753: inst = 32'h8220000;
      22754: inst = 32'h10408000;
      22755: inst = 32'hc40544b;
      22756: inst = 32'h8220000;
      22757: inst = 32'h10408000;
      22758: inst = 32'hc40544c;
      22759: inst = 32'h8220000;
      22760: inst = 32'h10408000;
      22761: inst = 32'hc40544d;
      22762: inst = 32'h8220000;
      22763: inst = 32'h10408000;
      22764: inst = 32'hc40544e;
      22765: inst = 32'h8220000;
      22766: inst = 32'h10408000;
      22767: inst = 32'hc40544f;
      22768: inst = 32'h8220000;
      22769: inst = 32'h10408000;
      22770: inst = 32'hc405450;
      22771: inst = 32'h8220000;
      22772: inst = 32'h10408000;
      22773: inst = 32'hc405451;
      22774: inst = 32'h8220000;
      22775: inst = 32'h10408000;
      22776: inst = 32'hc405452;
      22777: inst = 32'h8220000;
      22778: inst = 32'h10408000;
      22779: inst = 32'hc405453;
      22780: inst = 32'h8220000;
      22781: inst = 32'h10408000;
      22782: inst = 32'hc405454;
      22783: inst = 32'h8220000;
      22784: inst = 32'h10408000;
      22785: inst = 32'hc405455;
      22786: inst = 32'h8220000;
      22787: inst = 32'h10408000;
      22788: inst = 32'hc405456;
      22789: inst = 32'h8220000;
      22790: inst = 32'h10408000;
      22791: inst = 32'hc405457;
      22792: inst = 32'h8220000;
      22793: inst = 32'h10408000;
      22794: inst = 32'hc405458;
      22795: inst = 32'h8220000;
      22796: inst = 32'h10408000;
      22797: inst = 32'hc405459;
      22798: inst = 32'h8220000;
      22799: inst = 32'h10408000;
      22800: inst = 32'hc40545a;
      22801: inst = 32'h8220000;
      22802: inst = 32'h10408000;
      22803: inst = 32'hc40545b;
      22804: inst = 32'h8220000;
      22805: inst = 32'h10408000;
      22806: inst = 32'hc40545c;
      22807: inst = 32'h8220000;
      22808: inst = 32'h10408000;
      22809: inst = 32'hc40545d;
      22810: inst = 32'h8220000;
      22811: inst = 32'h10408000;
      22812: inst = 32'hc40545e;
      22813: inst = 32'h8220000;
      22814: inst = 32'h10408000;
      22815: inst = 32'hc40545f;
      22816: inst = 32'h8220000;
      22817: inst = 32'h10408000;
      22818: inst = 32'hc405460;
      22819: inst = 32'h8220000;
      22820: inst = 32'h10408000;
      22821: inst = 32'hc405461;
      22822: inst = 32'h8220000;
      22823: inst = 32'h10408000;
      22824: inst = 32'hc405462;
      22825: inst = 32'h8220000;
      22826: inst = 32'h10408000;
      22827: inst = 32'hc405463;
      22828: inst = 32'h8220000;
      22829: inst = 32'h10408000;
      22830: inst = 32'hc405464;
      22831: inst = 32'h8220000;
      22832: inst = 32'h10408000;
      22833: inst = 32'hc405465;
      22834: inst = 32'h8220000;
      22835: inst = 32'h10408000;
      22836: inst = 32'hc405466;
      22837: inst = 32'h8220000;
      22838: inst = 32'h10408000;
      22839: inst = 32'hc405467;
      22840: inst = 32'h8220000;
      22841: inst = 32'h10408000;
      22842: inst = 32'hc405468;
      22843: inst = 32'h8220000;
      22844: inst = 32'h10408000;
      22845: inst = 32'hc405469;
      22846: inst = 32'h8220000;
      22847: inst = 32'h10408000;
      22848: inst = 32'hc40546a;
      22849: inst = 32'h8220000;
      22850: inst = 32'h10408000;
      22851: inst = 32'hc40546b;
      22852: inst = 32'h8220000;
      22853: inst = 32'h10408000;
      22854: inst = 32'hc40546c;
      22855: inst = 32'h8220000;
      22856: inst = 32'h10408000;
      22857: inst = 32'hc40546d;
      22858: inst = 32'h8220000;
      22859: inst = 32'h10408000;
      22860: inst = 32'hc40546e;
      22861: inst = 32'h8220000;
      22862: inst = 32'h10408000;
      22863: inst = 32'hc40546f;
      22864: inst = 32'h8220000;
      22865: inst = 32'h10408000;
      22866: inst = 32'hc405470;
      22867: inst = 32'h8220000;
      22868: inst = 32'h10408000;
      22869: inst = 32'hc405471;
      22870: inst = 32'h8220000;
      22871: inst = 32'h10408000;
      22872: inst = 32'hc405472;
      22873: inst = 32'h8220000;
      22874: inst = 32'h10408000;
      22875: inst = 32'hc405473;
      22876: inst = 32'h8220000;
      22877: inst = 32'h10408000;
      22878: inst = 32'hc405474;
      22879: inst = 32'h8220000;
      22880: inst = 32'h10408000;
      22881: inst = 32'hc405475;
      22882: inst = 32'h8220000;
      22883: inst = 32'h10408000;
      22884: inst = 32'hc405476;
      22885: inst = 32'h8220000;
      22886: inst = 32'hc202106;
      22887: inst = 32'h10408000;
      22888: inst = 32'hc404347;
      22889: inst = 32'h8220000;
      22890: inst = 32'h10408000;
      22891: inst = 32'hc404398;
      22892: inst = 32'h8220000;
      22893: inst = 32'h10408000;
      22894: inst = 32'hc4053c7;
      22895: inst = 32'h8220000;
      22896: inst = 32'h10408000;
      22897: inst = 32'hc405418;
      22898: inst = 32'h8220000;
      22899: inst = 32'hc2018c3;
      22900: inst = 32'h10408000;
      22901: inst = 32'hc404348;
      22902: inst = 32'h8220000;
      22903: inst = 32'h10408000;
      22904: inst = 32'hc404349;
      22905: inst = 32'h8220000;
      22906: inst = 32'h10408000;
      22907: inst = 32'hc40434a;
      22908: inst = 32'h8220000;
      22909: inst = 32'h10408000;
      22910: inst = 32'hc40434b;
      22911: inst = 32'h8220000;
      22912: inst = 32'h10408000;
      22913: inst = 32'hc40434c;
      22914: inst = 32'h8220000;
      22915: inst = 32'h10408000;
      22916: inst = 32'hc40434d;
      22917: inst = 32'h8220000;
      22918: inst = 32'h10408000;
      22919: inst = 32'hc40434e;
      22920: inst = 32'h8220000;
      22921: inst = 32'h10408000;
      22922: inst = 32'hc40434f;
      22923: inst = 32'h8220000;
      22924: inst = 32'h10408000;
      22925: inst = 32'hc404350;
      22926: inst = 32'h8220000;
      22927: inst = 32'h10408000;
      22928: inst = 32'hc404351;
      22929: inst = 32'h8220000;
      22930: inst = 32'h10408000;
      22931: inst = 32'hc404352;
      22932: inst = 32'h8220000;
      22933: inst = 32'h10408000;
      22934: inst = 32'hc404353;
      22935: inst = 32'h8220000;
      22936: inst = 32'h10408000;
      22937: inst = 32'hc404354;
      22938: inst = 32'h8220000;
      22939: inst = 32'h10408000;
      22940: inst = 32'hc404355;
      22941: inst = 32'h8220000;
      22942: inst = 32'h10408000;
      22943: inst = 32'hc404356;
      22944: inst = 32'h8220000;
      22945: inst = 32'h10408000;
      22946: inst = 32'hc404357;
      22947: inst = 32'h8220000;
      22948: inst = 32'h10408000;
      22949: inst = 32'hc404358;
      22950: inst = 32'h8220000;
      22951: inst = 32'h10408000;
      22952: inst = 32'hc404359;
      22953: inst = 32'h8220000;
      22954: inst = 32'h10408000;
      22955: inst = 32'hc40435a;
      22956: inst = 32'h8220000;
      22957: inst = 32'h10408000;
      22958: inst = 32'hc40435b;
      22959: inst = 32'h8220000;
      22960: inst = 32'h10408000;
      22961: inst = 32'hc40435c;
      22962: inst = 32'h8220000;
      22963: inst = 32'h10408000;
      22964: inst = 32'hc40435d;
      22965: inst = 32'h8220000;
      22966: inst = 32'h10408000;
      22967: inst = 32'hc40435e;
      22968: inst = 32'h8220000;
      22969: inst = 32'h10408000;
      22970: inst = 32'hc40435f;
      22971: inst = 32'h8220000;
      22972: inst = 32'h10408000;
      22973: inst = 32'hc404360;
      22974: inst = 32'h8220000;
      22975: inst = 32'h10408000;
      22976: inst = 32'hc404361;
      22977: inst = 32'h8220000;
      22978: inst = 32'h10408000;
      22979: inst = 32'hc404362;
      22980: inst = 32'h8220000;
      22981: inst = 32'h10408000;
      22982: inst = 32'hc404363;
      22983: inst = 32'h8220000;
      22984: inst = 32'h10408000;
      22985: inst = 32'hc404364;
      22986: inst = 32'h8220000;
      22987: inst = 32'h10408000;
      22988: inst = 32'hc404365;
      22989: inst = 32'h8220000;
      22990: inst = 32'h10408000;
      22991: inst = 32'hc404366;
      22992: inst = 32'h8220000;
      22993: inst = 32'h10408000;
      22994: inst = 32'hc404367;
      22995: inst = 32'h8220000;
      22996: inst = 32'h10408000;
      22997: inst = 32'hc404368;
      22998: inst = 32'h8220000;
      22999: inst = 32'h10408000;
      23000: inst = 32'hc404369;
      23001: inst = 32'h8220000;
      23002: inst = 32'h10408000;
      23003: inst = 32'hc40436a;
      23004: inst = 32'h8220000;
      23005: inst = 32'h10408000;
      23006: inst = 32'hc40436b;
      23007: inst = 32'h8220000;
      23008: inst = 32'h10408000;
      23009: inst = 32'hc40436c;
      23010: inst = 32'h8220000;
      23011: inst = 32'h10408000;
      23012: inst = 32'hc40436d;
      23013: inst = 32'h8220000;
      23014: inst = 32'h10408000;
      23015: inst = 32'hc40436e;
      23016: inst = 32'h8220000;
      23017: inst = 32'h10408000;
      23018: inst = 32'hc40436f;
      23019: inst = 32'h8220000;
      23020: inst = 32'h10408000;
      23021: inst = 32'hc404370;
      23022: inst = 32'h8220000;
      23023: inst = 32'h10408000;
      23024: inst = 32'hc404371;
      23025: inst = 32'h8220000;
      23026: inst = 32'h10408000;
      23027: inst = 32'hc404372;
      23028: inst = 32'h8220000;
      23029: inst = 32'h10408000;
      23030: inst = 32'hc404373;
      23031: inst = 32'h8220000;
      23032: inst = 32'h10408000;
      23033: inst = 32'hc404374;
      23034: inst = 32'h8220000;
      23035: inst = 32'h10408000;
      23036: inst = 32'hc404375;
      23037: inst = 32'h8220000;
      23038: inst = 32'h10408000;
      23039: inst = 32'hc404376;
      23040: inst = 32'h8220000;
      23041: inst = 32'h10408000;
      23042: inst = 32'hc404377;
      23043: inst = 32'h8220000;
      23044: inst = 32'h10408000;
      23045: inst = 32'hc404378;
      23046: inst = 32'h8220000;
      23047: inst = 32'h10408000;
      23048: inst = 32'hc404379;
      23049: inst = 32'h8220000;
      23050: inst = 32'h10408000;
      23051: inst = 32'hc40437a;
      23052: inst = 32'h8220000;
      23053: inst = 32'h10408000;
      23054: inst = 32'hc40437b;
      23055: inst = 32'h8220000;
      23056: inst = 32'h10408000;
      23057: inst = 32'hc40437c;
      23058: inst = 32'h8220000;
      23059: inst = 32'h10408000;
      23060: inst = 32'hc40437d;
      23061: inst = 32'h8220000;
      23062: inst = 32'h10408000;
      23063: inst = 32'hc40437e;
      23064: inst = 32'h8220000;
      23065: inst = 32'h10408000;
      23066: inst = 32'hc40437f;
      23067: inst = 32'h8220000;
      23068: inst = 32'h10408000;
      23069: inst = 32'hc404380;
      23070: inst = 32'h8220000;
      23071: inst = 32'h10408000;
      23072: inst = 32'hc404381;
      23073: inst = 32'h8220000;
      23074: inst = 32'h10408000;
      23075: inst = 32'hc404382;
      23076: inst = 32'h8220000;
      23077: inst = 32'h10408000;
      23078: inst = 32'hc404383;
      23079: inst = 32'h8220000;
      23080: inst = 32'h10408000;
      23081: inst = 32'hc404384;
      23082: inst = 32'h8220000;
      23083: inst = 32'h10408000;
      23084: inst = 32'hc404385;
      23085: inst = 32'h8220000;
      23086: inst = 32'h10408000;
      23087: inst = 32'hc404386;
      23088: inst = 32'h8220000;
      23089: inst = 32'h10408000;
      23090: inst = 32'hc404387;
      23091: inst = 32'h8220000;
      23092: inst = 32'h10408000;
      23093: inst = 32'hc404388;
      23094: inst = 32'h8220000;
      23095: inst = 32'h10408000;
      23096: inst = 32'hc404389;
      23097: inst = 32'h8220000;
      23098: inst = 32'h10408000;
      23099: inst = 32'hc40438a;
      23100: inst = 32'h8220000;
      23101: inst = 32'h10408000;
      23102: inst = 32'hc40438b;
      23103: inst = 32'h8220000;
      23104: inst = 32'h10408000;
      23105: inst = 32'hc40438c;
      23106: inst = 32'h8220000;
      23107: inst = 32'h10408000;
      23108: inst = 32'hc40438d;
      23109: inst = 32'h8220000;
      23110: inst = 32'h10408000;
      23111: inst = 32'hc40438e;
      23112: inst = 32'h8220000;
      23113: inst = 32'h10408000;
      23114: inst = 32'hc40438f;
      23115: inst = 32'h8220000;
      23116: inst = 32'h10408000;
      23117: inst = 32'hc404390;
      23118: inst = 32'h8220000;
      23119: inst = 32'h10408000;
      23120: inst = 32'hc404391;
      23121: inst = 32'h8220000;
      23122: inst = 32'h10408000;
      23123: inst = 32'hc404392;
      23124: inst = 32'h8220000;
      23125: inst = 32'h10408000;
      23126: inst = 32'hc404393;
      23127: inst = 32'h8220000;
      23128: inst = 32'h10408000;
      23129: inst = 32'hc404394;
      23130: inst = 32'h8220000;
      23131: inst = 32'h10408000;
      23132: inst = 32'hc404395;
      23133: inst = 32'h8220000;
      23134: inst = 32'h10408000;
      23135: inst = 32'hc404396;
      23136: inst = 32'h8220000;
      23137: inst = 32'h10408000;
      23138: inst = 32'hc404397;
      23139: inst = 32'h8220000;
      23140: inst = 32'h10408000;
      23141: inst = 32'hc4043a7;
      23142: inst = 32'h8220000;
      23143: inst = 32'h10408000;
      23144: inst = 32'hc4043a8;
      23145: inst = 32'h8220000;
      23146: inst = 32'h10408000;
      23147: inst = 32'hc4043a9;
      23148: inst = 32'h8220000;
      23149: inst = 32'h10408000;
      23150: inst = 32'hc4043aa;
      23151: inst = 32'h8220000;
      23152: inst = 32'h10408000;
      23153: inst = 32'hc4043ab;
      23154: inst = 32'h8220000;
      23155: inst = 32'h10408000;
      23156: inst = 32'hc4043ac;
      23157: inst = 32'h8220000;
      23158: inst = 32'h10408000;
      23159: inst = 32'hc4043ad;
      23160: inst = 32'h8220000;
      23161: inst = 32'h10408000;
      23162: inst = 32'hc4043ae;
      23163: inst = 32'h8220000;
      23164: inst = 32'h10408000;
      23165: inst = 32'hc4043af;
      23166: inst = 32'h8220000;
      23167: inst = 32'h10408000;
      23168: inst = 32'hc4043b0;
      23169: inst = 32'h8220000;
      23170: inst = 32'h10408000;
      23171: inst = 32'hc4043b1;
      23172: inst = 32'h8220000;
      23173: inst = 32'h10408000;
      23174: inst = 32'hc4043b2;
      23175: inst = 32'h8220000;
      23176: inst = 32'h10408000;
      23177: inst = 32'hc4043b3;
      23178: inst = 32'h8220000;
      23179: inst = 32'h10408000;
      23180: inst = 32'hc4043b4;
      23181: inst = 32'h8220000;
      23182: inst = 32'h10408000;
      23183: inst = 32'hc4043b5;
      23184: inst = 32'h8220000;
      23185: inst = 32'h10408000;
      23186: inst = 32'hc4043b6;
      23187: inst = 32'h8220000;
      23188: inst = 32'h10408000;
      23189: inst = 32'hc4043b7;
      23190: inst = 32'h8220000;
      23191: inst = 32'h10408000;
      23192: inst = 32'hc4043b8;
      23193: inst = 32'h8220000;
      23194: inst = 32'h10408000;
      23195: inst = 32'hc4043b9;
      23196: inst = 32'h8220000;
      23197: inst = 32'h10408000;
      23198: inst = 32'hc4043ba;
      23199: inst = 32'h8220000;
      23200: inst = 32'h10408000;
      23201: inst = 32'hc4043bb;
      23202: inst = 32'h8220000;
      23203: inst = 32'h10408000;
      23204: inst = 32'hc4043bc;
      23205: inst = 32'h8220000;
      23206: inst = 32'h10408000;
      23207: inst = 32'hc4043bd;
      23208: inst = 32'h8220000;
      23209: inst = 32'h10408000;
      23210: inst = 32'hc4043be;
      23211: inst = 32'h8220000;
      23212: inst = 32'h10408000;
      23213: inst = 32'hc4043bf;
      23214: inst = 32'h8220000;
      23215: inst = 32'h10408000;
      23216: inst = 32'hc4043c0;
      23217: inst = 32'h8220000;
      23218: inst = 32'h10408000;
      23219: inst = 32'hc4043c1;
      23220: inst = 32'h8220000;
      23221: inst = 32'h10408000;
      23222: inst = 32'hc4043c2;
      23223: inst = 32'h8220000;
      23224: inst = 32'h10408000;
      23225: inst = 32'hc4043c3;
      23226: inst = 32'h8220000;
      23227: inst = 32'h10408000;
      23228: inst = 32'hc4043c4;
      23229: inst = 32'h8220000;
      23230: inst = 32'h10408000;
      23231: inst = 32'hc4043c5;
      23232: inst = 32'h8220000;
      23233: inst = 32'h10408000;
      23234: inst = 32'hc4043c6;
      23235: inst = 32'h8220000;
      23236: inst = 32'h10408000;
      23237: inst = 32'hc4043c7;
      23238: inst = 32'h8220000;
      23239: inst = 32'h10408000;
      23240: inst = 32'hc4043c8;
      23241: inst = 32'h8220000;
      23242: inst = 32'h10408000;
      23243: inst = 32'hc4043c9;
      23244: inst = 32'h8220000;
      23245: inst = 32'h10408000;
      23246: inst = 32'hc4043ca;
      23247: inst = 32'h8220000;
      23248: inst = 32'h10408000;
      23249: inst = 32'hc4043cb;
      23250: inst = 32'h8220000;
      23251: inst = 32'h10408000;
      23252: inst = 32'hc4043cc;
      23253: inst = 32'h8220000;
      23254: inst = 32'h10408000;
      23255: inst = 32'hc4043cd;
      23256: inst = 32'h8220000;
      23257: inst = 32'h10408000;
      23258: inst = 32'hc4043ce;
      23259: inst = 32'h8220000;
      23260: inst = 32'h10408000;
      23261: inst = 32'hc4043cf;
      23262: inst = 32'h8220000;
      23263: inst = 32'h10408000;
      23264: inst = 32'hc4043d0;
      23265: inst = 32'h8220000;
      23266: inst = 32'h10408000;
      23267: inst = 32'hc4043d1;
      23268: inst = 32'h8220000;
      23269: inst = 32'h10408000;
      23270: inst = 32'hc4043d2;
      23271: inst = 32'h8220000;
      23272: inst = 32'h10408000;
      23273: inst = 32'hc4043d3;
      23274: inst = 32'h8220000;
      23275: inst = 32'h10408000;
      23276: inst = 32'hc4043d4;
      23277: inst = 32'h8220000;
      23278: inst = 32'h10408000;
      23279: inst = 32'hc4043d5;
      23280: inst = 32'h8220000;
      23281: inst = 32'h10408000;
      23282: inst = 32'hc4043d6;
      23283: inst = 32'h8220000;
      23284: inst = 32'h10408000;
      23285: inst = 32'hc4043d7;
      23286: inst = 32'h8220000;
      23287: inst = 32'h10408000;
      23288: inst = 32'hc4043d8;
      23289: inst = 32'h8220000;
      23290: inst = 32'h10408000;
      23291: inst = 32'hc4043d9;
      23292: inst = 32'h8220000;
      23293: inst = 32'h10408000;
      23294: inst = 32'hc4043da;
      23295: inst = 32'h8220000;
      23296: inst = 32'h10408000;
      23297: inst = 32'hc4043db;
      23298: inst = 32'h8220000;
      23299: inst = 32'h10408000;
      23300: inst = 32'hc4043dc;
      23301: inst = 32'h8220000;
      23302: inst = 32'h10408000;
      23303: inst = 32'hc4043dd;
      23304: inst = 32'h8220000;
      23305: inst = 32'h10408000;
      23306: inst = 32'hc4043de;
      23307: inst = 32'h8220000;
      23308: inst = 32'h10408000;
      23309: inst = 32'hc4043df;
      23310: inst = 32'h8220000;
      23311: inst = 32'h10408000;
      23312: inst = 32'hc4043e0;
      23313: inst = 32'h8220000;
      23314: inst = 32'h10408000;
      23315: inst = 32'hc4043e1;
      23316: inst = 32'h8220000;
      23317: inst = 32'h10408000;
      23318: inst = 32'hc4043e2;
      23319: inst = 32'h8220000;
      23320: inst = 32'h10408000;
      23321: inst = 32'hc4043e3;
      23322: inst = 32'h8220000;
      23323: inst = 32'h10408000;
      23324: inst = 32'hc4043e4;
      23325: inst = 32'h8220000;
      23326: inst = 32'h10408000;
      23327: inst = 32'hc4043e5;
      23328: inst = 32'h8220000;
      23329: inst = 32'h10408000;
      23330: inst = 32'hc4043e6;
      23331: inst = 32'h8220000;
      23332: inst = 32'h10408000;
      23333: inst = 32'hc4043e7;
      23334: inst = 32'h8220000;
      23335: inst = 32'h10408000;
      23336: inst = 32'hc4043e8;
      23337: inst = 32'h8220000;
      23338: inst = 32'h10408000;
      23339: inst = 32'hc4043e9;
      23340: inst = 32'h8220000;
      23341: inst = 32'h10408000;
      23342: inst = 32'hc4043ea;
      23343: inst = 32'h8220000;
      23344: inst = 32'h10408000;
      23345: inst = 32'hc4043eb;
      23346: inst = 32'h8220000;
      23347: inst = 32'h10408000;
      23348: inst = 32'hc4043ec;
      23349: inst = 32'h8220000;
      23350: inst = 32'h10408000;
      23351: inst = 32'hc4043ed;
      23352: inst = 32'h8220000;
      23353: inst = 32'h10408000;
      23354: inst = 32'hc4043ee;
      23355: inst = 32'h8220000;
      23356: inst = 32'h10408000;
      23357: inst = 32'hc4043ef;
      23358: inst = 32'h8220000;
      23359: inst = 32'h10408000;
      23360: inst = 32'hc4043f0;
      23361: inst = 32'h8220000;
      23362: inst = 32'h10408000;
      23363: inst = 32'hc4043f1;
      23364: inst = 32'h8220000;
      23365: inst = 32'h10408000;
      23366: inst = 32'hc4043f2;
      23367: inst = 32'h8220000;
      23368: inst = 32'h10408000;
      23369: inst = 32'hc4043f3;
      23370: inst = 32'h8220000;
      23371: inst = 32'h10408000;
      23372: inst = 32'hc4043f4;
      23373: inst = 32'h8220000;
      23374: inst = 32'h10408000;
      23375: inst = 32'hc4043f5;
      23376: inst = 32'h8220000;
      23377: inst = 32'h10408000;
      23378: inst = 32'hc4043f6;
      23379: inst = 32'h8220000;
      23380: inst = 32'h10408000;
      23381: inst = 32'hc4043f7;
      23382: inst = 32'h8220000;
      23383: inst = 32'h10408000;
      23384: inst = 32'hc4043f8;
      23385: inst = 32'h8220000;
      23386: inst = 32'h10408000;
      23387: inst = 32'hc404407;
      23388: inst = 32'h8220000;
      23389: inst = 32'h10408000;
      23390: inst = 32'hc404408;
      23391: inst = 32'h8220000;
      23392: inst = 32'h10408000;
      23393: inst = 32'hc404409;
      23394: inst = 32'h8220000;
      23395: inst = 32'h10408000;
      23396: inst = 32'hc40440a;
      23397: inst = 32'h8220000;
      23398: inst = 32'h10408000;
      23399: inst = 32'hc40440b;
      23400: inst = 32'h8220000;
      23401: inst = 32'h10408000;
      23402: inst = 32'hc40440c;
      23403: inst = 32'h8220000;
      23404: inst = 32'h10408000;
      23405: inst = 32'hc40440d;
      23406: inst = 32'h8220000;
      23407: inst = 32'h10408000;
      23408: inst = 32'hc40440e;
      23409: inst = 32'h8220000;
      23410: inst = 32'h10408000;
      23411: inst = 32'hc40440f;
      23412: inst = 32'h8220000;
      23413: inst = 32'h10408000;
      23414: inst = 32'hc404410;
      23415: inst = 32'h8220000;
      23416: inst = 32'h10408000;
      23417: inst = 32'hc404411;
      23418: inst = 32'h8220000;
      23419: inst = 32'h10408000;
      23420: inst = 32'hc404412;
      23421: inst = 32'h8220000;
      23422: inst = 32'h10408000;
      23423: inst = 32'hc404413;
      23424: inst = 32'h8220000;
      23425: inst = 32'h10408000;
      23426: inst = 32'hc404414;
      23427: inst = 32'h8220000;
      23428: inst = 32'h10408000;
      23429: inst = 32'hc404415;
      23430: inst = 32'h8220000;
      23431: inst = 32'h10408000;
      23432: inst = 32'hc404416;
      23433: inst = 32'h8220000;
      23434: inst = 32'h10408000;
      23435: inst = 32'hc404417;
      23436: inst = 32'h8220000;
      23437: inst = 32'h10408000;
      23438: inst = 32'hc404418;
      23439: inst = 32'h8220000;
      23440: inst = 32'h10408000;
      23441: inst = 32'hc404419;
      23442: inst = 32'h8220000;
      23443: inst = 32'h10408000;
      23444: inst = 32'hc40441a;
      23445: inst = 32'h8220000;
      23446: inst = 32'h10408000;
      23447: inst = 32'hc40441b;
      23448: inst = 32'h8220000;
      23449: inst = 32'h10408000;
      23450: inst = 32'hc40441c;
      23451: inst = 32'h8220000;
      23452: inst = 32'h10408000;
      23453: inst = 32'hc40441d;
      23454: inst = 32'h8220000;
      23455: inst = 32'h10408000;
      23456: inst = 32'hc40441e;
      23457: inst = 32'h8220000;
      23458: inst = 32'h10408000;
      23459: inst = 32'hc40441f;
      23460: inst = 32'h8220000;
      23461: inst = 32'h10408000;
      23462: inst = 32'hc404420;
      23463: inst = 32'h8220000;
      23464: inst = 32'h10408000;
      23465: inst = 32'hc404421;
      23466: inst = 32'h8220000;
      23467: inst = 32'h10408000;
      23468: inst = 32'hc404422;
      23469: inst = 32'h8220000;
      23470: inst = 32'h10408000;
      23471: inst = 32'hc404423;
      23472: inst = 32'h8220000;
      23473: inst = 32'h10408000;
      23474: inst = 32'hc404424;
      23475: inst = 32'h8220000;
      23476: inst = 32'h10408000;
      23477: inst = 32'hc404425;
      23478: inst = 32'h8220000;
      23479: inst = 32'h10408000;
      23480: inst = 32'hc404426;
      23481: inst = 32'h8220000;
      23482: inst = 32'h10408000;
      23483: inst = 32'hc404427;
      23484: inst = 32'h8220000;
      23485: inst = 32'h10408000;
      23486: inst = 32'hc404428;
      23487: inst = 32'h8220000;
      23488: inst = 32'h10408000;
      23489: inst = 32'hc404429;
      23490: inst = 32'h8220000;
      23491: inst = 32'h10408000;
      23492: inst = 32'hc40442a;
      23493: inst = 32'h8220000;
      23494: inst = 32'h10408000;
      23495: inst = 32'hc40442b;
      23496: inst = 32'h8220000;
      23497: inst = 32'h10408000;
      23498: inst = 32'hc40442c;
      23499: inst = 32'h8220000;
      23500: inst = 32'h10408000;
      23501: inst = 32'hc40442d;
      23502: inst = 32'h8220000;
      23503: inst = 32'h10408000;
      23504: inst = 32'hc40442e;
      23505: inst = 32'h8220000;
      23506: inst = 32'h10408000;
      23507: inst = 32'hc40442f;
      23508: inst = 32'h8220000;
      23509: inst = 32'h10408000;
      23510: inst = 32'hc404430;
      23511: inst = 32'h8220000;
      23512: inst = 32'h10408000;
      23513: inst = 32'hc404431;
      23514: inst = 32'h8220000;
      23515: inst = 32'h10408000;
      23516: inst = 32'hc404432;
      23517: inst = 32'h8220000;
      23518: inst = 32'h10408000;
      23519: inst = 32'hc404433;
      23520: inst = 32'h8220000;
      23521: inst = 32'h10408000;
      23522: inst = 32'hc404434;
      23523: inst = 32'h8220000;
      23524: inst = 32'h10408000;
      23525: inst = 32'hc404435;
      23526: inst = 32'h8220000;
      23527: inst = 32'h10408000;
      23528: inst = 32'hc404436;
      23529: inst = 32'h8220000;
      23530: inst = 32'h10408000;
      23531: inst = 32'hc404437;
      23532: inst = 32'h8220000;
      23533: inst = 32'h10408000;
      23534: inst = 32'hc404438;
      23535: inst = 32'h8220000;
      23536: inst = 32'h10408000;
      23537: inst = 32'hc404439;
      23538: inst = 32'h8220000;
      23539: inst = 32'h10408000;
      23540: inst = 32'hc40443a;
      23541: inst = 32'h8220000;
      23542: inst = 32'h10408000;
      23543: inst = 32'hc40443b;
      23544: inst = 32'h8220000;
      23545: inst = 32'h10408000;
      23546: inst = 32'hc40443c;
      23547: inst = 32'h8220000;
      23548: inst = 32'h10408000;
      23549: inst = 32'hc40443d;
      23550: inst = 32'h8220000;
      23551: inst = 32'h10408000;
      23552: inst = 32'hc40443e;
      23553: inst = 32'h8220000;
      23554: inst = 32'h10408000;
      23555: inst = 32'hc40443f;
      23556: inst = 32'h8220000;
      23557: inst = 32'h10408000;
      23558: inst = 32'hc404440;
      23559: inst = 32'h8220000;
      23560: inst = 32'h10408000;
      23561: inst = 32'hc404441;
      23562: inst = 32'h8220000;
      23563: inst = 32'h10408000;
      23564: inst = 32'hc404442;
      23565: inst = 32'h8220000;
      23566: inst = 32'h10408000;
      23567: inst = 32'hc404443;
      23568: inst = 32'h8220000;
      23569: inst = 32'h10408000;
      23570: inst = 32'hc404444;
      23571: inst = 32'h8220000;
      23572: inst = 32'h10408000;
      23573: inst = 32'hc404445;
      23574: inst = 32'h8220000;
      23575: inst = 32'h10408000;
      23576: inst = 32'hc404446;
      23577: inst = 32'h8220000;
      23578: inst = 32'h10408000;
      23579: inst = 32'hc404447;
      23580: inst = 32'h8220000;
      23581: inst = 32'h10408000;
      23582: inst = 32'hc404448;
      23583: inst = 32'h8220000;
      23584: inst = 32'h10408000;
      23585: inst = 32'hc404449;
      23586: inst = 32'h8220000;
      23587: inst = 32'h10408000;
      23588: inst = 32'hc40444a;
      23589: inst = 32'h8220000;
      23590: inst = 32'h10408000;
      23591: inst = 32'hc40444b;
      23592: inst = 32'h8220000;
      23593: inst = 32'h10408000;
      23594: inst = 32'hc40444c;
      23595: inst = 32'h8220000;
      23596: inst = 32'h10408000;
      23597: inst = 32'hc40444d;
      23598: inst = 32'h8220000;
      23599: inst = 32'h10408000;
      23600: inst = 32'hc40444e;
      23601: inst = 32'h8220000;
      23602: inst = 32'h10408000;
      23603: inst = 32'hc40444f;
      23604: inst = 32'h8220000;
      23605: inst = 32'h10408000;
      23606: inst = 32'hc404450;
      23607: inst = 32'h8220000;
      23608: inst = 32'h10408000;
      23609: inst = 32'hc404451;
      23610: inst = 32'h8220000;
      23611: inst = 32'h10408000;
      23612: inst = 32'hc404452;
      23613: inst = 32'h8220000;
      23614: inst = 32'h10408000;
      23615: inst = 32'hc404453;
      23616: inst = 32'h8220000;
      23617: inst = 32'h10408000;
      23618: inst = 32'hc404454;
      23619: inst = 32'h8220000;
      23620: inst = 32'h10408000;
      23621: inst = 32'hc404455;
      23622: inst = 32'h8220000;
      23623: inst = 32'h10408000;
      23624: inst = 32'hc404456;
      23625: inst = 32'h8220000;
      23626: inst = 32'h10408000;
      23627: inst = 32'hc404457;
      23628: inst = 32'h8220000;
      23629: inst = 32'h10408000;
      23630: inst = 32'hc404458;
      23631: inst = 32'h8220000;
      23632: inst = 32'h10408000;
      23633: inst = 32'hc404467;
      23634: inst = 32'h8220000;
      23635: inst = 32'h10408000;
      23636: inst = 32'hc404468;
      23637: inst = 32'h8220000;
      23638: inst = 32'h10408000;
      23639: inst = 32'hc404469;
      23640: inst = 32'h8220000;
      23641: inst = 32'h10408000;
      23642: inst = 32'hc40446a;
      23643: inst = 32'h8220000;
      23644: inst = 32'h10408000;
      23645: inst = 32'hc40446b;
      23646: inst = 32'h8220000;
      23647: inst = 32'h10408000;
      23648: inst = 32'hc40446c;
      23649: inst = 32'h8220000;
      23650: inst = 32'h10408000;
      23651: inst = 32'hc40446d;
      23652: inst = 32'h8220000;
      23653: inst = 32'h10408000;
      23654: inst = 32'hc40446e;
      23655: inst = 32'h8220000;
      23656: inst = 32'h10408000;
      23657: inst = 32'hc40446f;
      23658: inst = 32'h8220000;
      23659: inst = 32'h10408000;
      23660: inst = 32'hc404470;
      23661: inst = 32'h8220000;
      23662: inst = 32'h10408000;
      23663: inst = 32'hc404471;
      23664: inst = 32'h8220000;
      23665: inst = 32'h10408000;
      23666: inst = 32'hc404472;
      23667: inst = 32'h8220000;
      23668: inst = 32'h10408000;
      23669: inst = 32'hc404473;
      23670: inst = 32'h8220000;
      23671: inst = 32'h10408000;
      23672: inst = 32'hc404474;
      23673: inst = 32'h8220000;
      23674: inst = 32'h10408000;
      23675: inst = 32'hc404475;
      23676: inst = 32'h8220000;
      23677: inst = 32'h10408000;
      23678: inst = 32'hc404476;
      23679: inst = 32'h8220000;
      23680: inst = 32'h10408000;
      23681: inst = 32'hc404477;
      23682: inst = 32'h8220000;
      23683: inst = 32'h10408000;
      23684: inst = 32'hc404478;
      23685: inst = 32'h8220000;
      23686: inst = 32'h10408000;
      23687: inst = 32'hc404479;
      23688: inst = 32'h8220000;
      23689: inst = 32'h10408000;
      23690: inst = 32'hc40447a;
      23691: inst = 32'h8220000;
      23692: inst = 32'h10408000;
      23693: inst = 32'hc40447b;
      23694: inst = 32'h8220000;
      23695: inst = 32'h10408000;
      23696: inst = 32'hc40447c;
      23697: inst = 32'h8220000;
      23698: inst = 32'h10408000;
      23699: inst = 32'hc40447d;
      23700: inst = 32'h8220000;
      23701: inst = 32'h10408000;
      23702: inst = 32'hc40447e;
      23703: inst = 32'h8220000;
      23704: inst = 32'h10408000;
      23705: inst = 32'hc40447f;
      23706: inst = 32'h8220000;
      23707: inst = 32'h10408000;
      23708: inst = 32'hc404480;
      23709: inst = 32'h8220000;
      23710: inst = 32'h10408000;
      23711: inst = 32'hc404481;
      23712: inst = 32'h8220000;
      23713: inst = 32'h10408000;
      23714: inst = 32'hc404482;
      23715: inst = 32'h8220000;
      23716: inst = 32'h10408000;
      23717: inst = 32'hc404483;
      23718: inst = 32'h8220000;
      23719: inst = 32'h10408000;
      23720: inst = 32'hc404484;
      23721: inst = 32'h8220000;
      23722: inst = 32'h10408000;
      23723: inst = 32'hc404485;
      23724: inst = 32'h8220000;
      23725: inst = 32'h10408000;
      23726: inst = 32'hc404486;
      23727: inst = 32'h8220000;
      23728: inst = 32'h10408000;
      23729: inst = 32'hc404487;
      23730: inst = 32'h8220000;
      23731: inst = 32'h10408000;
      23732: inst = 32'hc404488;
      23733: inst = 32'h8220000;
      23734: inst = 32'h10408000;
      23735: inst = 32'hc404489;
      23736: inst = 32'h8220000;
      23737: inst = 32'h10408000;
      23738: inst = 32'hc40448a;
      23739: inst = 32'h8220000;
      23740: inst = 32'h10408000;
      23741: inst = 32'hc40448b;
      23742: inst = 32'h8220000;
      23743: inst = 32'h10408000;
      23744: inst = 32'hc40448c;
      23745: inst = 32'h8220000;
      23746: inst = 32'h10408000;
      23747: inst = 32'hc40448d;
      23748: inst = 32'h8220000;
      23749: inst = 32'h10408000;
      23750: inst = 32'hc40448e;
      23751: inst = 32'h8220000;
      23752: inst = 32'h10408000;
      23753: inst = 32'hc40448f;
      23754: inst = 32'h8220000;
      23755: inst = 32'h10408000;
      23756: inst = 32'hc404490;
      23757: inst = 32'h8220000;
      23758: inst = 32'h10408000;
      23759: inst = 32'hc404491;
      23760: inst = 32'h8220000;
      23761: inst = 32'h10408000;
      23762: inst = 32'hc404492;
      23763: inst = 32'h8220000;
      23764: inst = 32'h10408000;
      23765: inst = 32'hc404493;
      23766: inst = 32'h8220000;
      23767: inst = 32'h10408000;
      23768: inst = 32'hc404494;
      23769: inst = 32'h8220000;
      23770: inst = 32'h10408000;
      23771: inst = 32'hc404495;
      23772: inst = 32'h8220000;
      23773: inst = 32'h10408000;
      23774: inst = 32'hc404496;
      23775: inst = 32'h8220000;
      23776: inst = 32'h10408000;
      23777: inst = 32'hc404497;
      23778: inst = 32'h8220000;
      23779: inst = 32'h10408000;
      23780: inst = 32'hc404498;
      23781: inst = 32'h8220000;
      23782: inst = 32'h10408000;
      23783: inst = 32'hc404499;
      23784: inst = 32'h8220000;
      23785: inst = 32'h10408000;
      23786: inst = 32'hc40449a;
      23787: inst = 32'h8220000;
      23788: inst = 32'h10408000;
      23789: inst = 32'hc40449b;
      23790: inst = 32'h8220000;
      23791: inst = 32'h10408000;
      23792: inst = 32'hc40449c;
      23793: inst = 32'h8220000;
      23794: inst = 32'h10408000;
      23795: inst = 32'hc40449d;
      23796: inst = 32'h8220000;
      23797: inst = 32'h10408000;
      23798: inst = 32'hc40449e;
      23799: inst = 32'h8220000;
      23800: inst = 32'h10408000;
      23801: inst = 32'hc40449f;
      23802: inst = 32'h8220000;
      23803: inst = 32'h10408000;
      23804: inst = 32'hc4044a0;
      23805: inst = 32'h8220000;
      23806: inst = 32'h10408000;
      23807: inst = 32'hc4044a1;
      23808: inst = 32'h8220000;
      23809: inst = 32'h10408000;
      23810: inst = 32'hc4044a2;
      23811: inst = 32'h8220000;
      23812: inst = 32'h10408000;
      23813: inst = 32'hc4044a3;
      23814: inst = 32'h8220000;
      23815: inst = 32'h10408000;
      23816: inst = 32'hc4044a4;
      23817: inst = 32'h8220000;
      23818: inst = 32'h10408000;
      23819: inst = 32'hc4044a5;
      23820: inst = 32'h8220000;
      23821: inst = 32'h10408000;
      23822: inst = 32'hc4044a6;
      23823: inst = 32'h8220000;
      23824: inst = 32'h10408000;
      23825: inst = 32'hc4044a7;
      23826: inst = 32'h8220000;
      23827: inst = 32'h10408000;
      23828: inst = 32'hc4044a8;
      23829: inst = 32'h8220000;
      23830: inst = 32'h10408000;
      23831: inst = 32'hc4044a9;
      23832: inst = 32'h8220000;
      23833: inst = 32'h10408000;
      23834: inst = 32'hc4044aa;
      23835: inst = 32'h8220000;
      23836: inst = 32'h10408000;
      23837: inst = 32'hc4044ab;
      23838: inst = 32'h8220000;
      23839: inst = 32'h10408000;
      23840: inst = 32'hc4044ac;
      23841: inst = 32'h8220000;
      23842: inst = 32'h10408000;
      23843: inst = 32'hc4044ad;
      23844: inst = 32'h8220000;
      23845: inst = 32'h10408000;
      23846: inst = 32'hc4044ae;
      23847: inst = 32'h8220000;
      23848: inst = 32'h10408000;
      23849: inst = 32'hc4044af;
      23850: inst = 32'h8220000;
      23851: inst = 32'h10408000;
      23852: inst = 32'hc4044b0;
      23853: inst = 32'h8220000;
      23854: inst = 32'h10408000;
      23855: inst = 32'hc4044b1;
      23856: inst = 32'h8220000;
      23857: inst = 32'h10408000;
      23858: inst = 32'hc4044b2;
      23859: inst = 32'h8220000;
      23860: inst = 32'h10408000;
      23861: inst = 32'hc4044b3;
      23862: inst = 32'h8220000;
      23863: inst = 32'h10408000;
      23864: inst = 32'hc4044b4;
      23865: inst = 32'h8220000;
      23866: inst = 32'h10408000;
      23867: inst = 32'hc4044b5;
      23868: inst = 32'h8220000;
      23869: inst = 32'h10408000;
      23870: inst = 32'hc4044b6;
      23871: inst = 32'h8220000;
      23872: inst = 32'h10408000;
      23873: inst = 32'hc4044b7;
      23874: inst = 32'h8220000;
      23875: inst = 32'h10408000;
      23876: inst = 32'hc4044b8;
      23877: inst = 32'h8220000;
      23878: inst = 32'h10408000;
      23879: inst = 32'hc4044c7;
      23880: inst = 32'h8220000;
      23881: inst = 32'h10408000;
      23882: inst = 32'hc4044c8;
      23883: inst = 32'h8220000;
      23884: inst = 32'h10408000;
      23885: inst = 32'hc4044c9;
      23886: inst = 32'h8220000;
      23887: inst = 32'h10408000;
      23888: inst = 32'hc4044ca;
      23889: inst = 32'h8220000;
      23890: inst = 32'h10408000;
      23891: inst = 32'hc4044cb;
      23892: inst = 32'h8220000;
      23893: inst = 32'h10408000;
      23894: inst = 32'hc4044cc;
      23895: inst = 32'h8220000;
      23896: inst = 32'h10408000;
      23897: inst = 32'hc4044cd;
      23898: inst = 32'h8220000;
      23899: inst = 32'h10408000;
      23900: inst = 32'hc4044ce;
      23901: inst = 32'h8220000;
      23902: inst = 32'h10408000;
      23903: inst = 32'hc4044cf;
      23904: inst = 32'h8220000;
      23905: inst = 32'h10408000;
      23906: inst = 32'hc4044d0;
      23907: inst = 32'h8220000;
      23908: inst = 32'h10408000;
      23909: inst = 32'hc4044d1;
      23910: inst = 32'h8220000;
      23911: inst = 32'h10408000;
      23912: inst = 32'hc4044d2;
      23913: inst = 32'h8220000;
      23914: inst = 32'h10408000;
      23915: inst = 32'hc4044d3;
      23916: inst = 32'h8220000;
      23917: inst = 32'h10408000;
      23918: inst = 32'hc4044d4;
      23919: inst = 32'h8220000;
      23920: inst = 32'h10408000;
      23921: inst = 32'hc4044d5;
      23922: inst = 32'h8220000;
      23923: inst = 32'h10408000;
      23924: inst = 32'hc4044d6;
      23925: inst = 32'h8220000;
      23926: inst = 32'h10408000;
      23927: inst = 32'hc4044d7;
      23928: inst = 32'h8220000;
      23929: inst = 32'h10408000;
      23930: inst = 32'hc4044d8;
      23931: inst = 32'h8220000;
      23932: inst = 32'h10408000;
      23933: inst = 32'hc4044d9;
      23934: inst = 32'h8220000;
      23935: inst = 32'h10408000;
      23936: inst = 32'hc4044da;
      23937: inst = 32'h8220000;
      23938: inst = 32'h10408000;
      23939: inst = 32'hc4044db;
      23940: inst = 32'h8220000;
      23941: inst = 32'h10408000;
      23942: inst = 32'hc4044dc;
      23943: inst = 32'h8220000;
      23944: inst = 32'h10408000;
      23945: inst = 32'hc4044dd;
      23946: inst = 32'h8220000;
      23947: inst = 32'h10408000;
      23948: inst = 32'hc4044de;
      23949: inst = 32'h8220000;
      23950: inst = 32'h10408000;
      23951: inst = 32'hc4044df;
      23952: inst = 32'h8220000;
      23953: inst = 32'h10408000;
      23954: inst = 32'hc4044e0;
      23955: inst = 32'h8220000;
      23956: inst = 32'h10408000;
      23957: inst = 32'hc4044e1;
      23958: inst = 32'h8220000;
      23959: inst = 32'h10408000;
      23960: inst = 32'hc4044e2;
      23961: inst = 32'h8220000;
      23962: inst = 32'h10408000;
      23963: inst = 32'hc4044e3;
      23964: inst = 32'h8220000;
      23965: inst = 32'h10408000;
      23966: inst = 32'hc4044e4;
      23967: inst = 32'h8220000;
      23968: inst = 32'h10408000;
      23969: inst = 32'hc4044e5;
      23970: inst = 32'h8220000;
      23971: inst = 32'h10408000;
      23972: inst = 32'hc4044e6;
      23973: inst = 32'h8220000;
      23974: inst = 32'h10408000;
      23975: inst = 32'hc4044e7;
      23976: inst = 32'h8220000;
      23977: inst = 32'h10408000;
      23978: inst = 32'hc4044e8;
      23979: inst = 32'h8220000;
      23980: inst = 32'h10408000;
      23981: inst = 32'hc4044e9;
      23982: inst = 32'h8220000;
      23983: inst = 32'h10408000;
      23984: inst = 32'hc4044ea;
      23985: inst = 32'h8220000;
      23986: inst = 32'h10408000;
      23987: inst = 32'hc4044eb;
      23988: inst = 32'h8220000;
      23989: inst = 32'h10408000;
      23990: inst = 32'hc4044ec;
      23991: inst = 32'h8220000;
      23992: inst = 32'h10408000;
      23993: inst = 32'hc4044ed;
      23994: inst = 32'h8220000;
      23995: inst = 32'h10408000;
      23996: inst = 32'hc4044ee;
      23997: inst = 32'h8220000;
      23998: inst = 32'h10408000;
      23999: inst = 32'hc4044ef;
      24000: inst = 32'h8220000;
      24001: inst = 32'h10408000;
      24002: inst = 32'hc4044f0;
      24003: inst = 32'h8220000;
      24004: inst = 32'h10408000;
      24005: inst = 32'hc4044f1;
      24006: inst = 32'h8220000;
      24007: inst = 32'h10408000;
      24008: inst = 32'hc4044f2;
      24009: inst = 32'h8220000;
      24010: inst = 32'h10408000;
      24011: inst = 32'hc4044f3;
      24012: inst = 32'h8220000;
      24013: inst = 32'h10408000;
      24014: inst = 32'hc4044f4;
      24015: inst = 32'h8220000;
      24016: inst = 32'h10408000;
      24017: inst = 32'hc4044f5;
      24018: inst = 32'h8220000;
      24019: inst = 32'h10408000;
      24020: inst = 32'hc4044f6;
      24021: inst = 32'h8220000;
      24022: inst = 32'h10408000;
      24023: inst = 32'hc4044f7;
      24024: inst = 32'h8220000;
      24025: inst = 32'h10408000;
      24026: inst = 32'hc4044f8;
      24027: inst = 32'h8220000;
      24028: inst = 32'h10408000;
      24029: inst = 32'hc4044f9;
      24030: inst = 32'h8220000;
      24031: inst = 32'h10408000;
      24032: inst = 32'hc4044fa;
      24033: inst = 32'h8220000;
      24034: inst = 32'h10408000;
      24035: inst = 32'hc4044fb;
      24036: inst = 32'h8220000;
      24037: inst = 32'h10408000;
      24038: inst = 32'hc4044fc;
      24039: inst = 32'h8220000;
      24040: inst = 32'h10408000;
      24041: inst = 32'hc4044fd;
      24042: inst = 32'h8220000;
      24043: inst = 32'h10408000;
      24044: inst = 32'hc4044fe;
      24045: inst = 32'h8220000;
      24046: inst = 32'h10408000;
      24047: inst = 32'hc4044ff;
      24048: inst = 32'h8220000;
      24049: inst = 32'h10408000;
      24050: inst = 32'hc404500;
      24051: inst = 32'h8220000;
      24052: inst = 32'h10408000;
      24053: inst = 32'hc404501;
      24054: inst = 32'h8220000;
      24055: inst = 32'h10408000;
      24056: inst = 32'hc404502;
      24057: inst = 32'h8220000;
      24058: inst = 32'h10408000;
      24059: inst = 32'hc404503;
      24060: inst = 32'h8220000;
      24061: inst = 32'h10408000;
      24062: inst = 32'hc404504;
      24063: inst = 32'h8220000;
      24064: inst = 32'h10408000;
      24065: inst = 32'hc404505;
      24066: inst = 32'h8220000;
      24067: inst = 32'h10408000;
      24068: inst = 32'hc404506;
      24069: inst = 32'h8220000;
      24070: inst = 32'h10408000;
      24071: inst = 32'hc404507;
      24072: inst = 32'h8220000;
      24073: inst = 32'h10408000;
      24074: inst = 32'hc404508;
      24075: inst = 32'h8220000;
      24076: inst = 32'h10408000;
      24077: inst = 32'hc404509;
      24078: inst = 32'h8220000;
      24079: inst = 32'h10408000;
      24080: inst = 32'hc40450a;
      24081: inst = 32'h8220000;
      24082: inst = 32'h10408000;
      24083: inst = 32'hc40450b;
      24084: inst = 32'h8220000;
      24085: inst = 32'h10408000;
      24086: inst = 32'hc40450c;
      24087: inst = 32'h8220000;
      24088: inst = 32'h10408000;
      24089: inst = 32'hc40450d;
      24090: inst = 32'h8220000;
      24091: inst = 32'h10408000;
      24092: inst = 32'hc40450e;
      24093: inst = 32'h8220000;
      24094: inst = 32'h10408000;
      24095: inst = 32'hc40450f;
      24096: inst = 32'h8220000;
      24097: inst = 32'h10408000;
      24098: inst = 32'hc404510;
      24099: inst = 32'h8220000;
      24100: inst = 32'h10408000;
      24101: inst = 32'hc404511;
      24102: inst = 32'h8220000;
      24103: inst = 32'h10408000;
      24104: inst = 32'hc404512;
      24105: inst = 32'h8220000;
      24106: inst = 32'h10408000;
      24107: inst = 32'hc404513;
      24108: inst = 32'h8220000;
      24109: inst = 32'h10408000;
      24110: inst = 32'hc404514;
      24111: inst = 32'h8220000;
      24112: inst = 32'h10408000;
      24113: inst = 32'hc404515;
      24114: inst = 32'h8220000;
      24115: inst = 32'h10408000;
      24116: inst = 32'hc404516;
      24117: inst = 32'h8220000;
      24118: inst = 32'h10408000;
      24119: inst = 32'hc404517;
      24120: inst = 32'h8220000;
      24121: inst = 32'h10408000;
      24122: inst = 32'hc404518;
      24123: inst = 32'h8220000;
      24124: inst = 32'h10408000;
      24125: inst = 32'hc404527;
      24126: inst = 32'h8220000;
      24127: inst = 32'h10408000;
      24128: inst = 32'hc404528;
      24129: inst = 32'h8220000;
      24130: inst = 32'h10408000;
      24131: inst = 32'hc404529;
      24132: inst = 32'h8220000;
      24133: inst = 32'h10408000;
      24134: inst = 32'hc40452a;
      24135: inst = 32'h8220000;
      24136: inst = 32'h10408000;
      24137: inst = 32'hc40452b;
      24138: inst = 32'h8220000;
      24139: inst = 32'h10408000;
      24140: inst = 32'hc40452c;
      24141: inst = 32'h8220000;
      24142: inst = 32'h10408000;
      24143: inst = 32'hc40452d;
      24144: inst = 32'h8220000;
      24145: inst = 32'h10408000;
      24146: inst = 32'hc40452e;
      24147: inst = 32'h8220000;
      24148: inst = 32'h10408000;
      24149: inst = 32'hc40452f;
      24150: inst = 32'h8220000;
      24151: inst = 32'h10408000;
      24152: inst = 32'hc404530;
      24153: inst = 32'h8220000;
      24154: inst = 32'h10408000;
      24155: inst = 32'hc404531;
      24156: inst = 32'h8220000;
      24157: inst = 32'h10408000;
      24158: inst = 32'hc404532;
      24159: inst = 32'h8220000;
      24160: inst = 32'h10408000;
      24161: inst = 32'hc404533;
      24162: inst = 32'h8220000;
      24163: inst = 32'h10408000;
      24164: inst = 32'hc404534;
      24165: inst = 32'h8220000;
      24166: inst = 32'h10408000;
      24167: inst = 32'hc404535;
      24168: inst = 32'h8220000;
      24169: inst = 32'h10408000;
      24170: inst = 32'hc404536;
      24171: inst = 32'h8220000;
      24172: inst = 32'h10408000;
      24173: inst = 32'hc404537;
      24174: inst = 32'h8220000;
      24175: inst = 32'h10408000;
      24176: inst = 32'hc404538;
      24177: inst = 32'h8220000;
      24178: inst = 32'h10408000;
      24179: inst = 32'hc404539;
      24180: inst = 32'h8220000;
      24181: inst = 32'h10408000;
      24182: inst = 32'hc40453a;
      24183: inst = 32'h8220000;
      24184: inst = 32'h10408000;
      24185: inst = 32'hc40453b;
      24186: inst = 32'h8220000;
      24187: inst = 32'h10408000;
      24188: inst = 32'hc40453c;
      24189: inst = 32'h8220000;
      24190: inst = 32'h10408000;
      24191: inst = 32'hc40453d;
      24192: inst = 32'h8220000;
      24193: inst = 32'h10408000;
      24194: inst = 32'hc40453e;
      24195: inst = 32'h8220000;
      24196: inst = 32'h10408000;
      24197: inst = 32'hc40453f;
      24198: inst = 32'h8220000;
      24199: inst = 32'h10408000;
      24200: inst = 32'hc404540;
      24201: inst = 32'h8220000;
      24202: inst = 32'h10408000;
      24203: inst = 32'hc404541;
      24204: inst = 32'h8220000;
      24205: inst = 32'h10408000;
      24206: inst = 32'hc404542;
      24207: inst = 32'h8220000;
      24208: inst = 32'h10408000;
      24209: inst = 32'hc404543;
      24210: inst = 32'h8220000;
      24211: inst = 32'h10408000;
      24212: inst = 32'hc404544;
      24213: inst = 32'h8220000;
      24214: inst = 32'h10408000;
      24215: inst = 32'hc404545;
      24216: inst = 32'h8220000;
      24217: inst = 32'h10408000;
      24218: inst = 32'hc404546;
      24219: inst = 32'h8220000;
      24220: inst = 32'h10408000;
      24221: inst = 32'hc404547;
      24222: inst = 32'h8220000;
      24223: inst = 32'h10408000;
      24224: inst = 32'hc404548;
      24225: inst = 32'h8220000;
      24226: inst = 32'h10408000;
      24227: inst = 32'hc404549;
      24228: inst = 32'h8220000;
      24229: inst = 32'h10408000;
      24230: inst = 32'hc40454a;
      24231: inst = 32'h8220000;
      24232: inst = 32'h10408000;
      24233: inst = 32'hc40454b;
      24234: inst = 32'h8220000;
      24235: inst = 32'h10408000;
      24236: inst = 32'hc40454c;
      24237: inst = 32'h8220000;
      24238: inst = 32'h10408000;
      24239: inst = 32'hc40454d;
      24240: inst = 32'h8220000;
      24241: inst = 32'h10408000;
      24242: inst = 32'hc40454e;
      24243: inst = 32'h8220000;
      24244: inst = 32'h10408000;
      24245: inst = 32'hc40454f;
      24246: inst = 32'h8220000;
      24247: inst = 32'h10408000;
      24248: inst = 32'hc404550;
      24249: inst = 32'h8220000;
      24250: inst = 32'h10408000;
      24251: inst = 32'hc404551;
      24252: inst = 32'h8220000;
      24253: inst = 32'h10408000;
      24254: inst = 32'hc404552;
      24255: inst = 32'h8220000;
      24256: inst = 32'h10408000;
      24257: inst = 32'hc404553;
      24258: inst = 32'h8220000;
      24259: inst = 32'h10408000;
      24260: inst = 32'hc404554;
      24261: inst = 32'h8220000;
      24262: inst = 32'h10408000;
      24263: inst = 32'hc404555;
      24264: inst = 32'h8220000;
      24265: inst = 32'h10408000;
      24266: inst = 32'hc404556;
      24267: inst = 32'h8220000;
      24268: inst = 32'h10408000;
      24269: inst = 32'hc404557;
      24270: inst = 32'h8220000;
      24271: inst = 32'h10408000;
      24272: inst = 32'hc404558;
      24273: inst = 32'h8220000;
      24274: inst = 32'h10408000;
      24275: inst = 32'hc404559;
      24276: inst = 32'h8220000;
      24277: inst = 32'h10408000;
      24278: inst = 32'hc40455a;
      24279: inst = 32'h8220000;
      24280: inst = 32'h10408000;
      24281: inst = 32'hc40455b;
      24282: inst = 32'h8220000;
      24283: inst = 32'h10408000;
      24284: inst = 32'hc40455c;
      24285: inst = 32'h8220000;
      24286: inst = 32'h10408000;
      24287: inst = 32'hc40455d;
      24288: inst = 32'h8220000;
      24289: inst = 32'h10408000;
      24290: inst = 32'hc40455e;
      24291: inst = 32'h8220000;
      24292: inst = 32'h10408000;
      24293: inst = 32'hc40455f;
      24294: inst = 32'h8220000;
      24295: inst = 32'h10408000;
      24296: inst = 32'hc404560;
      24297: inst = 32'h8220000;
      24298: inst = 32'h10408000;
      24299: inst = 32'hc404561;
      24300: inst = 32'h8220000;
      24301: inst = 32'h10408000;
      24302: inst = 32'hc404562;
      24303: inst = 32'h8220000;
      24304: inst = 32'h10408000;
      24305: inst = 32'hc404563;
      24306: inst = 32'h8220000;
      24307: inst = 32'h10408000;
      24308: inst = 32'hc404564;
      24309: inst = 32'h8220000;
      24310: inst = 32'h10408000;
      24311: inst = 32'hc404565;
      24312: inst = 32'h8220000;
      24313: inst = 32'h10408000;
      24314: inst = 32'hc404566;
      24315: inst = 32'h8220000;
      24316: inst = 32'h10408000;
      24317: inst = 32'hc404567;
      24318: inst = 32'h8220000;
      24319: inst = 32'h10408000;
      24320: inst = 32'hc404568;
      24321: inst = 32'h8220000;
      24322: inst = 32'h10408000;
      24323: inst = 32'hc404569;
      24324: inst = 32'h8220000;
      24325: inst = 32'h10408000;
      24326: inst = 32'hc40456a;
      24327: inst = 32'h8220000;
      24328: inst = 32'h10408000;
      24329: inst = 32'hc40456b;
      24330: inst = 32'h8220000;
      24331: inst = 32'h10408000;
      24332: inst = 32'hc40456c;
      24333: inst = 32'h8220000;
      24334: inst = 32'h10408000;
      24335: inst = 32'hc40456d;
      24336: inst = 32'h8220000;
      24337: inst = 32'h10408000;
      24338: inst = 32'hc40456e;
      24339: inst = 32'h8220000;
      24340: inst = 32'h10408000;
      24341: inst = 32'hc40456f;
      24342: inst = 32'h8220000;
      24343: inst = 32'h10408000;
      24344: inst = 32'hc404570;
      24345: inst = 32'h8220000;
      24346: inst = 32'h10408000;
      24347: inst = 32'hc404571;
      24348: inst = 32'h8220000;
      24349: inst = 32'h10408000;
      24350: inst = 32'hc404572;
      24351: inst = 32'h8220000;
      24352: inst = 32'h10408000;
      24353: inst = 32'hc404573;
      24354: inst = 32'h8220000;
      24355: inst = 32'h10408000;
      24356: inst = 32'hc404574;
      24357: inst = 32'h8220000;
      24358: inst = 32'h10408000;
      24359: inst = 32'hc404575;
      24360: inst = 32'h8220000;
      24361: inst = 32'h10408000;
      24362: inst = 32'hc404576;
      24363: inst = 32'h8220000;
      24364: inst = 32'h10408000;
      24365: inst = 32'hc404577;
      24366: inst = 32'h8220000;
      24367: inst = 32'h10408000;
      24368: inst = 32'hc404578;
      24369: inst = 32'h8220000;
      24370: inst = 32'h10408000;
      24371: inst = 32'hc404587;
      24372: inst = 32'h8220000;
      24373: inst = 32'h10408000;
      24374: inst = 32'hc404588;
      24375: inst = 32'h8220000;
      24376: inst = 32'h10408000;
      24377: inst = 32'hc404589;
      24378: inst = 32'h8220000;
      24379: inst = 32'h10408000;
      24380: inst = 32'hc40458a;
      24381: inst = 32'h8220000;
      24382: inst = 32'h10408000;
      24383: inst = 32'hc40458b;
      24384: inst = 32'h8220000;
      24385: inst = 32'h10408000;
      24386: inst = 32'hc40458c;
      24387: inst = 32'h8220000;
      24388: inst = 32'h10408000;
      24389: inst = 32'hc40458d;
      24390: inst = 32'h8220000;
      24391: inst = 32'h10408000;
      24392: inst = 32'hc40458e;
      24393: inst = 32'h8220000;
      24394: inst = 32'h10408000;
      24395: inst = 32'hc40458f;
      24396: inst = 32'h8220000;
      24397: inst = 32'h10408000;
      24398: inst = 32'hc404590;
      24399: inst = 32'h8220000;
      24400: inst = 32'h10408000;
      24401: inst = 32'hc404591;
      24402: inst = 32'h8220000;
      24403: inst = 32'h10408000;
      24404: inst = 32'hc404592;
      24405: inst = 32'h8220000;
      24406: inst = 32'h10408000;
      24407: inst = 32'hc404593;
      24408: inst = 32'h8220000;
      24409: inst = 32'h10408000;
      24410: inst = 32'hc404594;
      24411: inst = 32'h8220000;
      24412: inst = 32'h10408000;
      24413: inst = 32'hc404595;
      24414: inst = 32'h8220000;
      24415: inst = 32'h10408000;
      24416: inst = 32'hc404596;
      24417: inst = 32'h8220000;
      24418: inst = 32'h10408000;
      24419: inst = 32'hc404597;
      24420: inst = 32'h8220000;
      24421: inst = 32'h10408000;
      24422: inst = 32'hc404598;
      24423: inst = 32'h8220000;
      24424: inst = 32'h10408000;
      24425: inst = 32'hc404599;
      24426: inst = 32'h8220000;
      24427: inst = 32'h10408000;
      24428: inst = 32'hc40459a;
      24429: inst = 32'h8220000;
      24430: inst = 32'h10408000;
      24431: inst = 32'hc40459b;
      24432: inst = 32'h8220000;
      24433: inst = 32'h10408000;
      24434: inst = 32'hc40459c;
      24435: inst = 32'h8220000;
      24436: inst = 32'h10408000;
      24437: inst = 32'hc40459d;
      24438: inst = 32'h8220000;
      24439: inst = 32'h10408000;
      24440: inst = 32'hc40459e;
      24441: inst = 32'h8220000;
      24442: inst = 32'h10408000;
      24443: inst = 32'hc40459f;
      24444: inst = 32'h8220000;
      24445: inst = 32'h10408000;
      24446: inst = 32'hc4045a0;
      24447: inst = 32'h8220000;
      24448: inst = 32'h10408000;
      24449: inst = 32'hc4045a1;
      24450: inst = 32'h8220000;
      24451: inst = 32'h10408000;
      24452: inst = 32'hc4045a2;
      24453: inst = 32'h8220000;
      24454: inst = 32'h10408000;
      24455: inst = 32'hc4045a3;
      24456: inst = 32'h8220000;
      24457: inst = 32'h10408000;
      24458: inst = 32'hc4045a4;
      24459: inst = 32'h8220000;
      24460: inst = 32'h10408000;
      24461: inst = 32'hc4045a5;
      24462: inst = 32'h8220000;
      24463: inst = 32'h10408000;
      24464: inst = 32'hc4045a6;
      24465: inst = 32'h8220000;
      24466: inst = 32'h10408000;
      24467: inst = 32'hc4045a7;
      24468: inst = 32'h8220000;
      24469: inst = 32'h10408000;
      24470: inst = 32'hc4045a8;
      24471: inst = 32'h8220000;
      24472: inst = 32'h10408000;
      24473: inst = 32'hc4045a9;
      24474: inst = 32'h8220000;
      24475: inst = 32'h10408000;
      24476: inst = 32'hc4045aa;
      24477: inst = 32'h8220000;
      24478: inst = 32'h10408000;
      24479: inst = 32'hc4045ab;
      24480: inst = 32'h8220000;
      24481: inst = 32'h10408000;
      24482: inst = 32'hc4045ac;
      24483: inst = 32'h8220000;
      24484: inst = 32'h10408000;
      24485: inst = 32'hc4045ad;
      24486: inst = 32'h8220000;
      24487: inst = 32'h10408000;
      24488: inst = 32'hc4045ae;
      24489: inst = 32'h8220000;
      24490: inst = 32'h10408000;
      24491: inst = 32'hc4045af;
      24492: inst = 32'h8220000;
      24493: inst = 32'h10408000;
      24494: inst = 32'hc4045b0;
      24495: inst = 32'h8220000;
      24496: inst = 32'h10408000;
      24497: inst = 32'hc4045b1;
      24498: inst = 32'h8220000;
      24499: inst = 32'h10408000;
      24500: inst = 32'hc4045b2;
      24501: inst = 32'h8220000;
      24502: inst = 32'h10408000;
      24503: inst = 32'hc4045b3;
      24504: inst = 32'h8220000;
      24505: inst = 32'h10408000;
      24506: inst = 32'hc4045b4;
      24507: inst = 32'h8220000;
      24508: inst = 32'h10408000;
      24509: inst = 32'hc4045b5;
      24510: inst = 32'h8220000;
      24511: inst = 32'h10408000;
      24512: inst = 32'hc4045b6;
      24513: inst = 32'h8220000;
      24514: inst = 32'h10408000;
      24515: inst = 32'hc4045b7;
      24516: inst = 32'h8220000;
      24517: inst = 32'h10408000;
      24518: inst = 32'hc4045b8;
      24519: inst = 32'h8220000;
      24520: inst = 32'h10408000;
      24521: inst = 32'hc4045b9;
      24522: inst = 32'h8220000;
      24523: inst = 32'h10408000;
      24524: inst = 32'hc4045ba;
      24525: inst = 32'h8220000;
      24526: inst = 32'h10408000;
      24527: inst = 32'hc4045bb;
      24528: inst = 32'h8220000;
      24529: inst = 32'h10408000;
      24530: inst = 32'hc4045bc;
      24531: inst = 32'h8220000;
      24532: inst = 32'h10408000;
      24533: inst = 32'hc4045bd;
      24534: inst = 32'h8220000;
      24535: inst = 32'h10408000;
      24536: inst = 32'hc4045be;
      24537: inst = 32'h8220000;
      24538: inst = 32'h10408000;
      24539: inst = 32'hc4045bf;
      24540: inst = 32'h8220000;
      24541: inst = 32'h10408000;
      24542: inst = 32'hc4045c0;
      24543: inst = 32'h8220000;
      24544: inst = 32'h10408000;
      24545: inst = 32'hc4045c1;
      24546: inst = 32'h8220000;
      24547: inst = 32'h10408000;
      24548: inst = 32'hc4045c2;
      24549: inst = 32'h8220000;
      24550: inst = 32'h10408000;
      24551: inst = 32'hc4045c3;
      24552: inst = 32'h8220000;
      24553: inst = 32'h10408000;
      24554: inst = 32'hc4045c4;
      24555: inst = 32'h8220000;
      24556: inst = 32'h10408000;
      24557: inst = 32'hc4045c5;
      24558: inst = 32'h8220000;
      24559: inst = 32'h10408000;
      24560: inst = 32'hc4045c6;
      24561: inst = 32'h8220000;
      24562: inst = 32'h10408000;
      24563: inst = 32'hc4045c7;
      24564: inst = 32'h8220000;
      24565: inst = 32'h10408000;
      24566: inst = 32'hc4045c8;
      24567: inst = 32'h8220000;
      24568: inst = 32'h10408000;
      24569: inst = 32'hc4045c9;
      24570: inst = 32'h8220000;
      24571: inst = 32'h10408000;
      24572: inst = 32'hc4045ca;
      24573: inst = 32'h8220000;
      24574: inst = 32'h10408000;
      24575: inst = 32'hc4045cb;
      24576: inst = 32'h8220000;
      24577: inst = 32'h10408000;
      24578: inst = 32'hc4045cc;
      24579: inst = 32'h8220000;
      24580: inst = 32'h10408000;
      24581: inst = 32'hc4045cd;
      24582: inst = 32'h8220000;
      24583: inst = 32'h10408000;
      24584: inst = 32'hc4045ce;
      24585: inst = 32'h8220000;
      24586: inst = 32'h10408000;
      24587: inst = 32'hc4045cf;
      24588: inst = 32'h8220000;
      24589: inst = 32'h10408000;
      24590: inst = 32'hc4045d0;
      24591: inst = 32'h8220000;
      24592: inst = 32'h10408000;
      24593: inst = 32'hc4045d1;
      24594: inst = 32'h8220000;
      24595: inst = 32'h10408000;
      24596: inst = 32'hc4045d2;
      24597: inst = 32'h8220000;
      24598: inst = 32'h10408000;
      24599: inst = 32'hc4045d3;
      24600: inst = 32'h8220000;
      24601: inst = 32'h10408000;
      24602: inst = 32'hc4045d4;
      24603: inst = 32'h8220000;
      24604: inst = 32'h10408000;
      24605: inst = 32'hc4045d5;
      24606: inst = 32'h8220000;
      24607: inst = 32'h10408000;
      24608: inst = 32'hc4045d6;
      24609: inst = 32'h8220000;
      24610: inst = 32'h10408000;
      24611: inst = 32'hc4045d7;
      24612: inst = 32'h8220000;
      24613: inst = 32'h10408000;
      24614: inst = 32'hc4045d8;
      24615: inst = 32'h8220000;
      24616: inst = 32'h10408000;
      24617: inst = 32'hc4045e7;
      24618: inst = 32'h8220000;
      24619: inst = 32'h10408000;
      24620: inst = 32'hc4045e8;
      24621: inst = 32'h8220000;
      24622: inst = 32'h10408000;
      24623: inst = 32'hc4045e9;
      24624: inst = 32'h8220000;
      24625: inst = 32'h10408000;
      24626: inst = 32'hc4045ea;
      24627: inst = 32'h8220000;
      24628: inst = 32'h10408000;
      24629: inst = 32'hc4045eb;
      24630: inst = 32'h8220000;
      24631: inst = 32'h10408000;
      24632: inst = 32'hc4045ec;
      24633: inst = 32'h8220000;
      24634: inst = 32'h10408000;
      24635: inst = 32'hc4045ed;
      24636: inst = 32'h8220000;
      24637: inst = 32'h10408000;
      24638: inst = 32'hc4045ee;
      24639: inst = 32'h8220000;
      24640: inst = 32'h10408000;
      24641: inst = 32'hc4045ef;
      24642: inst = 32'h8220000;
      24643: inst = 32'h10408000;
      24644: inst = 32'hc4045f0;
      24645: inst = 32'h8220000;
      24646: inst = 32'h10408000;
      24647: inst = 32'hc4045f1;
      24648: inst = 32'h8220000;
      24649: inst = 32'h10408000;
      24650: inst = 32'hc4045f2;
      24651: inst = 32'h8220000;
      24652: inst = 32'h10408000;
      24653: inst = 32'hc4045f3;
      24654: inst = 32'h8220000;
      24655: inst = 32'h10408000;
      24656: inst = 32'hc4045f4;
      24657: inst = 32'h8220000;
      24658: inst = 32'h10408000;
      24659: inst = 32'hc4045f5;
      24660: inst = 32'h8220000;
      24661: inst = 32'h10408000;
      24662: inst = 32'hc4045f6;
      24663: inst = 32'h8220000;
      24664: inst = 32'h10408000;
      24665: inst = 32'hc4045f7;
      24666: inst = 32'h8220000;
      24667: inst = 32'h10408000;
      24668: inst = 32'hc4045f8;
      24669: inst = 32'h8220000;
      24670: inst = 32'h10408000;
      24671: inst = 32'hc4045f9;
      24672: inst = 32'h8220000;
      24673: inst = 32'h10408000;
      24674: inst = 32'hc4045fa;
      24675: inst = 32'h8220000;
      24676: inst = 32'h10408000;
      24677: inst = 32'hc4045fb;
      24678: inst = 32'h8220000;
      24679: inst = 32'h10408000;
      24680: inst = 32'hc4045fc;
      24681: inst = 32'h8220000;
      24682: inst = 32'h10408000;
      24683: inst = 32'hc4045fd;
      24684: inst = 32'h8220000;
      24685: inst = 32'h10408000;
      24686: inst = 32'hc4045fe;
      24687: inst = 32'h8220000;
      24688: inst = 32'h10408000;
      24689: inst = 32'hc4045ff;
      24690: inst = 32'h8220000;
      24691: inst = 32'h10408000;
      24692: inst = 32'hc404600;
      24693: inst = 32'h8220000;
      24694: inst = 32'h10408000;
      24695: inst = 32'hc404601;
      24696: inst = 32'h8220000;
      24697: inst = 32'h10408000;
      24698: inst = 32'hc404602;
      24699: inst = 32'h8220000;
      24700: inst = 32'h10408000;
      24701: inst = 32'hc404603;
      24702: inst = 32'h8220000;
      24703: inst = 32'h10408000;
      24704: inst = 32'hc404604;
      24705: inst = 32'h8220000;
      24706: inst = 32'h10408000;
      24707: inst = 32'hc404605;
      24708: inst = 32'h8220000;
      24709: inst = 32'h10408000;
      24710: inst = 32'hc404606;
      24711: inst = 32'h8220000;
      24712: inst = 32'h10408000;
      24713: inst = 32'hc404607;
      24714: inst = 32'h8220000;
      24715: inst = 32'h10408000;
      24716: inst = 32'hc404608;
      24717: inst = 32'h8220000;
      24718: inst = 32'h10408000;
      24719: inst = 32'hc404609;
      24720: inst = 32'h8220000;
      24721: inst = 32'h10408000;
      24722: inst = 32'hc40460a;
      24723: inst = 32'h8220000;
      24724: inst = 32'h10408000;
      24725: inst = 32'hc40460b;
      24726: inst = 32'h8220000;
      24727: inst = 32'h10408000;
      24728: inst = 32'hc40460c;
      24729: inst = 32'h8220000;
      24730: inst = 32'h10408000;
      24731: inst = 32'hc40460d;
      24732: inst = 32'h8220000;
      24733: inst = 32'h10408000;
      24734: inst = 32'hc40460e;
      24735: inst = 32'h8220000;
      24736: inst = 32'h10408000;
      24737: inst = 32'hc40460f;
      24738: inst = 32'h8220000;
      24739: inst = 32'h10408000;
      24740: inst = 32'hc404610;
      24741: inst = 32'h8220000;
      24742: inst = 32'h10408000;
      24743: inst = 32'hc404611;
      24744: inst = 32'h8220000;
      24745: inst = 32'h10408000;
      24746: inst = 32'hc404612;
      24747: inst = 32'h8220000;
      24748: inst = 32'h10408000;
      24749: inst = 32'hc404613;
      24750: inst = 32'h8220000;
      24751: inst = 32'h10408000;
      24752: inst = 32'hc404614;
      24753: inst = 32'h8220000;
      24754: inst = 32'h10408000;
      24755: inst = 32'hc404615;
      24756: inst = 32'h8220000;
      24757: inst = 32'h10408000;
      24758: inst = 32'hc404616;
      24759: inst = 32'h8220000;
      24760: inst = 32'h10408000;
      24761: inst = 32'hc404617;
      24762: inst = 32'h8220000;
      24763: inst = 32'h10408000;
      24764: inst = 32'hc404618;
      24765: inst = 32'h8220000;
      24766: inst = 32'h10408000;
      24767: inst = 32'hc404619;
      24768: inst = 32'h8220000;
      24769: inst = 32'h10408000;
      24770: inst = 32'hc40461a;
      24771: inst = 32'h8220000;
      24772: inst = 32'h10408000;
      24773: inst = 32'hc40461b;
      24774: inst = 32'h8220000;
      24775: inst = 32'h10408000;
      24776: inst = 32'hc40461c;
      24777: inst = 32'h8220000;
      24778: inst = 32'h10408000;
      24779: inst = 32'hc40461d;
      24780: inst = 32'h8220000;
      24781: inst = 32'h10408000;
      24782: inst = 32'hc40461e;
      24783: inst = 32'h8220000;
      24784: inst = 32'h10408000;
      24785: inst = 32'hc40461f;
      24786: inst = 32'h8220000;
      24787: inst = 32'h10408000;
      24788: inst = 32'hc404620;
      24789: inst = 32'h8220000;
      24790: inst = 32'h10408000;
      24791: inst = 32'hc404621;
      24792: inst = 32'h8220000;
      24793: inst = 32'h10408000;
      24794: inst = 32'hc404622;
      24795: inst = 32'h8220000;
      24796: inst = 32'h10408000;
      24797: inst = 32'hc404623;
      24798: inst = 32'h8220000;
      24799: inst = 32'h10408000;
      24800: inst = 32'hc404624;
      24801: inst = 32'h8220000;
      24802: inst = 32'h10408000;
      24803: inst = 32'hc404625;
      24804: inst = 32'h8220000;
      24805: inst = 32'h10408000;
      24806: inst = 32'hc404626;
      24807: inst = 32'h8220000;
      24808: inst = 32'h10408000;
      24809: inst = 32'hc404627;
      24810: inst = 32'h8220000;
      24811: inst = 32'h10408000;
      24812: inst = 32'hc404628;
      24813: inst = 32'h8220000;
      24814: inst = 32'h10408000;
      24815: inst = 32'hc404629;
      24816: inst = 32'h8220000;
      24817: inst = 32'h10408000;
      24818: inst = 32'hc40462a;
      24819: inst = 32'h8220000;
      24820: inst = 32'h10408000;
      24821: inst = 32'hc40462b;
      24822: inst = 32'h8220000;
      24823: inst = 32'h10408000;
      24824: inst = 32'hc40462c;
      24825: inst = 32'h8220000;
      24826: inst = 32'h10408000;
      24827: inst = 32'hc40462d;
      24828: inst = 32'h8220000;
      24829: inst = 32'h10408000;
      24830: inst = 32'hc40462e;
      24831: inst = 32'h8220000;
      24832: inst = 32'h10408000;
      24833: inst = 32'hc40462f;
      24834: inst = 32'h8220000;
      24835: inst = 32'h10408000;
      24836: inst = 32'hc404630;
      24837: inst = 32'h8220000;
      24838: inst = 32'h10408000;
      24839: inst = 32'hc404631;
      24840: inst = 32'h8220000;
      24841: inst = 32'h10408000;
      24842: inst = 32'hc404632;
      24843: inst = 32'h8220000;
      24844: inst = 32'h10408000;
      24845: inst = 32'hc404633;
      24846: inst = 32'h8220000;
      24847: inst = 32'h10408000;
      24848: inst = 32'hc404634;
      24849: inst = 32'h8220000;
      24850: inst = 32'h10408000;
      24851: inst = 32'hc404635;
      24852: inst = 32'h8220000;
      24853: inst = 32'h10408000;
      24854: inst = 32'hc404636;
      24855: inst = 32'h8220000;
      24856: inst = 32'h10408000;
      24857: inst = 32'hc404637;
      24858: inst = 32'h8220000;
      24859: inst = 32'h10408000;
      24860: inst = 32'hc404638;
      24861: inst = 32'h8220000;
      24862: inst = 32'h10408000;
      24863: inst = 32'hc404647;
      24864: inst = 32'h8220000;
      24865: inst = 32'h10408000;
      24866: inst = 32'hc404648;
      24867: inst = 32'h8220000;
      24868: inst = 32'h10408000;
      24869: inst = 32'hc404649;
      24870: inst = 32'h8220000;
      24871: inst = 32'h10408000;
      24872: inst = 32'hc40464a;
      24873: inst = 32'h8220000;
      24874: inst = 32'h10408000;
      24875: inst = 32'hc40464b;
      24876: inst = 32'h8220000;
      24877: inst = 32'h10408000;
      24878: inst = 32'hc40464c;
      24879: inst = 32'h8220000;
      24880: inst = 32'h10408000;
      24881: inst = 32'hc40464d;
      24882: inst = 32'h8220000;
      24883: inst = 32'h10408000;
      24884: inst = 32'hc404651;
      24885: inst = 32'h8220000;
      24886: inst = 32'h10408000;
      24887: inst = 32'hc404652;
      24888: inst = 32'h8220000;
      24889: inst = 32'h10408000;
      24890: inst = 32'hc404653;
      24891: inst = 32'h8220000;
      24892: inst = 32'h10408000;
      24893: inst = 32'hc404654;
      24894: inst = 32'h8220000;
      24895: inst = 32'h10408000;
      24896: inst = 32'hc404655;
      24897: inst = 32'h8220000;
      24898: inst = 32'h10408000;
      24899: inst = 32'hc404656;
      24900: inst = 32'h8220000;
      24901: inst = 32'h10408000;
      24902: inst = 32'hc404657;
      24903: inst = 32'h8220000;
      24904: inst = 32'h10408000;
      24905: inst = 32'hc404658;
      24906: inst = 32'h8220000;
      24907: inst = 32'h10408000;
      24908: inst = 32'hc404659;
      24909: inst = 32'h8220000;
      24910: inst = 32'h10408000;
      24911: inst = 32'hc40465a;
      24912: inst = 32'h8220000;
      24913: inst = 32'h10408000;
      24914: inst = 32'hc40465b;
      24915: inst = 32'h8220000;
      24916: inst = 32'h10408000;
      24917: inst = 32'hc40465c;
      24918: inst = 32'h8220000;
      24919: inst = 32'h10408000;
      24920: inst = 32'hc40465d;
      24921: inst = 32'h8220000;
      24922: inst = 32'h10408000;
      24923: inst = 32'hc40465e;
      24924: inst = 32'h8220000;
      24925: inst = 32'h10408000;
      24926: inst = 32'hc40465f;
      24927: inst = 32'h8220000;
      24928: inst = 32'h10408000;
      24929: inst = 32'hc404660;
      24930: inst = 32'h8220000;
      24931: inst = 32'h10408000;
      24932: inst = 32'hc404661;
      24933: inst = 32'h8220000;
      24934: inst = 32'h10408000;
      24935: inst = 32'hc404662;
      24936: inst = 32'h8220000;
      24937: inst = 32'h10408000;
      24938: inst = 32'hc404663;
      24939: inst = 32'h8220000;
      24940: inst = 32'h10408000;
      24941: inst = 32'hc404664;
      24942: inst = 32'h8220000;
      24943: inst = 32'h10408000;
      24944: inst = 32'hc404665;
      24945: inst = 32'h8220000;
      24946: inst = 32'h10408000;
      24947: inst = 32'hc404666;
      24948: inst = 32'h8220000;
      24949: inst = 32'h10408000;
      24950: inst = 32'hc404667;
      24951: inst = 32'h8220000;
      24952: inst = 32'h10408000;
      24953: inst = 32'hc404668;
      24954: inst = 32'h8220000;
      24955: inst = 32'h10408000;
      24956: inst = 32'hc404669;
      24957: inst = 32'h8220000;
      24958: inst = 32'h10408000;
      24959: inst = 32'hc40466a;
      24960: inst = 32'h8220000;
      24961: inst = 32'h10408000;
      24962: inst = 32'hc40466b;
      24963: inst = 32'h8220000;
      24964: inst = 32'h10408000;
      24965: inst = 32'hc40466c;
      24966: inst = 32'h8220000;
      24967: inst = 32'h10408000;
      24968: inst = 32'hc40466d;
      24969: inst = 32'h8220000;
      24970: inst = 32'h10408000;
      24971: inst = 32'hc40466e;
      24972: inst = 32'h8220000;
      24973: inst = 32'h10408000;
      24974: inst = 32'hc40466f;
      24975: inst = 32'h8220000;
      24976: inst = 32'h10408000;
      24977: inst = 32'hc404670;
      24978: inst = 32'h8220000;
      24979: inst = 32'h10408000;
      24980: inst = 32'hc404671;
      24981: inst = 32'h8220000;
      24982: inst = 32'h10408000;
      24983: inst = 32'hc404672;
      24984: inst = 32'h8220000;
      24985: inst = 32'h10408000;
      24986: inst = 32'hc404673;
      24987: inst = 32'h8220000;
      24988: inst = 32'h10408000;
      24989: inst = 32'hc404674;
      24990: inst = 32'h8220000;
      24991: inst = 32'h10408000;
      24992: inst = 32'hc404675;
      24993: inst = 32'h8220000;
      24994: inst = 32'h10408000;
      24995: inst = 32'hc404676;
      24996: inst = 32'h8220000;
      24997: inst = 32'h10408000;
      24998: inst = 32'hc404677;
      24999: inst = 32'h8220000;
      25000: inst = 32'h10408000;
      25001: inst = 32'hc404678;
      25002: inst = 32'h8220000;
      25003: inst = 32'h10408000;
      25004: inst = 32'hc404679;
      25005: inst = 32'h8220000;
      25006: inst = 32'h10408000;
      25007: inst = 32'hc40467a;
      25008: inst = 32'h8220000;
      25009: inst = 32'h10408000;
      25010: inst = 32'hc40467b;
      25011: inst = 32'h8220000;
      25012: inst = 32'h10408000;
      25013: inst = 32'hc40467c;
      25014: inst = 32'h8220000;
      25015: inst = 32'h10408000;
      25016: inst = 32'hc40467d;
      25017: inst = 32'h8220000;
      25018: inst = 32'h10408000;
      25019: inst = 32'hc40467e;
      25020: inst = 32'h8220000;
      25021: inst = 32'h10408000;
      25022: inst = 32'hc40467f;
      25023: inst = 32'h8220000;
      25024: inst = 32'h10408000;
      25025: inst = 32'hc404680;
      25026: inst = 32'h8220000;
      25027: inst = 32'h10408000;
      25028: inst = 32'hc404681;
      25029: inst = 32'h8220000;
      25030: inst = 32'h10408000;
      25031: inst = 32'hc404682;
      25032: inst = 32'h8220000;
      25033: inst = 32'h10408000;
      25034: inst = 32'hc404683;
      25035: inst = 32'h8220000;
      25036: inst = 32'h10408000;
      25037: inst = 32'hc404684;
      25038: inst = 32'h8220000;
      25039: inst = 32'h10408000;
      25040: inst = 32'hc404685;
      25041: inst = 32'h8220000;
      25042: inst = 32'h10408000;
      25043: inst = 32'hc404686;
      25044: inst = 32'h8220000;
      25045: inst = 32'h10408000;
      25046: inst = 32'hc404687;
      25047: inst = 32'h8220000;
      25048: inst = 32'h10408000;
      25049: inst = 32'hc404688;
      25050: inst = 32'h8220000;
      25051: inst = 32'h10408000;
      25052: inst = 32'hc404689;
      25053: inst = 32'h8220000;
      25054: inst = 32'h10408000;
      25055: inst = 32'hc40468a;
      25056: inst = 32'h8220000;
      25057: inst = 32'h10408000;
      25058: inst = 32'hc40468b;
      25059: inst = 32'h8220000;
      25060: inst = 32'h10408000;
      25061: inst = 32'hc40468c;
      25062: inst = 32'h8220000;
      25063: inst = 32'h10408000;
      25064: inst = 32'hc40468d;
      25065: inst = 32'h8220000;
      25066: inst = 32'h10408000;
      25067: inst = 32'hc40468e;
      25068: inst = 32'h8220000;
      25069: inst = 32'h10408000;
      25070: inst = 32'hc40468f;
      25071: inst = 32'h8220000;
      25072: inst = 32'h10408000;
      25073: inst = 32'hc404693;
      25074: inst = 32'h8220000;
      25075: inst = 32'h10408000;
      25076: inst = 32'hc404694;
      25077: inst = 32'h8220000;
      25078: inst = 32'h10408000;
      25079: inst = 32'hc404695;
      25080: inst = 32'h8220000;
      25081: inst = 32'h10408000;
      25082: inst = 32'hc404696;
      25083: inst = 32'h8220000;
      25084: inst = 32'h10408000;
      25085: inst = 32'hc404697;
      25086: inst = 32'h8220000;
      25087: inst = 32'h10408000;
      25088: inst = 32'hc404698;
      25089: inst = 32'h8220000;
      25090: inst = 32'h10408000;
      25091: inst = 32'hc4046a7;
      25092: inst = 32'h8220000;
      25093: inst = 32'h10408000;
      25094: inst = 32'hc4046a8;
      25095: inst = 32'h8220000;
      25096: inst = 32'h10408000;
      25097: inst = 32'hc4046a9;
      25098: inst = 32'h8220000;
      25099: inst = 32'h10408000;
      25100: inst = 32'hc4046aa;
      25101: inst = 32'h8220000;
      25102: inst = 32'h10408000;
      25103: inst = 32'hc4046ab;
      25104: inst = 32'h8220000;
      25105: inst = 32'h10408000;
      25106: inst = 32'hc4046ac;
      25107: inst = 32'h8220000;
      25108: inst = 32'h10408000;
      25109: inst = 32'hc4046ad;
      25110: inst = 32'h8220000;
      25111: inst = 32'h10408000;
      25112: inst = 32'hc4046b1;
      25113: inst = 32'h8220000;
      25114: inst = 32'h10408000;
      25115: inst = 32'hc4046b2;
      25116: inst = 32'h8220000;
      25117: inst = 32'h10408000;
      25118: inst = 32'hc4046b3;
      25119: inst = 32'h8220000;
      25120: inst = 32'h10408000;
      25121: inst = 32'hc4046b4;
      25122: inst = 32'h8220000;
      25123: inst = 32'h10408000;
      25124: inst = 32'hc4046b5;
      25125: inst = 32'h8220000;
      25126: inst = 32'h10408000;
      25127: inst = 32'hc4046b6;
      25128: inst = 32'h8220000;
      25129: inst = 32'h10408000;
      25130: inst = 32'hc4046b7;
      25131: inst = 32'h8220000;
      25132: inst = 32'h10408000;
      25133: inst = 32'hc4046b8;
      25134: inst = 32'h8220000;
      25135: inst = 32'h10408000;
      25136: inst = 32'hc4046b9;
      25137: inst = 32'h8220000;
      25138: inst = 32'h10408000;
      25139: inst = 32'hc4046ba;
      25140: inst = 32'h8220000;
      25141: inst = 32'h10408000;
      25142: inst = 32'hc4046bb;
      25143: inst = 32'h8220000;
      25144: inst = 32'h10408000;
      25145: inst = 32'hc4046bc;
      25146: inst = 32'h8220000;
      25147: inst = 32'h10408000;
      25148: inst = 32'hc4046bd;
      25149: inst = 32'h8220000;
      25150: inst = 32'h10408000;
      25151: inst = 32'hc4046be;
      25152: inst = 32'h8220000;
      25153: inst = 32'h10408000;
      25154: inst = 32'hc4046bf;
      25155: inst = 32'h8220000;
      25156: inst = 32'h10408000;
      25157: inst = 32'hc4046c0;
      25158: inst = 32'h8220000;
      25159: inst = 32'h10408000;
      25160: inst = 32'hc4046c1;
      25161: inst = 32'h8220000;
      25162: inst = 32'h10408000;
      25163: inst = 32'hc4046c2;
      25164: inst = 32'h8220000;
      25165: inst = 32'h10408000;
      25166: inst = 32'hc4046c3;
      25167: inst = 32'h8220000;
      25168: inst = 32'h10408000;
      25169: inst = 32'hc4046c4;
      25170: inst = 32'h8220000;
      25171: inst = 32'h10408000;
      25172: inst = 32'hc4046c5;
      25173: inst = 32'h8220000;
      25174: inst = 32'h10408000;
      25175: inst = 32'hc4046c6;
      25176: inst = 32'h8220000;
      25177: inst = 32'h10408000;
      25178: inst = 32'hc4046c7;
      25179: inst = 32'h8220000;
      25180: inst = 32'h10408000;
      25181: inst = 32'hc4046c8;
      25182: inst = 32'h8220000;
      25183: inst = 32'h10408000;
      25184: inst = 32'hc4046c9;
      25185: inst = 32'h8220000;
      25186: inst = 32'h10408000;
      25187: inst = 32'hc4046ca;
      25188: inst = 32'h8220000;
      25189: inst = 32'h10408000;
      25190: inst = 32'hc4046cb;
      25191: inst = 32'h8220000;
      25192: inst = 32'h10408000;
      25193: inst = 32'hc4046cc;
      25194: inst = 32'h8220000;
      25195: inst = 32'h10408000;
      25196: inst = 32'hc4046cd;
      25197: inst = 32'h8220000;
      25198: inst = 32'h10408000;
      25199: inst = 32'hc4046ce;
      25200: inst = 32'h8220000;
      25201: inst = 32'h10408000;
      25202: inst = 32'hc4046cf;
      25203: inst = 32'h8220000;
      25204: inst = 32'h10408000;
      25205: inst = 32'hc4046d0;
      25206: inst = 32'h8220000;
      25207: inst = 32'h10408000;
      25208: inst = 32'hc4046d1;
      25209: inst = 32'h8220000;
      25210: inst = 32'h10408000;
      25211: inst = 32'hc4046d2;
      25212: inst = 32'h8220000;
      25213: inst = 32'h10408000;
      25214: inst = 32'hc4046d3;
      25215: inst = 32'h8220000;
      25216: inst = 32'h10408000;
      25217: inst = 32'hc4046d4;
      25218: inst = 32'h8220000;
      25219: inst = 32'h10408000;
      25220: inst = 32'hc4046d5;
      25221: inst = 32'h8220000;
      25222: inst = 32'h10408000;
      25223: inst = 32'hc4046d6;
      25224: inst = 32'h8220000;
      25225: inst = 32'h10408000;
      25226: inst = 32'hc4046d7;
      25227: inst = 32'h8220000;
      25228: inst = 32'h10408000;
      25229: inst = 32'hc4046d8;
      25230: inst = 32'h8220000;
      25231: inst = 32'h10408000;
      25232: inst = 32'hc4046d9;
      25233: inst = 32'h8220000;
      25234: inst = 32'h10408000;
      25235: inst = 32'hc4046da;
      25236: inst = 32'h8220000;
      25237: inst = 32'h10408000;
      25238: inst = 32'hc4046db;
      25239: inst = 32'h8220000;
      25240: inst = 32'h10408000;
      25241: inst = 32'hc4046dc;
      25242: inst = 32'h8220000;
      25243: inst = 32'h10408000;
      25244: inst = 32'hc4046dd;
      25245: inst = 32'h8220000;
      25246: inst = 32'h10408000;
      25247: inst = 32'hc4046de;
      25248: inst = 32'h8220000;
      25249: inst = 32'h10408000;
      25250: inst = 32'hc4046df;
      25251: inst = 32'h8220000;
      25252: inst = 32'h10408000;
      25253: inst = 32'hc4046e0;
      25254: inst = 32'h8220000;
      25255: inst = 32'h10408000;
      25256: inst = 32'hc4046e1;
      25257: inst = 32'h8220000;
      25258: inst = 32'h10408000;
      25259: inst = 32'hc4046e2;
      25260: inst = 32'h8220000;
      25261: inst = 32'h10408000;
      25262: inst = 32'hc4046e3;
      25263: inst = 32'h8220000;
      25264: inst = 32'h10408000;
      25265: inst = 32'hc4046e4;
      25266: inst = 32'h8220000;
      25267: inst = 32'h10408000;
      25268: inst = 32'hc4046e5;
      25269: inst = 32'h8220000;
      25270: inst = 32'h10408000;
      25271: inst = 32'hc4046e6;
      25272: inst = 32'h8220000;
      25273: inst = 32'h10408000;
      25274: inst = 32'hc4046e7;
      25275: inst = 32'h8220000;
      25276: inst = 32'h10408000;
      25277: inst = 32'hc4046e8;
      25278: inst = 32'h8220000;
      25279: inst = 32'h10408000;
      25280: inst = 32'hc4046e9;
      25281: inst = 32'h8220000;
      25282: inst = 32'h10408000;
      25283: inst = 32'hc4046ea;
      25284: inst = 32'h8220000;
      25285: inst = 32'h10408000;
      25286: inst = 32'hc4046eb;
      25287: inst = 32'h8220000;
      25288: inst = 32'h10408000;
      25289: inst = 32'hc4046ec;
      25290: inst = 32'h8220000;
      25291: inst = 32'h10408000;
      25292: inst = 32'hc4046ed;
      25293: inst = 32'h8220000;
      25294: inst = 32'h10408000;
      25295: inst = 32'hc4046ee;
      25296: inst = 32'h8220000;
      25297: inst = 32'h10408000;
      25298: inst = 32'hc4046ef;
      25299: inst = 32'h8220000;
      25300: inst = 32'h10408000;
      25301: inst = 32'hc4046f3;
      25302: inst = 32'h8220000;
      25303: inst = 32'h10408000;
      25304: inst = 32'hc4046f4;
      25305: inst = 32'h8220000;
      25306: inst = 32'h10408000;
      25307: inst = 32'hc4046f5;
      25308: inst = 32'h8220000;
      25309: inst = 32'h10408000;
      25310: inst = 32'hc4046f6;
      25311: inst = 32'h8220000;
      25312: inst = 32'h10408000;
      25313: inst = 32'hc4046f7;
      25314: inst = 32'h8220000;
      25315: inst = 32'h10408000;
      25316: inst = 32'hc4046f8;
      25317: inst = 32'h8220000;
      25318: inst = 32'h10408000;
      25319: inst = 32'hc404707;
      25320: inst = 32'h8220000;
      25321: inst = 32'h10408000;
      25322: inst = 32'hc404708;
      25323: inst = 32'h8220000;
      25324: inst = 32'h10408000;
      25325: inst = 32'hc404709;
      25326: inst = 32'h8220000;
      25327: inst = 32'h10408000;
      25328: inst = 32'hc40470a;
      25329: inst = 32'h8220000;
      25330: inst = 32'h10408000;
      25331: inst = 32'hc40470b;
      25332: inst = 32'h8220000;
      25333: inst = 32'h10408000;
      25334: inst = 32'hc40470c;
      25335: inst = 32'h8220000;
      25336: inst = 32'h10408000;
      25337: inst = 32'hc40470d;
      25338: inst = 32'h8220000;
      25339: inst = 32'h10408000;
      25340: inst = 32'hc40470e;
      25341: inst = 32'h8220000;
      25342: inst = 32'h10408000;
      25343: inst = 32'hc404711;
      25344: inst = 32'h8220000;
      25345: inst = 32'h10408000;
      25346: inst = 32'hc404712;
      25347: inst = 32'h8220000;
      25348: inst = 32'h10408000;
      25349: inst = 32'hc404713;
      25350: inst = 32'h8220000;
      25351: inst = 32'h10408000;
      25352: inst = 32'hc404714;
      25353: inst = 32'h8220000;
      25354: inst = 32'h10408000;
      25355: inst = 32'hc404717;
      25356: inst = 32'h8220000;
      25357: inst = 32'h10408000;
      25358: inst = 32'hc404718;
      25359: inst = 32'h8220000;
      25360: inst = 32'h10408000;
      25361: inst = 32'hc404719;
      25362: inst = 32'h8220000;
      25363: inst = 32'h10408000;
      25364: inst = 32'hc40471a;
      25365: inst = 32'h8220000;
      25366: inst = 32'h10408000;
      25367: inst = 32'hc40471b;
      25368: inst = 32'h8220000;
      25369: inst = 32'h10408000;
      25370: inst = 32'hc40471c;
      25371: inst = 32'h8220000;
      25372: inst = 32'h10408000;
      25373: inst = 32'hc40471d;
      25374: inst = 32'h8220000;
      25375: inst = 32'h10408000;
      25376: inst = 32'hc40471e;
      25377: inst = 32'h8220000;
      25378: inst = 32'h10408000;
      25379: inst = 32'hc40471f;
      25380: inst = 32'h8220000;
      25381: inst = 32'h10408000;
      25382: inst = 32'hc404720;
      25383: inst = 32'h8220000;
      25384: inst = 32'h10408000;
      25385: inst = 32'hc404721;
      25386: inst = 32'h8220000;
      25387: inst = 32'h10408000;
      25388: inst = 32'hc404722;
      25389: inst = 32'h8220000;
      25390: inst = 32'h10408000;
      25391: inst = 32'hc404723;
      25392: inst = 32'h8220000;
      25393: inst = 32'h10408000;
      25394: inst = 32'hc404726;
      25395: inst = 32'h8220000;
      25396: inst = 32'h10408000;
      25397: inst = 32'hc404727;
      25398: inst = 32'h8220000;
      25399: inst = 32'h10408000;
      25400: inst = 32'hc404728;
      25401: inst = 32'h8220000;
      25402: inst = 32'h10408000;
      25403: inst = 32'hc404729;
      25404: inst = 32'h8220000;
      25405: inst = 32'h10408000;
      25406: inst = 32'hc40472a;
      25407: inst = 32'h8220000;
      25408: inst = 32'h10408000;
      25409: inst = 32'hc40472b;
      25410: inst = 32'h8220000;
      25411: inst = 32'h10408000;
      25412: inst = 32'hc40472c;
      25413: inst = 32'h8220000;
      25414: inst = 32'h10408000;
      25415: inst = 32'hc40472d;
      25416: inst = 32'h8220000;
      25417: inst = 32'h10408000;
      25418: inst = 32'hc40472e;
      25419: inst = 32'h8220000;
      25420: inst = 32'h10408000;
      25421: inst = 32'hc40472f;
      25422: inst = 32'h8220000;
      25423: inst = 32'h10408000;
      25424: inst = 32'hc404730;
      25425: inst = 32'h8220000;
      25426: inst = 32'h10408000;
      25427: inst = 32'hc404731;
      25428: inst = 32'h8220000;
      25429: inst = 32'h10408000;
      25430: inst = 32'hc404732;
      25431: inst = 32'h8220000;
      25432: inst = 32'h10408000;
      25433: inst = 32'hc404733;
      25434: inst = 32'h8220000;
      25435: inst = 32'h10408000;
      25436: inst = 32'hc404734;
      25437: inst = 32'h8220000;
      25438: inst = 32'h10408000;
      25439: inst = 32'hc404735;
      25440: inst = 32'h8220000;
      25441: inst = 32'h10408000;
      25442: inst = 32'hc404736;
      25443: inst = 32'h8220000;
      25444: inst = 32'h10408000;
      25445: inst = 32'hc404737;
      25446: inst = 32'h8220000;
      25447: inst = 32'h10408000;
      25448: inst = 32'hc404738;
      25449: inst = 32'h8220000;
      25450: inst = 32'h10408000;
      25451: inst = 32'hc404739;
      25452: inst = 32'h8220000;
      25453: inst = 32'h10408000;
      25454: inst = 32'hc40473a;
      25455: inst = 32'h8220000;
      25456: inst = 32'h10408000;
      25457: inst = 32'hc40473b;
      25458: inst = 32'h8220000;
      25459: inst = 32'h10408000;
      25460: inst = 32'hc40473c;
      25461: inst = 32'h8220000;
      25462: inst = 32'h10408000;
      25463: inst = 32'hc40473d;
      25464: inst = 32'h8220000;
      25465: inst = 32'h10408000;
      25466: inst = 32'hc40473e;
      25467: inst = 32'h8220000;
      25468: inst = 32'h10408000;
      25469: inst = 32'hc40473f;
      25470: inst = 32'h8220000;
      25471: inst = 32'h10408000;
      25472: inst = 32'hc404740;
      25473: inst = 32'h8220000;
      25474: inst = 32'h10408000;
      25475: inst = 32'hc404741;
      25476: inst = 32'h8220000;
      25477: inst = 32'h10408000;
      25478: inst = 32'hc404744;
      25479: inst = 32'h8220000;
      25480: inst = 32'h10408000;
      25481: inst = 32'hc404745;
      25482: inst = 32'h8220000;
      25483: inst = 32'h10408000;
      25484: inst = 32'hc404746;
      25485: inst = 32'h8220000;
      25486: inst = 32'h10408000;
      25487: inst = 32'hc404747;
      25488: inst = 32'h8220000;
      25489: inst = 32'h10408000;
      25490: inst = 32'hc404748;
      25491: inst = 32'h8220000;
      25492: inst = 32'h10408000;
      25493: inst = 32'hc404749;
      25494: inst = 32'h8220000;
      25495: inst = 32'h10408000;
      25496: inst = 32'hc40474a;
      25497: inst = 32'h8220000;
      25498: inst = 32'h10408000;
      25499: inst = 32'hc40474b;
      25500: inst = 32'h8220000;
      25501: inst = 32'h10408000;
      25502: inst = 32'hc40474c;
      25503: inst = 32'h8220000;
      25504: inst = 32'h10408000;
      25505: inst = 32'hc40474d;
      25506: inst = 32'h8220000;
      25507: inst = 32'h10408000;
      25508: inst = 32'hc40474e;
      25509: inst = 32'h8220000;
      25510: inst = 32'h10408000;
      25511: inst = 32'hc40474f;
      25512: inst = 32'h8220000;
      25513: inst = 32'h10408000;
      25514: inst = 32'hc404750;
      25515: inst = 32'h8220000;
      25516: inst = 32'h10408000;
      25517: inst = 32'hc404753;
      25518: inst = 32'h8220000;
      25519: inst = 32'h10408000;
      25520: inst = 32'hc404754;
      25521: inst = 32'h8220000;
      25522: inst = 32'h10408000;
      25523: inst = 32'hc404755;
      25524: inst = 32'h8220000;
      25525: inst = 32'h10408000;
      25526: inst = 32'hc404756;
      25527: inst = 32'h8220000;
      25528: inst = 32'h10408000;
      25529: inst = 32'hc404757;
      25530: inst = 32'h8220000;
      25531: inst = 32'h10408000;
      25532: inst = 32'hc404758;
      25533: inst = 32'h8220000;
      25534: inst = 32'h10408000;
      25535: inst = 32'hc404767;
      25536: inst = 32'h8220000;
      25537: inst = 32'h10408000;
      25538: inst = 32'hc404768;
      25539: inst = 32'h8220000;
      25540: inst = 32'h10408000;
      25541: inst = 32'hc404769;
      25542: inst = 32'h8220000;
      25543: inst = 32'h10408000;
      25544: inst = 32'hc40476a;
      25545: inst = 32'h8220000;
      25546: inst = 32'h10408000;
      25547: inst = 32'hc40476b;
      25548: inst = 32'h8220000;
      25549: inst = 32'h10408000;
      25550: inst = 32'hc40476c;
      25551: inst = 32'h8220000;
      25552: inst = 32'h10408000;
      25553: inst = 32'hc40476d;
      25554: inst = 32'h8220000;
      25555: inst = 32'h10408000;
      25556: inst = 32'hc40476e;
      25557: inst = 32'h8220000;
      25558: inst = 32'h10408000;
      25559: inst = 32'hc404773;
      25560: inst = 32'h8220000;
      25561: inst = 32'h10408000;
      25562: inst = 32'hc404778;
      25563: inst = 32'h8220000;
      25564: inst = 32'h10408000;
      25565: inst = 32'hc40477d;
      25566: inst = 32'h8220000;
      25567: inst = 32'h10408000;
      25568: inst = 32'hc40477e;
      25569: inst = 32'h8220000;
      25570: inst = 32'h10408000;
      25571: inst = 32'hc40477f;
      25572: inst = 32'h8220000;
      25573: inst = 32'h10408000;
      25574: inst = 32'hc404780;
      25575: inst = 32'h8220000;
      25576: inst = 32'h10408000;
      25577: inst = 32'hc404781;
      25578: inst = 32'h8220000;
      25579: inst = 32'h10408000;
      25580: inst = 32'hc404782;
      25581: inst = 32'h8220000;
      25582: inst = 32'h10408000;
      25583: inst = 32'hc404787;
      25584: inst = 32'h8220000;
      25585: inst = 32'h10408000;
      25586: inst = 32'hc404788;
      25587: inst = 32'h8220000;
      25588: inst = 32'h10408000;
      25589: inst = 32'hc40478c;
      25590: inst = 32'h8220000;
      25591: inst = 32'h10408000;
      25592: inst = 32'hc40478d;
      25593: inst = 32'h8220000;
      25594: inst = 32'h10408000;
      25595: inst = 32'hc40478e;
      25596: inst = 32'h8220000;
      25597: inst = 32'h10408000;
      25598: inst = 32'hc40478f;
      25599: inst = 32'h8220000;
      25600: inst = 32'h10408000;
      25601: inst = 32'hc404790;
      25602: inst = 32'h8220000;
      25603: inst = 32'h10408000;
      25604: inst = 32'hc404791;
      25605: inst = 32'h8220000;
      25606: inst = 32'h10408000;
      25607: inst = 32'hc404792;
      25608: inst = 32'h8220000;
      25609: inst = 32'h10408000;
      25610: inst = 32'hc404796;
      25611: inst = 32'h8220000;
      25612: inst = 32'h10408000;
      25613: inst = 32'hc404797;
      25614: inst = 32'h8220000;
      25615: inst = 32'h10408000;
      25616: inst = 32'hc40479b;
      25617: inst = 32'h8220000;
      25618: inst = 32'h10408000;
      25619: inst = 32'hc4047a0;
      25620: inst = 32'h8220000;
      25621: inst = 32'h10408000;
      25622: inst = 32'hc4047a5;
      25623: inst = 32'h8220000;
      25624: inst = 32'h10408000;
      25625: inst = 32'hc4047a8;
      25626: inst = 32'h8220000;
      25627: inst = 32'h10408000;
      25628: inst = 32'hc4047ab;
      25629: inst = 32'h8220000;
      25630: inst = 32'h10408000;
      25631: inst = 32'hc4047af;
      25632: inst = 32'h8220000;
      25633: inst = 32'h10408000;
      25634: inst = 32'hc4047b0;
      25635: inst = 32'h8220000;
      25636: inst = 32'h10408000;
      25637: inst = 32'hc4047b3;
      25638: inst = 32'h8220000;
      25639: inst = 32'h10408000;
      25640: inst = 32'hc4047b4;
      25641: inst = 32'h8220000;
      25642: inst = 32'h10408000;
      25643: inst = 32'hc4047b5;
      25644: inst = 32'h8220000;
      25645: inst = 32'h10408000;
      25646: inst = 32'hc4047b6;
      25647: inst = 32'h8220000;
      25648: inst = 32'h10408000;
      25649: inst = 32'hc4047b7;
      25650: inst = 32'h8220000;
      25651: inst = 32'h10408000;
      25652: inst = 32'hc4047b8;
      25653: inst = 32'h8220000;
      25654: inst = 32'h10408000;
      25655: inst = 32'hc4047c7;
      25656: inst = 32'h8220000;
      25657: inst = 32'h10408000;
      25658: inst = 32'hc4047c8;
      25659: inst = 32'h8220000;
      25660: inst = 32'h10408000;
      25661: inst = 32'hc4047c9;
      25662: inst = 32'h8220000;
      25663: inst = 32'h10408000;
      25664: inst = 32'hc4047ca;
      25665: inst = 32'h8220000;
      25666: inst = 32'h10408000;
      25667: inst = 32'hc4047cb;
      25668: inst = 32'h8220000;
      25669: inst = 32'h10408000;
      25670: inst = 32'hc4047cc;
      25671: inst = 32'h8220000;
      25672: inst = 32'h10408000;
      25673: inst = 32'hc4047cd;
      25674: inst = 32'h8220000;
      25675: inst = 32'h10408000;
      25676: inst = 32'hc4047ce;
      25677: inst = 32'h8220000;
      25678: inst = 32'h10408000;
      25679: inst = 32'hc4047de;
      25680: inst = 32'h8220000;
      25681: inst = 32'h10408000;
      25682: inst = 32'hc4047df;
      25683: inst = 32'h8220000;
      25684: inst = 32'h10408000;
      25685: inst = 32'hc4047e0;
      25686: inst = 32'h8220000;
      25687: inst = 32'h10408000;
      25688: inst = 32'hc4047e1;
      25689: inst = 32'h8220000;
      25690: inst = 32'h10408000;
      25691: inst = 32'hc4047e2;
      25692: inst = 32'h8220000;
      25693: inst = 32'h10408000;
      25694: inst = 32'hc4047e7;
      25695: inst = 32'h8220000;
      25696: inst = 32'h10408000;
      25697: inst = 32'hc4047ed;
      25698: inst = 32'h8220000;
      25699: inst = 32'h10408000;
      25700: inst = 32'hc4047ee;
      25701: inst = 32'h8220000;
      25702: inst = 32'h10408000;
      25703: inst = 32'hc4047ef;
      25704: inst = 32'h8220000;
      25705: inst = 32'h10408000;
      25706: inst = 32'hc4047f0;
      25707: inst = 32'h8220000;
      25708: inst = 32'h10408000;
      25709: inst = 32'hc4047f1;
      25710: inst = 32'h8220000;
      25711: inst = 32'h10408000;
      25712: inst = 32'hc404810;
      25713: inst = 32'h8220000;
      25714: inst = 32'h10408000;
      25715: inst = 32'hc404813;
      25716: inst = 32'h8220000;
      25717: inst = 32'h10408000;
      25718: inst = 32'hc404814;
      25719: inst = 32'h8220000;
      25720: inst = 32'h10408000;
      25721: inst = 32'hc404815;
      25722: inst = 32'h8220000;
      25723: inst = 32'h10408000;
      25724: inst = 32'hc404816;
      25725: inst = 32'h8220000;
      25726: inst = 32'h10408000;
      25727: inst = 32'hc404817;
      25728: inst = 32'h8220000;
      25729: inst = 32'h10408000;
      25730: inst = 32'hc404818;
      25731: inst = 32'h8220000;
      25732: inst = 32'h10408000;
      25733: inst = 32'hc404827;
      25734: inst = 32'h8220000;
      25735: inst = 32'h10408000;
      25736: inst = 32'hc404828;
      25737: inst = 32'h8220000;
      25738: inst = 32'h10408000;
      25739: inst = 32'hc404829;
      25740: inst = 32'h8220000;
      25741: inst = 32'h10408000;
      25742: inst = 32'hc40482a;
      25743: inst = 32'h8220000;
      25744: inst = 32'h10408000;
      25745: inst = 32'hc40482b;
      25746: inst = 32'h8220000;
      25747: inst = 32'h10408000;
      25748: inst = 32'hc40482c;
      25749: inst = 32'h8220000;
      25750: inst = 32'h10408000;
      25751: inst = 32'hc40482d;
      25752: inst = 32'h8220000;
      25753: inst = 32'h10408000;
      25754: inst = 32'hc40482e;
      25755: inst = 32'h8220000;
      25756: inst = 32'h10408000;
      25757: inst = 32'hc404831;
      25758: inst = 32'h8220000;
      25759: inst = 32'h10408000;
      25760: inst = 32'hc404834;
      25761: inst = 32'h8220000;
      25762: inst = 32'h10408000;
      25763: inst = 32'hc404837;
      25764: inst = 32'h8220000;
      25765: inst = 32'h10408000;
      25766: inst = 32'hc404838;
      25767: inst = 32'h8220000;
      25768: inst = 32'h10408000;
      25769: inst = 32'hc40483b;
      25770: inst = 32'h8220000;
      25771: inst = 32'h10408000;
      25772: inst = 32'hc40483e;
      25773: inst = 32'h8220000;
      25774: inst = 32'h10408000;
      25775: inst = 32'hc40483f;
      25776: inst = 32'h8220000;
      25777: inst = 32'h10408000;
      25778: inst = 32'hc404840;
      25779: inst = 32'h8220000;
      25780: inst = 32'h10408000;
      25781: inst = 32'hc404841;
      25782: inst = 32'h8220000;
      25783: inst = 32'h10408000;
      25784: inst = 32'hc404842;
      25785: inst = 32'h8220000;
      25786: inst = 32'h10408000;
      25787: inst = 32'hc404843;
      25788: inst = 32'h8220000;
      25789: inst = 32'h10408000;
      25790: inst = 32'hc404846;
      25791: inst = 32'h8220000;
      25792: inst = 32'h10408000;
      25793: inst = 32'hc404849;
      25794: inst = 32'h8220000;
      25795: inst = 32'h10408000;
      25796: inst = 32'hc40484a;
      25797: inst = 32'h8220000;
      25798: inst = 32'h10408000;
      25799: inst = 32'hc40484d;
      25800: inst = 32'h8220000;
      25801: inst = 32'h10408000;
      25802: inst = 32'hc40484e;
      25803: inst = 32'h8220000;
      25804: inst = 32'h10408000;
      25805: inst = 32'hc40484f;
      25806: inst = 32'h8220000;
      25807: inst = 32'h10408000;
      25808: inst = 32'hc404850;
      25809: inst = 32'h8220000;
      25810: inst = 32'h10408000;
      25811: inst = 32'hc404851;
      25812: inst = 32'h8220000;
      25813: inst = 32'h10408000;
      25814: inst = 32'hc404854;
      25815: inst = 32'h8220000;
      25816: inst = 32'h10408000;
      25817: inst = 32'hc404858;
      25818: inst = 32'h8220000;
      25819: inst = 32'h10408000;
      25820: inst = 32'hc404859;
      25821: inst = 32'h8220000;
      25822: inst = 32'h10408000;
      25823: inst = 32'hc40485e;
      25824: inst = 32'h8220000;
      25825: inst = 32'h10408000;
      25826: inst = 32'hc404861;
      25827: inst = 32'h8220000;
      25828: inst = 32'h10408000;
      25829: inst = 32'hc404864;
      25830: inst = 32'h8220000;
      25831: inst = 32'h10408000;
      25832: inst = 32'hc404865;
      25833: inst = 32'h8220000;
      25834: inst = 32'h10408000;
      25835: inst = 32'hc404869;
      25836: inst = 32'h8220000;
      25837: inst = 32'h10408000;
      25838: inst = 32'hc40486c;
      25839: inst = 32'h8220000;
      25840: inst = 32'h10408000;
      25841: inst = 32'hc40486d;
      25842: inst = 32'h8220000;
      25843: inst = 32'h10408000;
      25844: inst = 32'hc404870;
      25845: inst = 32'h8220000;
      25846: inst = 32'h10408000;
      25847: inst = 32'hc404873;
      25848: inst = 32'h8220000;
      25849: inst = 32'h10408000;
      25850: inst = 32'hc404874;
      25851: inst = 32'h8220000;
      25852: inst = 32'h10408000;
      25853: inst = 32'hc404875;
      25854: inst = 32'h8220000;
      25855: inst = 32'h10408000;
      25856: inst = 32'hc404876;
      25857: inst = 32'h8220000;
      25858: inst = 32'h10408000;
      25859: inst = 32'hc404877;
      25860: inst = 32'h8220000;
      25861: inst = 32'h10408000;
      25862: inst = 32'hc404878;
      25863: inst = 32'h8220000;
      25864: inst = 32'h10408000;
      25865: inst = 32'hc404887;
      25866: inst = 32'h8220000;
      25867: inst = 32'h10408000;
      25868: inst = 32'hc404888;
      25869: inst = 32'h8220000;
      25870: inst = 32'h10408000;
      25871: inst = 32'hc404889;
      25872: inst = 32'h8220000;
      25873: inst = 32'h10408000;
      25874: inst = 32'hc40488a;
      25875: inst = 32'h8220000;
      25876: inst = 32'h10408000;
      25877: inst = 32'hc40488b;
      25878: inst = 32'h8220000;
      25879: inst = 32'h10408000;
      25880: inst = 32'hc40488c;
      25881: inst = 32'h8220000;
      25882: inst = 32'h10408000;
      25883: inst = 32'hc40488d;
      25884: inst = 32'h8220000;
      25885: inst = 32'h10408000;
      25886: inst = 32'hc40488e;
      25887: inst = 32'h8220000;
      25888: inst = 32'h10408000;
      25889: inst = 32'hc404891;
      25890: inst = 32'h8220000;
      25891: inst = 32'h10408000;
      25892: inst = 32'hc404894;
      25893: inst = 32'h8220000;
      25894: inst = 32'h10408000;
      25895: inst = 32'hc404897;
      25896: inst = 32'h8220000;
      25897: inst = 32'h10408000;
      25898: inst = 32'hc404898;
      25899: inst = 32'h8220000;
      25900: inst = 32'h10408000;
      25901: inst = 32'hc40489b;
      25902: inst = 32'h8220000;
      25903: inst = 32'h10408000;
      25904: inst = 32'hc40489e;
      25905: inst = 32'h8220000;
      25906: inst = 32'h10408000;
      25907: inst = 32'hc40489f;
      25908: inst = 32'h8220000;
      25909: inst = 32'h10408000;
      25910: inst = 32'hc4048a0;
      25911: inst = 32'h8220000;
      25912: inst = 32'h10408000;
      25913: inst = 32'hc4048a1;
      25914: inst = 32'h8220000;
      25915: inst = 32'h10408000;
      25916: inst = 32'hc4048a2;
      25917: inst = 32'h8220000;
      25918: inst = 32'h10408000;
      25919: inst = 32'hc4048a3;
      25920: inst = 32'h8220000;
      25921: inst = 32'h10408000;
      25922: inst = 32'hc4048a6;
      25923: inst = 32'h8220000;
      25924: inst = 32'h10408000;
      25925: inst = 32'hc4048a9;
      25926: inst = 32'h8220000;
      25927: inst = 32'h10408000;
      25928: inst = 32'hc4048aa;
      25929: inst = 32'h8220000;
      25930: inst = 32'h10408000;
      25931: inst = 32'hc4048ad;
      25932: inst = 32'h8220000;
      25933: inst = 32'h10408000;
      25934: inst = 32'hc4048ae;
      25935: inst = 32'h8220000;
      25936: inst = 32'h10408000;
      25937: inst = 32'hc4048af;
      25938: inst = 32'h8220000;
      25939: inst = 32'h10408000;
      25940: inst = 32'hc4048b0;
      25941: inst = 32'h8220000;
      25942: inst = 32'h10408000;
      25943: inst = 32'hc4048b3;
      25944: inst = 32'h8220000;
      25945: inst = 32'h10408000;
      25946: inst = 32'hc4048b4;
      25947: inst = 32'h8220000;
      25948: inst = 32'h10408000;
      25949: inst = 32'hc4048b5;
      25950: inst = 32'h8220000;
      25951: inst = 32'h10408000;
      25952: inst = 32'hc4048b8;
      25953: inst = 32'h8220000;
      25954: inst = 32'h10408000;
      25955: inst = 32'hc4048b9;
      25956: inst = 32'h8220000;
      25957: inst = 32'h10408000;
      25958: inst = 32'hc4048be;
      25959: inst = 32'h8220000;
      25960: inst = 32'h10408000;
      25961: inst = 32'hc4048c1;
      25962: inst = 32'h8220000;
      25963: inst = 32'h10408000;
      25964: inst = 32'hc4048c4;
      25965: inst = 32'h8220000;
      25966: inst = 32'h10408000;
      25967: inst = 32'hc4048c5;
      25968: inst = 32'h8220000;
      25969: inst = 32'h10408000;
      25970: inst = 32'hc4048c8;
      25971: inst = 32'h8220000;
      25972: inst = 32'h10408000;
      25973: inst = 32'hc4048c9;
      25974: inst = 32'h8220000;
      25975: inst = 32'h10408000;
      25976: inst = 32'hc4048cc;
      25977: inst = 32'h8220000;
      25978: inst = 32'h10408000;
      25979: inst = 32'hc4048cd;
      25980: inst = 32'h8220000;
      25981: inst = 32'h10408000;
      25982: inst = 32'hc4048d0;
      25983: inst = 32'h8220000;
      25984: inst = 32'h10408000;
      25985: inst = 32'hc4048d3;
      25986: inst = 32'h8220000;
      25987: inst = 32'h10408000;
      25988: inst = 32'hc4048d4;
      25989: inst = 32'h8220000;
      25990: inst = 32'h10408000;
      25991: inst = 32'hc4048d5;
      25992: inst = 32'h8220000;
      25993: inst = 32'h10408000;
      25994: inst = 32'hc4048d6;
      25995: inst = 32'h8220000;
      25996: inst = 32'h10408000;
      25997: inst = 32'hc4048d7;
      25998: inst = 32'h8220000;
      25999: inst = 32'h10408000;
      26000: inst = 32'hc4048d8;
      26001: inst = 32'h8220000;
      26002: inst = 32'h10408000;
      26003: inst = 32'hc4048e7;
      26004: inst = 32'h8220000;
      26005: inst = 32'h10408000;
      26006: inst = 32'hc4048e8;
      26007: inst = 32'h8220000;
      26008: inst = 32'h10408000;
      26009: inst = 32'hc4048e9;
      26010: inst = 32'h8220000;
      26011: inst = 32'h10408000;
      26012: inst = 32'hc4048ea;
      26013: inst = 32'h8220000;
      26014: inst = 32'h10408000;
      26015: inst = 32'hc4048eb;
      26016: inst = 32'h8220000;
      26017: inst = 32'h10408000;
      26018: inst = 32'hc4048ec;
      26019: inst = 32'h8220000;
      26020: inst = 32'h10408000;
      26021: inst = 32'hc4048ed;
      26022: inst = 32'h8220000;
      26023: inst = 32'h10408000;
      26024: inst = 32'hc4048ee;
      26025: inst = 32'h8220000;
      26026: inst = 32'h10408000;
      26027: inst = 32'hc4048f1;
      26028: inst = 32'h8220000;
      26029: inst = 32'h10408000;
      26030: inst = 32'hc4048f4;
      26031: inst = 32'h8220000;
      26032: inst = 32'h10408000;
      26033: inst = 32'hc4048f7;
      26034: inst = 32'h8220000;
      26035: inst = 32'h10408000;
      26036: inst = 32'hc4048f8;
      26037: inst = 32'h8220000;
      26038: inst = 32'h10408000;
      26039: inst = 32'hc4048fb;
      26040: inst = 32'h8220000;
      26041: inst = 32'h10408000;
      26042: inst = 32'hc4048fe;
      26043: inst = 32'h8220000;
      26044: inst = 32'h10408000;
      26045: inst = 32'hc4048ff;
      26046: inst = 32'h8220000;
      26047: inst = 32'h10408000;
      26048: inst = 32'hc404900;
      26049: inst = 32'h8220000;
      26050: inst = 32'h10408000;
      26051: inst = 32'hc404901;
      26052: inst = 32'h8220000;
      26053: inst = 32'h10408000;
      26054: inst = 32'hc404902;
      26055: inst = 32'h8220000;
      26056: inst = 32'h10408000;
      26057: inst = 32'hc404903;
      26058: inst = 32'h8220000;
      26059: inst = 32'h10408000;
      26060: inst = 32'hc404906;
      26061: inst = 32'h8220000;
      26062: inst = 32'h10408000;
      26063: inst = 32'hc404909;
      26064: inst = 32'h8220000;
      26065: inst = 32'h10408000;
      26066: inst = 32'hc40490a;
      26067: inst = 32'h8220000;
      26068: inst = 32'h10408000;
      26069: inst = 32'hc40490d;
      26070: inst = 32'h8220000;
      26071: inst = 32'h10408000;
      26072: inst = 32'hc40490e;
      26073: inst = 32'h8220000;
      26074: inst = 32'h10408000;
      26075: inst = 32'hc40490f;
      26076: inst = 32'h8220000;
      26077: inst = 32'h10408000;
      26078: inst = 32'hc404910;
      26079: inst = 32'h8220000;
      26080: inst = 32'h10408000;
      26081: inst = 32'hc404913;
      26082: inst = 32'h8220000;
      26083: inst = 32'h10408000;
      26084: inst = 32'hc404914;
      26085: inst = 32'h8220000;
      26086: inst = 32'h10408000;
      26087: inst = 32'hc404915;
      26088: inst = 32'h8220000;
      26089: inst = 32'h10408000;
      26090: inst = 32'hc404918;
      26091: inst = 32'h8220000;
      26092: inst = 32'h10408000;
      26093: inst = 32'hc404919;
      26094: inst = 32'h8220000;
      26095: inst = 32'h10408000;
      26096: inst = 32'hc40491e;
      26097: inst = 32'h8220000;
      26098: inst = 32'h10408000;
      26099: inst = 32'hc404921;
      26100: inst = 32'h8220000;
      26101: inst = 32'h10408000;
      26102: inst = 32'hc404924;
      26103: inst = 32'h8220000;
      26104: inst = 32'h10408000;
      26105: inst = 32'hc404925;
      26106: inst = 32'h8220000;
      26107: inst = 32'h10408000;
      26108: inst = 32'hc404928;
      26109: inst = 32'h8220000;
      26110: inst = 32'h10408000;
      26111: inst = 32'hc404929;
      26112: inst = 32'h8220000;
      26113: inst = 32'h10408000;
      26114: inst = 32'hc40492c;
      26115: inst = 32'h8220000;
      26116: inst = 32'h10408000;
      26117: inst = 32'hc40492d;
      26118: inst = 32'h8220000;
      26119: inst = 32'h10408000;
      26120: inst = 32'hc404930;
      26121: inst = 32'h8220000;
      26122: inst = 32'h10408000;
      26123: inst = 32'hc404933;
      26124: inst = 32'h8220000;
      26125: inst = 32'h10408000;
      26126: inst = 32'hc404934;
      26127: inst = 32'h8220000;
      26128: inst = 32'h10408000;
      26129: inst = 32'hc404935;
      26130: inst = 32'h8220000;
      26131: inst = 32'h10408000;
      26132: inst = 32'hc404936;
      26133: inst = 32'h8220000;
      26134: inst = 32'h10408000;
      26135: inst = 32'hc404937;
      26136: inst = 32'h8220000;
      26137: inst = 32'h10408000;
      26138: inst = 32'hc404938;
      26139: inst = 32'h8220000;
      26140: inst = 32'h10408000;
      26141: inst = 32'hc404947;
      26142: inst = 32'h8220000;
      26143: inst = 32'h10408000;
      26144: inst = 32'hc404948;
      26145: inst = 32'h8220000;
      26146: inst = 32'h10408000;
      26147: inst = 32'hc404949;
      26148: inst = 32'h8220000;
      26149: inst = 32'h10408000;
      26150: inst = 32'hc40494a;
      26151: inst = 32'h8220000;
      26152: inst = 32'h10408000;
      26153: inst = 32'hc40494b;
      26154: inst = 32'h8220000;
      26155: inst = 32'h10408000;
      26156: inst = 32'hc40494c;
      26157: inst = 32'h8220000;
      26158: inst = 32'h10408000;
      26159: inst = 32'hc40494d;
      26160: inst = 32'h8220000;
      26161: inst = 32'h10408000;
      26162: inst = 32'hc40494e;
      26163: inst = 32'h8220000;
      26164: inst = 32'h10408000;
      26165: inst = 32'hc404951;
      26166: inst = 32'h8220000;
      26167: inst = 32'h10408000;
      26168: inst = 32'hc404954;
      26169: inst = 32'h8220000;
      26170: inst = 32'h10408000;
      26171: inst = 32'hc404957;
      26172: inst = 32'h8220000;
      26173: inst = 32'h10408000;
      26174: inst = 32'hc40495b;
      26175: inst = 32'h8220000;
      26176: inst = 32'h10408000;
      26177: inst = 32'hc40495e;
      26178: inst = 32'h8220000;
      26179: inst = 32'h10408000;
      26180: inst = 32'hc40495f;
      26181: inst = 32'h8220000;
      26182: inst = 32'h10408000;
      26183: inst = 32'hc404960;
      26184: inst = 32'h8220000;
      26185: inst = 32'h10408000;
      26186: inst = 32'hc404961;
      26187: inst = 32'h8220000;
      26188: inst = 32'h10408000;
      26189: inst = 32'hc404962;
      26190: inst = 32'h8220000;
      26191: inst = 32'h10408000;
      26192: inst = 32'hc404963;
      26193: inst = 32'h8220000;
      26194: inst = 32'h10408000;
      26195: inst = 32'hc404966;
      26196: inst = 32'h8220000;
      26197: inst = 32'h10408000;
      26198: inst = 32'hc404969;
      26199: inst = 32'h8220000;
      26200: inst = 32'h10408000;
      26201: inst = 32'hc40496a;
      26202: inst = 32'h8220000;
      26203: inst = 32'h10408000;
      26204: inst = 32'hc40496d;
      26205: inst = 32'h8220000;
      26206: inst = 32'h10408000;
      26207: inst = 32'hc40496e;
      26208: inst = 32'h8220000;
      26209: inst = 32'h10408000;
      26210: inst = 32'hc40496f;
      26211: inst = 32'h8220000;
      26212: inst = 32'h10408000;
      26213: inst = 32'hc404970;
      26214: inst = 32'h8220000;
      26215: inst = 32'h10408000;
      26216: inst = 32'hc404974;
      26217: inst = 32'h8220000;
      26218: inst = 32'h10408000;
      26219: inst = 32'hc404975;
      26220: inst = 32'h8220000;
      26221: inst = 32'h10408000;
      26222: inst = 32'hc404978;
      26223: inst = 32'h8220000;
      26224: inst = 32'h10408000;
      26225: inst = 32'hc404979;
      26226: inst = 32'h8220000;
      26227: inst = 32'h10408000;
      26228: inst = 32'hc40497e;
      26229: inst = 32'h8220000;
      26230: inst = 32'h10408000;
      26231: inst = 32'hc404981;
      26232: inst = 32'h8220000;
      26233: inst = 32'h10408000;
      26234: inst = 32'hc404984;
      26235: inst = 32'h8220000;
      26236: inst = 32'h10408000;
      26237: inst = 32'hc404988;
      26238: inst = 32'h8220000;
      26239: inst = 32'h10408000;
      26240: inst = 32'hc404989;
      26241: inst = 32'h8220000;
      26242: inst = 32'h10408000;
      26243: inst = 32'hc40498c;
      26244: inst = 32'h8220000;
      26245: inst = 32'h10408000;
      26246: inst = 32'hc40498d;
      26247: inst = 32'h8220000;
      26248: inst = 32'h10408000;
      26249: inst = 32'hc404990;
      26250: inst = 32'h8220000;
      26251: inst = 32'h10408000;
      26252: inst = 32'hc404993;
      26253: inst = 32'h8220000;
      26254: inst = 32'h10408000;
      26255: inst = 32'hc404994;
      26256: inst = 32'h8220000;
      26257: inst = 32'h10408000;
      26258: inst = 32'hc404995;
      26259: inst = 32'h8220000;
      26260: inst = 32'h10408000;
      26261: inst = 32'hc404996;
      26262: inst = 32'h8220000;
      26263: inst = 32'h10408000;
      26264: inst = 32'hc404997;
      26265: inst = 32'h8220000;
      26266: inst = 32'h10408000;
      26267: inst = 32'hc404998;
      26268: inst = 32'h8220000;
      26269: inst = 32'h10408000;
      26270: inst = 32'hc4049a7;
      26271: inst = 32'h8220000;
      26272: inst = 32'h10408000;
      26273: inst = 32'hc4049a8;
      26274: inst = 32'h8220000;
      26275: inst = 32'h10408000;
      26276: inst = 32'hc4049a9;
      26277: inst = 32'h8220000;
      26278: inst = 32'h10408000;
      26279: inst = 32'hc4049aa;
      26280: inst = 32'h8220000;
      26281: inst = 32'h10408000;
      26282: inst = 32'hc4049ab;
      26283: inst = 32'h8220000;
      26284: inst = 32'h10408000;
      26285: inst = 32'hc4049ac;
      26286: inst = 32'h8220000;
      26287: inst = 32'h10408000;
      26288: inst = 32'hc4049ad;
      26289: inst = 32'h8220000;
      26290: inst = 32'h10408000;
      26291: inst = 32'hc4049ae;
      26292: inst = 32'h8220000;
      26293: inst = 32'h10408000;
      26294: inst = 32'hc4049b4;
      26295: inst = 32'h8220000;
      26296: inst = 32'h10408000;
      26297: inst = 32'hc4049bb;
      26298: inst = 32'h8220000;
      26299: inst = 32'h10408000;
      26300: inst = 32'hc4049be;
      26301: inst = 32'h8220000;
      26302: inst = 32'h10408000;
      26303: inst = 32'hc4049bf;
      26304: inst = 32'h8220000;
      26305: inst = 32'h10408000;
      26306: inst = 32'hc4049c0;
      26307: inst = 32'h8220000;
      26308: inst = 32'h10408000;
      26309: inst = 32'hc4049c1;
      26310: inst = 32'h8220000;
      26311: inst = 32'h10408000;
      26312: inst = 32'hc4049c2;
      26313: inst = 32'h8220000;
      26314: inst = 32'h10408000;
      26315: inst = 32'hc4049c3;
      26316: inst = 32'h8220000;
      26317: inst = 32'h10408000;
      26318: inst = 32'hc4049cd;
      26319: inst = 32'h8220000;
      26320: inst = 32'h10408000;
      26321: inst = 32'hc4049ce;
      26322: inst = 32'h8220000;
      26323: inst = 32'h10408000;
      26324: inst = 32'hc4049cf;
      26325: inst = 32'h8220000;
      26326: inst = 32'h10408000;
      26327: inst = 32'hc4049d0;
      26328: inst = 32'h8220000;
      26329: inst = 32'h10408000;
      26330: inst = 32'hc4049d1;
      26331: inst = 32'h8220000;
      26332: inst = 32'h10408000;
      26333: inst = 32'hc4049de;
      26334: inst = 32'h8220000;
      26335: inst = 32'h10408000;
      26336: inst = 32'hc4049e1;
      26337: inst = 32'h8220000;
      26338: inst = 32'h10408000;
      26339: inst = 32'hc4049ea;
      26340: inst = 32'h8220000;
      26341: inst = 32'h10408000;
      26342: inst = 32'hc4049f5;
      26343: inst = 32'h8220000;
      26344: inst = 32'h10408000;
      26345: inst = 32'hc4049f6;
      26346: inst = 32'h8220000;
      26347: inst = 32'h10408000;
      26348: inst = 32'hc4049f7;
      26349: inst = 32'h8220000;
      26350: inst = 32'h10408000;
      26351: inst = 32'hc4049f8;
      26352: inst = 32'h8220000;
      26353: inst = 32'h10408000;
      26354: inst = 32'hc404a07;
      26355: inst = 32'h8220000;
      26356: inst = 32'h10408000;
      26357: inst = 32'hc404a08;
      26358: inst = 32'h8220000;
      26359: inst = 32'h10408000;
      26360: inst = 32'hc404a09;
      26361: inst = 32'h8220000;
      26362: inst = 32'h10408000;
      26363: inst = 32'hc404a0a;
      26364: inst = 32'h8220000;
      26365: inst = 32'h10408000;
      26366: inst = 32'hc404a0b;
      26367: inst = 32'h8220000;
      26368: inst = 32'h10408000;
      26369: inst = 32'hc404a0c;
      26370: inst = 32'h8220000;
      26371: inst = 32'h10408000;
      26372: inst = 32'hc404a0d;
      26373: inst = 32'h8220000;
      26374: inst = 32'h10408000;
      26375: inst = 32'hc404a0e;
      26376: inst = 32'h8220000;
      26377: inst = 32'h10408000;
      26378: inst = 32'hc404a0f;
      26379: inst = 32'h8220000;
      26380: inst = 32'h10408000;
      26381: inst = 32'hc404a12;
      26382: inst = 32'h8220000;
      26383: inst = 32'h10408000;
      26384: inst = 32'hc404a13;
      26385: inst = 32'h8220000;
      26386: inst = 32'h10408000;
      26387: inst = 32'hc404a14;
      26388: inst = 32'h8220000;
      26389: inst = 32'h10408000;
      26390: inst = 32'hc404a15;
      26391: inst = 32'h8220000;
      26392: inst = 32'h10408000;
      26393: inst = 32'hc404a1b;
      26394: inst = 32'h8220000;
      26395: inst = 32'h10408000;
      26396: inst = 32'hc404a1e;
      26397: inst = 32'h8220000;
      26398: inst = 32'h10408000;
      26399: inst = 32'hc404a1f;
      26400: inst = 32'h8220000;
      26401: inst = 32'h10408000;
      26402: inst = 32'hc404a20;
      26403: inst = 32'h8220000;
      26404: inst = 32'h10408000;
      26405: inst = 32'hc404a21;
      26406: inst = 32'h8220000;
      26407: inst = 32'h10408000;
      26408: inst = 32'hc404a22;
      26409: inst = 32'h8220000;
      26410: inst = 32'h10408000;
      26411: inst = 32'hc404a23;
      26412: inst = 32'h8220000;
      26413: inst = 32'h10408000;
      26414: inst = 32'hc404a24;
      26415: inst = 32'h8220000;
      26416: inst = 32'h10408000;
      26417: inst = 32'hc404a27;
      26418: inst = 32'h8220000;
      26419: inst = 32'h10408000;
      26420: inst = 32'hc404a28;
      26421: inst = 32'h8220000;
      26422: inst = 32'h10408000;
      26423: inst = 32'hc404a2b;
      26424: inst = 32'h8220000;
      26425: inst = 32'h10408000;
      26426: inst = 32'hc404a2c;
      26427: inst = 32'h8220000;
      26428: inst = 32'h10408000;
      26429: inst = 32'hc404a2d;
      26430: inst = 32'h8220000;
      26431: inst = 32'h10408000;
      26432: inst = 32'hc404a2e;
      26433: inst = 32'h8220000;
      26434: inst = 32'h10408000;
      26435: inst = 32'hc404a2f;
      26436: inst = 32'h8220000;
      26437: inst = 32'h10408000;
      26438: inst = 32'hc404a30;
      26439: inst = 32'h8220000;
      26440: inst = 32'h10408000;
      26441: inst = 32'hc404a31;
      26442: inst = 32'h8220000;
      26443: inst = 32'h10408000;
      26444: inst = 32'hc404a32;
      26445: inst = 32'h8220000;
      26446: inst = 32'h10408000;
      26447: inst = 32'hc404a36;
      26448: inst = 32'h8220000;
      26449: inst = 32'h10408000;
      26450: inst = 32'hc404a37;
      26451: inst = 32'h8220000;
      26452: inst = 32'h10408000;
      26453: inst = 32'hc404a3a;
      26454: inst = 32'h8220000;
      26455: inst = 32'h10408000;
      26456: inst = 32'hc404a3e;
      26457: inst = 32'h8220000;
      26458: inst = 32'h10408000;
      26459: inst = 32'hc404a41;
      26460: inst = 32'h8220000;
      26461: inst = 32'h10408000;
      26462: inst = 32'hc404a42;
      26463: inst = 32'h8220000;
      26464: inst = 32'h10408000;
      26465: inst = 32'hc404a49;
      26466: inst = 32'h8220000;
      26467: inst = 32'h10408000;
      26468: inst = 32'hc404a4a;
      26469: inst = 32'h8220000;
      26470: inst = 32'h10408000;
      26471: inst = 32'hc404a4b;
      26472: inst = 32'h8220000;
      26473: inst = 32'h10408000;
      26474: inst = 32'hc404a4e;
      26475: inst = 32'h8220000;
      26476: inst = 32'h10408000;
      26477: inst = 32'hc404a4f;
      26478: inst = 32'h8220000;
      26479: inst = 32'h10408000;
      26480: inst = 32'hc404a54;
      26481: inst = 32'h8220000;
      26482: inst = 32'h10408000;
      26483: inst = 32'hc404a55;
      26484: inst = 32'h8220000;
      26485: inst = 32'h10408000;
      26486: inst = 32'hc404a56;
      26487: inst = 32'h8220000;
      26488: inst = 32'h10408000;
      26489: inst = 32'hc404a57;
      26490: inst = 32'h8220000;
      26491: inst = 32'h10408000;
      26492: inst = 32'hc404a58;
      26493: inst = 32'h8220000;
      26494: inst = 32'h10408000;
      26495: inst = 32'hc404a67;
      26496: inst = 32'h8220000;
      26497: inst = 32'h10408000;
      26498: inst = 32'hc404a68;
      26499: inst = 32'h8220000;
      26500: inst = 32'h10408000;
      26501: inst = 32'hc404a69;
      26502: inst = 32'h8220000;
      26503: inst = 32'h10408000;
      26504: inst = 32'hc404a6a;
      26505: inst = 32'h8220000;
      26506: inst = 32'h10408000;
      26507: inst = 32'hc404a6b;
      26508: inst = 32'h8220000;
      26509: inst = 32'h10408000;
      26510: inst = 32'hc404a6c;
      26511: inst = 32'h8220000;
      26512: inst = 32'h10408000;
      26513: inst = 32'hc404a6d;
      26514: inst = 32'h8220000;
      26515: inst = 32'h10408000;
      26516: inst = 32'hc404a6e;
      26517: inst = 32'h8220000;
      26518: inst = 32'h10408000;
      26519: inst = 32'hc404a6f;
      26520: inst = 32'h8220000;
      26521: inst = 32'h10408000;
      26522: inst = 32'hc404a70;
      26523: inst = 32'h8220000;
      26524: inst = 32'h10408000;
      26525: inst = 32'hc404a71;
      26526: inst = 32'h8220000;
      26527: inst = 32'h10408000;
      26528: inst = 32'hc404a72;
      26529: inst = 32'h8220000;
      26530: inst = 32'h10408000;
      26531: inst = 32'hc404a73;
      26532: inst = 32'h8220000;
      26533: inst = 32'h10408000;
      26534: inst = 32'hc404a74;
      26535: inst = 32'h8220000;
      26536: inst = 32'h10408000;
      26537: inst = 32'hc404a75;
      26538: inst = 32'h8220000;
      26539: inst = 32'h10408000;
      26540: inst = 32'hc404a76;
      26541: inst = 32'h8220000;
      26542: inst = 32'h10408000;
      26543: inst = 32'hc404a77;
      26544: inst = 32'h8220000;
      26545: inst = 32'h10408000;
      26546: inst = 32'hc404a78;
      26547: inst = 32'h8220000;
      26548: inst = 32'h10408000;
      26549: inst = 32'hc404a79;
      26550: inst = 32'h8220000;
      26551: inst = 32'h10408000;
      26552: inst = 32'hc404a7a;
      26553: inst = 32'h8220000;
      26554: inst = 32'h10408000;
      26555: inst = 32'hc404a7b;
      26556: inst = 32'h8220000;
      26557: inst = 32'h10408000;
      26558: inst = 32'hc404a7c;
      26559: inst = 32'h8220000;
      26560: inst = 32'h10408000;
      26561: inst = 32'hc404a7d;
      26562: inst = 32'h8220000;
      26563: inst = 32'h10408000;
      26564: inst = 32'hc404a7e;
      26565: inst = 32'h8220000;
      26566: inst = 32'h10408000;
      26567: inst = 32'hc404a7f;
      26568: inst = 32'h8220000;
      26569: inst = 32'h10408000;
      26570: inst = 32'hc404a80;
      26571: inst = 32'h8220000;
      26572: inst = 32'h10408000;
      26573: inst = 32'hc404a81;
      26574: inst = 32'h8220000;
      26575: inst = 32'h10408000;
      26576: inst = 32'hc404a82;
      26577: inst = 32'h8220000;
      26578: inst = 32'h10408000;
      26579: inst = 32'hc404a83;
      26580: inst = 32'h8220000;
      26581: inst = 32'h10408000;
      26582: inst = 32'hc404a84;
      26583: inst = 32'h8220000;
      26584: inst = 32'h10408000;
      26585: inst = 32'hc404a85;
      26586: inst = 32'h8220000;
      26587: inst = 32'h10408000;
      26588: inst = 32'hc404a86;
      26589: inst = 32'h8220000;
      26590: inst = 32'h10408000;
      26591: inst = 32'hc404a87;
      26592: inst = 32'h8220000;
      26593: inst = 32'h10408000;
      26594: inst = 32'hc404a88;
      26595: inst = 32'h8220000;
      26596: inst = 32'h10408000;
      26597: inst = 32'hc404a89;
      26598: inst = 32'h8220000;
      26599: inst = 32'h10408000;
      26600: inst = 32'hc404a8a;
      26601: inst = 32'h8220000;
      26602: inst = 32'h10408000;
      26603: inst = 32'hc404a8b;
      26604: inst = 32'h8220000;
      26605: inst = 32'h10408000;
      26606: inst = 32'hc404a8c;
      26607: inst = 32'h8220000;
      26608: inst = 32'h10408000;
      26609: inst = 32'hc404a8d;
      26610: inst = 32'h8220000;
      26611: inst = 32'h10408000;
      26612: inst = 32'hc404a8e;
      26613: inst = 32'h8220000;
      26614: inst = 32'h10408000;
      26615: inst = 32'hc404a8f;
      26616: inst = 32'h8220000;
      26617: inst = 32'h10408000;
      26618: inst = 32'hc404a90;
      26619: inst = 32'h8220000;
      26620: inst = 32'h10408000;
      26621: inst = 32'hc404a91;
      26622: inst = 32'h8220000;
      26623: inst = 32'h10408000;
      26624: inst = 32'hc404a92;
      26625: inst = 32'h8220000;
      26626: inst = 32'h10408000;
      26627: inst = 32'hc404a93;
      26628: inst = 32'h8220000;
      26629: inst = 32'h10408000;
      26630: inst = 32'hc404a94;
      26631: inst = 32'h8220000;
      26632: inst = 32'h10408000;
      26633: inst = 32'hc404a95;
      26634: inst = 32'h8220000;
      26635: inst = 32'h10408000;
      26636: inst = 32'hc404a96;
      26637: inst = 32'h8220000;
      26638: inst = 32'h10408000;
      26639: inst = 32'hc404a97;
      26640: inst = 32'h8220000;
      26641: inst = 32'h10408000;
      26642: inst = 32'hc404a98;
      26643: inst = 32'h8220000;
      26644: inst = 32'h10408000;
      26645: inst = 32'hc404a99;
      26646: inst = 32'h8220000;
      26647: inst = 32'h10408000;
      26648: inst = 32'hc404a9a;
      26649: inst = 32'h8220000;
      26650: inst = 32'h10408000;
      26651: inst = 32'hc404a9b;
      26652: inst = 32'h8220000;
      26653: inst = 32'h10408000;
      26654: inst = 32'hc404a9c;
      26655: inst = 32'h8220000;
      26656: inst = 32'h10408000;
      26657: inst = 32'hc404a9d;
      26658: inst = 32'h8220000;
      26659: inst = 32'h10408000;
      26660: inst = 32'hc404a9e;
      26661: inst = 32'h8220000;
      26662: inst = 32'h10408000;
      26663: inst = 32'hc404a9f;
      26664: inst = 32'h8220000;
      26665: inst = 32'h10408000;
      26666: inst = 32'hc404aa0;
      26667: inst = 32'h8220000;
      26668: inst = 32'h10408000;
      26669: inst = 32'hc404aa1;
      26670: inst = 32'h8220000;
      26671: inst = 32'h10408000;
      26672: inst = 32'hc404aa2;
      26673: inst = 32'h8220000;
      26674: inst = 32'h10408000;
      26675: inst = 32'hc404aa3;
      26676: inst = 32'h8220000;
      26677: inst = 32'h10408000;
      26678: inst = 32'hc404aa4;
      26679: inst = 32'h8220000;
      26680: inst = 32'h10408000;
      26681: inst = 32'hc404aa5;
      26682: inst = 32'h8220000;
      26683: inst = 32'h10408000;
      26684: inst = 32'hc404aa6;
      26685: inst = 32'h8220000;
      26686: inst = 32'h10408000;
      26687: inst = 32'hc404aa7;
      26688: inst = 32'h8220000;
      26689: inst = 32'h10408000;
      26690: inst = 32'hc404aa8;
      26691: inst = 32'h8220000;
      26692: inst = 32'h10408000;
      26693: inst = 32'hc404aa9;
      26694: inst = 32'h8220000;
      26695: inst = 32'h10408000;
      26696: inst = 32'hc404aaa;
      26697: inst = 32'h8220000;
      26698: inst = 32'h10408000;
      26699: inst = 32'hc404aab;
      26700: inst = 32'h8220000;
      26701: inst = 32'h10408000;
      26702: inst = 32'hc404aac;
      26703: inst = 32'h8220000;
      26704: inst = 32'h10408000;
      26705: inst = 32'hc404aad;
      26706: inst = 32'h8220000;
      26707: inst = 32'h10408000;
      26708: inst = 32'hc404aae;
      26709: inst = 32'h8220000;
      26710: inst = 32'h10408000;
      26711: inst = 32'hc404aaf;
      26712: inst = 32'h8220000;
      26713: inst = 32'h10408000;
      26714: inst = 32'hc404ab0;
      26715: inst = 32'h8220000;
      26716: inst = 32'h10408000;
      26717: inst = 32'hc404ab1;
      26718: inst = 32'h8220000;
      26719: inst = 32'h10408000;
      26720: inst = 32'hc404ab2;
      26721: inst = 32'h8220000;
      26722: inst = 32'h10408000;
      26723: inst = 32'hc404ab3;
      26724: inst = 32'h8220000;
      26725: inst = 32'h10408000;
      26726: inst = 32'hc404ab4;
      26727: inst = 32'h8220000;
      26728: inst = 32'h10408000;
      26729: inst = 32'hc404ab5;
      26730: inst = 32'h8220000;
      26731: inst = 32'h10408000;
      26732: inst = 32'hc404ab6;
      26733: inst = 32'h8220000;
      26734: inst = 32'h10408000;
      26735: inst = 32'hc404ab7;
      26736: inst = 32'h8220000;
      26737: inst = 32'h10408000;
      26738: inst = 32'hc404ab8;
      26739: inst = 32'h8220000;
      26740: inst = 32'h10408000;
      26741: inst = 32'hc404ac7;
      26742: inst = 32'h8220000;
      26743: inst = 32'h10408000;
      26744: inst = 32'hc404ac8;
      26745: inst = 32'h8220000;
      26746: inst = 32'h10408000;
      26747: inst = 32'hc404ac9;
      26748: inst = 32'h8220000;
      26749: inst = 32'h10408000;
      26750: inst = 32'hc404aca;
      26751: inst = 32'h8220000;
      26752: inst = 32'h10408000;
      26753: inst = 32'hc404acb;
      26754: inst = 32'h8220000;
      26755: inst = 32'h10408000;
      26756: inst = 32'hc404acc;
      26757: inst = 32'h8220000;
      26758: inst = 32'h10408000;
      26759: inst = 32'hc404acd;
      26760: inst = 32'h8220000;
      26761: inst = 32'h10408000;
      26762: inst = 32'hc404ace;
      26763: inst = 32'h8220000;
      26764: inst = 32'h10408000;
      26765: inst = 32'hc404acf;
      26766: inst = 32'h8220000;
      26767: inst = 32'h10408000;
      26768: inst = 32'hc404ad0;
      26769: inst = 32'h8220000;
      26770: inst = 32'h10408000;
      26771: inst = 32'hc404ad1;
      26772: inst = 32'h8220000;
      26773: inst = 32'h10408000;
      26774: inst = 32'hc404ad2;
      26775: inst = 32'h8220000;
      26776: inst = 32'h10408000;
      26777: inst = 32'hc404ad3;
      26778: inst = 32'h8220000;
      26779: inst = 32'h10408000;
      26780: inst = 32'hc404ad4;
      26781: inst = 32'h8220000;
      26782: inst = 32'h10408000;
      26783: inst = 32'hc404ad5;
      26784: inst = 32'h8220000;
      26785: inst = 32'h10408000;
      26786: inst = 32'hc404ad6;
      26787: inst = 32'h8220000;
      26788: inst = 32'h10408000;
      26789: inst = 32'hc404ad7;
      26790: inst = 32'h8220000;
      26791: inst = 32'h10408000;
      26792: inst = 32'hc404ad8;
      26793: inst = 32'h8220000;
      26794: inst = 32'h10408000;
      26795: inst = 32'hc404ad9;
      26796: inst = 32'h8220000;
      26797: inst = 32'h10408000;
      26798: inst = 32'hc404ada;
      26799: inst = 32'h8220000;
      26800: inst = 32'h10408000;
      26801: inst = 32'hc404adb;
      26802: inst = 32'h8220000;
      26803: inst = 32'h10408000;
      26804: inst = 32'hc404adc;
      26805: inst = 32'h8220000;
      26806: inst = 32'h10408000;
      26807: inst = 32'hc404add;
      26808: inst = 32'h8220000;
      26809: inst = 32'h10408000;
      26810: inst = 32'hc404ade;
      26811: inst = 32'h8220000;
      26812: inst = 32'h10408000;
      26813: inst = 32'hc404adf;
      26814: inst = 32'h8220000;
      26815: inst = 32'h10408000;
      26816: inst = 32'hc404ae0;
      26817: inst = 32'h8220000;
      26818: inst = 32'h10408000;
      26819: inst = 32'hc404ae1;
      26820: inst = 32'h8220000;
      26821: inst = 32'h10408000;
      26822: inst = 32'hc404ae2;
      26823: inst = 32'h8220000;
      26824: inst = 32'h10408000;
      26825: inst = 32'hc404ae3;
      26826: inst = 32'h8220000;
      26827: inst = 32'h10408000;
      26828: inst = 32'hc404ae4;
      26829: inst = 32'h8220000;
      26830: inst = 32'h10408000;
      26831: inst = 32'hc404ae5;
      26832: inst = 32'h8220000;
      26833: inst = 32'h10408000;
      26834: inst = 32'hc404ae6;
      26835: inst = 32'h8220000;
      26836: inst = 32'h10408000;
      26837: inst = 32'hc404ae7;
      26838: inst = 32'h8220000;
      26839: inst = 32'h10408000;
      26840: inst = 32'hc404ae8;
      26841: inst = 32'h8220000;
      26842: inst = 32'h10408000;
      26843: inst = 32'hc404ae9;
      26844: inst = 32'h8220000;
      26845: inst = 32'h10408000;
      26846: inst = 32'hc404aea;
      26847: inst = 32'h8220000;
      26848: inst = 32'h10408000;
      26849: inst = 32'hc404aeb;
      26850: inst = 32'h8220000;
      26851: inst = 32'h10408000;
      26852: inst = 32'hc404aec;
      26853: inst = 32'h8220000;
      26854: inst = 32'h10408000;
      26855: inst = 32'hc404aed;
      26856: inst = 32'h8220000;
      26857: inst = 32'h10408000;
      26858: inst = 32'hc404aee;
      26859: inst = 32'h8220000;
      26860: inst = 32'h10408000;
      26861: inst = 32'hc404aef;
      26862: inst = 32'h8220000;
      26863: inst = 32'h10408000;
      26864: inst = 32'hc404af0;
      26865: inst = 32'h8220000;
      26866: inst = 32'h10408000;
      26867: inst = 32'hc404af1;
      26868: inst = 32'h8220000;
      26869: inst = 32'h10408000;
      26870: inst = 32'hc404af2;
      26871: inst = 32'h8220000;
      26872: inst = 32'h10408000;
      26873: inst = 32'hc404af3;
      26874: inst = 32'h8220000;
      26875: inst = 32'h10408000;
      26876: inst = 32'hc404af4;
      26877: inst = 32'h8220000;
      26878: inst = 32'h10408000;
      26879: inst = 32'hc404af5;
      26880: inst = 32'h8220000;
      26881: inst = 32'h10408000;
      26882: inst = 32'hc404af6;
      26883: inst = 32'h8220000;
      26884: inst = 32'h10408000;
      26885: inst = 32'hc404af7;
      26886: inst = 32'h8220000;
      26887: inst = 32'h10408000;
      26888: inst = 32'hc404af8;
      26889: inst = 32'h8220000;
      26890: inst = 32'h10408000;
      26891: inst = 32'hc404af9;
      26892: inst = 32'h8220000;
      26893: inst = 32'h10408000;
      26894: inst = 32'hc404afa;
      26895: inst = 32'h8220000;
      26896: inst = 32'h10408000;
      26897: inst = 32'hc404afb;
      26898: inst = 32'h8220000;
      26899: inst = 32'h10408000;
      26900: inst = 32'hc404afc;
      26901: inst = 32'h8220000;
      26902: inst = 32'h10408000;
      26903: inst = 32'hc404afd;
      26904: inst = 32'h8220000;
      26905: inst = 32'h10408000;
      26906: inst = 32'hc404afe;
      26907: inst = 32'h8220000;
      26908: inst = 32'h10408000;
      26909: inst = 32'hc404aff;
      26910: inst = 32'h8220000;
      26911: inst = 32'h10408000;
      26912: inst = 32'hc404b00;
      26913: inst = 32'h8220000;
      26914: inst = 32'h10408000;
      26915: inst = 32'hc404b01;
      26916: inst = 32'h8220000;
      26917: inst = 32'h10408000;
      26918: inst = 32'hc404b02;
      26919: inst = 32'h8220000;
      26920: inst = 32'h10408000;
      26921: inst = 32'hc404b03;
      26922: inst = 32'h8220000;
      26923: inst = 32'h10408000;
      26924: inst = 32'hc404b04;
      26925: inst = 32'h8220000;
      26926: inst = 32'h10408000;
      26927: inst = 32'hc404b05;
      26928: inst = 32'h8220000;
      26929: inst = 32'h10408000;
      26930: inst = 32'hc404b06;
      26931: inst = 32'h8220000;
      26932: inst = 32'h10408000;
      26933: inst = 32'hc404b07;
      26934: inst = 32'h8220000;
      26935: inst = 32'h10408000;
      26936: inst = 32'hc404b08;
      26937: inst = 32'h8220000;
      26938: inst = 32'h10408000;
      26939: inst = 32'hc404b09;
      26940: inst = 32'h8220000;
      26941: inst = 32'h10408000;
      26942: inst = 32'hc404b0a;
      26943: inst = 32'h8220000;
      26944: inst = 32'h10408000;
      26945: inst = 32'hc404b0b;
      26946: inst = 32'h8220000;
      26947: inst = 32'h10408000;
      26948: inst = 32'hc404b0c;
      26949: inst = 32'h8220000;
      26950: inst = 32'h10408000;
      26951: inst = 32'hc404b0d;
      26952: inst = 32'h8220000;
      26953: inst = 32'h10408000;
      26954: inst = 32'hc404b0e;
      26955: inst = 32'h8220000;
      26956: inst = 32'h10408000;
      26957: inst = 32'hc404b0f;
      26958: inst = 32'h8220000;
      26959: inst = 32'h10408000;
      26960: inst = 32'hc404b10;
      26961: inst = 32'h8220000;
      26962: inst = 32'h10408000;
      26963: inst = 32'hc404b11;
      26964: inst = 32'h8220000;
      26965: inst = 32'h10408000;
      26966: inst = 32'hc404b12;
      26967: inst = 32'h8220000;
      26968: inst = 32'h10408000;
      26969: inst = 32'hc404b13;
      26970: inst = 32'h8220000;
      26971: inst = 32'h10408000;
      26972: inst = 32'hc404b14;
      26973: inst = 32'h8220000;
      26974: inst = 32'h10408000;
      26975: inst = 32'hc404b15;
      26976: inst = 32'h8220000;
      26977: inst = 32'h10408000;
      26978: inst = 32'hc404b16;
      26979: inst = 32'h8220000;
      26980: inst = 32'h10408000;
      26981: inst = 32'hc404b17;
      26982: inst = 32'h8220000;
      26983: inst = 32'h10408000;
      26984: inst = 32'hc404b18;
      26985: inst = 32'h8220000;
      26986: inst = 32'h10408000;
      26987: inst = 32'hc404b27;
      26988: inst = 32'h8220000;
      26989: inst = 32'h10408000;
      26990: inst = 32'hc404b28;
      26991: inst = 32'h8220000;
      26992: inst = 32'h10408000;
      26993: inst = 32'hc404b29;
      26994: inst = 32'h8220000;
      26995: inst = 32'h10408000;
      26996: inst = 32'hc404b2a;
      26997: inst = 32'h8220000;
      26998: inst = 32'h10408000;
      26999: inst = 32'hc404b2b;
      27000: inst = 32'h8220000;
      27001: inst = 32'h10408000;
      27002: inst = 32'hc404b2c;
      27003: inst = 32'h8220000;
      27004: inst = 32'h10408000;
      27005: inst = 32'hc404b2d;
      27006: inst = 32'h8220000;
      27007: inst = 32'h10408000;
      27008: inst = 32'hc404b2e;
      27009: inst = 32'h8220000;
      27010: inst = 32'h10408000;
      27011: inst = 32'hc404b2f;
      27012: inst = 32'h8220000;
      27013: inst = 32'h10408000;
      27014: inst = 32'hc404b30;
      27015: inst = 32'h8220000;
      27016: inst = 32'h10408000;
      27017: inst = 32'hc404b31;
      27018: inst = 32'h8220000;
      27019: inst = 32'h10408000;
      27020: inst = 32'hc404b32;
      27021: inst = 32'h8220000;
      27022: inst = 32'h10408000;
      27023: inst = 32'hc404b33;
      27024: inst = 32'h8220000;
      27025: inst = 32'h10408000;
      27026: inst = 32'hc404b34;
      27027: inst = 32'h8220000;
      27028: inst = 32'h10408000;
      27029: inst = 32'hc404b35;
      27030: inst = 32'h8220000;
      27031: inst = 32'h10408000;
      27032: inst = 32'hc404b36;
      27033: inst = 32'h8220000;
      27034: inst = 32'h10408000;
      27035: inst = 32'hc404b37;
      27036: inst = 32'h8220000;
      27037: inst = 32'h10408000;
      27038: inst = 32'hc404b38;
      27039: inst = 32'h8220000;
      27040: inst = 32'h10408000;
      27041: inst = 32'hc404b39;
      27042: inst = 32'h8220000;
      27043: inst = 32'h10408000;
      27044: inst = 32'hc404b3a;
      27045: inst = 32'h8220000;
      27046: inst = 32'h10408000;
      27047: inst = 32'hc404b3b;
      27048: inst = 32'h8220000;
      27049: inst = 32'h10408000;
      27050: inst = 32'hc404b3c;
      27051: inst = 32'h8220000;
      27052: inst = 32'h10408000;
      27053: inst = 32'hc404b3d;
      27054: inst = 32'h8220000;
      27055: inst = 32'h10408000;
      27056: inst = 32'hc404b3e;
      27057: inst = 32'h8220000;
      27058: inst = 32'h10408000;
      27059: inst = 32'hc404b3f;
      27060: inst = 32'h8220000;
      27061: inst = 32'h10408000;
      27062: inst = 32'hc404b40;
      27063: inst = 32'h8220000;
      27064: inst = 32'h10408000;
      27065: inst = 32'hc404b41;
      27066: inst = 32'h8220000;
      27067: inst = 32'h10408000;
      27068: inst = 32'hc404b42;
      27069: inst = 32'h8220000;
      27070: inst = 32'h10408000;
      27071: inst = 32'hc404b43;
      27072: inst = 32'h8220000;
      27073: inst = 32'h10408000;
      27074: inst = 32'hc404b44;
      27075: inst = 32'h8220000;
      27076: inst = 32'h10408000;
      27077: inst = 32'hc404b45;
      27078: inst = 32'h8220000;
      27079: inst = 32'h10408000;
      27080: inst = 32'hc404b46;
      27081: inst = 32'h8220000;
      27082: inst = 32'h10408000;
      27083: inst = 32'hc404b47;
      27084: inst = 32'h8220000;
      27085: inst = 32'h10408000;
      27086: inst = 32'hc404b48;
      27087: inst = 32'h8220000;
      27088: inst = 32'h10408000;
      27089: inst = 32'hc404b49;
      27090: inst = 32'h8220000;
      27091: inst = 32'h10408000;
      27092: inst = 32'hc404b4a;
      27093: inst = 32'h8220000;
      27094: inst = 32'h10408000;
      27095: inst = 32'hc404b4b;
      27096: inst = 32'h8220000;
      27097: inst = 32'h10408000;
      27098: inst = 32'hc404b4c;
      27099: inst = 32'h8220000;
      27100: inst = 32'h10408000;
      27101: inst = 32'hc404b4d;
      27102: inst = 32'h8220000;
      27103: inst = 32'h10408000;
      27104: inst = 32'hc404b4e;
      27105: inst = 32'h8220000;
      27106: inst = 32'h10408000;
      27107: inst = 32'hc404b4f;
      27108: inst = 32'h8220000;
      27109: inst = 32'h10408000;
      27110: inst = 32'hc404b50;
      27111: inst = 32'h8220000;
      27112: inst = 32'h10408000;
      27113: inst = 32'hc404b51;
      27114: inst = 32'h8220000;
      27115: inst = 32'h10408000;
      27116: inst = 32'hc404b52;
      27117: inst = 32'h8220000;
      27118: inst = 32'h10408000;
      27119: inst = 32'hc404b53;
      27120: inst = 32'h8220000;
      27121: inst = 32'h10408000;
      27122: inst = 32'hc404b54;
      27123: inst = 32'h8220000;
      27124: inst = 32'h10408000;
      27125: inst = 32'hc404b55;
      27126: inst = 32'h8220000;
      27127: inst = 32'h10408000;
      27128: inst = 32'hc404b56;
      27129: inst = 32'h8220000;
      27130: inst = 32'h10408000;
      27131: inst = 32'hc404b57;
      27132: inst = 32'h8220000;
      27133: inst = 32'h10408000;
      27134: inst = 32'hc404b58;
      27135: inst = 32'h8220000;
      27136: inst = 32'h10408000;
      27137: inst = 32'hc404b59;
      27138: inst = 32'h8220000;
      27139: inst = 32'h10408000;
      27140: inst = 32'hc404b5a;
      27141: inst = 32'h8220000;
      27142: inst = 32'h10408000;
      27143: inst = 32'hc404b5b;
      27144: inst = 32'h8220000;
      27145: inst = 32'h10408000;
      27146: inst = 32'hc404b5c;
      27147: inst = 32'h8220000;
      27148: inst = 32'h10408000;
      27149: inst = 32'hc404b5d;
      27150: inst = 32'h8220000;
      27151: inst = 32'h10408000;
      27152: inst = 32'hc404b5e;
      27153: inst = 32'h8220000;
      27154: inst = 32'h10408000;
      27155: inst = 32'hc404b5f;
      27156: inst = 32'h8220000;
      27157: inst = 32'h10408000;
      27158: inst = 32'hc404b60;
      27159: inst = 32'h8220000;
      27160: inst = 32'h10408000;
      27161: inst = 32'hc404b61;
      27162: inst = 32'h8220000;
      27163: inst = 32'h10408000;
      27164: inst = 32'hc404b62;
      27165: inst = 32'h8220000;
      27166: inst = 32'h10408000;
      27167: inst = 32'hc404b63;
      27168: inst = 32'h8220000;
      27169: inst = 32'h10408000;
      27170: inst = 32'hc404b64;
      27171: inst = 32'h8220000;
      27172: inst = 32'h10408000;
      27173: inst = 32'hc404b65;
      27174: inst = 32'h8220000;
      27175: inst = 32'h10408000;
      27176: inst = 32'hc404b66;
      27177: inst = 32'h8220000;
      27178: inst = 32'h10408000;
      27179: inst = 32'hc404b67;
      27180: inst = 32'h8220000;
      27181: inst = 32'h10408000;
      27182: inst = 32'hc404b68;
      27183: inst = 32'h8220000;
      27184: inst = 32'h10408000;
      27185: inst = 32'hc404b69;
      27186: inst = 32'h8220000;
      27187: inst = 32'h10408000;
      27188: inst = 32'hc404b6a;
      27189: inst = 32'h8220000;
      27190: inst = 32'h10408000;
      27191: inst = 32'hc404b6b;
      27192: inst = 32'h8220000;
      27193: inst = 32'h10408000;
      27194: inst = 32'hc404b6c;
      27195: inst = 32'h8220000;
      27196: inst = 32'h10408000;
      27197: inst = 32'hc404b6d;
      27198: inst = 32'h8220000;
      27199: inst = 32'h10408000;
      27200: inst = 32'hc404b6e;
      27201: inst = 32'h8220000;
      27202: inst = 32'h10408000;
      27203: inst = 32'hc404b6f;
      27204: inst = 32'h8220000;
      27205: inst = 32'h10408000;
      27206: inst = 32'hc404b70;
      27207: inst = 32'h8220000;
      27208: inst = 32'h10408000;
      27209: inst = 32'hc404b71;
      27210: inst = 32'h8220000;
      27211: inst = 32'h10408000;
      27212: inst = 32'hc404b72;
      27213: inst = 32'h8220000;
      27214: inst = 32'h10408000;
      27215: inst = 32'hc404b73;
      27216: inst = 32'h8220000;
      27217: inst = 32'h10408000;
      27218: inst = 32'hc404b74;
      27219: inst = 32'h8220000;
      27220: inst = 32'h10408000;
      27221: inst = 32'hc404b75;
      27222: inst = 32'h8220000;
      27223: inst = 32'h10408000;
      27224: inst = 32'hc404b76;
      27225: inst = 32'h8220000;
      27226: inst = 32'h10408000;
      27227: inst = 32'hc404b77;
      27228: inst = 32'h8220000;
      27229: inst = 32'h10408000;
      27230: inst = 32'hc404b78;
      27231: inst = 32'h8220000;
      27232: inst = 32'h10408000;
      27233: inst = 32'hc404b87;
      27234: inst = 32'h8220000;
      27235: inst = 32'h10408000;
      27236: inst = 32'hc404b88;
      27237: inst = 32'h8220000;
      27238: inst = 32'h10408000;
      27239: inst = 32'hc404b89;
      27240: inst = 32'h8220000;
      27241: inst = 32'h10408000;
      27242: inst = 32'hc404b8a;
      27243: inst = 32'h8220000;
      27244: inst = 32'h10408000;
      27245: inst = 32'hc404b8b;
      27246: inst = 32'h8220000;
      27247: inst = 32'h10408000;
      27248: inst = 32'hc404b8c;
      27249: inst = 32'h8220000;
      27250: inst = 32'h10408000;
      27251: inst = 32'hc404b8d;
      27252: inst = 32'h8220000;
      27253: inst = 32'h10408000;
      27254: inst = 32'hc404b8e;
      27255: inst = 32'h8220000;
      27256: inst = 32'h10408000;
      27257: inst = 32'hc404b8f;
      27258: inst = 32'h8220000;
      27259: inst = 32'h10408000;
      27260: inst = 32'hc404b90;
      27261: inst = 32'h8220000;
      27262: inst = 32'h10408000;
      27263: inst = 32'hc404b91;
      27264: inst = 32'h8220000;
      27265: inst = 32'h10408000;
      27266: inst = 32'hc404b92;
      27267: inst = 32'h8220000;
      27268: inst = 32'h10408000;
      27269: inst = 32'hc404b93;
      27270: inst = 32'h8220000;
      27271: inst = 32'h10408000;
      27272: inst = 32'hc404b94;
      27273: inst = 32'h8220000;
      27274: inst = 32'h10408000;
      27275: inst = 32'hc404b95;
      27276: inst = 32'h8220000;
      27277: inst = 32'h10408000;
      27278: inst = 32'hc404b96;
      27279: inst = 32'h8220000;
      27280: inst = 32'h10408000;
      27281: inst = 32'hc404b97;
      27282: inst = 32'h8220000;
      27283: inst = 32'h10408000;
      27284: inst = 32'hc404b98;
      27285: inst = 32'h8220000;
      27286: inst = 32'h10408000;
      27287: inst = 32'hc404b99;
      27288: inst = 32'h8220000;
      27289: inst = 32'h10408000;
      27290: inst = 32'hc404b9a;
      27291: inst = 32'h8220000;
      27292: inst = 32'h10408000;
      27293: inst = 32'hc404b9b;
      27294: inst = 32'h8220000;
      27295: inst = 32'h10408000;
      27296: inst = 32'hc404b9c;
      27297: inst = 32'h8220000;
      27298: inst = 32'h10408000;
      27299: inst = 32'hc404b9d;
      27300: inst = 32'h8220000;
      27301: inst = 32'h10408000;
      27302: inst = 32'hc404b9e;
      27303: inst = 32'h8220000;
      27304: inst = 32'h10408000;
      27305: inst = 32'hc404b9f;
      27306: inst = 32'h8220000;
      27307: inst = 32'h10408000;
      27308: inst = 32'hc404ba0;
      27309: inst = 32'h8220000;
      27310: inst = 32'h10408000;
      27311: inst = 32'hc404ba1;
      27312: inst = 32'h8220000;
      27313: inst = 32'h10408000;
      27314: inst = 32'hc404ba2;
      27315: inst = 32'h8220000;
      27316: inst = 32'h10408000;
      27317: inst = 32'hc404ba3;
      27318: inst = 32'h8220000;
      27319: inst = 32'h10408000;
      27320: inst = 32'hc404ba4;
      27321: inst = 32'h8220000;
      27322: inst = 32'h10408000;
      27323: inst = 32'hc404ba5;
      27324: inst = 32'h8220000;
      27325: inst = 32'h10408000;
      27326: inst = 32'hc404ba6;
      27327: inst = 32'h8220000;
      27328: inst = 32'h10408000;
      27329: inst = 32'hc404ba7;
      27330: inst = 32'h8220000;
      27331: inst = 32'h10408000;
      27332: inst = 32'hc404ba8;
      27333: inst = 32'h8220000;
      27334: inst = 32'h10408000;
      27335: inst = 32'hc404ba9;
      27336: inst = 32'h8220000;
      27337: inst = 32'h10408000;
      27338: inst = 32'hc404baa;
      27339: inst = 32'h8220000;
      27340: inst = 32'h10408000;
      27341: inst = 32'hc404bab;
      27342: inst = 32'h8220000;
      27343: inst = 32'h10408000;
      27344: inst = 32'hc404bac;
      27345: inst = 32'h8220000;
      27346: inst = 32'h10408000;
      27347: inst = 32'hc404bad;
      27348: inst = 32'h8220000;
      27349: inst = 32'h10408000;
      27350: inst = 32'hc404bae;
      27351: inst = 32'h8220000;
      27352: inst = 32'h10408000;
      27353: inst = 32'hc404baf;
      27354: inst = 32'h8220000;
      27355: inst = 32'h10408000;
      27356: inst = 32'hc404bb0;
      27357: inst = 32'h8220000;
      27358: inst = 32'h10408000;
      27359: inst = 32'hc404bb1;
      27360: inst = 32'h8220000;
      27361: inst = 32'h10408000;
      27362: inst = 32'hc404bb2;
      27363: inst = 32'h8220000;
      27364: inst = 32'h10408000;
      27365: inst = 32'hc404bb3;
      27366: inst = 32'h8220000;
      27367: inst = 32'h10408000;
      27368: inst = 32'hc404bb4;
      27369: inst = 32'h8220000;
      27370: inst = 32'h10408000;
      27371: inst = 32'hc404bb5;
      27372: inst = 32'h8220000;
      27373: inst = 32'h10408000;
      27374: inst = 32'hc404bb6;
      27375: inst = 32'h8220000;
      27376: inst = 32'h10408000;
      27377: inst = 32'hc404bb7;
      27378: inst = 32'h8220000;
      27379: inst = 32'h10408000;
      27380: inst = 32'hc404bb8;
      27381: inst = 32'h8220000;
      27382: inst = 32'h10408000;
      27383: inst = 32'hc404bb9;
      27384: inst = 32'h8220000;
      27385: inst = 32'h10408000;
      27386: inst = 32'hc404bba;
      27387: inst = 32'h8220000;
      27388: inst = 32'h10408000;
      27389: inst = 32'hc404bbb;
      27390: inst = 32'h8220000;
      27391: inst = 32'h10408000;
      27392: inst = 32'hc404bbc;
      27393: inst = 32'h8220000;
      27394: inst = 32'h10408000;
      27395: inst = 32'hc404bbd;
      27396: inst = 32'h8220000;
      27397: inst = 32'h10408000;
      27398: inst = 32'hc404bbe;
      27399: inst = 32'h8220000;
      27400: inst = 32'h10408000;
      27401: inst = 32'hc404bbf;
      27402: inst = 32'h8220000;
      27403: inst = 32'h10408000;
      27404: inst = 32'hc404bc0;
      27405: inst = 32'h8220000;
      27406: inst = 32'h10408000;
      27407: inst = 32'hc404bc1;
      27408: inst = 32'h8220000;
      27409: inst = 32'h10408000;
      27410: inst = 32'hc404bc2;
      27411: inst = 32'h8220000;
      27412: inst = 32'h10408000;
      27413: inst = 32'hc404bc3;
      27414: inst = 32'h8220000;
      27415: inst = 32'h10408000;
      27416: inst = 32'hc404bc4;
      27417: inst = 32'h8220000;
      27418: inst = 32'h10408000;
      27419: inst = 32'hc404bc5;
      27420: inst = 32'h8220000;
      27421: inst = 32'h10408000;
      27422: inst = 32'hc404bc6;
      27423: inst = 32'h8220000;
      27424: inst = 32'h10408000;
      27425: inst = 32'hc404bc7;
      27426: inst = 32'h8220000;
      27427: inst = 32'h10408000;
      27428: inst = 32'hc404bc8;
      27429: inst = 32'h8220000;
      27430: inst = 32'h10408000;
      27431: inst = 32'hc404bc9;
      27432: inst = 32'h8220000;
      27433: inst = 32'h10408000;
      27434: inst = 32'hc404bca;
      27435: inst = 32'h8220000;
      27436: inst = 32'h10408000;
      27437: inst = 32'hc404bcb;
      27438: inst = 32'h8220000;
      27439: inst = 32'h10408000;
      27440: inst = 32'hc404bcc;
      27441: inst = 32'h8220000;
      27442: inst = 32'h10408000;
      27443: inst = 32'hc404bcd;
      27444: inst = 32'h8220000;
      27445: inst = 32'h10408000;
      27446: inst = 32'hc404bce;
      27447: inst = 32'h8220000;
      27448: inst = 32'h10408000;
      27449: inst = 32'hc404bcf;
      27450: inst = 32'h8220000;
      27451: inst = 32'h10408000;
      27452: inst = 32'hc404bd0;
      27453: inst = 32'h8220000;
      27454: inst = 32'h10408000;
      27455: inst = 32'hc404bd1;
      27456: inst = 32'h8220000;
      27457: inst = 32'h10408000;
      27458: inst = 32'hc404bd2;
      27459: inst = 32'h8220000;
      27460: inst = 32'h10408000;
      27461: inst = 32'hc404bd3;
      27462: inst = 32'h8220000;
      27463: inst = 32'h10408000;
      27464: inst = 32'hc404bd4;
      27465: inst = 32'h8220000;
      27466: inst = 32'h10408000;
      27467: inst = 32'hc404bd5;
      27468: inst = 32'h8220000;
      27469: inst = 32'h10408000;
      27470: inst = 32'hc404bd6;
      27471: inst = 32'h8220000;
      27472: inst = 32'h10408000;
      27473: inst = 32'hc404bd7;
      27474: inst = 32'h8220000;
      27475: inst = 32'h10408000;
      27476: inst = 32'hc404bd8;
      27477: inst = 32'h8220000;
      27478: inst = 32'h10408000;
      27479: inst = 32'hc404be7;
      27480: inst = 32'h8220000;
      27481: inst = 32'h10408000;
      27482: inst = 32'hc404be8;
      27483: inst = 32'h8220000;
      27484: inst = 32'h10408000;
      27485: inst = 32'hc404be9;
      27486: inst = 32'h8220000;
      27487: inst = 32'h10408000;
      27488: inst = 32'hc404bea;
      27489: inst = 32'h8220000;
      27490: inst = 32'h10408000;
      27491: inst = 32'hc404beb;
      27492: inst = 32'h8220000;
      27493: inst = 32'h10408000;
      27494: inst = 32'hc404bec;
      27495: inst = 32'h8220000;
      27496: inst = 32'h10408000;
      27497: inst = 32'hc404bed;
      27498: inst = 32'h8220000;
      27499: inst = 32'h10408000;
      27500: inst = 32'hc404bee;
      27501: inst = 32'h8220000;
      27502: inst = 32'h10408000;
      27503: inst = 32'hc404bef;
      27504: inst = 32'h8220000;
      27505: inst = 32'h10408000;
      27506: inst = 32'hc404bf0;
      27507: inst = 32'h8220000;
      27508: inst = 32'h10408000;
      27509: inst = 32'hc404bf1;
      27510: inst = 32'h8220000;
      27511: inst = 32'h10408000;
      27512: inst = 32'hc404bf2;
      27513: inst = 32'h8220000;
      27514: inst = 32'h10408000;
      27515: inst = 32'hc404bf3;
      27516: inst = 32'h8220000;
      27517: inst = 32'h10408000;
      27518: inst = 32'hc404bf4;
      27519: inst = 32'h8220000;
      27520: inst = 32'h10408000;
      27521: inst = 32'hc404bf5;
      27522: inst = 32'h8220000;
      27523: inst = 32'h10408000;
      27524: inst = 32'hc404bf6;
      27525: inst = 32'h8220000;
      27526: inst = 32'h10408000;
      27527: inst = 32'hc404bf7;
      27528: inst = 32'h8220000;
      27529: inst = 32'h10408000;
      27530: inst = 32'hc404bf8;
      27531: inst = 32'h8220000;
      27532: inst = 32'h10408000;
      27533: inst = 32'hc404bf9;
      27534: inst = 32'h8220000;
      27535: inst = 32'h10408000;
      27536: inst = 32'hc404bfa;
      27537: inst = 32'h8220000;
      27538: inst = 32'h10408000;
      27539: inst = 32'hc404bfb;
      27540: inst = 32'h8220000;
      27541: inst = 32'h10408000;
      27542: inst = 32'hc404bfc;
      27543: inst = 32'h8220000;
      27544: inst = 32'h10408000;
      27545: inst = 32'hc404bfd;
      27546: inst = 32'h8220000;
      27547: inst = 32'h10408000;
      27548: inst = 32'hc404bfe;
      27549: inst = 32'h8220000;
      27550: inst = 32'h10408000;
      27551: inst = 32'hc404bff;
      27552: inst = 32'h8220000;
      27553: inst = 32'h10408000;
      27554: inst = 32'hc404c00;
      27555: inst = 32'h8220000;
      27556: inst = 32'h10408000;
      27557: inst = 32'hc404c01;
      27558: inst = 32'h8220000;
      27559: inst = 32'h10408000;
      27560: inst = 32'hc404c02;
      27561: inst = 32'h8220000;
      27562: inst = 32'h10408000;
      27563: inst = 32'hc404c03;
      27564: inst = 32'h8220000;
      27565: inst = 32'h10408000;
      27566: inst = 32'hc404c04;
      27567: inst = 32'h8220000;
      27568: inst = 32'h10408000;
      27569: inst = 32'hc404c05;
      27570: inst = 32'h8220000;
      27571: inst = 32'h10408000;
      27572: inst = 32'hc404c06;
      27573: inst = 32'h8220000;
      27574: inst = 32'h10408000;
      27575: inst = 32'hc404c07;
      27576: inst = 32'h8220000;
      27577: inst = 32'h10408000;
      27578: inst = 32'hc404c08;
      27579: inst = 32'h8220000;
      27580: inst = 32'h10408000;
      27581: inst = 32'hc404c09;
      27582: inst = 32'h8220000;
      27583: inst = 32'h10408000;
      27584: inst = 32'hc404c0a;
      27585: inst = 32'h8220000;
      27586: inst = 32'h10408000;
      27587: inst = 32'hc404c0b;
      27588: inst = 32'h8220000;
      27589: inst = 32'h10408000;
      27590: inst = 32'hc404c0c;
      27591: inst = 32'h8220000;
      27592: inst = 32'h10408000;
      27593: inst = 32'hc404c0d;
      27594: inst = 32'h8220000;
      27595: inst = 32'h10408000;
      27596: inst = 32'hc404c0e;
      27597: inst = 32'h8220000;
      27598: inst = 32'h10408000;
      27599: inst = 32'hc404c0f;
      27600: inst = 32'h8220000;
      27601: inst = 32'h10408000;
      27602: inst = 32'hc404c10;
      27603: inst = 32'h8220000;
      27604: inst = 32'h10408000;
      27605: inst = 32'hc404c11;
      27606: inst = 32'h8220000;
      27607: inst = 32'h10408000;
      27608: inst = 32'hc404c12;
      27609: inst = 32'h8220000;
      27610: inst = 32'h10408000;
      27611: inst = 32'hc404c13;
      27612: inst = 32'h8220000;
      27613: inst = 32'h10408000;
      27614: inst = 32'hc404c14;
      27615: inst = 32'h8220000;
      27616: inst = 32'h10408000;
      27617: inst = 32'hc404c15;
      27618: inst = 32'h8220000;
      27619: inst = 32'h10408000;
      27620: inst = 32'hc404c16;
      27621: inst = 32'h8220000;
      27622: inst = 32'h10408000;
      27623: inst = 32'hc404c17;
      27624: inst = 32'h8220000;
      27625: inst = 32'h10408000;
      27626: inst = 32'hc404c18;
      27627: inst = 32'h8220000;
      27628: inst = 32'h10408000;
      27629: inst = 32'hc404c19;
      27630: inst = 32'h8220000;
      27631: inst = 32'h10408000;
      27632: inst = 32'hc404c1a;
      27633: inst = 32'h8220000;
      27634: inst = 32'h10408000;
      27635: inst = 32'hc404c1b;
      27636: inst = 32'h8220000;
      27637: inst = 32'h10408000;
      27638: inst = 32'hc404c1c;
      27639: inst = 32'h8220000;
      27640: inst = 32'h10408000;
      27641: inst = 32'hc404c1d;
      27642: inst = 32'h8220000;
      27643: inst = 32'h10408000;
      27644: inst = 32'hc404c1e;
      27645: inst = 32'h8220000;
      27646: inst = 32'h10408000;
      27647: inst = 32'hc404c1f;
      27648: inst = 32'h8220000;
      27649: inst = 32'h10408000;
      27650: inst = 32'hc404c20;
      27651: inst = 32'h8220000;
      27652: inst = 32'h10408000;
      27653: inst = 32'hc404c21;
      27654: inst = 32'h8220000;
      27655: inst = 32'h10408000;
      27656: inst = 32'hc404c22;
      27657: inst = 32'h8220000;
      27658: inst = 32'h10408000;
      27659: inst = 32'hc404c23;
      27660: inst = 32'h8220000;
      27661: inst = 32'h10408000;
      27662: inst = 32'hc404c24;
      27663: inst = 32'h8220000;
      27664: inst = 32'h10408000;
      27665: inst = 32'hc404c25;
      27666: inst = 32'h8220000;
      27667: inst = 32'h10408000;
      27668: inst = 32'hc404c26;
      27669: inst = 32'h8220000;
      27670: inst = 32'h10408000;
      27671: inst = 32'hc404c27;
      27672: inst = 32'h8220000;
      27673: inst = 32'h10408000;
      27674: inst = 32'hc404c28;
      27675: inst = 32'h8220000;
      27676: inst = 32'h10408000;
      27677: inst = 32'hc404c29;
      27678: inst = 32'h8220000;
      27679: inst = 32'h10408000;
      27680: inst = 32'hc404c2a;
      27681: inst = 32'h8220000;
      27682: inst = 32'h10408000;
      27683: inst = 32'hc404c2b;
      27684: inst = 32'h8220000;
      27685: inst = 32'h10408000;
      27686: inst = 32'hc404c2c;
      27687: inst = 32'h8220000;
      27688: inst = 32'h10408000;
      27689: inst = 32'hc404c2d;
      27690: inst = 32'h8220000;
      27691: inst = 32'h10408000;
      27692: inst = 32'hc404c2e;
      27693: inst = 32'h8220000;
      27694: inst = 32'h10408000;
      27695: inst = 32'hc404c2f;
      27696: inst = 32'h8220000;
      27697: inst = 32'h10408000;
      27698: inst = 32'hc404c30;
      27699: inst = 32'h8220000;
      27700: inst = 32'h10408000;
      27701: inst = 32'hc404c31;
      27702: inst = 32'h8220000;
      27703: inst = 32'h10408000;
      27704: inst = 32'hc404c32;
      27705: inst = 32'h8220000;
      27706: inst = 32'h10408000;
      27707: inst = 32'hc404c33;
      27708: inst = 32'h8220000;
      27709: inst = 32'h10408000;
      27710: inst = 32'hc404c34;
      27711: inst = 32'h8220000;
      27712: inst = 32'h10408000;
      27713: inst = 32'hc404c35;
      27714: inst = 32'h8220000;
      27715: inst = 32'h10408000;
      27716: inst = 32'hc404c36;
      27717: inst = 32'h8220000;
      27718: inst = 32'h10408000;
      27719: inst = 32'hc404c37;
      27720: inst = 32'h8220000;
      27721: inst = 32'h10408000;
      27722: inst = 32'hc404c38;
      27723: inst = 32'h8220000;
      27724: inst = 32'h10408000;
      27725: inst = 32'hc404c47;
      27726: inst = 32'h8220000;
      27727: inst = 32'h10408000;
      27728: inst = 32'hc404c48;
      27729: inst = 32'h8220000;
      27730: inst = 32'h10408000;
      27731: inst = 32'hc404c49;
      27732: inst = 32'h8220000;
      27733: inst = 32'h10408000;
      27734: inst = 32'hc404c4a;
      27735: inst = 32'h8220000;
      27736: inst = 32'h10408000;
      27737: inst = 32'hc404c4b;
      27738: inst = 32'h8220000;
      27739: inst = 32'h10408000;
      27740: inst = 32'hc404c4c;
      27741: inst = 32'h8220000;
      27742: inst = 32'h10408000;
      27743: inst = 32'hc404c4d;
      27744: inst = 32'h8220000;
      27745: inst = 32'h10408000;
      27746: inst = 32'hc404c4e;
      27747: inst = 32'h8220000;
      27748: inst = 32'h10408000;
      27749: inst = 32'hc404c4f;
      27750: inst = 32'h8220000;
      27751: inst = 32'h10408000;
      27752: inst = 32'hc404c50;
      27753: inst = 32'h8220000;
      27754: inst = 32'h10408000;
      27755: inst = 32'hc404c51;
      27756: inst = 32'h8220000;
      27757: inst = 32'h10408000;
      27758: inst = 32'hc404c52;
      27759: inst = 32'h8220000;
      27760: inst = 32'h10408000;
      27761: inst = 32'hc404c53;
      27762: inst = 32'h8220000;
      27763: inst = 32'h10408000;
      27764: inst = 32'hc404c54;
      27765: inst = 32'h8220000;
      27766: inst = 32'h10408000;
      27767: inst = 32'hc404c55;
      27768: inst = 32'h8220000;
      27769: inst = 32'h10408000;
      27770: inst = 32'hc404c56;
      27771: inst = 32'h8220000;
      27772: inst = 32'h10408000;
      27773: inst = 32'hc404c57;
      27774: inst = 32'h8220000;
      27775: inst = 32'h10408000;
      27776: inst = 32'hc404c58;
      27777: inst = 32'h8220000;
      27778: inst = 32'h10408000;
      27779: inst = 32'hc404c59;
      27780: inst = 32'h8220000;
      27781: inst = 32'h10408000;
      27782: inst = 32'hc404c5a;
      27783: inst = 32'h8220000;
      27784: inst = 32'h10408000;
      27785: inst = 32'hc404c5b;
      27786: inst = 32'h8220000;
      27787: inst = 32'h10408000;
      27788: inst = 32'hc404c5c;
      27789: inst = 32'h8220000;
      27790: inst = 32'h10408000;
      27791: inst = 32'hc404c5d;
      27792: inst = 32'h8220000;
      27793: inst = 32'h10408000;
      27794: inst = 32'hc404c5e;
      27795: inst = 32'h8220000;
      27796: inst = 32'h10408000;
      27797: inst = 32'hc404c5f;
      27798: inst = 32'h8220000;
      27799: inst = 32'h10408000;
      27800: inst = 32'hc404c60;
      27801: inst = 32'h8220000;
      27802: inst = 32'h10408000;
      27803: inst = 32'hc404c61;
      27804: inst = 32'h8220000;
      27805: inst = 32'h10408000;
      27806: inst = 32'hc404c62;
      27807: inst = 32'h8220000;
      27808: inst = 32'h10408000;
      27809: inst = 32'hc404c63;
      27810: inst = 32'h8220000;
      27811: inst = 32'h10408000;
      27812: inst = 32'hc404c64;
      27813: inst = 32'h8220000;
      27814: inst = 32'h10408000;
      27815: inst = 32'hc404c65;
      27816: inst = 32'h8220000;
      27817: inst = 32'h10408000;
      27818: inst = 32'hc404c66;
      27819: inst = 32'h8220000;
      27820: inst = 32'h10408000;
      27821: inst = 32'hc404c67;
      27822: inst = 32'h8220000;
      27823: inst = 32'h10408000;
      27824: inst = 32'hc404c68;
      27825: inst = 32'h8220000;
      27826: inst = 32'h10408000;
      27827: inst = 32'hc404c69;
      27828: inst = 32'h8220000;
      27829: inst = 32'h10408000;
      27830: inst = 32'hc404c6a;
      27831: inst = 32'h8220000;
      27832: inst = 32'h10408000;
      27833: inst = 32'hc404c6b;
      27834: inst = 32'h8220000;
      27835: inst = 32'h10408000;
      27836: inst = 32'hc404c6c;
      27837: inst = 32'h8220000;
      27838: inst = 32'h10408000;
      27839: inst = 32'hc404c6d;
      27840: inst = 32'h8220000;
      27841: inst = 32'h10408000;
      27842: inst = 32'hc404c6e;
      27843: inst = 32'h8220000;
      27844: inst = 32'h10408000;
      27845: inst = 32'hc404c6f;
      27846: inst = 32'h8220000;
      27847: inst = 32'h10408000;
      27848: inst = 32'hc404c70;
      27849: inst = 32'h8220000;
      27850: inst = 32'h10408000;
      27851: inst = 32'hc404c71;
      27852: inst = 32'h8220000;
      27853: inst = 32'h10408000;
      27854: inst = 32'hc404c72;
      27855: inst = 32'h8220000;
      27856: inst = 32'h10408000;
      27857: inst = 32'hc404c73;
      27858: inst = 32'h8220000;
      27859: inst = 32'h10408000;
      27860: inst = 32'hc404c74;
      27861: inst = 32'h8220000;
      27862: inst = 32'h10408000;
      27863: inst = 32'hc404c75;
      27864: inst = 32'h8220000;
      27865: inst = 32'h10408000;
      27866: inst = 32'hc404c76;
      27867: inst = 32'h8220000;
      27868: inst = 32'h10408000;
      27869: inst = 32'hc404c77;
      27870: inst = 32'h8220000;
      27871: inst = 32'h10408000;
      27872: inst = 32'hc404c78;
      27873: inst = 32'h8220000;
      27874: inst = 32'h10408000;
      27875: inst = 32'hc404c79;
      27876: inst = 32'h8220000;
      27877: inst = 32'h10408000;
      27878: inst = 32'hc404c7a;
      27879: inst = 32'h8220000;
      27880: inst = 32'h10408000;
      27881: inst = 32'hc404c7b;
      27882: inst = 32'h8220000;
      27883: inst = 32'h10408000;
      27884: inst = 32'hc404c7c;
      27885: inst = 32'h8220000;
      27886: inst = 32'h10408000;
      27887: inst = 32'hc404c7d;
      27888: inst = 32'h8220000;
      27889: inst = 32'h10408000;
      27890: inst = 32'hc404c7e;
      27891: inst = 32'h8220000;
      27892: inst = 32'h10408000;
      27893: inst = 32'hc404c7f;
      27894: inst = 32'h8220000;
      27895: inst = 32'h10408000;
      27896: inst = 32'hc404c80;
      27897: inst = 32'h8220000;
      27898: inst = 32'h10408000;
      27899: inst = 32'hc404c81;
      27900: inst = 32'h8220000;
      27901: inst = 32'h10408000;
      27902: inst = 32'hc404c82;
      27903: inst = 32'h8220000;
      27904: inst = 32'h10408000;
      27905: inst = 32'hc404c83;
      27906: inst = 32'h8220000;
      27907: inst = 32'h10408000;
      27908: inst = 32'hc404c84;
      27909: inst = 32'h8220000;
      27910: inst = 32'h10408000;
      27911: inst = 32'hc404c85;
      27912: inst = 32'h8220000;
      27913: inst = 32'h10408000;
      27914: inst = 32'hc404c86;
      27915: inst = 32'h8220000;
      27916: inst = 32'h10408000;
      27917: inst = 32'hc404c87;
      27918: inst = 32'h8220000;
      27919: inst = 32'h10408000;
      27920: inst = 32'hc404c88;
      27921: inst = 32'h8220000;
      27922: inst = 32'h10408000;
      27923: inst = 32'hc404c89;
      27924: inst = 32'h8220000;
      27925: inst = 32'h10408000;
      27926: inst = 32'hc404c8a;
      27927: inst = 32'h8220000;
      27928: inst = 32'h10408000;
      27929: inst = 32'hc404c8b;
      27930: inst = 32'h8220000;
      27931: inst = 32'h10408000;
      27932: inst = 32'hc404c8c;
      27933: inst = 32'h8220000;
      27934: inst = 32'h10408000;
      27935: inst = 32'hc404c8d;
      27936: inst = 32'h8220000;
      27937: inst = 32'h10408000;
      27938: inst = 32'hc404c8e;
      27939: inst = 32'h8220000;
      27940: inst = 32'h10408000;
      27941: inst = 32'hc404c8f;
      27942: inst = 32'h8220000;
      27943: inst = 32'h10408000;
      27944: inst = 32'hc404c90;
      27945: inst = 32'h8220000;
      27946: inst = 32'h10408000;
      27947: inst = 32'hc404c91;
      27948: inst = 32'h8220000;
      27949: inst = 32'h10408000;
      27950: inst = 32'hc404c92;
      27951: inst = 32'h8220000;
      27952: inst = 32'h10408000;
      27953: inst = 32'hc404c93;
      27954: inst = 32'h8220000;
      27955: inst = 32'h10408000;
      27956: inst = 32'hc404c94;
      27957: inst = 32'h8220000;
      27958: inst = 32'h10408000;
      27959: inst = 32'hc404c95;
      27960: inst = 32'h8220000;
      27961: inst = 32'h10408000;
      27962: inst = 32'hc404c96;
      27963: inst = 32'h8220000;
      27964: inst = 32'h10408000;
      27965: inst = 32'hc404c97;
      27966: inst = 32'h8220000;
      27967: inst = 32'h10408000;
      27968: inst = 32'hc404c98;
      27969: inst = 32'h8220000;
      27970: inst = 32'h10408000;
      27971: inst = 32'hc404ca7;
      27972: inst = 32'h8220000;
      27973: inst = 32'h10408000;
      27974: inst = 32'hc404ca8;
      27975: inst = 32'h8220000;
      27976: inst = 32'h10408000;
      27977: inst = 32'hc404ca9;
      27978: inst = 32'h8220000;
      27979: inst = 32'h10408000;
      27980: inst = 32'hc404caa;
      27981: inst = 32'h8220000;
      27982: inst = 32'h10408000;
      27983: inst = 32'hc404cab;
      27984: inst = 32'h8220000;
      27985: inst = 32'h10408000;
      27986: inst = 32'hc404cac;
      27987: inst = 32'h8220000;
      27988: inst = 32'h10408000;
      27989: inst = 32'hc404cad;
      27990: inst = 32'h8220000;
      27991: inst = 32'h10408000;
      27992: inst = 32'hc404cae;
      27993: inst = 32'h8220000;
      27994: inst = 32'h10408000;
      27995: inst = 32'hc404cb2;
      27996: inst = 32'h8220000;
      27997: inst = 32'h10408000;
      27998: inst = 32'hc404cb3;
      27999: inst = 32'h8220000;
      28000: inst = 32'h10408000;
      28001: inst = 32'hc404cb4;
      28002: inst = 32'h8220000;
      28003: inst = 32'h10408000;
      28004: inst = 32'hc404cb5;
      28005: inst = 32'h8220000;
      28006: inst = 32'h10408000;
      28007: inst = 32'hc404cb6;
      28008: inst = 32'h8220000;
      28009: inst = 32'h10408000;
      28010: inst = 32'hc404cb7;
      28011: inst = 32'h8220000;
      28012: inst = 32'h10408000;
      28013: inst = 32'hc404cb8;
      28014: inst = 32'h8220000;
      28015: inst = 32'h10408000;
      28016: inst = 32'hc404cb9;
      28017: inst = 32'h8220000;
      28018: inst = 32'h10408000;
      28019: inst = 32'hc404cba;
      28020: inst = 32'h8220000;
      28021: inst = 32'h10408000;
      28022: inst = 32'hc404cbb;
      28023: inst = 32'h8220000;
      28024: inst = 32'h10408000;
      28025: inst = 32'hc404cbc;
      28026: inst = 32'h8220000;
      28027: inst = 32'h10408000;
      28028: inst = 32'hc404cbd;
      28029: inst = 32'h8220000;
      28030: inst = 32'h10408000;
      28031: inst = 32'hc404cbe;
      28032: inst = 32'h8220000;
      28033: inst = 32'h10408000;
      28034: inst = 32'hc404cbf;
      28035: inst = 32'h8220000;
      28036: inst = 32'h10408000;
      28037: inst = 32'hc404cc0;
      28038: inst = 32'h8220000;
      28039: inst = 32'h10408000;
      28040: inst = 32'hc404cc1;
      28041: inst = 32'h8220000;
      28042: inst = 32'h10408000;
      28043: inst = 32'hc404cc2;
      28044: inst = 32'h8220000;
      28045: inst = 32'h10408000;
      28046: inst = 32'hc404cc3;
      28047: inst = 32'h8220000;
      28048: inst = 32'h10408000;
      28049: inst = 32'hc404cc4;
      28050: inst = 32'h8220000;
      28051: inst = 32'h10408000;
      28052: inst = 32'hc404cc5;
      28053: inst = 32'h8220000;
      28054: inst = 32'h10408000;
      28055: inst = 32'hc404cc6;
      28056: inst = 32'h8220000;
      28057: inst = 32'h10408000;
      28058: inst = 32'hc404cc7;
      28059: inst = 32'h8220000;
      28060: inst = 32'h10408000;
      28061: inst = 32'hc404cc8;
      28062: inst = 32'h8220000;
      28063: inst = 32'h10408000;
      28064: inst = 32'hc404cc9;
      28065: inst = 32'h8220000;
      28066: inst = 32'h10408000;
      28067: inst = 32'hc404cca;
      28068: inst = 32'h8220000;
      28069: inst = 32'h10408000;
      28070: inst = 32'hc404ccb;
      28071: inst = 32'h8220000;
      28072: inst = 32'h10408000;
      28073: inst = 32'hc404ccc;
      28074: inst = 32'h8220000;
      28075: inst = 32'h10408000;
      28076: inst = 32'hc404ccd;
      28077: inst = 32'h8220000;
      28078: inst = 32'h10408000;
      28079: inst = 32'hc404cce;
      28080: inst = 32'h8220000;
      28081: inst = 32'h10408000;
      28082: inst = 32'hc404ccf;
      28083: inst = 32'h8220000;
      28084: inst = 32'h10408000;
      28085: inst = 32'hc404cd0;
      28086: inst = 32'h8220000;
      28087: inst = 32'h10408000;
      28088: inst = 32'hc404cd1;
      28089: inst = 32'h8220000;
      28090: inst = 32'h10408000;
      28091: inst = 32'hc404cd2;
      28092: inst = 32'h8220000;
      28093: inst = 32'h10408000;
      28094: inst = 32'hc404cd3;
      28095: inst = 32'h8220000;
      28096: inst = 32'h10408000;
      28097: inst = 32'hc404cd4;
      28098: inst = 32'h8220000;
      28099: inst = 32'h10408000;
      28100: inst = 32'hc404cd5;
      28101: inst = 32'h8220000;
      28102: inst = 32'h10408000;
      28103: inst = 32'hc404cd6;
      28104: inst = 32'h8220000;
      28105: inst = 32'h10408000;
      28106: inst = 32'hc404cd7;
      28107: inst = 32'h8220000;
      28108: inst = 32'h10408000;
      28109: inst = 32'hc404cd8;
      28110: inst = 32'h8220000;
      28111: inst = 32'h10408000;
      28112: inst = 32'hc404cd9;
      28113: inst = 32'h8220000;
      28114: inst = 32'h10408000;
      28115: inst = 32'hc404cda;
      28116: inst = 32'h8220000;
      28117: inst = 32'h10408000;
      28118: inst = 32'hc404cdb;
      28119: inst = 32'h8220000;
      28120: inst = 32'h10408000;
      28121: inst = 32'hc404cdc;
      28122: inst = 32'h8220000;
      28123: inst = 32'h10408000;
      28124: inst = 32'hc404cdd;
      28125: inst = 32'h8220000;
      28126: inst = 32'h10408000;
      28127: inst = 32'hc404cde;
      28128: inst = 32'h8220000;
      28129: inst = 32'h10408000;
      28130: inst = 32'hc404cdf;
      28131: inst = 32'h8220000;
      28132: inst = 32'h10408000;
      28133: inst = 32'hc404ce0;
      28134: inst = 32'h8220000;
      28135: inst = 32'h10408000;
      28136: inst = 32'hc404ce1;
      28137: inst = 32'h8220000;
      28138: inst = 32'h10408000;
      28139: inst = 32'hc404ce2;
      28140: inst = 32'h8220000;
      28141: inst = 32'h10408000;
      28142: inst = 32'hc404ce3;
      28143: inst = 32'h8220000;
      28144: inst = 32'h10408000;
      28145: inst = 32'hc404ce4;
      28146: inst = 32'h8220000;
      28147: inst = 32'h10408000;
      28148: inst = 32'hc404ce5;
      28149: inst = 32'h8220000;
      28150: inst = 32'h10408000;
      28151: inst = 32'hc404ce6;
      28152: inst = 32'h8220000;
      28153: inst = 32'h10408000;
      28154: inst = 32'hc404ce7;
      28155: inst = 32'h8220000;
      28156: inst = 32'h10408000;
      28157: inst = 32'hc404ce8;
      28158: inst = 32'h8220000;
      28159: inst = 32'h10408000;
      28160: inst = 32'hc404ce9;
      28161: inst = 32'h8220000;
      28162: inst = 32'h10408000;
      28163: inst = 32'hc404cea;
      28164: inst = 32'h8220000;
      28165: inst = 32'h10408000;
      28166: inst = 32'hc404ceb;
      28167: inst = 32'h8220000;
      28168: inst = 32'h10408000;
      28169: inst = 32'hc404cec;
      28170: inst = 32'h8220000;
      28171: inst = 32'h10408000;
      28172: inst = 32'hc404ced;
      28173: inst = 32'h8220000;
      28174: inst = 32'h10408000;
      28175: inst = 32'hc404cee;
      28176: inst = 32'h8220000;
      28177: inst = 32'h10408000;
      28178: inst = 32'hc404cef;
      28179: inst = 32'h8220000;
      28180: inst = 32'h10408000;
      28181: inst = 32'hc404cf3;
      28182: inst = 32'h8220000;
      28183: inst = 32'h10408000;
      28184: inst = 32'hc404cf4;
      28185: inst = 32'h8220000;
      28186: inst = 32'h10408000;
      28187: inst = 32'hc404cf5;
      28188: inst = 32'h8220000;
      28189: inst = 32'h10408000;
      28190: inst = 32'hc404cf6;
      28191: inst = 32'h8220000;
      28192: inst = 32'h10408000;
      28193: inst = 32'hc404cf7;
      28194: inst = 32'h8220000;
      28195: inst = 32'h10408000;
      28196: inst = 32'hc404cf8;
      28197: inst = 32'h8220000;
      28198: inst = 32'h10408000;
      28199: inst = 32'hc404d07;
      28200: inst = 32'h8220000;
      28201: inst = 32'h10408000;
      28202: inst = 32'hc404d08;
      28203: inst = 32'h8220000;
      28204: inst = 32'h10408000;
      28205: inst = 32'hc404d09;
      28206: inst = 32'h8220000;
      28207: inst = 32'h10408000;
      28208: inst = 32'hc404d0a;
      28209: inst = 32'h8220000;
      28210: inst = 32'h10408000;
      28211: inst = 32'hc404d0b;
      28212: inst = 32'h8220000;
      28213: inst = 32'h10408000;
      28214: inst = 32'hc404d0c;
      28215: inst = 32'h8220000;
      28216: inst = 32'h10408000;
      28217: inst = 32'hc404d0d;
      28218: inst = 32'h8220000;
      28219: inst = 32'h10408000;
      28220: inst = 32'hc404d0e;
      28221: inst = 32'h8220000;
      28222: inst = 32'h10408000;
      28223: inst = 32'hc404d12;
      28224: inst = 32'h8220000;
      28225: inst = 32'h10408000;
      28226: inst = 32'hc404d13;
      28227: inst = 32'h8220000;
      28228: inst = 32'h10408000;
      28229: inst = 32'hc404d14;
      28230: inst = 32'h8220000;
      28231: inst = 32'h10408000;
      28232: inst = 32'hc404d15;
      28233: inst = 32'h8220000;
      28234: inst = 32'h10408000;
      28235: inst = 32'hc404d16;
      28236: inst = 32'h8220000;
      28237: inst = 32'h10408000;
      28238: inst = 32'hc404d17;
      28239: inst = 32'h8220000;
      28240: inst = 32'h10408000;
      28241: inst = 32'hc404d18;
      28242: inst = 32'h8220000;
      28243: inst = 32'h10408000;
      28244: inst = 32'hc404d19;
      28245: inst = 32'h8220000;
      28246: inst = 32'h10408000;
      28247: inst = 32'hc404d1a;
      28248: inst = 32'h8220000;
      28249: inst = 32'h10408000;
      28250: inst = 32'hc404d1b;
      28251: inst = 32'h8220000;
      28252: inst = 32'h10408000;
      28253: inst = 32'hc404d1c;
      28254: inst = 32'h8220000;
      28255: inst = 32'h10408000;
      28256: inst = 32'hc404d1d;
      28257: inst = 32'h8220000;
      28258: inst = 32'h10408000;
      28259: inst = 32'hc404d1e;
      28260: inst = 32'h8220000;
      28261: inst = 32'h10408000;
      28262: inst = 32'hc404d1f;
      28263: inst = 32'h8220000;
      28264: inst = 32'h10408000;
      28265: inst = 32'hc404d20;
      28266: inst = 32'h8220000;
      28267: inst = 32'h10408000;
      28268: inst = 32'hc404d22;
      28269: inst = 32'h8220000;
      28270: inst = 32'h10408000;
      28271: inst = 32'hc404d23;
      28272: inst = 32'h8220000;
      28273: inst = 32'h10408000;
      28274: inst = 32'hc404d24;
      28275: inst = 32'h8220000;
      28276: inst = 32'h10408000;
      28277: inst = 32'hc404d25;
      28278: inst = 32'h8220000;
      28279: inst = 32'h10408000;
      28280: inst = 32'hc404d26;
      28281: inst = 32'h8220000;
      28282: inst = 32'h10408000;
      28283: inst = 32'hc404d27;
      28284: inst = 32'h8220000;
      28285: inst = 32'h10408000;
      28286: inst = 32'hc404d28;
      28287: inst = 32'h8220000;
      28288: inst = 32'h10408000;
      28289: inst = 32'hc404d29;
      28290: inst = 32'h8220000;
      28291: inst = 32'h10408000;
      28292: inst = 32'hc404d2a;
      28293: inst = 32'h8220000;
      28294: inst = 32'h10408000;
      28295: inst = 32'hc404d2c;
      28296: inst = 32'h8220000;
      28297: inst = 32'h10408000;
      28298: inst = 32'hc404d2d;
      28299: inst = 32'h8220000;
      28300: inst = 32'h10408000;
      28301: inst = 32'hc404d2e;
      28302: inst = 32'h8220000;
      28303: inst = 32'h10408000;
      28304: inst = 32'hc404d2f;
      28305: inst = 32'h8220000;
      28306: inst = 32'h10408000;
      28307: inst = 32'hc404d30;
      28308: inst = 32'h8220000;
      28309: inst = 32'h10408000;
      28310: inst = 32'hc404d31;
      28311: inst = 32'h8220000;
      28312: inst = 32'h10408000;
      28313: inst = 32'hc404d32;
      28314: inst = 32'h8220000;
      28315: inst = 32'h10408000;
      28316: inst = 32'hc404d33;
      28317: inst = 32'h8220000;
      28318: inst = 32'h10408000;
      28319: inst = 32'hc404d34;
      28320: inst = 32'h8220000;
      28321: inst = 32'h10408000;
      28322: inst = 32'hc404d35;
      28323: inst = 32'h8220000;
      28324: inst = 32'h10408000;
      28325: inst = 32'hc404d36;
      28326: inst = 32'h8220000;
      28327: inst = 32'h10408000;
      28328: inst = 32'hc404d37;
      28329: inst = 32'h8220000;
      28330: inst = 32'h10408000;
      28331: inst = 32'hc404d38;
      28332: inst = 32'h8220000;
      28333: inst = 32'h10408000;
      28334: inst = 32'hc404d39;
      28335: inst = 32'h8220000;
      28336: inst = 32'h10408000;
      28337: inst = 32'hc404d3a;
      28338: inst = 32'h8220000;
      28339: inst = 32'h10408000;
      28340: inst = 32'hc404d3b;
      28341: inst = 32'h8220000;
      28342: inst = 32'h10408000;
      28343: inst = 32'hc404d3c;
      28344: inst = 32'h8220000;
      28345: inst = 32'h10408000;
      28346: inst = 32'hc404d3d;
      28347: inst = 32'h8220000;
      28348: inst = 32'h10408000;
      28349: inst = 32'hc404d3e;
      28350: inst = 32'h8220000;
      28351: inst = 32'h10408000;
      28352: inst = 32'hc404d40;
      28353: inst = 32'h8220000;
      28354: inst = 32'h10408000;
      28355: inst = 32'hc404d41;
      28356: inst = 32'h8220000;
      28357: inst = 32'h10408000;
      28358: inst = 32'hc404d42;
      28359: inst = 32'h8220000;
      28360: inst = 32'h10408000;
      28361: inst = 32'hc404d43;
      28362: inst = 32'h8220000;
      28363: inst = 32'h10408000;
      28364: inst = 32'hc404d45;
      28365: inst = 32'h8220000;
      28366: inst = 32'h10408000;
      28367: inst = 32'hc404d46;
      28368: inst = 32'h8220000;
      28369: inst = 32'h10408000;
      28370: inst = 32'hc404d47;
      28371: inst = 32'h8220000;
      28372: inst = 32'h10408000;
      28373: inst = 32'hc404d48;
      28374: inst = 32'h8220000;
      28375: inst = 32'h10408000;
      28376: inst = 32'hc404d49;
      28377: inst = 32'h8220000;
      28378: inst = 32'h10408000;
      28379: inst = 32'hc404d4a;
      28380: inst = 32'h8220000;
      28381: inst = 32'h10408000;
      28382: inst = 32'hc404d4b;
      28383: inst = 32'h8220000;
      28384: inst = 32'h10408000;
      28385: inst = 32'hc404d4c;
      28386: inst = 32'h8220000;
      28387: inst = 32'h10408000;
      28388: inst = 32'hc404d4d;
      28389: inst = 32'h8220000;
      28390: inst = 32'h10408000;
      28391: inst = 32'hc404d4e;
      28392: inst = 32'h8220000;
      28393: inst = 32'h10408000;
      28394: inst = 32'hc404d4f;
      28395: inst = 32'h8220000;
      28396: inst = 32'h10408000;
      28397: inst = 32'hc404d53;
      28398: inst = 32'h8220000;
      28399: inst = 32'h10408000;
      28400: inst = 32'hc404d54;
      28401: inst = 32'h8220000;
      28402: inst = 32'h10408000;
      28403: inst = 32'hc404d55;
      28404: inst = 32'h8220000;
      28405: inst = 32'h10408000;
      28406: inst = 32'hc404d56;
      28407: inst = 32'h8220000;
      28408: inst = 32'h10408000;
      28409: inst = 32'hc404d57;
      28410: inst = 32'h8220000;
      28411: inst = 32'h10408000;
      28412: inst = 32'hc404d58;
      28413: inst = 32'h8220000;
      28414: inst = 32'h10408000;
      28415: inst = 32'hc404d67;
      28416: inst = 32'h8220000;
      28417: inst = 32'h10408000;
      28418: inst = 32'hc404d68;
      28419: inst = 32'h8220000;
      28420: inst = 32'h10408000;
      28421: inst = 32'hc404d69;
      28422: inst = 32'h8220000;
      28423: inst = 32'h10408000;
      28424: inst = 32'hc404d6a;
      28425: inst = 32'h8220000;
      28426: inst = 32'h10408000;
      28427: inst = 32'hc404d6b;
      28428: inst = 32'h8220000;
      28429: inst = 32'h10408000;
      28430: inst = 32'hc404d6c;
      28431: inst = 32'h8220000;
      28432: inst = 32'h10408000;
      28433: inst = 32'hc404d6d;
      28434: inst = 32'h8220000;
      28435: inst = 32'h10408000;
      28436: inst = 32'hc404d6e;
      28437: inst = 32'h8220000;
      28438: inst = 32'h10408000;
      28439: inst = 32'hc404d6f;
      28440: inst = 32'h8220000;
      28441: inst = 32'h10408000;
      28442: inst = 32'hc404d72;
      28443: inst = 32'h8220000;
      28444: inst = 32'h10408000;
      28445: inst = 32'hc404d73;
      28446: inst = 32'h8220000;
      28447: inst = 32'h10408000;
      28448: inst = 32'hc404d74;
      28449: inst = 32'h8220000;
      28450: inst = 32'h10408000;
      28451: inst = 32'hc404d75;
      28452: inst = 32'h8220000;
      28453: inst = 32'h10408000;
      28454: inst = 32'hc404d76;
      28455: inst = 32'h8220000;
      28456: inst = 32'h10408000;
      28457: inst = 32'hc404d77;
      28458: inst = 32'h8220000;
      28459: inst = 32'h10408000;
      28460: inst = 32'hc404d78;
      28461: inst = 32'h8220000;
      28462: inst = 32'h10408000;
      28463: inst = 32'hc404d79;
      28464: inst = 32'h8220000;
      28465: inst = 32'h10408000;
      28466: inst = 32'hc404d7a;
      28467: inst = 32'h8220000;
      28468: inst = 32'h10408000;
      28469: inst = 32'hc404d7b;
      28470: inst = 32'h8220000;
      28471: inst = 32'h10408000;
      28472: inst = 32'hc404d7c;
      28473: inst = 32'h8220000;
      28474: inst = 32'h10408000;
      28475: inst = 32'hc404d7d;
      28476: inst = 32'h8220000;
      28477: inst = 32'h10408000;
      28478: inst = 32'hc404d7e;
      28479: inst = 32'h8220000;
      28480: inst = 32'h10408000;
      28481: inst = 32'hc404d7f;
      28482: inst = 32'h8220000;
      28483: inst = 32'h10408000;
      28484: inst = 32'hc404d82;
      28485: inst = 32'h8220000;
      28486: inst = 32'h10408000;
      28487: inst = 32'hc404d83;
      28488: inst = 32'h8220000;
      28489: inst = 32'h10408000;
      28490: inst = 32'hc404d84;
      28491: inst = 32'h8220000;
      28492: inst = 32'h10408000;
      28493: inst = 32'hc404d85;
      28494: inst = 32'h8220000;
      28495: inst = 32'h10408000;
      28496: inst = 32'hc404d86;
      28497: inst = 32'h8220000;
      28498: inst = 32'h10408000;
      28499: inst = 32'hc404d87;
      28500: inst = 32'h8220000;
      28501: inst = 32'h10408000;
      28502: inst = 32'hc404d88;
      28503: inst = 32'h8220000;
      28504: inst = 32'h10408000;
      28505: inst = 32'hc404d89;
      28506: inst = 32'h8220000;
      28507: inst = 32'h10408000;
      28508: inst = 32'hc404d8c;
      28509: inst = 32'h8220000;
      28510: inst = 32'h10408000;
      28511: inst = 32'hc404d8d;
      28512: inst = 32'h8220000;
      28513: inst = 32'h10408000;
      28514: inst = 32'hc404d8e;
      28515: inst = 32'h8220000;
      28516: inst = 32'h10408000;
      28517: inst = 32'hc404d8f;
      28518: inst = 32'h8220000;
      28519: inst = 32'h10408000;
      28520: inst = 32'hc404d90;
      28521: inst = 32'h8220000;
      28522: inst = 32'h10408000;
      28523: inst = 32'hc404d91;
      28524: inst = 32'h8220000;
      28525: inst = 32'h10408000;
      28526: inst = 32'hc404d92;
      28527: inst = 32'h8220000;
      28528: inst = 32'h10408000;
      28529: inst = 32'hc404d93;
      28530: inst = 32'h8220000;
      28531: inst = 32'h10408000;
      28532: inst = 32'hc404d94;
      28533: inst = 32'h8220000;
      28534: inst = 32'h10408000;
      28535: inst = 32'hc404d95;
      28536: inst = 32'h8220000;
      28537: inst = 32'h10408000;
      28538: inst = 32'hc404d96;
      28539: inst = 32'h8220000;
      28540: inst = 32'h10408000;
      28541: inst = 32'hc404d97;
      28542: inst = 32'h8220000;
      28543: inst = 32'h10408000;
      28544: inst = 32'hc404d98;
      28545: inst = 32'h8220000;
      28546: inst = 32'h10408000;
      28547: inst = 32'hc404d99;
      28548: inst = 32'h8220000;
      28549: inst = 32'h10408000;
      28550: inst = 32'hc404d9a;
      28551: inst = 32'h8220000;
      28552: inst = 32'h10408000;
      28553: inst = 32'hc404d9b;
      28554: inst = 32'h8220000;
      28555: inst = 32'h10408000;
      28556: inst = 32'hc404d9c;
      28557: inst = 32'h8220000;
      28558: inst = 32'h10408000;
      28559: inst = 32'hc404d9d;
      28560: inst = 32'h8220000;
      28561: inst = 32'h10408000;
      28562: inst = 32'hc404da0;
      28563: inst = 32'h8220000;
      28564: inst = 32'h10408000;
      28565: inst = 32'hc404da1;
      28566: inst = 32'h8220000;
      28567: inst = 32'h10408000;
      28568: inst = 32'hc404da2;
      28569: inst = 32'h8220000;
      28570: inst = 32'h10408000;
      28571: inst = 32'hc404da5;
      28572: inst = 32'h8220000;
      28573: inst = 32'h10408000;
      28574: inst = 32'hc404da6;
      28575: inst = 32'h8220000;
      28576: inst = 32'h10408000;
      28577: inst = 32'hc404da7;
      28578: inst = 32'h8220000;
      28579: inst = 32'h10408000;
      28580: inst = 32'hc404da8;
      28581: inst = 32'h8220000;
      28582: inst = 32'h10408000;
      28583: inst = 32'hc404da9;
      28584: inst = 32'h8220000;
      28585: inst = 32'h10408000;
      28586: inst = 32'hc404daa;
      28587: inst = 32'h8220000;
      28588: inst = 32'h10408000;
      28589: inst = 32'hc404dab;
      28590: inst = 32'h8220000;
      28591: inst = 32'h10408000;
      28592: inst = 32'hc404dac;
      28593: inst = 32'h8220000;
      28594: inst = 32'h10408000;
      28595: inst = 32'hc404dad;
      28596: inst = 32'h8220000;
      28597: inst = 32'h10408000;
      28598: inst = 32'hc404dae;
      28599: inst = 32'h8220000;
      28600: inst = 32'h10408000;
      28601: inst = 32'hc404daf;
      28602: inst = 32'h8220000;
      28603: inst = 32'h10408000;
      28604: inst = 32'hc404db0;
      28605: inst = 32'h8220000;
      28606: inst = 32'h10408000;
      28607: inst = 32'hc404db3;
      28608: inst = 32'h8220000;
      28609: inst = 32'h10408000;
      28610: inst = 32'hc404db4;
      28611: inst = 32'h8220000;
      28612: inst = 32'h10408000;
      28613: inst = 32'hc404db5;
      28614: inst = 32'h8220000;
      28615: inst = 32'h10408000;
      28616: inst = 32'hc404db6;
      28617: inst = 32'h8220000;
      28618: inst = 32'h10408000;
      28619: inst = 32'hc404db7;
      28620: inst = 32'h8220000;
      28621: inst = 32'h10408000;
      28622: inst = 32'hc404db8;
      28623: inst = 32'h8220000;
      28624: inst = 32'h10408000;
      28625: inst = 32'hc404dc7;
      28626: inst = 32'h8220000;
      28627: inst = 32'h10408000;
      28628: inst = 32'hc404dc8;
      28629: inst = 32'h8220000;
      28630: inst = 32'h10408000;
      28631: inst = 32'hc404dc9;
      28632: inst = 32'h8220000;
      28633: inst = 32'h10408000;
      28634: inst = 32'hc404dca;
      28635: inst = 32'h8220000;
      28636: inst = 32'h10408000;
      28637: inst = 32'hc404dcb;
      28638: inst = 32'h8220000;
      28639: inst = 32'h10408000;
      28640: inst = 32'hc404dd4;
      28641: inst = 32'h8220000;
      28642: inst = 32'h10408000;
      28643: inst = 32'hc404dd5;
      28644: inst = 32'h8220000;
      28645: inst = 32'h10408000;
      28646: inst = 32'hc404dd9;
      28647: inst = 32'h8220000;
      28648: inst = 32'h10408000;
      28649: inst = 32'hc404ddc;
      28650: inst = 32'h8220000;
      28651: inst = 32'h10408000;
      28652: inst = 32'hc404de3;
      28653: inst = 32'h8220000;
      28654: inst = 32'h10408000;
      28655: inst = 32'hc404de4;
      28656: inst = 32'h8220000;
      28657: inst = 32'h10408000;
      28658: inst = 32'hc404de5;
      28659: inst = 32'h8220000;
      28660: inst = 32'h10408000;
      28661: inst = 32'hc404de6;
      28662: inst = 32'h8220000;
      28663: inst = 32'h10408000;
      28664: inst = 32'hc404de7;
      28665: inst = 32'h8220000;
      28666: inst = 32'h10408000;
      28667: inst = 32'hc404de8;
      28668: inst = 32'h8220000;
      28669: inst = 32'h10408000;
      28670: inst = 32'hc404ded;
      28671: inst = 32'h8220000;
      28672: inst = 32'h10408000;
      28673: inst = 32'hc404dee;
      28674: inst = 32'h8220000;
      28675: inst = 32'h10408000;
      28676: inst = 32'hc404df2;
      28677: inst = 32'h8220000;
      28678: inst = 32'h10408000;
      28679: inst = 32'hc404df3;
      28680: inst = 32'h8220000;
      28681: inst = 32'h10408000;
      28682: inst = 32'hc404df4;
      28683: inst = 32'h8220000;
      28684: inst = 32'h10408000;
      28685: inst = 32'hc404df5;
      28686: inst = 32'h8220000;
      28687: inst = 32'h10408000;
      28688: inst = 32'hc404df6;
      28689: inst = 32'h8220000;
      28690: inst = 32'h10408000;
      28691: inst = 32'hc404df7;
      28692: inst = 32'h8220000;
      28693: inst = 32'h10408000;
      28694: inst = 32'hc404df8;
      28695: inst = 32'h8220000;
      28696: inst = 32'h10408000;
      28697: inst = 32'hc404dfc;
      28698: inst = 32'h8220000;
      28699: inst = 32'h10408000;
      28700: inst = 32'hc404e01;
      28701: inst = 32'h8220000;
      28702: inst = 32'h10408000;
      28703: inst = 32'hc404e06;
      28704: inst = 32'h8220000;
      28705: inst = 32'h10408000;
      28706: inst = 32'hc404e07;
      28707: inst = 32'h8220000;
      28708: inst = 32'h10408000;
      28709: inst = 32'hc404e0b;
      28710: inst = 32'h8220000;
      28711: inst = 32'h10408000;
      28712: inst = 32'hc404e0c;
      28713: inst = 32'h8220000;
      28714: inst = 32'h10408000;
      28715: inst = 32'hc404e0d;
      28716: inst = 32'h8220000;
      28717: inst = 32'h10408000;
      28718: inst = 32'hc404e10;
      28719: inst = 32'h8220000;
      28720: inst = 32'h10408000;
      28721: inst = 32'hc404e13;
      28722: inst = 32'h8220000;
      28723: inst = 32'h10408000;
      28724: inst = 32'hc404e16;
      28725: inst = 32'h8220000;
      28726: inst = 32'h10408000;
      28727: inst = 32'hc404e17;
      28728: inst = 32'h8220000;
      28729: inst = 32'h10408000;
      28730: inst = 32'hc404e18;
      28731: inst = 32'h8220000;
      28732: inst = 32'h10408000;
      28733: inst = 32'hc404e27;
      28734: inst = 32'h8220000;
      28735: inst = 32'h10408000;
      28736: inst = 32'hc404e28;
      28737: inst = 32'h8220000;
      28738: inst = 32'h10408000;
      28739: inst = 32'hc404e29;
      28740: inst = 32'h8220000;
      28741: inst = 32'h10408000;
      28742: inst = 32'hc404e2a;
      28743: inst = 32'h8220000;
      28744: inst = 32'h10408000;
      28745: inst = 32'hc404e3c;
      28746: inst = 32'h8220000;
      28747: inst = 32'h10408000;
      28748: inst = 32'hc404e44;
      28749: inst = 32'h8220000;
      28750: inst = 32'h10408000;
      28751: inst = 32'hc404e45;
      28752: inst = 32'h8220000;
      28753: inst = 32'h10408000;
      28754: inst = 32'hc404e46;
      28755: inst = 32'h8220000;
      28756: inst = 32'h10408000;
      28757: inst = 32'hc404e47;
      28758: inst = 32'h8220000;
      28759: inst = 32'h10408000;
      28760: inst = 32'hc404e48;
      28761: inst = 32'h8220000;
      28762: inst = 32'h10408000;
      28763: inst = 32'hc404e53;
      28764: inst = 32'h8220000;
      28765: inst = 32'h10408000;
      28766: inst = 32'hc404e54;
      28767: inst = 32'h8220000;
      28768: inst = 32'h10408000;
      28769: inst = 32'hc404e55;
      28770: inst = 32'h8220000;
      28771: inst = 32'h10408000;
      28772: inst = 32'hc404e56;
      28773: inst = 32'h8220000;
      28774: inst = 32'h10408000;
      28775: inst = 32'hc404e57;
      28776: inst = 32'h8220000;
      28777: inst = 32'h10408000;
      28778: inst = 32'hc404e76;
      28779: inst = 32'h8220000;
      28780: inst = 32'h10408000;
      28781: inst = 32'hc404e77;
      28782: inst = 32'h8220000;
      28783: inst = 32'h10408000;
      28784: inst = 32'hc404e78;
      28785: inst = 32'h8220000;
      28786: inst = 32'h10408000;
      28787: inst = 32'hc404e87;
      28788: inst = 32'h8220000;
      28789: inst = 32'h10408000;
      28790: inst = 32'hc404e88;
      28791: inst = 32'h8220000;
      28792: inst = 32'h10408000;
      28793: inst = 32'hc404e89;
      28794: inst = 32'h8220000;
      28795: inst = 32'h10408000;
      28796: inst = 32'hc404e8a;
      28797: inst = 32'h8220000;
      28798: inst = 32'h10408000;
      28799: inst = 32'hc404e8d;
      28800: inst = 32'h8220000;
      28801: inst = 32'h10408000;
      28802: inst = 32'hc404e8e;
      28803: inst = 32'h8220000;
      28804: inst = 32'h10408000;
      28805: inst = 32'hc404e92;
      28806: inst = 32'h8220000;
      28807: inst = 32'h10408000;
      28808: inst = 32'hc404e97;
      28809: inst = 32'h8220000;
      28810: inst = 32'h10408000;
      28811: inst = 32'hc404e9c;
      28812: inst = 32'h8220000;
      28813: inst = 32'h10408000;
      28814: inst = 32'hc404e9f;
      28815: inst = 32'h8220000;
      28816: inst = 32'h10408000;
      28817: inst = 32'hc404ea2;
      28818: inst = 32'h8220000;
      28819: inst = 32'h10408000;
      28820: inst = 32'hc404ea3;
      28821: inst = 32'h8220000;
      28822: inst = 32'h10408000;
      28823: inst = 32'hc404ea4;
      28824: inst = 32'h8220000;
      28825: inst = 32'h10408000;
      28826: inst = 32'hc404ea5;
      28827: inst = 32'h8220000;
      28828: inst = 32'h10408000;
      28829: inst = 32'hc404ea6;
      28830: inst = 32'h8220000;
      28831: inst = 32'h10408000;
      28832: inst = 32'hc404ea7;
      28833: inst = 32'h8220000;
      28834: inst = 32'h10408000;
      28835: inst = 32'hc404ea8;
      28836: inst = 32'h8220000;
      28837: inst = 32'h10408000;
      28838: inst = 32'hc404ea9;
      28839: inst = 32'h8220000;
      28840: inst = 32'h10408000;
      28841: inst = 32'hc404eac;
      28842: inst = 32'h8220000;
      28843: inst = 32'h10408000;
      28844: inst = 32'hc404ead;
      28845: inst = 32'h8220000;
      28846: inst = 32'h10408000;
      28847: inst = 32'hc404eb0;
      28848: inst = 32'h8220000;
      28849: inst = 32'h10408000;
      28850: inst = 32'hc404eb3;
      28851: inst = 32'h8220000;
      28852: inst = 32'h10408000;
      28853: inst = 32'hc404eb4;
      28854: inst = 32'h8220000;
      28855: inst = 32'h10408000;
      28856: inst = 32'hc404eb5;
      28857: inst = 32'h8220000;
      28858: inst = 32'h10408000;
      28859: inst = 32'hc404eb6;
      28860: inst = 32'h8220000;
      28861: inst = 32'h10408000;
      28862: inst = 32'hc404eb7;
      28863: inst = 32'h8220000;
      28864: inst = 32'h10408000;
      28865: inst = 32'hc404eba;
      28866: inst = 32'h8220000;
      28867: inst = 32'h10408000;
      28868: inst = 32'hc404ebd;
      28869: inst = 32'h8220000;
      28870: inst = 32'h10408000;
      28871: inst = 32'hc404ec0;
      28872: inst = 32'h8220000;
      28873: inst = 32'h10408000;
      28874: inst = 32'hc404ec1;
      28875: inst = 32'h8220000;
      28876: inst = 32'h10408000;
      28877: inst = 32'hc404ec2;
      28878: inst = 32'h8220000;
      28879: inst = 32'h10408000;
      28880: inst = 32'hc404ec5;
      28881: inst = 32'h8220000;
      28882: inst = 32'h10408000;
      28883: inst = 32'hc404ec6;
      28884: inst = 32'h8220000;
      28885: inst = 32'h10408000;
      28886: inst = 32'hc404ec9;
      28887: inst = 32'h8220000;
      28888: inst = 32'h10408000;
      28889: inst = 32'hc404ece;
      28890: inst = 32'h8220000;
      28891: inst = 32'h10408000;
      28892: inst = 32'hc404ed5;
      28893: inst = 32'h8220000;
      28894: inst = 32'h10408000;
      28895: inst = 32'hc404ed6;
      28896: inst = 32'h8220000;
      28897: inst = 32'h10408000;
      28898: inst = 32'hc404ed7;
      28899: inst = 32'h8220000;
      28900: inst = 32'h10408000;
      28901: inst = 32'hc404ed8;
      28902: inst = 32'h8220000;
      28903: inst = 32'h10408000;
      28904: inst = 32'hc404ee7;
      28905: inst = 32'h8220000;
      28906: inst = 32'h10408000;
      28907: inst = 32'hc404ee8;
      28908: inst = 32'h8220000;
      28909: inst = 32'h10408000;
      28910: inst = 32'hc404ee9;
      28911: inst = 32'h8220000;
      28912: inst = 32'h10408000;
      28913: inst = 32'hc404eea;
      28914: inst = 32'h8220000;
      28915: inst = 32'h10408000;
      28916: inst = 32'hc404eef;
      28917: inst = 32'h8220000;
      28918: inst = 32'h10408000;
      28919: inst = 32'hc404ef2;
      28920: inst = 32'h8220000;
      28921: inst = 32'h10408000;
      28922: inst = 32'hc404ef6;
      28923: inst = 32'h8220000;
      28924: inst = 32'h10408000;
      28925: inst = 32'hc404ef7;
      28926: inst = 32'h8220000;
      28927: inst = 32'h10408000;
      28928: inst = 32'hc404ef8;
      28929: inst = 32'h8220000;
      28930: inst = 32'h10408000;
      28931: inst = 32'hc404efc;
      28932: inst = 32'h8220000;
      28933: inst = 32'h10408000;
      28934: inst = 32'hc404eff;
      28935: inst = 32'h8220000;
      28936: inst = 32'h10408000;
      28937: inst = 32'hc404f02;
      28938: inst = 32'h8220000;
      28939: inst = 32'h10408000;
      28940: inst = 32'hc404f03;
      28941: inst = 32'h8220000;
      28942: inst = 32'h10408000;
      28943: inst = 32'hc404f04;
      28944: inst = 32'h8220000;
      28945: inst = 32'h10408000;
      28946: inst = 32'hc404f05;
      28947: inst = 32'h8220000;
      28948: inst = 32'h10408000;
      28949: inst = 32'hc404f06;
      28950: inst = 32'h8220000;
      28951: inst = 32'h10408000;
      28952: inst = 32'hc404f07;
      28953: inst = 32'h8220000;
      28954: inst = 32'h10408000;
      28955: inst = 32'hc404f08;
      28956: inst = 32'h8220000;
      28957: inst = 32'h10408000;
      28958: inst = 32'hc404f09;
      28959: inst = 32'h8220000;
      28960: inst = 32'h10408000;
      28961: inst = 32'hc404f0c;
      28962: inst = 32'h8220000;
      28963: inst = 32'h10408000;
      28964: inst = 32'hc404f0f;
      28965: inst = 32'h8220000;
      28966: inst = 32'h10408000;
      28967: inst = 32'hc404f10;
      28968: inst = 32'h8220000;
      28969: inst = 32'h10408000;
      28970: inst = 32'hc404f11;
      28971: inst = 32'h8220000;
      28972: inst = 32'h10408000;
      28973: inst = 32'hc404f14;
      28974: inst = 32'h8220000;
      28975: inst = 32'h10408000;
      28976: inst = 32'hc404f15;
      28977: inst = 32'h8220000;
      28978: inst = 32'h10408000;
      28979: inst = 32'hc404f16;
      28980: inst = 32'h8220000;
      28981: inst = 32'h10408000;
      28982: inst = 32'hc404f17;
      28983: inst = 32'h8220000;
      28984: inst = 32'h10408000;
      28985: inst = 32'hc404f1d;
      28986: inst = 32'h8220000;
      28987: inst = 32'h10408000;
      28988: inst = 32'hc404f20;
      28989: inst = 32'h8220000;
      28990: inst = 32'h10408000;
      28991: inst = 32'hc404f21;
      28992: inst = 32'h8220000;
      28993: inst = 32'h10408000;
      28994: inst = 32'hc404f22;
      28995: inst = 32'h8220000;
      28996: inst = 32'h10408000;
      28997: inst = 32'hc404f25;
      28998: inst = 32'h8220000;
      28999: inst = 32'h10408000;
      29000: inst = 32'hc404f26;
      29001: inst = 32'h8220000;
      29002: inst = 32'h10408000;
      29003: inst = 32'hc404f2e;
      29004: inst = 32'h8220000;
      29005: inst = 32'h10408000;
      29006: inst = 32'hc404f2f;
      29007: inst = 32'h8220000;
      29008: inst = 32'h10408000;
      29009: inst = 32'hc404f30;
      29010: inst = 32'h8220000;
      29011: inst = 32'h10408000;
      29012: inst = 32'hc404f35;
      29013: inst = 32'h8220000;
      29014: inst = 32'h10408000;
      29015: inst = 32'hc404f36;
      29016: inst = 32'h8220000;
      29017: inst = 32'h10408000;
      29018: inst = 32'hc404f37;
      29019: inst = 32'h8220000;
      29020: inst = 32'h10408000;
      29021: inst = 32'hc404f38;
      29022: inst = 32'h8220000;
      29023: inst = 32'h10408000;
      29024: inst = 32'hc404f47;
      29025: inst = 32'h8220000;
      29026: inst = 32'h10408000;
      29027: inst = 32'hc404f48;
      29028: inst = 32'h8220000;
      29029: inst = 32'h10408000;
      29030: inst = 32'hc404f49;
      29031: inst = 32'h8220000;
      29032: inst = 32'h10408000;
      29033: inst = 32'hc404f4a;
      29034: inst = 32'h8220000;
      29035: inst = 32'h10408000;
      29036: inst = 32'hc404f4b;
      29037: inst = 32'h8220000;
      29038: inst = 32'h10408000;
      29039: inst = 32'hc404f4c;
      29040: inst = 32'h8220000;
      29041: inst = 32'h10408000;
      29042: inst = 32'hc404f52;
      29043: inst = 32'h8220000;
      29044: inst = 32'h10408000;
      29045: inst = 32'hc404f56;
      29046: inst = 32'h8220000;
      29047: inst = 32'h10408000;
      29048: inst = 32'hc404f57;
      29049: inst = 32'h8220000;
      29050: inst = 32'h10408000;
      29051: inst = 32'hc404f58;
      29052: inst = 32'h8220000;
      29053: inst = 32'h10408000;
      29054: inst = 32'hc404f5c;
      29055: inst = 32'h8220000;
      29056: inst = 32'h10408000;
      29057: inst = 32'hc404f5f;
      29058: inst = 32'h8220000;
      29059: inst = 32'h10408000;
      29060: inst = 32'hc404f62;
      29061: inst = 32'h8220000;
      29062: inst = 32'h10408000;
      29063: inst = 32'hc404f63;
      29064: inst = 32'h8220000;
      29065: inst = 32'h10408000;
      29066: inst = 32'hc404f64;
      29067: inst = 32'h8220000;
      29068: inst = 32'h10408000;
      29069: inst = 32'hc404f65;
      29070: inst = 32'h8220000;
      29071: inst = 32'h10408000;
      29072: inst = 32'hc404f66;
      29073: inst = 32'h8220000;
      29074: inst = 32'h10408000;
      29075: inst = 32'hc404f67;
      29076: inst = 32'h8220000;
      29077: inst = 32'h10408000;
      29078: inst = 32'hc404f68;
      29079: inst = 32'h8220000;
      29080: inst = 32'h10408000;
      29081: inst = 32'hc404f69;
      29082: inst = 32'h8220000;
      29083: inst = 32'h10408000;
      29084: inst = 32'hc404f6c;
      29085: inst = 32'h8220000;
      29086: inst = 32'h10408000;
      29087: inst = 32'hc404f6f;
      29088: inst = 32'h8220000;
      29089: inst = 32'h10408000;
      29090: inst = 32'hc404f70;
      29091: inst = 32'h8220000;
      29092: inst = 32'h10408000;
      29093: inst = 32'hc404f71;
      29094: inst = 32'h8220000;
      29095: inst = 32'h10408000;
      29096: inst = 32'hc404f74;
      29097: inst = 32'h8220000;
      29098: inst = 32'h10408000;
      29099: inst = 32'hc404f75;
      29100: inst = 32'h8220000;
      29101: inst = 32'h10408000;
      29102: inst = 32'hc404f76;
      29103: inst = 32'h8220000;
      29104: inst = 32'h10408000;
      29105: inst = 32'hc404f77;
      29106: inst = 32'h8220000;
      29107: inst = 32'h10408000;
      29108: inst = 32'hc404f7a;
      29109: inst = 32'h8220000;
      29110: inst = 32'h10408000;
      29111: inst = 32'hc404f7d;
      29112: inst = 32'h8220000;
      29113: inst = 32'h10408000;
      29114: inst = 32'hc404f80;
      29115: inst = 32'h8220000;
      29116: inst = 32'h10408000;
      29117: inst = 32'hc404f81;
      29118: inst = 32'h8220000;
      29119: inst = 32'h10408000;
      29120: inst = 32'hc404f82;
      29121: inst = 32'h8220000;
      29122: inst = 32'h10408000;
      29123: inst = 32'hc404f85;
      29124: inst = 32'h8220000;
      29125: inst = 32'h10408000;
      29126: inst = 32'hc404f86;
      29127: inst = 32'h8220000;
      29128: inst = 32'h10408000;
      29129: inst = 32'hc404f89;
      29130: inst = 32'h8220000;
      29131: inst = 32'h10408000;
      29132: inst = 32'hc404f8e;
      29133: inst = 32'h8220000;
      29134: inst = 32'h10408000;
      29135: inst = 32'hc404f8f;
      29136: inst = 32'h8220000;
      29137: inst = 32'h10408000;
      29138: inst = 32'hc404f90;
      29139: inst = 32'h8220000;
      29140: inst = 32'h10408000;
      29141: inst = 32'hc404f95;
      29142: inst = 32'h8220000;
      29143: inst = 32'h10408000;
      29144: inst = 32'hc404f96;
      29145: inst = 32'h8220000;
      29146: inst = 32'h10408000;
      29147: inst = 32'hc404f97;
      29148: inst = 32'h8220000;
      29149: inst = 32'h10408000;
      29150: inst = 32'hc404f98;
      29151: inst = 32'h8220000;
      29152: inst = 32'h10408000;
      29153: inst = 32'hc404fa7;
      29154: inst = 32'h8220000;
      29155: inst = 32'h10408000;
      29156: inst = 32'hc404fa8;
      29157: inst = 32'h8220000;
      29158: inst = 32'h10408000;
      29159: inst = 32'hc404fa9;
      29160: inst = 32'h8220000;
      29161: inst = 32'h10408000;
      29162: inst = 32'hc404faa;
      29163: inst = 32'h8220000;
      29164: inst = 32'h10408000;
      29165: inst = 32'hc404fad;
      29166: inst = 32'h8220000;
      29167: inst = 32'h10408000;
      29168: inst = 32'hc404fae;
      29169: inst = 32'h8220000;
      29170: inst = 32'h10408000;
      29171: inst = 32'hc404fb2;
      29172: inst = 32'h8220000;
      29173: inst = 32'h10408000;
      29174: inst = 32'hc404fb7;
      29175: inst = 32'h8220000;
      29176: inst = 32'h10408000;
      29177: inst = 32'hc404fbc;
      29178: inst = 32'h8220000;
      29179: inst = 32'h10408000;
      29180: inst = 32'hc404fbf;
      29181: inst = 32'h8220000;
      29182: inst = 32'h10408000;
      29183: inst = 32'hc404fc2;
      29184: inst = 32'h8220000;
      29185: inst = 32'h10408000;
      29186: inst = 32'hc404fc4;
      29187: inst = 32'h8220000;
      29188: inst = 32'h10408000;
      29189: inst = 32'hc404fc5;
      29190: inst = 32'h8220000;
      29191: inst = 32'h10408000;
      29192: inst = 32'hc404fc6;
      29193: inst = 32'h8220000;
      29194: inst = 32'h10408000;
      29195: inst = 32'hc404fc7;
      29196: inst = 32'h8220000;
      29197: inst = 32'h10408000;
      29198: inst = 32'hc404fc8;
      29199: inst = 32'h8220000;
      29200: inst = 32'h10408000;
      29201: inst = 32'hc404fc9;
      29202: inst = 32'h8220000;
      29203: inst = 32'h10408000;
      29204: inst = 32'hc404fcc;
      29205: inst = 32'h8220000;
      29206: inst = 32'h10408000;
      29207: inst = 32'hc404fd0;
      29208: inst = 32'h8220000;
      29209: inst = 32'h10408000;
      29210: inst = 32'hc404fd4;
      29211: inst = 32'h8220000;
      29212: inst = 32'h10408000;
      29213: inst = 32'hc404fd5;
      29214: inst = 32'h8220000;
      29215: inst = 32'h10408000;
      29216: inst = 32'hc404fd6;
      29217: inst = 32'h8220000;
      29218: inst = 32'h10408000;
      29219: inst = 32'hc404fd9;
      29220: inst = 32'h8220000;
      29221: inst = 32'h10408000;
      29222: inst = 32'hc404fda;
      29223: inst = 32'h8220000;
      29224: inst = 32'h10408000;
      29225: inst = 32'hc404fe0;
      29226: inst = 32'h8220000;
      29227: inst = 32'h10408000;
      29228: inst = 32'hc404fe2;
      29229: inst = 32'h8220000;
      29230: inst = 32'h10408000;
      29231: inst = 32'hc404fe5;
      29232: inst = 32'h8220000;
      29233: inst = 32'h10408000;
      29234: inst = 32'hc404fe8;
      29235: inst = 32'h8220000;
      29236: inst = 32'h10408000;
      29237: inst = 32'hc404fe9;
      29238: inst = 32'h8220000;
      29239: inst = 32'h10408000;
      29240: inst = 32'hc404fee;
      29241: inst = 32'h8220000;
      29242: inst = 32'h10408000;
      29243: inst = 32'hc404fef;
      29244: inst = 32'h8220000;
      29245: inst = 32'h10408000;
      29246: inst = 32'hc404ff3;
      29247: inst = 32'h8220000;
      29248: inst = 32'h10408000;
      29249: inst = 32'hc404ff6;
      29250: inst = 32'h8220000;
      29251: inst = 32'h10408000;
      29252: inst = 32'hc404ff7;
      29253: inst = 32'h8220000;
      29254: inst = 32'h10408000;
      29255: inst = 32'hc404ff8;
      29256: inst = 32'h8220000;
      29257: inst = 32'h10408000;
      29258: inst = 32'hc405007;
      29259: inst = 32'h8220000;
      29260: inst = 32'h10408000;
      29261: inst = 32'hc405008;
      29262: inst = 32'h8220000;
      29263: inst = 32'h10408000;
      29264: inst = 32'hc405009;
      29265: inst = 32'h8220000;
      29266: inst = 32'h10408000;
      29267: inst = 32'hc40500a;
      29268: inst = 32'h8220000;
      29269: inst = 32'h10408000;
      29270: inst = 32'hc405012;
      29271: inst = 32'h8220000;
      29272: inst = 32'h10408000;
      29273: inst = 32'hc405024;
      29274: inst = 32'h8220000;
      29275: inst = 32'h10408000;
      29276: inst = 32'hc405025;
      29277: inst = 32'h8220000;
      29278: inst = 32'h10408000;
      29279: inst = 32'hc405026;
      29280: inst = 32'h8220000;
      29281: inst = 32'h10408000;
      29282: inst = 32'hc405027;
      29283: inst = 32'h8220000;
      29284: inst = 32'h10408000;
      29285: inst = 32'hc405028;
      29286: inst = 32'h8220000;
      29287: inst = 32'h10408000;
      29288: inst = 32'hc405029;
      29289: inst = 32'h8220000;
      29290: inst = 32'h10408000;
      29291: inst = 32'hc405033;
      29292: inst = 32'h8220000;
      29293: inst = 32'h10408000;
      29294: inst = 32'hc405034;
      29295: inst = 32'h8220000;
      29296: inst = 32'h10408000;
      29297: inst = 32'hc405035;
      29298: inst = 32'h8220000;
      29299: inst = 32'h10408000;
      29300: inst = 32'hc405036;
      29301: inst = 32'h8220000;
      29302: inst = 32'h10408000;
      29303: inst = 32'hc405037;
      29304: inst = 32'h8220000;
      29305: inst = 32'h10408000;
      29306: inst = 32'hc405042;
      29307: inst = 32'h8220000;
      29308: inst = 32'h10408000;
      29309: inst = 32'hc405053;
      29310: inst = 32'h8220000;
      29311: inst = 32'h10408000;
      29312: inst = 32'hc405057;
      29313: inst = 32'h8220000;
      29314: inst = 32'h10408000;
      29315: inst = 32'hc405058;
      29316: inst = 32'h8220000;
      29317: inst = 32'h10408000;
      29318: inst = 32'hc405067;
      29319: inst = 32'h8220000;
      29320: inst = 32'h10408000;
      29321: inst = 32'hc405068;
      29322: inst = 32'h8220000;
      29323: inst = 32'h10408000;
      29324: inst = 32'hc405069;
      29325: inst = 32'h8220000;
      29326: inst = 32'h10408000;
      29327: inst = 32'hc40506a;
      29328: inst = 32'h8220000;
      29329: inst = 32'h10408000;
      29330: inst = 32'hc40506c;
      29331: inst = 32'h8220000;
      29332: inst = 32'h10408000;
      29333: inst = 32'hc40506f;
      29334: inst = 32'h8220000;
      29335: inst = 32'h10408000;
      29336: inst = 32'hc405072;
      29337: inst = 32'h8220000;
      29338: inst = 32'h10408000;
      29339: inst = 32'hc405075;
      29340: inst = 32'h8220000;
      29341: inst = 32'h10408000;
      29342: inst = 32'hc405079;
      29343: inst = 32'h8220000;
      29344: inst = 32'h10408000;
      29345: inst = 32'hc40507a;
      29346: inst = 32'h8220000;
      29347: inst = 32'h10408000;
      29348: inst = 32'hc40507d;
      29349: inst = 32'h8220000;
      29350: inst = 32'h10408000;
      29351: inst = 32'hc40507e;
      29352: inst = 32'h8220000;
      29353: inst = 32'h10408000;
      29354: inst = 32'hc40507f;
      29355: inst = 32'h8220000;
      29356: inst = 32'h10408000;
      29357: inst = 32'hc405080;
      29358: inst = 32'h8220000;
      29359: inst = 32'h10408000;
      29360: inst = 32'hc405083;
      29361: inst = 32'h8220000;
      29362: inst = 32'h10408000;
      29363: inst = 32'hc405084;
      29364: inst = 32'h8220000;
      29365: inst = 32'h10408000;
      29366: inst = 32'hc405085;
      29367: inst = 32'h8220000;
      29368: inst = 32'h10408000;
      29369: inst = 32'hc405086;
      29370: inst = 32'h8220000;
      29371: inst = 32'h10408000;
      29372: inst = 32'hc405087;
      29373: inst = 32'h8220000;
      29374: inst = 32'h10408000;
      29375: inst = 32'hc405088;
      29376: inst = 32'h8220000;
      29377: inst = 32'h10408000;
      29378: inst = 32'hc405089;
      29379: inst = 32'h8220000;
      29380: inst = 32'h10408000;
      29381: inst = 32'hc40508a;
      29382: inst = 32'h8220000;
      29383: inst = 32'h10408000;
      29384: inst = 32'hc40508d;
      29385: inst = 32'h8220000;
      29386: inst = 32'h10408000;
      29387: inst = 32'hc40508e;
      29388: inst = 32'h8220000;
      29389: inst = 32'h10408000;
      29390: inst = 32'hc405092;
      29391: inst = 32'h8220000;
      29392: inst = 32'h10408000;
      29393: inst = 32'hc405093;
      29394: inst = 32'h8220000;
      29395: inst = 32'h10408000;
      29396: inst = 32'hc405094;
      29397: inst = 32'h8220000;
      29398: inst = 32'h10408000;
      29399: inst = 32'hc405095;
      29400: inst = 32'h8220000;
      29401: inst = 32'h10408000;
      29402: inst = 32'hc405096;
      29403: inst = 32'h8220000;
      29404: inst = 32'h10408000;
      29405: inst = 32'hc405097;
      29406: inst = 32'h8220000;
      29407: inst = 32'h10408000;
      29408: inst = 32'hc405098;
      29409: inst = 32'h8220000;
      29410: inst = 32'h10408000;
      29411: inst = 32'hc40509b;
      29412: inst = 32'h8220000;
      29413: inst = 32'h10408000;
      29414: inst = 32'hc40509d;
      29415: inst = 32'h8220000;
      29416: inst = 32'h10408000;
      29417: inst = 32'hc40509e;
      29418: inst = 32'h8220000;
      29419: inst = 32'h10408000;
      29420: inst = 32'hc4050a1;
      29421: inst = 32'h8220000;
      29422: inst = 32'h10408000;
      29423: inst = 32'hc4050a2;
      29424: inst = 32'h8220000;
      29425: inst = 32'h10408000;
      29426: inst = 32'hc4050a3;
      29427: inst = 32'h8220000;
      29428: inst = 32'h10408000;
      29429: inst = 32'hc4050a6;
      29430: inst = 32'h8220000;
      29431: inst = 32'h10408000;
      29432: inst = 32'hc4050a7;
      29433: inst = 32'h8220000;
      29434: inst = 32'h10408000;
      29435: inst = 32'hc4050aa;
      29436: inst = 32'h8220000;
      29437: inst = 32'h10408000;
      29438: inst = 32'hc4050ac;
      29439: inst = 32'h8220000;
      29440: inst = 32'h10408000;
      29441: inst = 32'hc4050b0;
      29442: inst = 32'h8220000;
      29443: inst = 32'h10408000;
      29444: inst = 32'hc4050b3;
      29445: inst = 32'h8220000;
      29446: inst = 32'h10408000;
      29447: inst = 32'hc4050b6;
      29448: inst = 32'h8220000;
      29449: inst = 32'h10408000;
      29450: inst = 32'hc4050b7;
      29451: inst = 32'h8220000;
      29452: inst = 32'h10408000;
      29453: inst = 32'hc4050b8;
      29454: inst = 32'h8220000;
      29455: inst = 32'h10408000;
      29456: inst = 32'hc4050c7;
      29457: inst = 32'h8220000;
      29458: inst = 32'h10408000;
      29459: inst = 32'hc4050c8;
      29460: inst = 32'h8220000;
      29461: inst = 32'h10408000;
      29462: inst = 32'hc4050c9;
      29463: inst = 32'h8220000;
      29464: inst = 32'h10408000;
      29465: inst = 32'hc4050ca;
      29466: inst = 32'h8220000;
      29467: inst = 32'h10408000;
      29468: inst = 32'hc4050cb;
      29469: inst = 32'h8220000;
      29470: inst = 32'h10408000;
      29471: inst = 32'hc4050cc;
      29472: inst = 32'h8220000;
      29473: inst = 32'h10408000;
      29474: inst = 32'hc4050cd;
      29475: inst = 32'h8220000;
      29476: inst = 32'h10408000;
      29477: inst = 32'hc4050ce;
      29478: inst = 32'h8220000;
      29479: inst = 32'h10408000;
      29480: inst = 32'hc4050cf;
      29481: inst = 32'h8220000;
      29482: inst = 32'h10408000;
      29483: inst = 32'hc4050d0;
      29484: inst = 32'h8220000;
      29485: inst = 32'h10408000;
      29486: inst = 32'hc4050d1;
      29487: inst = 32'h8220000;
      29488: inst = 32'h10408000;
      29489: inst = 32'hc4050d2;
      29490: inst = 32'h8220000;
      29491: inst = 32'h10408000;
      29492: inst = 32'hc4050d3;
      29493: inst = 32'h8220000;
      29494: inst = 32'h10408000;
      29495: inst = 32'hc4050d4;
      29496: inst = 32'h8220000;
      29497: inst = 32'h10408000;
      29498: inst = 32'hc4050d5;
      29499: inst = 32'h8220000;
      29500: inst = 32'h10408000;
      29501: inst = 32'hc4050d6;
      29502: inst = 32'h8220000;
      29503: inst = 32'h10408000;
      29504: inst = 32'hc4050d7;
      29505: inst = 32'h8220000;
      29506: inst = 32'h10408000;
      29507: inst = 32'hc4050d8;
      29508: inst = 32'h8220000;
      29509: inst = 32'h10408000;
      29510: inst = 32'hc4050d9;
      29511: inst = 32'h8220000;
      29512: inst = 32'h10408000;
      29513: inst = 32'hc4050da;
      29514: inst = 32'h8220000;
      29515: inst = 32'h10408000;
      29516: inst = 32'hc4050db;
      29517: inst = 32'h8220000;
      29518: inst = 32'h10408000;
      29519: inst = 32'hc4050dc;
      29520: inst = 32'h8220000;
      29521: inst = 32'h10408000;
      29522: inst = 32'hc4050dd;
      29523: inst = 32'h8220000;
      29524: inst = 32'h10408000;
      29525: inst = 32'hc4050de;
      29526: inst = 32'h8220000;
      29527: inst = 32'h10408000;
      29528: inst = 32'hc4050df;
      29529: inst = 32'h8220000;
      29530: inst = 32'h10408000;
      29531: inst = 32'hc4050e0;
      29532: inst = 32'h8220000;
      29533: inst = 32'h10408000;
      29534: inst = 32'hc4050e1;
      29535: inst = 32'h8220000;
      29536: inst = 32'h10408000;
      29537: inst = 32'hc4050e2;
      29538: inst = 32'h8220000;
      29539: inst = 32'h10408000;
      29540: inst = 32'hc4050e3;
      29541: inst = 32'h8220000;
      29542: inst = 32'h10408000;
      29543: inst = 32'hc4050e4;
      29544: inst = 32'h8220000;
      29545: inst = 32'h10408000;
      29546: inst = 32'hc4050e5;
      29547: inst = 32'h8220000;
      29548: inst = 32'h10408000;
      29549: inst = 32'hc4050e6;
      29550: inst = 32'h8220000;
      29551: inst = 32'h10408000;
      29552: inst = 32'hc4050e7;
      29553: inst = 32'h8220000;
      29554: inst = 32'h10408000;
      29555: inst = 32'hc4050e8;
      29556: inst = 32'h8220000;
      29557: inst = 32'h10408000;
      29558: inst = 32'hc4050e9;
      29559: inst = 32'h8220000;
      29560: inst = 32'h10408000;
      29561: inst = 32'hc4050ea;
      29562: inst = 32'h8220000;
      29563: inst = 32'h10408000;
      29564: inst = 32'hc4050eb;
      29565: inst = 32'h8220000;
      29566: inst = 32'h10408000;
      29567: inst = 32'hc4050ec;
      29568: inst = 32'h8220000;
      29569: inst = 32'h10408000;
      29570: inst = 32'hc4050ed;
      29571: inst = 32'h8220000;
      29572: inst = 32'h10408000;
      29573: inst = 32'hc4050ee;
      29574: inst = 32'h8220000;
      29575: inst = 32'h10408000;
      29576: inst = 32'hc4050ef;
      29577: inst = 32'h8220000;
      29578: inst = 32'h10408000;
      29579: inst = 32'hc4050f0;
      29580: inst = 32'h8220000;
      29581: inst = 32'h10408000;
      29582: inst = 32'hc4050f1;
      29583: inst = 32'h8220000;
      29584: inst = 32'h10408000;
      29585: inst = 32'hc4050f2;
      29586: inst = 32'h8220000;
      29587: inst = 32'h10408000;
      29588: inst = 32'hc4050f3;
      29589: inst = 32'h8220000;
      29590: inst = 32'h10408000;
      29591: inst = 32'hc4050f4;
      29592: inst = 32'h8220000;
      29593: inst = 32'h10408000;
      29594: inst = 32'hc4050f5;
      29595: inst = 32'h8220000;
      29596: inst = 32'h10408000;
      29597: inst = 32'hc4050f6;
      29598: inst = 32'h8220000;
      29599: inst = 32'h10408000;
      29600: inst = 32'hc4050f7;
      29601: inst = 32'h8220000;
      29602: inst = 32'h10408000;
      29603: inst = 32'hc4050f8;
      29604: inst = 32'h8220000;
      29605: inst = 32'h10408000;
      29606: inst = 32'hc4050f9;
      29607: inst = 32'h8220000;
      29608: inst = 32'h10408000;
      29609: inst = 32'hc4050fa;
      29610: inst = 32'h8220000;
      29611: inst = 32'h10408000;
      29612: inst = 32'hc4050fb;
      29613: inst = 32'h8220000;
      29614: inst = 32'h10408000;
      29615: inst = 32'hc4050fc;
      29616: inst = 32'h8220000;
      29617: inst = 32'h10408000;
      29618: inst = 32'hc4050fd;
      29619: inst = 32'h8220000;
      29620: inst = 32'h10408000;
      29621: inst = 32'hc4050fe;
      29622: inst = 32'h8220000;
      29623: inst = 32'h10408000;
      29624: inst = 32'hc4050ff;
      29625: inst = 32'h8220000;
      29626: inst = 32'h10408000;
      29627: inst = 32'hc405100;
      29628: inst = 32'h8220000;
      29629: inst = 32'h10408000;
      29630: inst = 32'hc405101;
      29631: inst = 32'h8220000;
      29632: inst = 32'h10408000;
      29633: inst = 32'hc405102;
      29634: inst = 32'h8220000;
      29635: inst = 32'h10408000;
      29636: inst = 32'hc405103;
      29637: inst = 32'h8220000;
      29638: inst = 32'h10408000;
      29639: inst = 32'hc405104;
      29640: inst = 32'h8220000;
      29641: inst = 32'h10408000;
      29642: inst = 32'hc405105;
      29643: inst = 32'h8220000;
      29644: inst = 32'h10408000;
      29645: inst = 32'hc405106;
      29646: inst = 32'h8220000;
      29647: inst = 32'h10408000;
      29648: inst = 32'hc405107;
      29649: inst = 32'h8220000;
      29650: inst = 32'h10408000;
      29651: inst = 32'hc405108;
      29652: inst = 32'h8220000;
      29653: inst = 32'h10408000;
      29654: inst = 32'hc405109;
      29655: inst = 32'h8220000;
      29656: inst = 32'h10408000;
      29657: inst = 32'hc40510a;
      29658: inst = 32'h8220000;
      29659: inst = 32'h10408000;
      29660: inst = 32'hc40510b;
      29661: inst = 32'h8220000;
      29662: inst = 32'h10408000;
      29663: inst = 32'hc40510c;
      29664: inst = 32'h8220000;
      29665: inst = 32'h10408000;
      29666: inst = 32'hc40510d;
      29667: inst = 32'h8220000;
      29668: inst = 32'h10408000;
      29669: inst = 32'hc40510e;
      29670: inst = 32'h8220000;
      29671: inst = 32'h10408000;
      29672: inst = 32'hc40510f;
      29673: inst = 32'h8220000;
      29674: inst = 32'h10408000;
      29675: inst = 32'hc405110;
      29676: inst = 32'h8220000;
      29677: inst = 32'h10408000;
      29678: inst = 32'hc405111;
      29679: inst = 32'h8220000;
      29680: inst = 32'h10408000;
      29681: inst = 32'hc405112;
      29682: inst = 32'h8220000;
      29683: inst = 32'h10408000;
      29684: inst = 32'hc405113;
      29685: inst = 32'h8220000;
      29686: inst = 32'h10408000;
      29687: inst = 32'hc405114;
      29688: inst = 32'h8220000;
      29689: inst = 32'h10408000;
      29690: inst = 32'hc405115;
      29691: inst = 32'h8220000;
      29692: inst = 32'h10408000;
      29693: inst = 32'hc405116;
      29694: inst = 32'h8220000;
      29695: inst = 32'h10408000;
      29696: inst = 32'hc405117;
      29697: inst = 32'h8220000;
      29698: inst = 32'h10408000;
      29699: inst = 32'hc405118;
      29700: inst = 32'h8220000;
      29701: inst = 32'h10408000;
      29702: inst = 32'hc405127;
      29703: inst = 32'h8220000;
      29704: inst = 32'h10408000;
      29705: inst = 32'hc405128;
      29706: inst = 32'h8220000;
      29707: inst = 32'h10408000;
      29708: inst = 32'hc405129;
      29709: inst = 32'h8220000;
      29710: inst = 32'h10408000;
      29711: inst = 32'hc40512a;
      29712: inst = 32'h8220000;
      29713: inst = 32'h10408000;
      29714: inst = 32'hc40512b;
      29715: inst = 32'h8220000;
      29716: inst = 32'h10408000;
      29717: inst = 32'hc40512c;
      29718: inst = 32'h8220000;
      29719: inst = 32'h10408000;
      29720: inst = 32'hc40512d;
      29721: inst = 32'h8220000;
      29722: inst = 32'h10408000;
      29723: inst = 32'hc40512e;
      29724: inst = 32'h8220000;
      29725: inst = 32'h10408000;
      29726: inst = 32'hc40512f;
      29727: inst = 32'h8220000;
      29728: inst = 32'h10408000;
      29729: inst = 32'hc405130;
      29730: inst = 32'h8220000;
      29731: inst = 32'h10408000;
      29732: inst = 32'hc405131;
      29733: inst = 32'h8220000;
      29734: inst = 32'h10408000;
      29735: inst = 32'hc405132;
      29736: inst = 32'h8220000;
      29737: inst = 32'h10408000;
      29738: inst = 32'hc405133;
      29739: inst = 32'h8220000;
      29740: inst = 32'h10408000;
      29741: inst = 32'hc405134;
      29742: inst = 32'h8220000;
      29743: inst = 32'h10408000;
      29744: inst = 32'hc405135;
      29745: inst = 32'h8220000;
      29746: inst = 32'h10408000;
      29747: inst = 32'hc405136;
      29748: inst = 32'h8220000;
      29749: inst = 32'h10408000;
      29750: inst = 32'hc405137;
      29751: inst = 32'h8220000;
      29752: inst = 32'h10408000;
      29753: inst = 32'hc405138;
      29754: inst = 32'h8220000;
      29755: inst = 32'h10408000;
      29756: inst = 32'hc405139;
      29757: inst = 32'h8220000;
      29758: inst = 32'h10408000;
      29759: inst = 32'hc40513a;
      29760: inst = 32'h8220000;
      29761: inst = 32'h10408000;
      29762: inst = 32'hc40513b;
      29763: inst = 32'h8220000;
      29764: inst = 32'h10408000;
      29765: inst = 32'hc40513c;
      29766: inst = 32'h8220000;
      29767: inst = 32'h10408000;
      29768: inst = 32'hc40513d;
      29769: inst = 32'h8220000;
      29770: inst = 32'h10408000;
      29771: inst = 32'hc40513e;
      29772: inst = 32'h8220000;
      29773: inst = 32'h10408000;
      29774: inst = 32'hc40513f;
      29775: inst = 32'h8220000;
      29776: inst = 32'h10408000;
      29777: inst = 32'hc405140;
      29778: inst = 32'h8220000;
      29779: inst = 32'h10408000;
      29780: inst = 32'hc405141;
      29781: inst = 32'h8220000;
      29782: inst = 32'h10408000;
      29783: inst = 32'hc405142;
      29784: inst = 32'h8220000;
      29785: inst = 32'h10408000;
      29786: inst = 32'hc405143;
      29787: inst = 32'h8220000;
      29788: inst = 32'h10408000;
      29789: inst = 32'hc405144;
      29790: inst = 32'h8220000;
      29791: inst = 32'h10408000;
      29792: inst = 32'hc405145;
      29793: inst = 32'h8220000;
      29794: inst = 32'h10408000;
      29795: inst = 32'hc405146;
      29796: inst = 32'h8220000;
      29797: inst = 32'h10408000;
      29798: inst = 32'hc405147;
      29799: inst = 32'h8220000;
      29800: inst = 32'h10408000;
      29801: inst = 32'hc405148;
      29802: inst = 32'h8220000;
      29803: inst = 32'h10408000;
      29804: inst = 32'hc405149;
      29805: inst = 32'h8220000;
      29806: inst = 32'h10408000;
      29807: inst = 32'hc40514a;
      29808: inst = 32'h8220000;
      29809: inst = 32'h10408000;
      29810: inst = 32'hc40514b;
      29811: inst = 32'h8220000;
      29812: inst = 32'h10408000;
      29813: inst = 32'hc40514c;
      29814: inst = 32'h8220000;
      29815: inst = 32'h10408000;
      29816: inst = 32'hc40514d;
      29817: inst = 32'h8220000;
      29818: inst = 32'h10408000;
      29819: inst = 32'hc40514e;
      29820: inst = 32'h8220000;
      29821: inst = 32'h10408000;
      29822: inst = 32'hc40514f;
      29823: inst = 32'h8220000;
      29824: inst = 32'h10408000;
      29825: inst = 32'hc405150;
      29826: inst = 32'h8220000;
      29827: inst = 32'h10408000;
      29828: inst = 32'hc405151;
      29829: inst = 32'h8220000;
      29830: inst = 32'h10408000;
      29831: inst = 32'hc405152;
      29832: inst = 32'h8220000;
      29833: inst = 32'h10408000;
      29834: inst = 32'hc405153;
      29835: inst = 32'h8220000;
      29836: inst = 32'h10408000;
      29837: inst = 32'hc405154;
      29838: inst = 32'h8220000;
      29839: inst = 32'h10408000;
      29840: inst = 32'hc405155;
      29841: inst = 32'h8220000;
      29842: inst = 32'h10408000;
      29843: inst = 32'hc405156;
      29844: inst = 32'h8220000;
      29845: inst = 32'h10408000;
      29846: inst = 32'hc405157;
      29847: inst = 32'h8220000;
      29848: inst = 32'h10408000;
      29849: inst = 32'hc405158;
      29850: inst = 32'h8220000;
      29851: inst = 32'h10408000;
      29852: inst = 32'hc405159;
      29853: inst = 32'h8220000;
      29854: inst = 32'h10408000;
      29855: inst = 32'hc40515a;
      29856: inst = 32'h8220000;
      29857: inst = 32'h10408000;
      29858: inst = 32'hc40515b;
      29859: inst = 32'h8220000;
      29860: inst = 32'h10408000;
      29861: inst = 32'hc40515c;
      29862: inst = 32'h8220000;
      29863: inst = 32'h10408000;
      29864: inst = 32'hc40515d;
      29865: inst = 32'h8220000;
      29866: inst = 32'h10408000;
      29867: inst = 32'hc40515e;
      29868: inst = 32'h8220000;
      29869: inst = 32'h10408000;
      29870: inst = 32'hc40515f;
      29871: inst = 32'h8220000;
      29872: inst = 32'h10408000;
      29873: inst = 32'hc405160;
      29874: inst = 32'h8220000;
      29875: inst = 32'h10408000;
      29876: inst = 32'hc405161;
      29877: inst = 32'h8220000;
      29878: inst = 32'h10408000;
      29879: inst = 32'hc405162;
      29880: inst = 32'h8220000;
      29881: inst = 32'h10408000;
      29882: inst = 32'hc405163;
      29883: inst = 32'h8220000;
      29884: inst = 32'h10408000;
      29885: inst = 32'hc405164;
      29886: inst = 32'h8220000;
      29887: inst = 32'h10408000;
      29888: inst = 32'hc405165;
      29889: inst = 32'h8220000;
      29890: inst = 32'h10408000;
      29891: inst = 32'hc405166;
      29892: inst = 32'h8220000;
      29893: inst = 32'h10408000;
      29894: inst = 32'hc405167;
      29895: inst = 32'h8220000;
      29896: inst = 32'h10408000;
      29897: inst = 32'hc405168;
      29898: inst = 32'h8220000;
      29899: inst = 32'h10408000;
      29900: inst = 32'hc405169;
      29901: inst = 32'h8220000;
      29902: inst = 32'h10408000;
      29903: inst = 32'hc40516a;
      29904: inst = 32'h8220000;
      29905: inst = 32'h10408000;
      29906: inst = 32'hc40516b;
      29907: inst = 32'h8220000;
      29908: inst = 32'h10408000;
      29909: inst = 32'hc40516c;
      29910: inst = 32'h8220000;
      29911: inst = 32'h10408000;
      29912: inst = 32'hc40516d;
      29913: inst = 32'h8220000;
      29914: inst = 32'h10408000;
      29915: inst = 32'hc40516e;
      29916: inst = 32'h8220000;
      29917: inst = 32'h10408000;
      29918: inst = 32'hc40516f;
      29919: inst = 32'h8220000;
      29920: inst = 32'h10408000;
      29921: inst = 32'hc405170;
      29922: inst = 32'h8220000;
      29923: inst = 32'h10408000;
      29924: inst = 32'hc405171;
      29925: inst = 32'h8220000;
      29926: inst = 32'h10408000;
      29927: inst = 32'hc405172;
      29928: inst = 32'h8220000;
      29929: inst = 32'h10408000;
      29930: inst = 32'hc405173;
      29931: inst = 32'h8220000;
      29932: inst = 32'h10408000;
      29933: inst = 32'hc405174;
      29934: inst = 32'h8220000;
      29935: inst = 32'h10408000;
      29936: inst = 32'hc405175;
      29937: inst = 32'h8220000;
      29938: inst = 32'h10408000;
      29939: inst = 32'hc405176;
      29940: inst = 32'h8220000;
      29941: inst = 32'h10408000;
      29942: inst = 32'hc405177;
      29943: inst = 32'h8220000;
      29944: inst = 32'h10408000;
      29945: inst = 32'hc405178;
      29946: inst = 32'h8220000;
      29947: inst = 32'h10408000;
      29948: inst = 32'hc405187;
      29949: inst = 32'h8220000;
      29950: inst = 32'h10408000;
      29951: inst = 32'hc405188;
      29952: inst = 32'h8220000;
      29953: inst = 32'h10408000;
      29954: inst = 32'hc405189;
      29955: inst = 32'h8220000;
      29956: inst = 32'h10408000;
      29957: inst = 32'hc40518a;
      29958: inst = 32'h8220000;
      29959: inst = 32'h10408000;
      29960: inst = 32'hc40518b;
      29961: inst = 32'h8220000;
      29962: inst = 32'h10408000;
      29963: inst = 32'hc40518c;
      29964: inst = 32'h8220000;
      29965: inst = 32'h10408000;
      29966: inst = 32'hc40518d;
      29967: inst = 32'h8220000;
      29968: inst = 32'h10408000;
      29969: inst = 32'hc40518e;
      29970: inst = 32'h8220000;
      29971: inst = 32'h10408000;
      29972: inst = 32'hc40518f;
      29973: inst = 32'h8220000;
      29974: inst = 32'h10408000;
      29975: inst = 32'hc405190;
      29976: inst = 32'h8220000;
      29977: inst = 32'h10408000;
      29978: inst = 32'hc405191;
      29979: inst = 32'h8220000;
      29980: inst = 32'h10408000;
      29981: inst = 32'hc405192;
      29982: inst = 32'h8220000;
      29983: inst = 32'h10408000;
      29984: inst = 32'hc405193;
      29985: inst = 32'h8220000;
      29986: inst = 32'h10408000;
      29987: inst = 32'hc405194;
      29988: inst = 32'h8220000;
      29989: inst = 32'h10408000;
      29990: inst = 32'hc405195;
      29991: inst = 32'h8220000;
      29992: inst = 32'h10408000;
      29993: inst = 32'hc405196;
      29994: inst = 32'h8220000;
      29995: inst = 32'h10408000;
      29996: inst = 32'hc405197;
      29997: inst = 32'h8220000;
      29998: inst = 32'h10408000;
      29999: inst = 32'hc405198;
      30000: inst = 32'h8220000;
      30001: inst = 32'h10408000;
      30002: inst = 32'hc405199;
      30003: inst = 32'h8220000;
      30004: inst = 32'h10408000;
      30005: inst = 32'hc40519a;
      30006: inst = 32'h8220000;
      30007: inst = 32'h10408000;
      30008: inst = 32'hc40519b;
      30009: inst = 32'h8220000;
      30010: inst = 32'h10408000;
      30011: inst = 32'hc40519c;
      30012: inst = 32'h8220000;
      30013: inst = 32'h10408000;
      30014: inst = 32'hc40519d;
      30015: inst = 32'h8220000;
      30016: inst = 32'h10408000;
      30017: inst = 32'hc40519e;
      30018: inst = 32'h8220000;
      30019: inst = 32'h10408000;
      30020: inst = 32'hc40519f;
      30021: inst = 32'h8220000;
      30022: inst = 32'h10408000;
      30023: inst = 32'hc4051a0;
      30024: inst = 32'h8220000;
      30025: inst = 32'h10408000;
      30026: inst = 32'hc4051a1;
      30027: inst = 32'h8220000;
      30028: inst = 32'h10408000;
      30029: inst = 32'hc4051a2;
      30030: inst = 32'h8220000;
      30031: inst = 32'h10408000;
      30032: inst = 32'hc4051a3;
      30033: inst = 32'h8220000;
      30034: inst = 32'h10408000;
      30035: inst = 32'hc4051a4;
      30036: inst = 32'h8220000;
      30037: inst = 32'h10408000;
      30038: inst = 32'hc4051a5;
      30039: inst = 32'h8220000;
      30040: inst = 32'h10408000;
      30041: inst = 32'hc4051a6;
      30042: inst = 32'h8220000;
      30043: inst = 32'h10408000;
      30044: inst = 32'hc4051a7;
      30045: inst = 32'h8220000;
      30046: inst = 32'h10408000;
      30047: inst = 32'hc4051a8;
      30048: inst = 32'h8220000;
      30049: inst = 32'h10408000;
      30050: inst = 32'hc4051a9;
      30051: inst = 32'h8220000;
      30052: inst = 32'h10408000;
      30053: inst = 32'hc4051aa;
      30054: inst = 32'h8220000;
      30055: inst = 32'h10408000;
      30056: inst = 32'hc4051ab;
      30057: inst = 32'h8220000;
      30058: inst = 32'h10408000;
      30059: inst = 32'hc4051ac;
      30060: inst = 32'h8220000;
      30061: inst = 32'h10408000;
      30062: inst = 32'hc4051ad;
      30063: inst = 32'h8220000;
      30064: inst = 32'h10408000;
      30065: inst = 32'hc4051ae;
      30066: inst = 32'h8220000;
      30067: inst = 32'h10408000;
      30068: inst = 32'hc4051af;
      30069: inst = 32'h8220000;
      30070: inst = 32'h10408000;
      30071: inst = 32'hc4051b0;
      30072: inst = 32'h8220000;
      30073: inst = 32'h10408000;
      30074: inst = 32'hc4051b1;
      30075: inst = 32'h8220000;
      30076: inst = 32'h10408000;
      30077: inst = 32'hc4051b2;
      30078: inst = 32'h8220000;
      30079: inst = 32'h10408000;
      30080: inst = 32'hc4051b3;
      30081: inst = 32'h8220000;
      30082: inst = 32'h10408000;
      30083: inst = 32'hc4051b4;
      30084: inst = 32'h8220000;
      30085: inst = 32'h10408000;
      30086: inst = 32'hc4051b5;
      30087: inst = 32'h8220000;
      30088: inst = 32'h10408000;
      30089: inst = 32'hc4051b6;
      30090: inst = 32'h8220000;
      30091: inst = 32'h10408000;
      30092: inst = 32'hc4051b7;
      30093: inst = 32'h8220000;
      30094: inst = 32'h10408000;
      30095: inst = 32'hc4051b8;
      30096: inst = 32'h8220000;
      30097: inst = 32'h10408000;
      30098: inst = 32'hc4051b9;
      30099: inst = 32'h8220000;
      30100: inst = 32'h10408000;
      30101: inst = 32'hc4051ba;
      30102: inst = 32'h8220000;
      30103: inst = 32'h10408000;
      30104: inst = 32'hc4051bb;
      30105: inst = 32'h8220000;
      30106: inst = 32'h10408000;
      30107: inst = 32'hc4051bc;
      30108: inst = 32'h8220000;
      30109: inst = 32'h10408000;
      30110: inst = 32'hc4051bd;
      30111: inst = 32'h8220000;
      30112: inst = 32'h10408000;
      30113: inst = 32'hc4051be;
      30114: inst = 32'h8220000;
      30115: inst = 32'h10408000;
      30116: inst = 32'hc4051bf;
      30117: inst = 32'h8220000;
      30118: inst = 32'h10408000;
      30119: inst = 32'hc4051c0;
      30120: inst = 32'h8220000;
      30121: inst = 32'h10408000;
      30122: inst = 32'hc4051c1;
      30123: inst = 32'h8220000;
      30124: inst = 32'h10408000;
      30125: inst = 32'hc4051c2;
      30126: inst = 32'h8220000;
      30127: inst = 32'h10408000;
      30128: inst = 32'hc4051c3;
      30129: inst = 32'h8220000;
      30130: inst = 32'h10408000;
      30131: inst = 32'hc4051c4;
      30132: inst = 32'h8220000;
      30133: inst = 32'h10408000;
      30134: inst = 32'hc4051c5;
      30135: inst = 32'h8220000;
      30136: inst = 32'h10408000;
      30137: inst = 32'hc4051c6;
      30138: inst = 32'h8220000;
      30139: inst = 32'h10408000;
      30140: inst = 32'hc4051c7;
      30141: inst = 32'h8220000;
      30142: inst = 32'h10408000;
      30143: inst = 32'hc4051c8;
      30144: inst = 32'h8220000;
      30145: inst = 32'h10408000;
      30146: inst = 32'hc4051c9;
      30147: inst = 32'h8220000;
      30148: inst = 32'h10408000;
      30149: inst = 32'hc4051ca;
      30150: inst = 32'h8220000;
      30151: inst = 32'h10408000;
      30152: inst = 32'hc4051cb;
      30153: inst = 32'h8220000;
      30154: inst = 32'h10408000;
      30155: inst = 32'hc4051cc;
      30156: inst = 32'h8220000;
      30157: inst = 32'h10408000;
      30158: inst = 32'hc4051cd;
      30159: inst = 32'h8220000;
      30160: inst = 32'h10408000;
      30161: inst = 32'hc4051ce;
      30162: inst = 32'h8220000;
      30163: inst = 32'h10408000;
      30164: inst = 32'hc4051cf;
      30165: inst = 32'h8220000;
      30166: inst = 32'h10408000;
      30167: inst = 32'hc4051d0;
      30168: inst = 32'h8220000;
      30169: inst = 32'h10408000;
      30170: inst = 32'hc4051d1;
      30171: inst = 32'h8220000;
      30172: inst = 32'h10408000;
      30173: inst = 32'hc4051d2;
      30174: inst = 32'h8220000;
      30175: inst = 32'h10408000;
      30176: inst = 32'hc4051d3;
      30177: inst = 32'h8220000;
      30178: inst = 32'h10408000;
      30179: inst = 32'hc4051d4;
      30180: inst = 32'h8220000;
      30181: inst = 32'h10408000;
      30182: inst = 32'hc4051d5;
      30183: inst = 32'h8220000;
      30184: inst = 32'h10408000;
      30185: inst = 32'hc4051d6;
      30186: inst = 32'h8220000;
      30187: inst = 32'h10408000;
      30188: inst = 32'hc4051d7;
      30189: inst = 32'h8220000;
      30190: inst = 32'h10408000;
      30191: inst = 32'hc4051d8;
      30192: inst = 32'h8220000;
      30193: inst = 32'h10408000;
      30194: inst = 32'hc4051e7;
      30195: inst = 32'h8220000;
      30196: inst = 32'h10408000;
      30197: inst = 32'hc4051e8;
      30198: inst = 32'h8220000;
      30199: inst = 32'h10408000;
      30200: inst = 32'hc4051e9;
      30201: inst = 32'h8220000;
      30202: inst = 32'h10408000;
      30203: inst = 32'hc4051ea;
      30204: inst = 32'h8220000;
      30205: inst = 32'h10408000;
      30206: inst = 32'hc4051eb;
      30207: inst = 32'h8220000;
      30208: inst = 32'h10408000;
      30209: inst = 32'hc4051ec;
      30210: inst = 32'h8220000;
      30211: inst = 32'h10408000;
      30212: inst = 32'hc4051ed;
      30213: inst = 32'h8220000;
      30214: inst = 32'h10408000;
      30215: inst = 32'hc4051ee;
      30216: inst = 32'h8220000;
      30217: inst = 32'h10408000;
      30218: inst = 32'hc4051ef;
      30219: inst = 32'h8220000;
      30220: inst = 32'h10408000;
      30221: inst = 32'hc4051f0;
      30222: inst = 32'h8220000;
      30223: inst = 32'h10408000;
      30224: inst = 32'hc4051f1;
      30225: inst = 32'h8220000;
      30226: inst = 32'h10408000;
      30227: inst = 32'hc4051f2;
      30228: inst = 32'h8220000;
      30229: inst = 32'h10408000;
      30230: inst = 32'hc4051f3;
      30231: inst = 32'h8220000;
      30232: inst = 32'h10408000;
      30233: inst = 32'hc4051f4;
      30234: inst = 32'h8220000;
      30235: inst = 32'h10408000;
      30236: inst = 32'hc4051f5;
      30237: inst = 32'h8220000;
      30238: inst = 32'h10408000;
      30239: inst = 32'hc4051f6;
      30240: inst = 32'h8220000;
      30241: inst = 32'h10408000;
      30242: inst = 32'hc4051f7;
      30243: inst = 32'h8220000;
      30244: inst = 32'h10408000;
      30245: inst = 32'hc4051f8;
      30246: inst = 32'h8220000;
      30247: inst = 32'h10408000;
      30248: inst = 32'hc4051f9;
      30249: inst = 32'h8220000;
      30250: inst = 32'h10408000;
      30251: inst = 32'hc4051fa;
      30252: inst = 32'h8220000;
      30253: inst = 32'h10408000;
      30254: inst = 32'hc4051fb;
      30255: inst = 32'h8220000;
      30256: inst = 32'h10408000;
      30257: inst = 32'hc4051fc;
      30258: inst = 32'h8220000;
      30259: inst = 32'h10408000;
      30260: inst = 32'hc4051fd;
      30261: inst = 32'h8220000;
      30262: inst = 32'h10408000;
      30263: inst = 32'hc4051fe;
      30264: inst = 32'h8220000;
      30265: inst = 32'h10408000;
      30266: inst = 32'hc4051ff;
      30267: inst = 32'h8220000;
      30268: inst = 32'h10408000;
      30269: inst = 32'hc405200;
      30270: inst = 32'h8220000;
      30271: inst = 32'h10408000;
      30272: inst = 32'hc405201;
      30273: inst = 32'h8220000;
      30274: inst = 32'h10408000;
      30275: inst = 32'hc405202;
      30276: inst = 32'h8220000;
      30277: inst = 32'h10408000;
      30278: inst = 32'hc405203;
      30279: inst = 32'h8220000;
      30280: inst = 32'h10408000;
      30281: inst = 32'hc405204;
      30282: inst = 32'h8220000;
      30283: inst = 32'h10408000;
      30284: inst = 32'hc405205;
      30285: inst = 32'h8220000;
      30286: inst = 32'h10408000;
      30287: inst = 32'hc405206;
      30288: inst = 32'h8220000;
      30289: inst = 32'h10408000;
      30290: inst = 32'hc405207;
      30291: inst = 32'h8220000;
      30292: inst = 32'h10408000;
      30293: inst = 32'hc405208;
      30294: inst = 32'h8220000;
      30295: inst = 32'h10408000;
      30296: inst = 32'hc405209;
      30297: inst = 32'h8220000;
      30298: inst = 32'h10408000;
      30299: inst = 32'hc40520a;
      30300: inst = 32'h8220000;
      30301: inst = 32'h10408000;
      30302: inst = 32'hc40520b;
      30303: inst = 32'h8220000;
      30304: inst = 32'h10408000;
      30305: inst = 32'hc40520c;
      30306: inst = 32'h8220000;
      30307: inst = 32'h10408000;
      30308: inst = 32'hc40520d;
      30309: inst = 32'h8220000;
      30310: inst = 32'h10408000;
      30311: inst = 32'hc40520e;
      30312: inst = 32'h8220000;
      30313: inst = 32'h10408000;
      30314: inst = 32'hc40520f;
      30315: inst = 32'h8220000;
      30316: inst = 32'h10408000;
      30317: inst = 32'hc405210;
      30318: inst = 32'h8220000;
      30319: inst = 32'h10408000;
      30320: inst = 32'hc405211;
      30321: inst = 32'h8220000;
      30322: inst = 32'h10408000;
      30323: inst = 32'hc405212;
      30324: inst = 32'h8220000;
      30325: inst = 32'h10408000;
      30326: inst = 32'hc405213;
      30327: inst = 32'h8220000;
      30328: inst = 32'h10408000;
      30329: inst = 32'hc405214;
      30330: inst = 32'h8220000;
      30331: inst = 32'h10408000;
      30332: inst = 32'hc405215;
      30333: inst = 32'h8220000;
      30334: inst = 32'h10408000;
      30335: inst = 32'hc405216;
      30336: inst = 32'h8220000;
      30337: inst = 32'h10408000;
      30338: inst = 32'hc405217;
      30339: inst = 32'h8220000;
      30340: inst = 32'h10408000;
      30341: inst = 32'hc405218;
      30342: inst = 32'h8220000;
      30343: inst = 32'h10408000;
      30344: inst = 32'hc405219;
      30345: inst = 32'h8220000;
      30346: inst = 32'h10408000;
      30347: inst = 32'hc40521a;
      30348: inst = 32'h8220000;
      30349: inst = 32'h10408000;
      30350: inst = 32'hc40521b;
      30351: inst = 32'h8220000;
      30352: inst = 32'h10408000;
      30353: inst = 32'hc40521c;
      30354: inst = 32'h8220000;
      30355: inst = 32'h10408000;
      30356: inst = 32'hc40521d;
      30357: inst = 32'h8220000;
      30358: inst = 32'h10408000;
      30359: inst = 32'hc40521e;
      30360: inst = 32'h8220000;
      30361: inst = 32'h10408000;
      30362: inst = 32'hc40521f;
      30363: inst = 32'h8220000;
      30364: inst = 32'h10408000;
      30365: inst = 32'hc405220;
      30366: inst = 32'h8220000;
      30367: inst = 32'h10408000;
      30368: inst = 32'hc405221;
      30369: inst = 32'h8220000;
      30370: inst = 32'h10408000;
      30371: inst = 32'hc405222;
      30372: inst = 32'h8220000;
      30373: inst = 32'h10408000;
      30374: inst = 32'hc405223;
      30375: inst = 32'h8220000;
      30376: inst = 32'h10408000;
      30377: inst = 32'hc405224;
      30378: inst = 32'h8220000;
      30379: inst = 32'h10408000;
      30380: inst = 32'hc405225;
      30381: inst = 32'h8220000;
      30382: inst = 32'h10408000;
      30383: inst = 32'hc405226;
      30384: inst = 32'h8220000;
      30385: inst = 32'h10408000;
      30386: inst = 32'hc405227;
      30387: inst = 32'h8220000;
      30388: inst = 32'h10408000;
      30389: inst = 32'hc405228;
      30390: inst = 32'h8220000;
      30391: inst = 32'h10408000;
      30392: inst = 32'hc405229;
      30393: inst = 32'h8220000;
      30394: inst = 32'h10408000;
      30395: inst = 32'hc40522a;
      30396: inst = 32'h8220000;
      30397: inst = 32'h10408000;
      30398: inst = 32'hc40522b;
      30399: inst = 32'h8220000;
      30400: inst = 32'h10408000;
      30401: inst = 32'hc40522c;
      30402: inst = 32'h8220000;
      30403: inst = 32'h10408000;
      30404: inst = 32'hc40522d;
      30405: inst = 32'h8220000;
      30406: inst = 32'h10408000;
      30407: inst = 32'hc40522e;
      30408: inst = 32'h8220000;
      30409: inst = 32'h10408000;
      30410: inst = 32'hc40522f;
      30411: inst = 32'h8220000;
      30412: inst = 32'h10408000;
      30413: inst = 32'hc405230;
      30414: inst = 32'h8220000;
      30415: inst = 32'h10408000;
      30416: inst = 32'hc405231;
      30417: inst = 32'h8220000;
      30418: inst = 32'h10408000;
      30419: inst = 32'hc405232;
      30420: inst = 32'h8220000;
      30421: inst = 32'h10408000;
      30422: inst = 32'hc405233;
      30423: inst = 32'h8220000;
      30424: inst = 32'h10408000;
      30425: inst = 32'hc405234;
      30426: inst = 32'h8220000;
      30427: inst = 32'h10408000;
      30428: inst = 32'hc405235;
      30429: inst = 32'h8220000;
      30430: inst = 32'h10408000;
      30431: inst = 32'hc405236;
      30432: inst = 32'h8220000;
      30433: inst = 32'h10408000;
      30434: inst = 32'hc405237;
      30435: inst = 32'h8220000;
      30436: inst = 32'h10408000;
      30437: inst = 32'hc405238;
      30438: inst = 32'h8220000;
      30439: inst = 32'h10408000;
      30440: inst = 32'hc405247;
      30441: inst = 32'h8220000;
      30442: inst = 32'h10408000;
      30443: inst = 32'hc405248;
      30444: inst = 32'h8220000;
      30445: inst = 32'h10408000;
      30446: inst = 32'hc405249;
      30447: inst = 32'h8220000;
      30448: inst = 32'h10408000;
      30449: inst = 32'hc40524a;
      30450: inst = 32'h8220000;
      30451: inst = 32'h10408000;
      30452: inst = 32'hc40524b;
      30453: inst = 32'h8220000;
      30454: inst = 32'h10408000;
      30455: inst = 32'hc40524c;
      30456: inst = 32'h8220000;
      30457: inst = 32'h10408000;
      30458: inst = 32'hc40524d;
      30459: inst = 32'h8220000;
      30460: inst = 32'h10408000;
      30461: inst = 32'hc40524e;
      30462: inst = 32'h8220000;
      30463: inst = 32'h10408000;
      30464: inst = 32'hc40524f;
      30465: inst = 32'h8220000;
      30466: inst = 32'h10408000;
      30467: inst = 32'hc405250;
      30468: inst = 32'h8220000;
      30469: inst = 32'h10408000;
      30470: inst = 32'hc405251;
      30471: inst = 32'h8220000;
      30472: inst = 32'h10408000;
      30473: inst = 32'hc405252;
      30474: inst = 32'h8220000;
      30475: inst = 32'h10408000;
      30476: inst = 32'hc405253;
      30477: inst = 32'h8220000;
      30478: inst = 32'h10408000;
      30479: inst = 32'hc405254;
      30480: inst = 32'h8220000;
      30481: inst = 32'h10408000;
      30482: inst = 32'hc405255;
      30483: inst = 32'h8220000;
      30484: inst = 32'h10408000;
      30485: inst = 32'hc405256;
      30486: inst = 32'h8220000;
      30487: inst = 32'h10408000;
      30488: inst = 32'hc405257;
      30489: inst = 32'h8220000;
      30490: inst = 32'h10408000;
      30491: inst = 32'hc405258;
      30492: inst = 32'h8220000;
      30493: inst = 32'h10408000;
      30494: inst = 32'hc405259;
      30495: inst = 32'h8220000;
      30496: inst = 32'h10408000;
      30497: inst = 32'hc40525a;
      30498: inst = 32'h8220000;
      30499: inst = 32'h10408000;
      30500: inst = 32'hc40525b;
      30501: inst = 32'h8220000;
      30502: inst = 32'h10408000;
      30503: inst = 32'hc40525c;
      30504: inst = 32'h8220000;
      30505: inst = 32'h10408000;
      30506: inst = 32'hc40525d;
      30507: inst = 32'h8220000;
      30508: inst = 32'h10408000;
      30509: inst = 32'hc40525e;
      30510: inst = 32'h8220000;
      30511: inst = 32'h10408000;
      30512: inst = 32'hc40525f;
      30513: inst = 32'h8220000;
      30514: inst = 32'h10408000;
      30515: inst = 32'hc405260;
      30516: inst = 32'h8220000;
      30517: inst = 32'h10408000;
      30518: inst = 32'hc405261;
      30519: inst = 32'h8220000;
      30520: inst = 32'h10408000;
      30521: inst = 32'hc405262;
      30522: inst = 32'h8220000;
      30523: inst = 32'h10408000;
      30524: inst = 32'hc405263;
      30525: inst = 32'h8220000;
      30526: inst = 32'h10408000;
      30527: inst = 32'hc405264;
      30528: inst = 32'h8220000;
      30529: inst = 32'h10408000;
      30530: inst = 32'hc405265;
      30531: inst = 32'h8220000;
      30532: inst = 32'h10408000;
      30533: inst = 32'hc405266;
      30534: inst = 32'h8220000;
      30535: inst = 32'h10408000;
      30536: inst = 32'hc405267;
      30537: inst = 32'h8220000;
      30538: inst = 32'h10408000;
      30539: inst = 32'hc405268;
      30540: inst = 32'h8220000;
      30541: inst = 32'h10408000;
      30542: inst = 32'hc405269;
      30543: inst = 32'h8220000;
      30544: inst = 32'h10408000;
      30545: inst = 32'hc40526a;
      30546: inst = 32'h8220000;
      30547: inst = 32'h10408000;
      30548: inst = 32'hc40526b;
      30549: inst = 32'h8220000;
      30550: inst = 32'h10408000;
      30551: inst = 32'hc40526c;
      30552: inst = 32'h8220000;
      30553: inst = 32'h10408000;
      30554: inst = 32'hc40526d;
      30555: inst = 32'h8220000;
      30556: inst = 32'h10408000;
      30557: inst = 32'hc40526e;
      30558: inst = 32'h8220000;
      30559: inst = 32'h10408000;
      30560: inst = 32'hc40526f;
      30561: inst = 32'h8220000;
      30562: inst = 32'h10408000;
      30563: inst = 32'hc405270;
      30564: inst = 32'h8220000;
      30565: inst = 32'h10408000;
      30566: inst = 32'hc405271;
      30567: inst = 32'h8220000;
      30568: inst = 32'h10408000;
      30569: inst = 32'hc405272;
      30570: inst = 32'h8220000;
      30571: inst = 32'h10408000;
      30572: inst = 32'hc405273;
      30573: inst = 32'h8220000;
      30574: inst = 32'h10408000;
      30575: inst = 32'hc405274;
      30576: inst = 32'h8220000;
      30577: inst = 32'h10408000;
      30578: inst = 32'hc405275;
      30579: inst = 32'h8220000;
      30580: inst = 32'h10408000;
      30581: inst = 32'hc405276;
      30582: inst = 32'h8220000;
      30583: inst = 32'h10408000;
      30584: inst = 32'hc405277;
      30585: inst = 32'h8220000;
      30586: inst = 32'h10408000;
      30587: inst = 32'hc405278;
      30588: inst = 32'h8220000;
      30589: inst = 32'h10408000;
      30590: inst = 32'hc405279;
      30591: inst = 32'h8220000;
      30592: inst = 32'h10408000;
      30593: inst = 32'hc40527a;
      30594: inst = 32'h8220000;
      30595: inst = 32'h10408000;
      30596: inst = 32'hc40527b;
      30597: inst = 32'h8220000;
      30598: inst = 32'h10408000;
      30599: inst = 32'hc40527c;
      30600: inst = 32'h8220000;
      30601: inst = 32'h10408000;
      30602: inst = 32'hc40527d;
      30603: inst = 32'h8220000;
      30604: inst = 32'h10408000;
      30605: inst = 32'hc40527e;
      30606: inst = 32'h8220000;
      30607: inst = 32'h10408000;
      30608: inst = 32'hc40527f;
      30609: inst = 32'h8220000;
      30610: inst = 32'h10408000;
      30611: inst = 32'hc405280;
      30612: inst = 32'h8220000;
      30613: inst = 32'h10408000;
      30614: inst = 32'hc405281;
      30615: inst = 32'h8220000;
      30616: inst = 32'h10408000;
      30617: inst = 32'hc405282;
      30618: inst = 32'h8220000;
      30619: inst = 32'h10408000;
      30620: inst = 32'hc405283;
      30621: inst = 32'h8220000;
      30622: inst = 32'h10408000;
      30623: inst = 32'hc405284;
      30624: inst = 32'h8220000;
      30625: inst = 32'h10408000;
      30626: inst = 32'hc405285;
      30627: inst = 32'h8220000;
      30628: inst = 32'h10408000;
      30629: inst = 32'hc405286;
      30630: inst = 32'h8220000;
      30631: inst = 32'h10408000;
      30632: inst = 32'hc405287;
      30633: inst = 32'h8220000;
      30634: inst = 32'h10408000;
      30635: inst = 32'hc405288;
      30636: inst = 32'h8220000;
      30637: inst = 32'h10408000;
      30638: inst = 32'hc405289;
      30639: inst = 32'h8220000;
      30640: inst = 32'h10408000;
      30641: inst = 32'hc40528a;
      30642: inst = 32'h8220000;
      30643: inst = 32'h10408000;
      30644: inst = 32'hc40528b;
      30645: inst = 32'h8220000;
      30646: inst = 32'h10408000;
      30647: inst = 32'hc40528c;
      30648: inst = 32'h8220000;
      30649: inst = 32'h10408000;
      30650: inst = 32'hc40528d;
      30651: inst = 32'h8220000;
      30652: inst = 32'h10408000;
      30653: inst = 32'hc40528e;
      30654: inst = 32'h8220000;
      30655: inst = 32'h10408000;
      30656: inst = 32'hc40528f;
      30657: inst = 32'h8220000;
      30658: inst = 32'h10408000;
      30659: inst = 32'hc405290;
      30660: inst = 32'h8220000;
      30661: inst = 32'h10408000;
      30662: inst = 32'hc405291;
      30663: inst = 32'h8220000;
      30664: inst = 32'h10408000;
      30665: inst = 32'hc405292;
      30666: inst = 32'h8220000;
      30667: inst = 32'h10408000;
      30668: inst = 32'hc405293;
      30669: inst = 32'h8220000;
      30670: inst = 32'h10408000;
      30671: inst = 32'hc405294;
      30672: inst = 32'h8220000;
      30673: inst = 32'h10408000;
      30674: inst = 32'hc405295;
      30675: inst = 32'h8220000;
      30676: inst = 32'h10408000;
      30677: inst = 32'hc405296;
      30678: inst = 32'h8220000;
      30679: inst = 32'h10408000;
      30680: inst = 32'hc405297;
      30681: inst = 32'h8220000;
      30682: inst = 32'h10408000;
      30683: inst = 32'hc405298;
      30684: inst = 32'h8220000;
      30685: inst = 32'h10408000;
      30686: inst = 32'hc4052a7;
      30687: inst = 32'h8220000;
      30688: inst = 32'h10408000;
      30689: inst = 32'hc4052a8;
      30690: inst = 32'h8220000;
      30691: inst = 32'h10408000;
      30692: inst = 32'hc4052a9;
      30693: inst = 32'h8220000;
      30694: inst = 32'h10408000;
      30695: inst = 32'hc4052aa;
      30696: inst = 32'h8220000;
      30697: inst = 32'h10408000;
      30698: inst = 32'hc4052ab;
      30699: inst = 32'h8220000;
      30700: inst = 32'h10408000;
      30701: inst = 32'hc4052ac;
      30702: inst = 32'h8220000;
      30703: inst = 32'h10408000;
      30704: inst = 32'hc4052ad;
      30705: inst = 32'h8220000;
      30706: inst = 32'h10408000;
      30707: inst = 32'hc4052ae;
      30708: inst = 32'h8220000;
      30709: inst = 32'h10408000;
      30710: inst = 32'hc4052af;
      30711: inst = 32'h8220000;
      30712: inst = 32'h10408000;
      30713: inst = 32'hc4052b0;
      30714: inst = 32'h8220000;
      30715: inst = 32'h10408000;
      30716: inst = 32'hc4052b1;
      30717: inst = 32'h8220000;
      30718: inst = 32'h10408000;
      30719: inst = 32'hc4052b2;
      30720: inst = 32'h8220000;
      30721: inst = 32'h10408000;
      30722: inst = 32'hc4052b3;
      30723: inst = 32'h8220000;
      30724: inst = 32'h10408000;
      30725: inst = 32'hc4052b4;
      30726: inst = 32'h8220000;
      30727: inst = 32'h10408000;
      30728: inst = 32'hc4052b5;
      30729: inst = 32'h8220000;
      30730: inst = 32'h10408000;
      30731: inst = 32'hc4052b6;
      30732: inst = 32'h8220000;
      30733: inst = 32'h10408000;
      30734: inst = 32'hc4052b7;
      30735: inst = 32'h8220000;
      30736: inst = 32'h10408000;
      30737: inst = 32'hc4052b8;
      30738: inst = 32'h8220000;
      30739: inst = 32'h10408000;
      30740: inst = 32'hc4052b9;
      30741: inst = 32'h8220000;
      30742: inst = 32'h10408000;
      30743: inst = 32'hc4052ba;
      30744: inst = 32'h8220000;
      30745: inst = 32'h10408000;
      30746: inst = 32'hc4052bb;
      30747: inst = 32'h8220000;
      30748: inst = 32'h10408000;
      30749: inst = 32'hc4052bc;
      30750: inst = 32'h8220000;
      30751: inst = 32'h10408000;
      30752: inst = 32'hc4052bd;
      30753: inst = 32'h8220000;
      30754: inst = 32'h10408000;
      30755: inst = 32'hc4052be;
      30756: inst = 32'h8220000;
      30757: inst = 32'h10408000;
      30758: inst = 32'hc4052bf;
      30759: inst = 32'h8220000;
      30760: inst = 32'h10408000;
      30761: inst = 32'hc4052c0;
      30762: inst = 32'h8220000;
      30763: inst = 32'h10408000;
      30764: inst = 32'hc4052c1;
      30765: inst = 32'h8220000;
      30766: inst = 32'h10408000;
      30767: inst = 32'hc4052c2;
      30768: inst = 32'h8220000;
      30769: inst = 32'h10408000;
      30770: inst = 32'hc4052c3;
      30771: inst = 32'h8220000;
      30772: inst = 32'h10408000;
      30773: inst = 32'hc4052c4;
      30774: inst = 32'h8220000;
      30775: inst = 32'h10408000;
      30776: inst = 32'hc4052c5;
      30777: inst = 32'h8220000;
      30778: inst = 32'h10408000;
      30779: inst = 32'hc4052c6;
      30780: inst = 32'h8220000;
      30781: inst = 32'h10408000;
      30782: inst = 32'hc4052c7;
      30783: inst = 32'h8220000;
      30784: inst = 32'h10408000;
      30785: inst = 32'hc4052c8;
      30786: inst = 32'h8220000;
      30787: inst = 32'h10408000;
      30788: inst = 32'hc4052c9;
      30789: inst = 32'h8220000;
      30790: inst = 32'h10408000;
      30791: inst = 32'hc4052ca;
      30792: inst = 32'h8220000;
      30793: inst = 32'h10408000;
      30794: inst = 32'hc4052cb;
      30795: inst = 32'h8220000;
      30796: inst = 32'h10408000;
      30797: inst = 32'hc4052cc;
      30798: inst = 32'h8220000;
      30799: inst = 32'h10408000;
      30800: inst = 32'hc4052cd;
      30801: inst = 32'h8220000;
      30802: inst = 32'h10408000;
      30803: inst = 32'hc4052ce;
      30804: inst = 32'h8220000;
      30805: inst = 32'h10408000;
      30806: inst = 32'hc4052cf;
      30807: inst = 32'h8220000;
      30808: inst = 32'h10408000;
      30809: inst = 32'hc4052d0;
      30810: inst = 32'h8220000;
      30811: inst = 32'h10408000;
      30812: inst = 32'hc4052d1;
      30813: inst = 32'h8220000;
      30814: inst = 32'h10408000;
      30815: inst = 32'hc4052d2;
      30816: inst = 32'h8220000;
      30817: inst = 32'h10408000;
      30818: inst = 32'hc4052d3;
      30819: inst = 32'h8220000;
      30820: inst = 32'h10408000;
      30821: inst = 32'hc4052d4;
      30822: inst = 32'h8220000;
      30823: inst = 32'h10408000;
      30824: inst = 32'hc4052d5;
      30825: inst = 32'h8220000;
      30826: inst = 32'h10408000;
      30827: inst = 32'hc4052d6;
      30828: inst = 32'h8220000;
      30829: inst = 32'h10408000;
      30830: inst = 32'hc4052d7;
      30831: inst = 32'h8220000;
      30832: inst = 32'h10408000;
      30833: inst = 32'hc4052d8;
      30834: inst = 32'h8220000;
      30835: inst = 32'h10408000;
      30836: inst = 32'hc4052d9;
      30837: inst = 32'h8220000;
      30838: inst = 32'h10408000;
      30839: inst = 32'hc4052da;
      30840: inst = 32'h8220000;
      30841: inst = 32'h10408000;
      30842: inst = 32'hc4052db;
      30843: inst = 32'h8220000;
      30844: inst = 32'h10408000;
      30845: inst = 32'hc4052dc;
      30846: inst = 32'h8220000;
      30847: inst = 32'h10408000;
      30848: inst = 32'hc4052dd;
      30849: inst = 32'h8220000;
      30850: inst = 32'h10408000;
      30851: inst = 32'hc4052de;
      30852: inst = 32'h8220000;
      30853: inst = 32'h10408000;
      30854: inst = 32'hc4052df;
      30855: inst = 32'h8220000;
      30856: inst = 32'h10408000;
      30857: inst = 32'hc4052e0;
      30858: inst = 32'h8220000;
      30859: inst = 32'h10408000;
      30860: inst = 32'hc4052e1;
      30861: inst = 32'h8220000;
      30862: inst = 32'h10408000;
      30863: inst = 32'hc4052e2;
      30864: inst = 32'h8220000;
      30865: inst = 32'h10408000;
      30866: inst = 32'hc4052e3;
      30867: inst = 32'h8220000;
      30868: inst = 32'h10408000;
      30869: inst = 32'hc4052e4;
      30870: inst = 32'h8220000;
      30871: inst = 32'h10408000;
      30872: inst = 32'hc4052e5;
      30873: inst = 32'h8220000;
      30874: inst = 32'h10408000;
      30875: inst = 32'hc4052e6;
      30876: inst = 32'h8220000;
      30877: inst = 32'h10408000;
      30878: inst = 32'hc4052e7;
      30879: inst = 32'h8220000;
      30880: inst = 32'h10408000;
      30881: inst = 32'hc4052e8;
      30882: inst = 32'h8220000;
      30883: inst = 32'h10408000;
      30884: inst = 32'hc4052e9;
      30885: inst = 32'h8220000;
      30886: inst = 32'h10408000;
      30887: inst = 32'hc4052ea;
      30888: inst = 32'h8220000;
      30889: inst = 32'h10408000;
      30890: inst = 32'hc4052eb;
      30891: inst = 32'h8220000;
      30892: inst = 32'h10408000;
      30893: inst = 32'hc4052ec;
      30894: inst = 32'h8220000;
      30895: inst = 32'h10408000;
      30896: inst = 32'hc4052ed;
      30897: inst = 32'h8220000;
      30898: inst = 32'h10408000;
      30899: inst = 32'hc4052ee;
      30900: inst = 32'h8220000;
      30901: inst = 32'h10408000;
      30902: inst = 32'hc4052ef;
      30903: inst = 32'h8220000;
      30904: inst = 32'h10408000;
      30905: inst = 32'hc4052f0;
      30906: inst = 32'h8220000;
      30907: inst = 32'h10408000;
      30908: inst = 32'hc4052f1;
      30909: inst = 32'h8220000;
      30910: inst = 32'h10408000;
      30911: inst = 32'hc4052f2;
      30912: inst = 32'h8220000;
      30913: inst = 32'h10408000;
      30914: inst = 32'hc4052f3;
      30915: inst = 32'h8220000;
      30916: inst = 32'h10408000;
      30917: inst = 32'hc4052f4;
      30918: inst = 32'h8220000;
      30919: inst = 32'h10408000;
      30920: inst = 32'hc4052f5;
      30921: inst = 32'h8220000;
      30922: inst = 32'h10408000;
      30923: inst = 32'hc4052f6;
      30924: inst = 32'h8220000;
      30925: inst = 32'h10408000;
      30926: inst = 32'hc4052f7;
      30927: inst = 32'h8220000;
      30928: inst = 32'h10408000;
      30929: inst = 32'hc4052f8;
      30930: inst = 32'h8220000;
      30931: inst = 32'h10408000;
      30932: inst = 32'hc405307;
      30933: inst = 32'h8220000;
      30934: inst = 32'h10408000;
      30935: inst = 32'hc405308;
      30936: inst = 32'h8220000;
      30937: inst = 32'h10408000;
      30938: inst = 32'hc405309;
      30939: inst = 32'h8220000;
      30940: inst = 32'h10408000;
      30941: inst = 32'hc40530a;
      30942: inst = 32'h8220000;
      30943: inst = 32'h10408000;
      30944: inst = 32'hc40530b;
      30945: inst = 32'h8220000;
      30946: inst = 32'h10408000;
      30947: inst = 32'hc40530c;
      30948: inst = 32'h8220000;
      30949: inst = 32'h10408000;
      30950: inst = 32'hc40530d;
      30951: inst = 32'h8220000;
      30952: inst = 32'h10408000;
      30953: inst = 32'hc40530e;
      30954: inst = 32'h8220000;
      30955: inst = 32'h10408000;
      30956: inst = 32'hc40530f;
      30957: inst = 32'h8220000;
      30958: inst = 32'h10408000;
      30959: inst = 32'hc405310;
      30960: inst = 32'h8220000;
      30961: inst = 32'h10408000;
      30962: inst = 32'hc405311;
      30963: inst = 32'h8220000;
      30964: inst = 32'h10408000;
      30965: inst = 32'hc405312;
      30966: inst = 32'h8220000;
      30967: inst = 32'h10408000;
      30968: inst = 32'hc405313;
      30969: inst = 32'h8220000;
      30970: inst = 32'h10408000;
      30971: inst = 32'hc405314;
      30972: inst = 32'h8220000;
      30973: inst = 32'h10408000;
      30974: inst = 32'hc405315;
      30975: inst = 32'h8220000;
      30976: inst = 32'h10408000;
      30977: inst = 32'hc405316;
      30978: inst = 32'h8220000;
      30979: inst = 32'h10408000;
      30980: inst = 32'hc405317;
      30981: inst = 32'h8220000;
      30982: inst = 32'h10408000;
      30983: inst = 32'hc405318;
      30984: inst = 32'h8220000;
      30985: inst = 32'h10408000;
      30986: inst = 32'hc405319;
      30987: inst = 32'h8220000;
      30988: inst = 32'h10408000;
      30989: inst = 32'hc40531a;
      30990: inst = 32'h8220000;
      30991: inst = 32'h10408000;
      30992: inst = 32'hc40531b;
      30993: inst = 32'h8220000;
      30994: inst = 32'h10408000;
      30995: inst = 32'hc40531c;
      30996: inst = 32'h8220000;
      30997: inst = 32'h10408000;
      30998: inst = 32'hc40531d;
      30999: inst = 32'h8220000;
      31000: inst = 32'h10408000;
      31001: inst = 32'hc40531e;
      31002: inst = 32'h8220000;
      31003: inst = 32'h10408000;
      31004: inst = 32'hc40531f;
      31005: inst = 32'h8220000;
      31006: inst = 32'h10408000;
      31007: inst = 32'hc405320;
      31008: inst = 32'h8220000;
      31009: inst = 32'h10408000;
      31010: inst = 32'hc405321;
      31011: inst = 32'h8220000;
      31012: inst = 32'h10408000;
      31013: inst = 32'hc405322;
      31014: inst = 32'h8220000;
      31015: inst = 32'h10408000;
      31016: inst = 32'hc405323;
      31017: inst = 32'h8220000;
      31018: inst = 32'h10408000;
      31019: inst = 32'hc405324;
      31020: inst = 32'h8220000;
      31021: inst = 32'h10408000;
      31022: inst = 32'hc405325;
      31023: inst = 32'h8220000;
      31024: inst = 32'h10408000;
      31025: inst = 32'hc405326;
      31026: inst = 32'h8220000;
      31027: inst = 32'h10408000;
      31028: inst = 32'hc405327;
      31029: inst = 32'h8220000;
      31030: inst = 32'h10408000;
      31031: inst = 32'hc405328;
      31032: inst = 32'h8220000;
      31033: inst = 32'h10408000;
      31034: inst = 32'hc405329;
      31035: inst = 32'h8220000;
      31036: inst = 32'h10408000;
      31037: inst = 32'hc40532a;
      31038: inst = 32'h8220000;
      31039: inst = 32'h10408000;
      31040: inst = 32'hc40532b;
      31041: inst = 32'h8220000;
      31042: inst = 32'h10408000;
      31043: inst = 32'hc40532c;
      31044: inst = 32'h8220000;
      31045: inst = 32'h10408000;
      31046: inst = 32'hc40532d;
      31047: inst = 32'h8220000;
      31048: inst = 32'h10408000;
      31049: inst = 32'hc40532e;
      31050: inst = 32'h8220000;
      31051: inst = 32'h10408000;
      31052: inst = 32'hc40532f;
      31053: inst = 32'h8220000;
      31054: inst = 32'h10408000;
      31055: inst = 32'hc405330;
      31056: inst = 32'h8220000;
      31057: inst = 32'h10408000;
      31058: inst = 32'hc405331;
      31059: inst = 32'h8220000;
      31060: inst = 32'h10408000;
      31061: inst = 32'hc405332;
      31062: inst = 32'h8220000;
      31063: inst = 32'h10408000;
      31064: inst = 32'hc405333;
      31065: inst = 32'h8220000;
      31066: inst = 32'h10408000;
      31067: inst = 32'hc405334;
      31068: inst = 32'h8220000;
      31069: inst = 32'h10408000;
      31070: inst = 32'hc405335;
      31071: inst = 32'h8220000;
      31072: inst = 32'h10408000;
      31073: inst = 32'hc405336;
      31074: inst = 32'h8220000;
      31075: inst = 32'h10408000;
      31076: inst = 32'hc405337;
      31077: inst = 32'h8220000;
      31078: inst = 32'h10408000;
      31079: inst = 32'hc405338;
      31080: inst = 32'h8220000;
      31081: inst = 32'h10408000;
      31082: inst = 32'hc405339;
      31083: inst = 32'h8220000;
      31084: inst = 32'h10408000;
      31085: inst = 32'hc40533a;
      31086: inst = 32'h8220000;
      31087: inst = 32'h10408000;
      31088: inst = 32'hc40533b;
      31089: inst = 32'h8220000;
      31090: inst = 32'h10408000;
      31091: inst = 32'hc40533c;
      31092: inst = 32'h8220000;
      31093: inst = 32'h10408000;
      31094: inst = 32'hc40533d;
      31095: inst = 32'h8220000;
      31096: inst = 32'h10408000;
      31097: inst = 32'hc40533e;
      31098: inst = 32'h8220000;
      31099: inst = 32'h10408000;
      31100: inst = 32'hc40533f;
      31101: inst = 32'h8220000;
      31102: inst = 32'h10408000;
      31103: inst = 32'hc405340;
      31104: inst = 32'h8220000;
      31105: inst = 32'h10408000;
      31106: inst = 32'hc405341;
      31107: inst = 32'h8220000;
      31108: inst = 32'h10408000;
      31109: inst = 32'hc405342;
      31110: inst = 32'h8220000;
      31111: inst = 32'h10408000;
      31112: inst = 32'hc405343;
      31113: inst = 32'h8220000;
      31114: inst = 32'h10408000;
      31115: inst = 32'hc405344;
      31116: inst = 32'h8220000;
      31117: inst = 32'h10408000;
      31118: inst = 32'hc405345;
      31119: inst = 32'h8220000;
      31120: inst = 32'h10408000;
      31121: inst = 32'hc405346;
      31122: inst = 32'h8220000;
      31123: inst = 32'h10408000;
      31124: inst = 32'hc405347;
      31125: inst = 32'h8220000;
      31126: inst = 32'h10408000;
      31127: inst = 32'hc405348;
      31128: inst = 32'h8220000;
      31129: inst = 32'h10408000;
      31130: inst = 32'hc405349;
      31131: inst = 32'h8220000;
      31132: inst = 32'h10408000;
      31133: inst = 32'hc40534a;
      31134: inst = 32'h8220000;
      31135: inst = 32'h10408000;
      31136: inst = 32'hc40534b;
      31137: inst = 32'h8220000;
      31138: inst = 32'h10408000;
      31139: inst = 32'hc40534c;
      31140: inst = 32'h8220000;
      31141: inst = 32'h10408000;
      31142: inst = 32'hc40534d;
      31143: inst = 32'h8220000;
      31144: inst = 32'h10408000;
      31145: inst = 32'hc40534e;
      31146: inst = 32'h8220000;
      31147: inst = 32'h10408000;
      31148: inst = 32'hc40534f;
      31149: inst = 32'h8220000;
      31150: inst = 32'h10408000;
      31151: inst = 32'hc405350;
      31152: inst = 32'h8220000;
      31153: inst = 32'h10408000;
      31154: inst = 32'hc405351;
      31155: inst = 32'h8220000;
      31156: inst = 32'h10408000;
      31157: inst = 32'hc405352;
      31158: inst = 32'h8220000;
      31159: inst = 32'h10408000;
      31160: inst = 32'hc405353;
      31161: inst = 32'h8220000;
      31162: inst = 32'h10408000;
      31163: inst = 32'hc405354;
      31164: inst = 32'h8220000;
      31165: inst = 32'h10408000;
      31166: inst = 32'hc405355;
      31167: inst = 32'h8220000;
      31168: inst = 32'h10408000;
      31169: inst = 32'hc405356;
      31170: inst = 32'h8220000;
      31171: inst = 32'h10408000;
      31172: inst = 32'hc405357;
      31173: inst = 32'h8220000;
      31174: inst = 32'h10408000;
      31175: inst = 32'hc405358;
      31176: inst = 32'h8220000;
      31177: inst = 32'h10408000;
      31178: inst = 32'hc405367;
      31179: inst = 32'h8220000;
      31180: inst = 32'h10408000;
      31181: inst = 32'hc405368;
      31182: inst = 32'h8220000;
      31183: inst = 32'h10408000;
      31184: inst = 32'hc405369;
      31185: inst = 32'h8220000;
      31186: inst = 32'h10408000;
      31187: inst = 32'hc40536a;
      31188: inst = 32'h8220000;
      31189: inst = 32'h10408000;
      31190: inst = 32'hc40536b;
      31191: inst = 32'h8220000;
      31192: inst = 32'h10408000;
      31193: inst = 32'hc40536c;
      31194: inst = 32'h8220000;
      31195: inst = 32'h10408000;
      31196: inst = 32'hc40536d;
      31197: inst = 32'h8220000;
      31198: inst = 32'h10408000;
      31199: inst = 32'hc40536e;
      31200: inst = 32'h8220000;
      31201: inst = 32'h10408000;
      31202: inst = 32'hc40536f;
      31203: inst = 32'h8220000;
      31204: inst = 32'h10408000;
      31205: inst = 32'hc405370;
      31206: inst = 32'h8220000;
      31207: inst = 32'h10408000;
      31208: inst = 32'hc405371;
      31209: inst = 32'h8220000;
      31210: inst = 32'h10408000;
      31211: inst = 32'hc405372;
      31212: inst = 32'h8220000;
      31213: inst = 32'h10408000;
      31214: inst = 32'hc405373;
      31215: inst = 32'h8220000;
      31216: inst = 32'h10408000;
      31217: inst = 32'hc405374;
      31218: inst = 32'h8220000;
      31219: inst = 32'h10408000;
      31220: inst = 32'hc405375;
      31221: inst = 32'h8220000;
      31222: inst = 32'h10408000;
      31223: inst = 32'hc405376;
      31224: inst = 32'h8220000;
      31225: inst = 32'h10408000;
      31226: inst = 32'hc405377;
      31227: inst = 32'h8220000;
      31228: inst = 32'h10408000;
      31229: inst = 32'hc405378;
      31230: inst = 32'h8220000;
      31231: inst = 32'h10408000;
      31232: inst = 32'hc405379;
      31233: inst = 32'h8220000;
      31234: inst = 32'h10408000;
      31235: inst = 32'hc40537a;
      31236: inst = 32'h8220000;
      31237: inst = 32'h10408000;
      31238: inst = 32'hc40537b;
      31239: inst = 32'h8220000;
      31240: inst = 32'h10408000;
      31241: inst = 32'hc40537c;
      31242: inst = 32'h8220000;
      31243: inst = 32'h10408000;
      31244: inst = 32'hc40537d;
      31245: inst = 32'h8220000;
      31246: inst = 32'h10408000;
      31247: inst = 32'hc40537e;
      31248: inst = 32'h8220000;
      31249: inst = 32'h10408000;
      31250: inst = 32'hc40537f;
      31251: inst = 32'h8220000;
      31252: inst = 32'h10408000;
      31253: inst = 32'hc405380;
      31254: inst = 32'h8220000;
      31255: inst = 32'h10408000;
      31256: inst = 32'hc405381;
      31257: inst = 32'h8220000;
      31258: inst = 32'h10408000;
      31259: inst = 32'hc405382;
      31260: inst = 32'h8220000;
      31261: inst = 32'h10408000;
      31262: inst = 32'hc405383;
      31263: inst = 32'h8220000;
      31264: inst = 32'h10408000;
      31265: inst = 32'hc405384;
      31266: inst = 32'h8220000;
      31267: inst = 32'h10408000;
      31268: inst = 32'hc405385;
      31269: inst = 32'h8220000;
      31270: inst = 32'h10408000;
      31271: inst = 32'hc405386;
      31272: inst = 32'h8220000;
      31273: inst = 32'h10408000;
      31274: inst = 32'hc405387;
      31275: inst = 32'h8220000;
      31276: inst = 32'h10408000;
      31277: inst = 32'hc405388;
      31278: inst = 32'h8220000;
      31279: inst = 32'h10408000;
      31280: inst = 32'hc405389;
      31281: inst = 32'h8220000;
      31282: inst = 32'h10408000;
      31283: inst = 32'hc40538a;
      31284: inst = 32'h8220000;
      31285: inst = 32'h10408000;
      31286: inst = 32'hc40538b;
      31287: inst = 32'h8220000;
      31288: inst = 32'h10408000;
      31289: inst = 32'hc40538c;
      31290: inst = 32'h8220000;
      31291: inst = 32'h10408000;
      31292: inst = 32'hc40538d;
      31293: inst = 32'h8220000;
      31294: inst = 32'h10408000;
      31295: inst = 32'hc40538e;
      31296: inst = 32'h8220000;
      31297: inst = 32'h10408000;
      31298: inst = 32'hc40538f;
      31299: inst = 32'h8220000;
      31300: inst = 32'h10408000;
      31301: inst = 32'hc405390;
      31302: inst = 32'h8220000;
      31303: inst = 32'h10408000;
      31304: inst = 32'hc405391;
      31305: inst = 32'h8220000;
      31306: inst = 32'h10408000;
      31307: inst = 32'hc405392;
      31308: inst = 32'h8220000;
      31309: inst = 32'h10408000;
      31310: inst = 32'hc405393;
      31311: inst = 32'h8220000;
      31312: inst = 32'h10408000;
      31313: inst = 32'hc405394;
      31314: inst = 32'h8220000;
      31315: inst = 32'h10408000;
      31316: inst = 32'hc405395;
      31317: inst = 32'h8220000;
      31318: inst = 32'h10408000;
      31319: inst = 32'hc405396;
      31320: inst = 32'h8220000;
      31321: inst = 32'h10408000;
      31322: inst = 32'hc405397;
      31323: inst = 32'h8220000;
      31324: inst = 32'h10408000;
      31325: inst = 32'hc405398;
      31326: inst = 32'h8220000;
      31327: inst = 32'h10408000;
      31328: inst = 32'hc405399;
      31329: inst = 32'h8220000;
      31330: inst = 32'h10408000;
      31331: inst = 32'hc40539a;
      31332: inst = 32'h8220000;
      31333: inst = 32'h10408000;
      31334: inst = 32'hc40539b;
      31335: inst = 32'h8220000;
      31336: inst = 32'h10408000;
      31337: inst = 32'hc40539c;
      31338: inst = 32'h8220000;
      31339: inst = 32'h10408000;
      31340: inst = 32'hc40539d;
      31341: inst = 32'h8220000;
      31342: inst = 32'h10408000;
      31343: inst = 32'hc40539e;
      31344: inst = 32'h8220000;
      31345: inst = 32'h10408000;
      31346: inst = 32'hc40539f;
      31347: inst = 32'h8220000;
      31348: inst = 32'h10408000;
      31349: inst = 32'hc4053a0;
      31350: inst = 32'h8220000;
      31351: inst = 32'h10408000;
      31352: inst = 32'hc4053a1;
      31353: inst = 32'h8220000;
      31354: inst = 32'h10408000;
      31355: inst = 32'hc4053a2;
      31356: inst = 32'h8220000;
      31357: inst = 32'h10408000;
      31358: inst = 32'hc4053a3;
      31359: inst = 32'h8220000;
      31360: inst = 32'h10408000;
      31361: inst = 32'hc4053a4;
      31362: inst = 32'h8220000;
      31363: inst = 32'h10408000;
      31364: inst = 32'hc4053a5;
      31365: inst = 32'h8220000;
      31366: inst = 32'h10408000;
      31367: inst = 32'hc4053a6;
      31368: inst = 32'h8220000;
      31369: inst = 32'h10408000;
      31370: inst = 32'hc4053a7;
      31371: inst = 32'h8220000;
      31372: inst = 32'h10408000;
      31373: inst = 32'hc4053a8;
      31374: inst = 32'h8220000;
      31375: inst = 32'h10408000;
      31376: inst = 32'hc4053a9;
      31377: inst = 32'h8220000;
      31378: inst = 32'h10408000;
      31379: inst = 32'hc4053aa;
      31380: inst = 32'h8220000;
      31381: inst = 32'h10408000;
      31382: inst = 32'hc4053ab;
      31383: inst = 32'h8220000;
      31384: inst = 32'h10408000;
      31385: inst = 32'hc4053ac;
      31386: inst = 32'h8220000;
      31387: inst = 32'h10408000;
      31388: inst = 32'hc4053ad;
      31389: inst = 32'h8220000;
      31390: inst = 32'h10408000;
      31391: inst = 32'hc4053ae;
      31392: inst = 32'h8220000;
      31393: inst = 32'h10408000;
      31394: inst = 32'hc4053af;
      31395: inst = 32'h8220000;
      31396: inst = 32'h10408000;
      31397: inst = 32'hc4053b0;
      31398: inst = 32'h8220000;
      31399: inst = 32'h10408000;
      31400: inst = 32'hc4053b1;
      31401: inst = 32'h8220000;
      31402: inst = 32'h10408000;
      31403: inst = 32'hc4053b2;
      31404: inst = 32'h8220000;
      31405: inst = 32'h10408000;
      31406: inst = 32'hc4053b3;
      31407: inst = 32'h8220000;
      31408: inst = 32'h10408000;
      31409: inst = 32'hc4053b4;
      31410: inst = 32'h8220000;
      31411: inst = 32'h10408000;
      31412: inst = 32'hc4053b5;
      31413: inst = 32'h8220000;
      31414: inst = 32'h10408000;
      31415: inst = 32'hc4053b6;
      31416: inst = 32'h8220000;
      31417: inst = 32'h10408000;
      31418: inst = 32'hc4053b7;
      31419: inst = 32'h8220000;
      31420: inst = 32'h10408000;
      31421: inst = 32'hc4053b8;
      31422: inst = 32'h8220000;
      31423: inst = 32'h10408000;
      31424: inst = 32'hc4053c8;
      31425: inst = 32'h8220000;
      31426: inst = 32'h10408000;
      31427: inst = 32'hc4053c9;
      31428: inst = 32'h8220000;
      31429: inst = 32'h10408000;
      31430: inst = 32'hc4053ca;
      31431: inst = 32'h8220000;
      31432: inst = 32'h10408000;
      31433: inst = 32'hc4053cb;
      31434: inst = 32'h8220000;
      31435: inst = 32'h10408000;
      31436: inst = 32'hc4053cc;
      31437: inst = 32'h8220000;
      31438: inst = 32'h10408000;
      31439: inst = 32'hc4053cd;
      31440: inst = 32'h8220000;
      31441: inst = 32'h10408000;
      31442: inst = 32'hc4053ce;
      31443: inst = 32'h8220000;
      31444: inst = 32'h10408000;
      31445: inst = 32'hc4053cf;
      31446: inst = 32'h8220000;
      31447: inst = 32'h10408000;
      31448: inst = 32'hc4053d0;
      31449: inst = 32'h8220000;
      31450: inst = 32'h10408000;
      31451: inst = 32'hc4053d1;
      31452: inst = 32'h8220000;
      31453: inst = 32'h10408000;
      31454: inst = 32'hc4053d2;
      31455: inst = 32'h8220000;
      31456: inst = 32'h10408000;
      31457: inst = 32'hc4053d3;
      31458: inst = 32'h8220000;
      31459: inst = 32'h10408000;
      31460: inst = 32'hc4053d4;
      31461: inst = 32'h8220000;
      31462: inst = 32'h10408000;
      31463: inst = 32'hc4053d5;
      31464: inst = 32'h8220000;
      31465: inst = 32'h10408000;
      31466: inst = 32'hc4053d6;
      31467: inst = 32'h8220000;
      31468: inst = 32'h10408000;
      31469: inst = 32'hc4053d7;
      31470: inst = 32'h8220000;
      31471: inst = 32'h10408000;
      31472: inst = 32'hc4053d8;
      31473: inst = 32'h8220000;
      31474: inst = 32'h10408000;
      31475: inst = 32'hc4053d9;
      31476: inst = 32'h8220000;
      31477: inst = 32'h10408000;
      31478: inst = 32'hc4053da;
      31479: inst = 32'h8220000;
      31480: inst = 32'h10408000;
      31481: inst = 32'hc4053db;
      31482: inst = 32'h8220000;
      31483: inst = 32'h10408000;
      31484: inst = 32'hc4053dc;
      31485: inst = 32'h8220000;
      31486: inst = 32'h10408000;
      31487: inst = 32'hc4053dd;
      31488: inst = 32'h8220000;
      31489: inst = 32'h10408000;
      31490: inst = 32'hc4053de;
      31491: inst = 32'h8220000;
      31492: inst = 32'h10408000;
      31493: inst = 32'hc4053df;
      31494: inst = 32'h8220000;
      31495: inst = 32'h10408000;
      31496: inst = 32'hc4053e0;
      31497: inst = 32'h8220000;
      31498: inst = 32'h10408000;
      31499: inst = 32'hc4053e1;
      31500: inst = 32'h8220000;
      31501: inst = 32'h10408000;
      31502: inst = 32'hc4053e2;
      31503: inst = 32'h8220000;
      31504: inst = 32'h10408000;
      31505: inst = 32'hc4053e3;
      31506: inst = 32'h8220000;
      31507: inst = 32'h10408000;
      31508: inst = 32'hc4053e4;
      31509: inst = 32'h8220000;
      31510: inst = 32'h10408000;
      31511: inst = 32'hc4053e5;
      31512: inst = 32'h8220000;
      31513: inst = 32'h10408000;
      31514: inst = 32'hc4053e6;
      31515: inst = 32'h8220000;
      31516: inst = 32'h10408000;
      31517: inst = 32'hc4053e7;
      31518: inst = 32'h8220000;
      31519: inst = 32'h10408000;
      31520: inst = 32'hc4053e8;
      31521: inst = 32'h8220000;
      31522: inst = 32'h10408000;
      31523: inst = 32'hc4053e9;
      31524: inst = 32'h8220000;
      31525: inst = 32'h10408000;
      31526: inst = 32'hc4053ea;
      31527: inst = 32'h8220000;
      31528: inst = 32'h10408000;
      31529: inst = 32'hc4053eb;
      31530: inst = 32'h8220000;
      31531: inst = 32'h10408000;
      31532: inst = 32'hc4053ec;
      31533: inst = 32'h8220000;
      31534: inst = 32'h10408000;
      31535: inst = 32'hc4053ed;
      31536: inst = 32'h8220000;
      31537: inst = 32'h10408000;
      31538: inst = 32'hc4053ee;
      31539: inst = 32'h8220000;
      31540: inst = 32'h10408000;
      31541: inst = 32'hc4053ef;
      31542: inst = 32'h8220000;
      31543: inst = 32'h10408000;
      31544: inst = 32'hc4053f0;
      31545: inst = 32'h8220000;
      31546: inst = 32'h10408000;
      31547: inst = 32'hc4053f1;
      31548: inst = 32'h8220000;
      31549: inst = 32'h10408000;
      31550: inst = 32'hc4053f2;
      31551: inst = 32'h8220000;
      31552: inst = 32'h10408000;
      31553: inst = 32'hc4053f3;
      31554: inst = 32'h8220000;
      31555: inst = 32'h10408000;
      31556: inst = 32'hc4053f4;
      31557: inst = 32'h8220000;
      31558: inst = 32'h10408000;
      31559: inst = 32'hc4053f5;
      31560: inst = 32'h8220000;
      31561: inst = 32'h10408000;
      31562: inst = 32'hc4053f6;
      31563: inst = 32'h8220000;
      31564: inst = 32'h10408000;
      31565: inst = 32'hc4053f7;
      31566: inst = 32'h8220000;
      31567: inst = 32'h10408000;
      31568: inst = 32'hc4053f8;
      31569: inst = 32'h8220000;
      31570: inst = 32'h10408000;
      31571: inst = 32'hc4053f9;
      31572: inst = 32'h8220000;
      31573: inst = 32'h10408000;
      31574: inst = 32'hc4053fa;
      31575: inst = 32'h8220000;
      31576: inst = 32'h10408000;
      31577: inst = 32'hc4053fb;
      31578: inst = 32'h8220000;
      31579: inst = 32'h10408000;
      31580: inst = 32'hc4053fc;
      31581: inst = 32'h8220000;
      31582: inst = 32'h10408000;
      31583: inst = 32'hc4053fd;
      31584: inst = 32'h8220000;
      31585: inst = 32'h10408000;
      31586: inst = 32'hc4053fe;
      31587: inst = 32'h8220000;
      31588: inst = 32'h10408000;
      31589: inst = 32'hc4053ff;
      31590: inst = 32'h8220000;
      31591: inst = 32'h10408000;
      31592: inst = 32'hc405400;
      31593: inst = 32'h8220000;
      31594: inst = 32'h10408000;
      31595: inst = 32'hc405401;
      31596: inst = 32'h8220000;
      31597: inst = 32'h10408000;
      31598: inst = 32'hc405402;
      31599: inst = 32'h8220000;
      31600: inst = 32'h10408000;
      31601: inst = 32'hc405403;
      31602: inst = 32'h8220000;
      31603: inst = 32'h10408000;
      31604: inst = 32'hc405404;
      31605: inst = 32'h8220000;
      31606: inst = 32'h10408000;
      31607: inst = 32'hc405405;
      31608: inst = 32'h8220000;
      31609: inst = 32'h10408000;
      31610: inst = 32'hc405406;
      31611: inst = 32'h8220000;
      31612: inst = 32'h10408000;
      31613: inst = 32'hc405407;
      31614: inst = 32'h8220000;
      31615: inst = 32'h10408000;
      31616: inst = 32'hc405408;
      31617: inst = 32'h8220000;
      31618: inst = 32'h10408000;
      31619: inst = 32'hc405409;
      31620: inst = 32'h8220000;
      31621: inst = 32'h10408000;
      31622: inst = 32'hc40540a;
      31623: inst = 32'h8220000;
      31624: inst = 32'h10408000;
      31625: inst = 32'hc40540b;
      31626: inst = 32'h8220000;
      31627: inst = 32'h10408000;
      31628: inst = 32'hc40540c;
      31629: inst = 32'h8220000;
      31630: inst = 32'h10408000;
      31631: inst = 32'hc40540d;
      31632: inst = 32'h8220000;
      31633: inst = 32'h10408000;
      31634: inst = 32'hc40540e;
      31635: inst = 32'h8220000;
      31636: inst = 32'h10408000;
      31637: inst = 32'hc40540f;
      31638: inst = 32'h8220000;
      31639: inst = 32'h10408000;
      31640: inst = 32'hc405410;
      31641: inst = 32'h8220000;
      31642: inst = 32'h10408000;
      31643: inst = 32'hc405411;
      31644: inst = 32'h8220000;
      31645: inst = 32'h10408000;
      31646: inst = 32'hc405412;
      31647: inst = 32'h8220000;
      31648: inst = 32'h10408000;
      31649: inst = 32'hc405413;
      31650: inst = 32'h8220000;
      31651: inst = 32'h10408000;
      31652: inst = 32'hc405414;
      31653: inst = 32'h8220000;
      31654: inst = 32'h10408000;
      31655: inst = 32'hc405415;
      31656: inst = 32'h8220000;
      31657: inst = 32'h10408000;
      31658: inst = 32'hc405416;
      31659: inst = 32'h8220000;
      31660: inst = 32'h10408000;
      31661: inst = 32'hc405417;
      31662: inst = 32'h8220000;
      31663: inst = 32'hc20296c;
      31664: inst = 32'h10408000;
      31665: inst = 32'hc404406;
      31666: inst = 32'h8220000;
      31667: inst = 32'h10408000;
      31668: inst = 32'hc404459;
      31669: inst = 32'h8220000;
      31670: inst = 32'h10408000;
      31671: inst = 32'hc404466;
      31672: inst = 32'h8220000;
      31673: inst = 32'h10408000;
      31674: inst = 32'hc4044b9;
      31675: inst = 32'h8220000;
      31676: inst = 32'h10408000;
      31677: inst = 32'hc4044c6;
      31678: inst = 32'h8220000;
      31679: inst = 32'h10408000;
      31680: inst = 32'hc404519;
      31681: inst = 32'h8220000;
      31682: inst = 32'h10408000;
      31683: inst = 32'hc404526;
      31684: inst = 32'h8220000;
      31685: inst = 32'h10408000;
      31686: inst = 32'hc404579;
      31687: inst = 32'h8220000;
      31688: inst = 32'h10408000;
      31689: inst = 32'hc404586;
      31690: inst = 32'h8220000;
      31691: inst = 32'h10408000;
      31692: inst = 32'hc4045d9;
      31693: inst = 32'h8220000;
      31694: inst = 32'h10408000;
      31695: inst = 32'hc4045e6;
      31696: inst = 32'h8220000;
      31697: inst = 32'h10408000;
      31698: inst = 32'hc404639;
      31699: inst = 32'h8220000;
      31700: inst = 32'h10408000;
      31701: inst = 32'hc404646;
      31702: inst = 32'h8220000;
      31703: inst = 32'h10408000;
      31704: inst = 32'hc404699;
      31705: inst = 32'h8220000;
      31706: inst = 32'h10408000;
      31707: inst = 32'hc4046a6;
      31708: inst = 32'h8220000;
      31709: inst = 32'h10408000;
      31710: inst = 32'hc4046f9;
      31711: inst = 32'h8220000;
      31712: inst = 32'h10408000;
      31713: inst = 32'hc404706;
      31714: inst = 32'h8220000;
      31715: inst = 32'h10408000;
      31716: inst = 32'hc404759;
      31717: inst = 32'h8220000;
      31718: inst = 32'h10408000;
      31719: inst = 32'hc404766;
      31720: inst = 32'h8220000;
      31721: inst = 32'h10408000;
      31722: inst = 32'hc4047b9;
      31723: inst = 32'h8220000;
      31724: inst = 32'h10408000;
      31725: inst = 32'hc4047c6;
      31726: inst = 32'h8220000;
      31727: inst = 32'h10408000;
      31728: inst = 32'hc404819;
      31729: inst = 32'h8220000;
      31730: inst = 32'h10408000;
      31731: inst = 32'hc404826;
      31732: inst = 32'h8220000;
      31733: inst = 32'h10408000;
      31734: inst = 32'hc404879;
      31735: inst = 32'h8220000;
      31736: inst = 32'h10408000;
      31737: inst = 32'hc404886;
      31738: inst = 32'h8220000;
      31739: inst = 32'h10408000;
      31740: inst = 32'hc4048d9;
      31741: inst = 32'h8220000;
      31742: inst = 32'h10408000;
      31743: inst = 32'hc4048e6;
      31744: inst = 32'h8220000;
      31745: inst = 32'h10408000;
      31746: inst = 32'hc404939;
      31747: inst = 32'h8220000;
      31748: inst = 32'h10408000;
      31749: inst = 32'hc404946;
      31750: inst = 32'h8220000;
      31751: inst = 32'h10408000;
      31752: inst = 32'hc404999;
      31753: inst = 32'h8220000;
      31754: inst = 32'h10408000;
      31755: inst = 32'hc4049a6;
      31756: inst = 32'h8220000;
      31757: inst = 32'h10408000;
      31758: inst = 32'hc4049f9;
      31759: inst = 32'h8220000;
      31760: inst = 32'h10408000;
      31761: inst = 32'hc404a06;
      31762: inst = 32'h8220000;
      31763: inst = 32'h10408000;
      31764: inst = 32'hc404a59;
      31765: inst = 32'h8220000;
      31766: inst = 32'h10408000;
      31767: inst = 32'hc404a66;
      31768: inst = 32'h8220000;
      31769: inst = 32'h10408000;
      31770: inst = 32'hc404ab9;
      31771: inst = 32'h8220000;
      31772: inst = 32'h10408000;
      31773: inst = 32'hc404ac6;
      31774: inst = 32'h8220000;
      31775: inst = 32'h10408000;
      31776: inst = 32'hc404b19;
      31777: inst = 32'h8220000;
      31778: inst = 32'h10408000;
      31779: inst = 32'hc404b26;
      31780: inst = 32'h8220000;
      31781: inst = 32'h10408000;
      31782: inst = 32'hc404b79;
      31783: inst = 32'h8220000;
      31784: inst = 32'h10408000;
      31785: inst = 32'hc404b86;
      31786: inst = 32'h8220000;
      31787: inst = 32'h10408000;
      31788: inst = 32'hc404bd9;
      31789: inst = 32'h8220000;
      31790: inst = 32'h10408000;
      31791: inst = 32'hc404be6;
      31792: inst = 32'h8220000;
      31793: inst = 32'h10408000;
      31794: inst = 32'hc404c39;
      31795: inst = 32'h8220000;
      31796: inst = 32'h10408000;
      31797: inst = 32'hc404c46;
      31798: inst = 32'h8220000;
      31799: inst = 32'h10408000;
      31800: inst = 32'hc404c99;
      31801: inst = 32'h8220000;
      31802: inst = 32'h10408000;
      31803: inst = 32'hc404ca6;
      31804: inst = 32'h8220000;
      31805: inst = 32'h10408000;
      31806: inst = 32'hc404cf9;
      31807: inst = 32'h8220000;
      31808: inst = 32'h10408000;
      31809: inst = 32'hc404d06;
      31810: inst = 32'h8220000;
      31811: inst = 32'h10408000;
      31812: inst = 32'hc404d59;
      31813: inst = 32'h8220000;
      31814: inst = 32'h10408000;
      31815: inst = 32'hc404d66;
      31816: inst = 32'h8220000;
      31817: inst = 32'h10408000;
      31818: inst = 32'hc404db9;
      31819: inst = 32'h8220000;
      31820: inst = 32'h10408000;
      31821: inst = 32'hc404dc6;
      31822: inst = 32'h8220000;
      31823: inst = 32'h10408000;
      31824: inst = 32'hc404e19;
      31825: inst = 32'h8220000;
      31826: inst = 32'h10408000;
      31827: inst = 32'hc404e26;
      31828: inst = 32'h8220000;
      31829: inst = 32'h10408000;
      31830: inst = 32'hc404e79;
      31831: inst = 32'h8220000;
      31832: inst = 32'h10408000;
      31833: inst = 32'hc404e86;
      31834: inst = 32'h8220000;
      31835: inst = 32'h10408000;
      31836: inst = 32'hc404ed9;
      31837: inst = 32'h8220000;
      31838: inst = 32'h10408000;
      31839: inst = 32'hc404ee6;
      31840: inst = 32'h8220000;
      31841: inst = 32'h10408000;
      31842: inst = 32'hc404f39;
      31843: inst = 32'h8220000;
      31844: inst = 32'h10408000;
      31845: inst = 32'hc404f46;
      31846: inst = 32'h8220000;
      31847: inst = 32'h10408000;
      31848: inst = 32'hc404f99;
      31849: inst = 32'h8220000;
      31850: inst = 32'h10408000;
      31851: inst = 32'hc404fa6;
      31852: inst = 32'h8220000;
      31853: inst = 32'h10408000;
      31854: inst = 32'hc404ff9;
      31855: inst = 32'h8220000;
      31856: inst = 32'h10408000;
      31857: inst = 32'hc405006;
      31858: inst = 32'h8220000;
      31859: inst = 32'h10408000;
      31860: inst = 32'hc405059;
      31861: inst = 32'h8220000;
      31862: inst = 32'h10408000;
      31863: inst = 32'hc405066;
      31864: inst = 32'h8220000;
      31865: inst = 32'h10408000;
      31866: inst = 32'hc4050b9;
      31867: inst = 32'h8220000;
      31868: inst = 32'h10408000;
      31869: inst = 32'hc4050c6;
      31870: inst = 32'h8220000;
      31871: inst = 32'h10408000;
      31872: inst = 32'hc405119;
      31873: inst = 32'h8220000;
      31874: inst = 32'h10408000;
      31875: inst = 32'hc405126;
      31876: inst = 32'h8220000;
      31877: inst = 32'h10408000;
      31878: inst = 32'hc405179;
      31879: inst = 32'h8220000;
      31880: inst = 32'h10408000;
      31881: inst = 32'hc405186;
      31882: inst = 32'h8220000;
      31883: inst = 32'h10408000;
      31884: inst = 32'hc4051d9;
      31885: inst = 32'h8220000;
      31886: inst = 32'h10408000;
      31887: inst = 32'hc4051e6;
      31888: inst = 32'h8220000;
      31889: inst = 32'h10408000;
      31890: inst = 32'hc405239;
      31891: inst = 32'h8220000;
      31892: inst = 32'h10408000;
      31893: inst = 32'hc405246;
      31894: inst = 32'h8220000;
      31895: inst = 32'h10408000;
      31896: inst = 32'hc405299;
      31897: inst = 32'h8220000;
      31898: inst = 32'h10408000;
      31899: inst = 32'hc4052a6;
      31900: inst = 32'h8220000;
      31901: inst = 32'h10408000;
      31902: inst = 32'hc4052f9;
      31903: inst = 32'h8220000;
      31904: inst = 32'h10408000;
      31905: inst = 32'hc405306;
      31906: inst = 32'h8220000;
      31907: inst = 32'h10408000;
      31908: inst = 32'hc405359;
      31909: inst = 32'h8220000;
      31910: inst = 32'hc20738e;
      31911: inst = 32'h10408000;
      31912: inst = 32'hc40464e;
      31913: inst = 32'h8220000;
      31914: inst = 32'h10408000;
      31915: inst = 32'hc404690;
      31916: inst = 32'h8220000;
      31917: inst = 32'h10408000;
      31918: inst = 32'hc4046ae;
      31919: inst = 32'h8220000;
      31920: inst = 32'h10408000;
      31921: inst = 32'hc4046f0;
      31922: inst = 32'h8220000;
      31923: inst = 32'h10408000;
      31924: inst = 32'hc4047d3;
      31925: inst = 32'h8220000;
      31926: inst = 32'h10408000;
      31927: inst = 32'hc4047dd;
      31928: inst = 32'h8220000;
      31929: inst = 32'h10408000;
      31930: inst = 32'hc404800;
      31931: inst = 32'h8220000;
      31932: inst = 32'h10408000;
      31933: inst = 32'hc40483a;
      31934: inst = 32'h8220000;
      31935: inst = 32'h10408000;
      31936: inst = 32'hc40485d;
      31937: inst = 32'h8220000;
      31938: inst = 32'h10408000;
      31939: inst = 32'hc4049b8;
      31940: inst = 32'h8220000;
      31941: inst = 32'h10408000;
      31942: inst = 32'hc4049c7;
      31943: inst = 32'h8220000;
      31944: inst = 32'h10408000;
      31945: inst = 32'hc4049e5;
      31946: inst = 32'h8220000;
      31947: inst = 32'h10408000;
      31948: inst = 32'hc4049f0;
      31949: inst = 32'h8220000;
      31950: inst = 32'h10408000;
      31951: inst = 32'hc404cb1;
      31952: inst = 32'h8220000;
      31953: inst = 32'h10408000;
      31954: inst = 32'hc404cf2;
      31955: inst = 32'h8220000;
      31956: inst = 32'h10408000;
      31957: inst = 32'hc404dda;
      31958: inst = 32'h8220000;
      31959: inst = 32'h10408000;
      31960: inst = 32'hc404e5c;
      31961: inst = 32'h8220000;
      31962: inst = 32'h10408000;
      31963: inst = 32'hc404e6b;
      31964: inst = 32'h8220000;
      31965: inst = 32'h10408000;
      31966: inst = 32'hc404e96;
      31967: inst = 32'h8220000;
      31968: inst = 32'h10408000;
      31969: inst = 32'hc404eaf;
      31970: inst = 32'h8220000;
      31971: inst = 32'h10408000;
      31972: inst = 32'hc404fb6;
      31973: inst = 32'h8220000;
      31974: inst = 32'h10408000;
      31975: inst = 32'hc404fcf;
      31976: inst = 32'h8220000;
      31977: inst = 32'h10408000;
      31978: inst = 32'hc40501a;
      31979: inst = 32'h8220000;
      31980: inst = 32'hc20ad75;
      31981: inst = 32'h10408000;
      31982: inst = 32'hc40464f;
      31983: inst = 32'h8220000;
      31984: inst = 32'h10408000;
      31985: inst = 32'hc404692;
      31986: inst = 32'h8220000;
      31987: inst = 32'h10408000;
      31988: inst = 32'hc404809;
      31989: inst = 32'h8220000;
      31990: inst = 32'h10408000;
      31991: inst = 32'hc40483d;
      31992: inst = 32'h8220000;
      31993: inst = 32'h10408000;
      31994: inst = 32'hc404860;
      31995: inst = 32'h8220000;
      31996: inst = 32'h10408000;
      31997: inst = 32'hc404e58;
      31998: inst = 32'h8220000;
      31999: inst = 32'h10408000;
      32000: inst = 32'hc404e59;
      32001: inst = 32'h8220000;
      32002: inst = 32'h10408000;
      32003: inst = 32'hc404e67;
      32004: inst = 32'h8220000;
      32005: inst = 32'h10408000;
      32006: inst = 32'hc404e68;
      32007: inst = 32'h8220000;
      32008: inst = 32'h10408000;
      32009: inst = 32'hc404f19;
      32010: inst = 32'h8220000;
      32011: inst = 32'h10408000;
      32012: inst = 32'hc404f28;
      32013: inst = 32'h8220000;
      32014: inst = 32'h10408000;
      32015: inst = 32'hc404f4f;
      32016: inst = 32'h8220000;
      32017: inst = 32'h10408000;
      32018: inst = 32'hc404fc3;
      32019: inst = 32'h8220000;
      32020: inst = 32'h10408000;
      32021: inst = 32'hc404fcd;
      32022: inst = 32'h8220000;
      32023: inst = 32'h10408000;
      32024: inst = 32'hc404fe1;
      32025: inst = 32'h8220000;
      32026: inst = 32'h10408000;
      32027: inst = 32'hc404ff0;
      32028: inst = 32'h8220000;
      32029: inst = 32'h10408000;
      32030: inst = 32'hc40500e;
      32031: inst = 32'h8220000;
      32032: inst = 32'h10408000;
      32033: inst = 32'hc405054;
      32034: inst = 32'h8220000;
      32035: inst = 32'hc2031a6;
      32036: inst = 32'h10408000;
      32037: inst = 32'hc404650;
      32038: inst = 32'h8220000;
      32039: inst = 32'h10408000;
      32040: inst = 32'hc404772;
      32041: inst = 32'h8220000;
      32042: inst = 32'h10408000;
      32043: inst = 32'hc40477a;
      32044: inst = 32'h8220000;
      32045: inst = 32'h10408000;
      32046: inst = 32'hc40478b;
      32047: inst = 32'h8220000;
      32048: inst = 32'h10408000;
      32049: inst = 32'hc404793;
      32050: inst = 32'h8220000;
      32051: inst = 32'h10408000;
      32052: inst = 32'hc404795;
      32053: inst = 32'h8220000;
      32054: inst = 32'h10408000;
      32055: inst = 32'hc40479a;
      32056: inst = 32'h8220000;
      32057: inst = 32'h10408000;
      32058: inst = 32'hc40479d;
      32059: inst = 32'h8220000;
      32060: inst = 32'h10408000;
      32061: inst = 32'hc4047ae;
      32062: inst = 32'h8220000;
      32063: inst = 32'h10408000;
      32064: inst = 32'hc404847;
      32065: inst = 32'h8220000;
      32066: inst = 32'h10408000;
      32067: inst = 32'hc404971;
      32068: inst = 32'h8220000;
      32069: inst = 32'h10408000;
      32070: inst = 32'hc40498a;
      32071: inst = 32'h8220000;
      32072: inst = 32'h10408000;
      32073: inst = 32'hc404a10;
      32074: inst = 32'h8220000;
      32075: inst = 32'h10408000;
      32076: inst = 32'hc404a18;
      32077: inst = 32'h8220000;
      32078: inst = 32'h10408000;
      32079: inst = 32'hc404a35;
      32080: inst = 32'h8220000;
      32081: inst = 32'h10408000;
      32082: inst = 32'hc404a3b;
      32083: inst = 32'h8220000;
      32084: inst = 32'h10408000;
      32085: inst = 32'hc404a45;
      32086: inst = 32'h8220000;
      32087: inst = 32'h10408000;
      32088: inst = 32'hc404a50;
      32089: inst = 32'h8220000;
      32090: inst = 32'h10408000;
      32091: inst = 32'hc404d21;
      32092: inst = 32'h8220000;
      32093: inst = 32'h10408000;
      32094: inst = 32'hc404d2b;
      32095: inst = 32'h8220000;
      32096: inst = 32'h10408000;
      32097: inst = 32'hc404d3f;
      32098: inst = 32'h8220000;
      32099: inst = 32'h10408000;
      32100: inst = 32'hc404d44;
      32101: inst = 32'h8220000;
      32102: inst = 32'h10408000;
      32103: inst = 32'hc404dcc;
      32104: inst = 32'h8220000;
      32105: inst = 32'h10408000;
      32106: inst = 32'hc404dcf;
      32107: inst = 32'h8220000;
      32108: inst = 32'h10408000;
      32109: inst = 32'hc404dd6;
      32110: inst = 32'h8220000;
      32111: inst = 32'h10408000;
      32112: inst = 32'hc404def;
      32113: inst = 32'h8220000;
      32114: inst = 32'h10408000;
      32115: inst = 32'hc404e98;
      32116: inst = 32'h8220000;
      32117: inst = 32'h10408000;
      32118: inst = 32'hc404eb1;
      32119: inst = 32'h8220000;
      32120: inst = 32'h10408000;
      32121: inst = 32'hc404fac;
      32122: inst = 32'h8220000;
      32123: inst = 32'h10408000;
      32124: inst = 32'hc404fb8;
      32125: inst = 32'h8220000;
      32126: inst = 32'h10408000;
      32127: inst = 32'hc404fd1;
      32128: inst = 32'h8220000;
      32129: inst = 32'h10408000;
      32130: inst = 32'hc404fd3;
      32131: inst = 32'h8220000;
      32132: inst = 32'h10408000;
      32133: inst = 32'hc40506b;
      32134: inst = 32'h8220000;
      32135: inst = 32'h10408000;
      32136: inst = 32'hc405076;
      32137: inst = 32'h8220000;
      32138: inst = 32'h10408000;
      32139: inst = 32'hc405078;
      32140: inst = 32'h8220000;
      32141: inst = 32'h10408000;
      32142: inst = 32'hc405081;
      32143: inst = 32'h8220000;
      32144: inst = 32'h10408000;
      32145: inst = 32'hc40508b;
      32146: inst = 32'h8220000;
      32147: inst = 32'h10408000;
      32148: inst = 32'hc40508f;
      32149: inst = 32'h8220000;
      32150: inst = 32'h10408000;
      32151: inst = 32'hc405091;
      32152: inst = 32'h8220000;
      32153: inst = 32'h10408000;
      32154: inst = 32'hc40509f;
      32155: inst = 32'h8220000;
      32156: inst = 32'h10408000;
      32157: inst = 32'hc4050a4;
      32158: inst = 32'h8220000;
      32159: inst = 32'h10408000;
      32160: inst = 32'hc4050ad;
      32161: inst = 32'h8220000;
      32162: inst = 32'hc20a514;
      32163: inst = 32'h10408000;
      32164: inst = 32'hc404691;
      32165: inst = 32'h8220000;
      32166: inst = 32'h10408000;
      32167: inst = 32'hc4046f1;
      32168: inst = 32'h8220000;
      32169: inst = 32'h10408000;
      32170: inst = 32'hc404715;
      32171: inst = 32'h8220000;
      32172: inst = 32'h10408000;
      32173: inst = 32'hc404716;
      32174: inst = 32'h8220000;
      32175: inst = 32'h10408000;
      32176: inst = 32'hc404724;
      32177: inst = 32'h8220000;
      32178: inst = 32'h10408000;
      32179: inst = 32'hc404725;
      32180: inst = 32'h8220000;
      32181: inst = 32'h10408000;
      32182: inst = 32'hc404742;
      32183: inst = 32'h8220000;
      32184: inst = 32'h10408000;
      32185: inst = 32'hc404743;
      32186: inst = 32'h8220000;
      32187: inst = 32'h10408000;
      32188: inst = 32'hc404776;
      32189: inst = 32'h8220000;
      32190: inst = 32'h10408000;
      32191: inst = 32'hc404785;
      32192: inst = 32'h8220000;
      32193: inst = 32'h10408000;
      32194: inst = 32'hc4047a3;
      32195: inst = 32'h8220000;
      32196: inst = 32'h10408000;
      32197: inst = 32'hc4047d4;
      32198: inst = 32'h8220000;
      32199: inst = 32'h10408000;
      32200: inst = 32'hc4047d7;
      32201: inst = 32'h8220000;
      32202: inst = 32'h10408000;
      32203: inst = 32'hc4047db;
      32204: inst = 32'h8220000;
      32205: inst = 32'h10408000;
      32206: inst = 32'hc4047e3;
      32207: inst = 32'h8220000;
      32208: inst = 32'h10408000;
      32209: inst = 32'hc4047e6;
      32210: inst = 32'h8220000;
      32211: inst = 32'h10408000;
      32212: inst = 32'hc4047ea;
      32213: inst = 32'h8220000;
      32214: inst = 32'h10408000;
      32215: inst = 32'hc4047f4;
      32216: inst = 32'h8220000;
      32217: inst = 32'h10408000;
      32218: inst = 32'hc4047f9;
      32219: inst = 32'h8220000;
      32220: inst = 32'h10408000;
      32221: inst = 32'hc4047fe;
      32222: inst = 32'h8220000;
      32223: inst = 32'h10408000;
      32224: inst = 32'hc404801;
      32225: inst = 32'h8220000;
      32226: inst = 32'h10408000;
      32227: inst = 32'hc404804;
      32228: inst = 32'h8220000;
      32229: inst = 32'h10408000;
      32230: inst = 32'hc404806;
      32231: inst = 32'h8220000;
      32232: inst = 32'h10408000;
      32233: inst = 32'hc404808;
      32234: inst = 32'h8220000;
      32235: inst = 32'h10408000;
      32236: inst = 32'hc40480d;
      32237: inst = 32'h8220000;
      32238: inst = 32'h10408000;
      32239: inst = 32'hc404836;
      32240: inst = 32'h8220000;
      32241: inst = 32'h10408000;
      32242: inst = 32'hc40483c;
      32243: inst = 32'h8220000;
      32244: inst = 32'h10408000;
      32245: inst = 32'hc404845;
      32246: inst = 32'h8220000;
      32247: inst = 32'h10408000;
      32248: inst = 32'hc404856;
      32249: inst = 32'h8220000;
      32250: inst = 32'h10408000;
      32251: inst = 32'hc40485f;
      32252: inst = 32'h8220000;
      32253: inst = 32'h10408000;
      32254: inst = 32'hc404863;
      32255: inst = 32'h8220000;
      32256: inst = 32'h10408000;
      32257: inst = 32'hc40486a;
      32258: inst = 32'h8220000;
      32259: inst = 32'h10408000;
      32260: inst = 32'hc404896;
      32261: inst = 32'h8220000;
      32262: inst = 32'h10408000;
      32263: inst = 32'hc40489c;
      32264: inst = 32'h8220000;
      32265: inst = 32'h10408000;
      32266: inst = 32'hc4048a5;
      32267: inst = 32'h8220000;
      32268: inst = 32'h10408000;
      32269: inst = 32'hc4048bf;
      32270: inst = 32'h8220000;
      32271: inst = 32'h10408000;
      32272: inst = 32'hc4048c3;
      32273: inst = 32'h8220000;
      32274: inst = 32'h10408000;
      32275: inst = 32'hc4048f6;
      32276: inst = 32'h8220000;
      32277: inst = 32'h10408000;
      32278: inst = 32'hc4048fc;
      32279: inst = 32'h8220000;
      32280: inst = 32'h10408000;
      32281: inst = 32'hc404905;
      32282: inst = 32'h8220000;
      32283: inst = 32'h10408000;
      32284: inst = 32'hc40491f;
      32285: inst = 32'h8220000;
      32286: inst = 32'h10408000;
      32287: inst = 32'hc404923;
      32288: inst = 32'h8220000;
      32289: inst = 32'h10408000;
      32290: inst = 32'hc404956;
      32291: inst = 32'h8220000;
      32292: inst = 32'h10408000;
      32293: inst = 32'hc404958;
      32294: inst = 32'h8220000;
      32295: inst = 32'h10408000;
      32296: inst = 32'hc40495c;
      32297: inst = 32'h8220000;
      32298: inst = 32'h10408000;
      32299: inst = 32'hc404965;
      32300: inst = 32'h8220000;
      32301: inst = 32'h10408000;
      32302: inst = 32'hc404967;
      32303: inst = 32'h8220000;
      32304: inst = 32'h10408000;
      32305: inst = 32'hc404976;
      32306: inst = 32'h8220000;
      32307: inst = 32'h10408000;
      32308: inst = 32'hc40497f;
      32309: inst = 32'h8220000;
      32310: inst = 32'h10408000;
      32311: inst = 32'hc404983;
      32312: inst = 32'h8220000;
      32313: inst = 32'h10408000;
      32314: inst = 32'hc404985;
      32315: inst = 32'h8220000;
      32316: inst = 32'h10408000;
      32317: inst = 32'hc4049b1;
      32318: inst = 32'h8220000;
      32319: inst = 32'h10408000;
      32320: inst = 32'hc4049b5;
      32321: inst = 32'h8220000;
      32322: inst = 32'h10408000;
      32323: inst = 32'hc4049ba;
      32324: inst = 32'h8220000;
      32325: inst = 32'h10408000;
      32326: inst = 32'hc4049c4;
      32327: inst = 32'h8220000;
      32328: inst = 32'h10408000;
      32329: inst = 32'hc4049ca;
      32330: inst = 32'h8220000;
      32331: inst = 32'h10408000;
      32332: inst = 32'hc4049d4;
      32333: inst = 32'h8220000;
      32334: inst = 32'h10408000;
      32335: inst = 32'hc4049d9;
      32336: inst = 32'h8220000;
      32337: inst = 32'h10408000;
      32338: inst = 32'hc4049dd;
      32339: inst = 32'h8220000;
      32340: inst = 32'h10408000;
      32341: inst = 32'hc4049e2;
      32342: inst = 32'h8220000;
      32343: inst = 32'h10408000;
      32344: inst = 32'hc4049e6;
      32345: inst = 32'h8220000;
      32346: inst = 32'h10408000;
      32347: inst = 32'hc4049e8;
      32348: inst = 32'h8220000;
      32349: inst = 32'h10408000;
      32350: inst = 32'hc4049ed;
      32351: inst = 32'h8220000;
      32352: inst = 32'h10408000;
      32353: inst = 32'hc4049f1;
      32354: inst = 32'h8220000;
      32355: inst = 32'h10408000;
      32356: inst = 32'hc4049f3;
      32357: inst = 32'h8220000;
      32358: inst = 32'h10408000;
      32359: inst = 32'hc404cb0;
      32360: inst = 32'h8220000;
      32361: inst = 32'h10408000;
      32362: inst = 32'hc404cf1;
      32363: inst = 32'h8220000;
      32364: inst = 32'h10408000;
      32365: inst = 32'hc404d11;
      32366: inst = 32'h8220000;
      32367: inst = 32'h10408000;
      32368: inst = 32'hc404d52;
      32369: inst = 32'h8220000;
      32370: inst = 32'h10408000;
      32371: inst = 32'hc404d71;
      32372: inst = 32'h8220000;
      32373: inst = 32'h10408000;
      32374: inst = 32'hc404db2;
      32375: inst = 32'h8220000;
      32376: inst = 32'h10408000;
      32377: inst = 32'hc404dd1;
      32378: inst = 32'h8220000;
      32379: inst = 32'h10408000;
      32380: inst = 32'hc404e12;
      32381: inst = 32'h8220000;
      32382: inst = 32'h10408000;
      32383: inst = 32'hc404e2d;
      32384: inst = 32'h8220000;
      32385: inst = 32'h10408000;
      32386: inst = 32'hc404e34;
      32387: inst = 32'h8220000;
      32388: inst = 32'h10408000;
      32389: inst = 32'hc404e37;
      32390: inst = 32'h8220000;
      32391: inst = 32'h10408000;
      32392: inst = 32'hc404e39;
      32393: inst = 32'h8220000;
      32394: inst = 32'h10408000;
      32395: inst = 32'hc404e3b;
      32396: inst = 32'h8220000;
      32397: inst = 32'h10408000;
      32398: inst = 32'hc404e3d;
      32399: inst = 32'h8220000;
      32400: inst = 32'h10408000;
      32401: inst = 32'hc404e42;
      32402: inst = 32'h8220000;
      32403: inst = 32'h10408000;
      32404: inst = 32'hc404e4c;
      32405: inst = 32'h8220000;
      32406: inst = 32'h10408000;
      32407: inst = 32'hc404e50;
      32408: inst = 32'h8220000;
      32409: inst = 32'h10408000;
      32410: inst = 32'hc404e5a;
      32411: inst = 32'h8220000;
      32412: inst = 32'h10408000;
      32413: inst = 32'hc404e60;
      32414: inst = 32'h8220000;
      32415: inst = 32'h10408000;
      32416: inst = 32'hc404e65;
      32417: inst = 32'h8220000;
      32418: inst = 32'h10408000;
      32419: inst = 32'hc404e69;
      32420: inst = 32'h8220000;
      32421: inst = 32'h10408000;
      32422: inst = 32'hc404e6e;
      32423: inst = 32'h8220000;
      32424: inst = 32'h10408000;
      32425: inst = 32'hc404e70;
      32426: inst = 32'h8220000;
      32427: inst = 32'h10408000;
      32428: inst = 32'hc404e72;
      32429: inst = 32'h8220000;
      32430: inst = 32'h10408000;
      32431: inst = 32'hc404e75;
      32432: inst = 32'h8220000;
      32433: inst = 32'h10408000;
      32434: inst = 32'hc404e8b;
      32435: inst = 32'h8220000;
      32436: inst = 32'h10408000;
      32437: inst = 32'hc404e8c;
      32438: inst = 32'h8220000;
      32439: inst = 32'h10408000;
      32440: inst = 32'hc404e91;
      32441: inst = 32'h8220000;
      32442: inst = 32'h10408000;
      32443: inst = 32'hc404e9b;
      32444: inst = 32'h8220000;
      32445: inst = 32'h10408000;
      32446: inst = 32'hc404ea0;
      32447: inst = 32'h8220000;
      32448: inst = 32'h10408000;
      32449: inst = 32'hc404eaa;
      32450: inst = 32'h8220000;
      32451: inst = 32'h10408000;
      32452: inst = 32'hc404ebb;
      32453: inst = 32'h8220000;
      32454: inst = 32'h10408000;
      32455: inst = 32'hc404ebe;
      32456: inst = 32'h8220000;
      32457: inst = 32'h10408000;
      32458: inst = 32'hc404ec3;
      32459: inst = 32'h8220000;
      32460: inst = 32'h10408000;
      32461: inst = 32'hc404eca;
      32462: inst = 32'h8220000;
      32463: inst = 32'h10408000;
      32464: inst = 32'hc404ecd;
      32465: inst = 32'h8220000;
      32466: inst = 32'h10408000;
      32467: inst = 32'hc404ed2;
      32468: inst = 32'h8220000;
      32469: inst = 32'h10408000;
      32470: inst = 32'hc404ed3;
      32471: inst = 32'h8220000;
      32472: inst = 32'h10408000;
      32473: inst = 32'hc404ed4;
      32474: inst = 32'h8220000;
      32475: inst = 32'h10408000;
      32476: inst = 32'hc404ef1;
      32477: inst = 32'h8220000;
      32478: inst = 32'h10408000;
      32479: inst = 32'hc404efb;
      32480: inst = 32'h8220000;
      32481: inst = 32'h10408000;
      32482: inst = 32'hc404f00;
      32483: inst = 32'h8220000;
      32484: inst = 32'h10408000;
      32485: inst = 32'hc404f0a;
      32486: inst = 32'h8220000;
      32487: inst = 32'h10408000;
      32488: inst = 32'hc404f1e;
      32489: inst = 32'h8220000;
      32490: inst = 32'h10408000;
      32491: inst = 32'hc404f23;
      32492: inst = 32'h8220000;
      32493: inst = 32'h10408000;
      32494: inst = 32'hc404f4d;
      32495: inst = 32'h8220000;
      32496: inst = 32'h10408000;
      32497: inst = 32'hc404f51;
      32498: inst = 32'h8220000;
      32499: inst = 32'h10408000;
      32500: inst = 32'hc404f5b;
      32501: inst = 32'h8220000;
      32502: inst = 32'h10408000;
      32503: inst = 32'hc404f60;
      32504: inst = 32'h8220000;
      32505: inst = 32'h10408000;
      32506: inst = 32'hc404f6a;
      32507: inst = 32'h8220000;
      32508: inst = 32'h10408000;
      32509: inst = 32'hc404f7b;
      32510: inst = 32'h8220000;
      32511: inst = 32'h10408000;
      32512: inst = 32'hc404f7e;
      32513: inst = 32'h8220000;
      32514: inst = 32'h10408000;
      32515: inst = 32'hc404f83;
      32516: inst = 32'h8220000;
      32517: inst = 32'h10408000;
      32518: inst = 32'hc404f8a;
      32519: inst = 32'h8220000;
      32520: inst = 32'h10408000;
      32521: inst = 32'hc404f93;
      32522: inst = 32'h8220000;
      32523: inst = 32'h10408000;
      32524: inst = 32'hc404fb1;
      32525: inst = 32'h8220000;
      32526: inst = 32'h10408000;
      32527: inst = 32'hc404fbb;
      32528: inst = 32'h8220000;
      32529: inst = 32'h10408000;
      32530: inst = 32'hc404fbd;
      32531: inst = 32'h8220000;
      32532: inst = 32'h10408000;
      32533: inst = 32'hc404fc0;
      32534: inst = 32'h8220000;
      32535: inst = 32'h10408000;
      32536: inst = 32'hc404fca;
      32537: inst = 32'h8220000;
      32538: inst = 32'h10408000;
      32539: inst = 32'hc404fdb;
      32540: inst = 32'h8220000;
      32541: inst = 32'h10408000;
      32542: inst = 32'hc404fde;
      32543: inst = 32'h8220000;
      32544: inst = 32'h10408000;
      32545: inst = 32'hc404fe3;
      32546: inst = 32'h8220000;
      32547: inst = 32'h10408000;
      32548: inst = 32'hc404fea;
      32549: inst = 32'h8220000;
      32550: inst = 32'h10408000;
      32551: inst = 32'hc404ff2;
      32552: inst = 32'h8220000;
      32553: inst = 32'h10408000;
      32554: inst = 32'hc40500d;
      32555: inst = 32'h8220000;
      32556: inst = 32'h10408000;
      32557: inst = 32'hc40500f;
      32558: inst = 32'h8220000;
      32559: inst = 32'h10408000;
      32560: inst = 32'hc405013;
      32561: inst = 32'h8220000;
      32562: inst = 32'h10408000;
      32563: inst = 32'hc405017;
      32564: inst = 32'h8220000;
      32565: inst = 32'h10408000;
      32566: inst = 32'hc405023;
      32567: inst = 32'h8220000;
      32568: inst = 32'h10408000;
      32569: inst = 32'hc40502d;
      32570: inst = 32'h8220000;
      32571: inst = 32'h10408000;
      32572: inst = 32'hc405030;
      32573: inst = 32'h8220000;
      32574: inst = 32'h10408000;
      32575: inst = 32'hc40503a;
      32576: inst = 32'h8220000;
      32577: inst = 32'h10408000;
      32578: inst = 32'hc40503d;
      32579: inst = 32'h8220000;
      32580: inst = 32'h10408000;
      32581: inst = 32'hc405041;
      32582: inst = 32'h8220000;
      32583: inst = 32'h10408000;
      32584: inst = 32'hc405046;
      32585: inst = 32'h8220000;
      32586: inst = 32'h10408000;
      32587: inst = 32'hc405049;
      32588: inst = 32'h8220000;
      32589: inst = 32'h10408000;
      32590: inst = 32'hc40504c;
      32591: inst = 32'h8220000;
      32592: inst = 32'h10408000;
      32593: inst = 32'hc40504e;
      32594: inst = 32'h8220000;
      32595: inst = 32'hc20f7be;
      32596: inst = 32'h10408000;
      32597: inst = 32'hc4046af;
      32598: inst = 32'h8220000;
      32599: inst = 32'h10408000;
      32600: inst = 32'hc4046f2;
      32601: inst = 32'h8220000;
      32602: inst = 32'h10408000;
      32603: inst = 32'hc40470f;
      32604: inst = 32'h8220000;
      32605: inst = 32'h10408000;
      32606: inst = 32'hc404752;
      32607: inst = 32'h8220000;
      32608: inst = 32'h10408000;
      32609: inst = 32'hc40476f;
      32610: inst = 32'h8220000;
      32611: inst = 32'h10408000;
      32612: inst = 32'hc4047b2;
      32613: inst = 32'h8220000;
      32614: inst = 32'h10408000;
      32615: inst = 32'hc4047cf;
      32616: inst = 32'h8220000;
      32617: inst = 32'h10408000;
      32618: inst = 32'hc4047d9;
      32619: inst = 32'h8220000;
      32620: inst = 32'h10408000;
      32621: inst = 32'hc4047fc;
      32622: inst = 32'h8220000;
      32623: inst = 32'h10408000;
      32624: inst = 32'hc404807;
      32625: inst = 32'h8220000;
      32626: inst = 32'h10408000;
      32627: inst = 32'hc40480a;
      32628: inst = 32'h8220000;
      32629: inst = 32'h10408000;
      32630: inst = 32'hc404812;
      32631: inst = 32'h8220000;
      32632: inst = 32'h10408000;
      32633: inst = 32'hc40482f;
      32634: inst = 32'h8220000;
      32635: inst = 32'h10408000;
      32636: inst = 32'hc404839;
      32637: inst = 32'h8220000;
      32638: inst = 32'h10408000;
      32639: inst = 32'hc40485c;
      32640: inst = 32'h8220000;
      32641: inst = 32'h10408000;
      32642: inst = 32'hc404867;
      32643: inst = 32'h8220000;
      32644: inst = 32'h10408000;
      32645: inst = 32'hc404872;
      32646: inst = 32'h8220000;
      32647: inst = 32'h10408000;
      32648: inst = 32'hc40488f;
      32649: inst = 32'h8220000;
      32650: inst = 32'h10408000;
      32651: inst = 32'hc404893;
      32652: inst = 32'h8220000;
      32653: inst = 32'h10408000;
      32654: inst = 32'hc404899;
      32655: inst = 32'h8220000;
      32656: inst = 32'h10408000;
      32657: inst = 32'hc4048ac;
      32658: inst = 32'h8220000;
      32659: inst = 32'h10408000;
      32660: inst = 32'hc4048b2;
      32661: inst = 32'h8220000;
      32662: inst = 32'h10408000;
      32663: inst = 32'hc4048bb;
      32664: inst = 32'h8220000;
      32665: inst = 32'h10408000;
      32666: inst = 32'hc4048bc;
      32667: inst = 32'h8220000;
      32668: inst = 32'h10408000;
      32669: inst = 32'hc4048c7;
      32670: inst = 32'h8220000;
      32671: inst = 32'h10408000;
      32672: inst = 32'hc4048cf;
      32673: inst = 32'h8220000;
      32674: inst = 32'h10408000;
      32675: inst = 32'hc4048d2;
      32676: inst = 32'h8220000;
      32677: inst = 32'h10408000;
      32678: inst = 32'hc4048ef;
      32679: inst = 32'h8220000;
      32680: inst = 32'h10408000;
      32681: inst = 32'hc4048f3;
      32682: inst = 32'h8220000;
      32683: inst = 32'h10408000;
      32684: inst = 32'hc4048f9;
      32685: inst = 32'h8220000;
      32686: inst = 32'h10408000;
      32687: inst = 32'hc40490c;
      32688: inst = 32'h8220000;
      32689: inst = 32'h10408000;
      32690: inst = 32'hc404912;
      32691: inst = 32'h8220000;
      32692: inst = 32'h10408000;
      32693: inst = 32'hc40491b;
      32694: inst = 32'h8220000;
      32695: inst = 32'h10408000;
      32696: inst = 32'hc40491c;
      32697: inst = 32'h8220000;
      32698: inst = 32'h10408000;
      32699: inst = 32'hc404927;
      32700: inst = 32'h8220000;
      32701: inst = 32'h10408000;
      32702: inst = 32'hc40492f;
      32703: inst = 32'h8220000;
      32704: inst = 32'h10408000;
      32705: inst = 32'hc404932;
      32706: inst = 32'h8220000;
      32707: inst = 32'h10408000;
      32708: inst = 32'hc40494f;
      32709: inst = 32'h8220000;
      32710: inst = 32'h10408000;
      32711: inst = 32'hc404959;
      32712: inst = 32'h8220000;
      32713: inst = 32'h10408000;
      32714: inst = 32'hc404972;
      32715: inst = 32'h8220000;
      32716: inst = 32'h10408000;
      32717: inst = 32'hc40497c;
      32718: inst = 32'h8220000;
      32719: inst = 32'h10408000;
      32720: inst = 32'hc404987;
      32721: inst = 32'h8220000;
      32722: inst = 32'h10408000;
      32723: inst = 32'hc404992;
      32724: inst = 32'h8220000;
      32725: inst = 32'h10408000;
      32726: inst = 32'hc4049b9;
      32727: inst = 32'h8220000;
      32728: inst = 32'h10408000;
      32729: inst = 32'hc4049dc;
      32730: inst = 32'h8220000;
      32731: inst = 32'h10408000;
      32732: inst = 32'hc4049e7;
      32733: inst = 32'h8220000;
      32734: inst = 32'h10408000;
      32735: inst = 32'hc4049f2;
      32736: inst = 32'h8220000;
      32737: inst = 32'h10408000;
      32738: inst = 32'hc404e74;
      32739: inst = 32'h8220000;
      32740: inst = 32'h10408000;
      32741: inst = 32'hc404ef4;
      32742: inst = 32'h8220000;
      32743: inst = 32'h10408000;
      32744: inst = 32'hc404ef5;
      32745: inst = 32'h8220000;
      32746: inst = 32'h10408000;
      32747: inst = 32'hc404ef9;
      32748: inst = 32'h8220000;
      32749: inst = 32'h10408000;
      32750: inst = 32'hc404f0e;
      32751: inst = 32'h8220000;
      32752: inst = 32'h10408000;
      32753: inst = 32'hc404f12;
      32754: inst = 32'h8220000;
      32755: inst = 32'h10408000;
      32756: inst = 32'hc404f2c;
      32757: inst = 32'h8220000;
      32758: inst = 32'h10408000;
      32759: inst = 32'hc404f33;
      32760: inst = 32'h8220000;
      32761: inst = 32'h10408000;
      32762: inst = 32'hc404f54;
      32763: inst = 32'h8220000;
      32764: inst = 32'h10408000;
      32765: inst = 32'hc404f59;
      32766: inst = 32'h8220000;
      32767: inst = 32'h10408000;
      32768: inst = 32'hc404f72;
      32769: inst = 32'h8220000;
      32770: inst = 32'h10408000;
      32771: inst = 32'hc404f8c;
      32772: inst = 32'h8220000;
      32773: inst = 32'h10408000;
      32774: inst = 32'hc404fb4;
      32775: inst = 32'h8220000;
      32776: inst = 32'h10408000;
      32777: inst = 32'hc404fb9;
      32778: inst = 32'h8220000;
      32779: inst = 32'h10408000;
      32780: inst = 32'hc404fd2;
      32781: inst = 32'h8220000;
      32782: inst = 32'h10408000;
      32783: inst = 32'hc404fd8;
      32784: inst = 32'h8220000;
      32785: inst = 32'h10408000;
      32786: inst = 32'hc404fe7;
      32787: inst = 32'h8220000;
      32788: inst = 32'h10408000;
      32789: inst = 32'hc405014;
      32790: inst = 32'h8220000;
      32791: inst = 32'hc20630c;
      32792: inst = 32'h10408000;
      32793: inst = 32'hc4046b0;
      32794: inst = 32'h8220000;
      32795: inst = 32'h10408000;
      32796: inst = 32'hc404710;
      32797: inst = 32'h8220000;
      32798: inst = 32'h10408000;
      32799: inst = 32'hc404751;
      32800: inst = 32'h8220000;
      32801: inst = 32'h10408000;
      32802: inst = 32'hc404770;
      32803: inst = 32'h8220000;
      32804: inst = 32'h10408000;
      32805: inst = 32'hc404771;
      32806: inst = 32'h8220000;
      32807: inst = 32'h10408000;
      32808: inst = 32'hc404774;
      32809: inst = 32'h8220000;
      32810: inst = 32'h10408000;
      32811: inst = 32'hc404777;
      32812: inst = 32'h8220000;
      32813: inst = 32'h10408000;
      32814: inst = 32'hc40477b;
      32815: inst = 32'h8220000;
      32816: inst = 32'h10408000;
      32817: inst = 32'hc404783;
      32818: inst = 32'h8220000;
      32819: inst = 32'h10408000;
      32820: inst = 32'hc404786;
      32821: inst = 32'h8220000;
      32822: inst = 32'h10408000;
      32823: inst = 32'hc40478a;
      32824: inst = 32'h8220000;
      32825: inst = 32'h10408000;
      32826: inst = 32'hc404794;
      32827: inst = 32'h8220000;
      32828: inst = 32'h10408000;
      32829: inst = 32'hc404799;
      32830: inst = 32'h8220000;
      32831: inst = 32'h10408000;
      32832: inst = 32'hc40479e;
      32833: inst = 32'h8220000;
      32834: inst = 32'h10408000;
      32835: inst = 32'hc4047a1;
      32836: inst = 32'h8220000;
      32837: inst = 32'h10408000;
      32838: inst = 32'hc4047a4;
      32839: inst = 32'h8220000;
      32840: inst = 32'h10408000;
      32841: inst = 32'hc4047a6;
      32842: inst = 32'h8220000;
      32843: inst = 32'h10408000;
      32844: inst = 32'hc4047a9;
      32845: inst = 32'h8220000;
      32846: inst = 32'h10408000;
      32847: inst = 32'hc4047ad;
      32848: inst = 32'h8220000;
      32849: inst = 32'h10408000;
      32850: inst = 32'hc4047b1;
      32851: inst = 32'h8220000;
      32852: inst = 32'h10408000;
      32853: inst = 32'hc4047f6;
      32854: inst = 32'h8220000;
      32855: inst = 32'h10408000;
      32856: inst = 32'hc404811;
      32857: inst = 32'h8220000;
      32858: inst = 32'h10408000;
      32859: inst = 32'hc404853;
      32860: inst = 32'h8220000;
      32861: inst = 32'h10408000;
      32862: inst = 32'hc404866;
      32863: inst = 32'h8220000;
      32864: inst = 32'h10408000;
      32865: inst = 32'hc404871;
      32866: inst = 32'h8220000;
      32867: inst = 32'h10408000;
      32868: inst = 32'hc404890;
      32869: inst = 32'h8220000;
      32870: inst = 32'h10408000;
      32871: inst = 32'hc404892;
      32872: inst = 32'h8220000;
      32873: inst = 32'h10408000;
      32874: inst = 32'hc40489a;
      32875: inst = 32'h8220000;
      32876: inst = 32'h10408000;
      32877: inst = 32'hc4048ab;
      32878: inst = 32'h8220000;
      32879: inst = 32'h10408000;
      32880: inst = 32'hc4048b1;
      32881: inst = 32'h8220000;
      32882: inst = 32'h10408000;
      32883: inst = 32'hc4048ba;
      32884: inst = 32'h8220000;
      32885: inst = 32'h10408000;
      32886: inst = 32'hc4048bd;
      32887: inst = 32'h8220000;
      32888: inst = 32'h10408000;
      32889: inst = 32'hc4048c6;
      32890: inst = 32'h8220000;
      32891: inst = 32'h10408000;
      32892: inst = 32'hc4048ce;
      32893: inst = 32'h8220000;
      32894: inst = 32'h10408000;
      32895: inst = 32'hc4048d1;
      32896: inst = 32'h8220000;
      32897: inst = 32'h10408000;
      32898: inst = 32'hc4048f0;
      32899: inst = 32'h8220000;
      32900: inst = 32'h10408000;
      32901: inst = 32'hc4048f2;
      32902: inst = 32'h8220000;
      32903: inst = 32'h10408000;
      32904: inst = 32'hc4048fa;
      32905: inst = 32'h8220000;
      32906: inst = 32'h10408000;
      32907: inst = 32'hc40490b;
      32908: inst = 32'h8220000;
      32909: inst = 32'h10408000;
      32910: inst = 32'hc404911;
      32911: inst = 32'h8220000;
      32912: inst = 32'h10408000;
      32913: inst = 32'hc40491a;
      32914: inst = 32'h8220000;
      32915: inst = 32'h10408000;
      32916: inst = 32'hc40491d;
      32917: inst = 32'h8220000;
      32918: inst = 32'h10408000;
      32919: inst = 32'hc404926;
      32920: inst = 32'h8220000;
      32921: inst = 32'h10408000;
      32922: inst = 32'hc40492e;
      32923: inst = 32'h8220000;
      32924: inst = 32'h10408000;
      32925: inst = 32'hc404931;
      32926: inst = 32'h8220000;
      32927: inst = 32'h10408000;
      32928: inst = 32'hc404950;
      32929: inst = 32'h8220000;
      32930: inst = 32'h10408000;
      32931: inst = 32'hc40495a;
      32932: inst = 32'h8220000;
      32933: inst = 32'h10408000;
      32934: inst = 32'hc40497d;
      32935: inst = 32'h8220000;
      32936: inst = 32'h10408000;
      32937: inst = 32'hc404986;
      32938: inst = 32'h8220000;
      32939: inst = 32'h10408000;
      32940: inst = 32'hc404991;
      32941: inst = 32'h8220000;
      32942: inst = 32'h10408000;
      32943: inst = 32'hc404a11;
      32944: inst = 32'h8220000;
      32945: inst = 32'h10408000;
      32946: inst = 32'hc404a19;
      32947: inst = 32'h8220000;
      32948: inst = 32'h10408000;
      32949: inst = 32'hc404a1c;
      32950: inst = 32'h8220000;
      32951: inst = 32'h10408000;
      32952: inst = 32'hc404a1d;
      32953: inst = 32'h8220000;
      32954: inst = 32'h10408000;
      32955: inst = 32'hc404a2a;
      32956: inst = 32'h8220000;
      32957: inst = 32'h10408000;
      32958: inst = 32'hc404a34;
      32959: inst = 32'h8220000;
      32960: inst = 32'h10408000;
      32961: inst = 32'hc404a39;
      32962: inst = 32'h8220000;
      32963: inst = 32'h10408000;
      32964: inst = 32'hc404a3c;
      32965: inst = 32'h8220000;
      32966: inst = 32'h10408000;
      32967: inst = 32'hc404a3f;
      32968: inst = 32'h8220000;
      32969: inst = 32'h10408000;
      32970: inst = 32'hc404a40;
      32971: inst = 32'h8220000;
      32972: inst = 32'h10408000;
      32973: inst = 32'hc404a46;
      32974: inst = 32'h8220000;
      32975: inst = 32'h10408000;
      32976: inst = 32'hc404a47;
      32977: inst = 32'h8220000;
      32978: inst = 32'h10408000;
      32979: inst = 32'hc404a48;
      32980: inst = 32'h8220000;
      32981: inst = 32'h10408000;
      32982: inst = 32'hc404a4d;
      32983: inst = 32'h8220000;
      32984: inst = 32'h10408000;
      32985: inst = 32'hc404a51;
      32986: inst = 32'h8220000;
      32987: inst = 32'h10408000;
      32988: inst = 32'hc404a52;
      32989: inst = 32'h8220000;
      32990: inst = 32'h10408000;
      32991: inst = 32'hc404a53;
      32992: inst = 32'h8220000;
      32993: inst = 32'h10408000;
      32994: inst = 32'hc404d80;
      32995: inst = 32'h8220000;
      32996: inst = 32'h10408000;
      32997: inst = 32'hc404d8a;
      32998: inst = 32'h8220000;
      32999: inst = 32'h10408000;
      33000: inst = 32'hc404d9e;
      33001: inst = 32'h8220000;
      33002: inst = 32'h10408000;
      33003: inst = 32'hc404da3;
      33004: inst = 32'h8220000;
      33005: inst = 32'h10408000;
      33006: inst = 32'hc404dcd;
      33007: inst = 32'h8220000;
      33008: inst = 32'h10408000;
      33009: inst = 32'hc404dd2;
      33010: inst = 32'h8220000;
      33011: inst = 32'h10408000;
      33012: inst = 32'hc404dd3;
      33013: inst = 32'h8220000;
      33014: inst = 32'h10408000;
      33015: inst = 32'hc404dd7;
      33016: inst = 32'h8220000;
      33017: inst = 32'h10408000;
      33018: inst = 32'hc404dde;
      33019: inst = 32'h8220000;
      33020: inst = 32'h10408000;
      33021: inst = 32'hc404de2;
      33022: inst = 32'h8220000;
      33023: inst = 32'h10408000;
      33024: inst = 32'hc404dec;
      33025: inst = 32'h8220000;
      33026: inst = 32'h10408000;
      33027: inst = 32'hc404df0;
      33028: inst = 32'h8220000;
      33029: inst = 32'h10408000;
      33030: inst = 32'hc404dfa;
      33031: inst = 32'h8220000;
      33032: inst = 32'h10408000;
      33033: inst = 32'hc404e00;
      33034: inst = 32'h8220000;
      33035: inst = 32'h10408000;
      33036: inst = 32'hc404e05;
      33037: inst = 32'h8220000;
      33038: inst = 32'h10408000;
      33039: inst = 32'hc404e09;
      33040: inst = 32'h8220000;
      33041: inst = 32'h10408000;
      33042: inst = 32'hc404e0e;
      33043: inst = 32'h8220000;
      33044: inst = 32'h10408000;
      33045: inst = 32'hc404e14;
      33046: inst = 32'h8220000;
      33047: inst = 32'h10408000;
      33048: inst = 32'hc404e15;
      33049: inst = 32'h8220000;
      33050: inst = 32'h10408000;
      33051: inst = 32'hc404e93;
      33052: inst = 32'h8220000;
      33053: inst = 32'h10408000;
      33054: inst = 32'hc404e9d;
      33055: inst = 32'h8220000;
      33056: inst = 32'h10408000;
      33057: inst = 32'hc404eb9;
      33058: inst = 32'h8220000;
      33059: inst = 32'h10408000;
      33060: inst = 32'hc404ec8;
      33061: inst = 32'h8220000;
      33062: inst = 32'h10408000;
      33063: inst = 32'hc404ef3;
      33064: inst = 32'h8220000;
      33065: inst = 32'h10408000;
      33066: inst = 32'hc404efd;
      33067: inst = 32'h8220000;
      33068: inst = 32'h10408000;
      33069: inst = 32'hc404f13;
      33070: inst = 32'h8220000;
      33071: inst = 32'h10408000;
      33072: inst = 32'hc404f2d;
      33073: inst = 32'h8220000;
      33074: inst = 32'h10408000;
      33075: inst = 32'hc404f53;
      33076: inst = 32'h8220000;
      33077: inst = 32'h10408000;
      33078: inst = 32'hc404f5d;
      33079: inst = 32'h8220000;
      33080: inst = 32'h10408000;
      33081: inst = 32'hc404f73;
      33082: inst = 32'h8220000;
      33083: inst = 32'h10408000;
      33084: inst = 32'hc404f8d;
      33085: inst = 32'h8220000;
      33086: inst = 32'h10408000;
      33087: inst = 32'hc404fb3;
      33088: inst = 32'h8220000;
      33089: inst = 32'h10408000;
      33090: inst = 32'hc404fd7;
      33091: inst = 32'h8220000;
      33092: inst = 32'h10408000;
      33093: inst = 32'hc404fdd;
      33094: inst = 32'h8220000;
      33095: inst = 32'h10408000;
      33096: inst = 32'hc405020;
      33097: inst = 32'h8220000;
      33098: inst = 32'h10408000;
      33099: inst = 32'hc40502a;
      33100: inst = 32'h8220000;
      33101: inst = 32'h10408000;
      33102: inst = 32'hc40503e;
      33103: inst = 32'h8220000;
      33104: inst = 32'h10408000;
      33105: inst = 32'hc405043;
      33106: inst = 32'h8220000;
      33107: inst = 32'h10408000;
      33108: inst = 32'hc40506d;
      33109: inst = 32'h8220000;
      33110: inst = 32'h10408000;
      33111: inst = 32'hc405070;
      33112: inst = 32'h8220000;
      33113: inst = 32'h10408000;
      33114: inst = 32'hc405071;
      33115: inst = 32'h8220000;
      33116: inst = 32'h10408000;
      33117: inst = 32'hc405074;
      33118: inst = 32'h8220000;
      33119: inst = 32'h10408000;
      33120: inst = 32'hc405077;
      33121: inst = 32'h8220000;
      33122: inst = 32'h10408000;
      33123: inst = 32'hc40507c;
      33124: inst = 32'h8220000;
      33125: inst = 32'h10408000;
      33126: inst = 32'hc405082;
      33127: inst = 32'h8220000;
      33128: inst = 32'h10408000;
      33129: inst = 32'hc40508c;
      33130: inst = 32'h8220000;
      33131: inst = 32'h10408000;
      33132: inst = 32'hc405090;
      33133: inst = 32'h8220000;
      33134: inst = 32'h10408000;
      33135: inst = 32'hc405099;
      33136: inst = 32'h8220000;
      33137: inst = 32'h10408000;
      33138: inst = 32'hc40509c;
      33139: inst = 32'h8220000;
      33140: inst = 32'h10408000;
      33141: inst = 32'hc4050a0;
      33142: inst = 32'h8220000;
      33143: inst = 32'h10408000;
      33144: inst = 32'hc4050a5;
      33145: inst = 32'h8220000;
      33146: inst = 32'h10408000;
      33147: inst = 32'hc4050a8;
      33148: inst = 32'h8220000;
      33149: inst = 32'h10408000;
      33150: inst = 32'hc4050ab;
      33151: inst = 32'h8220000;
      33152: inst = 32'h10408000;
      33153: inst = 32'hc4050ae;
      33154: inst = 32'h8220000;
      33155: inst = 32'h10408000;
      33156: inst = 32'hc4050b1;
      33157: inst = 32'h8220000;
      33158: inst = 32'h10408000;
      33159: inst = 32'hc4050b2;
      33160: inst = 32'h8220000;
      33161: inst = 32'h10408000;
      33162: inst = 32'hc4050b5;
      33163: inst = 32'h8220000;
      33164: inst = 32'hc20defb;
      33165: inst = 32'h10408000;
      33166: inst = 32'hc404775;
      33167: inst = 32'h8220000;
      33168: inst = 32'h10408000;
      33169: inst = 32'hc404784;
      33170: inst = 32'h8220000;
      33171: inst = 32'h10408000;
      33172: inst = 32'hc4047a2;
      33173: inst = 32'h8220000;
      33174: inst = 32'h10408000;
      33175: inst = 32'hc4047d2;
      33176: inst = 32'h8220000;
      33177: inst = 32'h10408000;
      33178: inst = 32'hc4047d5;
      33179: inst = 32'h8220000;
      33180: inst = 32'h10408000;
      33181: inst = 32'hc4047e4;
      33182: inst = 32'h8220000;
      33183: inst = 32'h10408000;
      33184: inst = 32'hc4047eb;
      33185: inst = 32'h8220000;
      33186: inst = 32'h10408000;
      33187: inst = 32'hc4047fa;
      33188: inst = 32'h8220000;
      33189: inst = 32'h10408000;
      33190: inst = 32'hc404802;
      33191: inst = 32'h8220000;
      33192: inst = 32'h10408000;
      33193: inst = 32'hc40480e;
      33194: inst = 32'h8220000;
      33195: inst = 32'h10408000;
      33196: inst = 32'hc404833;
      33197: inst = 32'h8220000;
      33198: inst = 32'h10408000;
      33199: inst = 32'hc40496c;
      33200: inst = 32'h8220000;
      33201: inst = 32'h10408000;
      33202: inst = 32'hc40497b;
      33203: inst = 32'h8220000;
      33204: inst = 32'h10408000;
      33205: inst = 32'hc40498f;
      33206: inst = 32'h8220000;
      33207: inst = 32'h10408000;
      33208: inst = 32'hc4049af;
      33209: inst = 32'h8220000;
      33210: inst = 32'h10408000;
      33211: inst = 32'hc4049b6;
      33212: inst = 32'h8220000;
      33213: inst = 32'h10408000;
      33214: inst = 32'hc4049bd;
      33215: inst = 32'h8220000;
      33216: inst = 32'h10408000;
      33217: inst = 32'hc4049c5;
      33218: inst = 32'h8220000;
      33219: inst = 32'h10408000;
      33220: inst = 32'hc4049d3;
      33221: inst = 32'h8220000;
      33222: inst = 32'h10408000;
      33223: inst = 32'hc4049e0;
      33224: inst = 32'h8220000;
      33225: inst = 32'h10408000;
      33226: inst = 32'hc4049e3;
      33227: inst = 32'h8220000;
      33228: inst = 32'h10408000;
      33229: inst = 32'hc404d10;
      33230: inst = 32'h8220000;
      33231: inst = 32'h10408000;
      33232: inst = 32'hc404d51;
      33233: inst = 32'h8220000;
      33234: inst = 32'h10408000;
      33235: inst = 32'hc404e31;
      33236: inst = 32'h8220000;
      33237: inst = 32'h10408000;
      33238: inst = 32'hc404e3a;
      33239: inst = 32'h8220000;
      33240: inst = 32'h10408000;
      33241: inst = 32'hc404e41;
      33242: inst = 32'h8220000;
      33243: inst = 32'h10408000;
      33244: inst = 32'hc404e4b;
      33245: inst = 32'h8220000;
      33246: inst = 32'h10408000;
      33247: inst = 32'hc404e5f;
      33248: inst = 32'h8220000;
      33249: inst = 32'h10408000;
      33250: inst = 32'hc404e64;
      33251: inst = 32'h8220000;
      33252: inst = 32'h10408000;
      33253: inst = 32'hc404e94;
      33254: inst = 32'h8220000;
      33255: inst = 32'h10408000;
      33256: inst = 32'hc404e95;
      33257: inst = 32'h8220000;
      33258: inst = 32'h10408000;
      33259: inst = 32'hc404e99;
      33260: inst = 32'h8220000;
      33261: inst = 32'h10408000;
      33262: inst = 32'hc404eae;
      33263: inst = 32'h8220000;
      33264: inst = 32'h10408000;
      33265: inst = 32'hc404eb2;
      33266: inst = 32'h8220000;
      33267: inst = 32'h10408000;
      33268: inst = 32'hc404f4e;
      33269: inst = 32'h8220000;
      33270: inst = 32'h10408000;
      33271: inst = 32'hc404fb5;
      33272: inst = 32'h8220000;
      33273: inst = 32'h10408000;
      33274: inst = 32'hc404fce;
      33275: inst = 32'h8220000;
      33276: inst = 32'h10408000;
      33277: inst = 32'hc405010;
      33278: inst = 32'h8220000;
      33279: inst = 32'h10408000;
      33280: inst = 32'hc40504d;
      33281: inst = 32'h8220000;
      33282: inst = 32'h10408000;
      33283: inst = 32'hc405051;
      33284: inst = 32'h8220000;
      33285: inst = 32'hc208410;
      33286: inst = 32'h10408000;
      33287: inst = 32'hc404779;
      33288: inst = 32'h8220000;
      33289: inst = 32'h10408000;
      33290: inst = 32'hc40479c;
      33291: inst = 32'h8220000;
      33292: inst = 32'h10408000;
      33293: inst = 32'hc4047e8;
      33294: inst = 32'h8220000;
      33295: inst = 32'h10408000;
      33296: inst = 32'hc4047f2;
      33297: inst = 32'h8220000;
      33298: inst = 32'h10408000;
      33299: inst = 32'hc4047f7;
      33300: inst = 32'h8220000;
      33301: inst = 32'h10408000;
      33302: inst = 32'hc40480b;
      33303: inst = 32'h8220000;
      33304: inst = 32'h10408000;
      33305: inst = 32'hc404830;
      33306: inst = 32'h8220000;
      33307: inst = 32'h10408000;
      33308: inst = 32'hc40484b;
      33309: inst = 32'h8220000;
      33310: inst = 32'h10408000;
      33311: inst = 32'hc40485a;
      33312: inst = 32'h8220000;
      33313: inst = 32'h10408000;
      33314: inst = 32'hc40486e;
      33315: inst = 32'h8220000;
      33316: inst = 32'h10408000;
      33317: inst = 32'hc40496b;
      33318: inst = 32'h8220000;
      33319: inst = 32'h10408000;
      33320: inst = 32'hc40497a;
      33321: inst = 32'h8220000;
      33322: inst = 32'h10408000;
      33323: inst = 32'hc40498e;
      33324: inst = 32'h8220000;
      33325: inst = 32'h10408000;
      33326: inst = 32'hc4049c8;
      33327: inst = 32'h8220000;
      33328: inst = 32'h10408000;
      33329: inst = 32'hc4049d2;
      33330: inst = 32'h8220000;
      33331: inst = 32'h10408000;
      33332: inst = 32'hc4049d7;
      33333: inst = 32'h8220000;
      33334: inst = 32'h10408000;
      33335: inst = 32'hc4049eb;
      33336: inst = 32'h8220000;
      33337: inst = 32'h10408000;
      33338: inst = 32'hc404e52;
      33339: inst = 32'h8220000;
      33340: inst = 32'h10408000;
      33341: inst = 32'hc404eee;
      33342: inst = 32'h8220000;
      33343: inst = 32'h10408000;
      33344: inst = 32'hc404ff5;
      33345: inst = 32'h8220000;
      33346: inst = 32'h10408000;
      33347: inst = 32'hc405019;
      33348: inst = 32'h8220000;
      33349: inst = 32'h10408000;
      33350: inst = 32'hc40501f;
      33351: inst = 32'h8220000;
      33352: inst = 32'h10408000;
      33353: inst = 32'hc405032;
      33354: inst = 32'h8220000;
      33355: inst = 32'h10408000;
      33356: inst = 32'hc405050;
      33357: inst = 32'h8220000;
      33358: inst = 32'hc204a69;
      33359: inst = 32'h10408000;
      33360: inst = 32'hc40477c;
      33361: inst = 32'h8220000;
      33362: inst = 32'h10408000;
      33363: inst = 32'hc404789;
      33364: inst = 32'h8220000;
      33365: inst = 32'h10408000;
      33366: inst = 32'hc404798;
      33367: inst = 32'h8220000;
      33368: inst = 32'h10408000;
      33369: inst = 32'hc40479f;
      33370: inst = 32'h8220000;
      33371: inst = 32'h10408000;
      33372: inst = 32'hc4047aa;
      33373: inst = 32'h8220000;
      33374: inst = 32'h10408000;
      33375: inst = 32'hc4047ac;
      33376: inst = 32'h8220000;
      33377: inst = 32'h10408000;
      33378: inst = 32'hc4047d8;
      33379: inst = 32'h8220000;
      33380: inst = 32'h10408000;
      33381: inst = 32'hc4047ec;
      33382: inst = 32'h8220000;
      33383: inst = 32'h10408000;
      33384: inst = 32'hc4047fb;
      33385: inst = 32'h8220000;
      33386: inst = 32'h10408000;
      33387: inst = 32'hc404805;
      33388: inst = 32'h8220000;
      33389: inst = 32'h10408000;
      33390: inst = 32'hc40480f;
      33391: inst = 32'h8220000;
      33392: inst = 32'h10408000;
      33393: inst = 32'hc404973;
      33394: inst = 32'h8220000;
      33395: inst = 32'h10408000;
      33396: inst = 32'hc4049b3;
      33397: inst = 32'h8220000;
      33398: inst = 32'h10408000;
      33399: inst = 32'hc4049cc;
      33400: inst = 32'h8220000;
      33401: inst = 32'h10408000;
      33402: inst = 32'hc4049d6;
      33403: inst = 32'h8220000;
      33404: inst = 32'h10408000;
      33405: inst = 32'hc4049e9;
      33406: inst = 32'h8220000;
      33407: inst = 32'h10408000;
      33408: inst = 32'hc4049ef;
      33409: inst = 32'h8220000;
      33410: inst = 32'h10408000;
      33411: inst = 32'hc4049f4;
      33412: inst = 32'h8220000;
      33413: inst = 32'h10408000;
      33414: inst = 32'hc404a16;
      33415: inst = 32'h8220000;
      33416: inst = 32'h10408000;
      33417: inst = 32'hc404a17;
      33418: inst = 32'h8220000;
      33419: inst = 32'h10408000;
      33420: inst = 32'hc404a1a;
      33421: inst = 32'h8220000;
      33422: inst = 32'h10408000;
      33423: inst = 32'hc404a25;
      33424: inst = 32'h8220000;
      33425: inst = 32'h10408000;
      33426: inst = 32'hc404a26;
      33427: inst = 32'h8220000;
      33428: inst = 32'h10408000;
      33429: inst = 32'hc404a29;
      33430: inst = 32'h8220000;
      33431: inst = 32'h10408000;
      33432: inst = 32'hc404a33;
      33433: inst = 32'h8220000;
      33434: inst = 32'h10408000;
      33435: inst = 32'hc404a38;
      33436: inst = 32'h8220000;
      33437: inst = 32'h10408000;
      33438: inst = 32'hc404a3d;
      33439: inst = 32'h8220000;
      33440: inst = 32'h10408000;
      33441: inst = 32'hc404a43;
      33442: inst = 32'h8220000;
      33443: inst = 32'h10408000;
      33444: inst = 32'hc404a44;
      33445: inst = 32'h8220000;
      33446: inst = 32'h10408000;
      33447: inst = 32'hc404a4c;
      33448: inst = 32'h8220000;
      33449: inst = 32'h10408000;
      33450: inst = 32'hc404caf;
      33451: inst = 32'h8220000;
      33452: inst = 32'h10408000;
      33453: inst = 32'hc404cf0;
      33454: inst = 32'h8220000;
      33455: inst = 32'h10408000;
      33456: inst = 32'hc404d0f;
      33457: inst = 32'h8220000;
      33458: inst = 32'h10408000;
      33459: inst = 32'hc404d50;
      33460: inst = 32'h8220000;
      33461: inst = 32'h10408000;
      33462: inst = 32'hc404dce;
      33463: inst = 32'h8220000;
      33464: inst = 32'h10408000;
      33465: inst = 32'hc404dd8;
      33466: inst = 32'h8220000;
      33467: inst = 32'h10408000;
      33468: inst = 32'hc404ddb;
      33469: inst = 32'h8220000;
      33470: inst = 32'h10408000;
      33471: inst = 32'hc404ddd;
      33472: inst = 32'h8220000;
      33473: inst = 32'h10408000;
      33474: inst = 32'hc404ddf;
      33475: inst = 32'h8220000;
      33476: inst = 32'h10408000;
      33477: inst = 32'hc404de9;
      33478: inst = 32'h8220000;
      33479: inst = 32'h10408000;
      33480: inst = 32'hc404df1;
      33481: inst = 32'h8220000;
      33482: inst = 32'h10408000;
      33483: inst = 32'hc404df9;
      33484: inst = 32'h8220000;
      33485: inst = 32'h10408000;
      33486: inst = 32'hc404dfb;
      33487: inst = 32'h8220000;
      33488: inst = 32'h10408000;
      33489: inst = 32'hc404dfd;
      33490: inst = 32'h8220000;
      33491: inst = 32'h10408000;
      33492: inst = 32'hc404e02;
      33493: inst = 32'h8220000;
      33494: inst = 32'h10408000;
      33495: inst = 32'hc404e08;
      33496: inst = 32'h8220000;
      33497: inst = 32'h10408000;
      33498: inst = 32'hc404e0a;
      33499: inst = 32'h8220000;
      33500: inst = 32'h10408000;
      33501: inst = 32'hc404e0f;
      33502: inst = 32'h8220000;
      33503: inst = 32'h10408000;
      33504: inst = 32'hc404e2b;
      33505: inst = 32'h8220000;
      33506: inst = 32'h10408000;
      33507: inst = 32'hc404e35;
      33508: inst = 32'h8220000;
      33509: inst = 32'h10408000;
      33510: inst = 32'hc404e43;
      33511: inst = 32'h8220000;
      33512: inst = 32'h10408000;
      33513: inst = 32'hc404e4d;
      33514: inst = 32'h8220000;
      33515: inst = 32'h10408000;
      33516: inst = 32'hc404e4e;
      33517: inst = 32'h8220000;
      33518: inst = 32'h10408000;
      33519: inst = 32'hc404e61;
      33520: inst = 32'h8220000;
      33521: inst = 32'h10408000;
      33522: inst = 32'hc404e66;
      33523: inst = 32'h8220000;
      33524: inst = 32'h10408000;
      33525: inst = 32'hc404e6c;
      33526: inst = 32'h8220000;
      33527: inst = 32'h10408000;
      33528: inst = 32'hc404e73;
      33529: inst = 32'h8220000;
      33530: inst = 32'h10408000;
      33531: inst = 32'hc404eeb;
      33532: inst = 32'h8220000;
      33533: inst = 32'h10408000;
      33534: inst = 32'hc404f0d;
      33535: inst = 32'h8220000;
      33536: inst = 32'h10408000;
      33537: inst = 32'hc404f18;
      33538: inst = 32'h8220000;
      33539: inst = 32'h10408000;
      33540: inst = 32'hc404f27;
      33541: inst = 32'h8220000;
      33542: inst = 32'h10408000;
      33543: inst = 32'hc404f34;
      33544: inst = 32'h8220000;
      33545: inst = 32'h10408000;
      33546: inst = 32'hc404f6d;
      33547: inst = 32'h8220000;
      33548: inst = 32'h10408000;
      33549: inst = 32'hc405015;
      33550: inst = 32'h8220000;
      33551: inst = 32'h10408000;
      33552: inst = 32'hc40502e;
      33553: inst = 32'h8220000;
      33554: inst = 32'h10408000;
      33555: inst = 32'hc405056;
      33556: inst = 32'h8220000;
      33557: inst = 32'h10408000;
      33558: inst = 32'hc40506e;
      33559: inst = 32'h8220000;
      33560: inst = 32'h10408000;
      33561: inst = 32'hc405073;
      33562: inst = 32'h8220000;
      33563: inst = 32'h10408000;
      33564: inst = 32'hc40507b;
      33565: inst = 32'h8220000;
      33566: inst = 32'h10408000;
      33567: inst = 32'hc40509a;
      33568: inst = 32'h8220000;
      33569: inst = 32'h10408000;
      33570: inst = 32'hc4050a9;
      33571: inst = 32'h8220000;
      33572: inst = 32'h10408000;
      33573: inst = 32'hc4050af;
      33574: inst = 32'h8220000;
      33575: inst = 32'h10408000;
      33576: inst = 32'hc4050b4;
      33577: inst = 32'h8220000;
      33578: inst = 32'hc209492;
      33579: inst = 32'h10408000;
      33580: inst = 32'hc4047a7;
      33581: inst = 32'h8220000;
      33582: inst = 32'h10408000;
      33583: inst = 32'hc404832;
      33584: inst = 32'h8220000;
      33585: inst = 32'h10408000;
      33586: inst = 32'hc404868;
      33587: inst = 32'h8220000;
      33588: inst = 32'h10408000;
      33589: inst = 32'hc4048a7;
      33590: inst = 32'h8220000;
      33591: inst = 32'h10408000;
      33592: inst = 32'hc4048b6;
      33593: inst = 32'h8220000;
      33594: inst = 32'h10408000;
      33595: inst = 32'hc4048ca;
      33596: inst = 32'h8220000;
      33597: inst = 32'h10408000;
      33598: inst = 32'hc404907;
      33599: inst = 32'h8220000;
      33600: inst = 32'h10408000;
      33601: inst = 32'hc404916;
      33602: inst = 32'h8220000;
      33603: inst = 32'h10408000;
      33604: inst = 32'hc40492a;
      33605: inst = 32'h8220000;
      33606: inst = 32'h10408000;
      33607: inst = 32'hc404952;
      33608: inst = 32'h8220000;
      33609: inst = 32'h10408000;
      33610: inst = 32'hc4049db;
      33611: inst = 32'h8220000;
      33612: inst = 32'h10408000;
      33613: inst = 32'hc404e3f;
      33614: inst = 32'h8220000;
      33615: inst = 32'h10408000;
      33616: inst = 32'hc404e49;
      33617: inst = 32'h8220000;
      33618: inst = 32'h10408000;
      33619: inst = 32'hc404e5d;
      33620: inst = 32'h8220000;
      33621: inst = 32'h10408000;
      33622: inst = 32'hc404e62;
      33623: inst = 32'h8220000;
      33624: inst = 32'h10408000;
      33625: inst = 32'hc404ecf;
      33626: inst = 32'h8220000;
      33627: inst = 32'h10408000;
      33628: inst = 32'hc404f79;
      33629: inst = 32'h8220000;
      33630: inst = 32'h10408000;
      33631: inst = 32'hc404f88;
      33632: inst = 32'h8220000;
      33633: inst = 32'h10408000;
      33634: inst = 32'hc404fed;
      33635: inst = 32'h8220000;
      33636: inst = 32'hc20d69a;
      33637: inst = 32'h10408000;
      33638: inst = 32'hc4047d0;
      33639: inst = 32'h8220000;
      33640: inst = 32'h10408000;
      33641: inst = 32'hc4047da;
      33642: inst = 32'h8220000;
      33643: inst = 32'h10408000;
      33644: inst = 32'hc4047f5;
      33645: inst = 32'h8220000;
      33646: inst = 32'h10408000;
      33647: inst = 32'hc4047fd;
      33648: inst = 32'h8220000;
      33649: inst = 32'h10408000;
      33650: inst = 32'hc4048a8;
      33651: inst = 32'h8220000;
      33652: inst = 32'h10408000;
      33653: inst = 32'hc4048b7;
      33654: inst = 32'h8220000;
      33655: inst = 32'h10408000;
      33656: inst = 32'hc4048cb;
      33657: inst = 32'h8220000;
      33658: inst = 32'h10408000;
      33659: inst = 32'hc404953;
      33660: inst = 32'h8220000;
      33661: inst = 32'h10408000;
      33662: inst = 32'hc4049b2;
      33663: inst = 32'h8220000;
      33664: inst = 32'h10408000;
      33665: inst = 32'hc4049cb;
      33666: inst = 32'h8220000;
      33667: inst = 32'h10408000;
      33668: inst = 32'hc4049da;
      33669: inst = 32'h8220000;
      33670: inst = 32'h10408000;
      33671: inst = 32'hc4049ee;
      33672: inst = 32'h8220000;
      33673: inst = 32'h10408000;
      33674: inst = 32'hc404e33;
      33675: inst = 32'h8220000;
      33676: inst = 32'h10408000;
      33677: inst = 32'hc404e36;
      33678: inst = 32'h8220000;
      33679: inst = 32'h10408000;
      33680: inst = 32'hc404e38;
      33681: inst = 32'h8220000;
      33682: inst = 32'h10408000;
      33683: inst = 32'hc404e4f;
      33684: inst = 32'h8220000;
      33685: inst = 32'h10408000;
      33686: inst = 32'hc404e51;
      33687: inst = 32'h8220000;
      33688: inst = 32'h10408000;
      33689: inst = 32'hc404e5b;
      33690: inst = 32'h8220000;
      33691: inst = 32'h10408000;
      33692: inst = 32'hc404e6a;
      33693: inst = 32'h8220000;
      33694: inst = 32'h10408000;
      33695: inst = 32'hc404e6d;
      33696: inst = 32'h8220000;
      33697: inst = 32'h10408000;
      33698: inst = 32'hc404eed;
      33699: inst = 32'h8220000;
      33700: inst = 32'h10408000;
      33701: inst = 32'hc404efa;
      33702: inst = 32'h8220000;
      33703: inst = 32'h10408000;
      33704: inst = 32'hc404f1a;
      33705: inst = 32'h8220000;
      33706: inst = 32'h10408000;
      33707: inst = 32'hc404f1b;
      33708: inst = 32'h8220000;
      33709: inst = 32'h10408000;
      33710: inst = 32'hc404f29;
      33711: inst = 32'h8220000;
      33712: inst = 32'h10408000;
      33713: inst = 32'hc404f2a;
      33714: inst = 32'h8220000;
      33715: inst = 32'h10408000;
      33716: inst = 32'hc404f5a;
      33717: inst = 32'h8220000;
      33718: inst = 32'h10408000;
      33719: inst = 32'hc404fba;
      33720: inst = 32'h8220000;
      33721: inst = 32'h10408000;
      33722: inst = 32'hc404fe6;
      33723: inst = 32'h8220000;
      33724: inst = 32'h10408000;
      33725: inst = 32'hc40500c;
      33726: inst = 32'h8220000;
      33727: inst = 32'h10408000;
      33728: inst = 32'hc405038;
      33729: inst = 32'h8220000;
      33730: inst = 32'h10408000;
      33731: inst = 32'hc40503b;
      33732: inst = 32'h8220000;
      33733: inst = 32'h10408000;
      33734: inst = 32'hc405047;
      33735: inst = 32'h8220000;
      33736: inst = 32'h10408000;
      33737: inst = 32'hc40504a;
      33738: inst = 32'h8220000;
      33739: inst = 32'hc20bdd7;
      33740: inst = 32'h10408000;
      33741: inst = 32'hc4047d1;
      33742: inst = 32'h8220000;
      33743: inst = 32'h10408000;
      33744: inst = 32'hc4047d6;
      33745: inst = 32'h8220000;
      33746: inst = 32'h10408000;
      33747: inst = 32'hc4047e5;
      33748: inst = 32'h8220000;
      33749: inst = 32'h10408000;
      33750: inst = 32'hc404803;
      33751: inst = 32'h8220000;
      33752: inst = 32'h10408000;
      33753: inst = 32'hc404855;
      33754: inst = 32'h8220000;
      33755: inst = 32'h10408000;
      33756: inst = 32'hc4049c9;
      33757: inst = 32'h8220000;
      33758: inst = 32'h10408000;
      33759: inst = 32'hc4049d8;
      33760: inst = 32'h8220000;
      33761: inst = 32'h10408000;
      33762: inst = 32'hc4049ec;
      33763: inst = 32'h8220000;
      33764: inst = 32'h10408000;
      33765: inst = 32'hc404de0;
      33766: inst = 32'h8220000;
      33767: inst = 32'h10408000;
      33768: inst = 32'hc404dea;
      33769: inst = 32'h8220000;
      33770: inst = 32'h10408000;
      33771: inst = 32'hc404dfe;
      33772: inst = 32'h8220000;
      33773: inst = 32'h10408000;
      33774: inst = 32'hc404e03;
      33775: inst = 32'h8220000;
      33776: inst = 32'h10408000;
      33777: inst = 32'hc404e2c;
      33778: inst = 32'h8220000;
      33779: inst = 32'h10408000;
      33780: inst = 32'hc404e2e;
      33781: inst = 32'h8220000;
      33782: inst = 32'h10408000;
      33783: inst = 32'hc404e32;
      33784: inst = 32'h8220000;
      33785: inst = 32'h10408000;
      33786: inst = 32'hc404e40;
      33787: inst = 32'h8220000;
      33788: inst = 32'h10408000;
      33789: inst = 32'hc404e4a;
      33790: inst = 32'h8220000;
      33791: inst = 32'h10408000;
      33792: inst = 32'hc404e5e;
      33793: inst = 32'h8220000;
      33794: inst = 32'h10408000;
      33795: inst = 32'hc404e63;
      33796: inst = 32'h8220000;
      33797: inst = 32'h10408000;
      33798: inst = 32'hc404e6f;
      33799: inst = 32'h8220000;
      33800: inst = 32'h10408000;
      33801: inst = 32'hc404e8f;
      33802: inst = 32'h8220000;
      33803: inst = 32'h10408000;
      33804: inst = 32'hc404ed0;
      33805: inst = 32'h8220000;
      33806: inst = 32'h10408000;
      33807: inst = 32'hc404fab;
      33808: inst = 32'h8220000;
      33809: inst = 32'h10408000;
      33810: inst = 32'hc405039;
      33811: inst = 32'h8220000;
      33812: inst = 32'h10408000;
      33813: inst = 32'hc405048;
      33814: inst = 32'h8220000;
      33815: inst = 32'h10408000;
      33816: inst = 32'hc40504f;
      33817: inst = 32'h8220000;
      33818: inst = 32'hc20ef5d;
      33819: inst = 32'h10408000;
      33820: inst = 32'hc4047dc;
      33821: inst = 32'h8220000;
      33822: inst = 32'h10408000;
      33823: inst = 32'hc4047ff;
      33824: inst = 32'h8220000;
      33825: inst = 32'h10408000;
      33826: inst = 32'hc404848;
      33827: inst = 32'h8220000;
      33828: inst = 32'h10408000;
      33829: inst = 32'hc404852;
      33830: inst = 32'h8220000;
      33831: inst = 32'h10408000;
      33832: inst = 32'hc404857;
      33833: inst = 32'h8220000;
      33834: inst = 32'h10408000;
      33835: inst = 32'hc40486b;
      33836: inst = 32'h8220000;
      33837: inst = 32'h10408000;
      33838: inst = 32'hc404968;
      33839: inst = 32'h8220000;
      33840: inst = 32'h10408000;
      33841: inst = 32'hc404977;
      33842: inst = 32'h8220000;
      33843: inst = 32'h10408000;
      33844: inst = 32'hc40498b;
      33845: inst = 32'h8220000;
      33846: inst = 32'h10408000;
      33847: inst = 32'hc404eec;
      33848: inst = 32'h8220000;
      33849: inst = 32'h10408000;
      33850: inst = 32'hc404f55;
      33851: inst = 32'h8220000;
      33852: inst = 32'h10408000;
      33853: inst = 32'hc404f6e;
      33854: inst = 32'h8220000;
      33855: inst = 32'h10408000;
      33856: inst = 32'hc404f78;
      33857: inst = 32'h8220000;
      33858: inst = 32'h10408000;
      33859: inst = 32'hc404f87;
      33860: inst = 32'h8220000;
      33861: inst = 32'h10408000;
      33862: inst = 32'hc404faf;
      33863: inst = 32'h8220000;
      33864: inst = 32'h10408000;
      33865: inst = 32'hc404ff4;
      33866: inst = 32'h8220000;
      33867: inst = 32'h10408000;
      33868: inst = 32'hc40501b;
      33869: inst = 32'h8220000;
      33870: inst = 32'h10408000;
      33871: inst = 32'hc40501e;
      33872: inst = 32'h8220000;
      33873: inst = 32'h10408000;
      33874: inst = 32'hc405021;
      33875: inst = 32'h8220000;
      33876: inst = 32'h10408000;
      33877: inst = 32'hc40502b;
      33878: inst = 32'h8220000;
      33879: inst = 32'h10408000;
      33880: inst = 32'hc40503c;
      33881: inst = 32'h8220000;
      33882: inst = 32'h10408000;
      33883: inst = 32'hc40503f;
      33884: inst = 32'h8220000;
      33885: inst = 32'h10408000;
      33886: inst = 32'hc405044;
      33887: inst = 32'h8220000;
      33888: inst = 32'h10408000;
      33889: inst = 32'hc40504b;
      33890: inst = 32'h8220000;
      33891: inst = 32'h10408000;
      33892: inst = 32'hc405055;
      33893: inst = 32'h8220000;
      33894: inst = 32'hc20c638;
      33895: inst = 32'h10408000;
      33896: inst = 32'hc4047e9;
      33897: inst = 32'h8220000;
      33898: inst = 32'h10408000;
      33899: inst = 32'hc4047f3;
      33900: inst = 32'h8220000;
      33901: inst = 32'h10408000;
      33902: inst = 32'hc4047f8;
      33903: inst = 32'h8220000;
      33904: inst = 32'h10408000;
      33905: inst = 32'hc40480c;
      33906: inst = 32'h8220000;
      33907: inst = 32'h10408000;
      33908: inst = 32'hc404835;
      33909: inst = 32'h8220000;
      33910: inst = 32'h10408000;
      33911: inst = 32'hc404844;
      33912: inst = 32'h8220000;
      33913: inst = 32'h10408000;
      33914: inst = 32'hc40484c;
      33915: inst = 32'h8220000;
      33916: inst = 32'h10408000;
      33917: inst = 32'hc40485b;
      33918: inst = 32'h8220000;
      33919: inst = 32'h10408000;
      33920: inst = 32'hc404862;
      33921: inst = 32'h8220000;
      33922: inst = 32'h10408000;
      33923: inst = 32'hc40486f;
      33924: inst = 32'h8220000;
      33925: inst = 32'h10408000;
      33926: inst = 32'hc404895;
      33927: inst = 32'h8220000;
      33928: inst = 32'h10408000;
      33929: inst = 32'hc40489d;
      33930: inst = 32'h8220000;
      33931: inst = 32'h10408000;
      33932: inst = 32'hc4048a4;
      33933: inst = 32'h8220000;
      33934: inst = 32'h10408000;
      33935: inst = 32'hc4048c0;
      33936: inst = 32'h8220000;
      33937: inst = 32'h10408000;
      33938: inst = 32'hc4048c2;
      33939: inst = 32'h8220000;
      33940: inst = 32'h10408000;
      33941: inst = 32'hc4048f5;
      33942: inst = 32'h8220000;
      33943: inst = 32'h10408000;
      33944: inst = 32'hc4048fd;
      33945: inst = 32'h8220000;
      33946: inst = 32'h10408000;
      33947: inst = 32'hc404904;
      33948: inst = 32'h8220000;
      33949: inst = 32'h10408000;
      33950: inst = 32'hc404908;
      33951: inst = 32'h8220000;
      33952: inst = 32'h10408000;
      33953: inst = 32'hc404917;
      33954: inst = 32'h8220000;
      33955: inst = 32'h10408000;
      33956: inst = 32'hc404920;
      33957: inst = 32'h8220000;
      33958: inst = 32'h10408000;
      33959: inst = 32'hc404922;
      33960: inst = 32'h8220000;
      33961: inst = 32'h10408000;
      33962: inst = 32'hc40492b;
      33963: inst = 32'h8220000;
      33964: inst = 32'h10408000;
      33965: inst = 32'hc404955;
      33966: inst = 32'h8220000;
      33967: inst = 32'h10408000;
      33968: inst = 32'hc40495d;
      33969: inst = 32'h8220000;
      33970: inst = 32'h10408000;
      33971: inst = 32'hc404964;
      33972: inst = 32'h8220000;
      33973: inst = 32'h10408000;
      33974: inst = 32'hc404980;
      33975: inst = 32'h8220000;
      33976: inst = 32'h10408000;
      33977: inst = 32'hc404982;
      33978: inst = 32'h8220000;
      33979: inst = 32'h10408000;
      33980: inst = 32'hc4049b0;
      33981: inst = 32'h8220000;
      33982: inst = 32'h10408000;
      33983: inst = 32'hc4049b7;
      33984: inst = 32'h8220000;
      33985: inst = 32'h10408000;
      33986: inst = 32'hc4049bc;
      33987: inst = 32'h8220000;
      33988: inst = 32'h10408000;
      33989: inst = 32'hc4049c6;
      33990: inst = 32'h8220000;
      33991: inst = 32'h10408000;
      33992: inst = 32'hc4049d5;
      33993: inst = 32'h8220000;
      33994: inst = 32'h10408000;
      33995: inst = 32'hc4049df;
      33996: inst = 32'h8220000;
      33997: inst = 32'h10408000;
      33998: inst = 32'hc4049e4;
      33999: inst = 32'h8220000;
      34000: inst = 32'h10408000;
      34001: inst = 32'hc404d70;
      34002: inst = 32'h8220000;
      34003: inst = 32'h10408000;
      34004: inst = 32'hc404d81;
      34005: inst = 32'h8220000;
      34006: inst = 32'h10408000;
      34007: inst = 32'hc404d8b;
      34008: inst = 32'h8220000;
      34009: inst = 32'h10408000;
      34010: inst = 32'hc404d9f;
      34011: inst = 32'h8220000;
      34012: inst = 32'h10408000;
      34013: inst = 32'hc404da4;
      34014: inst = 32'h8220000;
      34015: inst = 32'h10408000;
      34016: inst = 32'hc404db1;
      34017: inst = 32'h8220000;
      34018: inst = 32'h10408000;
      34019: inst = 32'hc404dd0;
      34020: inst = 32'h8220000;
      34021: inst = 32'h10408000;
      34022: inst = 32'hc404de1;
      34023: inst = 32'h8220000;
      34024: inst = 32'h10408000;
      34025: inst = 32'hc404deb;
      34026: inst = 32'h8220000;
      34027: inst = 32'h10408000;
      34028: inst = 32'hc404dff;
      34029: inst = 32'h8220000;
      34030: inst = 32'h10408000;
      34031: inst = 32'hc404e04;
      34032: inst = 32'h8220000;
      34033: inst = 32'h10408000;
      34034: inst = 32'hc404e11;
      34035: inst = 32'h8220000;
      34036: inst = 32'h10408000;
      34037: inst = 32'hc404e2f;
      34038: inst = 32'h8220000;
      34039: inst = 32'h10408000;
      34040: inst = 32'hc404e30;
      34041: inst = 32'h8220000;
      34042: inst = 32'h10408000;
      34043: inst = 32'hc404e3e;
      34044: inst = 32'h8220000;
      34045: inst = 32'h10408000;
      34046: inst = 32'hc404e71;
      34047: inst = 32'h8220000;
      34048: inst = 32'h10408000;
      34049: inst = 32'hc404e90;
      34050: inst = 32'h8220000;
      34051: inst = 32'h10408000;
      34052: inst = 32'hc404e9a;
      34053: inst = 32'h8220000;
      34054: inst = 32'h10408000;
      34055: inst = 32'hc404e9e;
      34056: inst = 32'h8220000;
      34057: inst = 32'h10408000;
      34058: inst = 32'hc404ea1;
      34059: inst = 32'h8220000;
      34060: inst = 32'h10408000;
      34061: inst = 32'hc404eab;
      34062: inst = 32'h8220000;
      34063: inst = 32'h10408000;
      34064: inst = 32'hc404eb8;
      34065: inst = 32'h8220000;
      34066: inst = 32'h10408000;
      34067: inst = 32'hc404ebc;
      34068: inst = 32'h8220000;
      34069: inst = 32'h10408000;
      34070: inst = 32'hc404ebf;
      34071: inst = 32'h8220000;
      34072: inst = 32'h10408000;
      34073: inst = 32'hc404ec4;
      34074: inst = 32'h8220000;
      34075: inst = 32'h10408000;
      34076: inst = 32'hc404ec7;
      34077: inst = 32'h8220000;
      34078: inst = 32'h10408000;
      34079: inst = 32'hc404ecb;
      34080: inst = 32'h8220000;
      34081: inst = 32'h10408000;
      34082: inst = 32'hc404ecc;
      34083: inst = 32'h8220000;
      34084: inst = 32'h10408000;
      34085: inst = 32'hc404ed1;
      34086: inst = 32'h8220000;
      34087: inst = 32'h10408000;
      34088: inst = 32'hc404ef0;
      34089: inst = 32'h8220000;
      34090: inst = 32'h10408000;
      34091: inst = 32'hc404efe;
      34092: inst = 32'h8220000;
      34093: inst = 32'h10408000;
      34094: inst = 32'hc404f01;
      34095: inst = 32'h8220000;
      34096: inst = 32'h10408000;
      34097: inst = 32'hc404f0b;
      34098: inst = 32'h8220000;
      34099: inst = 32'h10408000;
      34100: inst = 32'hc404f1c;
      34101: inst = 32'h8220000;
      34102: inst = 32'h10408000;
      34103: inst = 32'hc404f1f;
      34104: inst = 32'h8220000;
      34105: inst = 32'h10408000;
      34106: inst = 32'hc404f24;
      34107: inst = 32'h8220000;
      34108: inst = 32'h10408000;
      34109: inst = 32'hc404f2b;
      34110: inst = 32'h8220000;
      34111: inst = 32'h10408000;
      34112: inst = 32'hc404f31;
      34113: inst = 32'h8220000;
      34114: inst = 32'h10408000;
      34115: inst = 32'hc404f32;
      34116: inst = 32'h8220000;
      34117: inst = 32'h10408000;
      34118: inst = 32'hc404f50;
      34119: inst = 32'h8220000;
      34120: inst = 32'h10408000;
      34121: inst = 32'hc404f5e;
      34122: inst = 32'h8220000;
      34123: inst = 32'h10408000;
      34124: inst = 32'hc404f61;
      34125: inst = 32'h8220000;
      34126: inst = 32'h10408000;
      34127: inst = 32'hc404f6b;
      34128: inst = 32'h8220000;
      34129: inst = 32'h10408000;
      34130: inst = 32'hc404f7c;
      34131: inst = 32'h8220000;
      34132: inst = 32'h10408000;
      34133: inst = 32'hc404f7f;
      34134: inst = 32'h8220000;
      34135: inst = 32'h10408000;
      34136: inst = 32'hc404f84;
      34137: inst = 32'h8220000;
      34138: inst = 32'h10408000;
      34139: inst = 32'hc404f8b;
      34140: inst = 32'h8220000;
      34141: inst = 32'h10408000;
      34142: inst = 32'hc404f91;
      34143: inst = 32'h8220000;
      34144: inst = 32'h10408000;
      34145: inst = 32'hc404f92;
      34146: inst = 32'h8220000;
      34147: inst = 32'h10408000;
      34148: inst = 32'hc404f94;
      34149: inst = 32'h8220000;
      34150: inst = 32'h10408000;
      34151: inst = 32'hc404fb0;
      34152: inst = 32'h8220000;
      34153: inst = 32'h10408000;
      34154: inst = 32'hc404fbe;
      34155: inst = 32'h8220000;
      34156: inst = 32'h10408000;
      34157: inst = 32'hc404fc1;
      34158: inst = 32'h8220000;
      34159: inst = 32'h10408000;
      34160: inst = 32'hc404fcb;
      34161: inst = 32'h8220000;
      34162: inst = 32'h10408000;
      34163: inst = 32'hc404fdc;
      34164: inst = 32'h8220000;
      34165: inst = 32'h10408000;
      34166: inst = 32'hc404fdf;
      34167: inst = 32'h8220000;
      34168: inst = 32'h10408000;
      34169: inst = 32'hc404fe4;
      34170: inst = 32'h8220000;
      34171: inst = 32'h10408000;
      34172: inst = 32'hc404feb;
      34173: inst = 32'h8220000;
      34174: inst = 32'h10408000;
      34175: inst = 32'hc404ff1;
      34176: inst = 32'h8220000;
      34177: inst = 32'h10408000;
      34178: inst = 32'hc40500b;
      34179: inst = 32'h8220000;
      34180: inst = 32'h10408000;
      34181: inst = 32'hc405011;
      34182: inst = 32'h8220000;
      34183: inst = 32'h10408000;
      34184: inst = 32'hc405016;
      34185: inst = 32'h8220000;
      34186: inst = 32'h10408000;
      34187: inst = 32'hc405018;
      34188: inst = 32'h8220000;
      34189: inst = 32'h10408000;
      34190: inst = 32'hc40501c;
      34191: inst = 32'h8220000;
      34192: inst = 32'h10408000;
      34193: inst = 32'hc40501d;
      34194: inst = 32'h8220000;
      34195: inst = 32'h10408000;
      34196: inst = 32'hc405022;
      34197: inst = 32'h8220000;
      34198: inst = 32'h10408000;
      34199: inst = 32'hc40502c;
      34200: inst = 32'h8220000;
      34201: inst = 32'h10408000;
      34202: inst = 32'hc40502f;
      34203: inst = 32'h8220000;
      34204: inst = 32'h10408000;
      34205: inst = 32'hc405031;
      34206: inst = 32'h8220000;
      34207: inst = 32'h10408000;
      34208: inst = 32'hc405040;
      34209: inst = 32'h8220000;
      34210: inst = 32'h10408000;
      34211: inst = 32'hc405045;
      34212: inst = 32'h8220000;
      34213: inst = 32'h10408000;
      34214: inst = 32'hc405052;
      34215: inst = 32'h8220000;
      34216: inst = 32'hc20ffff;
      34217: inst = 32'h10408000;
      34218: inst = 32'hc404fec;
      34219: inst = 32'h8220000;
      34220: inst = 32'h58000000;
      34221: inst = 32'h13e0ffff;
      34222: inst = 32'h13e00000;
      34223: inst = 32'hfe085c4;
      34224: inst = 32'h5be00000;
      34225: inst = 32'h13e0ffff;
      34226: inst = 32'h13e00000;
      34227: inst = 32'hfe0882f;
      34228: inst = 32'h5be00000;
      34229: inst = 32'h13e0ffff;
      34230: inst = 32'h13e00000;
      34231: inst = 32'hfe0882f;
      34232: inst = 32'h5be00000;
      34233: inst = 32'h13e0ffff;
      34234: inst = 32'h13e00000;
      34235: inst = 32'hfe086ff;
      34236: inst = 32'h5be00000;
      34237: inst = 32'h13e0ffff;
      34238: inst = 32'h13e00000;
      34239: inst = 32'hfe086ff;
      34240: inst = 32'h5be00000;
      34241: inst = 32'h13e00000;
      34242: inst = 32'hfe085c4;
      34243: inst = 32'h5be00000;
      34244: inst = 32'hc6018c3;
      34245: inst = 32'h10408000;
      34246: inst = 32'hc40496b;
      34247: inst = 32'h8620000;
      34248: inst = 32'h10408000;
      34249: inst = 32'hc40496c;
      34250: inst = 32'h8620000;
      34251: inst = 32'h10408000;
      34252: inst = 32'hc40496d;
      34253: inst = 32'h8620000;
      34254: inst = 32'h10408000;
      34255: inst = 32'hc40496e;
      34256: inst = 32'h8620000;
      34257: inst = 32'h10408000;
      34258: inst = 32'hc40496f;
      34259: inst = 32'h8620000;
      34260: inst = 32'h10408000;
      34261: inst = 32'hc404970;
      34262: inst = 32'h8620000;
      34263: inst = 32'h10408000;
      34264: inst = 32'hc404971;
      34265: inst = 32'h8620000;
      34266: inst = 32'h10408000;
      34267: inst = 32'hc404972;
      34268: inst = 32'h8620000;
      34269: inst = 32'h10408000;
      34270: inst = 32'hc404973;
      34271: inst = 32'h8620000;
      34272: inst = 32'h10408000;
      34273: inst = 32'hc404974;
      34274: inst = 32'h8620000;
      34275: inst = 32'h10408000;
      34276: inst = 32'hc4049cb;
      34277: inst = 32'h8620000;
      34278: inst = 32'h10408000;
      34279: inst = 32'hc4049cc;
      34280: inst = 32'h8620000;
      34281: inst = 32'h10408000;
      34282: inst = 32'hc4049cd;
      34283: inst = 32'h8620000;
      34284: inst = 32'h10408000;
      34285: inst = 32'hc4049ce;
      34286: inst = 32'h8620000;
      34287: inst = 32'h10408000;
      34288: inst = 32'hc4049cf;
      34289: inst = 32'h8620000;
      34290: inst = 32'h10408000;
      34291: inst = 32'hc4049d0;
      34292: inst = 32'h8620000;
      34293: inst = 32'h10408000;
      34294: inst = 32'hc4049d1;
      34295: inst = 32'h8620000;
      34296: inst = 32'h10408000;
      34297: inst = 32'hc4049d2;
      34298: inst = 32'h8620000;
      34299: inst = 32'h10408000;
      34300: inst = 32'hc4049d3;
      34301: inst = 32'h8620000;
      34302: inst = 32'h10408000;
      34303: inst = 32'hc4049d4;
      34304: inst = 32'h8620000;
      34305: inst = 32'h10408000;
      34306: inst = 32'hc404a2b;
      34307: inst = 32'h8620000;
      34308: inst = 32'h10408000;
      34309: inst = 32'hc404a34;
      34310: inst = 32'h8620000;
      34311: inst = 32'h10408000;
      34312: inst = 32'hc404a8b;
      34313: inst = 32'h8620000;
      34314: inst = 32'h10408000;
      34315: inst = 32'hc404a8d;
      34316: inst = 32'h8620000;
      34317: inst = 32'h10408000;
      34318: inst = 32'hc404a92;
      34319: inst = 32'h8620000;
      34320: inst = 32'h10408000;
      34321: inst = 32'hc404a94;
      34322: inst = 32'h8620000;
      34323: inst = 32'h10408000;
      34324: inst = 32'hc404aeb;
      34325: inst = 32'h8620000;
      34326: inst = 32'h10408000;
      34327: inst = 32'hc404aed;
      34328: inst = 32'h8620000;
      34329: inst = 32'h10408000;
      34330: inst = 32'hc404af2;
      34331: inst = 32'h8620000;
      34332: inst = 32'h10408000;
      34333: inst = 32'hc404af4;
      34334: inst = 32'h8620000;
      34335: inst = 32'h10408000;
      34336: inst = 32'hc404b4b;
      34337: inst = 32'h8620000;
      34338: inst = 32'h10408000;
      34339: inst = 32'hc404b54;
      34340: inst = 32'h8620000;
      34341: inst = 32'h10408000;
      34342: inst = 32'hc404bab;
      34343: inst = 32'h8620000;
      34344: inst = 32'h10408000;
      34345: inst = 32'hc404bb4;
      34346: inst = 32'h8620000;
      34347: inst = 32'hc60f4ce;
      34348: inst = 32'h10408000;
      34349: inst = 32'hc404a2c;
      34350: inst = 32'h8620000;
      34351: inst = 32'h10408000;
      34352: inst = 32'hc404a2d;
      34353: inst = 32'h8620000;
      34354: inst = 32'h10408000;
      34355: inst = 32'hc404a2e;
      34356: inst = 32'h8620000;
      34357: inst = 32'h10408000;
      34358: inst = 32'hc404a2f;
      34359: inst = 32'h8620000;
      34360: inst = 32'h10408000;
      34361: inst = 32'hc404a30;
      34362: inst = 32'h8620000;
      34363: inst = 32'h10408000;
      34364: inst = 32'hc404a31;
      34365: inst = 32'h8620000;
      34366: inst = 32'h10408000;
      34367: inst = 32'hc404a32;
      34368: inst = 32'h8620000;
      34369: inst = 32'h10408000;
      34370: inst = 32'hc404a33;
      34371: inst = 32'h8620000;
      34372: inst = 32'h10408000;
      34373: inst = 32'hc404a8c;
      34374: inst = 32'h8620000;
      34375: inst = 32'h10408000;
      34376: inst = 32'hc404a8e;
      34377: inst = 32'h8620000;
      34378: inst = 32'h10408000;
      34379: inst = 32'hc404a8f;
      34380: inst = 32'h8620000;
      34381: inst = 32'h10408000;
      34382: inst = 32'hc404a90;
      34383: inst = 32'h8620000;
      34384: inst = 32'h10408000;
      34385: inst = 32'hc404a91;
      34386: inst = 32'h8620000;
      34387: inst = 32'h10408000;
      34388: inst = 32'hc404a93;
      34389: inst = 32'h8620000;
      34390: inst = 32'h10408000;
      34391: inst = 32'hc404aec;
      34392: inst = 32'h8620000;
      34393: inst = 32'h10408000;
      34394: inst = 32'hc404aee;
      34395: inst = 32'h8620000;
      34396: inst = 32'h10408000;
      34397: inst = 32'hc404aef;
      34398: inst = 32'h8620000;
      34399: inst = 32'h10408000;
      34400: inst = 32'hc404af0;
      34401: inst = 32'h8620000;
      34402: inst = 32'h10408000;
      34403: inst = 32'hc404af1;
      34404: inst = 32'h8620000;
      34405: inst = 32'h10408000;
      34406: inst = 32'hc404af3;
      34407: inst = 32'h8620000;
      34408: inst = 32'h10408000;
      34409: inst = 32'hc404b4c;
      34410: inst = 32'h8620000;
      34411: inst = 32'h10408000;
      34412: inst = 32'hc404b4d;
      34413: inst = 32'h8620000;
      34414: inst = 32'h10408000;
      34415: inst = 32'hc404b4e;
      34416: inst = 32'h8620000;
      34417: inst = 32'h10408000;
      34418: inst = 32'hc404b4f;
      34419: inst = 32'h8620000;
      34420: inst = 32'h10408000;
      34421: inst = 32'hc404b50;
      34422: inst = 32'h8620000;
      34423: inst = 32'h10408000;
      34424: inst = 32'hc404b51;
      34425: inst = 32'h8620000;
      34426: inst = 32'h10408000;
      34427: inst = 32'hc404b52;
      34428: inst = 32'h8620000;
      34429: inst = 32'h10408000;
      34430: inst = 32'hc404b53;
      34431: inst = 32'h8620000;
      34432: inst = 32'h10408000;
      34433: inst = 32'hc404bac;
      34434: inst = 32'h8620000;
      34435: inst = 32'h10408000;
      34436: inst = 32'hc404bad;
      34437: inst = 32'h8620000;
      34438: inst = 32'h10408000;
      34439: inst = 32'hc404bae;
      34440: inst = 32'h8620000;
      34441: inst = 32'h10408000;
      34442: inst = 32'hc404baf;
      34443: inst = 32'h8620000;
      34444: inst = 32'h10408000;
      34445: inst = 32'hc404bb0;
      34446: inst = 32'h8620000;
      34447: inst = 32'h10408000;
      34448: inst = 32'hc404bb1;
      34449: inst = 32'h8620000;
      34450: inst = 32'h10408000;
      34451: inst = 32'hc404bb2;
      34452: inst = 32'h8620000;
      34453: inst = 32'h10408000;
      34454: inst = 32'hc404bb3;
      34455: inst = 32'h8620000;
      34456: inst = 32'h10408000;
      34457: inst = 32'hc404c6b;
      34458: inst = 32'h8620000;
      34459: inst = 32'h10408000;
      34460: inst = 32'hc404c6c;
      34461: inst = 32'h8620000;
      34462: inst = 32'h10408000;
      34463: inst = 32'hc404c73;
      34464: inst = 32'h8620000;
      34465: inst = 32'h10408000;
      34466: inst = 32'hc404c74;
      34467: inst = 32'h8620000;
      34468: inst = 32'h10408000;
      34469: inst = 32'hc404dee;
      34470: inst = 32'h8620000;
      34471: inst = 32'h10408000;
      34472: inst = 32'hc404df1;
      34473: inst = 32'h8620000;
      34474: inst = 32'hc607800;
      34475: inst = 32'h10408000;
      34476: inst = 32'hc404c0d;
      34477: inst = 32'h8620000;
      34478: inst = 32'h10408000;
      34479: inst = 32'hc404c0e;
      34480: inst = 32'h8620000;
      34481: inst = 32'h10408000;
      34482: inst = 32'hc404c11;
      34483: inst = 32'h8620000;
      34484: inst = 32'h10408000;
      34485: inst = 32'hc404c12;
      34486: inst = 32'h8620000;
      34487: inst = 32'hc60a000;
      34488: inst = 32'h10408000;
      34489: inst = 32'hc404c0f;
      34490: inst = 32'h8620000;
      34491: inst = 32'h10408000;
      34492: inst = 32'hc404c10;
      34493: inst = 32'h8620000;
      34494: inst = 32'h10408000;
      34495: inst = 32'hc404c6d;
      34496: inst = 32'h8620000;
      34497: inst = 32'h10408000;
      34498: inst = 32'hc404c6e;
      34499: inst = 32'h8620000;
      34500: inst = 32'h10408000;
      34501: inst = 32'hc404c6f;
      34502: inst = 32'h8620000;
      34503: inst = 32'h10408000;
      34504: inst = 32'hc404c70;
      34505: inst = 32'h8620000;
      34506: inst = 32'h10408000;
      34507: inst = 32'hc404c71;
      34508: inst = 32'h8620000;
      34509: inst = 32'h10408000;
      34510: inst = 32'hc404c72;
      34511: inst = 32'h8620000;
      34512: inst = 32'h10408000;
      34513: inst = 32'hc404ccd;
      34514: inst = 32'h8620000;
      34515: inst = 32'h10408000;
      34516: inst = 32'hc404cce;
      34517: inst = 32'h8620000;
      34518: inst = 32'h10408000;
      34519: inst = 32'hc404ccf;
      34520: inst = 32'h8620000;
      34521: inst = 32'h10408000;
      34522: inst = 32'hc404cd0;
      34523: inst = 32'h8620000;
      34524: inst = 32'h10408000;
      34525: inst = 32'hc404cd1;
      34526: inst = 32'h8620000;
      34527: inst = 32'h10408000;
      34528: inst = 32'hc404cd2;
      34529: inst = 32'h8620000;
      34530: inst = 32'hc6010ac;
      34531: inst = 32'h10408000;
      34532: inst = 32'hc404d2d;
      34533: inst = 32'h8620000;
      34534: inst = 32'h10408000;
      34535: inst = 32'hc404d2e;
      34536: inst = 32'h8620000;
      34537: inst = 32'h10408000;
      34538: inst = 32'hc404d2f;
      34539: inst = 32'h8620000;
      34540: inst = 32'h10408000;
      34541: inst = 32'hc404d30;
      34542: inst = 32'h8620000;
      34543: inst = 32'h10408000;
      34544: inst = 32'hc404d31;
      34545: inst = 32'h8620000;
      34546: inst = 32'h10408000;
      34547: inst = 32'hc404d32;
      34548: inst = 32'h8620000;
      34549: inst = 32'hc60d42c;
      34550: inst = 32'h10408000;
      34551: inst = 32'hc404d8e;
      34552: inst = 32'h8620000;
      34553: inst = 32'h10408000;
      34554: inst = 32'hc404d91;
      34555: inst = 32'h8620000;
      34556: inst = 32'h13e00000;
      34557: inst = 32'hfe0895f;
      34558: inst = 32'h5be00000;
      34559: inst = 32'hc6018c3;
      34560: inst = 32'h10408000;
      34561: inst = 32'hc40496b;
      34562: inst = 32'h8620000;
      34563: inst = 32'h10408000;
      34564: inst = 32'hc40496c;
      34565: inst = 32'h8620000;
      34566: inst = 32'h10408000;
      34567: inst = 32'hc40496d;
      34568: inst = 32'h8620000;
      34569: inst = 32'h10408000;
      34570: inst = 32'hc40496e;
      34571: inst = 32'h8620000;
      34572: inst = 32'h10408000;
      34573: inst = 32'hc40496f;
      34574: inst = 32'h8620000;
      34575: inst = 32'h10408000;
      34576: inst = 32'hc404970;
      34577: inst = 32'h8620000;
      34578: inst = 32'h10408000;
      34579: inst = 32'hc404971;
      34580: inst = 32'h8620000;
      34581: inst = 32'h10408000;
      34582: inst = 32'hc404972;
      34583: inst = 32'h8620000;
      34584: inst = 32'h10408000;
      34585: inst = 32'hc404973;
      34586: inst = 32'h8620000;
      34587: inst = 32'h10408000;
      34588: inst = 32'hc404974;
      34589: inst = 32'h8620000;
      34590: inst = 32'h10408000;
      34591: inst = 32'hc4049cb;
      34592: inst = 32'h8620000;
      34593: inst = 32'h10408000;
      34594: inst = 32'hc4049cc;
      34595: inst = 32'h8620000;
      34596: inst = 32'h10408000;
      34597: inst = 32'hc4049cd;
      34598: inst = 32'h8620000;
      34599: inst = 32'h10408000;
      34600: inst = 32'hc4049ce;
      34601: inst = 32'h8620000;
      34602: inst = 32'h10408000;
      34603: inst = 32'hc4049cf;
      34604: inst = 32'h8620000;
      34605: inst = 32'h10408000;
      34606: inst = 32'hc4049d0;
      34607: inst = 32'h8620000;
      34608: inst = 32'h10408000;
      34609: inst = 32'hc4049d1;
      34610: inst = 32'h8620000;
      34611: inst = 32'h10408000;
      34612: inst = 32'hc4049d2;
      34613: inst = 32'h8620000;
      34614: inst = 32'h10408000;
      34615: inst = 32'hc4049d3;
      34616: inst = 32'h8620000;
      34617: inst = 32'h10408000;
      34618: inst = 32'hc4049d4;
      34619: inst = 32'h8620000;
      34620: inst = 32'h10408000;
      34621: inst = 32'hc404a2b;
      34622: inst = 32'h8620000;
      34623: inst = 32'h10408000;
      34624: inst = 32'hc404a2c;
      34625: inst = 32'h8620000;
      34626: inst = 32'h10408000;
      34627: inst = 32'hc404a8b;
      34628: inst = 32'h8620000;
      34629: inst = 32'h10408000;
      34630: inst = 32'hc404a93;
      34631: inst = 32'h8620000;
      34632: inst = 32'h10408000;
      34633: inst = 32'hc404aeb;
      34634: inst = 32'h8620000;
      34635: inst = 32'h10408000;
      34636: inst = 32'hc404af3;
      34637: inst = 32'h8620000;
      34638: inst = 32'h10408000;
      34639: inst = 32'hc404b4b;
      34640: inst = 32'h8620000;
      34641: inst = 32'h10408000;
      34642: inst = 32'hc404b4c;
      34643: inst = 32'h8620000;
      34644: inst = 32'h10408000;
      34645: inst = 32'hc404bab;
      34646: inst = 32'h8620000;
      34647: inst = 32'h10408000;
      34648: inst = 32'hc404bac;
      34649: inst = 32'h8620000;
      34650: inst = 32'hc60d42c;
      34651: inst = 32'h10408000;
      34652: inst = 32'hc404a2d;
      34653: inst = 32'h8620000;
      34654: inst = 32'h10408000;
      34655: inst = 32'hc404a2e;
      34656: inst = 32'h8620000;
      34657: inst = 32'h10408000;
      34658: inst = 32'hc404a2f;
      34659: inst = 32'h8620000;
      34660: inst = 32'h10408000;
      34661: inst = 32'hc404a30;
      34662: inst = 32'h8620000;
      34663: inst = 32'h10408000;
      34664: inst = 32'hc404a31;
      34665: inst = 32'h8620000;
      34666: inst = 32'h10408000;
      34667: inst = 32'hc404a32;
      34668: inst = 32'h8620000;
      34669: inst = 32'h10408000;
      34670: inst = 32'hc404a33;
      34671: inst = 32'h8620000;
      34672: inst = 32'h10408000;
      34673: inst = 32'hc404a34;
      34674: inst = 32'h8620000;
      34675: inst = 32'h10408000;
      34676: inst = 32'hc404b4d;
      34677: inst = 32'h8620000;
      34678: inst = 32'h10408000;
      34679: inst = 32'hc404bad;
      34680: inst = 32'h8620000;
      34681: inst = 32'h10408000;
      34682: inst = 32'hc404d8e;
      34683: inst = 32'h8620000;
      34684: inst = 32'h10408000;
      34685: inst = 32'hc404d91;
      34686: inst = 32'h8620000;
      34687: inst = 32'hc60f4ce;
      34688: inst = 32'h10408000;
      34689: inst = 32'hc404a8c;
      34690: inst = 32'h8620000;
      34691: inst = 32'h10408000;
      34692: inst = 32'hc404a8d;
      34693: inst = 32'h8620000;
      34694: inst = 32'h10408000;
      34695: inst = 32'hc404a8e;
      34696: inst = 32'h8620000;
      34697: inst = 32'h10408000;
      34698: inst = 32'hc404a8f;
      34699: inst = 32'h8620000;
      34700: inst = 32'h10408000;
      34701: inst = 32'hc404a90;
      34702: inst = 32'h8620000;
      34703: inst = 32'h10408000;
      34704: inst = 32'hc404a91;
      34705: inst = 32'h8620000;
      34706: inst = 32'h10408000;
      34707: inst = 32'hc404a92;
      34708: inst = 32'h8620000;
      34709: inst = 32'h10408000;
      34710: inst = 32'hc404a94;
      34711: inst = 32'h8620000;
      34712: inst = 32'h10408000;
      34713: inst = 32'hc404aec;
      34714: inst = 32'h8620000;
      34715: inst = 32'h10408000;
      34716: inst = 32'hc404aed;
      34717: inst = 32'h8620000;
      34718: inst = 32'h10408000;
      34719: inst = 32'hc404aee;
      34720: inst = 32'h8620000;
      34721: inst = 32'h10408000;
      34722: inst = 32'hc404aef;
      34723: inst = 32'h8620000;
      34724: inst = 32'h10408000;
      34725: inst = 32'hc404af0;
      34726: inst = 32'h8620000;
      34727: inst = 32'h10408000;
      34728: inst = 32'hc404af1;
      34729: inst = 32'h8620000;
      34730: inst = 32'h10408000;
      34731: inst = 32'hc404af2;
      34732: inst = 32'h8620000;
      34733: inst = 32'h10408000;
      34734: inst = 32'hc404af4;
      34735: inst = 32'h8620000;
      34736: inst = 32'h10408000;
      34737: inst = 32'hc404b4e;
      34738: inst = 32'h8620000;
      34739: inst = 32'h10408000;
      34740: inst = 32'hc404b4f;
      34741: inst = 32'h8620000;
      34742: inst = 32'h10408000;
      34743: inst = 32'hc404b50;
      34744: inst = 32'h8620000;
      34745: inst = 32'h10408000;
      34746: inst = 32'hc404b51;
      34747: inst = 32'h8620000;
      34748: inst = 32'h10408000;
      34749: inst = 32'hc404b52;
      34750: inst = 32'h8620000;
      34751: inst = 32'h10408000;
      34752: inst = 32'hc404b53;
      34753: inst = 32'h8620000;
      34754: inst = 32'h10408000;
      34755: inst = 32'hc404b54;
      34756: inst = 32'h8620000;
      34757: inst = 32'h10408000;
      34758: inst = 32'hc404bae;
      34759: inst = 32'h8620000;
      34760: inst = 32'h10408000;
      34761: inst = 32'hc404baf;
      34762: inst = 32'h8620000;
      34763: inst = 32'h10408000;
      34764: inst = 32'hc404bb0;
      34765: inst = 32'h8620000;
      34766: inst = 32'h10408000;
      34767: inst = 32'hc404bb1;
      34768: inst = 32'h8620000;
      34769: inst = 32'h10408000;
      34770: inst = 32'hc404bb2;
      34771: inst = 32'h8620000;
      34772: inst = 32'h10408000;
      34773: inst = 32'hc404bb3;
      34774: inst = 32'h8620000;
      34775: inst = 32'h10408000;
      34776: inst = 32'hc404bb4;
      34777: inst = 32'h8620000;
      34778: inst = 32'h10408000;
      34779: inst = 32'hc404c6f;
      34780: inst = 32'h8620000;
      34781: inst = 32'hc607841;
      34782: inst = 32'h10408000;
      34783: inst = 32'hc404c0d;
      34784: inst = 32'h8620000;
      34785: inst = 32'h10408000;
      34786: inst = 32'hc404c6d;
      34787: inst = 32'h8620000;
      34788: inst = 32'hc60a000;
      34789: inst = 32'h10408000;
      34790: inst = 32'hc404c0e;
      34791: inst = 32'h8620000;
      34792: inst = 32'h10408000;
      34793: inst = 32'hc404c0f;
      34794: inst = 32'h8620000;
      34795: inst = 32'h10408000;
      34796: inst = 32'hc404c10;
      34797: inst = 32'h8620000;
      34798: inst = 32'h10408000;
      34799: inst = 32'hc404c11;
      34800: inst = 32'h8620000;
      34801: inst = 32'h10408000;
      34802: inst = 32'hc404c12;
      34803: inst = 32'h8620000;
      34804: inst = 32'h10408000;
      34805: inst = 32'hc404c6e;
      34806: inst = 32'h8620000;
      34807: inst = 32'h10408000;
      34808: inst = 32'hc404c70;
      34809: inst = 32'h8620000;
      34810: inst = 32'h10408000;
      34811: inst = 32'hc404c71;
      34812: inst = 32'h8620000;
      34813: inst = 32'h10408000;
      34814: inst = 32'hc404c72;
      34815: inst = 32'h8620000;
      34816: inst = 32'h10408000;
      34817: inst = 32'hc404ccd;
      34818: inst = 32'h8620000;
      34819: inst = 32'h10408000;
      34820: inst = 32'hc404cce;
      34821: inst = 32'h8620000;
      34822: inst = 32'h10408000;
      34823: inst = 32'hc404ccf;
      34824: inst = 32'h8620000;
      34825: inst = 32'h10408000;
      34826: inst = 32'hc404cd0;
      34827: inst = 32'h8620000;
      34828: inst = 32'h10408000;
      34829: inst = 32'hc404cd1;
      34830: inst = 32'h8620000;
      34831: inst = 32'h10408000;
      34832: inst = 32'hc404cd2;
      34833: inst = 32'h8620000;
      34834: inst = 32'hc6010ac;
      34835: inst = 32'h10408000;
      34836: inst = 32'hc404d2d;
      34837: inst = 32'h8620000;
      34838: inst = 32'h10408000;
      34839: inst = 32'hc404d2e;
      34840: inst = 32'h8620000;
      34841: inst = 32'h10408000;
      34842: inst = 32'hc404d2f;
      34843: inst = 32'h8620000;
      34844: inst = 32'h10408000;
      34845: inst = 32'hc404d30;
      34846: inst = 32'h8620000;
      34847: inst = 32'h10408000;
      34848: inst = 32'hc404d31;
      34849: inst = 32'h8620000;
      34850: inst = 32'h10408000;
      34851: inst = 32'hc404d32;
      34852: inst = 32'h8620000;
      34853: inst = 32'h13e0ffff;
      34854: inst = 32'h13e00000;
      34855: inst = 32'hfe0882c;
      34856: inst = 32'h5be00000;
      34857: inst = 32'h13e00000;
      34858: inst = 32'hfe0895f;
      34859: inst = 32'h5be00000;
      34860: inst = 32'h13e00000;
      34861: inst = 32'hfe0895f;
      34862: inst = 32'h5be00000;
      34863: inst = 32'hc6018c3;
      34864: inst = 32'h10408000;
      34865: inst = 32'hc4049cb;
      34866: inst = 32'h8620000;
      34867: inst = 32'h10408000;
      34868: inst = 32'hc4049ca;
      34869: inst = 32'h8620000;
      34870: inst = 32'h10408000;
      34871: inst = 32'hc4049c9;
      34872: inst = 32'h8620000;
      34873: inst = 32'h10408000;
      34874: inst = 32'hc4049c8;
      34875: inst = 32'h8620000;
      34876: inst = 32'h10408000;
      34877: inst = 32'hc4049c7;
      34878: inst = 32'h8620000;
      34879: inst = 32'h10408000;
      34880: inst = 32'hc4049c6;
      34881: inst = 32'h8620000;
      34882: inst = 32'h10408000;
      34883: inst = 32'hc4049c5;
      34884: inst = 32'h8620000;
      34885: inst = 32'h10408000;
      34886: inst = 32'hc4049c4;
      34887: inst = 32'h8620000;
      34888: inst = 32'h10408000;
      34889: inst = 32'hc4049c3;
      34890: inst = 32'h8620000;
      34891: inst = 32'h10408000;
      34892: inst = 32'hc4049c2;
      34893: inst = 32'h8620000;
      34894: inst = 32'h10408000;
      34895: inst = 32'hc404a2b;
      34896: inst = 32'h8620000;
      34897: inst = 32'h10408000;
      34898: inst = 32'hc404a2a;
      34899: inst = 32'h8620000;
      34900: inst = 32'h10408000;
      34901: inst = 32'hc404a29;
      34902: inst = 32'h8620000;
      34903: inst = 32'h10408000;
      34904: inst = 32'hc404a28;
      34905: inst = 32'h8620000;
      34906: inst = 32'h10408000;
      34907: inst = 32'hc404a27;
      34908: inst = 32'h8620000;
      34909: inst = 32'h10408000;
      34910: inst = 32'hc404a26;
      34911: inst = 32'h8620000;
      34912: inst = 32'h10408000;
      34913: inst = 32'hc404a25;
      34914: inst = 32'h8620000;
      34915: inst = 32'h10408000;
      34916: inst = 32'hc404a24;
      34917: inst = 32'h8620000;
      34918: inst = 32'h10408000;
      34919: inst = 32'hc404a23;
      34920: inst = 32'h8620000;
      34921: inst = 32'h10408000;
      34922: inst = 32'hc404a22;
      34923: inst = 32'h8620000;
      34924: inst = 32'h10408000;
      34925: inst = 32'hc404a8b;
      34926: inst = 32'h8620000;
      34927: inst = 32'h10408000;
      34928: inst = 32'hc404a8a;
      34929: inst = 32'h8620000;
      34930: inst = 32'h10408000;
      34931: inst = 32'hc404aeb;
      34932: inst = 32'h8620000;
      34933: inst = 32'h10408000;
      34934: inst = 32'hc404ae3;
      34935: inst = 32'h8620000;
      34936: inst = 32'h10408000;
      34937: inst = 32'hc404b4b;
      34938: inst = 32'h8620000;
      34939: inst = 32'h10408000;
      34940: inst = 32'hc404b43;
      34941: inst = 32'h8620000;
      34942: inst = 32'h10408000;
      34943: inst = 32'hc404bab;
      34944: inst = 32'h8620000;
      34945: inst = 32'h10408000;
      34946: inst = 32'hc404baa;
      34947: inst = 32'h8620000;
      34948: inst = 32'h10408000;
      34949: inst = 32'hc404c0b;
      34950: inst = 32'h8620000;
      34951: inst = 32'h10408000;
      34952: inst = 32'hc404c0a;
      34953: inst = 32'h8620000;
      34954: inst = 32'hc60d42c;
      34955: inst = 32'h10408000;
      34956: inst = 32'hc404a89;
      34957: inst = 32'h8620000;
      34958: inst = 32'h10408000;
      34959: inst = 32'hc404a88;
      34960: inst = 32'h8620000;
      34961: inst = 32'h10408000;
      34962: inst = 32'hc404a87;
      34963: inst = 32'h8620000;
      34964: inst = 32'h10408000;
      34965: inst = 32'hc404a86;
      34966: inst = 32'h8620000;
      34967: inst = 32'h10408000;
      34968: inst = 32'hc404a85;
      34969: inst = 32'h8620000;
      34970: inst = 32'h10408000;
      34971: inst = 32'hc404a84;
      34972: inst = 32'h8620000;
      34973: inst = 32'h10408000;
      34974: inst = 32'hc404a83;
      34975: inst = 32'h8620000;
      34976: inst = 32'h10408000;
      34977: inst = 32'hc404a82;
      34978: inst = 32'h8620000;
      34979: inst = 32'h10408000;
      34980: inst = 32'hc404ba9;
      34981: inst = 32'h8620000;
      34982: inst = 32'h10408000;
      34983: inst = 32'hc404c09;
      34984: inst = 32'h8620000;
      34985: inst = 32'h10408000;
      34986: inst = 32'hc404de8;
      34987: inst = 32'h8620000;
      34988: inst = 32'h10408000;
      34989: inst = 32'hc404de5;
      34990: inst = 32'h8620000;
      34991: inst = 32'hc60f4ce;
      34992: inst = 32'h10408000;
      34993: inst = 32'hc404aea;
      34994: inst = 32'h8620000;
      34995: inst = 32'h10408000;
      34996: inst = 32'hc404ae9;
      34997: inst = 32'h8620000;
      34998: inst = 32'h10408000;
      34999: inst = 32'hc404ae8;
      35000: inst = 32'h8620000;
      35001: inst = 32'h10408000;
      35002: inst = 32'hc404ae7;
      35003: inst = 32'h8620000;
      35004: inst = 32'h10408000;
      35005: inst = 32'hc404ae6;
      35006: inst = 32'h8620000;
      35007: inst = 32'h10408000;
      35008: inst = 32'hc404ae5;
      35009: inst = 32'h8620000;
      35010: inst = 32'h10408000;
      35011: inst = 32'hc404ae4;
      35012: inst = 32'h8620000;
      35013: inst = 32'h10408000;
      35014: inst = 32'hc404ae2;
      35015: inst = 32'h8620000;
      35016: inst = 32'h10408000;
      35017: inst = 32'hc404b4a;
      35018: inst = 32'h8620000;
      35019: inst = 32'h10408000;
      35020: inst = 32'hc404b49;
      35021: inst = 32'h8620000;
      35022: inst = 32'h10408000;
      35023: inst = 32'hc404b48;
      35024: inst = 32'h8620000;
      35025: inst = 32'h10408000;
      35026: inst = 32'hc404b47;
      35027: inst = 32'h8620000;
      35028: inst = 32'h10408000;
      35029: inst = 32'hc404b46;
      35030: inst = 32'h8620000;
      35031: inst = 32'h10408000;
      35032: inst = 32'hc404b45;
      35033: inst = 32'h8620000;
      35034: inst = 32'h10408000;
      35035: inst = 32'hc404b44;
      35036: inst = 32'h8620000;
      35037: inst = 32'h10408000;
      35038: inst = 32'hc404b42;
      35039: inst = 32'h8620000;
      35040: inst = 32'h10408000;
      35041: inst = 32'hc404ba8;
      35042: inst = 32'h8620000;
      35043: inst = 32'h10408000;
      35044: inst = 32'hc404ba7;
      35045: inst = 32'h8620000;
      35046: inst = 32'h10408000;
      35047: inst = 32'hc404ba6;
      35048: inst = 32'h8620000;
      35049: inst = 32'h10408000;
      35050: inst = 32'hc404ba5;
      35051: inst = 32'h8620000;
      35052: inst = 32'h10408000;
      35053: inst = 32'hc404ba4;
      35054: inst = 32'h8620000;
      35055: inst = 32'h10408000;
      35056: inst = 32'hc404ba3;
      35057: inst = 32'h8620000;
      35058: inst = 32'h10408000;
      35059: inst = 32'hc404ba2;
      35060: inst = 32'h8620000;
      35061: inst = 32'h10408000;
      35062: inst = 32'hc404c08;
      35063: inst = 32'h8620000;
      35064: inst = 32'h10408000;
      35065: inst = 32'hc404c07;
      35066: inst = 32'h8620000;
      35067: inst = 32'h10408000;
      35068: inst = 32'hc404c06;
      35069: inst = 32'h8620000;
      35070: inst = 32'h10408000;
      35071: inst = 32'hc404c05;
      35072: inst = 32'h8620000;
      35073: inst = 32'h10408000;
      35074: inst = 32'hc404c04;
      35075: inst = 32'h8620000;
      35076: inst = 32'h10408000;
      35077: inst = 32'hc404c03;
      35078: inst = 32'h8620000;
      35079: inst = 32'h10408000;
      35080: inst = 32'hc404c02;
      35081: inst = 32'h8620000;
      35082: inst = 32'h10408000;
      35083: inst = 32'hc404cc7;
      35084: inst = 32'h8620000;
      35085: inst = 32'hc607841;
      35086: inst = 32'h10408000;
      35087: inst = 32'hc404c69;
      35088: inst = 32'h8620000;
      35089: inst = 32'h10408000;
      35090: inst = 32'hc404cc9;
      35091: inst = 32'h8620000;
      35092: inst = 32'hc60a000;
      35093: inst = 32'h10408000;
      35094: inst = 32'hc404c68;
      35095: inst = 32'h8620000;
      35096: inst = 32'h10408000;
      35097: inst = 32'hc404c67;
      35098: inst = 32'h8620000;
      35099: inst = 32'h10408000;
      35100: inst = 32'hc404c66;
      35101: inst = 32'h8620000;
      35102: inst = 32'h10408000;
      35103: inst = 32'hc404c65;
      35104: inst = 32'h8620000;
      35105: inst = 32'h10408000;
      35106: inst = 32'hc404c64;
      35107: inst = 32'h8620000;
      35108: inst = 32'h10408000;
      35109: inst = 32'hc404cc8;
      35110: inst = 32'h8620000;
      35111: inst = 32'h10408000;
      35112: inst = 32'hc404cc6;
      35113: inst = 32'h8620000;
      35114: inst = 32'h10408000;
      35115: inst = 32'hc404cc5;
      35116: inst = 32'h8620000;
      35117: inst = 32'h10408000;
      35118: inst = 32'hc404cc4;
      35119: inst = 32'h8620000;
      35120: inst = 32'h10408000;
      35121: inst = 32'hc404d29;
      35122: inst = 32'h8620000;
      35123: inst = 32'h10408000;
      35124: inst = 32'hc404d28;
      35125: inst = 32'h8620000;
      35126: inst = 32'h10408000;
      35127: inst = 32'hc404d27;
      35128: inst = 32'h8620000;
      35129: inst = 32'h10408000;
      35130: inst = 32'hc404d26;
      35131: inst = 32'h8620000;
      35132: inst = 32'h10408000;
      35133: inst = 32'hc404d25;
      35134: inst = 32'h8620000;
      35135: inst = 32'h10408000;
      35136: inst = 32'hc404d24;
      35137: inst = 32'h8620000;
      35138: inst = 32'hc6010ac;
      35139: inst = 32'h10408000;
      35140: inst = 32'hc404d89;
      35141: inst = 32'h8620000;
      35142: inst = 32'h10408000;
      35143: inst = 32'hc404d88;
      35144: inst = 32'h8620000;
      35145: inst = 32'h10408000;
      35146: inst = 32'hc404d87;
      35147: inst = 32'h8620000;
      35148: inst = 32'h10408000;
      35149: inst = 32'hc404d86;
      35150: inst = 32'h8620000;
      35151: inst = 32'h10408000;
      35152: inst = 32'hc404d85;
      35153: inst = 32'h8620000;
      35154: inst = 32'h10408000;
      35155: inst = 32'hc404d84;
      35156: inst = 32'h8620000;
      35157: inst = 32'h13e0ffff;
      35158: inst = 32'h13e00000;
      35159: inst = 32'hfe0895c;
      35160: inst = 32'h5be00000;
      35161: inst = 32'h13e00000;
      35162: inst = 32'hfe0895f;
      35163: inst = 32'h5be00000;
      35164: inst = 32'h13e00000;
      35165: inst = 32'hfe0895f;
      35166: inst = 32'h5be00000;
      35167: inst = 32'h58000000;
      35168: inst = 32'h10408000;
      35169: inst = 32'hc400002;
      35170: inst = 32'h4420000;
      35171: inst = 32'h10600000;
      35172: inst = 32'hc600010;
      35173: inst = 32'h38421800;
      35174: inst = 32'h4042000f;
      35175: inst = 32'h1c40000f;
      35176: inst = 32'h58000000;
      35177: inst = 32'h58200000;
      35178: inst = 32'h24612800;
      35179: inst = 32'h10a0ffff;
      35180: inst = 32'hca0ffe0;
      35181: inst = 32'h24822800;
      35182: inst = 32'h10a00000;
      35183: inst = 32'hca00004;
      35184: inst = 32'h38632800;
      35185: inst = 32'h38842800;
      35186: inst = 32'h10a00000;
      35187: inst = 32'hca08977;
      35188: inst = 32'h13e00001;
      35189: inst = 32'hfe0d96a;
      35190: inst = 32'h5be00000;
      35191: inst = 32'h8c50000;
      35192: inst = 32'h24612800;
      35193: inst = 32'h10a0ffff;
      35194: inst = 32'hca0ffe0;
      35195: inst = 32'h24822800;
      35196: inst = 32'h10a00000;
      35197: inst = 32'hca00004;
      35198: inst = 32'h38632800;
      35199: inst = 32'h38842800;
      35200: inst = 32'h10a00000;
      35201: inst = 32'hca08985;
      35202: inst = 32'h13e00001;
      35203: inst = 32'hfe0d96a;
      35204: inst = 32'h5be00000;
      35205: inst = 32'h8c50000;
      35206: inst = 32'h24612800;
      35207: inst = 32'h10a0ffff;
      35208: inst = 32'hca0ffe0;
      35209: inst = 32'h24822800;
      35210: inst = 32'h10a00000;
      35211: inst = 32'hca00004;
      35212: inst = 32'h38632800;
      35213: inst = 32'h38842800;
      35214: inst = 32'h10a00000;
      35215: inst = 32'hca08993;
      35216: inst = 32'h13e00001;
      35217: inst = 32'hfe0d96a;
      35218: inst = 32'h5be00000;
      35219: inst = 32'h8c50000;
      35220: inst = 32'h24612800;
      35221: inst = 32'h10a0ffff;
      35222: inst = 32'hca0ffe0;
      35223: inst = 32'h24822800;
      35224: inst = 32'h10a00000;
      35225: inst = 32'hca00004;
      35226: inst = 32'h38632800;
      35227: inst = 32'h38842800;
      35228: inst = 32'h10a00000;
      35229: inst = 32'hca089a1;
      35230: inst = 32'h13e00001;
      35231: inst = 32'hfe0d96a;
      35232: inst = 32'h5be00000;
      35233: inst = 32'h8c50000;
      35234: inst = 32'h24612800;
      35235: inst = 32'h10a0ffff;
      35236: inst = 32'hca0ffe0;
      35237: inst = 32'h24822800;
      35238: inst = 32'h10a00000;
      35239: inst = 32'hca00004;
      35240: inst = 32'h38632800;
      35241: inst = 32'h38842800;
      35242: inst = 32'h10a00000;
      35243: inst = 32'hca089af;
      35244: inst = 32'h13e00001;
      35245: inst = 32'hfe0d96a;
      35246: inst = 32'h5be00000;
      35247: inst = 32'h8c50000;
      35248: inst = 32'h24612800;
      35249: inst = 32'h10a0ffff;
      35250: inst = 32'hca0ffe0;
      35251: inst = 32'h24822800;
      35252: inst = 32'h10a00000;
      35253: inst = 32'hca00004;
      35254: inst = 32'h38632800;
      35255: inst = 32'h38842800;
      35256: inst = 32'h10a00000;
      35257: inst = 32'hca089bd;
      35258: inst = 32'h13e00001;
      35259: inst = 32'hfe0d96a;
      35260: inst = 32'h5be00000;
      35261: inst = 32'h8c50000;
      35262: inst = 32'h24612800;
      35263: inst = 32'h10a0ffff;
      35264: inst = 32'hca0ffe0;
      35265: inst = 32'h24822800;
      35266: inst = 32'h10a00000;
      35267: inst = 32'hca00004;
      35268: inst = 32'h38632800;
      35269: inst = 32'h38842800;
      35270: inst = 32'h10a00000;
      35271: inst = 32'hca089cb;
      35272: inst = 32'h13e00001;
      35273: inst = 32'hfe0d96a;
      35274: inst = 32'h5be00000;
      35275: inst = 32'h8c50000;
      35276: inst = 32'h24612800;
      35277: inst = 32'h10a0ffff;
      35278: inst = 32'hca0ffe0;
      35279: inst = 32'h24822800;
      35280: inst = 32'h10a00000;
      35281: inst = 32'hca00004;
      35282: inst = 32'h38632800;
      35283: inst = 32'h38842800;
      35284: inst = 32'h10a00000;
      35285: inst = 32'hca089d9;
      35286: inst = 32'h13e00001;
      35287: inst = 32'hfe0d96a;
      35288: inst = 32'h5be00000;
      35289: inst = 32'h8c50000;
      35290: inst = 32'h24612800;
      35291: inst = 32'h10a0ffff;
      35292: inst = 32'hca0ffe0;
      35293: inst = 32'h24822800;
      35294: inst = 32'h10a00000;
      35295: inst = 32'hca00004;
      35296: inst = 32'h38632800;
      35297: inst = 32'h38842800;
      35298: inst = 32'h10a00000;
      35299: inst = 32'hca089e7;
      35300: inst = 32'h13e00001;
      35301: inst = 32'hfe0d96a;
      35302: inst = 32'h5be00000;
      35303: inst = 32'h8c50000;
      35304: inst = 32'h24612800;
      35305: inst = 32'h10a0ffff;
      35306: inst = 32'hca0ffe0;
      35307: inst = 32'h24822800;
      35308: inst = 32'h10a00000;
      35309: inst = 32'hca00004;
      35310: inst = 32'h38632800;
      35311: inst = 32'h38842800;
      35312: inst = 32'h10a00000;
      35313: inst = 32'hca089f5;
      35314: inst = 32'h13e00001;
      35315: inst = 32'hfe0d96a;
      35316: inst = 32'h5be00000;
      35317: inst = 32'h8c50000;
      35318: inst = 32'h24612800;
      35319: inst = 32'h10a0ffff;
      35320: inst = 32'hca0ffe0;
      35321: inst = 32'h24822800;
      35322: inst = 32'h10a00000;
      35323: inst = 32'hca00004;
      35324: inst = 32'h38632800;
      35325: inst = 32'h38842800;
      35326: inst = 32'h10a00000;
      35327: inst = 32'hca08a03;
      35328: inst = 32'h13e00001;
      35329: inst = 32'hfe0d96a;
      35330: inst = 32'h5be00000;
      35331: inst = 32'h8c50000;
      35332: inst = 32'h24612800;
      35333: inst = 32'h10a0ffff;
      35334: inst = 32'hca0ffe0;
      35335: inst = 32'h24822800;
      35336: inst = 32'h10a00000;
      35337: inst = 32'hca00004;
      35338: inst = 32'h38632800;
      35339: inst = 32'h38842800;
      35340: inst = 32'h10a00000;
      35341: inst = 32'hca08a11;
      35342: inst = 32'h13e00001;
      35343: inst = 32'hfe0d96a;
      35344: inst = 32'h5be00000;
      35345: inst = 32'h8c50000;
      35346: inst = 32'h24612800;
      35347: inst = 32'h10a0ffff;
      35348: inst = 32'hca0ffe0;
      35349: inst = 32'h24822800;
      35350: inst = 32'h10a00000;
      35351: inst = 32'hca00004;
      35352: inst = 32'h38632800;
      35353: inst = 32'h38842800;
      35354: inst = 32'h10a00000;
      35355: inst = 32'hca08a1f;
      35356: inst = 32'h13e00001;
      35357: inst = 32'hfe0d96a;
      35358: inst = 32'h5be00000;
      35359: inst = 32'h8c50000;
      35360: inst = 32'h24612800;
      35361: inst = 32'h10a0ffff;
      35362: inst = 32'hca0ffe0;
      35363: inst = 32'h24822800;
      35364: inst = 32'h10a00000;
      35365: inst = 32'hca00004;
      35366: inst = 32'h38632800;
      35367: inst = 32'h38842800;
      35368: inst = 32'h10a00000;
      35369: inst = 32'hca08a2d;
      35370: inst = 32'h13e00001;
      35371: inst = 32'hfe0d96a;
      35372: inst = 32'h5be00000;
      35373: inst = 32'h8c50000;
      35374: inst = 32'h24612800;
      35375: inst = 32'h10a0ffff;
      35376: inst = 32'hca0ffe0;
      35377: inst = 32'h24822800;
      35378: inst = 32'h10a00000;
      35379: inst = 32'hca00004;
      35380: inst = 32'h38632800;
      35381: inst = 32'h38842800;
      35382: inst = 32'h10a00000;
      35383: inst = 32'hca08a3b;
      35384: inst = 32'h13e00001;
      35385: inst = 32'hfe0d96a;
      35386: inst = 32'h5be00000;
      35387: inst = 32'h8c50000;
      35388: inst = 32'h24612800;
      35389: inst = 32'h10a0ffff;
      35390: inst = 32'hca0ffe0;
      35391: inst = 32'h24822800;
      35392: inst = 32'h10a00000;
      35393: inst = 32'hca00004;
      35394: inst = 32'h38632800;
      35395: inst = 32'h38842800;
      35396: inst = 32'h10a00000;
      35397: inst = 32'hca08a49;
      35398: inst = 32'h13e00001;
      35399: inst = 32'hfe0d96a;
      35400: inst = 32'h5be00000;
      35401: inst = 32'h8c50000;
      35402: inst = 32'h24612800;
      35403: inst = 32'h10a0ffff;
      35404: inst = 32'hca0ffe0;
      35405: inst = 32'h24822800;
      35406: inst = 32'h10a00000;
      35407: inst = 32'hca00004;
      35408: inst = 32'h38632800;
      35409: inst = 32'h38842800;
      35410: inst = 32'h10a00000;
      35411: inst = 32'hca08a57;
      35412: inst = 32'h13e00001;
      35413: inst = 32'hfe0d96a;
      35414: inst = 32'h5be00000;
      35415: inst = 32'h8c50000;
      35416: inst = 32'h24612800;
      35417: inst = 32'h10a0ffff;
      35418: inst = 32'hca0ffe0;
      35419: inst = 32'h24822800;
      35420: inst = 32'h10a00000;
      35421: inst = 32'hca00004;
      35422: inst = 32'h38632800;
      35423: inst = 32'h38842800;
      35424: inst = 32'h10a00000;
      35425: inst = 32'hca08a65;
      35426: inst = 32'h13e00001;
      35427: inst = 32'hfe0d96a;
      35428: inst = 32'h5be00000;
      35429: inst = 32'h8c50000;
      35430: inst = 32'h24612800;
      35431: inst = 32'h10a0ffff;
      35432: inst = 32'hca0ffe0;
      35433: inst = 32'h24822800;
      35434: inst = 32'h10a00000;
      35435: inst = 32'hca00004;
      35436: inst = 32'h38632800;
      35437: inst = 32'h38842800;
      35438: inst = 32'h10a00000;
      35439: inst = 32'hca08a73;
      35440: inst = 32'h13e00001;
      35441: inst = 32'hfe0d96a;
      35442: inst = 32'h5be00000;
      35443: inst = 32'h8c50000;
      35444: inst = 32'h24612800;
      35445: inst = 32'h10a0ffff;
      35446: inst = 32'hca0ffe0;
      35447: inst = 32'h24822800;
      35448: inst = 32'h10a00000;
      35449: inst = 32'hca00004;
      35450: inst = 32'h38632800;
      35451: inst = 32'h38842800;
      35452: inst = 32'h10a00000;
      35453: inst = 32'hca08a81;
      35454: inst = 32'h13e00001;
      35455: inst = 32'hfe0d96a;
      35456: inst = 32'h5be00000;
      35457: inst = 32'h8c50000;
      35458: inst = 32'h24612800;
      35459: inst = 32'h10a0ffff;
      35460: inst = 32'hca0ffe0;
      35461: inst = 32'h24822800;
      35462: inst = 32'h10a00000;
      35463: inst = 32'hca00004;
      35464: inst = 32'h38632800;
      35465: inst = 32'h38842800;
      35466: inst = 32'h10a00000;
      35467: inst = 32'hca08a8f;
      35468: inst = 32'h13e00001;
      35469: inst = 32'hfe0d96a;
      35470: inst = 32'h5be00000;
      35471: inst = 32'h8c50000;
      35472: inst = 32'h24612800;
      35473: inst = 32'h10a0ffff;
      35474: inst = 32'hca0ffe0;
      35475: inst = 32'h24822800;
      35476: inst = 32'h10a00000;
      35477: inst = 32'hca00004;
      35478: inst = 32'h38632800;
      35479: inst = 32'h38842800;
      35480: inst = 32'h10a00000;
      35481: inst = 32'hca08a9d;
      35482: inst = 32'h13e00001;
      35483: inst = 32'hfe0d96a;
      35484: inst = 32'h5be00000;
      35485: inst = 32'h8c50000;
      35486: inst = 32'h24612800;
      35487: inst = 32'h10a0ffff;
      35488: inst = 32'hca0ffe0;
      35489: inst = 32'h24822800;
      35490: inst = 32'h10a00000;
      35491: inst = 32'hca00004;
      35492: inst = 32'h38632800;
      35493: inst = 32'h38842800;
      35494: inst = 32'h10a00000;
      35495: inst = 32'hca08aab;
      35496: inst = 32'h13e00001;
      35497: inst = 32'hfe0d96a;
      35498: inst = 32'h5be00000;
      35499: inst = 32'h8c50000;
      35500: inst = 32'h24612800;
      35501: inst = 32'h10a0ffff;
      35502: inst = 32'hca0ffe0;
      35503: inst = 32'h24822800;
      35504: inst = 32'h10a00000;
      35505: inst = 32'hca00004;
      35506: inst = 32'h38632800;
      35507: inst = 32'h38842800;
      35508: inst = 32'h10a00000;
      35509: inst = 32'hca08ab9;
      35510: inst = 32'h13e00001;
      35511: inst = 32'hfe0d96a;
      35512: inst = 32'h5be00000;
      35513: inst = 32'h8c50000;
      35514: inst = 32'h24612800;
      35515: inst = 32'h10a0ffff;
      35516: inst = 32'hca0ffe0;
      35517: inst = 32'h24822800;
      35518: inst = 32'h10a00000;
      35519: inst = 32'hca00004;
      35520: inst = 32'h38632800;
      35521: inst = 32'h38842800;
      35522: inst = 32'h10a00000;
      35523: inst = 32'hca08ac7;
      35524: inst = 32'h13e00001;
      35525: inst = 32'hfe0d96a;
      35526: inst = 32'h5be00000;
      35527: inst = 32'h8c50000;
      35528: inst = 32'h24612800;
      35529: inst = 32'h10a0ffff;
      35530: inst = 32'hca0ffe0;
      35531: inst = 32'h24822800;
      35532: inst = 32'h10a00000;
      35533: inst = 32'hca00004;
      35534: inst = 32'h38632800;
      35535: inst = 32'h38842800;
      35536: inst = 32'h10a00000;
      35537: inst = 32'hca08ad5;
      35538: inst = 32'h13e00001;
      35539: inst = 32'hfe0d96a;
      35540: inst = 32'h5be00000;
      35541: inst = 32'h8c50000;
      35542: inst = 32'h24612800;
      35543: inst = 32'h10a0ffff;
      35544: inst = 32'hca0ffe0;
      35545: inst = 32'h24822800;
      35546: inst = 32'h10a00000;
      35547: inst = 32'hca00004;
      35548: inst = 32'h38632800;
      35549: inst = 32'h38842800;
      35550: inst = 32'h10a00000;
      35551: inst = 32'hca08ae3;
      35552: inst = 32'h13e00001;
      35553: inst = 32'hfe0d96a;
      35554: inst = 32'h5be00000;
      35555: inst = 32'h8c50000;
      35556: inst = 32'h24612800;
      35557: inst = 32'h10a0ffff;
      35558: inst = 32'hca0ffe0;
      35559: inst = 32'h24822800;
      35560: inst = 32'h10a00000;
      35561: inst = 32'hca00004;
      35562: inst = 32'h38632800;
      35563: inst = 32'h38842800;
      35564: inst = 32'h10a00000;
      35565: inst = 32'hca08af1;
      35566: inst = 32'h13e00001;
      35567: inst = 32'hfe0d96a;
      35568: inst = 32'h5be00000;
      35569: inst = 32'h8c50000;
      35570: inst = 32'h24612800;
      35571: inst = 32'h10a0ffff;
      35572: inst = 32'hca0ffe0;
      35573: inst = 32'h24822800;
      35574: inst = 32'h10a00000;
      35575: inst = 32'hca00004;
      35576: inst = 32'h38632800;
      35577: inst = 32'h38842800;
      35578: inst = 32'h10a00000;
      35579: inst = 32'hca08aff;
      35580: inst = 32'h13e00001;
      35581: inst = 32'hfe0d96a;
      35582: inst = 32'h5be00000;
      35583: inst = 32'h8c50000;
      35584: inst = 32'h24612800;
      35585: inst = 32'h10a0ffff;
      35586: inst = 32'hca0ffe0;
      35587: inst = 32'h24822800;
      35588: inst = 32'h10a00000;
      35589: inst = 32'hca00004;
      35590: inst = 32'h38632800;
      35591: inst = 32'h38842800;
      35592: inst = 32'h10a00000;
      35593: inst = 32'hca08b0d;
      35594: inst = 32'h13e00001;
      35595: inst = 32'hfe0d96a;
      35596: inst = 32'h5be00000;
      35597: inst = 32'h8c50000;
      35598: inst = 32'h24612800;
      35599: inst = 32'h10a0ffff;
      35600: inst = 32'hca0ffe0;
      35601: inst = 32'h24822800;
      35602: inst = 32'h10a00000;
      35603: inst = 32'hca00004;
      35604: inst = 32'h38632800;
      35605: inst = 32'h38842800;
      35606: inst = 32'h10a00000;
      35607: inst = 32'hca08b1b;
      35608: inst = 32'h13e00001;
      35609: inst = 32'hfe0d96a;
      35610: inst = 32'h5be00000;
      35611: inst = 32'h8c50000;
      35612: inst = 32'h24612800;
      35613: inst = 32'h10a0ffff;
      35614: inst = 32'hca0ffe0;
      35615: inst = 32'h24822800;
      35616: inst = 32'h10a00000;
      35617: inst = 32'hca00004;
      35618: inst = 32'h38632800;
      35619: inst = 32'h38842800;
      35620: inst = 32'h10a00000;
      35621: inst = 32'hca08b29;
      35622: inst = 32'h13e00001;
      35623: inst = 32'hfe0d96a;
      35624: inst = 32'h5be00000;
      35625: inst = 32'h8c50000;
      35626: inst = 32'h24612800;
      35627: inst = 32'h10a0ffff;
      35628: inst = 32'hca0ffe0;
      35629: inst = 32'h24822800;
      35630: inst = 32'h10a00000;
      35631: inst = 32'hca00004;
      35632: inst = 32'h38632800;
      35633: inst = 32'h38842800;
      35634: inst = 32'h10a00000;
      35635: inst = 32'hca08b37;
      35636: inst = 32'h13e00001;
      35637: inst = 32'hfe0d96a;
      35638: inst = 32'h5be00000;
      35639: inst = 32'h8c50000;
      35640: inst = 32'h24612800;
      35641: inst = 32'h10a0ffff;
      35642: inst = 32'hca0ffe0;
      35643: inst = 32'h24822800;
      35644: inst = 32'h10a00000;
      35645: inst = 32'hca00004;
      35646: inst = 32'h38632800;
      35647: inst = 32'h38842800;
      35648: inst = 32'h10a00000;
      35649: inst = 32'hca08b45;
      35650: inst = 32'h13e00001;
      35651: inst = 32'hfe0d96a;
      35652: inst = 32'h5be00000;
      35653: inst = 32'h8c50000;
      35654: inst = 32'h24612800;
      35655: inst = 32'h10a0ffff;
      35656: inst = 32'hca0ffe0;
      35657: inst = 32'h24822800;
      35658: inst = 32'h10a00000;
      35659: inst = 32'hca00004;
      35660: inst = 32'h38632800;
      35661: inst = 32'h38842800;
      35662: inst = 32'h10a00000;
      35663: inst = 32'hca08b53;
      35664: inst = 32'h13e00001;
      35665: inst = 32'hfe0d96a;
      35666: inst = 32'h5be00000;
      35667: inst = 32'h8c50000;
      35668: inst = 32'h24612800;
      35669: inst = 32'h10a0ffff;
      35670: inst = 32'hca0ffe0;
      35671: inst = 32'h24822800;
      35672: inst = 32'h10a00000;
      35673: inst = 32'hca00004;
      35674: inst = 32'h38632800;
      35675: inst = 32'h38842800;
      35676: inst = 32'h10a00000;
      35677: inst = 32'hca08b61;
      35678: inst = 32'h13e00001;
      35679: inst = 32'hfe0d96a;
      35680: inst = 32'h5be00000;
      35681: inst = 32'h8c50000;
      35682: inst = 32'h24612800;
      35683: inst = 32'h10a0ffff;
      35684: inst = 32'hca0ffe0;
      35685: inst = 32'h24822800;
      35686: inst = 32'h10a00000;
      35687: inst = 32'hca00004;
      35688: inst = 32'h38632800;
      35689: inst = 32'h38842800;
      35690: inst = 32'h10a00000;
      35691: inst = 32'hca08b6f;
      35692: inst = 32'h13e00001;
      35693: inst = 32'hfe0d96a;
      35694: inst = 32'h5be00000;
      35695: inst = 32'h8c50000;
      35696: inst = 32'h24612800;
      35697: inst = 32'h10a0ffff;
      35698: inst = 32'hca0ffe0;
      35699: inst = 32'h24822800;
      35700: inst = 32'h10a00000;
      35701: inst = 32'hca00004;
      35702: inst = 32'h38632800;
      35703: inst = 32'h38842800;
      35704: inst = 32'h10a00000;
      35705: inst = 32'hca08b7d;
      35706: inst = 32'h13e00001;
      35707: inst = 32'hfe0d96a;
      35708: inst = 32'h5be00000;
      35709: inst = 32'h8c50000;
      35710: inst = 32'h24612800;
      35711: inst = 32'h10a0ffff;
      35712: inst = 32'hca0ffe0;
      35713: inst = 32'h24822800;
      35714: inst = 32'h10a00000;
      35715: inst = 32'hca00004;
      35716: inst = 32'h38632800;
      35717: inst = 32'h38842800;
      35718: inst = 32'h10a00000;
      35719: inst = 32'hca08b8b;
      35720: inst = 32'h13e00001;
      35721: inst = 32'hfe0d96a;
      35722: inst = 32'h5be00000;
      35723: inst = 32'h8c50000;
      35724: inst = 32'h24612800;
      35725: inst = 32'h10a0ffff;
      35726: inst = 32'hca0ffe0;
      35727: inst = 32'h24822800;
      35728: inst = 32'h10a00000;
      35729: inst = 32'hca00004;
      35730: inst = 32'h38632800;
      35731: inst = 32'h38842800;
      35732: inst = 32'h10a00000;
      35733: inst = 32'hca08b99;
      35734: inst = 32'h13e00001;
      35735: inst = 32'hfe0d96a;
      35736: inst = 32'h5be00000;
      35737: inst = 32'h8c50000;
      35738: inst = 32'h24612800;
      35739: inst = 32'h10a0ffff;
      35740: inst = 32'hca0ffe0;
      35741: inst = 32'h24822800;
      35742: inst = 32'h10a00000;
      35743: inst = 32'hca00004;
      35744: inst = 32'h38632800;
      35745: inst = 32'h38842800;
      35746: inst = 32'h10a00000;
      35747: inst = 32'hca08ba7;
      35748: inst = 32'h13e00001;
      35749: inst = 32'hfe0d96a;
      35750: inst = 32'h5be00000;
      35751: inst = 32'h8c50000;
      35752: inst = 32'h24612800;
      35753: inst = 32'h10a0ffff;
      35754: inst = 32'hca0ffe0;
      35755: inst = 32'h24822800;
      35756: inst = 32'h10a00000;
      35757: inst = 32'hca00004;
      35758: inst = 32'h38632800;
      35759: inst = 32'h38842800;
      35760: inst = 32'h10a00000;
      35761: inst = 32'hca08bb5;
      35762: inst = 32'h13e00001;
      35763: inst = 32'hfe0d96a;
      35764: inst = 32'h5be00000;
      35765: inst = 32'h8c50000;
      35766: inst = 32'h24612800;
      35767: inst = 32'h10a0ffff;
      35768: inst = 32'hca0ffe0;
      35769: inst = 32'h24822800;
      35770: inst = 32'h10a00000;
      35771: inst = 32'hca00004;
      35772: inst = 32'h38632800;
      35773: inst = 32'h38842800;
      35774: inst = 32'h10a00000;
      35775: inst = 32'hca08bc3;
      35776: inst = 32'h13e00001;
      35777: inst = 32'hfe0d96a;
      35778: inst = 32'h5be00000;
      35779: inst = 32'h8c50000;
      35780: inst = 32'h24612800;
      35781: inst = 32'h10a0ffff;
      35782: inst = 32'hca0ffe0;
      35783: inst = 32'h24822800;
      35784: inst = 32'h10a00000;
      35785: inst = 32'hca00004;
      35786: inst = 32'h38632800;
      35787: inst = 32'h38842800;
      35788: inst = 32'h10a00000;
      35789: inst = 32'hca08bd1;
      35790: inst = 32'h13e00001;
      35791: inst = 32'hfe0d96a;
      35792: inst = 32'h5be00000;
      35793: inst = 32'h8c50000;
      35794: inst = 32'h24612800;
      35795: inst = 32'h10a0ffff;
      35796: inst = 32'hca0ffe0;
      35797: inst = 32'h24822800;
      35798: inst = 32'h10a00000;
      35799: inst = 32'hca00004;
      35800: inst = 32'h38632800;
      35801: inst = 32'h38842800;
      35802: inst = 32'h10a00000;
      35803: inst = 32'hca08bdf;
      35804: inst = 32'h13e00001;
      35805: inst = 32'hfe0d96a;
      35806: inst = 32'h5be00000;
      35807: inst = 32'h8c50000;
      35808: inst = 32'h24612800;
      35809: inst = 32'h10a0ffff;
      35810: inst = 32'hca0ffe0;
      35811: inst = 32'h24822800;
      35812: inst = 32'h10a00000;
      35813: inst = 32'hca00004;
      35814: inst = 32'h38632800;
      35815: inst = 32'h38842800;
      35816: inst = 32'h10a00000;
      35817: inst = 32'hca08bed;
      35818: inst = 32'h13e00001;
      35819: inst = 32'hfe0d96a;
      35820: inst = 32'h5be00000;
      35821: inst = 32'h8c50000;
      35822: inst = 32'h24612800;
      35823: inst = 32'h10a0ffff;
      35824: inst = 32'hca0ffe0;
      35825: inst = 32'h24822800;
      35826: inst = 32'h10a00000;
      35827: inst = 32'hca00004;
      35828: inst = 32'h38632800;
      35829: inst = 32'h38842800;
      35830: inst = 32'h10a00000;
      35831: inst = 32'hca08bfb;
      35832: inst = 32'h13e00001;
      35833: inst = 32'hfe0d96a;
      35834: inst = 32'h5be00000;
      35835: inst = 32'h8c50000;
      35836: inst = 32'h24612800;
      35837: inst = 32'h10a0ffff;
      35838: inst = 32'hca0ffe0;
      35839: inst = 32'h24822800;
      35840: inst = 32'h10a00000;
      35841: inst = 32'hca00004;
      35842: inst = 32'h38632800;
      35843: inst = 32'h38842800;
      35844: inst = 32'h10a00000;
      35845: inst = 32'hca08c09;
      35846: inst = 32'h13e00001;
      35847: inst = 32'hfe0d96a;
      35848: inst = 32'h5be00000;
      35849: inst = 32'h8c50000;
      35850: inst = 32'h24612800;
      35851: inst = 32'h10a0ffff;
      35852: inst = 32'hca0ffe0;
      35853: inst = 32'h24822800;
      35854: inst = 32'h10a00000;
      35855: inst = 32'hca00004;
      35856: inst = 32'h38632800;
      35857: inst = 32'h38842800;
      35858: inst = 32'h10a00000;
      35859: inst = 32'hca08c17;
      35860: inst = 32'h13e00001;
      35861: inst = 32'hfe0d96a;
      35862: inst = 32'h5be00000;
      35863: inst = 32'h8c50000;
      35864: inst = 32'h24612800;
      35865: inst = 32'h10a0ffff;
      35866: inst = 32'hca0ffe0;
      35867: inst = 32'h24822800;
      35868: inst = 32'h10a00000;
      35869: inst = 32'hca00004;
      35870: inst = 32'h38632800;
      35871: inst = 32'h38842800;
      35872: inst = 32'h10a00000;
      35873: inst = 32'hca08c25;
      35874: inst = 32'h13e00001;
      35875: inst = 32'hfe0d96a;
      35876: inst = 32'h5be00000;
      35877: inst = 32'h8c50000;
      35878: inst = 32'h24612800;
      35879: inst = 32'h10a0ffff;
      35880: inst = 32'hca0ffe0;
      35881: inst = 32'h24822800;
      35882: inst = 32'h10a00000;
      35883: inst = 32'hca00004;
      35884: inst = 32'h38632800;
      35885: inst = 32'h38842800;
      35886: inst = 32'h10a00000;
      35887: inst = 32'hca08c33;
      35888: inst = 32'h13e00001;
      35889: inst = 32'hfe0d96a;
      35890: inst = 32'h5be00000;
      35891: inst = 32'h8c50000;
      35892: inst = 32'h24612800;
      35893: inst = 32'h10a0ffff;
      35894: inst = 32'hca0ffe0;
      35895: inst = 32'h24822800;
      35896: inst = 32'h10a00000;
      35897: inst = 32'hca00004;
      35898: inst = 32'h38632800;
      35899: inst = 32'h38842800;
      35900: inst = 32'h10a00000;
      35901: inst = 32'hca08c41;
      35902: inst = 32'h13e00001;
      35903: inst = 32'hfe0d96a;
      35904: inst = 32'h5be00000;
      35905: inst = 32'h8c50000;
      35906: inst = 32'h24612800;
      35907: inst = 32'h10a0ffff;
      35908: inst = 32'hca0ffe0;
      35909: inst = 32'h24822800;
      35910: inst = 32'h10a00000;
      35911: inst = 32'hca00004;
      35912: inst = 32'h38632800;
      35913: inst = 32'h38842800;
      35914: inst = 32'h10a00000;
      35915: inst = 32'hca08c4f;
      35916: inst = 32'h13e00001;
      35917: inst = 32'hfe0d96a;
      35918: inst = 32'h5be00000;
      35919: inst = 32'h8c50000;
      35920: inst = 32'h24612800;
      35921: inst = 32'h10a0ffff;
      35922: inst = 32'hca0ffe0;
      35923: inst = 32'h24822800;
      35924: inst = 32'h10a00000;
      35925: inst = 32'hca00004;
      35926: inst = 32'h38632800;
      35927: inst = 32'h38842800;
      35928: inst = 32'h10a00000;
      35929: inst = 32'hca08c5d;
      35930: inst = 32'h13e00001;
      35931: inst = 32'hfe0d96a;
      35932: inst = 32'h5be00000;
      35933: inst = 32'h8c50000;
      35934: inst = 32'h24612800;
      35935: inst = 32'h10a0ffff;
      35936: inst = 32'hca0ffe0;
      35937: inst = 32'h24822800;
      35938: inst = 32'h10a00000;
      35939: inst = 32'hca00004;
      35940: inst = 32'h38632800;
      35941: inst = 32'h38842800;
      35942: inst = 32'h10a00000;
      35943: inst = 32'hca08c6b;
      35944: inst = 32'h13e00001;
      35945: inst = 32'hfe0d96a;
      35946: inst = 32'h5be00000;
      35947: inst = 32'h8c50000;
      35948: inst = 32'h24612800;
      35949: inst = 32'h10a0ffff;
      35950: inst = 32'hca0ffe0;
      35951: inst = 32'h24822800;
      35952: inst = 32'h10a00000;
      35953: inst = 32'hca00004;
      35954: inst = 32'h38632800;
      35955: inst = 32'h38842800;
      35956: inst = 32'h10a00000;
      35957: inst = 32'hca08c79;
      35958: inst = 32'h13e00001;
      35959: inst = 32'hfe0d96a;
      35960: inst = 32'h5be00000;
      35961: inst = 32'h8c50000;
      35962: inst = 32'h24612800;
      35963: inst = 32'h10a0ffff;
      35964: inst = 32'hca0ffe0;
      35965: inst = 32'h24822800;
      35966: inst = 32'h10a00000;
      35967: inst = 32'hca00004;
      35968: inst = 32'h38632800;
      35969: inst = 32'h38842800;
      35970: inst = 32'h10a00000;
      35971: inst = 32'hca08c87;
      35972: inst = 32'h13e00001;
      35973: inst = 32'hfe0d96a;
      35974: inst = 32'h5be00000;
      35975: inst = 32'h8c50000;
      35976: inst = 32'h24612800;
      35977: inst = 32'h10a0ffff;
      35978: inst = 32'hca0ffe0;
      35979: inst = 32'h24822800;
      35980: inst = 32'h10a00000;
      35981: inst = 32'hca00004;
      35982: inst = 32'h38632800;
      35983: inst = 32'h38842800;
      35984: inst = 32'h10a00000;
      35985: inst = 32'hca08c95;
      35986: inst = 32'h13e00001;
      35987: inst = 32'hfe0d96a;
      35988: inst = 32'h5be00000;
      35989: inst = 32'h8c50000;
      35990: inst = 32'h24612800;
      35991: inst = 32'h10a0ffff;
      35992: inst = 32'hca0ffe0;
      35993: inst = 32'h24822800;
      35994: inst = 32'h10a00000;
      35995: inst = 32'hca00004;
      35996: inst = 32'h38632800;
      35997: inst = 32'h38842800;
      35998: inst = 32'h10a00000;
      35999: inst = 32'hca08ca3;
      36000: inst = 32'h13e00001;
      36001: inst = 32'hfe0d96a;
      36002: inst = 32'h5be00000;
      36003: inst = 32'h8c50000;
      36004: inst = 32'h24612800;
      36005: inst = 32'h10a0ffff;
      36006: inst = 32'hca0ffe0;
      36007: inst = 32'h24822800;
      36008: inst = 32'h10a00000;
      36009: inst = 32'hca00004;
      36010: inst = 32'h38632800;
      36011: inst = 32'h38842800;
      36012: inst = 32'h10a00000;
      36013: inst = 32'hca08cb1;
      36014: inst = 32'h13e00001;
      36015: inst = 32'hfe0d96a;
      36016: inst = 32'h5be00000;
      36017: inst = 32'h8c50000;
      36018: inst = 32'h24612800;
      36019: inst = 32'h10a0ffff;
      36020: inst = 32'hca0ffe0;
      36021: inst = 32'h24822800;
      36022: inst = 32'h10a00000;
      36023: inst = 32'hca00004;
      36024: inst = 32'h38632800;
      36025: inst = 32'h38842800;
      36026: inst = 32'h10a00000;
      36027: inst = 32'hca08cbf;
      36028: inst = 32'h13e00001;
      36029: inst = 32'hfe0d96a;
      36030: inst = 32'h5be00000;
      36031: inst = 32'h8c50000;
      36032: inst = 32'h24612800;
      36033: inst = 32'h10a0ffff;
      36034: inst = 32'hca0ffe0;
      36035: inst = 32'h24822800;
      36036: inst = 32'h10a00000;
      36037: inst = 32'hca00004;
      36038: inst = 32'h38632800;
      36039: inst = 32'h38842800;
      36040: inst = 32'h10a00000;
      36041: inst = 32'hca08ccd;
      36042: inst = 32'h13e00001;
      36043: inst = 32'hfe0d96a;
      36044: inst = 32'h5be00000;
      36045: inst = 32'h8c50000;
      36046: inst = 32'h24612800;
      36047: inst = 32'h10a0ffff;
      36048: inst = 32'hca0ffe0;
      36049: inst = 32'h24822800;
      36050: inst = 32'h10a00000;
      36051: inst = 32'hca00004;
      36052: inst = 32'h38632800;
      36053: inst = 32'h38842800;
      36054: inst = 32'h10a00000;
      36055: inst = 32'hca08cdb;
      36056: inst = 32'h13e00001;
      36057: inst = 32'hfe0d96a;
      36058: inst = 32'h5be00000;
      36059: inst = 32'h8c50000;
      36060: inst = 32'h24612800;
      36061: inst = 32'h10a0ffff;
      36062: inst = 32'hca0ffe0;
      36063: inst = 32'h24822800;
      36064: inst = 32'h10a00000;
      36065: inst = 32'hca00004;
      36066: inst = 32'h38632800;
      36067: inst = 32'h38842800;
      36068: inst = 32'h10a00000;
      36069: inst = 32'hca08ce9;
      36070: inst = 32'h13e00001;
      36071: inst = 32'hfe0d96a;
      36072: inst = 32'h5be00000;
      36073: inst = 32'h8c50000;
      36074: inst = 32'h24612800;
      36075: inst = 32'h10a0ffff;
      36076: inst = 32'hca0ffe0;
      36077: inst = 32'h24822800;
      36078: inst = 32'h10a00000;
      36079: inst = 32'hca00004;
      36080: inst = 32'h38632800;
      36081: inst = 32'h38842800;
      36082: inst = 32'h10a00000;
      36083: inst = 32'hca08cf7;
      36084: inst = 32'h13e00001;
      36085: inst = 32'hfe0d96a;
      36086: inst = 32'h5be00000;
      36087: inst = 32'h8c50000;
      36088: inst = 32'h24612800;
      36089: inst = 32'h10a0ffff;
      36090: inst = 32'hca0ffe0;
      36091: inst = 32'h24822800;
      36092: inst = 32'h10a00000;
      36093: inst = 32'hca00004;
      36094: inst = 32'h38632800;
      36095: inst = 32'h38842800;
      36096: inst = 32'h10a00000;
      36097: inst = 32'hca08d05;
      36098: inst = 32'h13e00001;
      36099: inst = 32'hfe0d96a;
      36100: inst = 32'h5be00000;
      36101: inst = 32'h8c50000;
      36102: inst = 32'h24612800;
      36103: inst = 32'h10a0ffff;
      36104: inst = 32'hca0ffe0;
      36105: inst = 32'h24822800;
      36106: inst = 32'h10a00000;
      36107: inst = 32'hca00004;
      36108: inst = 32'h38632800;
      36109: inst = 32'h38842800;
      36110: inst = 32'h10a00000;
      36111: inst = 32'hca08d13;
      36112: inst = 32'h13e00001;
      36113: inst = 32'hfe0d96a;
      36114: inst = 32'h5be00000;
      36115: inst = 32'h8c50000;
      36116: inst = 32'h24612800;
      36117: inst = 32'h10a0ffff;
      36118: inst = 32'hca0ffe0;
      36119: inst = 32'h24822800;
      36120: inst = 32'h10a00000;
      36121: inst = 32'hca00004;
      36122: inst = 32'h38632800;
      36123: inst = 32'h38842800;
      36124: inst = 32'h10a00000;
      36125: inst = 32'hca08d21;
      36126: inst = 32'h13e00001;
      36127: inst = 32'hfe0d96a;
      36128: inst = 32'h5be00000;
      36129: inst = 32'h8c50000;
      36130: inst = 32'h24612800;
      36131: inst = 32'h10a0ffff;
      36132: inst = 32'hca0ffe0;
      36133: inst = 32'h24822800;
      36134: inst = 32'h10a00000;
      36135: inst = 32'hca00004;
      36136: inst = 32'h38632800;
      36137: inst = 32'h38842800;
      36138: inst = 32'h10a00000;
      36139: inst = 32'hca08d2f;
      36140: inst = 32'h13e00001;
      36141: inst = 32'hfe0d96a;
      36142: inst = 32'h5be00000;
      36143: inst = 32'h8c50000;
      36144: inst = 32'h24612800;
      36145: inst = 32'h10a0ffff;
      36146: inst = 32'hca0ffe0;
      36147: inst = 32'h24822800;
      36148: inst = 32'h10a00000;
      36149: inst = 32'hca00004;
      36150: inst = 32'h38632800;
      36151: inst = 32'h38842800;
      36152: inst = 32'h10a00000;
      36153: inst = 32'hca08d3d;
      36154: inst = 32'h13e00001;
      36155: inst = 32'hfe0d96a;
      36156: inst = 32'h5be00000;
      36157: inst = 32'h8c50000;
      36158: inst = 32'h24612800;
      36159: inst = 32'h10a0ffff;
      36160: inst = 32'hca0ffe0;
      36161: inst = 32'h24822800;
      36162: inst = 32'h10a00000;
      36163: inst = 32'hca00004;
      36164: inst = 32'h38632800;
      36165: inst = 32'h38842800;
      36166: inst = 32'h10a00000;
      36167: inst = 32'hca08d4b;
      36168: inst = 32'h13e00001;
      36169: inst = 32'hfe0d96a;
      36170: inst = 32'h5be00000;
      36171: inst = 32'h8c50000;
      36172: inst = 32'h24612800;
      36173: inst = 32'h10a0ffff;
      36174: inst = 32'hca0ffe0;
      36175: inst = 32'h24822800;
      36176: inst = 32'h10a00000;
      36177: inst = 32'hca00004;
      36178: inst = 32'h38632800;
      36179: inst = 32'h38842800;
      36180: inst = 32'h10a00000;
      36181: inst = 32'hca08d59;
      36182: inst = 32'h13e00001;
      36183: inst = 32'hfe0d96a;
      36184: inst = 32'h5be00000;
      36185: inst = 32'h8c50000;
      36186: inst = 32'h24612800;
      36187: inst = 32'h10a0ffff;
      36188: inst = 32'hca0ffe0;
      36189: inst = 32'h24822800;
      36190: inst = 32'h10a00000;
      36191: inst = 32'hca00004;
      36192: inst = 32'h38632800;
      36193: inst = 32'h38842800;
      36194: inst = 32'h10a00000;
      36195: inst = 32'hca08d67;
      36196: inst = 32'h13e00001;
      36197: inst = 32'hfe0d96a;
      36198: inst = 32'h5be00000;
      36199: inst = 32'h8c50000;
      36200: inst = 32'h24612800;
      36201: inst = 32'h10a0ffff;
      36202: inst = 32'hca0ffe0;
      36203: inst = 32'h24822800;
      36204: inst = 32'h10a00000;
      36205: inst = 32'hca00004;
      36206: inst = 32'h38632800;
      36207: inst = 32'h38842800;
      36208: inst = 32'h10a00000;
      36209: inst = 32'hca08d75;
      36210: inst = 32'h13e00001;
      36211: inst = 32'hfe0d96a;
      36212: inst = 32'h5be00000;
      36213: inst = 32'h8c50000;
      36214: inst = 32'h24612800;
      36215: inst = 32'h10a0ffff;
      36216: inst = 32'hca0ffe0;
      36217: inst = 32'h24822800;
      36218: inst = 32'h10a00000;
      36219: inst = 32'hca00004;
      36220: inst = 32'h38632800;
      36221: inst = 32'h38842800;
      36222: inst = 32'h10a00000;
      36223: inst = 32'hca08d83;
      36224: inst = 32'h13e00001;
      36225: inst = 32'hfe0d96a;
      36226: inst = 32'h5be00000;
      36227: inst = 32'h8c50000;
      36228: inst = 32'h24612800;
      36229: inst = 32'h10a0ffff;
      36230: inst = 32'hca0ffe0;
      36231: inst = 32'h24822800;
      36232: inst = 32'h10a00000;
      36233: inst = 32'hca00004;
      36234: inst = 32'h38632800;
      36235: inst = 32'h38842800;
      36236: inst = 32'h10a00000;
      36237: inst = 32'hca08d91;
      36238: inst = 32'h13e00001;
      36239: inst = 32'hfe0d96a;
      36240: inst = 32'h5be00000;
      36241: inst = 32'h8c50000;
      36242: inst = 32'h24612800;
      36243: inst = 32'h10a0ffff;
      36244: inst = 32'hca0ffe0;
      36245: inst = 32'h24822800;
      36246: inst = 32'h10a00000;
      36247: inst = 32'hca00004;
      36248: inst = 32'h38632800;
      36249: inst = 32'h38842800;
      36250: inst = 32'h10a00000;
      36251: inst = 32'hca08d9f;
      36252: inst = 32'h13e00001;
      36253: inst = 32'hfe0d96a;
      36254: inst = 32'h5be00000;
      36255: inst = 32'h8c50000;
      36256: inst = 32'h24612800;
      36257: inst = 32'h10a0ffff;
      36258: inst = 32'hca0ffe0;
      36259: inst = 32'h24822800;
      36260: inst = 32'h10a00000;
      36261: inst = 32'hca00004;
      36262: inst = 32'h38632800;
      36263: inst = 32'h38842800;
      36264: inst = 32'h10a00000;
      36265: inst = 32'hca08dad;
      36266: inst = 32'h13e00001;
      36267: inst = 32'hfe0d96a;
      36268: inst = 32'h5be00000;
      36269: inst = 32'h8c50000;
      36270: inst = 32'h24612800;
      36271: inst = 32'h10a0ffff;
      36272: inst = 32'hca0ffe0;
      36273: inst = 32'h24822800;
      36274: inst = 32'h10a00000;
      36275: inst = 32'hca00004;
      36276: inst = 32'h38632800;
      36277: inst = 32'h38842800;
      36278: inst = 32'h10a00000;
      36279: inst = 32'hca08dbb;
      36280: inst = 32'h13e00001;
      36281: inst = 32'hfe0d96a;
      36282: inst = 32'h5be00000;
      36283: inst = 32'h8c50000;
      36284: inst = 32'h24612800;
      36285: inst = 32'h10a0ffff;
      36286: inst = 32'hca0ffe0;
      36287: inst = 32'h24822800;
      36288: inst = 32'h10a00000;
      36289: inst = 32'hca00004;
      36290: inst = 32'h38632800;
      36291: inst = 32'h38842800;
      36292: inst = 32'h10a00000;
      36293: inst = 32'hca08dc9;
      36294: inst = 32'h13e00001;
      36295: inst = 32'hfe0d96a;
      36296: inst = 32'h5be00000;
      36297: inst = 32'h8c50000;
      36298: inst = 32'h24612800;
      36299: inst = 32'h10a0ffff;
      36300: inst = 32'hca0ffe0;
      36301: inst = 32'h24822800;
      36302: inst = 32'h10a00000;
      36303: inst = 32'hca00004;
      36304: inst = 32'h38632800;
      36305: inst = 32'h38842800;
      36306: inst = 32'h10a00000;
      36307: inst = 32'hca08dd7;
      36308: inst = 32'h13e00001;
      36309: inst = 32'hfe0d96a;
      36310: inst = 32'h5be00000;
      36311: inst = 32'h8c50000;
      36312: inst = 32'h24612800;
      36313: inst = 32'h10a0ffff;
      36314: inst = 32'hca0ffe0;
      36315: inst = 32'h24822800;
      36316: inst = 32'h10a00000;
      36317: inst = 32'hca00004;
      36318: inst = 32'h38632800;
      36319: inst = 32'h38842800;
      36320: inst = 32'h10a00000;
      36321: inst = 32'hca08de5;
      36322: inst = 32'h13e00001;
      36323: inst = 32'hfe0d96a;
      36324: inst = 32'h5be00000;
      36325: inst = 32'h8c50000;
      36326: inst = 32'h24612800;
      36327: inst = 32'h10a0ffff;
      36328: inst = 32'hca0ffe0;
      36329: inst = 32'h24822800;
      36330: inst = 32'h10a00000;
      36331: inst = 32'hca00004;
      36332: inst = 32'h38632800;
      36333: inst = 32'h38842800;
      36334: inst = 32'h10a00000;
      36335: inst = 32'hca08df3;
      36336: inst = 32'h13e00001;
      36337: inst = 32'hfe0d96a;
      36338: inst = 32'h5be00000;
      36339: inst = 32'h8c50000;
      36340: inst = 32'h24612800;
      36341: inst = 32'h10a0ffff;
      36342: inst = 32'hca0ffe0;
      36343: inst = 32'h24822800;
      36344: inst = 32'h10a00000;
      36345: inst = 32'hca00004;
      36346: inst = 32'h38632800;
      36347: inst = 32'h38842800;
      36348: inst = 32'h10a00000;
      36349: inst = 32'hca08e01;
      36350: inst = 32'h13e00001;
      36351: inst = 32'hfe0d96a;
      36352: inst = 32'h5be00000;
      36353: inst = 32'h8c50000;
      36354: inst = 32'h24612800;
      36355: inst = 32'h10a0ffff;
      36356: inst = 32'hca0ffe0;
      36357: inst = 32'h24822800;
      36358: inst = 32'h10a00000;
      36359: inst = 32'hca00004;
      36360: inst = 32'h38632800;
      36361: inst = 32'h38842800;
      36362: inst = 32'h10a00000;
      36363: inst = 32'hca08e0f;
      36364: inst = 32'h13e00001;
      36365: inst = 32'hfe0d96a;
      36366: inst = 32'h5be00000;
      36367: inst = 32'h8c50000;
      36368: inst = 32'h24612800;
      36369: inst = 32'h10a0ffff;
      36370: inst = 32'hca0ffe0;
      36371: inst = 32'h24822800;
      36372: inst = 32'h10a00000;
      36373: inst = 32'hca00004;
      36374: inst = 32'h38632800;
      36375: inst = 32'h38842800;
      36376: inst = 32'h10a00000;
      36377: inst = 32'hca08e1d;
      36378: inst = 32'h13e00001;
      36379: inst = 32'hfe0d96a;
      36380: inst = 32'h5be00000;
      36381: inst = 32'h8c50000;
      36382: inst = 32'h24612800;
      36383: inst = 32'h10a0ffff;
      36384: inst = 32'hca0ffe0;
      36385: inst = 32'h24822800;
      36386: inst = 32'h10a00000;
      36387: inst = 32'hca00004;
      36388: inst = 32'h38632800;
      36389: inst = 32'h38842800;
      36390: inst = 32'h10a00000;
      36391: inst = 32'hca08e2b;
      36392: inst = 32'h13e00001;
      36393: inst = 32'hfe0d96a;
      36394: inst = 32'h5be00000;
      36395: inst = 32'h8c50000;
      36396: inst = 32'h24612800;
      36397: inst = 32'h10a0ffff;
      36398: inst = 32'hca0ffe0;
      36399: inst = 32'h24822800;
      36400: inst = 32'h10a00000;
      36401: inst = 32'hca00004;
      36402: inst = 32'h38632800;
      36403: inst = 32'h38842800;
      36404: inst = 32'h10a00000;
      36405: inst = 32'hca08e39;
      36406: inst = 32'h13e00001;
      36407: inst = 32'hfe0d96a;
      36408: inst = 32'h5be00000;
      36409: inst = 32'h8c50000;
      36410: inst = 32'h24612800;
      36411: inst = 32'h10a0ffff;
      36412: inst = 32'hca0ffe0;
      36413: inst = 32'h24822800;
      36414: inst = 32'h10a00000;
      36415: inst = 32'hca00004;
      36416: inst = 32'h38632800;
      36417: inst = 32'h38842800;
      36418: inst = 32'h10a00000;
      36419: inst = 32'hca08e47;
      36420: inst = 32'h13e00001;
      36421: inst = 32'hfe0d96a;
      36422: inst = 32'h5be00000;
      36423: inst = 32'h8c50000;
      36424: inst = 32'h24612800;
      36425: inst = 32'h10a0ffff;
      36426: inst = 32'hca0ffe0;
      36427: inst = 32'h24822800;
      36428: inst = 32'h10a00000;
      36429: inst = 32'hca00004;
      36430: inst = 32'h38632800;
      36431: inst = 32'h38842800;
      36432: inst = 32'h10a00000;
      36433: inst = 32'hca08e55;
      36434: inst = 32'h13e00001;
      36435: inst = 32'hfe0d96a;
      36436: inst = 32'h5be00000;
      36437: inst = 32'h8c50000;
      36438: inst = 32'h24612800;
      36439: inst = 32'h10a0ffff;
      36440: inst = 32'hca0ffe0;
      36441: inst = 32'h24822800;
      36442: inst = 32'h10a00000;
      36443: inst = 32'hca00004;
      36444: inst = 32'h38632800;
      36445: inst = 32'h38842800;
      36446: inst = 32'h10a00000;
      36447: inst = 32'hca08e63;
      36448: inst = 32'h13e00001;
      36449: inst = 32'hfe0d96a;
      36450: inst = 32'h5be00000;
      36451: inst = 32'h8c50000;
      36452: inst = 32'h24612800;
      36453: inst = 32'h10a0ffff;
      36454: inst = 32'hca0ffe0;
      36455: inst = 32'h24822800;
      36456: inst = 32'h10a00000;
      36457: inst = 32'hca00004;
      36458: inst = 32'h38632800;
      36459: inst = 32'h38842800;
      36460: inst = 32'h10a00000;
      36461: inst = 32'hca08e71;
      36462: inst = 32'h13e00001;
      36463: inst = 32'hfe0d96a;
      36464: inst = 32'h5be00000;
      36465: inst = 32'h8c50000;
      36466: inst = 32'h24612800;
      36467: inst = 32'h10a0ffff;
      36468: inst = 32'hca0ffe0;
      36469: inst = 32'h24822800;
      36470: inst = 32'h10a00000;
      36471: inst = 32'hca00004;
      36472: inst = 32'h38632800;
      36473: inst = 32'h38842800;
      36474: inst = 32'h10a00000;
      36475: inst = 32'hca08e7f;
      36476: inst = 32'h13e00001;
      36477: inst = 32'hfe0d96a;
      36478: inst = 32'h5be00000;
      36479: inst = 32'h8c50000;
      36480: inst = 32'h24612800;
      36481: inst = 32'h10a0ffff;
      36482: inst = 32'hca0ffe0;
      36483: inst = 32'h24822800;
      36484: inst = 32'h10a00000;
      36485: inst = 32'hca00004;
      36486: inst = 32'h38632800;
      36487: inst = 32'h38842800;
      36488: inst = 32'h10a00000;
      36489: inst = 32'hca08e8d;
      36490: inst = 32'h13e00001;
      36491: inst = 32'hfe0d96a;
      36492: inst = 32'h5be00000;
      36493: inst = 32'h8c50000;
      36494: inst = 32'h24612800;
      36495: inst = 32'h10a0ffff;
      36496: inst = 32'hca0ffe0;
      36497: inst = 32'h24822800;
      36498: inst = 32'h10a00000;
      36499: inst = 32'hca00004;
      36500: inst = 32'h38632800;
      36501: inst = 32'h38842800;
      36502: inst = 32'h10a00000;
      36503: inst = 32'hca08e9b;
      36504: inst = 32'h13e00001;
      36505: inst = 32'hfe0d96a;
      36506: inst = 32'h5be00000;
      36507: inst = 32'h8c50000;
      36508: inst = 32'h24612800;
      36509: inst = 32'h10a0ffff;
      36510: inst = 32'hca0ffe0;
      36511: inst = 32'h24822800;
      36512: inst = 32'h10a00000;
      36513: inst = 32'hca00004;
      36514: inst = 32'h38632800;
      36515: inst = 32'h38842800;
      36516: inst = 32'h10a00000;
      36517: inst = 32'hca08ea9;
      36518: inst = 32'h13e00001;
      36519: inst = 32'hfe0d96a;
      36520: inst = 32'h5be00000;
      36521: inst = 32'h8c50000;
      36522: inst = 32'h24612800;
      36523: inst = 32'h10a0ffff;
      36524: inst = 32'hca0ffe1;
      36525: inst = 32'h24822800;
      36526: inst = 32'h10a00000;
      36527: inst = 32'hca00004;
      36528: inst = 32'h38632800;
      36529: inst = 32'h38842800;
      36530: inst = 32'h10a00000;
      36531: inst = 32'hca08eb7;
      36532: inst = 32'h13e00001;
      36533: inst = 32'hfe0d96a;
      36534: inst = 32'h5be00000;
      36535: inst = 32'h8c50000;
      36536: inst = 32'h24612800;
      36537: inst = 32'h10a0ffff;
      36538: inst = 32'hca0ffe1;
      36539: inst = 32'h24822800;
      36540: inst = 32'h10a00000;
      36541: inst = 32'hca00004;
      36542: inst = 32'h38632800;
      36543: inst = 32'h38842800;
      36544: inst = 32'h10a00000;
      36545: inst = 32'hca08ec5;
      36546: inst = 32'h13e00001;
      36547: inst = 32'hfe0d96a;
      36548: inst = 32'h5be00000;
      36549: inst = 32'h8c50000;
      36550: inst = 32'h24612800;
      36551: inst = 32'h10a0ffff;
      36552: inst = 32'hca0ffe1;
      36553: inst = 32'h24822800;
      36554: inst = 32'h10a00000;
      36555: inst = 32'hca00004;
      36556: inst = 32'h38632800;
      36557: inst = 32'h38842800;
      36558: inst = 32'h10a00000;
      36559: inst = 32'hca08ed3;
      36560: inst = 32'h13e00001;
      36561: inst = 32'hfe0d96a;
      36562: inst = 32'h5be00000;
      36563: inst = 32'h8c50000;
      36564: inst = 32'h24612800;
      36565: inst = 32'h10a0ffff;
      36566: inst = 32'hca0ffe1;
      36567: inst = 32'h24822800;
      36568: inst = 32'h10a00000;
      36569: inst = 32'hca00004;
      36570: inst = 32'h38632800;
      36571: inst = 32'h38842800;
      36572: inst = 32'h10a00000;
      36573: inst = 32'hca08ee1;
      36574: inst = 32'h13e00001;
      36575: inst = 32'hfe0d96a;
      36576: inst = 32'h5be00000;
      36577: inst = 32'h8c50000;
      36578: inst = 32'h24612800;
      36579: inst = 32'h10a0ffff;
      36580: inst = 32'hca0ffe1;
      36581: inst = 32'h24822800;
      36582: inst = 32'h10a00000;
      36583: inst = 32'hca00004;
      36584: inst = 32'h38632800;
      36585: inst = 32'h38842800;
      36586: inst = 32'h10a00000;
      36587: inst = 32'hca08eef;
      36588: inst = 32'h13e00001;
      36589: inst = 32'hfe0d96a;
      36590: inst = 32'h5be00000;
      36591: inst = 32'h8c50000;
      36592: inst = 32'h24612800;
      36593: inst = 32'h10a0ffff;
      36594: inst = 32'hca0ffe1;
      36595: inst = 32'h24822800;
      36596: inst = 32'h10a00000;
      36597: inst = 32'hca00004;
      36598: inst = 32'h38632800;
      36599: inst = 32'h38842800;
      36600: inst = 32'h10a00000;
      36601: inst = 32'hca08efd;
      36602: inst = 32'h13e00001;
      36603: inst = 32'hfe0d96a;
      36604: inst = 32'h5be00000;
      36605: inst = 32'h8c50000;
      36606: inst = 32'h24612800;
      36607: inst = 32'h10a0ffff;
      36608: inst = 32'hca0ffe1;
      36609: inst = 32'h24822800;
      36610: inst = 32'h10a00000;
      36611: inst = 32'hca00004;
      36612: inst = 32'h38632800;
      36613: inst = 32'h38842800;
      36614: inst = 32'h10a00000;
      36615: inst = 32'hca08f0b;
      36616: inst = 32'h13e00001;
      36617: inst = 32'hfe0d96a;
      36618: inst = 32'h5be00000;
      36619: inst = 32'h8c50000;
      36620: inst = 32'h24612800;
      36621: inst = 32'h10a0ffff;
      36622: inst = 32'hca0ffe1;
      36623: inst = 32'h24822800;
      36624: inst = 32'h10a00000;
      36625: inst = 32'hca00004;
      36626: inst = 32'h38632800;
      36627: inst = 32'h38842800;
      36628: inst = 32'h10a00000;
      36629: inst = 32'hca08f19;
      36630: inst = 32'h13e00001;
      36631: inst = 32'hfe0d96a;
      36632: inst = 32'h5be00000;
      36633: inst = 32'h8c50000;
      36634: inst = 32'h24612800;
      36635: inst = 32'h10a0ffff;
      36636: inst = 32'hca0ffe1;
      36637: inst = 32'h24822800;
      36638: inst = 32'h10a00000;
      36639: inst = 32'hca00004;
      36640: inst = 32'h38632800;
      36641: inst = 32'h38842800;
      36642: inst = 32'h10a00000;
      36643: inst = 32'hca08f27;
      36644: inst = 32'h13e00001;
      36645: inst = 32'hfe0d96a;
      36646: inst = 32'h5be00000;
      36647: inst = 32'h8c50000;
      36648: inst = 32'h24612800;
      36649: inst = 32'h10a0ffff;
      36650: inst = 32'hca0ffe1;
      36651: inst = 32'h24822800;
      36652: inst = 32'h10a00000;
      36653: inst = 32'hca00004;
      36654: inst = 32'h38632800;
      36655: inst = 32'h38842800;
      36656: inst = 32'h10a00000;
      36657: inst = 32'hca08f35;
      36658: inst = 32'h13e00001;
      36659: inst = 32'hfe0d96a;
      36660: inst = 32'h5be00000;
      36661: inst = 32'h8c50000;
      36662: inst = 32'h24612800;
      36663: inst = 32'h10a0ffff;
      36664: inst = 32'hca0ffe1;
      36665: inst = 32'h24822800;
      36666: inst = 32'h10a00000;
      36667: inst = 32'hca00004;
      36668: inst = 32'h38632800;
      36669: inst = 32'h38842800;
      36670: inst = 32'h10a00000;
      36671: inst = 32'hca08f43;
      36672: inst = 32'h13e00001;
      36673: inst = 32'hfe0d96a;
      36674: inst = 32'h5be00000;
      36675: inst = 32'h8c50000;
      36676: inst = 32'h24612800;
      36677: inst = 32'h10a0ffff;
      36678: inst = 32'hca0ffe1;
      36679: inst = 32'h24822800;
      36680: inst = 32'h10a00000;
      36681: inst = 32'hca00004;
      36682: inst = 32'h38632800;
      36683: inst = 32'h38842800;
      36684: inst = 32'h10a00000;
      36685: inst = 32'hca08f51;
      36686: inst = 32'h13e00001;
      36687: inst = 32'hfe0d96a;
      36688: inst = 32'h5be00000;
      36689: inst = 32'h8c50000;
      36690: inst = 32'h24612800;
      36691: inst = 32'h10a0ffff;
      36692: inst = 32'hca0ffe1;
      36693: inst = 32'h24822800;
      36694: inst = 32'h10a00000;
      36695: inst = 32'hca00004;
      36696: inst = 32'h38632800;
      36697: inst = 32'h38842800;
      36698: inst = 32'h10a00000;
      36699: inst = 32'hca08f5f;
      36700: inst = 32'h13e00001;
      36701: inst = 32'hfe0d96a;
      36702: inst = 32'h5be00000;
      36703: inst = 32'h8c50000;
      36704: inst = 32'h24612800;
      36705: inst = 32'h10a0ffff;
      36706: inst = 32'hca0ffe1;
      36707: inst = 32'h24822800;
      36708: inst = 32'h10a00000;
      36709: inst = 32'hca00004;
      36710: inst = 32'h38632800;
      36711: inst = 32'h38842800;
      36712: inst = 32'h10a00000;
      36713: inst = 32'hca08f6d;
      36714: inst = 32'h13e00001;
      36715: inst = 32'hfe0d96a;
      36716: inst = 32'h5be00000;
      36717: inst = 32'h8c50000;
      36718: inst = 32'h24612800;
      36719: inst = 32'h10a0ffff;
      36720: inst = 32'hca0ffe1;
      36721: inst = 32'h24822800;
      36722: inst = 32'h10a00000;
      36723: inst = 32'hca00004;
      36724: inst = 32'h38632800;
      36725: inst = 32'h38842800;
      36726: inst = 32'h10a00000;
      36727: inst = 32'hca08f7b;
      36728: inst = 32'h13e00001;
      36729: inst = 32'hfe0d96a;
      36730: inst = 32'h5be00000;
      36731: inst = 32'h8c50000;
      36732: inst = 32'h24612800;
      36733: inst = 32'h10a0ffff;
      36734: inst = 32'hca0ffe1;
      36735: inst = 32'h24822800;
      36736: inst = 32'h10a00000;
      36737: inst = 32'hca00004;
      36738: inst = 32'h38632800;
      36739: inst = 32'h38842800;
      36740: inst = 32'h10a00000;
      36741: inst = 32'hca08f89;
      36742: inst = 32'h13e00001;
      36743: inst = 32'hfe0d96a;
      36744: inst = 32'h5be00000;
      36745: inst = 32'h8c50000;
      36746: inst = 32'h24612800;
      36747: inst = 32'h10a0ffff;
      36748: inst = 32'hca0ffe1;
      36749: inst = 32'h24822800;
      36750: inst = 32'h10a00000;
      36751: inst = 32'hca00004;
      36752: inst = 32'h38632800;
      36753: inst = 32'h38842800;
      36754: inst = 32'h10a00000;
      36755: inst = 32'hca08f97;
      36756: inst = 32'h13e00001;
      36757: inst = 32'hfe0d96a;
      36758: inst = 32'h5be00000;
      36759: inst = 32'h8c50000;
      36760: inst = 32'h24612800;
      36761: inst = 32'h10a0ffff;
      36762: inst = 32'hca0ffe1;
      36763: inst = 32'h24822800;
      36764: inst = 32'h10a00000;
      36765: inst = 32'hca00004;
      36766: inst = 32'h38632800;
      36767: inst = 32'h38842800;
      36768: inst = 32'h10a00000;
      36769: inst = 32'hca08fa5;
      36770: inst = 32'h13e00001;
      36771: inst = 32'hfe0d96a;
      36772: inst = 32'h5be00000;
      36773: inst = 32'h8c50000;
      36774: inst = 32'h24612800;
      36775: inst = 32'h10a0ffff;
      36776: inst = 32'hca0ffe1;
      36777: inst = 32'h24822800;
      36778: inst = 32'h10a00000;
      36779: inst = 32'hca00004;
      36780: inst = 32'h38632800;
      36781: inst = 32'h38842800;
      36782: inst = 32'h10a00000;
      36783: inst = 32'hca08fb3;
      36784: inst = 32'h13e00001;
      36785: inst = 32'hfe0d96a;
      36786: inst = 32'h5be00000;
      36787: inst = 32'h8c50000;
      36788: inst = 32'h24612800;
      36789: inst = 32'h10a0ffff;
      36790: inst = 32'hca0ffe1;
      36791: inst = 32'h24822800;
      36792: inst = 32'h10a00000;
      36793: inst = 32'hca00004;
      36794: inst = 32'h38632800;
      36795: inst = 32'h38842800;
      36796: inst = 32'h10a00000;
      36797: inst = 32'hca08fc1;
      36798: inst = 32'h13e00001;
      36799: inst = 32'hfe0d96a;
      36800: inst = 32'h5be00000;
      36801: inst = 32'h8c50000;
      36802: inst = 32'h24612800;
      36803: inst = 32'h10a0ffff;
      36804: inst = 32'hca0ffe1;
      36805: inst = 32'h24822800;
      36806: inst = 32'h10a00000;
      36807: inst = 32'hca00004;
      36808: inst = 32'h38632800;
      36809: inst = 32'h38842800;
      36810: inst = 32'h10a00000;
      36811: inst = 32'hca08fcf;
      36812: inst = 32'h13e00001;
      36813: inst = 32'hfe0d96a;
      36814: inst = 32'h5be00000;
      36815: inst = 32'h8c50000;
      36816: inst = 32'h24612800;
      36817: inst = 32'h10a0ffff;
      36818: inst = 32'hca0ffe1;
      36819: inst = 32'h24822800;
      36820: inst = 32'h10a00000;
      36821: inst = 32'hca00004;
      36822: inst = 32'h38632800;
      36823: inst = 32'h38842800;
      36824: inst = 32'h10a00000;
      36825: inst = 32'hca08fdd;
      36826: inst = 32'h13e00001;
      36827: inst = 32'hfe0d96a;
      36828: inst = 32'h5be00000;
      36829: inst = 32'h8c50000;
      36830: inst = 32'h24612800;
      36831: inst = 32'h10a0ffff;
      36832: inst = 32'hca0ffe1;
      36833: inst = 32'h24822800;
      36834: inst = 32'h10a00000;
      36835: inst = 32'hca00004;
      36836: inst = 32'h38632800;
      36837: inst = 32'h38842800;
      36838: inst = 32'h10a00000;
      36839: inst = 32'hca08feb;
      36840: inst = 32'h13e00001;
      36841: inst = 32'hfe0d96a;
      36842: inst = 32'h5be00000;
      36843: inst = 32'h8c50000;
      36844: inst = 32'h24612800;
      36845: inst = 32'h10a0ffff;
      36846: inst = 32'hca0ffe1;
      36847: inst = 32'h24822800;
      36848: inst = 32'h10a00000;
      36849: inst = 32'hca00004;
      36850: inst = 32'h38632800;
      36851: inst = 32'h38842800;
      36852: inst = 32'h10a00000;
      36853: inst = 32'hca08ff9;
      36854: inst = 32'h13e00001;
      36855: inst = 32'hfe0d96a;
      36856: inst = 32'h5be00000;
      36857: inst = 32'h8c50000;
      36858: inst = 32'h24612800;
      36859: inst = 32'h10a0ffff;
      36860: inst = 32'hca0ffe1;
      36861: inst = 32'h24822800;
      36862: inst = 32'h10a00000;
      36863: inst = 32'hca00004;
      36864: inst = 32'h38632800;
      36865: inst = 32'h38842800;
      36866: inst = 32'h10a00000;
      36867: inst = 32'hca09007;
      36868: inst = 32'h13e00001;
      36869: inst = 32'hfe0d96a;
      36870: inst = 32'h5be00000;
      36871: inst = 32'h8c50000;
      36872: inst = 32'h24612800;
      36873: inst = 32'h10a0ffff;
      36874: inst = 32'hca0ffe1;
      36875: inst = 32'h24822800;
      36876: inst = 32'h10a00000;
      36877: inst = 32'hca00004;
      36878: inst = 32'h38632800;
      36879: inst = 32'h38842800;
      36880: inst = 32'h10a00000;
      36881: inst = 32'hca09015;
      36882: inst = 32'h13e00001;
      36883: inst = 32'hfe0d96a;
      36884: inst = 32'h5be00000;
      36885: inst = 32'h8c50000;
      36886: inst = 32'h24612800;
      36887: inst = 32'h10a0ffff;
      36888: inst = 32'hca0ffe1;
      36889: inst = 32'h24822800;
      36890: inst = 32'h10a00000;
      36891: inst = 32'hca00004;
      36892: inst = 32'h38632800;
      36893: inst = 32'h38842800;
      36894: inst = 32'h10a00000;
      36895: inst = 32'hca09023;
      36896: inst = 32'h13e00001;
      36897: inst = 32'hfe0d96a;
      36898: inst = 32'h5be00000;
      36899: inst = 32'h8c50000;
      36900: inst = 32'h24612800;
      36901: inst = 32'h10a0ffff;
      36902: inst = 32'hca0ffe1;
      36903: inst = 32'h24822800;
      36904: inst = 32'h10a00000;
      36905: inst = 32'hca00004;
      36906: inst = 32'h38632800;
      36907: inst = 32'h38842800;
      36908: inst = 32'h10a00000;
      36909: inst = 32'hca09031;
      36910: inst = 32'h13e00001;
      36911: inst = 32'hfe0d96a;
      36912: inst = 32'h5be00000;
      36913: inst = 32'h8c50000;
      36914: inst = 32'h24612800;
      36915: inst = 32'h10a0ffff;
      36916: inst = 32'hca0ffe1;
      36917: inst = 32'h24822800;
      36918: inst = 32'h10a00000;
      36919: inst = 32'hca00004;
      36920: inst = 32'h38632800;
      36921: inst = 32'h38842800;
      36922: inst = 32'h10a00000;
      36923: inst = 32'hca0903f;
      36924: inst = 32'h13e00001;
      36925: inst = 32'hfe0d96a;
      36926: inst = 32'h5be00000;
      36927: inst = 32'h8c50000;
      36928: inst = 32'h24612800;
      36929: inst = 32'h10a0ffff;
      36930: inst = 32'hca0ffe1;
      36931: inst = 32'h24822800;
      36932: inst = 32'h10a00000;
      36933: inst = 32'hca00004;
      36934: inst = 32'h38632800;
      36935: inst = 32'h38842800;
      36936: inst = 32'h10a00000;
      36937: inst = 32'hca0904d;
      36938: inst = 32'h13e00001;
      36939: inst = 32'hfe0d96a;
      36940: inst = 32'h5be00000;
      36941: inst = 32'h8c50000;
      36942: inst = 32'h24612800;
      36943: inst = 32'h10a0ffff;
      36944: inst = 32'hca0ffe1;
      36945: inst = 32'h24822800;
      36946: inst = 32'h10a00000;
      36947: inst = 32'hca00004;
      36948: inst = 32'h38632800;
      36949: inst = 32'h38842800;
      36950: inst = 32'h10a00000;
      36951: inst = 32'hca0905b;
      36952: inst = 32'h13e00001;
      36953: inst = 32'hfe0d96a;
      36954: inst = 32'h5be00000;
      36955: inst = 32'h8c50000;
      36956: inst = 32'h24612800;
      36957: inst = 32'h10a0ffff;
      36958: inst = 32'hca0ffe1;
      36959: inst = 32'h24822800;
      36960: inst = 32'h10a00000;
      36961: inst = 32'hca00004;
      36962: inst = 32'h38632800;
      36963: inst = 32'h38842800;
      36964: inst = 32'h10a00000;
      36965: inst = 32'hca09069;
      36966: inst = 32'h13e00001;
      36967: inst = 32'hfe0d96a;
      36968: inst = 32'h5be00000;
      36969: inst = 32'h8c50000;
      36970: inst = 32'h24612800;
      36971: inst = 32'h10a0ffff;
      36972: inst = 32'hca0ffe1;
      36973: inst = 32'h24822800;
      36974: inst = 32'h10a00000;
      36975: inst = 32'hca00004;
      36976: inst = 32'h38632800;
      36977: inst = 32'h38842800;
      36978: inst = 32'h10a00000;
      36979: inst = 32'hca09077;
      36980: inst = 32'h13e00001;
      36981: inst = 32'hfe0d96a;
      36982: inst = 32'h5be00000;
      36983: inst = 32'h8c50000;
      36984: inst = 32'h24612800;
      36985: inst = 32'h10a0ffff;
      36986: inst = 32'hca0ffe1;
      36987: inst = 32'h24822800;
      36988: inst = 32'h10a00000;
      36989: inst = 32'hca00004;
      36990: inst = 32'h38632800;
      36991: inst = 32'h38842800;
      36992: inst = 32'h10a00000;
      36993: inst = 32'hca09085;
      36994: inst = 32'h13e00001;
      36995: inst = 32'hfe0d96a;
      36996: inst = 32'h5be00000;
      36997: inst = 32'h8c50000;
      36998: inst = 32'h24612800;
      36999: inst = 32'h10a0ffff;
      37000: inst = 32'hca0ffe1;
      37001: inst = 32'h24822800;
      37002: inst = 32'h10a00000;
      37003: inst = 32'hca00004;
      37004: inst = 32'h38632800;
      37005: inst = 32'h38842800;
      37006: inst = 32'h10a00000;
      37007: inst = 32'hca09093;
      37008: inst = 32'h13e00001;
      37009: inst = 32'hfe0d96a;
      37010: inst = 32'h5be00000;
      37011: inst = 32'h8c50000;
      37012: inst = 32'h24612800;
      37013: inst = 32'h10a0ffff;
      37014: inst = 32'hca0ffe1;
      37015: inst = 32'h24822800;
      37016: inst = 32'h10a00000;
      37017: inst = 32'hca00004;
      37018: inst = 32'h38632800;
      37019: inst = 32'h38842800;
      37020: inst = 32'h10a00000;
      37021: inst = 32'hca090a1;
      37022: inst = 32'h13e00001;
      37023: inst = 32'hfe0d96a;
      37024: inst = 32'h5be00000;
      37025: inst = 32'h8c50000;
      37026: inst = 32'h24612800;
      37027: inst = 32'h10a0ffff;
      37028: inst = 32'hca0ffe1;
      37029: inst = 32'h24822800;
      37030: inst = 32'h10a00000;
      37031: inst = 32'hca00004;
      37032: inst = 32'h38632800;
      37033: inst = 32'h38842800;
      37034: inst = 32'h10a00000;
      37035: inst = 32'hca090af;
      37036: inst = 32'h13e00001;
      37037: inst = 32'hfe0d96a;
      37038: inst = 32'h5be00000;
      37039: inst = 32'h8c50000;
      37040: inst = 32'h24612800;
      37041: inst = 32'h10a0ffff;
      37042: inst = 32'hca0ffe1;
      37043: inst = 32'h24822800;
      37044: inst = 32'h10a00000;
      37045: inst = 32'hca00004;
      37046: inst = 32'h38632800;
      37047: inst = 32'h38842800;
      37048: inst = 32'h10a00000;
      37049: inst = 32'hca090bd;
      37050: inst = 32'h13e00001;
      37051: inst = 32'hfe0d96a;
      37052: inst = 32'h5be00000;
      37053: inst = 32'h8c50000;
      37054: inst = 32'h24612800;
      37055: inst = 32'h10a0ffff;
      37056: inst = 32'hca0ffe1;
      37057: inst = 32'h24822800;
      37058: inst = 32'h10a00000;
      37059: inst = 32'hca00004;
      37060: inst = 32'h38632800;
      37061: inst = 32'h38842800;
      37062: inst = 32'h10a00000;
      37063: inst = 32'hca090cb;
      37064: inst = 32'h13e00001;
      37065: inst = 32'hfe0d96a;
      37066: inst = 32'h5be00000;
      37067: inst = 32'h8c50000;
      37068: inst = 32'h24612800;
      37069: inst = 32'h10a0ffff;
      37070: inst = 32'hca0ffe1;
      37071: inst = 32'h24822800;
      37072: inst = 32'h10a00000;
      37073: inst = 32'hca00004;
      37074: inst = 32'h38632800;
      37075: inst = 32'h38842800;
      37076: inst = 32'h10a00000;
      37077: inst = 32'hca090d9;
      37078: inst = 32'h13e00001;
      37079: inst = 32'hfe0d96a;
      37080: inst = 32'h5be00000;
      37081: inst = 32'h8c50000;
      37082: inst = 32'h24612800;
      37083: inst = 32'h10a0ffff;
      37084: inst = 32'hca0ffe1;
      37085: inst = 32'h24822800;
      37086: inst = 32'h10a00000;
      37087: inst = 32'hca00004;
      37088: inst = 32'h38632800;
      37089: inst = 32'h38842800;
      37090: inst = 32'h10a00000;
      37091: inst = 32'hca090e7;
      37092: inst = 32'h13e00001;
      37093: inst = 32'hfe0d96a;
      37094: inst = 32'h5be00000;
      37095: inst = 32'h8c50000;
      37096: inst = 32'h24612800;
      37097: inst = 32'h10a0ffff;
      37098: inst = 32'hca0ffe1;
      37099: inst = 32'h24822800;
      37100: inst = 32'h10a00000;
      37101: inst = 32'hca00004;
      37102: inst = 32'h38632800;
      37103: inst = 32'h38842800;
      37104: inst = 32'h10a00000;
      37105: inst = 32'hca090f5;
      37106: inst = 32'h13e00001;
      37107: inst = 32'hfe0d96a;
      37108: inst = 32'h5be00000;
      37109: inst = 32'h8c50000;
      37110: inst = 32'h24612800;
      37111: inst = 32'h10a0ffff;
      37112: inst = 32'hca0ffe1;
      37113: inst = 32'h24822800;
      37114: inst = 32'h10a00000;
      37115: inst = 32'hca00004;
      37116: inst = 32'h38632800;
      37117: inst = 32'h38842800;
      37118: inst = 32'h10a00000;
      37119: inst = 32'hca09103;
      37120: inst = 32'h13e00001;
      37121: inst = 32'hfe0d96a;
      37122: inst = 32'h5be00000;
      37123: inst = 32'h8c50000;
      37124: inst = 32'h24612800;
      37125: inst = 32'h10a0ffff;
      37126: inst = 32'hca0ffe1;
      37127: inst = 32'h24822800;
      37128: inst = 32'h10a00000;
      37129: inst = 32'hca00004;
      37130: inst = 32'h38632800;
      37131: inst = 32'h38842800;
      37132: inst = 32'h10a00000;
      37133: inst = 32'hca09111;
      37134: inst = 32'h13e00001;
      37135: inst = 32'hfe0d96a;
      37136: inst = 32'h5be00000;
      37137: inst = 32'h8c50000;
      37138: inst = 32'h24612800;
      37139: inst = 32'h10a0ffff;
      37140: inst = 32'hca0ffe1;
      37141: inst = 32'h24822800;
      37142: inst = 32'h10a00000;
      37143: inst = 32'hca00004;
      37144: inst = 32'h38632800;
      37145: inst = 32'h38842800;
      37146: inst = 32'h10a00000;
      37147: inst = 32'hca0911f;
      37148: inst = 32'h13e00001;
      37149: inst = 32'hfe0d96a;
      37150: inst = 32'h5be00000;
      37151: inst = 32'h8c50000;
      37152: inst = 32'h24612800;
      37153: inst = 32'h10a0ffff;
      37154: inst = 32'hca0ffe1;
      37155: inst = 32'h24822800;
      37156: inst = 32'h10a00000;
      37157: inst = 32'hca00004;
      37158: inst = 32'h38632800;
      37159: inst = 32'h38842800;
      37160: inst = 32'h10a00000;
      37161: inst = 32'hca0912d;
      37162: inst = 32'h13e00001;
      37163: inst = 32'hfe0d96a;
      37164: inst = 32'h5be00000;
      37165: inst = 32'h8c50000;
      37166: inst = 32'h24612800;
      37167: inst = 32'h10a0ffff;
      37168: inst = 32'hca0ffe1;
      37169: inst = 32'h24822800;
      37170: inst = 32'h10a00000;
      37171: inst = 32'hca00004;
      37172: inst = 32'h38632800;
      37173: inst = 32'h38842800;
      37174: inst = 32'h10a00000;
      37175: inst = 32'hca0913b;
      37176: inst = 32'h13e00001;
      37177: inst = 32'hfe0d96a;
      37178: inst = 32'h5be00000;
      37179: inst = 32'h8c50000;
      37180: inst = 32'h24612800;
      37181: inst = 32'h10a0ffff;
      37182: inst = 32'hca0ffe1;
      37183: inst = 32'h24822800;
      37184: inst = 32'h10a00000;
      37185: inst = 32'hca00004;
      37186: inst = 32'h38632800;
      37187: inst = 32'h38842800;
      37188: inst = 32'h10a00000;
      37189: inst = 32'hca09149;
      37190: inst = 32'h13e00001;
      37191: inst = 32'hfe0d96a;
      37192: inst = 32'h5be00000;
      37193: inst = 32'h8c50000;
      37194: inst = 32'h24612800;
      37195: inst = 32'h10a0ffff;
      37196: inst = 32'hca0ffe1;
      37197: inst = 32'h24822800;
      37198: inst = 32'h10a00000;
      37199: inst = 32'hca00004;
      37200: inst = 32'h38632800;
      37201: inst = 32'h38842800;
      37202: inst = 32'h10a00000;
      37203: inst = 32'hca09157;
      37204: inst = 32'h13e00001;
      37205: inst = 32'hfe0d96a;
      37206: inst = 32'h5be00000;
      37207: inst = 32'h8c50000;
      37208: inst = 32'h24612800;
      37209: inst = 32'h10a0ffff;
      37210: inst = 32'hca0ffe1;
      37211: inst = 32'h24822800;
      37212: inst = 32'h10a00000;
      37213: inst = 32'hca00004;
      37214: inst = 32'h38632800;
      37215: inst = 32'h38842800;
      37216: inst = 32'h10a00000;
      37217: inst = 32'hca09165;
      37218: inst = 32'h13e00001;
      37219: inst = 32'hfe0d96a;
      37220: inst = 32'h5be00000;
      37221: inst = 32'h8c50000;
      37222: inst = 32'h24612800;
      37223: inst = 32'h10a0ffff;
      37224: inst = 32'hca0ffe1;
      37225: inst = 32'h24822800;
      37226: inst = 32'h10a00000;
      37227: inst = 32'hca00004;
      37228: inst = 32'h38632800;
      37229: inst = 32'h38842800;
      37230: inst = 32'h10a00000;
      37231: inst = 32'hca09173;
      37232: inst = 32'h13e00001;
      37233: inst = 32'hfe0d96a;
      37234: inst = 32'h5be00000;
      37235: inst = 32'h8c50000;
      37236: inst = 32'h24612800;
      37237: inst = 32'h10a0ffff;
      37238: inst = 32'hca0ffe1;
      37239: inst = 32'h24822800;
      37240: inst = 32'h10a00000;
      37241: inst = 32'hca00004;
      37242: inst = 32'h38632800;
      37243: inst = 32'h38842800;
      37244: inst = 32'h10a00000;
      37245: inst = 32'hca09181;
      37246: inst = 32'h13e00001;
      37247: inst = 32'hfe0d96a;
      37248: inst = 32'h5be00000;
      37249: inst = 32'h8c50000;
      37250: inst = 32'h24612800;
      37251: inst = 32'h10a0ffff;
      37252: inst = 32'hca0ffe1;
      37253: inst = 32'h24822800;
      37254: inst = 32'h10a00000;
      37255: inst = 32'hca00004;
      37256: inst = 32'h38632800;
      37257: inst = 32'h38842800;
      37258: inst = 32'h10a00000;
      37259: inst = 32'hca0918f;
      37260: inst = 32'h13e00001;
      37261: inst = 32'hfe0d96a;
      37262: inst = 32'h5be00000;
      37263: inst = 32'h8c50000;
      37264: inst = 32'h24612800;
      37265: inst = 32'h10a0ffff;
      37266: inst = 32'hca0ffe1;
      37267: inst = 32'h24822800;
      37268: inst = 32'h10a00000;
      37269: inst = 32'hca00004;
      37270: inst = 32'h38632800;
      37271: inst = 32'h38842800;
      37272: inst = 32'h10a00000;
      37273: inst = 32'hca0919d;
      37274: inst = 32'h13e00001;
      37275: inst = 32'hfe0d96a;
      37276: inst = 32'h5be00000;
      37277: inst = 32'h8c50000;
      37278: inst = 32'h24612800;
      37279: inst = 32'h10a0ffff;
      37280: inst = 32'hca0ffe1;
      37281: inst = 32'h24822800;
      37282: inst = 32'h10a00000;
      37283: inst = 32'hca00004;
      37284: inst = 32'h38632800;
      37285: inst = 32'h38842800;
      37286: inst = 32'h10a00000;
      37287: inst = 32'hca091ab;
      37288: inst = 32'h13e00001;
      37289: inst = 32'hfe0d96a;
      37290: inst = 32'h5be00000;
      37291: inst = 32'h8c50000;
      37292: inst = 32'h24612800;
      37293: inst = 32'h10a0ffff;
      37294: inst = 32'hca0ffe1;
      37295: inst = 32'h24822800;
      37296: inst = 32'h10a00000;
      37297: inst = 32'hca00004;
      37298: inst = 32'h38632800;
      37299: inst = 32'h38842800;
      37300: inst = 32'h10a00000;
      37301: inst = 32'hca091b9;
      37302: inst = 32'h13e00001;
      37303: inst = 32'hfe0d96a;
      37304: inst = 32'h5be00000;
      37305: inst = 32'h8c50000;
      37306: inst = 32'h24612800;
      37307: inst = 32'h10a0ffff;
      37308: inst = 32'hca0ffe1;
      37309: inst = 32'h24822800;
      37310: inst = 32'h10a00000;
      37311: inst = 32'hca00004;
      37312: inst = 32'h38632800;
      37313: inst = 32'h38842800;
      37314: inst = 32'h10a00000;
      37315: inst = 32'hca091c7;
      37316: inst = 32'h13e00001;
      37317: inst = 32'hfe0d96a;
      37318: inst = 32'h5be00000;
      37319: inst = 32'h8c50000;
      37320: inst = 32'h24612800;
      37321: inst = 32'h10a0ffff;
      37322: inst = 32'hca0ffe1;
      37323: inst = 32'h24822800;
      37324: inst = 32'h10a00000;
      37325: inst = 32'hca00004;
      37326: inst = 32'h38632800;
      37327: inst = 32'h38842800;
      37328: inst = 32'h10a00000;
      37329: inst = 32'hca091d5;
      37330: inst = 32'h13e00001;
      37331: inst = 32'hfe0d96a;
      37332: inst = 32'h5be00000;
      37333: inst = 32'h8c50000;
      37334: inst = 32'h24612800;
      37335: inst = 32'h10a0ffff;
      37336: inst = 32'hca0ffe1;
      37337: inst = 32'h24822800;
      37338: inst = 32'h10a00000;
      37339: inst = 32'hca00004;
      37340: inst = 32'h38632800;
      37341: inst = 32'h38842800;
      37342: inst = 32'h10a00000;
      37343: inst = 32'hca091e3;
      37344: inst = 32'h13e00001;
      37345: inst = 32'hfe0d96a;
      37346: inst = 32'h5be00000;
      37347: inst = 32'h8c50000;
      37348: inst = 32'h24612800;
      37349: inst = 32'h10a0ffff;
      37350: inst = 32'hca0ffe1;
      37351: inst = 32'h24822800;
      37352: inst = 32'h10a00000;
      37353: inst = 32'hca00004;
      37354: inst = 32'h38632800;
      37355: inst = 32'h38842800;
      37356: inst = 32'h10a00000;
      37357: inst = 32'hca091f1;
      37358: inst = 32'h13e00001;
      37359: inst = 32'hfe0d96a;
      37360: inst = 32'h5be00000;
      37361: inst = 32'h8c50000;
      37362: inst = 32'h24612800;
      37363: inst = 32'h10a0ffff;
      37364: inst = 32'hca0ffe1;
      37365: inst = 32'h24822800;
      37366: inst = 32'h10a00000;
      37367: inst = 32'hca00004;
      37368: inst = 32'h38632800;
      37369: inst = 32'h38842800;
      37370: inst = 32'h10a00000;
      37371: inst = 32'hca091ff;
      37372: inst = 32'h13e00001;
      37373: inst = 32'hfe0d96a;
      37374: inst = 32'h5be00000;
      37375: inst = 32'h8c50000;
      37376: inst = 32'h24612800;
      37377: inst = 32'h10a0ffff;
      37378: inst = 32'hca0ffe1;
      37379: inst = 32'h24822800;
      37380: inst = 32'h10a00000;
      37381: inst = 32'hca00004;
      37382: inst = 32'h38632800;
      37383: inst = 32'h38842800;
      37384: inst = 32'h10a00000;
      37385: inst = 32'hca0920d;
      37386: inst = 32'h13e00001;
      37387: inst = 32'hfe0d96a;
      37388: inst = 32'h5be00000;
      37389: inst = 32'h8c50000;
      37390: inst = 32'h24612800;
      37391: inst = 32'h10a0ffff;
      37392: inst = 32'hca0ffe1;
      37393: inst = 32'h24822800;
      37394: inst = 32'h10a00000;
      37395: inst = 32'hca00004;
      37396: inst = 32'h38632800;
      37397: inst = 32'h38842800;
      37398: inst = 32'h10a00000;
      37399: inst = 32'hca0921b;
      37400: inst = 32'h13e00001;
      37401: inst = 32'hfe0d96a;
      37402: inst = 32'h5be00000;
      37403: inst = 32'h8c50000;
      37404: inst = 32'h24612800;
      37405: inst = 32'h10a0ffff;
      37406: inst = 32'hca0ffe1;
      37407: inst = 32'h24822800;
      37408: inst = 32'h10a00000;
      37409: inst = 32'hca00004;
      37410: inst = 32'h38632800;
      37411: inst = 32'h38842800;
      37412: inst = 32'h10a00000;
      37413: inst = 32'hca09229;
      37414: inst = 32'h13e00001;
      37415: inst = 32'hfe0d96a;
      37416: inst = 32'h5be00000;
      37417: inst = 32'h8c50000;
      37418: inst = 32'h24612800;
      37419: inst = 32'h10a0ffff;
      37420: inst = 32'hca0ffe1;
      37421: inst = 32'h24822800;
      37422: inst = 32'h10a00000;
      37423: inst = 32'hca00004;
      37424: inst = 32'h38632800;
      37425: inst = 32'h38842800;
      37426: inst = 32'h10a00000;
      37427: inst = 32'hca09237;
      37428: inst = 32'h13e00001;
      37429: inst = 32'hfe0d96a;
      37430: inst = 32'h5be00000;
      37431: inst = 32'h8c50000;
      37432: inst = 32'h24612800;
      37433: inst = 32'h10a0ffff;
      37434: inst = 32'hca0ffe1;
      37435: inst = 32'h24822800;
      37436: inst = 32'h10a00000;
      37437: inst = 32'hca00004;
      37438: inst = 32'h38632800;
      37439: inst = 32'h38842800;
      37440: inst = 32'h10a00000;
      37441: inst = 32'hca09245;
      37442: inst = 32'h13e00001;
      37443: inst = 32'hfe0d96a;
      37444: inst = 32'h5be00000;
      37445: inst = 32'h8c50000;
      37446: inst = 32'h24612800;
      37447: inst = 32'h10a0ffff;
      37448: inst = 32'hca0ffe1;
      37449: inst = 32'h24822800;
      37450: inst = 32'h10a00000;
      37451: inst = 32'hca00004;
      37452: inst = 32'h38632800;
      37453: inst = 32'h38842800;
      37454: inst = 32'h10a00000;
      37455: inst = 32'hca09253;
      37456: inst = 32'h13e00001;
      37457: inst = 32'hfe0d96a;
      37458: inst = 32'h5be00000;
      37459: inst = 32'h8c50000;
      37460: inst = 32'h24612800;
      37461: inst = 32'h10a0ffff;
      37462: inst = 32'hca0ffe1;
      37463: inst = 32'h24822800;
      37464: inst = 32'h10a00000;
      37465: inst = 32'hca00004;
      37466: inst = 32'h38632800;
      37467: inst = 32'h38842800;
      37468: inst = 32'h10a00000;
      37469: inst = 32'hca09261;
      37470: inst = 32'h13e00001;
      37471: inst = 32'hfe0d96a;
      37472: inst = 32'h5be00000;
      37473: inst = 32'h8c50000;
      37474: inst = 32'h24612800;
      37475: inst = 32'h10a0ffff;
      37476: inst = 32'hca0ffe1;
      37477: inst = 32'h24822800;
      37478: inst = 32'h10a00000;
      37479: inst = 32'hca00004;
      37480: inst = 32'h38632800;
      37481: inst = 32'h38842800;
      37482: inst = 32'h10a00000;
      37483: inst = 32'hca0926f;
      37484: inst = 32'h13e00001;
      37485: inst = 32'hfe0d96a;
      37486: inst = 32'h5be00000;
      37487: inst = 32'h8c50000;
      37488: inst = 32'h24612800;
      37489: inst = 32'h10a0ffff;
      37490: inst = 32'hca0ffe1;
      37491: inst = 32'h24822800;
      37492: inst = 32'h10a00000;
      37493: inst = 32'hca00004;
      37494: inst = 32'h38632800;
      37495: inst = 32'h38842800;
      37496: inst = 32'h10a00000;
      37497: inst = 32'hca0927d;
      37498: inst = 32'h13e00001;
      37499: inst = 32'hfe0d96a;
      37500: inst = 32'h5be00000;
      37501: inst = 32'h8c50000;
      37502: inst = 32'h24612800;
      37503: inst = 32'h10a0ffff;
      37504: inst = 32'hca0ffe1;
      37505: inst = 32'h24822800;
      37506: inst = 32'h10a00000;
      37507: inst = 32'hca00004;
      37508: inst = 32'h38632800;
      37509: inst = 32'h38842800;
      37510: inst = 32'h10a00000;
      37511: inst = 32'hca0928b;
      37512: inst = 32'h13e00001;
      37513: inst = 32'hfe0d96a;
      37514: inst = 32'h5be00000;
      37515: inst = 32'h8c50000;
      37516: inst = 32'h24612800;
      37517: inst = 32'h10a0ffff;
      37518: inst = 32'hca0ffe1;
      37519: inst = 32'h24822800;
      37520: inst = 32'h10a00000;
      37521: inst = 32'hca00004;
      37522: inst = 32'h38632800;
      37523: inst = 32'h38842800;
      37524: inst = 32'h10a00000;
      37525: inst = 32'hca09299;
      37526: inst = 32'h13e00001;
      37527: inst = 32'hfe0d96a;
      37528: inst = 32'h5be00000;
      37529: inst = 32'h8c50000;
      37530: inst = 32'h24612800;
      37531: inst = 32'h10a0ffff;
      37532: inst = 32'hca0ffe1;
      37533: inst = 32'h24822800;
      37534: inst = 32'h10a00000;
      37535: inst = 32'hca00004;
      37536: inst = 32'h38632800;
      37537: inst = 32'h38842800;
      37538: inst = 32'h10a00000;
      37539: inst = 32'hca092a7;
      37540: inst = 32'h13e00001;
      37541: inst = 32'hfe0d96a;
      37542: inst = 32'h5be00000;
      37543: inst = 32'h8c50000;
      37544: inst = 32'h24612800;
      37545: inst = 32'h10a0ffff;
      37546: inst = 32'hca0ffe1;
      37547: inst = 32'h24822800;
      37548: inst = 32'h10a00000;
      37549: inst = 32'hca00004;
      37550: inst = 32'h38632800;
      37551: inst = 32'h38842800;
      37552: inst = 32'h10a00000;
      37553: inst = 32'hca092b5;
      37554: inst = 32'h13e00001;
      37555: inst = 32'hfe0d96a;
      37556: inst = 32'h5be00000;
      37557: inst = 32'h8c50000;
      37558: inst = 32'h24612800;
      37559: inst = 32'h10a0ffff;
      37560: inst = 32'hca0ffe1;
      37561: inst = 32'h24822800;
      37562: inst = 32'h10a00000;
      37563: inst = 32'hca00004;
      37564: inst = 32'h38632800;
      37565: inst = 32'h38842800;
      37566: inst = 32'h10a00000;
      37567: inst = 32'hca092c3;
      37568: inst = 32'h13e00001;
      37569: inst = 32'hfe0d96a;
      37570: inst = 32'h5be00000;
      37571: inst = 32'h8c50000;
      37572: inst = 32'h24612800;
      37573: inst = 32'h10a0ffff;
      37574: inst = 32'hca0ffe1;
      37575: inst = 32'h24822800;
      37576: inst = 32'h10a00000;
      37577: inst = 32'hca00004;
      37578: inst = 32'h38632800;
      37579: inst = 32'h38842800;
      37580: inst = 32'h10a00000;
      37581: inst = 32'hca092d1;
      37582: inst = 32'h13e00001;
      37583: inst = 32'hfe0d96a;
      37584: inst = 32'h5be00000;
      37585: inst = 32'h8c50000;
      37586: inst = 32'h24612800;
      37587: inst = 32'h10a0ffff;
      37588: inst = 32'hca0ffe1;
      37589: inst = 32'h24822800;
      37590: inst = 32'h10a00000;
      37591: inst = 32'hca00004;
      37592: inst = 32'h38632800;
      37593: inst = 32'h38842800;
      37594: inst = 32'h10a00000;
      37595: inst = 32'hca092df;
      37596: inst = 32'h13e00001;
      37597: inst = 32'hfe0d96a;
      37598: inst = 32'h5be00000;
      37599: inst = 32'h8c50000;
      37600: inst = 32'h24612800;
      37601: inst = 32'h10a0ffff;
      37602: inst = 32'hca0ffe1;
      37603: inst = 32'h24822800;
      37604: inst = 32'h10a00000;
      37605: inst = 32'hca00004;
      37606: inst = 32'h38632800;
      37607: inst = 32'h38842800;
      37608: inst = 32'h10a00000;
      37609: inst = 32'hca092ed;
      37610: inst = 32'h13e00001;
      37611: inst = 32'hfe0d96a;
      37612: inst = 32'h5be00000;
      37613: inst = 32'h8c50000;
      37614: inst = 32'h24612800;
      37615: inst = 32'h10a0ffff;
      37616: inst = 32'hca0ffe1;
      37617: inst = 32'h24822800;
      37618: inst = 32'h10a00000;
      37619: inst = 32'hca00004;
      37620: inst = 32'h38632800;
      37621: inst = 32'h38842800;
      37622: inst = 32'h10a00000;
      37623: inst = 32'hca092fb;
      37624: inst = 32'h13e00001;
      37625: inst = 32'hfe0d96a;
      37626: inst = 32'h5be00000;
      37627: inst = 32'h8c50000;
      37628: inst = 32'h24612800;
      37629: inst = 32'h10a0ffff;
      37630: inst = 32'hca0ffe1;
      37631: inst = 32'h24822800;
      37632: inst = 32'h10a00000;
      37633: inst = 32'hca00004;
      37634: inst = 32'h38632800;
      37635: inst = 32'h38842800;
      37636: inst = 32'h10a00000;
      37637: inst = 32'hca09309;
      37638: inst = 32'h13e00001;
      37639: inst = 32'hfe0d96a;
      37640: inst = 32'h5be00000;
      37641: inst = 32'h8c50000;
      37642: inst = 32'h24612800;
      37643: inst = 32'h10a0ffff;
      37644: inst = 32'hca0ffe1;
      37645: inst = 32'h24822800;
      37646: inst = 32'h10a00000;
      37647: inst = 32'hca00004;
      37648: inst = 32'h38632800;
      37649: inst = 32'h38842800;
      37650: inst = 32'h10a00000;
      37651: inst = 32'hca09317;
      37652: inst = 32'h13e00001;
      37653: inst = 32'hfe0d96a;
      37654: inst = 32'h5be00000;
      37655: inst = 32'h8c50000;
      37656: inst = 32'h24612800;
      37657: inst = 32'h10a0ffff;
      37658: inst = 32'hca0ffe1;
      37659: inst = 32'h24822800;
      37660: inst = 32'h10a00000;
      37661: inst = 32'hca00004;
      37662: inst = 32'h38632800;
      37663: inst = 32'h38842800;
      37664: inst = 32'h10a00000;
      37665: inst = 32'hca09325;
      37666: inst = 32'h13e00001;
      37667: inst = 32'hfe0d96a;
      37668: inst = 32'h5be00000;
      37669: inst = 32'h8c50000;
      37670: inst = 32'h24612800;
      37671: inst = 32'h10a0ffff;
      37672: inst = 32'hca0ffe1;
      37673: inst = 32'h24822800;
      37674: inst = 32'h10a00000;
      37675: inst = 32'hca00004;
      37676: inst = 32'h38632800;
      37677: inst = 32'h38842800;
      37678: inst = 32'h10a00000;
      37679: inst = 32'hca09333;
      37680: inst = 32'h13e00001;
      37681: inst = 32'hfe0d96a;
      37682: inst = 32'h5be00000;
      37683: inst = 32'h8c50000;
      37684: inst = 32'h24612800;
      37685: inst = 32'h10a0ffff;
      37686: inst = 32'hca0ffe1;
      37687: inst = 32'h24822800;
      37688: inst = 32'h10a00000;
      37689: inst = 32'hca00004;
      37690: inst = 32'h38632800;
      37691: inst = 32'h38842800;
      37692: inst = 32'h10a00000;
      37693: inst = 32'hca09341;
      37694: inst = 32'h13e00001;
      37695: inst = 32'hfe0d96a;
      37696: inst = 32'h5be00000;
      37697: inst = 32'h8c50000;
      37698: inst = 32'h24612800;
      37699: inst = 32'h10a0ffff;
      37700: inst = 32'hca0ffe1;
      37701: inst = 32'h24822800;
      37702: inst = 32'h10a00000;
      37703: inst = 32'hca00004;
      37704: inst = 32'h38632800;
      37705: inst = 32'h38842800;
      37706: inst = 32'h10a00000;
      37707: inst = 32'hca0934f;
      37708: inst = 32'h13e00001;
      37709: inst = 32'hfe0d96a;
      37710: inst = 32'h5be00000;
      37711: inst = 32'h8c50000;
      37712: inst = 32'h24612800;
      37713: inst = 32'h10a0ffff;
      37714: inst = 32'hca0ffe1;
      37715: inst = 32'h24822800;
      37716: inst = 32'h10a00000;
      37717: inst = 32'hca00004;
      37718: inst = 32'h38632800;
      37719: inst = 32'h38842800;
      37720: inst = 32'h10a00000;
      37721: inst = 32'hca0935d;
      37722: inst = 32'h13e00001;
      37723: inst = 32'hfe0d96a;
      37724: inst = 32'h5be00000;
      37725: inst = 32'h8c50000;
      37726: inst = 32'h24612800;
      37727: inst = 32'h10a0ffff;
      37728: inst = 32'hca0ffe1;
      37729: inst = 32'h24822800;
      37730: inst = 32'h10a00000;
      37731: inst = 32'hca00004;
      37732: inst = 32'h38632800;
      37733: inst = 32'h38842800;
      37734: inst = 32'h10a00000;
      37735: inst = 32'hca0936b;
      37736: inst = 32'h13e00001;
      37737: inst = 32'hfe0d96a;
      37738: inst = 32'h5be00000;
      37739: inst = 32'h8c50000;
      37740: inst = 32'h24612800;
      37741: inst = 32'h10a0ffff;
      37742: inst = 32'hca0ffe1;
      37743: inst = 32'h24822800;
      37744: inst = 32'h10a00000;
      37745: inst = 32'hca00004;
      37746: inst = 32'h38632800;
      37747: inst = 32'h38842800;
      37748: inst = 32'h10a00000;
      37749: inst = 32'hca09379;
      37750: inst = 32'h13e00001;
      37751: inst = 32'hfe0d96a;
      37752: inst = 32'h5be00000;
      37753: inst = 32'h8c50000;
      37754: inst = 32'h24612800;
      37755: inst = 32'h10a0ffff;
      37756: inst = 32'hca0ffe1;
      37757: inst = 32'h24822800;
      37758: inst = 32'h10a00000;
      37759: inst = 32'hca00004;
      37760: inst = 32'h38632800;
      37761: inst = 32'h38842800;
      37762: inst = 32'h10a00000;
      37763: inst = 32'hca09387;
      37764: inst = 32'h13e00001;
      37765: inst = 32'hfe0d96a;
      37766: inst = 32'h5be00000;
      37767: inst = 32'h8c50000;
      37768: inst = 32'h24612800;
      37769: inst = 32'h10a0ffff;
      37770: inst = 32'hca0ffe1;
      37771: inst = 32'h24822800;
      37772: inst = 32'h10a00000;
      37773: inst = 32'hca00004;
      37774: inst = 32'h38632800;
      37775: inst = 32'h38842800;
      37776: inst = 32'h10a00000;
      37777: inst = 32'hca09395;
      37778: inst = 32'h13e00001;
      37779: inst = 32'hfe0d96a;
      37780: inst = 32'h5be00000;
      37781: inst = 32'h8c50000;
      37782: inst = 32'h24612800;
      37783: inst = 32'h10a0ffff;
      37784: inst = 32'hca0ffe1;
      37785: inst = 32'h24822800;
      37786: inst = 32'h10a00000;
      37787: inst = 32'hca00004;
      37788: inst = 32'h38632800;
      37789: inst = 32'h38842800;
      37790: inst = 32'h10a00000;
      37791: inst = 32'hca093a3;
      37792: inst = 32'h13e00001;
      37793: inst = 32'hfe0d96a;
      37794: inst = 32'h5be00000;
      37795: inst = 32'h8c50000;
      37796: inst = 32'h24612800;
      37797: inst = 32'h10a0ffff;
      37798: inst = 32'hca0ffe1;
      37799: inst = 32'h24822800;
      37800: inst = 32'h10a00000;
      37801: inst = 32'hca00004;
      37802: inst = 32'h38632800;
      37803: inst = 32'h38842800;
      37804: inst = 32'h10a00000;
      37805: inst = 32'hca093b1;
      37806: inst = 32'h13e00001;
      37807: inst = 32'hfe0d96a;
      37808: inst = 32'h5be00000;
      37809: inst = 32'h8c50000;
      37810: inst = 32'h24612800;
      37811: inst = 32'h10a0ffff;
      37812: inst = 32'hca0ffe1;
      37813: inst = 32'h24822800;
      37814: inst = 32'h10a00000;
      37815: inst = 32'hca00004;
      37816: inst = 32'h38632800;
      37817: inst = 32'h38842800;
      37818: inst = 32'h10a00000;
      37819: inst = 32'hca093bf;
      37820: inst = 32'h13e00001;
      37821: inst = 32'hfe0d96a;
      37822: inst = 32'h5be00000;
      37823: inst = 32'h8c50000;
      37824: inst = 32'h24612800;
      37825: inst = 32'h10a0ffff;
      37826: inst = 32'hca0ffe1;
      37827: inst = 32'h24822800;
      37828: inst = 32'h10a00000;
      37829: inst = 32'hca00004;
      37830: inst = 32'h38632800;
      37831: inst = 32'h38842800;
      37832: inst = 32'h10a00000;
      37833: inst = 32'hca093cd;
      37834: inst = 32'h13e00001;
      37835: inst = 32'hfe0d96a;
      37836: inst = 32'h5be00000;
      37837: inst = 32'h8c50000;
      37838: inst = 32'h24612800;
      37839: inst = 32'h10a0ffff;
      37840: inst = 32'hca0ffe1;
      37841: inst = 32'h24822800;
      37842: inst = 32'h10a00000;
      37843: inst = 32'hca00004;
      37844: inst = 32'h38632800;
      37845: inst = 32'h38842800;
      37846: inst = 32'h10a00000;
      37847: inst = 32'hca093db;
      37848: inst = 32'h13e00001;
      37849: inst = 32'hfe0d96a;
      37850: inst = 32'h5be00000;
      37851: inst = 32'h8c50000;
      37852: inst = 32'h24612800;
      37853: inst = 32'h10a0ffff;
      37854: inst = 32'hca0ffe1;
      37855: inst = 32'h24822800;
      37856: inst = 32'h10a00000;
      37857: inst = 32'hca00004;
      37858: inst = 32'h38632800;
      37859: inst = 32'h38842800;
      37860: inst = 32'h10a00000;
      37861: inst = 32'hca093e9;
      37862: inst = 32'h13e00001;
      37863: inst = 32'hfe0d96a;
      37864: inst = 32'h5be00000;
      37865: inst = 32'h8c50000;
      37866: inst = 32'h24612800;
      37867: inst = 32'h10a0ffff;
      37868: inst = 32'hca0ffe2;
      37869: inst = 32'h24822800;
      37870: inst = 32'h10a00000;
      37871: inst = 32'hca00004;
      37872: inst = 32'h38632800;
      37873: inst = 32'h38842800;
      37874: inst = 32'h10a00000;
      37875: inst = 32'hca093f7;
      37876: inst = 32'h13e00001;
      37877: inst = 32'hfe0d96a;
      37878: inst = 32'h5be00000;
      37879: inst = 32'h8c50000;
      37880: inst = 32'h24612800;
      37881: inst = 32'h10a0ffff;
      37882: inst = 32'hca0ffe2;
      37883: inst = 32'h24822800;
      37884: inst = 32'h10a00000;
      37885: inst = 32'hca00004;
      37886: inst = 32'h38632800;
      37887: inst = 32'h38842800;
      37888: inst = 32'h10a00000;
      37889: inst = 32'hca09405;
      37890: inst = 32'h13e00001;
      37891: inst = 32'hfe0d96a;
      37892: inst = 32'h5be00000;
      37893: inst = 32'h8c50000;
      37894: inst = 32'h24612800;
      37895: inst = 32'h10a0ffff;
      37896: inst = 32'hca0ffe2;
      37897: inst = 32'h24822800;
      37898: inst = 32'h10a00000;
      37899: inst = 32'hca00004;
      37900: inst = 32'h38632800;
      37901: inst = 32'h38842800;
      37902: inst = 32'h10a00000;
      37903: inst = 32'hca09413;
      37904: inst = 32'h13e00001;
      37905: inst = 32'hfe0d96a;
      37906: inst = 32'h5be00000;
      37907: inst = 32'h8c50000;
      37908: inst = 32'h24612800;
      37909: inst = 32'h10a0ffff;
      37910: inst = 32'hca0ffe2;
      37911: inst = 32'h24822800;
      37912: inst = 32'h10a00000;
      37913: inst = 32'hca00004;
      37914: inst = 32'h38632800;
      37915: inst = 32'h38842800;
      37916: inst = 32'h10a00000;
      37917: inst = 32'hca09421;
      37918: inst = 32'h13e00001;
      37919: inst = 32'hfe0d96a;
      37920: inst = 32'h5be00000;
      37921: inst = 32'h8c50000;
      37922: inst = 32'h24612800;
      37923: inst = 32'h10a0ffff;
      37924: inst = 32'hca0ffe2;
      37925: inst = 32'h24822800;
      37926: inst = 32'h10a00000;
      37927: inst = 32'hca00004;
      37928: inst = 32'h38632800;
      37929: inst = 32'h38842800;
      37930: inst = 32'h10a00000;
      37931: inst = 32'hca0942f;
      37932: inst = 32'h13e00001;
      37933: inst = 32'hfe0d96a;
      37934: inst = 32'h5be00000;
      37935: inst = 32'h8c50000;
      37936: inst = 32'h24612800;
      37937: inst = 32'h10a0ffff;
      37938: inst = 32'hca0ffe2;
      37939: inst = 32'h24822800;
      37940: inst = 32'h10a00000;
      37941: inst = 32'hca00004;
      37942: inst = 32'h38632800;
      37943: inst = 32'h38842800;
      37944: inst = 32'h10a00000;
      37945: inst = 32'hca0943d;
      37946: inst = 32'h13e00001;
      37947: inst = 32'hfe0d96a;
      37948: inst = 32'h5be00000;
      37949: inst = 32'h8c50000;
      37950: inst = 32'h24612800;
      37951: inst = 32'h10a0ffff;
      37952: inst = 32'hca0ffe2;
      37953: inst = 32'h24822800;
      37954: inst = 32'h10a00000;
      37955: inst = 32'hca00004;
      37956: inst = 32'h38632800;
      37957: inst = 32'h38842800;
      37958: inst = 32'h10a00000;
      37959: inst = 32'hca0944b;
      37960: inst = 32'h13e00001;
      37961: inst = 32'hfe0d96a;
      37962: inst = 32'h5be00000;
      37963: inst = 32'h8c50000;
      37964: inst = 32'h24612800;
      37965: inst = 32'h10a0ffff;
      37966: inst = 32'hca0ffe2;
      37967: inst = 32'h24822800;
      37968: inst = 32'h10a00000;
      37969: inst = 32'hca00004;
      37970: inst = 32'h38632800;
      37971: inst = 32'h38842800;
      37972: inst = 32'h10a00000;
      37973: inst = 32'hca09459;
      37974: inst = 32'h13e00001;
      37975: inst = 32'hfe0d96a;
      37976: inst = 32'h5be00000;
      37977: inst = 32'h8c50000;
      37978: inst = 32'h24612800;
      37979: inst = 32'h10a0ffff;
      37980: inst = 32'hca0ffe2;
      37981: inst = 32'h24822800;
      37982: inst = 32'h10a00000;
      37983: inst = 32'hca00004;
      37984: inst = 32'h38632800;
      37985: inst = 32'h38842800;
      37986: inst = 32'h10a00000;
      37987: inst = 32'hca09467;
      37988: inst = 32'h13e00001;
      37989: inst = 32'hfe0d96a;
      37990: inst = 32'h5be00000;
      37991: inst = 32'h8c50000;
      37992: inst = 32'h24612800;
      37993: inst = 32'h10a0ffff;
      37994: inst = 32'hca0ffe2;
      37995: inst = 32'h24822800;
      37996: inst = 32'h10a00000;
      37997: inst = 32'hca00004;
      37998: inst = 32'h38632800;
      37999: inst = 32'h38842800;
      38000: inst = 32'h10a00000;
      38001: inst = 32'hca09475;
      38002: inst = 32'h13e00001;
      38003: inst = 32'hfe0d96a;
      38004: inst = 32'h5be00000;
      38005: inst = 32'h8c50000;
      38006: inst = 32'h24612800;
      38007: inst = 32'h10a0ffff;
      38008: inst = 32'hca0ffe2;
      38009: inst = 32'h24822800;
      38010: inst = 32'h10a00000;
      38011: inst = 32'hca00004;
      38012: inst = 32'h38632800;
      38013: inst = 32'h38842800;
      38014: inst = 32'h10a00000;
      38015: inst = 32'hca09483;
      38016: inst = 32'h13e00001;
      38017: inst = 32'hfe0d96a;
      38018: inst = 32'h5be00000;
      38019: inst = 32'h8c50000;
      38020: inst = 32'h24612800;
      38021: inst = 32'h10a0ffff;
      38022: inst = 32'hca0ffe2;
      38023: inst = 32'h24822800;
      38024: inst = 32'h10a00000;
      38025: inst = 32'hca00004;
      38026: inst = 32'h38632800;
      38027: inst = 32'h38842800;
      38028: inst = 32'h10a00000;
      38029: inst = 32'hca09491;
      38030: inst = 32'h13e00001;
      38031: inst = 32'hfe0d96a;
      38032: inst = 32'h5be00000;
      38033: inst = 32'h8c50000;
      38034: inst = 32'h24612800;
      38035: inst = 32'h10a0ffff;
      38036: inst = 32'hca0ffe2;
      38037: inst = 32'h24822800;
      38038: inst = 32'h10a00000;
      38039: inst = 32'hca00004;
      38040: inst = 32'h38632800;
      38041: inst = 32'h38842800;
      38042: inst = 32'h10a00000;
      38043: inst = 32'hca0949f;
      38044: inst = 32'h13e00001;
      38045: inst = 32'hfe0d96a;
      38046: inst = 32'h5be00000;
      38047: inst = 32'h8c50000;
      38048: inst = 32'h24612800;
      38049: inst = 32'h10a0ffff;
      38050: inst = 32'hca0ffe2;
      38051: inst = 32'h24822800;
      38052: inst = 32'h10a00000;
      38053: inst = 32'hca00004;
      38054: inst = 32'h38632800;
      38055: inst = 32'h38842800;
      38056: inst = 32'h10a00000;
      38057: inst = 32'hca094ad;
      38058: inst = 32'h13e00001;
      38059: inst = 32'hfe0d96a;
      38060: inst = 32'h5be00000;
      38061: inst = 32'h8c50000;
      38062: inst = 32'h24612800;
      38063: inst = 32'h10a0ffff;
      38064: inst = 32'hca0ffe2;
      38065: inst = 32'h24822800;
      38066: inst = 32'h10a00000;
      38067: inst = 32'hca00004;
      38068: inst = 32'h38632800;
      38069: inst = 32'h38842800;
      38070: inst = 32'h10a00000;
      38071: inst = 32'hca094bb;
      38072: inst = 32'h13e00001;
      38073: inst = 32'hfe0d96a;
      38074: inst = 32'h5be00000;
      38075: inst = 32'h8c50000;
      38076: inst = 32'h24612800;
      38077: inst = 32'h10a0ffff;
      38078: inst = 32'hca0ffe2;
      38079: inst = 32'h24822800;
      38080: inst = 32'h10a00000;
      38081: inst = 32'hca00004;
      38082: inst = 32'h38632800;
      38083: inst = 32'h38842800;
      38084: inst = 32'h10a00000;
      38085: inst = 32'hca094c9;
      38086: inst = 32'h13e00001;
      38087: inst = 32'hfe0d96a;
      38088: inst = 32'h5be00000;
      38089: inst = 32'h8c50000;
      38090: inst = 32'h24612800;
      38091: inst = 32'h10a0ffff;
      38092: inst = 32'hca0ffe2;
      38093: inst = 32'h24822800;
      38094: inst = 32'h10a00000;
      38095: inst = 32'hca00004;
      38096: inst = 32'h38632800;
      38097: inst = 32'h38842800;
      38098: inst = 32'h10a00000;
      38099: inst = 32'hca094d7;
      38100: inst = 32'h13e00001;
      38101: inst = 32'hfe0d96a;
      38102: inst = 32'h5be00000;
      38103: inst = 32'h8c50000;
      38104: inst = 32'h24612800;
      38105: inst = 32'h10a0ffff;
      38106: inst = 32'hca0ffe2;
      38107: inst = 32'h24822800;
      38108: inst = 32'h10a00000;
      38109: inst = 32'hca00004;
      38110: inst = 32'h38632800;
      38111: inst = 32'h38842800;
      38112: inst = 32'h10a00000;
      38113: inst = 32'hca094e5;
      38114: inst = 32'h13e00001;
      38115: inst = 32'hfe0d96a;
      38116: inst = 32'h5be00000;
      38117: inst = 32'h8c50000;
      38118: inst = 32'h24612800;
      38119: inst = 32'h10a0ffff;
      38120: inst = 32'hca0ffe2;
      38121: inst = 32'h24822800;
      38122: inst = 32'h10a00000;
      38123: inst = 32'hca00004;
      38124: inst = 32'h38632800;
      38125: inst = 32'h38842800;
      38126: inst = 32'h10a00000;
      38127: inst = 32'hca094f3;
      38128: inst = 32'h13e00001;
      38129: inst = 32'hfe0d96a;
      38130: inst = 32'h5be00000;
      38131: inst = 32'h8c50000;
      38132: inst = 32'h24612800;
      38133: inst = 32'h10a0ffff;
      38134: inst = 32'hca0ffe2;
      38135: inst = 32'h24822800;
      38136: inst = 32'h10a00000;
      38137: inst = 32'hca00004;
      38138: inst = 32'h38632800;
      38139: inst = 32'h38842800;
      38140: inst = 32'h10a00000;
      38141: inst = 32'hca09501;
      38142: inst = 32'h13e00001;
      38143: inst = 32'hfe0d96a;
      38144: inst = 32'h5be00000;
      38145: inst = 32'h8c50000;
      38146: inst = 32'h24612800;
      38147: inst = 32'h10a0ffff;
      38148: inst = 32'hca0ffe2;
      38149: inst = 32'h24822800;
      38150: inst = 32'h10a00000;
      38151: inst = 32'hca00004;
      38152: inst = 32'h38632800;
      38153: inst = 32'h38842800;
      38154: inst = 32'h10a00000;
      38155: inst = 32'hca0950f;
      38156: inst = 32'h13e00001;
      38157: inst = 32'hfe0d96a;
      38158: inst = 32'h5be00000;
      38159: inst = 32'h8c50000;
      38160: inst = 32'h24612800;
      38161: inst = 32'h10a0ffff;
      38162: inst = 32'hca0ffe2;
      38163: inst = 32'h24822800;
      38164: inst = 32'h10a00000;
      38165: inst = 32'hca00004;
      38166: inst = 32'h38632800;
      38167: inst = 32'h38842800;
      38168: inst = 32'h10a00000;
      38169: inst = 32'hca0951d;
      38170: inst = 32'h13e00001;
      38171: inst = 32'hfe0d96a;
      38172: inst = 32'h5be00000;
      38173: inst = 32'h8c50000;
      38174: inst = 32'h24612800;
      38175: inst = 32'h10a0ffff;
      38176: inst = 32'hca0ffe2;
      38177: inst = 32'h24822800;
      38178: inst = 32'h10a00000;
      38179: inst = 32'hca00004;
      38180: inst = 32'h38632800;
      38181: inst = 32'h38842800;
      38182: inst = 32'h10a00000;
      38183: inst = 32'hca0952b;
      38184: inst = 32'h13e00001;
      38185: inst = 32'hfe0d96a;
      38186: inst = 32'h5be00000;
      38187: inst = 32'h8c50000;
      38188: inst = 32'h24612800;
      38189: inst = 32'h10a0ffff;
      38190: inst = 32'hca0ffe2;
      38191: inst = 32'h24822800;
      38192: inst = 32'h10a00000;
      38193: inst = 32'hca00004;
      38194: inst = 32'h38632800;
      38195: inst = 32'h38842800;
      38196: inst = 32'h10a00000;
      38197: inst = 32'hca09539;
      38198: inst = 32'h13e00001;
      38199: inst = 32'hfe0d96a;
      38200: inst = 32'h5be00000;
      38201: inst = 32'h8c50000;
      38202: inst = 32'h24612800;
      38203: inst = 32'h10a0ffff;
      38204: inst = 32'hca0ffe2;
      38205: inst = 32'h24822800;
      38206: inst = 32'h10a00000;
      38207: inst = 32'hca00004;
      38208: inst = 32'h38632800;
      38209: inst = 32'h38842800;
      38210: inst = 32'h10a00000;
      38211: inst = 32'hca09547;
      38212: inst = 32'h13e00001;
      38213: inst = 32'hfe0d96a;
      38214: inst = 32'h5be00000;
      38215: inst = 32'h8c50000;
      38216: inst = 32'h24612800;
      38217: inst = 32'h10a0ffff;
      38218: inst = 32'hca0ffe2;
      38219: inst = 32'h24822800;
      38220: inst = 32'h10a00000;
      38221: inst = 32'hca00004;
      38222: inst = 32'h38632800;
      38223: inst = 32'h38842800;
      38224: inst = 32'h10a00000;
      38225: inst = 32'hca09555;
      38226: inst = 32'h13e00001;
      38227: inst = 32'hfe0d96a;
      38228: inst = 32'h5be00000;
      38229: inst = 32'h8c50000;
      38230: inst = 32'h24612800;
      38231: inst = 32'h10a0ffff;
      38232: inst = 32'hca0ffe2;
      38233: inst = 32'h24822800;
      38234: inst = 32'h10a00000;
      38235: inst = 32'hca00004;
      38236: inst = 32'h38632800;
      38237: inst = 32'h38842800;
      38238: inst = 32'h10a00000;
      38239: inst = 32'hca09563;
      38240: inst = 32'h13e00001;
      38241: inst = 32'hfe0d96a;
      38242: inst = 32'h5be00000;
      38243: inst = 32'h8c50000;
      38244: inst = 32'h24612800;
      38245: inst = 32'h10a0ffff;
      38246: inst = 32'hca0ffe2;
      38247: inst = 32'h24822800;
      38248: inst = 32'h10a00000;
      38249: inst = 32'hca00004;
      38250: inst = 32'h38632800;
      38251: inst = 32'h38842800;
      38252: inst = 32'h10a00000;
      38253: inst = 32'hca09571;
      38254: inst = 32'h13e00001;
      38255: inst = 32'hfe0d96a;
      38256: inst = 32'h5be00000;
      38257: inst = 32'h8c50000;
      38258: inst = 32'h24612800;
      38259: inst = 32'h10a0ffff;
      38260: inst = 32'hca0ffe2;
      38261: inst = 32'h24822800;
      38262: inst = 32'h10a00000;
      38263: inst = 32'hca00004;
      38264: inst = 32'h38632800;
      38265: inst = 32'h38842800;
      38266: inst = 32'h10a00000;
      38267: inst = 32'hca0957f;
      38268: inst = 32'h13e00001;
      38269: inst = 32'hfe0d96a;
      38270: inst = 32'h5be00000;
      38271: inst = 32'h8c50000;
      38272: inst = 32'h24612800;
      38273: inst = 32'h10a0ffff;
      38274: inst = 32'hca0ffe2;
      38275: inst = 32'h24822800;
      38276: inst = 32'h10a00000;
      38277: inst = 32'hca00004;
      38278: inst = 32'h38632800;
      38279: inst = 32'h38842800;
      38280: inst = 32'h10a00000;
      38281: inst = 32'hca0958d;
      38282: inst = 32'h13e00001;
      38283: inst = 32'hfe0d96a;
      38284: inst = 32'h5be00000;
      38285: inst = 32'h8c50000;
      38286: inst = 32'h24612800;
      38287: inst = 32'h10a0ffff;
      38288: inst = 32'hca0ffe2;
      38289: inst = 32'h24822800;
      38290: inst = 32'h10a00000;
      38291: inst = 32'hca00004;
      38292: inst = 32'h38632800;
      38293: inst = 32'h38842800;
      38294: inst = 32'h10a00000;
      38295: inst = 32'hca0959b;
      38296: inst = 32'h13e00001;
      38297: inst = 32'hfe0d96a;
      38298: inst = 32'h5be00000;
      38299: inst = 32'h8c50000;
      38300: inst = 32'h24612800;
      38301: inst = 32'h10a0ffff;
      38302: inst = 32'hca0ffe2;
      38303: inst = 32'h24822800;
      38304: inst = 32'h10a00000;
      38305: inst = 32'hca00004;
      38306: inst = 32'h38632800;
      38307: inst = 32'h38842800;
      38308: inst = 32'h10a00000;
      38309: inst = 32'hca095a9;
      38310: inst = 32'h13e00001;
      38311: inst = 32'hfe0d96a;
      38312: inst = 32'h5be00000;
      38313: inst = 32'h8c50000;
      38314: inst = 32'h24612800;
      38315: inst = 32'h10a0ffff;
      38316: inst = 32'hca0ffe2;
      38317: inst = 32'h24822800;
      38318: inst = 32'h10a00000;
      38319: inst = 32'hca00004;
      38320: inst = 32'h38632800;
      38321: inst = 32'h38842800;
      38322: inst = 32'h10a00000;
      38323: inst = 32'hca095b7;
      38324: inst = 32'h13e00001;
      38325: inst = 32'hfe0d96a;
      38326: inst = 32'h5be00000;
      38327: inst = 32'h8c50000;
      38328: inst = 32'h24612800;
      38329: inst = 32'h10a0ffff;
      38330: inst = 32'hca0ffe2;
      38331: inst = 32'h24822800;
      38332: inst = 32'h10a00000;
      38333: inst = 32'hca00004;
      38334: inst = 32'h38632800;
      38335: inst = 32'h38842800;
      38336: inst = 32'h10a00000;
      38337: inst = 32'hca095c5;
      38338: inst = 32'h13e00001;
      38339: inst = 32'hfe0d96a;
      38340: inst = 32'h5be00000;
      38341: inst = 32'h8c50000;
      38342: inst = 32'h24612800;
      38343: inst = 32'h10a0ffff;
      38344: inst = 32'hca0ffe2;
      38345: inst = 32'h24822800;
      38346: inst = 32'h10a00000;
      38347: inst = 32'hca00004;
      38348: inst = 32'h38632800;
      38349: inst = 32'h38842800;
      38350: inst = 32'h10a00000;
      38351: inst = 32'hca095d3;
      38352: inst = 32'h13e00001;
      38353: inst = 32'hfe0d96a;
      38354: inst = 32'h5be00000;
      38355: inst = 32'h8c50000;
      38356: inst = 32'h24612800;
      38357: inst = 32'h10a0ffff;
      38358: inst = 32'hca0ffe2;
      38359: inst = 32'h24822800;
      38360: inst = 32'h10a00000;
      38361: inst = 32'hca00004;
      38362: inst = 32'h38632800;
      38363: inst = 32'h38842800;
      38364: inst = 32'h10a00000;
      38365: inst = 32'hca095e1;
      38366: inst = 32'h13e00001;
      38367: inst = 32'hfe0d96a;
      38368: inst = 32'h5be00000;
      38369: inst = 32'h8c50000;
      38370: inst = 32'h24612800;
      38371: inst = 32'h10a0ffff;
      38372: inst = 32'hca0ffe2;
      38373: inst = 32'h24822800;
      38374: inst = 32'h10a00000;
      38375: inst = 32'hca00004;
      38376: inst = 32'h38632800;
      38377: inst = 32'h38842800;
      38378: inst = 32'h10a00000;
      38379: inst = 32'hca095ef;
      38380: inst = 32'h13e00001;
      38381: inst = 32'hfe0d96a;
      38382: inst = 32'h5be00000;
      38383: inst = 32'h8c50000;
      38384: inst = 32'h24612800;
      38385: inst = 32'h10a0ffff;
      38386: inst = 32'hca0ffe2;
      38387: inst = 32'h24822800;
      38388: inst = 32'h10a00000;
      38389: inst = 32'hca00004;
      38390: inst = 32'h38632800;
      38391: inst = 32'h38842800;
      38392: inst = 32'h10a00000;
      38393: inst = 32'hca095fd;
      38394: inst = 32'h13e00001;
      38395: inst = 32'hfe0d96a;
      38396: inst = 32'h5be00000;
      38397: inst = 32'h8c50000;
      38398: inst = 32'h24612800;
      38399: inst = 32'h10a0ffff;
      38400: inst = 32'hca0ffe2;
      38401: inst = 32'h24822800;
      38402: inst = 32'h10a00000;
      38403: inst = 32'hca00004;
      38404: inst = 32'h38632800;
      38405: inst = 32'h38842800;
      38406: inst = 32'h10a00000;
      38407: inst = 32'hca0960b;
      38408: inst = 32'h13e00001;
      38409: inst = 32'hfe0d96a;
      38410: inst = 32'h5be00000;
      38411: inst = 32'h8c50000;
      38412: inst = 32'h24612800;
      38413: inst = 32'h10a0ffff;
      38414: inst = 32'hca0ffe2;
      38415: inst = 32'h24822800;
      38416: inst = 32'h10a00000;
      38417: inst = 32'hca00004;
      38418: inst = 32'h38632800;
      38419: inst = 32'h38842800;
      38420: inst = 32'h10a00000;
      38421: inst = 32'hca09619;
      38422: inst = 32'h13e00001;
      38423: inst = 32'hfe0d96a;
      38424: inst = 32'h5be00000;
      38425: inst = 32'h8c50000;
      38426: inst = 32'h24612800;
      38427: inst = 32'h10a0ffff;
      38428: inst = 32'hca0ffe2;
      38429: inst = 32'h24822800;
      38430: inst = 32'h10a00000;
      38431: inst = 32'hca00004;
      38432: inst = 32'h38632800;
      38433: inst = 32'h38842800;
      38434: inst = 32'h10a00000;
      38435: inst = 32'hca09627;
      38436: inst = 32'h13e00001;
      38437: inst = 32'hfe0d96a;
      38438: inst = 32'h5be00000;
      38439: inst = 32'h8c50000;
      38440: inst = 32'h24612800;
      38441: inst = 32'h10a0ffff;
      38442: inst = 32'hca0ffe2;
      38443: inst = 32'h24822800;
      38444: inst = 32'h10a00000;
      38445: inst = 32'hca00004;
      38446: inst = 32'h38632800;
      38447: inst = 32'h38842800;
      38448: inst = 32'h10a00000;
      38449: inst = 32'hca09635;
      38450: inst = 32'h13e00001;
      38451: inst = 32'hfe0d96a;
      38452: inst = 32'h5be00000;
      38453: inst = 32'h8c50000;
      38454: inst = 32'h24612800;
      38455: inst = 32'h10a0ffff;
      38456: inst = 32'hca0ffe2;
      38457: inst = 32'h24822800;
      38458: inst = 32'h10a00000;
      38459: inst = 32'hca00004;
      38460: inst = 32'h38632800;
      38461: inst = 32'h38842800;
      38462: inst = 32'h10a00000;
      38463: inst = 32'hca09643;
      38464: inst = 32'h13e00001;
      38465: inst = 32'hfe0d96a;
      38466: inst = 32'h5be00000;
      38467: inst = 32'h8c50000;
      38468: inst = 32'h24612800;
      38469: inst = 32'h10a0ffff;
      38470: inst = 32'hca0ffe2;
      38471: inst = 32'h24822800;
      38472: inst = 32'h10a00000;
      38473: inst = 32'hca00004;
      38474: inst = 32'h38632800;
      38475: inst = 32'h38842800;
      38476: inst = 32'h10a00000;
      38477: inst = 32'hca09651;
      38478: inst = 32'h13e00001;
      38479: inst = 32'hfe0d96a;
      38480: inst = 32'h5be00000;
      38481: inst = 32'h8c50000;
      38482: inst = 32'h24612800;
      38483: inst = 32'h10a0ffff;
      38484: inst = 32'hca0ffe2;
      38485: inst = 32'h24822800;
      38486: inst = 32'h10a00000;
      38487: inst = 32'hca00004;
      38488: inst = 32'h38632800;
      38489: inst = 32'h38842800;
      38490: inst = 32'h10a00000;
      38491: inst = 32'hca0965f;
      38492: inst = 32'h13e00001;
      38493: inst = 32'hfe0d96a;
      38494: inst = 32'h5be00000;
      38495: inst = 32'h8c50000;
      38496: inst = 32'h24612800;
      38497: inst = 32'h10a0ffff;
      38498: inst = 32'hca0ffe2;
      38499: inst = 32'h24822800;
      38500: inst = 32'h10a00000;
      38501: inst = 32'hca00004;
      38502: inst = 32'h38632800;
      38503: inst = 32'h38842800;
      38504: inst = 32'h10a00000;
      38505: inst = 32'hca0966d;
      38506: inst = 32'h13e00001;
      38507: inst = 32'hfe0d96a;
      38508: inst = 32'h5be00000;
      38509: inst = 32'h8c50000;
      38510: inst = 32'h24612800;
      38511: inst = 32'h10a0ffff;
      38512: inst = 32'hca0ffe2;
      38513: inst = 32'h24822800;
      38514: inst = 32'h10a00000;
      38515: inst = 32'hca00004;
      38516: inst = 32'h38632800;
      38517: inst = 32'h38842800;
      38518: inst = 32'h10a00000;
      38519: inst = 32'hca0967b;
      38520: inst = 32'h13e00001;
      38521: inst = 32'hfe0d96a;
      38522: inst = 32'h5be00000;
      38523: inst = 32'h8c50000;
      38524: inst = 32'h24612800;
      38525: inst = 32'h10a0ffff;
      38526: inst = 32'hca0ffe2;
      38527: inst = 32'h24822800;
      38528: inst = 32'h10a00000;
      38529: inst = 32'hca00004;
      38530: inst = 32'h38632800;
      38531: inst = 32'h38842800;
      38532: inst = 32'h10a00000;
      38533: inst = 32'hca09689;
      38534: inst = 32'h13e00001;
      38535: inst = 32'hfe0d96a;
      38536: inst = 32'h5be00000;
      38537: inst = 32'h8c50000;
      38538: inst = 32'h24612800;
      38539: inst = 32'h10a0ffff;
      38540: inst = 32'hca0ffe2;
      38541: inst = 32'h24822800;
      38542: inst = 32'h10a00000;
      38543: inst = 32'hca00004;
      38544: inst = 32'h38632800;
      38545: inst = 32'h38842800;
      38546: inst = 32'h10a00000;
      38547: inst = 32'hca09697;
      38548: inst = 32'h13e00001;
      38549: inst = 32'hfe0d96a;
      38550: inst = 32'h5be00000;
      38551: inst = 32'h8c50000;
      38552: inst = 32'h24612800;
      38553: inst = 32'h10a0ffff;
      38554: inst = 32'hca0ffe2;
      38555: inst = 32'h24822800;
      38556: inst = 32'h10a00000;
      38557: inst = 32'hca00004;
      38558: inst = 32'h38632800;
      38559: inst = 32'h38842800;
      38560: inst = 32'h10a00000;
      38561: inst = 32'hca096a5;
      38562: inst = 32'h13e00001;
      38563: inst = 32'hfe0d96a;
      38564: inst = 32'h5be00000;
      38565: inst = 32'h8c50000;
      38566: inst = 32'h24612800;
      38567: inst = 32'h10a0ffff;
      38568: inst = 32'hca0ffe2;
      38569: inst = 32'h24822800;
      38570: inst = 32'h10a00000;
      38571: inst = 32'hca00004;
      38572: inst = 32'h38632800;
      38573: inst = 32'h38842800;
      38574: inst = 32'h10a00000;
      38575: inst = 32'hca096b3;
      38576: inst = 32'h13e00001;
      38577: inst = 32'hfe0d96a;
      38578: inst = 32'h5be00000;
      38579: inst = 32'h8c50000;
      38580: inst = 32'h24612800;
      38581: inst = 32'h10a0ffff;
      38582: inst = 32'hca0ffe2;
      38583: inst = 32'h24822800;
      38584: inst = 32'h10a00000;
      38585: inst = 32'hca00004;
      38586: inst = 32'h38632800;
      38587: inst = 32'h38842800;
      38588: inst = 32'h10a00000;
      38589: inst = 32'hca096c1;
      38590: inst = 32'h13e00001;
      38591: inst = 32'hfe0d96a;
      38592: inst = 32'h5be00000;
      38593: inst = 32'h8c50000;
      38594: inst = 32'h24612800;
      38595: inst = 32'h10a0ffff;
      38596: inst = 32'hca0ffe2;
      38597: inst = 32'h24822800;
      38598: inst = 32'h10a00000;
      38599: inst = 32'hca00004;
      38600: inst = 32'h38632800;
      38601: inst = 32'h38842800;
      38602: inst = 32'h10a00000;
      38603: inst = 32'hca096cf;
      38604: inst = 32'h13e00001;
      38605: inst = 32'hfe0d96a;
      38606: inst = 32'h5be00000;
      38607: inst = 32'h8c50000;
      38608: inst = 32'h24612800;
      38609: inst = 32'h10a0ffff;
      38610: inst = 32'hca0ffe2;
      38611: inst = 32'h24822800;
      38612: inst = 32'h10a00000;
      38613: inst = 32'hca00004;
      38614: inst = 32'h38632800;
      38615: inst = 32'h38842800;
      38616: inst = 32'h10a00000;
      38617: inst = 32'hca096dd;
      38618: inst = 32'h13e00001;
      38619: inst = 32'hfe0d96a;
      38620: inst = 32'h5be00000;
      38621: inst = 32'h8c50000;
      38622: inst = 32'h24612800;
      38623: inst = 32'h10a0ffff;
      38624: inst = 32'hca0ffe2;
      38625: inst = 32'h24822800;
      38626: inst = 32'h10a00000;
      38627: inst = 32'hca00004;
      38628: inst = 32'h38632800;
      38629: inst = 32'h38842800;
      38630: inst = 32'h10a00000;
      38631: inst = 32'hca096eb;
      38632: inst = 32'h13e00001;
      38633: inst = 32'hfe0d96a;
      38634: inst = 32'h5be00000;
      38635: inst = 32'h8c50000;
      38636: inst = 32'h24612800;
      38637: inst = 32'h10a0ffff;
      38638: inst = 32'hca0ffe2;
      38639: inst = 32'h24822800;
      38640: inst = 32'h10a00000;
      38641: inst = 32'hca00004;
      38642: inst = 32'h38632800;
      38643: inst = 32'h38842800;
      38644: inst = 32'h10a00000;
      38645: inst = 32'hca096f9;
      38646: inst = 32'h13e00001;
      38647: inst = 32'hfe0d96a;
      38648: inst = 32'h5be00000;
      38649: inst = 32'h8c50000;
      38650: inst = 32'h24612800;
      38651: inst = 32'h10a0ffff;
      38652: inst = 32'hca0ffe2;
      38653: inst = 32'h24822800;
      38654: inst = 32'h10a00000;
      38655: inst = 32'hca00004;
      38656: inst = 32'h38632800;
      38657: inst = 32'h38842800;
      38658: inst = 32'h10a00000;
      38659: inst = 32'hca09707;
      38660: inst = 32'h13e00001;
      38661: inst = 32'hfe0d96a;
      38662: inst = 32'h5be00000;
      38663: inst = 32'h8c50000;
      38664: inst = 32'h24612800;
      38665: inst = 32'h10a0ffff;
      38666: inst = 32'hca0ffe2;
      38667: inst = 32'h24822800;
      38668: inst = 32'h10a00000;
      38669: inst = 32'hca00004;
      38670: inst = 32'h38632800;
      38671: inst = 32'h38842800;
      38672: inst = 32'h10a00000;
      38673: inst = 32'hca09715;
      38674: inst = 32'h13e00001;
      38675: inst = 32'hfe0d96a;
      38676: inst = 32'h5be00000;
      38677: inst = 32'h8c50000;
      38678: inst = 32'h24612800;
      38679: inst = 32'h10a0ffff;
      38680: inst = 32'hca0ffe2;
      38681: inst = 32'h24822800;
      38682: inst = 32'h10a00000;
      38683: inst = 32'hca00004;
      38684: inst = 32'h38632800;
      38685: inst = 32'h38842800;
      38686: inst = 32'h10a00000;
      38687: inst = 32'hca09723;
      38688: inst = 32'h13e00001;
      38689: inst = 32'hfe0d96a;
      38690: inst = 32'h5be00000;
      38691: inst = 32'h8c50000;
      38692: inst = 32'h24612800;
      38693: inst = 32'h10a0ffff;
      38694: inst = 32'hca0ffe2;
      38695: inst = 32'h24822800;
      38696: inst = 32'h10a00000;
      38697: inst = 32'hca00004;
      38698: inst = 32'h38632800;
      38699: inst = 32'h38842800;
      38700: inst = 32'h10a00000;
      38701: inst = 32'hca09731;
      38702: inst = 32'h13e00001;
      38703: inst = 32'hfe0d96a;
      38704: inst = 32'h5be00000;
      38705: inst = 32'h8c50000;
      38706: inst = 32'h24612800;
      38707: inst = 32'h10a0ffff;
      38708: inst = 32'hca0ffe2;
      38709: inst = 32'h24822800;
      38710: inst = 32'h10a00000;
      38711: inst = 32'hca00004;
      38712: inst = 32'h38632800;
      38713: inst = 32'h38842800;
      38714: inst = 32'h10a00000;
      38715: inst = 32'hca0973f;
      38716: inst = 32'h13e00001;
      38717: inst = 32'hfe0d96a;
      38718: inst = 32'h5be00000;
      38719: inst = 32'h8c50000;
      38720: inst = 32'h24612800;
      38721: inst = 32'h10a0ffff;
      38722: inst = 32'hca0ffe2;
      38723: inst = 32'h24822800;
      38724: inst = 32'h10a00000;
      38725: inst = 32'hca00004;
      38726: inst = 32'h38632800;
      38727: inst = 32'h38842800;
      38728: inst = 32'h10a00000;
      38729: inst = 32'hca0974d;
      38730: inst = 32'h13e00001;
      38731: inst = 32'hfe0d96a;
      38732: inst = 32'h5be00000;
      38733: inst = 32'h8c50000;
      38734: inst = 32'h24612800;
      38735: inst = 32'h10a0ffff;
      38736: inst = 32'hca0ffe2;
      38737: inst = 32'h24822800;
      38738: inst = 32'h10a00000;
      38739: inst = 32'hca00004;
      38740: inst = 32'h38632800;
      38741: inst = 32'h38842800;
      38742: inst = 32'h10a00000;
      38743: inst = 32'hca0975b;
      38744: inst = 32'h13e00001;
      38745: inst = 32'hfe0d96a;
      38746: inst = 32'h5be00000;
      38747: inst = 32'h8c50000;
      38748: inst = 32'h24612800;
      38749: inst = 32'h10a0ffff;
      38750: inst = 32'hca0ffe2;
      38751: inst = 32'h24822800;
      38752: inst = 32'h10a00000;
      38753: inst = 32'hca00004;
      38754: inst = 32'h38632800;
      38755: inst = 32'h38842800;
      38756: inst = 32'h10a00000;
      38757: inst = 32'hca09769;
      38758: inst = 32'h13e00001;
      38759: inst = 32'hfe0d96a;
      38760: inst = 32'h5be00000;
      38761: inst = 32'h8c50000;
      38762: inst = 32'h24612800;
      38763: inst = 32'h10a0ffff;
      38764: inst = 32'hca0ffe2;
      38765: inst = 32'h24822800;
      38766: inst = 32'h10a00000;
      38767: inst = 32'hca00004;
      38768: inst = 32'h38632800;
      38769: inst = 32'h38842800;
      38770: inst = 32'h10a00000;
      38771: inst = 32'hca09777;
      38772: inst = 32'h13e00001;
      38773: inst = 32'hfe0d96a;
      38774: inst = 32'h5be00000;
      38775: inst = 32'h8c50000;
      38776: inst = 32'h24612800;
      38777: inst = 32'h10a0ffff;
      38778: inst = 32'hca0ffe2;
      38779: inst = 32'h24822800;
      38780: inst = 32'h10a00000;
      38781: inst = 32'hca00004;
      38782: inst = 32'h38632800;
      38783: inst = 32'h38842800;
      38784: inst = 32'h10a00000;
      38785: inst = 32'hca09785;
      38786: inst = 32'h13e00001;
      38787: inst = 32'hfe0d96a;
      38788: inst = 32'h5be00000;
      38789: inst = 32'h8c50000;
      38790: inst = 32'h24612800;
      38791: inst = 32'h10a0ffff;
      38792: inst = 32'hca0ffe2;
      38793: inst = 32'h24822800;
      38794: inst = 32'h10a00000;
      38795: inst = 32'hca00004;
      38796: inst = 32'h38632800;
      38797: inst = 32'h38842800;
      38798: inst = 32'h10a00000;
      38799: inst = 32'hca09793;
      38800: inst = 32'h13e00001;
      38801: inst = 32'hfe0d96a;
      38802: inst = 32'h5be00000;
      38803: inst = 32'h8c50000;
      38804: inst = 32'h24612800;
      38805: inst = 32'h10a0ffff;
      38806: inst = 32'hca0ffe2;
      38807: inst = 32'h24822800;
      38808: inst = 32'h10a00000;
      38809: inst = 32'hca00004;
      38810: inst = 32'h38632800;
      38811: inst = 32'h38842800;
      38812: inst = 32'h10a00000;
      38813: inst = 32'hca097a1;
      38814: inst = 32'h13e00001;
      38815: inst = 32'hfe0d96a;
      38816: inst = 32'h5be00000;
      38817: inst = 32'h8c50000;
      38818: inst = 32'h24612800;
      38819: inst = 32'h10a0ffff;
      38820: inst = 32'hca0ffe2;
      38821: inst = 32'h24822800;
      38822: inst = 32'h10a00000;
      38823: inst = 32'hca00004;
      38824: inst = 32'h38632800;
      38825: inst = 32'h38842800;
      38826: inst = 32'h10a00000;
      38827: inst = 32'hca097af;
      38828: inst = 32'h13e00001;
      38829: inst = 32'hfe0d96a;
      38830: inst = 32'h5be00000;
      38831: inst = 32'h8c50000;
      38832: inst = 32'h24612800;
      38833: inst = 32'h10a0ffff;
      38834: inst = 32'hca0ffe2;
      38835: inst = 32'h24822800;
      38836: inst = 32'h10a00000;
      38837: inst = 32'hca00004;
      38838: inst = 32'h38632800;
      38839: inst = 32'h38842800;
      38840: inst = 32'h10a00000;
      38841: inst = 32'hca097bd;
      38842: inst = 32'h13e00001;
      38843: inst = 32'hfe0d96a;
      38844: inst = 32'h5be00000;
      38845: inst = 32'h8c50000;
      38846: inst = 32'h24612800;
      38847: inst = 32'h10a0ffff;
      38848: inst = 32'hca0ffe2;
      38849: inst = 32'h24822800;
      38850: inst = 32'h10a00000;
      38851: inst = 32'hca00004;
      38852: inst = 32'h38632800;
      38853: inst = 32'h38842800;
      38854: inst = 32'h10a00000;
      38855: inst = 32'hca097cb;
      38856: inst = 32'h13e00001;
      38857: inst = 32'hfe0d96a;
      38858: inst = 32'h5be00000;
      38859: inst = 32'h8c50000;
      38860: inst = 32'h24612800;
      38861: inst = 32'h10a0ffff;
      38862: inst = 32'hca0ffe2;
      38863: inst = 32'h24822800;
      38864: inst = 32'h10a00000;
      38865: inst = 32'hca00004;
      38866: inst = 32'h38632800;
      38867: inst = 32'h38842800;
      38868: inst = 32'h10a00000;
      38869: inst = 32'hca097d9;
      38870: inst = 32'h13e00001;
      38871: inst = 32'hfe0d96a;
      38872: inst = 32'h5be00000;
      38873: inst = 32'h8c50000;
      38874: inst = 32'h24612800;
      38875: inst = 32'h10a0ffff;
      38876: inst = 32'hca0ffe2;
      38877: inst = 32'h24822800;
      38878: inst = 32'h10a00000;
      38879: inst = 32'hca00004;
      38880: inst = 32'h38632800;
      38881: inst = 32'h38842800;
      38882: inst = 32'h10a00000;
      38883: inst = 32'hca097e7;
      38884: inst = 32'h13e00001;
      38885: inst = 32'hfe0d96a;
      38886: inst = 32'h5be00000;
      38887: inst = 32'h8c50000;
      38888: inst = 32'h24612800;
      38889: inst = 32'h10a0ffff;
      38890: inst = 32'hca0ffe2;
      38891: inst = 32'h24822800;
      38892: inst = 32'h10a00000;
      38893: inst = 32'hca00004;
      38894: inst = 32'h38632800;
      38895: inst = 32'h38842800;
      38896: inst = 32'h10a00000;
      38897: inst = 32'hca097f5;
      38898: inst = 32'h13e00001;
      38899: inst = 32'hfe0d96a;
      38900: inst = 32'h5be00000;
      38901: inst = 32'h8c50000;
      38902: inst = 32'h24612800;
      38903: inst = 32'h10a0ffff;
      38904: inst = 32'hca0ffe2;
      38905: inst = 32'h24822800;
      38906: inst = 32'h10a00000;
      38907: inst = 32'hca00004;
      38908: inst = 32'h38632800;
      38909: inst = 32'h38842800;
      38910: inst = 32'h10a00000;
      38911: inst = 32'hca09803;
      38912: inst = 32'h13e00001;
      38913: inst = 32'hfe0d96a;
      38914: inst = 32'h5be00000;
      38915: inst = 32'h8c50000;
      38916: inst = 32'h24612800;
      38917: inst = 32'h10a0ffff;
      38918: inst = 32'hca0ffe2;
      38919: inst = 32'h24822800;
      38920: inst = 32'h10a00000;
      38921: inst = 32'hca00004;
      38922: inst = 32'h38632800;
      38923: inst = 32'h38842800;
      38924: inst = 32'h10a00000;
      38925: inst = 32'hca09811;
      38926: inst = 32'h13e00001;
      38927: inst = 32'hfe0d96a;
      38928: inst = 32'h5be00000;
      38929: inst = 32'h8c50000;
      38930: inst = 32'h24612800;
      38931: inst = 32'h10a0ffff;
      38932: inst = 32'hca0ffe2;
      38933: inst = 32'h24822800;
      38934: inst = 32'h10a00000;
      38935: inst = 32'hca00004;
      38936: inst = 32'h38632800;
      38937: inst = 32'h38842800;
      38938: inst = 32'h10a00000;
      38939: inst = 32'hca0981f;
      38940: inst = 32'h13e00001;
      38941: inst = 32'hfe0d96a;
      38942: inst = 32'h5be00000;
      38943: inst = 32'h8c50000;
      38944: inst = 32'h24612800;
      38945: inst = 32'h10a0ffff;
      38946: inst = 32'hca0ffe2;
      38947: inst = 32'h24822800;
      38948: inst = 32'h10a00000;
      38949: inst = 32'hca00004;
      38950: inst = 32'h38632800;
      38951: inst = 32'h38842800;
      38952: inst = 32'h10a00000;
      38953: inst = 32'hca0982d;
      38954: inst = 32'h13e00001;
      38955: inst = 32'hfe0d96a;
      38956: inst = 32'h5be00000;
      38957: inst = 32'h8c50000;
      38958: inst = 32'h24612800;
      38959: inst = 32'h10a0ffff;
      38960: inst = 32'hca0ffe2;
      38961: inst = 32'h24822800;
      38962: inst = 32'h10a00000;
      38963: inst = 32'hca00004;
      38964: inst = 32'h38632800;
      38965: inst = 32'h38842800;
      38966: inst = 32'h10a00000;
      38967: inst = 32'hca0983b;
      38968: inst = 32'h13e00001;
      38969: inst = 32'hfe0d96a;
      38970: inst = 32'h5be00000;
      38971: inst = 32'h8c50000;
      38972: inst = 32'h24612800;
      38973: inst = 32'h10a0ffff;
      38974: inst = 32'hca0ffe2;
      38975: inst = 32'h24822800;
      38976: inst = 32'h10a00000;
      38977: inst = 32'hca00004;
      38978: inst = 32'h38632800;
      38979: inst = 32'h38842800;
      38980: inst = 32'h10a00000;
      38981: inst = 32'hca09849;
      38982: inst = 32'h13e00001;
      38983: inst = 32'hfe0d96a;
      38984: inst = 32'h5be00000;
      38985: inst = 32'h8c50000;
      38986: inst = 32'h24612800;
      38987: inst = 32'h10a0ffff;
      38988: inst = 32'hca0ffe2;
      38989: inst = 32'h24822800;
      38990: inst = 32'h10a00000;
      38991: inst = 32'hca00004;
      38992: inst = 32'h38632800;
      38993: inst = 32'h38842800;
      38994: inst = 32'h10a00000;
      38995: inst = 32'hca09857;
      38996: inst = 32'h13e00001;
      38997: inst = 32'hfe0d96a;
      38998: inst = 32'h5be00000;
      38999: inst = 32'h8c50000;
      39000: inst = 32'h24612800;
      39001: inst = 32'h10a0ffff;
      39002: inst = 32'hca0ffe2;
      39003: inst = 32'h24822800;
      39004: inst = 32'h10a00000;
      39005: inst = 32'hca00004;
      39006: inst = 32'h38632800;
      39007: inst = 32'h38842800;
      39008: inst = 32'h10a00000;
      39009: inst = 32'hca09865;
      39010: inst = 32'h13e00001;
      39011: inst = 32'hfe0d96a;
      39012: inst = 32'h5be00000;
      39013: inst = 32'h8c50000;
      39014: inst = 32'h24612800;
      39015: inst = 32'h10a0ffff;
      39016: inst = 32'hca0ffe2;
      39017: inst = 32'h24822800;
      39018: inst = 32'h10a00000;
      39019: inst = 32'hca00004;
      39020: inst = 32'h38632800;
      39021: inst = 32'h38842800;
      39022: inst = 32'h10a00000;
      39023: inst = 32'hca09873;
      39024: inst = 32'h13e00001;
      39025: inst = 32'hfe0d96a;
      39026: inst = 32'h5be00000;
      39027: inst = 32'h8c50000;
      39028: inst = 32'h24612800;
      39029: inst = 32'h10a0ffff;
      39030: inst = 32'hca0ffe2;
      39031: inst = 32'h24822800;
      39032: inst = 32'h10a00000;
      39033: inst = 32'hca00004;
      39034: inst = 32'h38632800;
      39035: inst = 32'h38842800;
      39036: inst = 32'h10a00000;
      39037: inst = 32'hca09881;
      39038: inst = 32'h13e00001;
      39039: inst = 32'hfe0d96a;
      39040: inst = 32'h5be00000;
      39041: inst = 32'h8c50000;
      39042: inst = 32'h24612800;
      39043: inst = 32'h10a0ffff;
      39044: inst = 32'hca0ffe2;
      39045: inst = 32'h24822800;
      39046: inst = 32'h10a00000;
      39047: inst = 32'hca00004;
      39048: inst = 32'h38632800;
      39049: inst = 32'h38842800;
      39050: inst = 32'h10a00000;
      39051: inst = 32'hca0988f;
      39052: inst = 32'h13e00001;
      39053: inst = 32'hfe0d96a;
      39054: inst = 32'h5be00000;
      39055: inst = 32'h8c50000;
      39056: inst = 32'h24612800;
      39057: inst = 32'h10a0ffff;
      39058: inst = 32'hca0ffe2;
      39059: inst = 32'h24822800;
      39060: inst = 32'h10a00000;
      39061: inst = 32'hca00004;
      39062: inst = 32'h38632800;
      39063: inst = 32'h38842800;
      39064: inst = 32'h10a00000;
      39065: inst = 32'hca0989d;
      39066: inst = 32'h13e00001;
      39067: inst = 32'hfe0d96a;
      39068: inst = 32'h5be00000;
      39069: inst = 32'h8c50000;
      39070: inst = 32'h24612800;
      39071: inst = 32'h10a0ffff;
      39072: inst = 32'hca0ffe2;
      39073: inst = 32'h24822800;
      39074: inst = 32'h10a00000;
      39075: inst = 32'hca00004;
      39076: inst = 32'h38632800;
      39077: inst = 32'h38842800;
      39078: inst = 32'h10a00000;
      39079: inst = 32'hca098ab;
      39080: inst = 32'h13e00001;
      39081: inst = 32'hfe0d96a;
      39082: inst = 32'h5be00000;
      39083: inst = 32'h8c50000;
      39084: inst = 32'h24612800;
      39085: inst = 32'h10a0ffff;
      39086: inst = 32'hca0ffe2;
      39087: inst = 32'h24822800;
      39088: inst = 32'h10a00000;
      39089: inst = 32'hca00004;
      39090: inst = 32'h38632800;
      39091: inst = 32'h38842800;
      39092: inst = 32'h10a00000;
      39093: inst = 32'hca098b9;
      39094: inst = 32'h13e00001;
      39095: inst = 32'hfe0d96a;
      39096: inst = 32'h5be00000;
      39097: inst = 32'h8c50000;
      39098: inst = 32'h24612800;
      39099: inst = 32'h10a0ffff;
      39100: inst = 32'hca0ffe2;
      39101: inst = 32'h24822800;
      39102: inst = 32'h10a00000;
      39103: inst = 32'hca00004;
      39104: inst = 32'h38632800;
      39105: inst = 32'h38842800;
      39106: inst = 32'h10a00000;
      39107: inst = 32'hca098c7;
      39108: inst = 32'h13e00001;
      39109: inst = 32'hfe0d96a;
      39110: inst = 32'h5be00000;
      39111: inst = 32'h8c50000;
      39112: inst = 32'h24612800;
      39113: inst = 32'h10a0ffff;
      39114: inst = 32'hca0ffe2;
      39115: inst = 32'h24822800;
      39116: inst = 32'h10a00000;
      39117: inst = 32'hca00004;
      39118: inst = 32'h38632800;
      39119: inst = 32'h38842800;
      39120: inst = 32'h10a00000;
      39121: inst = 32'hca098d5;
      39122: inst = 32'h13e00001;
      39123: inst = 32'hfe0d96a;
      39124: inst = 32'h5be00000;
      39125: inst = 32'h8c50000;
      39126: inst = 32'h24612800;
      39127: inst = 32'h10a0ffff;
      39128: inst = 32'hca0ffe2;
      39129: inst = 32'h24822800;
      39130: inst = 32'h10a00000;
      39131: inst = 32'hca00004;
      39132: inst = 32'h38632800;
      39133: inst = 32'h38842800;
      39134: inst = 32'h10a00000;
      39135: inst = 32'hca098e3;
      39136: inst = 32'h13e00001;
      39137: inst = 32'hfe0d96a;
      39138: inst = 32'h5be00000;
      39139: inst = 32'h8c50000;
      39140: inst = 32'h24612800;
      39141: inst = 32'h10a0ffff;
      39142: inst = 32'hca0ffe2;
      39143: inst = 32'h24822800;
      39144: inst = 32'h10a00000;
      39145: inst = 32'hca00004;
      39146: inst = 32'h38632800;
      39147: inst = 32'h38842800;
      39148: inst = 32'h10a00000;
      39149: inst = 32'hca098f1;
      39150: inst = 32'h13e00001;
      39151: inst = 32'hfe0d96a;
      39152: inst = 32'h5be00000;
      39153: inst = 32'h8c50000;
      39154: inst = 32'h24612800;
      39155: inst = 32'h10a0ffff;
      39156: inst = 32'hca0ffe2;
      39157: inst = 32'h24822800;
      39158: inst = 32'h10a00000;
      39159: inst = 32'hca00004;
      39160: inst = 32'h38632800;
      39161: inst = 32'h38842800;
      39162: inst = 32'h10a00000;
      39163: inst = 32'hca098ff;
      39164: inst = 32'h13e00001;
      39165: inst = 32'hfe0d96a;
      39166: inst = 32'h5be00000;
      39167: inst = 32'h8c50000;
      39168: inst = 32'h24612800;
      39169: inst = 32'h10a0ffff;
      39170: inst = 32'hca0ffe2;
      39171: inst = 32'h24822800;
      39172: inst = 32'h10a00000;
      39173: inst = 32'hca00004;
      39174: inst = 32'h38632800;
      39175: inst = 32'h38842800;
      39176: inst = 32'h10a00000;
      39177: inst = 32'hca0990d;
      39178: inst = 32'h13e00001;
      39179: inst = 32'hfe0d96a;
      39180: inst = 32'h5be00000;
      39181: inst = 32'h8c50000;
      39182: inst = 32'h24612800;
      39183: inst = 32'h10a0ffff;
      39184: inst = 32'hca0ffe2;
      39185: inst = 32'h24822800;
      39186: inst = 32'h10a00000;
      39187: inst = 32'hca00004;
      39188: inst = 32'h38632800;
      39189: inst = 32'h38842800;
      39190: inst = 32'h10a00000;
      39191: inst = 32'hca0991b;
      39192: inst = 32'h13e00001;
      39193: inst = 32'hfe0d96a;
      39194: inst = 32'h5be00000;
      39195: inst = 32'h8c50000;
      39196: inst = 32'h24612800;
      39197: inst = 32'h10a0ffff;
      39198: inst = 32'hca0ffe2;
      39199: inst = 32'h24822800;
      39200: inst = 32'h10a00000;
      39201: inst = 32'hca00004;
      39202: inst = 32'h38632800;
      39203: inst = 32'h38842800;
      39204: inst = 32'h10a00000;
      39205: inst = 32'hca09929;
      39206: inst = 32'h13e00001;
      39207: inst = 32'hfe0d96a;
      39208: inst = 32'h5be00000;
      39209: inst = 32'h8c50000;
      39210: inst = 32'h24612800;
      39211: inst = 32'h10a0ffff;
      39212: inst = 32'hca0ffe3;
      39213: inst = 32'h24822800;
      39214: inst = 32'h10a00000;
      39215: inst = 32'hca00004;
      39216: inst = 32'h38632800;
      39217: inst = 32'h38842800;
      39218: inst = 32'h10a00000;
      39219: inst = 32'hca09937;
      39220: inst = 32'h13e00001;
      39221: inst = 32'hfe0d96a;
      39222: inst = 32'h5be00000;
      39223: inst = 32'h8c50000;
      39224: inst = 32'h24612800;
      39225: inst = 32'h10a0ffff;
      39226: inst = 32'hca0ffe3;
      39227: inst = 32'h24822800;
      39228: inst = 32'h10a00000;
      39229: inst = 32'hca00004;
      39230: inst = 32'h38632800;
      39231: inst = 32'h38842800;
      39232: inst = 32'h10a00000;
      39233: inst = 32'hca09945;
      39234: inst = 32'h13e00001;
      39235: inst = 32'hfe0d96a;
      39236: inst = 32'h5be00000;
      39237: inst = 32'h8c50000;
      39238: inst = 32'h24612800;
      39239: inst = 32'h10a0ffff;
      39240: inst = 32'hca0ffe3;
      39241: inst = 32'h24822800;
      39242: inst = 32'h10a00000;
      39243: inst = 32'hca00004;
      39244: inst = 32'h38632800;
      39245: inst = 32'h38842800;
      39246: inst = 32'h10a00000;
      39247: inst = 32'hca09953;
      39248: inst = 32'h13e00001;
      39249: inst = 32'hfe0d96a;
      39250: inst = 32'h5be00000;
      39251: inst = 32'h8c50000;
      39252: inst = 32'h24612800;
      39253: inst = 32'h10a0ffff;
      39254: inst = 32'hca0ffe3;
      39255: inst = 32'h24822800;
      39256: inst = 32'h10a00000;
      39257: inst = 32'hca00004;
      39258: inst = 32'h38632800;
      39259: inst = 32'h38842800;
      39260: inst = 32'h10a00000;
      39261: inst = 32'hca09961;
      39262: inst = 32'h13e00001;
      39263: inst = 32'hfe0d96a;
      39264: inst = 32'h5be00000;
      39265: inst = 32'h8c50000;
      39266: inst = 32'h24612800;
      39267: inst = 32'h10a0ffff;
      39268: inst = 32'hca0ffe3;
      39269: inst = 32'h24822800;
      39270: inst = 32'h10a00000;
      39271: inst = 32'hca00004;
      39272: inst = 32'h38632800;
      39273: inst = 32'h38842800;
      39274: inst = 32'h10a00000;
      39275: inst = 32'hca0996f;
      39276: inst = 32'h13e00001;
      39277: inst = 32'hfe0d96a;
      39278: inst = 32'h5be00000;
      39279: inst = 32'h8c50000;
      39280: inst = 32'h24612800;
      39281: inst = 32'h10a0ffff;
      39282: inst = 32'hca0ffe3;
      39283: inst = 32'h24822800;
      39284: inst = 32'h10a00000;
      39285: inst = 32'hca00004;
      39286: inst = 32'h38632800;
      39287: inst = 32'h38842800;
      39288: inst = 32'h10a00000;
      39289: inst = 32'hca0997d;
      39290: inst = 32'h13e00001;
      39291: inst = 32'hfe0d96a;
      39292: inst = 32'h5be00000;
      39293: inst = 32'h8c50000;
      39294: inst = 32'h24612800;
      39295: inst = 32'h10a0ffff;
      39296: inst = 32'hca0ffe3;
      39297: inst = 32'h24822800;
      39298: inst = 32'h10a00000;
      39299: inst = 32'hca00004;
      39300: inst = 32'h38632800;
      39301: inst = 32'h38842800;
      39302: inst = 32'h10a00000;
      39303: inst = 32'hca0998b;
      39304: inst = 32'h13e00001;
      39305: inst = 32'hfe0d96a;
      39306: inst = 32'h5be00000;
      39307: inst = 32'h8c50000;
      39308: inst = 32'h24612800;
      39309: inst = 32'h10a0ffff;
      39310: inst = 32'hca0ffe3;
      39311: inst = 32'h24822800;
      39312: inst = 32'h10a00000;
      39313: inst = 32'hca00004;
      39314: inst = 32'h38632800;
      39315: inst = 32'h38842800;
      39316: inst = 32'h10a00000;
      39317: inst = 32'hca09999;
      39318: inst = 32'h13e00001;
      39319: inst = 32'hfe0d96a;
      39320: inst = 32'h5be00000;
      39321: inst = 32'h8c50000;
      39322: inst = 32'h24612800;
      39323: inst = 32'h10a0ffff;
      39324: inst = 32'hca0ffe3;
      39325: inst = 32'h24822800;
      39326: inst = 32'h10a00000;
      39327: inst = 32'hca00004;
      39328: inst = 32'h38632800;
      39329: inst = 32'h38842800;
      39330: inst = 32'h10a00000;
      39331: inst = 32'hca099a7;
      39332: inst = 32'h13e00001;
      39333: inst = 32'hfe0d96a;
      39334: inst = 32'h5be00000;
      39335: inst = 32'h8c50000;
      39336: inst = 32'h24612800;
      39337: inst = 32'h10a0ffff;
      39338: inst = 32'hca0ffe3;
      39339: inst = 32'h24822800;
      39340: inst = 32'h10a00000;
      39341: inst = 32'hca00004;
      39342: inst = 32'h38632800;
      39343: inst = 32'h38842800;
      39344: inst = 32'h10a00000;
      39345: inst = 32'hca099b5;
      39346: inst = 32'h13e00001;
      39347: inst = 32'hfe0d96a;
      39348: inst = 32'h5be00000;
      39349: inst = 32'h8c50000;
      39350: inst = 32'h24612800;
      39351: inst = 32'h10a0ffff;
      39352: inst = 32'hca0ffe3;
      39353: inst = 32'h24822800;
      39354: inst = 32'h10a00000;
      39355: inst = 32'hca00004;
      39356: inst = 32'h38632800;
      39357: inst = 32'h38842800;
      39358: inst = 32'h10a00000;
      39359: inst = 32'hca099c3;
      39360: inst = 32'h13e00001;
      39361: inst = 32'hfe0d96a;
      39362: inst = 32'h5be00000;
      39363: inst = 32'h8c50000;
      39364: inst = 32'h24612800;
      39365: inst = 32'h10a0ffff;
      39366: inst = 32'hca0ffe3;
      39367: inst = 32'h24822800;
      39368: inst = 32'h10a00000;
      39369: inst = 32'hca00004;
      39370: inst = 32'h38632800;
      39371: inst = 32'h38842800;
      39372: inst = 32'h10a00000;
      39373: inst = 32'hca099d1;
      39374: inst = 32'h13e00001;
      39375: inst = 32'hfe0d96a;
      39376: inst = 32'h5be00000;
      39377: inst = 32'h8c50000;
      39378: inst = 32'h24612800;
      39379: inst = 32'h10a0ffff;
      39380: inst = 32'hca0ffe3;
      39381: inst = 32'h24822800;
      39382: inst = 32'h10a00000;
      39383: inst = 32'hca00004;
      39384: inst = 32'h38632800;
      39385: inst = 32'h38842800;
      39386: inst = 32'h10a00000;
      39387: inst = 32'hca099df;
      39388: inst = 32'h13e00001;
      39389: inst = 32'hfe0d96a;
      39390: inst = 32'h5be00000;
      39391: inst = 32'h8c50000;
      39392: inst = 32'h24612800;
      39393: inst = 32'h10a0ffff;
      39394: inst = 32'hca0ffe3;
      39395: inst = 32'h24822800;
      39396: inst = 32'h10a00000;
      39397: inst = 32'hca00004;
      39398: inst = 32'h38632800;
      39399: inst = 32'h38842800;
      39400: inst = 32'h10a00000;
      39401: inst = 32'hca099ed;
      39402: inst = 32'h13e00001;
      39403: inst = 32'hfe0d96a;
      39404: inst = 32'h5be00000;
      39405: inst = 32'h8c50000;
      39406: inst = 32'h24612800;
      39407: inst = 32'h10a0ffff;
      39408: inst = 32'hca0ffe3;
      39409: inst = 32'h24822800;
      39410: inst = 32'h10a00000;
      39411: inst = 32'hca00004;
      39412: inst = 32'h38632800;
      39413: inst = 32'h38842800;
      39414: inst = 32'h10a00000;
      39415: inst = 32'hca099fb;
      39416: inst = 32'h13e00001;
      39417: inst = 32'hfe0d96a;
      39418: inst = 32'h5be00000;
      39419: inst = 32'h8c50000;
      39420: inst = 32'h24612800;
      39421: inst = 32'h10a0ffff;
      39422: inst = 32'hca0ffe3;
      39423: inst = 32'h24822800;
      39424: inst = 32'h10a00000;
      39425: inst = 32'hca00004;
      39426: inst = 32'h38632800;
      39427: inst = 32'h38842800;
      39428: inst = 32'h10a00000;
      39429: inst = 32'hca09a09;
      39430: inst = 32'h13e00001;
      39431: inst = 32'hfe0d96a;
      39432: inst = 32'h5be00000;
      39433: inst = 32'h8c50000;
      39434: inst = 32'h24612800;
      39435: inst = 32'h10a0ffff;
      39436: inst = 32'hca0ffe3;
      39437: inst = 32'h24822800;
      39438: inst = 32'h10a00000;
      39439: inst = 32'hca00004;
      39440: inst = 32'h38632800;
      39441: inst = 32'h38842800;
      39442: inst = 32'h10a00000;
      39443: inst = 32'hca09a17;
      39444: inst = 32'h13e00001;
      39445: inst = 32'hfe0d96a;
      39446: inst = 32'h5be00000;
      39447: inst = 32'h8c50000;
      39448: inst = 32'h24612800;
      39449: inst = 32'h10a0ffff;
      39450: inst = 32'hca0ffe3;
      39451: inst = 32'h24822800;
      39452: inst = 32'h10a00000;
      39453: inst = 32'hca00004;
      39454: inst = 32'h38632800;
      39455: inst = 32'h38842800;
      39456: inst = 32'h10a00000;
      39457: inst = 32'hca09a25;
      39458: inst = 32'h13e00001;
      39459: inst = 32'hfe0d96a;
      39460: inst = 32'h5be00000;
      39461: inst = 32'h8c50000;
      39462: inst = 32'h24612800;
      39463: inst = 32'h10a0ffff;
      39464: inst = 32'hca0ffe3;
      39465: inst = 32'h24822800;
      39466: inst = 32'h10a00000;
      39467: inst = 32'hca00004;
      39468: inst = 32'h38632800;
      39469: inst = 32'h38842800;
      39470: inst = 32'h10a00000;
      39471: inst = 32'hca09a33;
      39472: inst = 32'h13e00001;
      39473: inst = 32'hfe0d96a;
      39474: inst = 32'h5be00000;
      39475: inst = 32'h8c50000;
      39476: inst = 32'h24612800;
      39477: inst = 32'h10a0ffff;
      39478: inst = 32'hca0ffe3;
      39479: inst = 32'h24822800;
      39480: inst = 32'h10a00000;
      39481: inst = 32'hca00004;
      39482: inst = 32'h38632800;
      39483: inst = 32'h38842800;
      39484: inst = 32'h10a00000;
      39485: inst = 32'hca09a41;
      39486: inst = 32'h13e00001;
      39487: inst = 32'hfe0d96a;
      39488: inst = 32'h5be00000;
      39489: inst = 32'h8c50000;
      39490: inst = 32'h24612800;
      39491: inst = 32'h10a0ffff;
      39492: inst = 32'hca0ffe3;
      39493: inst = 32'h24822800;
      39494: inst = 32'h10a00000;
      39495: inst = 32'hca00004;
      39496: inst = 32'h38632800;
      39497: inst = 32'h38842800;
      39498: inst = 32'h10a00000;
      39499: inst = 32'hca09a4f;
      39500: inst = 32'h13e00001;
      39501: inst = 32'hfe0d96a;
      39502: inst = 32'h5be00000;
      39503: inst = 32'h8c50000;
      39504: inst = 32'h24612800;
      39505: inst = 32'h10a0ffff;
      39506: inst = 32'hca0ffe3;
      39507: inst = 32'h24822800;
      39508: inst = 32'h10a00000;
      39509: inst = 32'hca00004;
      39510: inst = 32'h38632800;
      39511: inst = 32'h38842800;
      39512: inst = 32'h10a00000;
      39513: inst = 32'hca09a5d;
      39514: inst = 32'h13e00001;
      39515: inst = 32'hfe0d96a;
      39516: inst = 32'h5be00000;
      39517: inst = 32'h8c50000;
      39518: inst = 32'h24612800;
      39519: inst = 32'h10a0ffff;
      39520: inst = 32'hca0ffe3;
      39521: inst = 32'h24822800;
      39522: inst = 32'h10a00000;
      39523: inst = 32'hca00004;
      39524: inst = 32'h38632800;
      39525: inst = 32'h38842800;
      39526: inst = 32'h10a00000;
      39527: inst = 32'hca09a6b;
      39528: inst = 32'h13e00001;
      39529: inst = 32'hfe0d96a;
      39530: inst = 32'h5be00000;
      39531: inst = 32'h8c50000;
      39532: inst = 32'h24612800;
      39533: inst = 32'h10a0ffff;
      39534: inst = 32'hca0ffe3;
      39535: inst = 32'h24822800;
      39536: inst = 32'h10a00000;
      39537: inst = 32'hca00004;
      39538: inst = 32'h38632800;
      39539: inst = 32'h38842800;
      39540: inst = 32'h10a00000;
      39541: inst = 32'hca09a79;
      39542: inst = 32'h13e00001;
      39543: inst = 32'hfe0d96a;
      39544: inst = 32'h5be00000;
      39545: inst = 32'h8c50000;
      39546: inst = 32'h24612800;
      39547: inst = 32'h10a0ffff;
      39548: inst = 32'hca0ffe3;
      39549: inst = 32'h24822800;
      39550: inst = 32'h10a00000;
      39551: inst = 32'hca00004;
      39552: inst = 32'h38632800;
      39553: inst = 32'h38842800;
      39554: inst = 32'h10a00000;
      39555: inst = 32'hca09a87;
      39556: inst = 32'h13e00001;
      39557: inst = 32'hfe0d96a;
      39558: inst = 32'h5be00000;
      39559: inst = 32'h8c50000;
      39560: inst = 32'h24612800;
      39561: inst = 32'h10a0ffff;
      39562: inst = 32'hca0ffe3;
      39563: inst = 32'h24822800;
      39564: inst = 32'h10a00000;
      39565: inst = 32'hca00004;
      39566: inst = 32'h38632800;
      39567: inst = 32'h38842800;
      39568: inst = 32'h10a00000;
      39569: inst = 32'hca09a95;
      39570: inst = 32'h13e00001;
      39571: inst = 32'hfe0d96a;
      39572: inst = 32'h5be00000;
      39573: inst = 32'h8c50000;
      39574: inst = 32'h24612800;
      39575: inst = 32'h10a0ffff;
      39576: inst = 32'hca0ffe3;
      39577: inst = 32'h24822800;
      39578: inst = 32'h10a00000;
      39579: inst = 32'hca00004;
      39580: inst = 32'h38632800;
      39581: inst = 32'h38842800;
      39582: inst = 32'h10a00000;
      39583: inst = 32'hca09aa3;
      39584: inst = 32'h13e00001;
      39585: inst = 32'hfe0d96a;
      39586: inst = 32'h5be00000;
      39587: inst = 32'h8c50000;
      39588: inst = 32'h24612800;
      39589: inst = 32'h10a0ffff;
      39590: inst = 32'hca0ffe3;
      39591: inst = 32'h24822800;
      39592: inst = 32'h10a00000;
      39593: inst = 32'hca00004;
      39594: inst = 32'h38632800;
      39595: inst = 32'h38842800;
      39596: inst = 32'h10a00000;
      39597: inst = 32'hca09ab1;
      39598: inst = 32'h13e00001;
      39599: inst = 32'hfe0d96a;
      39600: inst = 32'h5be00000;
      39601: inst = 32'h8c50000;
      39602: inst = 32'h24612800;
      39603: inst = 32'h10a0ffff;
      39604: inst = 32'hca0ffe3;
      39605: inst = 32'h24822800;
      39606: inst = 32'h10a00000;
      39607: inst = 32'hca00004;
      39608: inst = 32'h38632800;
      39609: inst = 32'h38842800;
      39610: inst = 32'h10a00000;
      39611: inst = 32'hca09abf;
      39612: inst = 32'h13e00001;
      39613: inst = 32'hfe0d96a;
      39614: inst = 32'h5be00000;
      39615: inst = 32'h8c50000;
      39616: inst = 32'h24612800;
      39617: inst = 32'h10a0ffff;
      39618: inst = 32'hca0ffe3;
      39619: inst = 32'h24822800;
      39620: inst = 32'h10a00000;
      39621: inst = 32'hca00004;
      39622: inst = 32'h38632800;
      39623: inst = 32'h38842800;
      39624: inst = 32'h10a00000;
      39625: inst = 32'hca09acd;
      39626: inst = 32'h13e00001;
      39627: inst = 32'hfe0d96a;
      39628: inst = 32'h5be00000;
      39629: inst = 32'h8c50000;
      39630: inst = 32'h24612800;
      39631: inst = 32'h10a0ffff;
      39632: inst = 32'hca0ffe3;
      39633: inst = 32'h24822800;
      39634: inst = 32'h10a00000;
      39635: inst = 32'hca00004;
      39636: inst = 32'h38632800;
      39637: inst = 32'h38842800;
      39638: inst = 32'h10a00000;
      39639: inst = 32'hca09adb;
      39640: inst = 32'h13e00001;
      39641: inst = 32'hfe0d96a;
      39642: inst = 32'h5be00000;
      39643: inst = 32'h8c50000;
      39644: inst = 32'h24612800;
      39645: inst = 32'h10a0ffff;
      39646: inst = 32'hca0ffe3;
      39647: inst = 32'h24822800;
      39648: inst = 32'h10a00000;
      39649: inst = 32'hca00004;
      39650: inst = 32'h38632800;
      39651: inst = 32'h38842800;
      39652: inst = 32'h10a00000;
      39653: inst = 32'hca09ae9;
      39654: inst = 32'h13e00001;
      39655: inst = 32'hfe0d96a;
      39656: inst = 32'h5be00000;
      39657: inst = 32'h8c50000;
      39658: inst = 32'h24612800;
      39659: inst = 32'h10a0ffff;
      39660: inst = 32'hca0ffe3;
      39661: inst = 32'h24822800;
      39662: inst = 32'h10a00000;
      39663: inst = 32'hca00004;
      39664: inst = 32'h38632800;
      39665: inst = 32'h38842800;
      39666: inst = 32'h10a00000;
      39667: inst = 32'hca09af7;
      39668: inst = 32'h13e00001;
      39669: inst = 32'hfe0d96a;
      39670: inst = 32'h5be00000;
      39671: inst = 32'h8c50000;
      39672: inst = 32'h24612800;
      39673: inst = 32'h10a0ffff;
      39674: inst = 32'hca0ffe3;
      39675: inst = 32'h24822800;
      39676: inst = 32'h10a00000;
      39677: inst = 32'hca00004;
      39678: inst = 32'h38632800;
      39679: inst = 32'h38842800;
      39680: inst = 32'h10a00000;
      39681: inst = 32'hca09b05;
      39682: inst = 32'h13e00001;
      39683: inst = 32'hfe0d96a;
      39684: inst = 32'h5be00000;
      39685: inst = 32'h8c50000;
      39686: inst = 32'h24612800;
      39687: inst = 32'h10a0ffff;
      39688: inst = 32'hca0ffe3;
      39689: inst = 32'h24822800;
      39690: inst = 32'h10a00000;
      39691: inst = 32'hca00004;
      39692: inst = 32'h38632800;
      39693: inst = 32'h38842800;
      39694: inst = 32'h10a00000;
      39695: inst = 32'hca09b13;
      39696: inst = 32'h13e00001;
      39697: inst = 32'hfe0d96a;
      39698: inst = 32'h5be00000;
      39699: inst = 32'h8c50000;
      39700: inst = 32'h24612800;
      39701: inst = 32'h10a0ffff;
      39702: inst = 32'hca0ffe3;
      39703: inst = 32'h24822800;
      39704: inst = 32'h10a00000;
      39705: inst = 32'hca00004;
      39706: inst = 32'h38632800;
      39707: inst = 32'h38842800;
      39708: inst = 32'h10a00000;
      39709: inst = 32'hca09b21;
      39710: inst = 32'h13e00001;
      39711: inst = 32'hfe0d96a;
      39712: inst = 32'h5be00000;
      39713: inst = 32'h8c50000;
      39714: inst = 32'h24612800;
      39715: inst = 32'h10a0ffff;
      39716: inst = 32'hca0ffe3;
      39717: inst = 32'h24822800;
      39718: inst = 32'h10a00000;
      39719: inst = 32'hca00004;
      39720: inst = 32'h38632800;
      39721: inst = 32'h38842800;
      39722: inst = 32'h10a00000;
      39723: inst = 32'hca09b2f;
      39724: inst = 32'h13e00001;
      39725: inst = 32'hfe0d96a;
      39726: inst = 32'h5be00000;
      39727: inst = 32'h8c50000;
      39728: inst = 32'h24612800;
      39729: inst = 32'h10a0ffff;
      39730: inst = 32'hca0ffe3;
      39731: inst = 32'h24822800;
      39732: inst = 32'h10a00000;
      39733: inst = 32'hca00004;
      39734: inst = 32'h38632800;
      39735: inst = 32'h38842800;
      39736: inst = 32'h10a00000;
      39737: inst = 32'hca09b3d;
      39738: inst = 32'h13e00001;
      39739: inst = 32'hfe0d96a;
      39740: inst = 32'h5be00000;
      39741: inst = 32'h8c50000;
      39742: inst = 32'h24612800;
      39743: inst = 32'h10a0ffff;
      39744: inst = 32'hca0ffe3;
      39745: inst = 32'h24822800;
      39746: inst = 32'h10a00000;
      39747: inst = 32'hca00004;
      39748: inst = 32'h38632800;
      39749: inst = 32'h38842800;
      39750: inst = 32'h10a00000;
      39751: inst = 32'hca09b4b;
      39752: inst = 32'h13e00001;
      39753: inst = 32'hfe0d96a;
      39754: inst = 32'h5be00000;
      39755: inst = 32'h8c50000;
      39756: inst = 32'h24612800;
      39757: inst = 32'h10a0ffff;
      39758: inst = 32'hca0ffe3;
      39759: inst = 32'h24822800;
      39760: inst = 32'h10a00000;
      39761: inst = 32'hca00004;
      39762: inst = 32'h38632800;
      39763: inst = 32'h38842800;
      39764: inst = 32'h10a00000;
      39765: inst = 32'hca09b59;
      39766: inst = 32'h13e00001;
      39767: inst = 32'hfe0d96a;
      39768: inst = 32'h5be00000;
      39769: inst = 32'h8c50000;
      39770: inst = 32'h24612800;
      39771: inst = 32'h10a0ffff;
      39772: inst = 32'hca0ffe3;
      39773: inst = 32'h24822800;
      39774: inst = 32'h10a00000;
      39775: inst = 32'hca00004;
      39776: inst = 32'h38632800;
      39777: inst = 32'h38842800;
      39778: inst = 32'h10a00000;
      39779: inst = 32'hca09b67;
      39780: inst = 32'h13e00001;
      39781: inst = 32'hfe0d96a;
      39782: inst = 32'h5be00000;
      39783: inst = 32'h8c50000;
      39784: inst = 32'h24612800;
      39785: inst = 32'h10a0ffff;
      39786: inst = 32'hca0ffe3;
      39787: inst = 32'h24822800;
      39788: inst = 32'h10a00000;
      39789: inst = 32'hca00004;
      39790: inst = 32'h38632800;
      39791: inst = 32'h38842800;
      39792: inst = 32'h10a00000;
      39793: inst = 32'hca09b75;
      39794: inst = 32'h13e00001;
      39795: inst = 32'hfe0d96a;
      39796: inst = 32'h5be00000;
      39797: inst = 32'h8c50000;
      39798: inst = 32'h24612800;
      39799: inst = 32'h10a0ffff;
      39800: inst = 32'hca0ffe3;
      39801: inst = 32'h24822800;
      39802: inst = 32'h10a00000;
      39803: inst = 32'hca00004;
      39804: inst = 32'h38632800;
      39805: inst = 32'h38842800;
      39806: inst = 32'h10a00000;
      39807: inst = 32'hca09b83;
      39808: inst = 32'h13e00001;
      39809: inst = 32'hfe0d96a;
      39810: inst = 32'h5be00000;
      39811: inst = 32'h8c50000;
      39812: inst = 32'h24612800;
      39813: inst = 32'h10a0ffff;
      39814: inst = 32'hca0ffe3;
      39815: inst = 32'h24822800;
      39816: inst = 32'h10a00000;
      39817: inst = 32'hca00004;
      39818: inst = 32'h38632800;
      39819: inst = 32'h38842800;
      39820: inst = 32'h10a00000;
      39821: inst = 32'hca09b91;
      39822: inst = 32'h13e00001;
      39823: inst = 32'hfe0d96a;
      39824: inst = 32'h5be00000;
      39825: inst = 32'h8c50000;
      39826: inst = 32'h24612800;
      39827: inst = 32'h10a0ffff;
      39828: inst = 32'hca0ffe3;
      39829: inst = 32'h24822800;
      39830: inst = 32'h10a00000;
      39831: inst = 32'hca00004;
      39832: inst = 32'h38632800;
      39833: inst = 32'h38842800;
      39834: inst = 32'h10a00000;
      39835: inst = 32'hca09b9f;
      39836: inst = 32'h13e00001;
      39837: inst = 32'hfe0d96a;
      39838: inst = 32'h5be00000;
      39839: inst = 32'h8c50000;
      39840: inst = 32'h24612800;
      39841: inst = 32'h10a0ffff;
      39842: inst = 32'hca0ffe3;
      39843: inst = 32'h24822800;
      39844: inst = 32'h10a00000;
      39845: inst = 32'hca00004;
      39846: inst = 32'h38632800;
      39847: inst = 32'h38842800;
      39848: inst = 32'h10a00000;
      39849: inst = 32'hca09bad;
      39850: inst = 32'h13e00001;
      39851: inst = 32'hfe0d96a;
      39852: inst = 32'h5be00000;
      39853: inst = 32'h8c50000;
      39854: inst = 32'h24612800;
      39855: inst = 32'h10a0ffff;
      39856: inst = 32'hca0ffe3;
      39857: inst = 32'h24822800;
      39858: inst = 32'h10a00000;
      39859: inst = 32'hca00004;
      39860: inst = 32'h38632800;
      39861: inst = 32'h38842800;
      39862: inst = 32'h10a00000;
      39863: inst = 32'hca09bbb;
      39864: inst = 32'h13e00001;
      39865: inst = 32'hfe0d96a;
      39866: inst = 32'h5be00000;
      39867: inst = 32'h8c50000;
      39868: inst = 32'h24612800;
      39869: inst = 32'h10a0ffff;
      39870: inst = 32'hca0ffe3;
      39871: inst = 32'h24822800;
      39872: inst = 32'h10a00000;
      39873: inst = 32'hca00004;
      39874: inst = 32'h38632800;
      39875: inst = 32'h38842800;
      39876: inst = 32'h10a00000;
      39877: inst = 32'hca09bc9;
      39878: inst = 32'h13e00001;
      39879: inst = 32'hfe0d96a;
      39880: inst = 32'h5be00000;
      39881: inst = 32'h8c50000;
      39882: inst = 32'h24612800;
      39883: inst = 32'h10a0ffff;
      39884: inst = 32'hca0ffe3;
      39885: inst = 32'h24822800;
      39886: inst = 32'h10a00000;
      39887: inst = 32'hca00004;
      39888: inst = 32'h38632800;
      39889: inst = 32'h38842800;
      39890: inst = 32'h10a00000;
      39891: inst = 32'hca09bd7;
      39892: inst = 32'h13e00001;
      39893: inst = 32'hfe0d96a;
      39894: inst = 32'h5be00000;
      39895: inst = 32'h8c50000;
      39896: inst = 32'h24612800;
      39897: inst = 32'h10a0ffff;
      39898: inst = 32'hca0ffe3;
      39899: inst = 32'h24822800;
      39900: inst = 32'h10a00000;
      39901: inst = 32'hca00004;
      39902: inst = 32'h38632800;
      39903: inst = 32'h38842800;
      39904: inst = 32'h10a00000;
      39905: inst = 32'hca09be5;
      39906: inst = 32'h13e00001;
      39907: inst = 32'hfe0d96a;
      39908: inst = 32'h5be00000;
      39909: inst = 32'h8c50000;
      39910: inst = 32'h24612800;
      39911: inst = 32'h10a0ffff;
      39912: inst = 32'hca0ffe3;
      39913: inst = 32'h24822800;
      39914: inst = 32'h10a00000;
      39915: inst = 32'hca00004;
      39916: inst = 32'h38632800;
      39917: inst = 32'h38842800;
      39918: inst = 32'h10a00000;
      39919: inst = 32'hca09bf3;
      39920: inst = 32'h13e00001;
      39921: inst = 32'hfe0d96a;
      39922: inst = 32'h5be00000;
      39923: inst = 32'h8c50000;
      39924: inst = 32'h24612800;
      39925: inst = 32'h10a0ffff;
      39926: inst = 32'hca0ffe3;
      39927: inst = 32'h24822800;
      39928: inst = 32'h10a00000;
      39929: inst = 32'hca00004;
      39930: inst = 32'h38632800;
      39931: inst = 32'h38842800;
      39932: inst = 32'h10a00000;
      39933: inst = 32'hca09c01;
      39934: inst = 32'h13e00001;
      39935: inst = 32'hfe0d96a;
      39936: inst = 32'h5be00000;
      39937: inst = 32'h8c50000;
      39938: inst = 32'h24612800;
      39939: inst = 32'h10a0ffff;
      39940: inst = 32'hca0ffe3;
      39941: inst = 32'h24822800;
      39942: inst = 32'h10a00000;
      39943: inst = 32'hca00004;
      39944: inst = 32'h38632800;
      39945: inst = 32'h38842800;
      39946: inst = 32'h10a00000;
      39947: inst = 32'hca09c0f;
      39948: inst = 32'h13e00001;
      39949: inst = 32'hfe0d96a;
      39950: inst = 32'h5be00000;
      39951: inst = 32'h8c50000;
      39952: inst = 32'h24612800;
      39953: inst = 32'h10a0ffff;
      39954: inst = 32'hca0ffe3;
      39955: inst = 32'h24822800;
      39956: inst = 32'h10a00000;
      39957: inst = 32'hca00004;
      39958: inst = 32'h38632800;
      39959: inst = 32'h38842800;
      39960: inst = 32'h10a00000;
      39961: inst = 32'hca09c1d;
      39962: inst = 32'h13e00001;
      39963: inst = 32'hfe0d96a;
      39964: inst = 32'h5be00000;
      39965: inst = 32'h8c50000;
      39966: inst = 32'h24612800;
      39967: inst = 32'h10a0ffff;
      39968: inst = 32'hca0ffe3;
      39969: inst = 32'h24822800;
      39970: inst = 32'h10a00000;
      39971: inst = 32'hca00004;
      39972: inst = 32'h38632800;
      39973: inst = 32'h38842800;
      39974: inst = 32'h10a00000;
      39975: inst = 32'hca09c2b;
      39976: inst = 32'h13e00001;
      39977: inst = 32'hfe0d96a;
      39978: inst = 32'h5be00000;
      39979: inst = 32'h8c50000;
      39980: inst = 32'h24612800;
      39981: inst = 32'h10a0ffff;
      39982: inst = 32'hca0ffe3;
      39983: inst = 32'h24822800;
      39984: inst = 32'h10a00000;
      39985: inst = 32'hca00004;
      39986: inst = 32'h38632800;
      39987: inst = 32'h38842800;
      39988: inst = 32'h10a00000;
      39989: inst = 32'hca09c39;
      39990: inst = 32'h13e00001;
      39991: inst = 32'hfe0d96a;
      39992: inst = 32'h5be00000;
      39993: inst = 32'h8c50000;
      39994: inst = 32'h24612800;
      39995: inst = 32'h10a0ffff;
      39996: inst = 32'hca0ffe3;
      39997: inst = 32'h24822800;
      39998: inst = 32'h10a00000;
      39999: inst = 32'hca00004;
      40000: inst = 32'h38632800;
      40001: inst = 32'h38842800;
      40002: inst = 32'h10a00000;
      40003: inst = 32'hca09c47;
      40004: inst = 32'h13e00001;
      40005: inst = 32'hfe0d96a;
      40006: inst = 32'h5be00000;
      40007: inst = 32'h8c50000;
      40008: inst = 32'h24612800;
      40009: inst = 32'h10a0ffff;
      40010: inst = 32'hca0ffe3;
      40011: inst = 32'h24822800;
      40012: inst = 32'h10a00000;
      40013: inst = 32'hca00004;
      40014: inst = 32'h38632800;
      40015: inst = 32'h38842800;
      40016: inst = 32'h10a00000;
      40017: inst = 32'hca09c55;
      40018: inst = 32'h13e00001;
      40019: inst = 32'hfe0d96a;
      40020: inst = 32'h5be00000;
      40021: inst = 32'h8c50000;
      40022: inst = 32'h24612800;
      40023: inst = 32'h10a0ffff;
      40024: inst = 32'hca0ffe3;
      40025: inst = 32'h24822800;
      40026: inst = 32'h10a00000;
      40027: inst = 32'hca00004;
      40028: inst = 32'h38632800;
      40029: inst = 32'h38842800;
      40030: inst = 32'h10a00000;
      40031: inst = 32'hca09c63;
      40032: inst = 32'h13e00001;
      40033: inst = 32'hfe0d96a;
      40034: inst = 32'h5be00000;
      40035: inst = 32'h8c50000;
      40036: inst = 32'h24612800;
      40037: inst = 32'h10a0ffff;
      40038: inst = 32'hca0ffe3;
      40039: inst = 32'h24822800;
      40040: inst = 32'h10a00000;
      40041: inst = 32'hca00004;
      40042: inst = 32'h38632800;
      40043: inst = 32'h38842800;
      40044: inst = 32'h10a00000;
      40045: inst = 32'hca09c71;
      40046: inst = 32'h13e00001;
      40047: inst = 32'hfe0d96a;
      40048: inst = 32'h5be00000;
      40049: inst = 32'h8c50000;
      40050: inst = 32'h24612800;
      40051: inst = 32'h10a0ffff;
      40052: inst = 32'hca0ffe3;
      40053: inst = 32'h24822800;
      40054: inst = 32'h10a00000;
      40055: inst = 32'hca00004;
      40056: inst = 32'h38632800;
      40057: inst = 32'h38842800;
      40058: inst = 32'h10a00000;
      40059: inst = 32'hca09c7f;
      40060: inst = 32'h13e00001;
      40061: inst = 32'hfe0d96a;
      40062: inst = 32'h5be00000;
      40063: inst = 32'h8c50000;
      40064: inst = 32'h24612800;
      40065: inst = 32'h10a0ffff;
      40066: inst = 32'hca0ffe3;
      40067: inst = 32'h24822800;
      40068: inst = 32'h10a00000;
      40069: inst = 32'hca00004;
      40070: inst = 32'h38632800;
      40071: inst = 32'h38842800;
      40072: inst = 32'h10a00000;
      40073: inst = 32'hca09c8d;
      40074: inst = 32'h13e00001;
      40075: inst = 32'hfe0d96a;
      40076: inst = 32'h5be00000;
      40077: inst = 32'h8c50000;
      40078: inst = 32'h24612800;
      40079: inst = 32'h10a0ffff;
      40080: inst = 32'hca0ffe3;
      40081: inst = 32'h24822800;
      40082: inst = 32'h10a00000;
      40083: inst = 32'hca00004;
      40084: inst = 32'h38632800;
      40085: inst = 32'h38842800;
      40086: inst = 32'h10a00000;
      40087: inst = 32'hca09c9b;
      40088: inst = 32'h13e00001;
      40089: inst = 32'hfe0d96a;
      40090: inst = 32'h5be00000;
      40091: inst = 32'h8c50000;
      40092: inst = 32'h24612800;
      40093: inst = 32'h10a0ffff;
      40094: inst = 32'hca0ffe3;
      40095: inst = 32'h24822800;
      40096: inst = 32'h10a00000;
      40097: inst = 32'hca00004;
      40098: inst = 32'h38632800;
      40099: inst = 32'h38842800;
      40100: inst = 32'h10a00000;
      40101: inst = 32'hca09ca9;
      40102: inst = 32'h13e00001;
      40103: inst = 32'hfe0d96a;
      40104: inst = 32'h5be00000;
      40105: inst = 32'h8c50000;
      40106: inst = 32'h24612800;
      40107: inst = 32'h10a0ffff;
      40108: inst = 32'hca0ffe3;
      40109: inst = 32'h24822800;
      40110: inst = 32'h10a00000;
      40111: inst = 32'hca00004;
      40112: inst = 32'h38632800;
      40113: inst = 32'h38842800;
      40114: inst = 32'h10a00000;
      40115: inst = 32'hca09cb7;
      40116: inst = 32'h13e00001;
      40117: inst = 32'hfe0d96a;
      40118: inst = 32'h5be00000;
      40119: inst = 32'h8c50000;
      40120: inst = 32'h24612800;
      40121: inst = 32'h10a0ffff;
      40122: inst = 32'hca0ffe3;
      40123: inst = 32'h24822800;
      40124: inst = 32'h10a00000;
      40125: inst = 32'hca00004;
      40126: inst = 32'h38632800;
      40127: inst = 32'h38842800;
      40128: inst = 32'h10a00000;
      40129: inst = 32'hca09cc5;
      40130: inst = 32'h13e00001;
      40131: inst = 32'hfe0d96a;
      40132: inst = 32'h5be00000;
      40133: inst = 32'h8c50000;
      40134: inst = 32'h24612800;
      40135: inst = 32'h10a0ffff;
      40136: inst = 32'hca0ffe3;
      40137: inst = 32'h24822800;
      40138: inst = 32'h10a00000;
      40139: inst = 32'hca00004;
      40140: inst = 32'h38632800;
      40141: inst = 32'h38842800;
      40142: inst = 32'h10a00000;
      40143: inst = 32'hca09cd3;
      40144: inst = 32'h13e00001;
      40145: inst = 32'hfe0d96a;
      40146: inst = 32'h5be00000;
      40147: inst = 32'h8c50000;
      40148: inst = 32'h24612800;
      40149: inst = 32'h10a0ffff;
      40150: inst = 32'hca0ffe3;
      40151: inst = 32'h24822800;
      40152: inst = 32'h10a00000;
      40153: inst = 32'hca00004;
      40154: inst = 32'h38632800;
      40155: inst = 32'h38842800;
      40156: inst = 32'h10a00000;
      40157: inst = 32'hca09ce1;
      40158: inst = 32'h13e00001;
      40159: inst = 32'hfe0d96a;
      40160: inst = 32'h5be00000;
      40161: inst = 32'h8c50000;
      40162: inst = 32'h24612800;
      40163: inst = 32'h10a0ffff;
      40164: inst = 32'hca0ffe3;
      40165: inst = 32'h24822800;
      40166: inst = 32'h10a00000;
      40167: inst = 32'hca00004;
      40168: inst = 32'h38632800;
      40169: inst = 32'h38842800;
      40170: inst = 32'h10a00000;
      40171: inst = 32'hca09cef;
      40172: inst = 32'h13e00001;
      40173: inst = 32'hfe0d96a;
      40174: inst = 32'h5be00000;
      40175: inst = 32'h8c50000;
      40176: inst = 32'h24612800;
      40177: inst = 32'h10a0ffff;
      40178: inst = 32'hca0ffe3;
      40179: inst = 32'h24822800;
      40180: inst = 32'h10a00000;
      40181: inst = 32'hca00004;
      40182: inst = 32'h38632800;
      40183: inst = 32'h38842800;
      40184: inst = 32'h10a00000;
      40185: inst = 32'hca09cfd;
      40186: inst = 32'h13e00001;
      40187: inst = 32'hfe0d96a;
      40188: inst = 32'h5be00000;
      40189: inst = 32'h8c50000;
      40190: inst = 32'h24612800;
      40191: inst = 32'h10a0ffff;
      40192: inst = 32'hca0ffe3;
      40193: inst = 32'h24822800;
      40194: inst = 32'h10a00000;
      40195: inst = 32'hca00004;
      40196: inst = 32'h38632800;
      40197: inst = 32'h38842800;
      40198: inst = 32'h10a00000;
      40199: inst = 32'hca09d0b;
      40200: inst = 32'h13e00001;
      40201: inst = 32'hfe0d96a;
      40202: inst = 32'h5be00000;
      40203: inst = 32'h8c50000;
      40204: inst = 32'h24612800;
      40205: inst = 32'h10a0ffff;
      40206: inst = 32'hca0ffe3;
      40207: inst = 32'h24822800;
      40208: inst = 32'h10a00000;
      40209: inst = 32'hca00004;
      40210: inst = 32'h38632800;
      40211: inst = 32'h38842800;
      40212: inst = 32'h10a00000;
      40213: inst = 32'hca09d19;
      40214: inst = 32'h13e00001;
      40215: inst = 32'hfe0d96a;
      40216: inst = 32'h5be00000;
      40217: inst = 32'h8c50000;
      40218: inst = 32'h24612800;
      40219: inst = 32'h10a0ffff;
      40220: inst = 32'hca0ffe3;
      40221: inst = 32'h24822800;
      40222: inst = 32'h10a00000;
      40223: inst = 32'hca00004;
      40224: inst = 32'h38632800;
      40225: inst = 32'h38842800;
      40226: inst = 32'h10a00000;
      40227: inst = 32'hca09d27;
      40228: inst = 32'h13e00001;
      40229: inst = 32'hfe0d96a;
      40230: inst = 32'h5be00000;
      40231: inst = 32'h8c50000;
      40232: inst = 32'h24612800;
      40233: inst = 32'h10a0ffff;
      40234: inst = 32'hca0ffe3;
      40235: inst = 32'h24822800;
      40236: inst = 32'h10a00000;
      40237: inst = 32'hca00004;
      40238: inst = 32'h38632800;
      40239: inst = 32'h38842800;
      40240: inst = 32'h10a00000;
      40241: inst = 32'hca09d35;
      40242: inst = 32'h13e00001;
      40243: inst = 32'hfe0d96a;
      40244: inst = 32'h5be00000;
      40245: inst = 32'h8c50000;
      40246: inst = 32'h24612800;
      40247: inst = 32'h10a0ffff;
      40248: inst = 32'hca0ffe3;
      40249: inst = 32'h24822800;
      40250: inst = 32'h10a00000;
      40251: inst = 32'hca00004;
      40252: inst = 32'h38632800;
      40253: inst = 32'h38842800;
      40254: inst = 32'h10a00000;
      40255: inst = 32'hca09d43;
      40256: inst = 32'h13e00001;
      40257: inst = 32'hfe0d96a;
      40258: inst = 32'h5be00000;
      40259: inst = 32'h8c50000;
      40260: inst = 32'h24612800;
      40261: inst = 32'h10a0ffff;
      40262: inst = 32'hca0ffe3;
      40263: inst = 32'h24822800;
      40264: inst = 32'h10a00000;
      40265: inst = 32'hca00004;
      40266: inst = 32'h38632800;
      40267: inst = 32'h38842800;
      40268: inst = 32'h10a00000;
      40269: inst = 32'hca09d51;
      40270: inst = 32'h13e00001;
      40271: inst = 32'hfe0d96a;
      40272: inst = 32'h5be00000;
      40273: inst = 32'h8c50000;
      40274: inst = 32'h24612800;
      40275: inst = 32'h10a0ffff;
      40276: inst = 32'hca0ffe3;
      40277: inst = 32'h24822800;
      40278: inst = 32'h10a00000;
      40279: inst = 32'hca00004;
      40280: inst = 32'h38632800;
      40281: inst = 32'h38842800;
      40282: inst = 32'h10a00000;
      40283: inst = 32'hca09d5f;
      40284: inst = 32'h13e00001;
      40285: inst = 32'hfe0d96a;
      40286: inst = 32'h5be00000;
      40287: inst = 32'h8c50000;
      40288: inst = 32'h24612800;
      40289: inst = 32'h10a0ffff;
      40290: inst = 32'hca0ffe3;
      40291: inst = 32'h24822800;
      40292: inst = 32'h10a00000;
      40293: inst = 32'hca00004;
      40294: inst = 32'h38632800;
      40295: inst = 32'h38842800;
      40296: inst = 32'h10a00000;
      40297: inst = 32'hca09d6d;
      40298: inst = 32'h13e00001;
      40299: inst = 32'hfe0d96a;
      40300: inst = 32'h5be00000;
      40301: inst = 32'h8c50000;
      40302: inst = 32'h24612800;
      40303: inst = 32'h10a0ffff;
      40304: inst = 32'hca0ffe3;
      40305: inst = 32'h24822800;
      40306: inst = 32'h10a00000;
      40307: inst = 32'hca00004;
      40308: inst = 32'h38632800;
      40309: inst = 32'h38842800;
      40310: inst = 32'h10a00000;
      40311: inst = 32'hca09d7b;
      40312: inst = 32'h13e00001;
      40313: inst = 32'hfe0d96a;
      40314: inst = 32'h5be00000;
      40315: inst = 32'h8c50000;
      40316: inst = 32'h24612800;
      40317: inst = 32'h10a0ffff;
      40318: inst = 32'hca0ffe3;
      40319: inst = 32'h24822800;
      40320: inst = 32'h10a00000;
      40321: inst = 32'hca00004;
      40322: inst = 32'h38632800;
      40323: inst = 32'h38842800;
      40324: inst = 32'h10a00000;
      40325: inst = 32'hca09d89;
      40326: inst = 32'h13e00001;
      40327: inst = 32'hfe0d96a;
      40328: inst = 32'h5be00000;
      40329: inst = 32'h8c50000;
      40330: inst = 32'h24612800;
      40331: inst = 32'h10a0ffff;
      40332: inst = 32'hca0ffe3;
      40333: inst = 32'h24822800;
      40334: inst = 32'h10a00000;
      40335: inst = 32'hca00004;
      40336: inst = 32'h38632800;
      40337: inst = 32'h38842800;
      40338: inst = 32'h10a00000;
      40339: inst = 32'hca09d97;
      40340: inst = 32'h13e00001;
      40341: inst = 32'hfe0d96a;
      40342: inst = 32'h5be00000;
      40343: inst = 32'h8c50000;
      40344: inst = 32'h24612800;
      40345: inst = 32'h10a0ffff;
      40346: inst = 32'hca0ffe3;
      40347: inst = 32'h24822800;
      40348: inst = 32'h10a00000;
      40349: inst = 32'hca00004;
      40350: inst = 32'h38632800;
      40351: inst = 32'h38842800;
      40352: inst = 32'h10a00000;
      40353: inst = 32'hca09da5;
      40354: inst = 32'h13e00001;
      40355: inst = 32'hfe0d96a;
      40356: inst = 32'h5be00000;
      40357: inst = 32'h8c50000;
      40358: inst = 32'h24612800;
      40359: inst = 32'h10a0ffff;
      40360: inst = 32'hca0ffe3;
      40361: inst = 32'h24822800;
      40362: inst = 32'h10a00000;
      40363: inst = 32'hca00004;
      40364: inst = 32'h38632800;
      40365: inst = 32'h38842800;
      40366: inst = 32'h10a00000;
      40367: inst = 32'hca09db3;
      40368: inst = 32'h13e00001;
      40369: inst = 32'hfe0d96a;
      40370: inst = 32'h5be00000;
      40371: inst = 32'h8c50000;
      40372: inst = 32'h24612800;
      40373: inst = 32'h10a0ffff;
      40374: inst = 32'hca0ffe3;
      40375: inst = 32'h24822800;
      40376: inst = 32'h10a00000;
      40377: inst = 32'hca00004;
      40378: inst = 32'h38632800;
      40379: inst = 32'h38842800;
      40380: inst = 32'h10a00000;
      40381: inst = 32'hca09dc1;
      40382: inst = 32'h13e00001;
      40383: inst = 32'hfe0d96a;
      40384: inst = 32'h5be00000;
      40385: inst = 32'h8c50000;
      40386: inst = 32'h24612800;
      40387: inst = 32'h10a0ffff;
      40388: inst = 32'hca0ffe3;
      40389: inst = 32'h24822800;
      40390: inst = 32'h10a00000;
      40391: inst = 32'hca00004;
      40392: inst = 32'h38632800;
      40393: inst = 32'h38842800;
      40394: inst = 32'h10a00000;
      40395: inst = 32'hca09dcf;
      40396: inst = 32'h13e00001;
      40397: inst = 32'hfe0d96a;
      40398: inst = 32'h5be00000;
      40399: inst = 32'h8c50000;
      40400: inst = 32'h24612800;
      40401: inst = 32'h10a0ffff;
      40402: inst = 32'hca0ffe3;
      40403: inst = 32'h24822800;
      40404: inst = 32'h10a00000;
      40405: inst = 32'hca00004;
      40406: inst = 32'h38632800;
      40407: inst = 32'h38842800;
      40408: inst = 32'h10a00000;
      40409: inst = 32'hca09ddd;
      40410: inst = 32'h13e00001;
      40411: inst = 32'hfe0d96a;
      40412: inst = 32'h5be00000;
      40413: inst = 32'h8c50000;
      40414: inst = 32'h24612800;
      40415: inst = 32'h10a0ffff;
      40416: inst = 32'hca0ffe3;
      40417: inst = 32'h24822800;
      40418: inst = 32'h10a00000;
      40419: inst = 32'hca00004;
      40420: inst = 32'h38632800;
      40421: inst = 32'h38842800;
      40422: inst = 32'h10a00000;
      40423: inst = 32'hca09deb;
      40424: inst = 32'h13e00001;
      40425: inst = 32'hfe0d96a;
      40426: inst = 32'h5be00000;
      40427: inst = 32'h8c50000;
      40428: inst = 32'h24612800;
      40429: inst = 32'h10a0ffff;
      40430: inst = 32'hca0ffe3;
      40431: inst = 32'h24822800;
      40432: inst = 32'h10a00000;
      40433: inst = 32'hca00004;
      40434: inst = 32'h38632800;
      40435: inst = 32'h38842800;
      40436: inst = 32'h10a00000;
      40437: inst = 32'hca09df9;
      40438: inst = 32'h13e00001;
      40439: inst = 32'hfe0d96a;
      40440: inst = 32'h5be00000;
      40441: inst = 32'h8c50000;
      40442: inst = 32'h24612800;
      40443: inst = 32'h10a0ffff;
      40444: inst = 32'hca0ffe3;
      40445: inst = 32'h24822800;
      40446: inst = 32'h10a00000;
      40447: inst = 32'hca00004;
      40448: inst = 32'h38632800;
      40449: inst = 32'h38842800;
      40450: inst = 32'h10a00000;
      40451: inst = 32'hca09e07;
      40452: inst = 32'h13e00001;
      40453: inst = 32'hfe0d96a;
      40454: inst = 32'h5be00000;
      40455: inst = 32'h8c50000;
      40456: inst = 32'h24612800;
      40457: inst = 32'h10a0ffff;
      40458: inst = 32'hca0ffe3;
      40459: inst = 32'h24822800;
      40460: inst = 32'h10a00000;
      40461: inst = 32'hca00004;
      40462: inst = 32'h38632800;
      40463: inst = 32'h38842800;
      40464: inst = 32'h10a00000;
      40465: inst = 32'hca09e15;
      40466: inst = 32'h13e00001;
      40467: inst = 32'hfe0d96a;
      40468: inst = 32'h5be00000;
      40469: inst = 32'h8c50000;
      40470: inst = 32'h24612800;
      40471: inst = 32'h10a0ffff;
      40472: inst = 32'hca0ffe3;
      40473: inst = 32'h24822800;
      40474: inst = 32'h10a00000;
      40475: inst = 32'hca00004;
      40476: inst = 32'h38632800;
      40477: inst = 32'h38842800;
      40478: inst = 32'h10a00000;
      40479: inst = 32'hca09e23;
      40480: inst = 32'h13e00001;
      40481: inst = 32'hfe0d96a;
      40482: inst = 32'h5be00000;
      40483: inst = 32'h8c50000;
      40484: inst = 32'h24612800;
      40485: inst = 32'h10a0ffff;
      40486: inst = 32'hca0ffe3;
      40487: inst = 32'h24822800;
      40488: inst = 32'h10a00000;
      40489: inst = 32'hca00004;
      40490: inst = 32'h38632800;
      40491: inst = 32'h38842800;
      40492: inst = 32'h10a00000;
      40493: inst = 32'hca09e31;
      40494: inst = 32'h13e00001;
      40495: inst = 32'hfe0d96a;
      40496: inst = 32'h5be00000;
      40497: inst = 32'h8c50000;
      40498: inst = 32'h24612800;
      40499: inst = 32'h10a0ffff;
      40500: inst = 32'hca0ffe3;
      40501: inst = 32'h24822800;
      40502: inst = 32'h10a00000;
      40503: inst = 32'hca00004;
      40504: inst = 32'h38632800;
      40505: inst = 32'h38842800;
      40506: inst = 32'h10a00000;
      40507: inst = 32'hca09e3f;
      40508: inst = 32'h13e00001;
      40509: inst = 32'hfe0d96a;
      40510: inst = 32'h5be00000;
      40511: inst = 32'h8c50000;
      40512: inst = 32'h24612800;
      40513: inst = 32'h10a0ffff;
      40514: inst = 32'hca0ffe3;
      40515: inst = 32'h24822800;
      40516: inst = 32'h10a00000;
      40517: inst = 32'hca00004;
      40518: inst = 32'h38632800;
      40519: inst = 32'h38842800;
      40520: inst = 32'h10a00000;
      40521: inst = 32'hca09e4d;
      40522: inst = 32'h13e00001;
      40523: inst = 32'hfe0d96a;
      40524: inst = 32'h5be00000;
      40525: inst = 32'h8c50000;
      40526: inst = 32'h24612800;
      40527: inst = 32'h10a0ffff;
      40528: inst = 32'hca0ffe3;
      40529: inst = 32'h24822800;
      40530: inst = 32'h10a00000;
      40531: inst = 32'hca00004;
      40532: inst = 32'h38632800;
      40533: inst = 32'h38842800;
      40534: inst = 32'h10a00000;
      40535: inst = 32'hca09e5b;
      40536: inst = 32'h13e00001;
      40537: inst = 32'hfe0d96a;
      40538: inst = 32'h5be00000;
      40539: inst = 32'h8c50000;
      40540: inst = 32'h24612800;
      40541: inst = 32'h10a0ffff;
      40542: inst = 32'hca0ffe3;
      40543: inst = 32'h24822800;
      40544: inst = 32'h10a00000;
      40545: inst = 32'hca00004;
      40546: inst = 32'h38632800;
      40547: inst = 32'h38842800;
      40548: inst = 32'h10a00000;
      40549: inst = 32'hca09e69;
      40550: inst = 32'h13e00001;
      40551: inst = 32'hfe0d96a;
      40552: inst = 32'h5be00000;
      40553: inst = 32'h8c50000;
      40554: inst = 32'h24612800;
      40555: inst = 32'h10a0ffff;
      40556: inst = 32'hca0ffe4;
      40557: inst = 32'h24822800;
      40558: inst = 32'h10a00000;
      40559: inst = 32'hca00004;
      40560: inst = 32'h38632800;
      40561: inst = 32'h38842800;
      40562: inst = 32'h10a00000;
      40563: inst = 32'hca09e77;
      40564: inst = 32'h13e00001;
      40565: inst = 32'hfe0d96a;
      40566: inst = 32'h5be00000;
      40567: inst = 32'h8c50000;
      40568: inst = 32'h24612800;
      40569: inst = 32'h10a0ffff;
      40570: inst = 32'hca0ffe4;
      40571: inst = 32'h24822800;
      40572: inst = 32'h10a00000;
      40573: inst = 32'hca00004;
      40574: inst = 32'h38632800;
      40575: inst = 32'h38842800;
      40576: inst = 32'h10a00000;
      40577: inst = 32'hca09e85;
      40578: inst = 32'h13e00001;
      40579: inst = 32'hfe0d96a;
      40580: inst = 32'h5be00000;
      40581: inst = 32'h8c50000;
      40582: inst = 32'h24612800;
      40583: inst = 32'h10a0ffff;
      40584: inst = 32'hca0ffe4;
      40585: inst = 32'h24822800;
      40586: inst = 32'h10a00000;
      40587: inst = 32'hca00004;
      40588: inst = 32'h38632800;
      40589: inst = 32'h38842800;
      40590: inst = 32'h10a00000;
      40591: inst = 32'hca09e93;
      40592: inst = 32'h13e00001;
      40593: inst = 32'hfe0d96a;
      40594: inst = 32'h5be00000;
      40595: inst = 32'h8c50000;
      40596: inst = 32'h24612800;
      40597: inst = 32'h10a0ffff;
      40598: inst = 32'hca0ffe4;
      40599: inst = 32'h24822800;
      40600: inst = 32'h10a00000;
      40601: inst = 32'hca00004;
      40602: inst = 32'h38632800;
      40603: inst = 32'h38842800;
      40604: inst = 32'h10a00000;
      40605: inst = 32'hca09ea1;
      40606: inst = 32'h13e00001;
      40607: inst = 32'hfe0d96a;
      40608: inst = 32'h5be00000;
      40609: inst = 32'h8c50000;
      40610: inst = 32'h24612800;
      40611: inst = 32'h10a0ffff;
      40612: inst = 32'hca0ffe4;
      40613: inst = 32'h24822800;
      40614: inst = 32'h10a00000;
      40615: inst = 32'hca00004;
      40616: inst = 32'h38632800;
      40617: inst = 32'h38842800;
      40618: inst = 32'h10a00000;
      40619: inst = 32'hca09eaf;
      40620: inst = 32'h13e00001;
      40621: inst = 32'hfe0d96a;
      40622: inst = 32'h5be00000;
      40623: inst = 32'h8c50000;
      40624: inst = 32'h24612800;
      40625: inst = 32'h10a0ffff;
      40626: inst = 32'hca0ffe4;
      40627: inst = 32'h24822800;
      40628: inst = 32'h10a00000;
      40629: inst = 32'hca00004;
      40630: inst = 32'h38632800;
      40631: inst = 32'h38842800;
      40632: inst = 32'h10a00000;
      40633: inst = 32'hca09ebd;
      40634: inst = 32'h13e00001;
      40635: inst = 32'hfe0d96a;
      40636: inst = 32'h5be00000;
      40637: inst = 32'h8c50000;
      40638: inst = 32'h24612800;
      40639: inst = 32'h10a0ffff;
      40640: inst = 32'hca0ffe4;
      40641: inst = 32'h24822800;
      40642: inst = 32'h10a00000;
      40643: inst = 32'hca00004;
      40644: inst = 32'h38632800;
      40645: inst = 32'h38842800;
      40646: inst = 32'h10a00000;
      40647: inst = 32'hca09ecb;
      40648: inst = 32'h13e00001;
      40649: inst = 32'hfe0d96a;
      40650: inst = 32'h5be00000;
      40651: inst = 32'h8c50000;
      40652: inst = 32'h24612800;
      40653: inst = 32'h10a0ffff;
      40654: inst = 32'hca0ffe4;
      40655: inst = 32'h24822800;
      40656: inst = 32'h10a00000;
      40657: inst = 32'hca00004;
      40658: inst = 32'h38632800;
      40659: inst = 32'h38842800;
      40660: inst = 32'h10a00000;
      40661: inst = 32'hca09ed9;
      40662: inst = 32'h13e00001;
      40663: inst = 32'hfe0d96a;
      40664: inst = 32'h5be00000;
      40665: inst = 32'h8c50000;
      40666: inst = 32'h24612800;
      40667: inst = 32'h10a0ffff;
      40668: inst = 32'hca0ffe4;
      40669: inst = 32'h24822800;
      40670: inst = 32'h10a00000;
      40671: inst = 32'hca00004;
      40672: inst = 32'h38632800;
      40673: inst = 32'h38842800;
      40674: inst = 32'h10a00000;
      40675: inst = 32'hca09ee7;
      40676: inst = 32'h13e00001;
      40677: inst = 32'hfe0d96a;
      40678: inst = 32'h5be00000;
      40679: inst = 32'h8c50000;
      40680: inst = 32'h24612800;
      40681: inst = 32'h10a0ffff;
      40682: inst = 32'hca0ffe4;
      40683: inst = 32'h24822800;
      40684: inst = 32'h10a00000;
      40685: inst = 32'hca00004;
      40686: inst = 32'h38632800;
      40687: inst = 32'h38842800;
      40688: inst = 32'h10a00000;
      40689: inst = 32'hca09ef5;
      40690: inst = 32'h13e00001;
      40691: inst = 32'hfe0d96a;
      40692: inst = 32'h5be00000;
      40693: inst = 32'h8c50000;
      40694: inst = 32'h24612800;
      40695: inst = 32'h10a0ffff;
      40696: inst = 32'hca0ffe4;
      40697: inst = 32'h24822800;
      40698: inst = 32'h10a00000;
      40699: inst = 32'hca00004;
      40700: inst = 32'h38632800;
      40701: inst = 32'h38842800;
      40702: inst = 32'h10a00000;
      40703: inst = 32'hca09f03;
      40704: inst = 32'h13e00001;
      40705: inst = 32'hfe0d96a;
      40706: inst = 32'h5be00000;
      40707: inst = 32'h8c50000;
      40708: inst = 32'h24612800;
      40709: inst = 32'h10a0ffff;
      40710: inst = 32'hca0ffe4;
      40711: inst = 32'h24822800;
      40712: inst = 32'h10a00000;
      40713: inst = 32'hca00004;
      40714: inst = 32'h38632800;
      40715: inst = 32'h38842800;
      40716: inst = 32'h10a00000;
      40717: inst = 32'hca09f11;
      40718: inst = 32'h13e00001;
      40719: inst = 32'hfe0d96a;
      40720: inst = 32'h5be00000;
      40721: inst = 32'h8c50000;
      40722: inst = 32'h24612800;
      40723: inst = 32'h10a0ffff;
      40724: inst = 32'hca0ffe4;
      40725: inst = 32'h24822800;
      40726: inst = 32'h10a00000;
      40727: inst = 32'hca00004;
      40728: inst = 32'h38632800;
      40729: inst = 32'h38842800;
      40730: inst = 32'h10a00000;
      40731: inst = 32'hca09f1f;
      40732: inst = 32'h13e00001;
      40733: inst = 32'hfe0d96a;
      40734: inst = 32'h5be00000;
      40735: inst = 32'h8c50000;
      40736: inst = 32'h24612800;
      40737: inst = 32'h10a0ffff;
      40738: inst = 32'hca0ffe4;
      40739: inst = 32'h24822800;
      40740: inst = 32'h10a00000;
      40741: inst = 32'hca00004;
      40742: inst = 32'h38632800;
      40743: inst = 32'h38842800;
      40744: inst = 32'h10a00000;
      40745: inst = 32'hca09f2d;
      40746: inst = 32'h13e00001;
      40747: inst = 32'hfe0d96a;
      40748: inst = 32'h5be00000;
      40749: inst = 32'h8c50000;
      40750: inst = 32'h24612800;
      40751: inst = 32'h10a0ffff;
      40752: inst = 32'hca0ffe4;
      40753: inst = 32'h24822800;
      40754: inst = 32'h10a00000;
      40755: inst = 32'hca00004;
      40756: inst = 32'h38632800;
      40757: inst = 32'h38842800;
      40758: inst = 32'h10a00000;
      40759: inst = 32'hca09f3b;
      40760: inst = 32'h13e00001;
      40761: inst = 32'hfe0d96a;
      40762: inst = 32'h5be00000;
      40763: inst = 32'h8c50000;
      40764: inst = 32'h24612800;
      40765: inst = 32'h10a0ffff;
      40766: inst = 32'hca0ffe4;
      40767: inst = 32'h24822800;
      40768: inst = 32'h10a00000;
      40769: inst = 32'hca00004;
      40770: inst = 32'h38632800;
      40771: inst = 32'h38842800;
      40772: inst = 32'h10a00000;
      40773: inst = 32'hca09f49;
      40774: inst = 32'h13e00001;
      40775: inst = 32'hfe0d96a;
      40776: inst = 32'h5be00000;
      40777: inst = 32'h8c50000;
      40778: inst = 32'h24612800;
      40779: inst = 32'h10a0ffff;
      40780: inst = 32'hca0ffe4;
      40781: inst = 32'h24822800;
      40782: inst = 32'h10a00000;
      40783: inst = 32'hca00004;
      40784: inst = 32'h38632800;
      40785: inst = 32'h38842800;
      40786: inst = 32'h10a00000;
      40787: inst = 32'hca09f57;
      40788: inst = 32'h13e00001;
      40789: inst = 32'hfe0d96a;
      40790: inst = 32'h5be00000;
      40791: inst = 32'h8c50000;
      40792: inst = 32'h24612800;
      40793: inst = 32'h10a0ffff;
      40794: inst = 32'hca0ffe4;
      40795: inst = 32'h24822800;
      40796: inst = 32'h10a00000;
      40797: inst = 32'hca00004;
      40798: inst = 32'h38632800;
      40799: inst = 32'h38842800;
      40800: inst = 32'h10a00000;
      40801: inst = 32'hca09f65;
      40802: inst = 32'h13e00001;
      40803: inst = 32'hfe0d96a;
      40804: inst = 32'h5be00000;
      40805: inst = 32'h8c50000;
      40806: inst = 32'h24612800;
      40807: inst = 32'h10a0ffff;
      40808: inst = 32'hca0ffe4;
      40809: inst = 32'h24822800;
      40810: inst = 32'h10a00000;
      40811: inst = 32'hca00004;
      40812: inst = 32'h38632800;
      40813: inst = 32'h38842800;
      40814: inst = 32'h10a00000;
      40815: inst = 32'hca09f73;
      40816: inst = 32'h13e00001;
      40817: inst = 32'hfe0d96a;
      40818: inst = 32'h5be00000;
      40819: inst = 32'h8c50000;
      40820: inst = 32'h24612800;
      40821: inst = 32'h10a0ffff;
      40822: inst = 32'hca0ffe4;
      40823: inst = 32'h24822800;
      40824: inst = 32'h10a00000;
      40825: inst = 32'hca00004;
      40826: inst = 32'h38632800;
      40827: inst = 32'h38842800;
      40828: inst = 32'h10a00000;
      40829: inst = 32'hca09f81;
      40830: inst = 32'h13e00001;
      40831: inst = 32'hfe0d96a;
      40832: inst = 32'h5be00000;
      40833: inst = 32'h8c50000;
      40834: inst = 32'h24612800;
      40835: inst = 32'h10a0ffff;
      40836: inst = 32'hca0ffe4;
      40837: inst = 32'h24822800;
      40838: inst = 32'h10a00000;
      40839: inst = 32'hca00004;
      40840: inst = 32'h38632800;
      40841: inst = 32'h38842800;
      40842: inst = 32'h10a00000;
      40843: inst = 32'hca09f8f;
      40844: inst = 32'h13e00001;
      40845: inst = 32'hfe0d96a;
      40846: inst = 32'h5be00000;
      40847: inst = 32'h8c50000;
      40848: inst = 32'h24612800;
      40849: inst = 32'h10a0ffff;
      40850: inst = 32'hca0ffe4;
      40851: inst = 32'h24822800;
      40852: inst = 32'h10a00000;
      40853: inst = 32'hca00004;
      40854: inst = 32'h38632800;
      40855: inst = 32'h38842800;
      40856: inst = 32'h10a00000;
      40857: inst = 32'hca09f9d;
      40858: inst = 32'h13e00001;
      40859: inst = 32'hfe0d96a;
      40860: inst = 32'h5be00000;
      40861: inst = 32'h8c50000;
      40862: inst = 32'h24612800;
      40863: inst = 32'h10a0ffff;
      40864: inst = 32'hca0ffe4;
      40865: inst = 32'h24822800;
      40866: inst = 32'h10a00000;
      40867: inst = 32'hca00004;
      40868: inst = 32'h38632800;
      40869: inst = 32'h38842800;
      40870: inst = 32'h10a00000;
      40871: inst = 32'hca09fab;
      40872: inst = 32'h13e00001;
      40873: inst = 32'hfe0d96a;
      40874: inst = 32'h5be00000;
      40875: inst = 32'h8c50000;
      40876: inst = 32'h24612800;
      40877: inst = 32'h10a0ffff;
      40878: inst = 32'hca0ffe4;
      40879: inst = 32'h24822800;
      40880: inst = 32'h10a00000;
      40881: inst = 32'hca00004;
      40882: inst = 32'h38632800;
      40883: inst = 32'h38842800;
      40884: inst = 32'h10a00000;
      40885: inst = 32'hca09fb9;
      40886: inst = 32'h13e00001;
      40887: inst = 32'hfe0d96a;
      40888: inst = 32'h5be00000;
      40889: inst = 32'h8c50000;
      40890: inst = 32'h24612800;
      40891: inst = 32'h10a0ffff;
      40892: inst = 32'hca0ffe4;
      40893: inst = 32'h24822800;
      40894: inst = 32'h10a00000;
      40895: inst = 32'hca00004;
      40896: inst = 32'h38632800;
      40897: inst = 32'h38842800;
      40898: inst = 32'h10a00000;
      40899: inst = 32'hca09fc7;
      40900: inst = 32'h13e00001;
      40901: inst = 32'hfe0d96a;
      40902: inst = 32'h5be00000;
      40903: inst = 32'h8c50000;
      40904: inst = 32'h24612800;
      40905: inst = 32'h10a0ffff;
      40906: inst = 32'hca0ffe4;
      40907: inst = 32'h24822800;
      40908: inst = 32'h10a00000;
      40909: inst = 32'hca00004;
      40910: inst = 32'h38632800;
      40911: inst = 32'h38842800;
      40912: inst = 32'h10a00000;
      40913: inst = 32'hca09fd5;
      40914: inst = 32'h13e00001;
      40915: inst = 32'hfe0d96a;
      40916: inst = 32'h5be00000;
      40917: inst = 32'h8c50000;
      40918: inst = 32'h24612800;
      40919: inst = 32'h10a0ffff;
      40920: inst = 32'hca0ffe4;
      40921: inst = 32'h24822800;
      40922: inst = 32'h10a00000;
      40923: inst = 32'hca00004;
      40924: inst = 32'h38632800;
      40925: inst = 32'h38842800;
      40926: inst = 32'h10a00000;
      40927: inst = 32'hca09fe3;
      40928: inst = 32'h13e00001;
      40929: inst = 32'hfe0d96a;
      40930: inst = 32'h5be00000;
      40931: inst = 32'h8c50000;
      40932: inst = 32'h24612800;
      40933: inst = 32'h10a0ffff;
      40934: inst = 32'hca0ffe4;
      40935: inst = 32'h24822800;
      40936: inst = 32'h10a00000;
      40937: inst = 32'hca00004;
      40938: inst = 32'h38632800;
      40939: inst = 32'h38842800;
      40940: inst = 32'h10a00000;
      40941: inst = 32'hca09ff1;
      40942: inst = 32'h13e00001;
      40943: inst = 32'hfe0d96a;
      40944: inst = 32'h5be00000;
      40945: inst = 32'h8c50000;
      40946: inst = 32'h24612800;
      40947: inst = 32'h10a0ffff;
      40948: inst = 32'hca0ffe4;
      40949: inst = 32'h24822800;
      40950: inst = 32'h10a00000;
      40951: inst = 32'hca00004;
      40952: inst = 32'h38632800;
      40953: inst = 32'h38842800;
      40954: inst = 32'h10a00000;
      40955: inst = 32'hca09fff;
      40956: inst = 32'h13e00001;
      40957: inst = 32'hfe0d96a;
      40958: inst = 32'h5be00000;
      40959: inst = 32'h8c50000;
      40960: inst = 32'h24612800;
      40961: inst = 32'h10a0ffff;
      40962: inst = 32'hca0ffe4;
      40963: inst = 32'h24822800;
      40964: inst = 32'h10a00000;
      40965: inst = 32'hca00004;
      40966: inst = 32'h38632800;
      40967: inst = 32'h38842800;
      40968: inst = 32'h10a00000;
      40969: inst = 32'hca0a00d;
      40970: inst = 32'h13e00001;
      40971: inst = 32'hfe0d96a;
      40972: inst = 32'h5be00000;
      40973: inst = 32'h8c50000;
      40974: inst = 32'h24612800;
      40975: inst = 32'h10a0ffff;
      40976: inst = 32'hca0ffe4;
      40977: inst = 32'h24822800;
      40978: inst = 32'h10a00000;
      40979: inst = 32'hca00004;
      40980: inst = 32'h38632800;
      40981: inst = 32'h38842800;
      40982: inst = 32'h10a00000;
      40983: inst = 32'hca0a01b;
      40984: inst = 32'h13e00001;
      40985: inst = 32'hfe0d96a;
      40986: inst = 32'h5be00000;
      40987: inst = 32'h8c50000;
      40988: inst = 32'h24612800;
      40989: inst = 32'h10a0ffff;
      40990: inst = 32'hca0ffe4;
      40991: inst = 32'h24822800;
      40992: inst = 32'h10a00000;
      40993: inst = 32'hca00004;
      40994: inst = 32'h38632800;
      40995: inst = 32'h38842800;
      40996: inst = 32'h10a00000;
      40997: inst = 32'hca0a029;
      40998: inst = 32'h13e00001;
      40999: inst = 32'hfe0d96a;
      41000: inst = 32'h5be00000;
      41001: inst = 32'h8c50000;
      41002: inst = 32'h24612800;
      41003: inst = 32'h10a0ffff;
      41004: inst = 32'hca0ffe4;
      41005: inst = 32'h24822800;
      41006: inst = 32'h10a00000;
      41007: inst = 32'hca00004;
      41008: inst = 32'h38632800;
      41009: inst = 32'h38842800;
      41010: inst = 32'h10a00000;
      41011: inst = 32'hca0a037;
      41012: inst = 32'h13e00001;
      41013: inst = 32'hfe0d96a;
      41014: inst = 32'h5be00000;
      41015: inst = 32'h8c50000;
      41016: inst = 32'h24612800;
      41017: inst = 32'h10a0ffff;
      41018: inst = 32'hca0ffe4;
      41019: inst = 32'h24822800;
      41020: inst = 32'h10a00000;
      41021: inst = 32'hca00004;
      41022: inst = 32'h38632800;
      41023: inst = 32'h38842800;
      41024: inst = 32'h10a00000;
      41025: inst = 32'hca0a045;
      41026: inst = 32'h13e00001;
      41027: inst = 32'hfe0d96a;
      41028: inst = 32'h5be00000;
      41029: inst = 32'h8c50000;
      41030: inst = 32'h24612800;
      41031: inst = 32'h10a0ffff;
      41032: inst = 32'hca0ffe4;
      41033: inst = 32'h24822800;
      41034: inst = 32'h10a00000;
      41035: inst = 32'hca00004;
      41036: inst = 32'h38632800;
      41037: inst = 32'h38842800;
      41038: inst = 32'h10a00000;
      41039: inst = 32'hca0a053;
      41040: inst = 32'h13e00001;
      41041: inst = 32'hfe0d96a;
      41042: inst = 32'h5be00000;
      41043: inst = 32'h8c50000;
      41044: inst = 32'h24612800;
      41045: inst = 32'h10a0ffff;
      41046: inst = 32'hca0ffe4;
      41047: inst = 32'h24822800;
      41048: inst = 32'h10a00000;
      41049: inst = 32'hca00004;
      41050: inst = 32'h38632800;
      41051: inst = 32'h38842800;
      41052: inst = 32'h10a00000;
      41053: inst = 32'hca0a061;
      41054: inst = 32'h13e00001;
      41055: inst = 32'hfe0d96a;
      41056: inst = 32'h5be00000;
      41057: inst = 32'h8c50000;
      41058: inst = 32'h24612800;
      41059: inst = 32'h10a0ffff;
      41060: inst = 32'hca0ffe4;
      41061: inst = 32'h24822800;
      41062: inst = 32'h10a00000;
      41063: inst = 32'hca00004;
      41064: inst = 32'h38632800;
      41065: inst = 32'h38842800;
      41066: inst = 32'h10a00000;
      41067: inst = 32'hca0a06f;
      41068: inst = 32'h13e00001;
      41069: inst = 32'hfe0d96a;
      41070: inst = 32'h5be00000;
      41071: inst = 32'h8c50000;
      41072: inst = 32'h24612800;
      41073: inst = 32'h10a0ffff;
      41074: inst = 32'hca0ffe4;
      41075: inst = 32'h24822800;
      41076: inst = 32'h10a00000;
      41077: inst = 32'hca00004;
      41078: inst = 32'h38632800;
      41079: inst = 32'h38842800;
      41080: inst = 32'h10a00000;
      41081: inst = 32'hca0a07d;
      41082: inst = 32'h13e00001;
      41083: inst = 32'hfe0d96a;
      41084: inst = 32'h5be00000;
      41085: inst = 32'h8c50000;
      41086: inst = 32'h24612800;
      41087: inst = 32'h10a0ffff;
      41088: inst = 32'hca0ffe4;
      41089: inst = 32'h24822800;
      41090: inst = 32'h10a00000;
      41091: inst = 32'hca00004;
      41092: inst = 32'h38632800;
      41093: inst = 32'h38842800;
      41094: inst = 32'h10a00000;
      41095: inst = 32'hca0a08b;
      41096: inst = 32'h13e00001;
      41097: inst = 32'hfe0d96a;
      41098: inst = 32'h5be00000;
      41099: inst = 32'h8c50000;
      41100: inst = 32'h24612800;
      41101: inst = 32'h10a0ffff;
      41102: inst = 32'hca0ffe4;
      41103: inst = 32'h24822800;
      41104: inst = 32'h10a00000;
      41105: inst = 32'hca00004;
      41106: inst = 32'h38632800;
      41107: inst = 32'h38842800;
      41108: inst = 32'h10a00000;
      41109: inst = 32'hca0a099;
      41110: inst = 32'h13e00001;
      41111: inst = 32'hfe0d96a;
      41112: inst = 32'h5be00000;
      41113: inst = 32'h8c50000;
      41114: inst = 32'h24612800;
      41115: inst = 32'h10a0ffff;
      41116: inst = 32'hca0ffe4;
      41117: inst = 32'h24822800;
      41118: inst = 32'h10a00000;
      41119: inst = 32'hca00004;
      41120: inst = 32'h38632800;
      41121: inst = 32'h38842800;
      41122: inst = 32'h10a00000;
      41123: inst = 32'hca0a0a7;
      41124: inst = 32'h13e00001;
      41125: inst = 32'hfe0d96a;
      41126: inst = 32'h5be00000;
      41127: inst = 32'h8c50000;
      41128: inst = 32'h24612800;
      41129: inst = 32'h10a0ffff;
      41130: inst = 32'hca0ffe4;
      41131: inst = 32'h24822800;
      41132: inst = 32'h10a00000;
      41133: inst = 32'hca00004;
      41134: inst = 32'h38632800;
      41135: inst = 32'h38842800;
      41136: inst = 32'h10a00000;
      41137: inst = 32'hca0a0b5;
      41138: inst = 32'h13e00001;
      41139: inst = 32'hfe0d96a;
      41140: inst = 32'h5be00000;
      41141: inst = 32'h8c50000;
      41142: inst = 32'h24612800;
      41143: inst = 32'h10a0ffff;
      41144: inst = 32'hca0ffe4;
      41145: inst = 32'h24822800;
      41146: inst = 32'h10a00000;
      41147: inst = 32'hca00004;
      41148: inst = 32'h38632800;
      41149: inst = 32'h38842800;
      41150: inst = 32'h10a00000;
      41151: inst = 32'hca0a0c3;
      41152: inst = 32'h13e00001;
      41153: inst = 32'hfe0d96a;
      41154: inst = 32'h5be00000;
      41155: inst = 32'h8c50000;
      41156: inst = 32'h24612800;
      41157: inst = 32'h10a0ffff;
      41158: inst = 32'hca0ffe4;
      41159: inst = 32'h24822800;
      41160: inst = 32'h10a00000;
      41161: inst = 32'hca00004;
      41162: inst = 32'h38632800;
      41163: inst = 32'h38842800;
      41164: inst = 32'h10a00000;
      41165: inst = 32'hca0a0d1;
      41166: inst = 32'h13e00001;
      41167: inst = 32'hfe0d96a;
      41168: inst = 32'h5be00000;
      41169: inst = 32'h8c50000;
      41170: inst = 32'h24612800;
      41171: inst = 32'h10a0ffff;
      41172: inst = 32'hca0ffe4;
      41173: inst = 32'h24822800;
      41174: inst = 32'h10a00000;
      41175: inst = 32'hca00004;
      41176: inst = 32'h38632800;
      41177: inst = 32'h38842800;
      41178: inst = 32'h10a00000;
      41179: inst = 32'hca0a0df;
      41180: inst = 32'h13e00001;
      41181: inst = 32'hfe0d96a;
      41182: inst = 32'h5be00000;
      41183: inst = 32'h8c50000;
      41184: inst = 32'h24612800;
      41185: inst = 32'h10a0ffff;
      41186: inst = 32'hca0ffe4;
      41187: inst = 32'h24822800;
      41188: inst = 32'h10a00000;
      41189: inst = 32'hca00004;
      41190: inst = 32'h38632800;
      41191: inst = 32'h38842800;
      41192: inst = 32'h10a00000;
      41193: inst = 32'hca0a0ed;
      41194: inst = 32'h13e00001;
      41195: inst = 32'hfe0d96a;
      41196: inst = 32'h5be00000;
      41197: inst = 32'h8c50000;
      41198: inst = 32'h24612800;
      41199: inst = 32'h10a0ffff;
      41200: inst = 32'hca0ffe4;
      41201: inst = 32'h24822800;
      41202: inst = 32'h10a00000;
      41203: inst = 32'hca00004;
      41204: inst = 32'h38632800;
      41205: inst = 32'h38842800;
      41206: inst = 32'h10a00000;
      41207: inst = 32'hca0a0fb;
      41208: inst = 32'h13e00001;
      41209: inst = 32'hfe0d96a;
      41210: inst = 32'h5be00000;
      41211: inst = 32'h8c50000;
      41212: inst = 32'h24612800;
      41213: inst = 32'h10a0ffff;
      41214: inst = 32'hca0ffe4;
      41215: inst = 32'h24822800;
      41216: inst = 32'h10a00000;
      41217: inst = 32'hca00004;
      41218: inst = 32'h38632800;
      41219: inst = 32'h38842800;
      41220: inst = 32'h10a00000;
      41221: inst = 32'hca0a109;
      41222: inst = 32'h13e00001;
      41223: inst = 32'hfe0d96a;
      41224: inst = 32'h5be00000;
      41225: inst = 32'h8c50000;
      41226: inst = 32'h24612800;
      41227: inst = 32'h10a0ffff;
      41228: inst = 32'hca0ffe4;
      41229: inst = 32'h24822800;
      41230: inst = 32'h10a00000;
      41231: inst = 32'hca00004;
      41232: inst = 32'h38632800;
      41233: inst = 32'h38842800;
      41234: inst = 32'h10a00000;
      41235: inst = 32'hca0a117;
      41236: inst = 32'h13e00001;
      41237: inst = 32'hfe0d96a;
      41238: inst = 32'h5be00000;
      41239: inst = 32'h8c50000;
      41240: inst = 32'h24612800;
      41241: inst = 32'h10a0ffff;
      41242: inst = 32'hca0ffe4;
      41243: inst = 32'h24822800;
      41244: inst = 32'h10a00000;
      41245: inst = 32'hca00004;
      41246: inst = 32'h38632800;
      41247: inst = 32'h38842800;
      41248: inst = 32'h10a00000;
      41249: inst = 32'hca0a125;
      41250: inst = 32'h13e00001;
      41251: inst = 32'hfe0d96a;
      41252: inst = 32'h5be00000;
      41253: inst = 32'h8c50000;
      41254: inst = 32'h24612800;
      41255: inst = 32'h10a0ffff;
      41256: inst = 32'hca0ffe4;
      41257: inst = 32'h24822800;
      41258: inst = 32'h10a00000;
      41259: inst = 32'hca00004;
      41260: inst = 32'h38632800;
      41261: inst = 32'h38842800;
      41262: inst = 32'h10a00000;
      41263: inst = 32'hca0a133;
      41264: inst = 32'h13e00001;
      41265: inst = 32'hfe0d96a;
      41266: inst = 32'h5be00000;
      41267: inst = 32'h8c50000;
      41268: inst = 32'h24612800;
      41269: inst = 32'h10a0ffff;
      41270: inst = 32'hca0ffe4;
      41271: inst = 32'h24822800;
      41272: inst = 32'h10a00000;
      41273: inst = 32'hca00004;
      41274: inst = 32'h38632800;
      41275: inst = 32'h38842800;
      41276: inst = 32'h10a00000;
      41277: inst = 32'hca0a141;
      41278: inst = 32'h13e00001;
      41279: inst = 32'hfe0d96a;
      41280: inst = 32'h5be00000;
      41281: inst = 32'h8c50000;
      41282: inst = 32'h24612800;
      41283: inst = 32'h10a0ffff;
      41284: inst = 32'hca0ffe4;
      41285: inst = 32'h24822800;
      41286: inst = 32'h10a00000;
      41287: inst = 32'hca00004;
      41288: inst = 32'h38632800;
      41289: inst = 32'h38842800;
      41290: inst = 32'h10a00000;
      41291: inst = 32'hca0a14f;
      41292: inst = 32'h13e00001;
      41293: inst = 32'hfe0d96a;
      41294: inst = 32'h5be00000;
      41295: inst = 32'h8c50000;
      41296: inst = 32'h24612800;
      41297: inst = 32'h10a0ffff;
      41298: inst = 32'hca0ffe4;
      41299: inst = 32'h24822800;
      41300: inst = 32'h10a00000;
      41301: inst = 32'hca00004;
      41302: inst = 32'h38632800;
      41303: inst = 32'h38842800;
      41304: inst = 32'h10a00000;
      41305: inst = 32'hca0a15d;
      41306: inst = 32'h13e00001;
      41307: inst = 32'hfe0d96a;
      41308: inst = 32'h5be00000;
      41309: inst = 32'h8c50000;
      41310: inst = 32'h24612800;
      41311: inst = 32'h10a0ffff;
      41312: inst = 32'hca0ffe4;
      41313: inst = 32'h24822800;
      41314: inst = 32'h10a00000;
      41315: inst = 32'hca00004;
      41316: inst = 32'h38632800;
      41317: inst = 32'h38842800;
      41318: inst = 32'h10a00000;
      41319: inst = 32'hca0a16b;
      41320: inst = 32'h13e00001;
      41321: inst = 32'hfe0d96a;
      41322: inst = 32'h5be00000;
      41323: inst = 32'h8c50000;
      41324: inst = 32'h24612800;
      41325: inst = 32'h10a0ffff;
      41326: inst = 32'hca0ffe4;
      41327: inst = 32'h24822800;
      41328: inst = 32'h10a00000;
      41329: inst = 32'hca00004;
      41330: inst = 32'h38632800;
      41331: inst = 32'h38842800;
      41332: inst = 32'h10a00000;
      41333: inst = 32'hca0a179;
      41334: inst = 32'h13e00001;
      41335: inst = 32'hfe0d96a;
      41336: inst = 32'h5be00000;
      41337: inst = 32'h8c50000;
      41338: inst = 32'h24612800;
      41339: inst = 32'h10a0ffff;
      41340: inst = 32'hca0ffe4;
      41341: inst = 32'h24822800;
      41342: inst = 32'h10a00000;
      41343: inst = 32'hca00004;
      41344: inst = 32'h38632800;
      41345: inst = 32'h38842800;
      41346: inst = 32'h10a00000;
      41347: inst = 32'hca0a187;
      41348: inst = 32'h13e00001;
      41349: inst = 32'hfe0d96a;
      41350: inst = 32'h5be00000;
      41351: inst = 32'h8c50000;
      41352: inst = 32'h24612800;
      41353: inst = 32'h10a0ffff;
      41354: inst = 32'hca0ffe4;
      41355: inst = 32'h24822800;
      41356: inst = 32'h10a00000;
      41357: inst = 32'hca00004;
      41358: inst = 32'h38632800;
      41359: inst = 32'h38842800;
      41360: inst = 32'h10a00000;
      41361: inst = 32'hca0a195;
      41362: inst = 32'h13e00001;
      41363: inst = 32'hfe0d96a;
      41364: inst = 32'h5be00000;
      41365: inst = 32'h8c50000;
      41366: inst = 32'h24612800;
      41367: inst = 32'h10a0ffff;
      41368: inst = 32'hca0ffe4;
      41369: inst = 32'h24822800;
      41370: inst = 32'h10a00000;
      41371: inst = 32'hca00004;
      41372: inst = 32'h38632800;
      41373: inst = 32'h38842800;
      41374: inst = 32'h10a00000;
      41375: inst = 32'hca0a1a3;
      41376: inst = 32'h13e00001;
      41377: inst = 32'hfe0d96a;
      41378: inst = 32'h5be00000;
      41379: inst = 32'h8c50000;
      41380: inst = 32'h24612800;
      41381: inst = 32'h10a0ffff;
      41382: inst = 32'hca0ffe4;
      41383: inst = 32'h24822800;
      41384: inst = 32'h10a00000;
      41385: inst = 32'hca00004;
      41386: inst = 32'h38632800;
      41387: inst = 32'h38842800;
      41388: inst = 32'h10a00000;
      41389: inst = 32'hca0a1b1;
      41390: inst = 32'h13e00001;
      41391: inst = 32'hfe0d96a;
      41392: inst = 32'h5be00000;
      41393: inst = 32'h8c50000;
      41394: inst = 32'h24612800;
      41395: inst = 32'h10a0ffff;
      41396: inst = 32'hca0ffe4;
      41397: inst = 32'h24822800;
      41398: inst = 32'h10a00000;
      41399: inst = 32'hca00004;
      41400: inst = 32'h38632800;
      41401: inst = 32'h38842800;
      41402: inst = 32'h10a00000;
      41403: inst = 32'hca0a1bf;
      41404: inst = 32'h13e00001;
      41405: inst = 32'hfe0d96a;
      41406: inst = 32'h5be00000;
      41407: inst = 32'h8c50000;
      41408: inst = 32'h24612800;
      41409: inst = 32'h10a0ffff;
      41410: inst = 32'hca0ffe4;
      41411: inst = 32'h24822800;
      41412: inst = 32'h10a00000;
      41413: inst = 32'hca00004;
      41414: inst = 32'h38632800;
      41415: inst = 32'h38842800;
      41416: inst = 32'h10a00000;
      41417: inst = 32'hca0a1cd;
      41418: inst = 32'h13e00001;
      41419: inst = 32'hfe0d96a;
      41420: inst = 32'h5be00000;
      41421: inst = 32'h8c50000;
      41422: inst = 32'h24612800;
      41423: inst = 32'h10a0ffff;
      41424: inst = 32'hca0ffe4;
      41425: inst = 32'h24822800;
      41426: inst = 32'h10a00000;
      41427: inst = 32'hca00004;
      41428: inst = 32'h38632800;
      41429: inst = 32'h38842800;
      41430: inst = 32'h10a00000;
      41431: inst = 32'hca0a1db;
      41432: inst = 32'h13e00001;
      41433: inst = 32'hfe0d96a;
      41434: inst = 32'h5be00000;
      41435: inst = 32'h8c50000;
      41436: inst = 32'h24612800;
      41437: inst = 32'h10a0ffff;
      41438: inst = 32'hca0ffe4;
      41439: inst = 32'h24822800;
      41440: inst = 32'h10a00000;
      41441: inst = 32'hca00004;
      41442: inst = 32'h38632800;
      41443: inst = 32'h38842800;
      41444: inst = 32'h10a00000;
      41445: inst = 32'hca0a1e9;
      41446: inst = 32'h13e00001;
      41447: inst = 32'hfe0d96a;
      41448: inst = 32'h5be00000;
      41449: inst = 32'h8c50000;
      41450: inst = 32'h24612800;
      41451: inst = 32'h10a0ffff;
      41452: inst = 32'hca0ffe4;
      41453: inst = 32'h24822800;
      41454: inst = 32'h10a00000;
      41455: inst = 32'hca00004;
      41456: inst = 32'h38632800;
      41457: inst = 32'h38842800;
      41458: inst = 32'h10a00000;
      41459: inst = 32'hca0a1f7;
      41460: inst = 32'h13e00001;
      41461: inst = 32'hfe0d96a;
      41462: inst = 32'h5be00000;
      41463: inst = 32'h8c50000;
      41464: inst = 32'h24612800;
      41465: inst = 32'h10a0ffff;
      41466: inst = 32'hca0ffe4;
      41467: inst = 32'h24822800;
      41468: inst = 32'h10a00000;
      41469: inst = 32'hca00004;
      41470: inst = 32'h38632800;
      41471: inst = 32'h38842800;
      41472: inst = 32'h10a00000;
      41473: inst = 32'hca0a205;
      41474: inst = 32'h13e00001;
      41475: inst = 32'hfe0d96a;
      41476: inst = 32'h5be00000;
      41477: inst = 32'h8c50000;
      41478: inst = 32'h24612800;
      41479: inst = 32'h10a0ffff;
      41480: inst = 32'hca0ffe4;
      41481: inst = 32'h24822800;
      41482: inst = 32'h10a00000;
      41483: inst = 32'hca00004;
      41484: inst = 32'h38632800;
      41485: inst = 32'h38842800;
      41486: inst = 32'h10a00000;
      41487: inst = 32'hca0a213;
      41488: inst = 32'h13e00001;
      41489: inst = 32'hfe0d96a;
      41490: inst = 32'h5be00000;
      41491: inst = 32'h8c50000;
      41492: inst = 32'h24612800;
      41493: inst = 32'h10a0ffff;
      41494: inst = 32'hca0ffe4;
      41495: inst = 32'h24822800;
      41496: inst = 32'h10a00000;
      41497: inst = 32'hca00004;
      41498: inst = 32'h38632800;
      41499: inst = 32'h38842800;
      41500: inst = 32'h10a00000;
      41501: inst = 32'hca0a221;
      41502: inst = 32'h13e00001;
      41503: inst = 32'hfe0d96a;
      41504: inst = 32'h5be00000;
      41505: inst = 32'h8c50000;
      41506: inst = 32'h24612800;
      41507: inst = 32'h10a0ffff;
      41508: inst = 32'hca0ffe4;
      41509: inst = 32'h24822800;
      41510: inst = 32'h10a00000;
      41511: inst = 32'hca00004;
      41512: inst = 32'h38632800;
      41513: inst = 32'h38842800;
      41514: inst = 32'h10a00000;
      41515: inst = 32'hca0a22f;
      41516: inst = 32'h13e00001;
      41517: inst = 32'hfe0d96a;
      41518: inst = 32'h5be00000;
      41519: inst = 32'h8c50000;
      41520: inst = 32'h24612800;
      41521: inst = 32'h10a0ffff;
      41522: inst = 32'hca0ffe4;
      41523: inst = 32'h24822800;
      41524: inst = 32'h10a00000;
      41525: inst = 32'hca00004;
      41526: inst = 32'h38632800;
      41527: inst = 32'h38842800;
      41528: inst = 32'h10a00000;
      41529: inst = 32'hca0a23d;
      41530: inst = 32'h13e00001;
      41531: inst = 32'hfe0d96a;
      41532: inst = 32'h5be00000;
      41533: inst = 32'h8c50000;
      41534: inst = 32'h24612800;
      41535: inst = 32'h10a0ffff;
      41536: inst = 32'hca0ffe4;
      41537: inst = 32'h24822800;
      41538: inst = 32'h10a00000;
      41539: inst = 32'hca00004;
      41540: inst = 32'h38632800;
      41541: inst = 32'h38842800;
      41542: inst = 32'h10a00000;
      41543: inst = 32'hca0a24b;
      41544: inst = 32'h13e00001;
      41545: inst = 32'hfe0d96a;
      41546: inst = 32'h5be00000;
      41547: inst = 32'h8c50000;
      41548: inst = 32'h24612800;
      41549: inst = 32'h10a0ffff;
      41550: inst = 32'hca0ffe4;
      41551: inst = 32'h24822800;
      41552: inst = 32'h10a00000;
      41553: inst = 32'hca00004;
      41554: inst = 32'h38632800;
      41555: inst = 32'h38842800;
      41556: inst = 32'h10a00000;
      41557: inst = 32'hca0a259;
      41558: inst = 32'h13e00001;
      41559: inst = 32'hfe0d96a;
      41560: inst = 32'h5be00000;
      41561: inst = 32'h8c50000;
      41562: inst = 32'h24612800;
      41563: inst = 32'h10a0ffff;
      41564: inst = 32'hca0ffe4;
      41565: inst = 32'h24822800;
      41566: inst = 32'h10a00000;
      41567: inst = 32'hca00004;
      41568: inst = 32'h38632800;
      41569: inst = 32'h38842800;
      41570: inst = 32'h10a00000;
      41571: inst = 32'hca0a267;
      41572: inst = 32'h13e00001;
      41573: inst = 32'hfe0d96a;
      41574: inst = 32'h5be00000;
      41575: inst = 32'h8c50000;
      41576: inst = 32'h24612800;
      41577: inst = 32'h10a0ffff;
      41578: inst = 32'hca0ffe4;
      41579: inst = 32'h24822800;
      41580: inst = 32'h10a00000;
      41581: inst = 32'hca00004;
      41582: inst = 32'h38632800;
      41583: inst = 32'h38842800;
      41584: inst = 32'h10a00000;
      41585: inst = 32'hca0a275;
      41586: inst = 32'h13e00001;
      41587: inst = 32'hfe0d96a;
      41588: inst = 32'h5be00000;
      41589: inst = 32'h8c50000;
      41590: inst = 32'h24612800;
      41591: inst = 32'h10a0ffff;
      41592: inst = 32'hca0ffe4;
      41593: inst = 32'h24822800;
      41594: inst = 32'h10a00000;
      41595: inst = 32'hca00004;
      41596: inst = 32'h38632800;
      41597: inst = 32'h38842800;
      41598: inst = 32'h10a00000;
      41599: inst = 32'hca0a283;
      41600: inst = 32'h13e00001;
      41601: inst = 32'hfe0d96a;
      41602: inst = 32'h5be00000;
      41603: inst = 32'h8c50000;
      41604: inst = 32'h24612800;
      41605: inst = 32'h10a0ffff;
      41606: inst = 32'hca0ffe4;
      41607: inst = 32'h24822800;
      41608: inst = 32'h10a00000;
      41609: inst = 32'hca00004;
      41610: inst = 32'h38632800;
      41611: inst = 32'h38842800;
      41612: inst = 32'h10a00000;
      41613: inst = 32'hca0a291;
      41614: inst = 32'h13e00001;
      41615: inst = 32'hfe0d96a;
      41616: inst = 32'h5be00000;
      41617: inst = 32'h8c50000;
      41618: inst = 32'h24612800;
      41619: inst = 32'h10a0ffff;
      41620: inst = 32'hca0ffe4;
      41621: inst = 32'h24822800;
      41622: inst = 32'h10a00000;
      41623: inst = 32'hca00004;
      41624: inst = 32'h38632800;
      41625: inst = 32'h38842800;
      41626: inst = 32'h10a00000;
      41627: inst = 32'hca0a29f;
      41628: inst = 32'h13e00001;
      41629: inst = 32'hfe0d96a;
      41630: inst = 32'h5be00000;
      41631: inst = 32'h8c50000;
      41632: inst = 32'h24612800;
      41633: inst = 32'h10a0ffff;
      41634: inst = 32'hca0ffe4;
      41635: inst = 32'h24822800;
      41636: inst = 32'h10a00000;
      41637: inst = 32'hca00004;
      41638: inst = 32'h38632800;
      41639: inst = 32'h38842800;
      41640: inst = 32'h10a00000;
      41641: inst = 32'hca0a2ad;
      41642: inst = 32'h13e00001;
      41643: inst = 32'hfe0d96a;
      41644: inst = 32'h5be00000;
      41645: inst = 32'h8c50000;
      41646: inst = 32'h24612800;
      41647: inst = 32'h10a0ffff;
      41648: inst = 32'hca0ffe4;
      41649: inst = 32'h24822800;
      41650: inst = 32'h10a00000;
      41651: inst = 32'hca00004;
      41652: inst = 32'h38632800;
      41653: inst = 32'h38842800;
      41654: inst = 32'h10a00000;
      41655: inst = 32'hca0a2bb;
      41656: inst = 32'h13e00001;
      41657: inst = 32'hfe0d96a;
      41658: inst = 32'h5be00000;
      41659: inst = 32'h8c50000;
      41660: inst = 32'h24612800;
      41661: inst = 32'h10a0ffff;
      41662: inst = 32'hca0ffe4;
      41663: inst = 32'h24822800;
      41664: inst = 32'h10a00000;
      41665: inst = 32'hca00004;
      41666: inst = 32'h38632800;
      41667: inst = 32'h38842800;
      41668: inst = 32'h10a00000;
      41669: inst = 32'hca0a2c9;
      41670: inst = 32'h13e00001;
      41671: inst = 32'hfe0d96a;
      41672: inst = 32'h5be00000;
      41673: inst = 32'h8c50000;
      41674: inst = 32'h24612800;
      41675: inst = 32'h10a0ffff;
      41676: inst = 32'hca0ffe4;
      41677: inst = 32'h24822800;
      41678: inst = 32'h10a00000;
      41679: inst = 32'hca00004;
      41680: inst = 32'h38632800;
      41681: inst = 32'h38842800;
      41682: inst = 32'h10a00000;
      41683: inst = 32'hca0a2d7;
      41684: inst = 32'h13e00001;
      41685: inst = 32'hfe0d96a;
      41686: inst = 32'h5be00000;
      41687: inst = 32'h8c50000;
      41688: inst = 32'h24612800;
      41689: inst = 32'h10a0ffff;
      41690: inst = 32'hca0ffe4;
      41691: inst = 32'h24822800;
      41692: inst = 32'h10a00000;
      41693: inst = 32'hca00004;
      41694: inst = 32'h38632800;
      41695: inst = 32'h38842800;
      41696: inst = 32'h10a00000;
      41697: inst = 32'hca0a2e5;
      41698: inst = 32'h13e00001;
      41699: inst = 32'hfe0d96a;
      41700: inst = 32'h5be00000;
      41701: inst = 32'h8c50000;
      41702: inst = 32'h24612800;
      41703: inst = 32'h10a0ffff;
      41704: inst = 32'hca0ffe4;
      41705: inst = 32'h24822800;
      41706: inst = 32'h10a00000;
      41707: inst = 32'hca00004;
      41708: inst = 32'h38632800;
      41709: inst = 32'h38842800;
      41710: inst = 32'h10a00000;
      41711: inst = 32'hca0a2f3;
      41712: inst = 32'h13e00001;
      41713: inst = 32'hfe0d96a;
      41714: inst = 32'h5be00000;
      41715: inst = 32'h8c50000;
      41716: inst = 32'h24612800;
      41717: inst = 32'h10a0ffff;
      41718: inst = 32'hca0ffe4;
      41719: inst = 32'h24822800;
      41720: inst = 32'h10a00000;
      41721: inst = 32'hca00004;
      41722: inst = 32'h38632800;
      41723: inst = 32'h38842800;
      41724: inst = 32'h10a00000;
      41725: inst = 32'hca0a301;
      41726: inst = 32'h13e00001;
      41727: inst = 32'hfe0d96a;
      41728: inst = 32'h5be00000;
      41729: inst = 32'h8c50000;
      41730: inst = 32'h24612800;
      41731: inst = 32'h10a0ffff;
      41732: inst = 32'hca0ffe4;
      41733: inst = 32'h24822800;
      41734: inst = 32'h10a00000;
      41735: inst = 32'hca00004;
      41736: inst = 32'h38632800;
      41737: inst = 32'h38842800;
      41738: inst = 32'h10a00000;
      41739: inst = 32'hca0a30f;
      41740: inst = 32'h13e00001;
      41741: inst = 32'hfe0d96a;
      41742: inst = 32'h5be00000;
      41743: inst = 32'h8c50000;
      41744: inst = 32'h24612800;
      41745: inst = 32'h10a0ffff;
      41746: inst = 32'hca0ffe4;
      41747: inst = 32'h24822800;
      41748: inst = 32'h10a00000;
      41749: inst = 32'hca00004;
      41750: inst = 32'h38632800;
      41751: inst = 32'h38842800;
      41752: inst = 32'h10a00000;
      41753: inst = 32'hca0a31d;
      41754: inst = 32'h13e00001;
      41755: inst = 32'hfe0d96a;
      41756: inst = 32'h5be00000;
      41757: inst = 32'h8c50000;
      41758: inst = 32'h24612800;
      41759: inst = 32'h10a0ffff;
      41760: inst = 32'hca0ffe4;
      41761: inst = 32'h24822800;
      41762: inst = 32'h10a00000;
      41763: inst = 32'hca00004;
      41764: inst = 32'h38632800;
      41765: inst = 32'h38842800;
      41766: inst = 32'h10a00000;
      41767: inst = 32'hca0a32b;
      41768: inst = 32'h13e00001;
      41769: inst = 32'hfe0d96a;
      41770: inst = 32'h5be00000;
      41771: inst = 32'h8c50000;
      41772: inst = 32'h24612800;
      41773: inst = 32'h10a0ffff;
      41774: inst = 32'hca0ffe4;
      41775: inst = 32'h24822800;
      41776: inst = 32'h10a00000;
      41777: inst = 32'hca00004;
      41778: inst = 32'h38632800;
      41779: inst = 32'h38842800;
      41780: inst = 32'h10a00000;
      41781: inst = 32'hca0a339;
      41782: inst = 32'h13e00001;
      41783: inst = 32'hfe0d96a;
      41784: inst = 32'h5be00000;
      41785: inst = 32'h8c50000;
      41786: inst = 32'h24612800;
      41787: inst = 32'h10a0ffff;
      41788: inst = 32'hca0ffe4;
      41789: inst = 32'h24822800;
      41790: inst = 32'h10a00000;
      41791: inst = 32'hca00004;
      41792: inst = 32'h38632800;
      41793: inst = 32'h38842800;
      41794: inst = 32'h10a00000;
      41795: inst = 32'hca0a347;
      41796: inst = 32'h13e00001;
      41797: inst = 32'hfe0d96a;
      41798: inst = 32'h5be00000;
      41799: inst = 32'h8c50000;
      41800: inst = 32'h24612800;
      41801: inst = 32'h10a0ffff;
      41802: inst = 32'hca0ffe4;
      41803: inst = 32'h24822800;
      41804: inst = 32'h10a00000;
      41805: inst = 32'hca00004;
      41806: inst = 32'h38632800;
      41807: inst = 32'h38842800;
      41808: inst = 32'h10a00000;
      41809: inst = 32'hca0a355;
      41810: inst = 32'h13e00001;
      41811: inst = 32'hfe0d96a;
      41812: inst = 32'h5be00000;
      41813: inst = 32'h8c50000;
      41814: inst = 32'h24612800;
      41815: inst = 32'h10a0ffff;
      41816: inst = 32'hca0ffe4;
      41817: inst = 32'h24822800;
      41818: inst = 32'h10a00000;
      41819: inst = 32'hca00004;
      41820: inst = 32'h38632800;
      41821: inst = 32'h38842800;
      41822: inst = 32'h10a00000;
      41823: inst = 32'hca0a363;
      41824: inst = 32'h13e00001;
      41825: inst = 32'hfe0d96a;
      41826: inst = 32'h5be00000;
      41827: inst = 32'h8c50000;
      41828: inst = 32'h24612800;
      41829: inst = 32'h10a0ffff;
      41830: inst = 32'hca0ffe4;
      41831: inst = 32'h24822800;
      41832: inst = 32'h10a00000;
      41833: inst = 32'hca00004;
      41834: inst = 32'h38632800;
      41835: inst = 32'h38842800;
      41836: inst = 32'h10a00000;
      41837: inst = 32'hca0a371;
      41838: inst = 32'h13e00001;
      41839: inst = 32'hfe0d96a;
      41840: inst = 32'h5be00000;
      41841: inst = 32'h8c50000;
      41842: inst = 32'h24612800;
      41843: inst = 32'h10a0ffff;
      41844: inst = 32'hca0ffe4;
      41845: inst = 32'h24822800;
      41846: inst = 32'h10a00000;
      41847: inst = 32'hca00004;
      41848: inst = 32'h38632800;
      41849: inst = 32'h38842800;
      41850: inst = 32'h10a00000;
      41851: inst = 32'hca0a37f;
      41852: inst = 32'h13e00001;
      41853: inst = 32'hfe0d96a;
      41854: inst = 32'h5be00000;
      41855: inst = 32'h8c50000;
      41856: inst = 32'h24612800;
      41857: inst = 32'h10a0ffff;
      41858: inst = 32'hca0ffe4;
      41859: inst = 32'h24822800;
      41860: inst = 32'h10a00000;
      41861: inst = 32'hca00004;
      41862: inst = 32'h38632800;
      41863: inst = 32'h38842800;
      41864: inst = 32'h10a00000;
      41865: inst = 32'hca0a38d;
      41866: inst = 32'h13e00001;
      41867: inst = 32'hfe0d96a;
      41868: inst = 32'h5be00000;
      41869: inst = 32'h8c50000;
      41870: inst = 32'h24612800;
      41871: inst = 32'h10a0ffff;
      41872: inst = 32'hca0ffe4;
      41873: inst = 32'h24822800;
      41874: inst = 32'h10a00000;
      41875: inst = 32'hca00004;
      41876: inst = 32'h38632800;
      41877: inst = 32'h38842800;
      41878: inst = 32'h10a00000;
      41879: inst = 32'hca0a39b;
      41880: inst = 32'h13e00001;
      41881: inst = 32'hfe0d96a;
      41882: inst = 32'h5be00000;
      41883: inst = 32'h8c50000;
      41884: inst = 32'h24612800;
      41885: inst = 32'h10a0ffff;
      41886: inst = 32'hca0ffe4;
      41887: inst = 32'h24822800;
      41888: inst = 32'h10a00000;
      41889: inst = 32'hca00004;
      41890: inst = 32'h38632800;
      41891: inst = 32'h38842800;
      41892: inst = 32'h10a00000;
      41893: inst = 32'hca0a3a9;
      41894: inst = 32'h13e00001;
      41895: inst = 32'hfe0d96a;
      41896: inst = 32'h5be00000;
      41897: inst = 32'h8c50000;
      41898: inst = 32'h24612800;
      41899: inst = 32'h10a0ffff;
      41900: inst = 32'hca0ffe5;
      41901: inst = 32'h24822800;
      41902: inst = 32'h10a00000;
      41903: inst = 32'hca00004;
      41904: inst = 32'h38632800;
      41905: inst = 32'h38842800;
      41906: inst = 32'h10a00000;
      41907: inst = 32'hca0a3b7;
      41908: inst = 32'h13e00001;
      41909: inst = 32'hfe0d96a;
      41910: inst = 32'h5be00000;
      41911: inst = 32'h8c50000;
      41912: inst = 32'h24612800;
      41913: inst = 32'h10a0ffff;
      41914: inst = 32'hca0ffe5;
      41915: inst = 32'h24822800;
      41916: inst = 32'h10a00000;
      41917: inst = 32'hca00004;
      41918: inst = 32'h38632800;
      41919: inst = 32'h38842800;
      41920: inst = 32'h10a00000;
      41921: inst = 32'hca0a3c5;
      41922: inst = 32'h13e00001;
      41923: inst = 32'hfe0d96a;
      41924: inst = 32'h5be00000;
      41925: inst = 32'h8c50000;
      41926: inst = 32'h24612800;
      41927: inst = 32'h10a0ffff;
      41928: inst = 32'hca0ffe5;
      41929: inst = 32'h24822800;
      41930: inst = 32'h10a00000;
      41931: inst = 32'hca00004;
      41932: inst = 32'h38632800;
      41933: inst = 32'h38842800;
      41934: inst = 32'h10a00000;
      41935: inst = 32'hca0a3d3;
      41936: inst = 32'h13e00001;
      41937: inst = 32'hfe0d96a;
      41938: inst = 32'h5be00000;
      41939: inst = 32'h8c50000;
      41940: inst = 32'h24612800;
      41941: inst = 32'h10a0ffff;
      41942: inst = 32'hca0ffe5;
      41943: inst = 32'h24822800;
      41944: inst = 32'h10a00000;
      41945: inst = 32'hca00004;
      41946: inst = 32'h38632800;
      41947: inst = 32'h38842800;
      41948: inst = 32'h10a00000;
      41949: inst = 32'hca0a3e1;
      41950: inst = 32'h13e00001;
      41951: inst = 32'hfe0d96a;
      41952: inst = 32'h5be00000;
      41953: inst = 32'h8c50000;
      41954: inst = 32'h24612800;
      41955: inst = 32'h10a0ffff;
      41956: inst = 32'hca0ffe5;
      41957: inst = 32'h24822800;
      41958: inst = 32'h10a00000;
      41959: inst = 32'hca00004;
      41960: inst = 32'h38632800;
      41961: inst = 32'h38842800;
      41962: inst = 32'h10a00000;
      41963: inst = 32'hca0a3ef;
      41964: inst = 32'h13e00001;
      41965: inst = 32'hfe0d96a;
      41966: inst = 32'h5be00000;
      41967: inst = 32'h8c50000;
      41968: inst = 32'h24612800;
      41969: inst = 32'h10a0ffff;
      41970: inst = 32'hca0ffe5;
      41971: inst = 32'h24822800;
      41972: inst = 32'h10a00000;
      41973: inst = 32'hca00004;
      41974: inst = 32'h38632800;
      41975: inst = 32'h38842800;
      41976: inst = 32'h10a00000;
      41977: inst = 32'hca0a3fd;
      41978: inst = 32'h13e00001;
      41979: inst = 32'hfe0d96a;
      41980: inst = 32'h5be00000;
      41981: inst = 32'h8c50000;
      41982: inst = 32'h24612800;
      41983: inst = 32'h10a0ffff;
      41984: inst = 32'hca0ffe5;
      41985: inst = 32'h24822800;
      41986: inst = 32'h10a00000;
      41987: inst = 32'hca00004;
      41988: inst = 32'h38632800;
      41989: inst = 32'h38842800;
      41990: inst = 32'h10a00000;
      41991: inst = 32'hca0a40b;
      41992: inst = 32'h13e00001;
      41993: inst = 32'hfe0d96a;
      41994: inst = 32'h5be00000;
      41995: inst = 32'h8c50000;
      41996: inst = 32'h24612800;
      41997: inst = 32'h10a0ffff;
      41998: inst = 32'hca0ffe5;
      41999: inst = 32'h24822800;
      42000: inst = 32'h10a00000;
      42001: inst = 32'hca00004;
      42002: inst = 32'h38632800;
      42003: inst = 32'h38842800;
      42004: inst = 32'h10a00000;
      42005: inst = 32'hca0a419;
      42006: inst = 32'h13e00001;
      42007: inst = 32'hfe0d96a;
      42008: inst = 32'h5be00000;
      42009: inst = 32'h8c50000;
      42010: inst = 32'h24612800;
      42011: inst = 32'h10a0ffff;
      42012: inst = 32'hca0ffe5;
      42013: inst = 32'h24822800;
      42014: inst = 32'h10a00000;
      42015: inst = 32'hca00004;
      42016: inst = 32'h38632800;
      42017: inst = 32'h38842800;
      42018: inst = 32'h10a00000;
      42019: inst = 32'hca0a427;
      42020: inst = 32'h13e00001;
      42021: inst = 32'hfe0d96a;
      42022: inst = 32'h5be00000;
      42023: inst = 32'h8c50000;
      42024: inst = 32'h24612800;
      42025: inst = 32'h10a0ffff;
      42026: inst = 32'hca0ffe5;
      42027: inst = 32'h24822800;
      42028: inst = 32'h10a00000;
      42029: inst = 32'hca00004;
      42030: inst = 32'h38632800;
      42031: inst = 32'h38842800;
      42032: inst = 32'h10a00000;
      42033: inst = 32'hca0a435;
      42034: inst = 32'h13e00001;
      42035: inst = 32'hfe0d96a;
      42036: inst = 32'h5be00000;
      42037: inst = 32'h8c50000;
      42038: inst = 32'h24612800;
      42039: inst = 32'h10a0ffff;
      42040: inst = 32'hca0ffe5;
      42041: inst = 32'h24822800;
      42042: inst = 32'h10a00000;
      42043: inst = 32'hca00004;
      42044: inst = 32'h38632800;
      42045: inst = 32'h38842800;
      42046: inst = 32'h10a00000;
      42047: inst = 32'hca0a443;
      42048: inst = 32'h13e00001;
      42049: inst = 32'hfe0d96a;
      42050: inst = 32'h5be00000;
      42051: inst = 32'h8c50000;
      42052: inst = 32'h24612800;
      42053: inst = 32'h10a0ffff;
      42054: inst = 32'hca0ffe5;
      42055: inst = 32'h24822800;
      42056: inst = 32'h10a00000;
      42057: inst = 32'hca00004;
      42058: inst = 32'h38632800;
      42059: inst = 32'h38842800;
      42060: inst = 32'h10a00000;
      42061: inst = 32'hca0a451;
      42062: inst = 32'h13e00001;
      42063: inst = 32'hfe0d96a;
      42064: inst = 32'h5be00000;
      42065: inst = 32'h8c50000;
      42066: inst = 32'h24612800;
      42067: inst = 32'h10a0ffff;
      42068: inst = 32'hca0ffe5;
      42069: inst = 32'h24822800;
      42070: inst = 32'h10a00000;
      42071: inst = 32'hca00004;
      42072: inst = 32'h38632800;
      42073: inst = 32'h38842800;
      42074: inst = 32'h10a00000;
      42075: inst = 32'hca0a45f;
      42076: inst = 32'h13e00001;
      42077: inst = 32'hfe0d96a;
      42078: inst = 32'h5be00000;
      42079: inst = 32'h8c50000;
      42080: inst = 32'h24612800;
      42081: inst = 32'h10a0ffff;
      42082: inst = 32'hca0ffe5;
      42083: inst = 32'h24822800;
      42084: inst = 32'h10a00000;
      42085: inst = 32'hca00004;
      42086: inst = 32'h38632800;
      42087: inst = 32'h38842800;
      42088: inst = 32'h10a00000;
      42089: inst = 32'hca0a46d;
      42090: inst = 32'h13e00001;
      42091: inst = 32'hfe0d96a;
      42092: inst = 32'h5be00000;
      42093: inst = 32'h8c50000;
      42094: inst = 32'h24612800;
      42095: inst = 32'h10a0ffff;
      42096: inst = 32'hca0ffe5;
      42097: inst = 32'h24822800;
      42098: inst = 32'h10a00000;
      42099: inst = 32'hca00004;
      42100: inst = 32'h38632800;
      42101: inst = 32'h38842800;
      42102: inst = 32'h10a00000;
      42103: inst = 32'hca0a47b;
      42104: inst = 32'h13e00001;
      42105: inst = 32'hfe0d96a;
      42106: inst = 32'h5be00000;
      42107: inst = 32'h8c50000;
      42108: inst = 32'h24612800;
      42109: inst = 32'h10a0ffff;
      42110: inst = 32'hca0ffe5;
      42111: inst = 32'h24822800;
      42112: inst = 32'h10a00000;
      42113: inst = 32'hca00004;
      42114: inst = 32'h38632800;
      42115: inst = 32'h38842800;
      42116: inst = 32'h10a00000;
      42117: inst = 32'hca0a489;
      42118: inst = 32'h13e00001;
      42119: inst = 32'hfe0d96a;
      42120: inst = 32'h5be00000;
      42121: inst = 32'h8c50000;
      42122: inst = 32'h24612800;
      42123: inst = 32'h10a0ffff;
      42124: inst = 32'hca0ffe5;
      42125: inst = 32'h24822800;
      42126: inst = 32'h10a00000;
      42127: inst = 32'hca00004;
      42128: inst = 32'h38632800;
      42129: inst = 32'h38842800;
      42130: inst = 32'h10a00000;
      42131: inst = 32'hca0a497;
      42132: inst = 32'h13e00001;
      42133: inst = 32'hfe0d96a;
      42134: inst = 32'h5be00000;
      42135: inst = 32'h8c50000;
      42136: inst = 32'h24612800;
      42137: inst = 32'h10a0ffff;
      42138: inst = 32'hca0ffe5;
      42139: inst = 32'h24822800;
      42140: inst = 32'h10a00000;
      42141: inst = 32'hca00004;
      42142: inst = 32'h38632800;
      42143: inst = 32'h38842800;
      42144: inst = 32'h10a00000;
      42145: inst = 32'hca0a4a5;
      42146: inst = 32'h13e00001;
      42147: inst = 32'hfe0d96a;
      42148: inst = 32'h5be00000;
      42149: inst = 32'h8c50000;
      42150: inst = 32'h24612800;
      42151: inst = 32'h10a0ffff;
      42152: inst = 32'hca0ffe5;
      42153: inst = 32'h24822800;
      42154: inst = 32'h10a00000;
      42155: inst = 32'hca00004;
      42156: inst = 32'h38632800;
      42157: inst = 32'h38842800;
      42158: inst = 32'h10a00000;
      42159: inst = 32'hca0a4b3;
      42160: inst = 32'h13e00001;
      42161: inst = 32'hfe0d96a;
      42162: inst = 32'h5be00000;
      42163: inst = 32'h8c50000;
      42164: inst = 32'h24612800;
      42165: inst = 32'h10a0ffff;
      42166: inst = 32'hca0ffe5;
      42167: inst = 32'h24822800;
      42168: inst = 32'h10a00000;
      42169: inst = 32'hca00004;
      42170: inst = 32'h38632800;
      42171: inst = 32'h38842800;
      42172: inst = 32'h10a00000;
      42173: inst = 32'hca0a4c1;
      42174: inst = 32'h13e00001;
      42175: inst = 32'hfe0d96a;
      42176: inst = 32'h5be00000;
      42177: inst = 32'h8c50000;
      42178: inst = 32'h24612800;
      42179: inst = 32'h10a0ffff;
      42180: inst = 32'hca0ffe5;
      42181: inst = 32'h24822800;
      42182: inst = 32'h10a00000;
      42183: inst = 32'hca00004;
      42184: inst = 32'h38632800;
      42185: inst = 32'h38842800;
      42186: inst = 32'h10a00000;
      42187: inst = 32'hca0a4cf;
      42188: inst = 32'h13e00001;
      42189: inst = 32'hfe0d96a;
      42190: inst = 32'h5be00000;
      42191: inst = 32'h8c50000;
      42192: inst = 32'h24612800;
      42193: inst = 32'h10a0ffff;
      42194: inst = 32'hca0ffe5;
      42195: inst = 32'h24822800;
      42196: inst = 32'h10a00000;
      42197: inst = 32'hca00004;
      42198: inst = 32'h38632800;
      42199: inst = 32'h38842800;
      42200: inst = 32'h10a00000;
      42201: inst = 32'hca0a4dd;
      42202: inst = 32'h13e00001;
      42203: inst = 32'hfe0d96a;
      42204: inst = 32'h5be00000;
      42205: inst = 32'h8c50000;
      42206: inst = 32'h24612800;
      42207: inst = 32'h10a0ffff;
      42208: inst = 32'hca0ffe5;
      42209: inst = 32'h24822800;
      42210: inst = 32'h10a00000;
      42211: inst = 32'hca00004;
      42212: inst = 32'h38632800;
      42213: inst = 32'h38842800;
      42214: inst = 32'h10a00000;
      42215: inst = 32'hca0a4eb;
      42216: inst = 32'h13e00001;
      42217: inst = 32'hfe0d96a;
      42218: inst = 32'h5be00000;
      42219: inst = 32'h8c50000;
      42220: inst = 32'h24612800;
      42221: inst = 32'h10a0ffff;
      42222: inst = 32'hca0ffe5;
      42223: inst = 32'h24822800;
      42224: inst = 32'h10a00000;
      42225: inst = 32'hca00004;
      42226: inst = 32'h38632800;
      42227: inst = 32'h38842800;
      42228: inst = 32'h10a00000;
      42229: inst = 32'hca0a4f9;
      42230: inst = 32'h13e00001;
      42231: inst = 32'hfe0d96a;
      42232: inst = 32'h5be00000;
      42233: inst = 32'h8c50000;
      42234: inst = 32'h24612800;
      42235: inst = 32'h10a0ffff;
      42236: inst = 32'hca0ffe5;
      42237: inst = 32'h24822800;
      42238: inst = 32'h10a00000;
      42239: inst = 32'hca00004;
      42240: inst = 32'h38632800;
      42241: inst = 32'h38842800;
      42242: inst = 32'h10a00000;
      42243: inst = 32'hca0a507;
      42244: inst = 32'h13e00001;
      42245: inst = 32'hfe0d96a;
      42246: inst = 32'h5be00000;
      42247: inst = 32'h8c50000;
      42248: inst = 32'h24612800;
      42249: inst = 32'h10a0ffff;
      42250: inst = 32'hca0ffe5;
      42251: inst = 32'h24822800;
      42252: inst = 32'h10a00000;
      42253: inst = 32'hca00004;
      42254: inst = 32'h38632800;
      42255: inst = 32'h38842800;
      42256: inst = 32'h10a00000;
      42257: inst = 32'hca0a515;
      42258: inst = 32'h13e00001;
      42259: inst = 32'hfe0d96a;
      42260: inst = 32'h5be00000;
      42261: inst = 32'h8c50000;
      42262: inst = 32'h24612800;
      42263: inst = 32'h10a0ffff;
      42264: inst = 32'hca0ffe5;
      42265: inst = 32'h24822800;
      42266: inst = 32'h10a00000;
      42267: inst = 32'hca00004;
      42268: inst = 32'h38632800;
      42269: inst = 32'h38842800;
      42270: inst = 32'h10a00000;
      42271: inst = 32'hca0a523;
      42272: inst = 32'h13e00001;
      42273: inst = 32'hfe0d96a;
      42274: inst = 32'h5be00000;
      42275: inst = 32'h8c50000;
      42276: inst = 32'h24612800;
      42277: inst = 32'h10a0ffff;
      42278: inst = 32'hca0ffe5;
      42279: inst = 32'h24822800;
      42280: inst = 32'h10a00000;
      42281: inst = 32'hca00004;
      42282: inst = 32'h38632800;
      42283: inst = 32'h38842800;
      42284: inst = 32'h10a00000;
      42285: inst = 32'hca0a531;
      42286: inst = 32'h13e00001;
      42287: inst = 32'hfe0d96a;
      42288: inst = 32'h5be00000;
      42289: inst = 32'h8c50000;
      42290: inst = 32'h24612800;
      42291: inst = 32'h10a0ffff;
      42292: inst = 32'hca0ffe5;
      42293: inst = 32'h24822800;
      42294: inst = 32'h10a00000;
      42295: inst = 32'hca00004;
      42296: inst = 32'h38632800;
      42297: inst = 32'h38842800;
      42298: inst = 32'h10a00000;
      42299: inst = 32'hca0a53f;
      42300: inst = 32'h13e00001;
      42301: inst = 32'hfe0d96a;
      42302: inst = 32'h5be00000;
      42303: inst = 32'h8c50000;
      42304: inst = 32'h24612800;
      42305: inst = 32'h10a0ffff;
      42306: inst = 32'hca0ffe5;
      42307: inst = 32'h24822800;
      42308: inst = 32'h10a00000;
      42309: inst = 32'hca00004;
      42310: inst = 32'h38632800;
      42311: inst = 32'h38842800;
      42312: inst = 32'h10a00000;
      42313: inst = 32'hca0a54d;
      42314: inst = 32'h13e00001;
      42315: inst = 32'hfe0d96a;
      42316: inst = 32'h5be00000;
      42317: inst = 32'h8c50000;
      42318: inst = 32'h24612800;
      42319: inst = 32'h10a0ffff;
      42320: inst = 32'hca0ffe5;
      42321: inst = 32'h24822800;
      42322: inst = 32'h10a00000;
      42323: inst = 32'hca00004;
      42324: inst = 32'h38632800;
      42325: inst = 32'h38842800;
      42326: inst = 32'h10a00000;
      42327: inst = 32'hca0a55b;
      42328: inst = 32'h13e00001;
      42329: inst = 32'hfe0d96a;
      42330: inst = 32'h5be00000;
      42331: inst = 32'h8c50000;
      42332: inst = 32'h24612800;
      42333: inst = 32'h10a0ffff;
      42334: inst = 32'hca0ffe5;
      42335: inst = 32'h24822800;
      42336: inst = 32'h10a00000;
      42337: inst = 32'hca00004;
      42338: inst = 32'h38632800;
      42339: inst = 32'h38842800;
      42340: inst = 32'h10a00000;
      42341: inst = 32'hca0a569;
      42342: inst = 32'h13e00001;
      42343: inst = 32'hfe0d96a;
      42344: inst = 32'h5be00000;
      42345: inst = 32'h8c50000;
      42346: inst = 32'h24612800;
      42347: inst = 32'h10a0ffff;
      42348: inst = 32'hca0ffe5;
      42349: inst = 32'h24822800;
      42350: inst = 32'h10a00000;
      42351: inst = 32'hca00004;
      42352: inst = 32'h38632800;
      42353: inst = 32'h38842800;
      42354: inst = 32'h10a00000;
      42355: inst = 32'hca0a577;
      42356: inst = 32'h13e00001;
      42357: inst = 32'hfe0d96a;
      42358: inst = 32'h5be00000;
      42359: inst = 32'h8c50000;
      42360: inst = 32'h24612800;
      42361: inst = 32'h10a0ffff;
      42362: inst = 32'hca0ffe5;
      42363: inst = 32'h24822800;
      42364: inst = 32'h10a00000;
      42365: inst = 32'hca00004;
      42366: inst = 32'h38632800;
      42367: inst = 32'h38842800;
      42368: inst = 32'h10a00000;
      42369: inst = 32'hca0a585;
      42370: inst = 32'h13e00001;
      42371: inst = 32'hfe0d96a;
      42372: inst = 32'h5be00000;
      42373: inst = 32'h8c50000;
      42374: inst = 32'h24612800;
      42375: inst = 32'h10a0ffff;
      42376: inst = 32'hca0ffe5;
      42377: inst = 32'h24822800;
      42378: inst = 32'h10a00000;
      42379: inst = 32'hca00004;
      42380: inst = 32'h38632800;
      42381: inst = 32'h38842800;
      42382: inst = 32'h10a00000;
      42383: inst = 32'hca0a593;
      42384: inst = 32'h13e00001;
      42385: inst = 32'hfe0d96a;
      42386: inst = 32'h5be00000;
      42387: inst = 32'h8c50000;
      42388: inst = 32'h24612800;
      42389: inst = 32'h10a0ffff;
      42390: inst = 32'hca0ffe5;
      42391: inst = 32'h24822800;
      42392: inst = 32'h10a00000;
      42393: inst = 32'hca00004;
      42394: inst = 32'h38632800;
      42395: inst = 32'h38842800;
      42396: inst = 32'h10a00000;
      42397: inst = 32'hca0a5a1;
      42398: inst = 32'h13e00001;
      42399: inst = 32'hfe0d96a;
      42400: inst = 32'h5be00000;
      42401: inst = 32'h8c50000;
      42402: inst = 32'h24612800;
      42403: inst = 32'h10a0ffff;
      42404: inst = 32'hca0ffe5;
      42405: inst = 32'h24822800;
      42406: inst = 32'h10a00000;
      42407: inst = 32'hca00004;
      42408: inst = 32'h38632800;
      42409: inst = 32'h38842800;
      42410: inst = 32'h10a00000;
      42411: inst = 32'hca0a5af;
      42412: inst = 32'h13e00001;
      42413: inst = 32'hfe0d96a;
      42414: inst = 32'h5be00000;
      42415: inst = 32'h8c50000;
      42416: inst = 32'h24612800;
      42417: inst = 32'h10a0ffff;
      42418: inst = 32'hca0ffe5;
      42419: inst = 32'h24822800;
      42420: inst = 32'h10a00000;
      42421: inst = 32'hca00004;
      42422: inst = 32'h38632800;
      42423: inst = 32'h38842800;
      42424: inst = 32'h10a00000;
      42425: inst = 32'hca0a5bd;
      42426: inst = 32'h13e00001;
      42427: inst = 32'hfe0d96a;
      42428: inst = 32'h5be00000;
      42429: inst = 32'h8c50000;
      42430: inst = 32'h24612800;
      42431: inst = 32'h10a0ffff;
      42432: inst = 32'hca0ffe5;
      42433: inst = 32'h24822800;
      42434: inst = 32'h10a00000;
      42435: inst = 32'hca00004;
      42436: inst = 32'h38632800;
      42437: inst = 32'h38842800;
      42438: inst = 32'h10a00000;
      42439: inst = 32'hca0a5cb;
      42440: inst = 32'h13e00001;
      42441: inst = 32'hfe0d96a;
      42442: inst = 32'h5be00000;
      42443: inst = 32'h8c50000;
      42444: inst = 32'h24612800;
      42445: inst = 32'h10a0ffff;
      42446: inst = 32'hca0ffe5;
      42447: inst = 32'h24822800;
      42448: inst = 32'h10a00000;
      42449: inst = 32'hca00004;
      42450: inst = 32'h38632800;
      42451: inst = 32'h38842800;
      42452: inst = 32'h10a00000;
      42453: inst = 32'hca0a5d9;
      42454: inst = 32'h13e00001;
      42455: inst = 32'hfe0d96a;
      42456: inst = 32'h5be00000;
      42457: inst = 32'h8c50000;
      42458: inst = 32'h24612800;
      42459: inst = 32'h10a0ffff;
      42460: inst = 32'hca0ffe5;
      42461: inst = 32'h24822800;
      42462: inst = 32'h10a00000;
      42463: inst = 32'hca00004;
      42464: inst = 32'h38632800;
      42465: inst = 32'h38842800;
      42466: inst = 32'h10a00000;
      42467: inst = 32'hca0a5e7;
      42468: inst = 32'h13e00001;
      42469: inst = 32'hfe0d96a;
      42470: inst = 32'h5be00000;
      42471: inst = 32'h8c50000;
      42472: inst = 32'h24612800;
      42473: inst = 32'h10a0ffff;
      42474: inst = 32'hca0ffe5;
      42475: inst = 32'h24822800;
      42476: inst = 32'h10a00000;
      42477: inst = 32'hca00004;
      42478: inst = 32'h38632800;
      42479: inst = 32'h38842800;
      42480: inst = 32'h10a00000;
      42481: inst = 32'hca0a5f5;
      42482: inst = 32'h13e00001;
      42483: inst = 32'hfe0d96a;
      42484: inst = 32'h5be00000;
      42485: inst = 32'h8c50000;
      42486: inst = 32'h24612800;
      42487: inst = 32'h10a0ffff;
      42488: inst = 32'hca0ffe5;
      42489: inst = 32'h24822800;
      42490: inst = 32'h10a00000;
      42491: inst = 32'hca00004;
      42492: inst = 32'h38632800;
      42493: inst = 32'h38842800;
      42494: inst = 32'h10a00000;
      42495: inst = 32'hca0a603;
      42496: inst = 32'h13e00001;
      42497: inst = 32'hfe0d96a;
      42498: inst = 32'h5be00000;
      42499: inst = 32'h8c50000;
      42500: inst = 32'h24612800;
      42501: inst = 32'h10a0ffff;
      42502: inst = 32'hca0ffe5;
      42503: inst = 32'h24822800;
      42504: inst = 32'h10a00000;
      42505: inst = 32'hca00004;
      42506: inst = 32'h38632800;
      42507: inst = 32'h38842800;
      42508: inst = 32'h10a00000;
      42509: inst = 32'hca0a611;
      42510: inst = 32'h13e00001;
      42511: inst = 32'hfe0d96a;
      42512: inst = 32'h5be00000;
      42513: inst = 32'h8c50000;
      42514: inst = 32'h24612800;
      42515: inst = 32'h10a0ffff;
      42516: inst = 32'hca0ffe5;
      42517: inst = 32'h24822800;
      42518: inst = 32'h10a00000;
      42519: inst = 32'hca00004;
      42520: inst = 32'h38632800;
      42521: inst = 32'h38842800;
      42522: inst = 32'h10a00000;
      42523: inst = 32'hca0a61f;
      42524: inst = 32'h13e00001;
      42525: inst = 32'hfe0d96a;
      42526: inst = 32'h5be00000;
      42527: inst = 32'h8c50000;
      42528: inst = 32'h24612800;
      42529: inst = 32'h10a0ffff;
      42530: inst = 32'hca0ffe5;
      42531: inst = 32'h24822800;
      42532: inst = 32'h10a00000;
      42533: inst = 32'hca00004;
      42534: inst = 32'h38632800;
      42535: inst = 32'h38842800;
      42536: inst = 32'h10a00000;
      42537: inst = 32'hca0a62d;
      42538: inst = 32'h13e00001;
      42539: inst = 32'hfe0d96a;
      42540: inst = 32'h5be00000;
      42541: inst = 32'h8c50000;
      42542: inst = 32'h24612800;
      42543: inst = 32'h10a0ffff;
      42544: inst = 32'hca0ffe5;
      42545: inst = 32'h24822800;
      42546: inst = 32'h10a00000;
      42547: inst = 32'hca00004;
      42548: inst = 32'h38632800;
      42549: inst = 32'h38842800;
      42550: inst = 32'h10a00000;
      42551: inst = 32'hca0a63b;
      42552: inst = 32'h13e00001;
      42553: inst = 32'hfe0d96a;
      42554: inst = 32'h5be00000;
      42555: inst = 32'h8c50000;
      42556: inst = 32'h24612800;
      42557: inst = 32'h10a0ffff;
      42558: inst = 32'hca0ffe5;
      42559: inst = 32'h24822800;
      42560: inst = 32'h10a00000;
      42561: inst = 32'hca00004;
      42562: inst = 32'h38632800;
      42563: inst = 32'h38842800;
      42564: inst = 32'h10a00000;
      42565: inst = 32'hca0a649;
      42566: inst = 32'h13e00001;
      42567: inst = 32'hfe0d96a;
      42568: inst = 32'h5be00000;
      42569: inst = 32'h8c50000;
      42570: inst = 32'h24612800;
      42571: inst = 32'h10a0ffff;
      42572: inst = 32'hca0ffe5;
      42573: inst = 32'h24822800;
      42574: inst = 32'h10a00000;
      42575: inst = 32'hca00004;
      42576: inst = 32'h38632800;
      42577: inst = 32'h38842800;
      42578: inst = 32'h10a00000;
      42579: inst = 32'hca0a657;
      42580: inst = 32'h13e00001;
      42581: inst = 32'hfe0d96a;
      42582: inst = 32'h5be00000;
      42583: inst = 32'h8c50000;
      42584: inst = 32'h24612800;
      42585: inst = 32'h10a0ffff;
      42586: inst = 32'hca0ffe5;
      42587: inst = 32'h24822800;
      42588: inst = 32'h10a00000;
      42589: inst = 32'hca00004;
      42590: inst = 32'h38632800;
      42591: inst = 32'h38842800;
      42592: inst = 32'h10a00000;
      42593: inst = 32'hca0a665;
      42594: inst = 32'h13e00001;
      42595: inst = 32'hfe0d96a;
      42596: inst = 32'h5be00000;
      42597: inst = 32'h8c50000;
      42598: inst = 32'h24612800;
      42599: inst = 32'h10a0ffff;
      42600: inst = 32'hca0ffe5;
      42601: inst = 32'h24822800;
      42602: inst = 32'h10a00000;
      42603: inst = 32'hca00004;
      42604: inst = 32'h38632800;
      42605: inst = 32'h38842800;
      42606: inst = 32'h10a00000;
      42607: inst = 32'hca0a673;
      42608: inst = 32'h13e00001;
      42609: inst = 32'hfe0d96a;
      42610: inst = 32'h5be00000;
      42611: inst = 32'h8c50000;
      42612: inst = 32'h24612800;
      42613: inst = 32'h10a0ffff;
      42614: inst = 32'hca0ffe5;
      42615: inst = 32'h24822800;
      42616: inst = 32'h10a00000;
      42617: inst = 32'hca00004;
      42618: inst = 32'h38632800;
      42619: inst = 32'h38842800;
      42620: inst = 32'h10a00000;
      42621: inst = 32'hca0a681;
      42622: inst = 32'h13e00001;
      42623: inst = 32'hfe0d96a;
      42624: inst = 32'h5be00000;
      42625: inst = 32'h8c50000;
      42626: inst = 32'h24612800;
      42627: inst = 32'h10a0ffff;
      42628: inst = 32'hca0ffe5;
      42629: inst = 32'h24822800;
      42630: inst = 32'h10a00000;
      42631: inst = 32'hca00004;
      42632: inst = 32'h38632800;
      42633: inst = 32'h38842800;
      42634: inst = 32'h10a00000;
      42635: inst = 32'hca0a68f;
      42636: inst = 32'h13e00001;
      42637: inst = 32'hfe0d96a;
      42638: inst = 32'h5be00000;
      42639: inst = 32'h8c50000;
      42640: inst = 32'h24612800;
      42641: inst = 32'h10a0ffff;
      42642: inst = 32'hca0ffe5;
      42643: inst = 32'h24822800;
      42644: inst = 32'h10a00000;
      42645: inst = 32'hca00004;
      42646: inst = 32'h38632800;
      42647: inst = 32'h38842800;
      42648: inst = 32'h10a00000;
      42649: inst = 32'hca0a69d;
      42650: inst = 32'h13e00001;
      42651: inst = 32'hfe0d96a;
      42652: inst = 32'h5be00000;
      42653: inst = 32'h8c50000;
      42654: inst = 32'h24612800;
      42655: inst = 32'h10a0ffff;
      42656: inst = 32'hca0ffe5;
      42657: inst = 32'h24822800;
      42658: inst = 32'h10a00000;
      42659: inst = 32'hca00004;
      42660: inst = 32'h38632800;
      42661: inst = 32'h38842800;
      42662: inst = 32'h10a00000;
      42663: inst = 32'hca0a6ab;
      42664: inst = 32'h13e00001;
      42665: inst = 32'hfe0d96a;
      42666: inst = 32'h5be00000;
      42667: inst = 32'h8c50000;
      42668: inst = 32'h24612800;
      42669: inst = 32'h10a0ffff;
      42670: inst = 32'hca0ffe5;
      42671: inst = 32'h24822800;
      42672: inst = 32'h10a00000;
      42673: inst = 32'hca00004;
      42674: inst = 32'h38632800;
      42675: inst = 32'h38842800;
      42676: inst = 32'h10a00000;
      42677: inst = 32'hca0a6b9;
      42678: inst = 32'h13e00001;
      42679: inst = 32'hfe0d96a;
      42680: inst = 32'h5be00000;
      42681: inst = 32'h8c50000;
      42682: inst = 32'h24612800;
      42683: inst = 32'h10a0ffff;
      42684: inst = 32'hca0ffe5;
      42685: inst = 32'h24822800;
      42686: inst = 32'h10a00000;
      42687: inst = 32'hca00004;
      42688: inst = 32'h38632800;
      42689: inst = 32'h38842800;
      42690: inst = 32'h10a00000;
      42691: inst = 32'hca0a6c7;
      42692: inst = 32'h13e00001;
      42693: inst = 32'hfe0d96a;
      42694: inst = 32'h5be00000;
      42695: inst = 32'h8c50000;
      42696: inst = 32'h24612800;
      42697: inst = 32'h10a0ffff;
      42698: inst = 32'hca0ffe5;
      42699: inst = 32'h24822800;
      42700: inst = 32'h10a00000;
      42701: inst = 32'hca00004;
      42702: inst = 32'h38632800;
      42703: inst = 32'h38842800;
      42704: inst = 32'h10a00000;
      42705: inst = 32'hca0a6d5;
      42706: inst = 32'h13e00001;
      42707: inst = 32'hfe0d96a;
      42708: inst = 32'h5be00000;
      42709: inst = 32'h8c50000;
      42710: inst = 32'h24612800;
      42711: inst = 32'h10a0ffff;
      42712: inst = 32'hca0ffe5;
      42713: inst = 32'h24822800;
      42714: inst = 32'h10a00000;
      42715: inst = 32'hca00004;
      42716: inst = 32'h38632800;
      42717: inst = 32'h38842800;
      42718: inst = 32'h10a00000;
      42719: inst = 32'hca0a6e3;
      42720: inst = 32'h13e00001;
      42721: inst = 32'hfe0d96a;
      42722: inst = 32'h5be00000;
      42723: inst = 32'h8c50000;
      42724: inst = 32'h24612800;
      42725: inst = 32'h10a0ffff;
      42726: inst = 32'hca0ffe5;
      42727: inst = 32'h24822800;
      42728: inst = 32'h10a00000;
      42729: inst = 32'hca00004;
      42730: inst = 32'h38632800;
      42731: inst = 32'h38842800;
      42732: inst = 32'h10a00000;
      42733: inst = 32'hca0a6f1;
      42734: inst = 32'h13e00001;
      42735: inst = 32'hfe0d96a;
      42736: inst = 32'h5be00000;
      42737: inst = 32'h8c50000;
      42738: inst = 32'h24612800;
      42739: inst = 32'h10a0ffff;
      42740: inst = 32'hca0ffe5;
      42741: inst = 32'h24822800;
      42742: inst = 32'h10a00000;
      42743: inst = 32'hca00004;
      42744: inst = 32'h38632800;
      42745: inst = 32'h38842800;
      42746: inst = 32'h10a00000;
      42747: inst = 32'hca0a6ff;
      42748: inst = 32'h13e00001;
      42749: inst = 32'hfe0d96a;
      42750: inst = 32'h5be00000;
      42751: inst = 32'h8c50000;
      42752: inst = 32'h24612800;
      42753: inst = 32'h10a0ffff;
      42754: inst = 32'hca0ffe5;
      42755: inst = 32'h24822800;
      42756: inst = 32'h10a00000;
      42757: inst = 32'hca00004;
      42758: inst = 32'h38632800;
      42759: inst = 32'h38842800;
      42760: inst = 32'h10a00000;
      42761: inst = 32'hca0a70d;
      42762: inst = 32'h13e00001;
      42763: inst = 32'hfe0d96a;
      42764: inst = 32'h5be00000;
      42765: inst = 32'h8c50000;
      42766: inst = 32'h24612800;
      42767: inst = 32'h10a0ffff;
      42768: inst = 32'hca0ffe5;
      42769: inst = 32'h24822800;
      42770: inst = 32'h10a00000;
      42771: inst = 32'hca00004;
      42772: inst = 32'h38632800;
      42773: inst = 32'h38842800;
      42774: inst = 32'h10a00000;
      42775: inst = 32'hca0a71b;
      42776: inst = 32'h13e00001;
      42777: inst = 32'hfe0d96a;
      42778: inst = 32'h5be00000;
      42779: inst = 32'h8c50000;
      42780: inst = 32'h24612800;
      42781: inst = 32'h10a0ffff;
      42782: inst = 32'hca0ffe5;
      42783: inst = 32'h24822800;
      42784: inst = 32'h10a00000;
      42785: inst = 32'hca00004;
      42786: inst = 32'h38632800;
      42787: inst = 32'h38842800;
      42788: inst = 32'h10a00000;
      42789: inst = 32'hca0a729;
      42790: inst = 32'h13e00001;
      42791: inst = 32'hfe0d96a;
      42792: inst = 32'h5be00000;
      42793: inst = 32'h8c50000;
      42794: inst = 32'h24612800;
      42795: inst = 32'h10a0ffff;
      42796: inst = 32'hca0ffe5;
      42797: inst = 32'h24822800;
      42798: inst = 32'h10a00000;
      42799: inst = 32'hca00004;
      42800: inst = 32'h38632800;
      42801: inst = 32'h38842800;
      42802: inst = 32'h10a00000;
      42803: inst = 32'hca0a737;
      42804: inst = 32'h13e00001;
      42805: inst = 32'hfe0d96a;
      42806: inst = 32'h5be00000;
      42807: inst = 32'h8c50000;
      42808: inst = 32'h24612800;
      42809: inst = 32'h10a0ffff;
      42810: inst = 32'hca0ffe5;
      42811: inst = 32'h24822800;
      42812: inst = 32'h10a00000;
      42813: inst = 32'hca00004;
      42814: inst = 32'h38632800;
      42815: inst = 32'h38842800;
      42816: inst = 32'h10a00000;
      42817: inst = 32'hca0a745;
      42818: inst = 32'h13e00001;
      42819: inst = 32'hfe0d96a;
      42820: inst = 32'h5be00000;
      42821: inst = 32'h8c50000;
      42822: inst = 32'h24612800;
      42823: inst = 32'h10a0ffff;
      42824: inst = 32'hca0ffe5;
      42825: inst = 32'h24822800;
      42826: inst = 32'h10a00000;
      42827: inst = 32'hca00004;
      42828: inst = 32'h38632800;
      42829: inst = 32'h38842800;
      42830: inst = 32'h10a00000;
      42831: inst = 32'hca0a753;
      42832: inst = 32'h13e00001;
      42833: inst = 32'hfe0d96a;
      42834: inst = 32'h5be00000;
      42835: inst = 32'h8c50000;
      42836: inst = 32'h24612800;
      42837: inst = 32'h10a0ffff;
      42838: inst = 32'hca0ffe5;
      42839: inst = 32'h24822800;
      42840: inst = 32'h10a00000;
      42841: inst = 32'hca00004;
      42842: inst = 32'h38632800;
      42843: inst = 32'h38842800;
      42844: inst = 32'h10a00000;
      42845: inst = 32'hca0a761;
      42846: inst = 32'h13e00001;
      42847: inst = 32'hfe0d96a;
      42848: inst = 32'h5be00000;
      42849: inst = 32'h8c50000;
      42850: inst = 32'h24612800;
      42851: inst = 32'h10a0ffff;
      42852: inst = 32'hca0ffe5;
      42853: inst = 32'h24822800;
      42854: inst = 32'h10a00000;
      42855: inst = 32'hca00004;
      42856: inst = 32'h38632800;
      42857: inst = 32'h38842800;
      42858: inst = 32'h10a00000;
      42859: inst = 32'hca0a76f;
      42860: inst = 32'h13e00001;
      42861: inst = 32'hfe0d96a;
      42862: inst = 32'h5be00000;
      42863: inst = 32'h8c50000;
      42864: inst = 32'h24612800;
      42865: inst = 32'h10a0ffff;
      42866: inst = 32'hca0ffe5;
      42867: inst = 32'h24822800;
      42868: inst = 32'h10a00000;
      42869: inst = 32'hca00004;
      42870: inst = 32'h38632800;
      42871: inst = 32'h38842800;
      42872: inst = 32'h10a00000;
      42873: inst = 32'hca0a77d;
      42874: inst = 32'h13e00001;
      42875: inst = 32'hfe0d96a;
      42876: inst = 32'h5be00000;
      42877: inst = 32'h8c50000;
      42878: inst = 32'h24612800;
      42879: inst = 32'h10a0ffff;
      42880: inst = 32'hca0ffe5;
      42881: inst = 32'h24822800;
      42882: inst = 32'h10a00000;
      42883: inst = 32'hca00004;
      42884: inst = 32'h38632800;
      42885: inst = 32'h38842800;
      42886: inst = 32'h10a00000;
      42887: inst = 32'hca0a78b;
      42888: inst = 32'h13e00001;
      42889: inst = 32'hfe0d96a;
      42890: inst = 32'h5be00000;
      42891: inst = 32'h8c50000;
      42892: inst = 32'h24612800;
      42893: inst = 32'h10a0ffff;
      42894: inst = 32'hca0ffe5;
      42895: inst = 32'h24822800;
      42896: inst = 32'h10a00000;
      42897: inst = 32'hca00004;
      42898: inst = 32'h38632800;
      42899: inst = 32'h38842800;
      42900: inst = 32'h10a00000;
      42901: inst = 32'hca0a799;
      42902: inst = 32'h13e00001;
      42903: inst = 32'hfe0d96a;
      42904: inst = 32'h5be00000;
      42905: inst = 32'h8c50000;
      42906: inst = 32'h24612800;
      42907: inst = 32'h10a0ffff;
      42908: inst = 32'hca0ffe5;
      42909: inst = 32'h24822800;
      42910: inst = 32'h10a00000;
      42911: inst = 32'hca00004;
      42912: inst = 32'h38632800;
      42913: inst = 32'h38842800;
      42914: inst = 32'h10a00000;
      42915: inst = 32'hca0a7a7;
      42916: inst = 32'h13e00001;
      42917: inst = 32'hfe0d96a;
      42918: inst = 32'h5be00000;
      42919: inst = 32'h8c50000;
      42920: inst = 32'h24612800;
      42921: inst = 32'h10a0ffff;
      42922: inst = 32'hca0ffe5;
      42923: inst = 32'h24822800;
      42924: inst = 32'h10a00000;
      42925: inst = 32'hca00004;
      42926: inst = 32'h38632800;
      42927: inst = 32'h38842800;
      42928: inst = 32'h10a00000;
      42929: inst = 32'hca0a7b5;
      42930: inst = 32'h13e00001;
      42931: inst = 32'hfe0d96a;
      42932: inst = 32'h5be00000;
      42933: inst = 32'h8c50000;
      42934: inst = 32'h24612800;
      42935: inst = 32'h10a0ffff;
      42936: inst = 32'hca0ffe5;
      42937: inst = 32'h24822800;
      42938: inst = 32'h10a00000;
      42939: inst = 32'hca00004;
      42940: inst = 32'h38632800;
      42941: inst = 32'h38842800;
      42942: inst = 32'h10a00000;
      42943: inst = 32'hca0a7c3;
      42944: inst = 32'h13e00001;
      42945: inst = 32'hfe0d96a;
      42946: inst = 32'h5be00000;
      42947: inst = 32'h8c50000;
      42948: inst = 32'h24612800;
      42949: inst = 32'h10a0ffff;
      42950: inst = 32'hca0ffe5;
      42951: inst = 32'h24822800;
      42952: inst = 32'h10a00000;
      42953: inst = 32'hca00004;
      42954: inst = 32'h38632800;
      42955: inst = 32'h38842800;
      42956: inst = 32'h10a00000;
      42957: inst = 32'hca0a7d1;
      42958: inst = 32'h13e00001;
      42959: inst = 32'hfe0d96a;
      42960: inst = 32'h5be00000;
      42961: inst = 32'h8c50000;
      42962: inst = 32'h24612800;
      42963: inst = 32'h10a0ffff;
      42964: inst = 32'hca0ffe5;
      42965: inst = 32'h24822800;
      42966: inst = 32'h10a00000;
      42967: inst = 32'hca00004;
      42968: inst = 32'h38632800;
      42969: inst = 32'h38842800;
      42970: inst = 32'h10a00000;
      42971: inst = 32'hca0a7df;
      42972: inst = 32'h13e00001;
      42973: inst = 32'hfe0d96a;
      42974: inst = 32'h5be00000;
      42975: inst = 32'h8c50000;
      42976: inst = 32'h24612800;
      42977: inst = 32'h10a0ffff;
      42978: inst = 32'hca0ffe5;
      42979: inst = 32'h24822800;
      42980: inst = 32'h10a00000;
      42981: inst = 32'hca00004;
      42982: inst = 32'h38632800;
      42983: inst = 32'h38842800;
      42984: inst = 32'h10a00000;
      42985: inst = 32'hca0a7ed;
      42986: inst = 32'h13e00001;
      42987: inst = 32'hfe0d96a;
      42988: inst = 32'h5be00000;
      42989: inst = 32'h8c50000;
      42990: inst = 32'h24612800;
      42991: inst = 32'h10a0ffff;
      42992: inst = 32'hca0ffe5;
      42993: inst = 32'h24822800;
      42994: inst = 32'h10a00000;
      42995: inst = 32'hca00004;
      42996: inst = 32'h38632800;
      42997: inst = 32'h38842800;
      42998: inst = 32'h10a00000;
      42999: inst = 32'hca0a7fb;
      43000: inst = 32'h13e00001;
      43001: inst = 32'hfe0d96a;
      43002: inst = 32'h5be00000;
      43003: inst = 32'h8c50000;
      43004: inst = 32'h24612800;
      43005: inst = 32'h10a0ffff;
      43006: inst = 32'hca0ffe5;
      43007: inst = 32'h24822800;
      43008: inst = 32'h10a00000;
      43009: inst = 32'hca00004;
      43010: inst = 32'h38632800;
      43011: inst = 32'h38842800;
      43012: inst = 32'h10a00000;
      43013: inst = 32'hca0a809;
      43014: inst = 32'h13e00001;
      43015: inst = 32'hfe0d96a;
      43016: inst = 32'h5be00000;
      43017: inst = 32'h8c50000;
      43018: inst = 32'h24612800;
      43019: inst = 32'h10a0ffff;
      43020: inst = 32'hca0ffe5;
      43021: inst = 32'h24822800;
      43022: inst = 32'h10a00000;
      43023: inst = 32'hca00004;
      43024: inst = 32'h38632800;
      43025: inst = 32'h38842800;
      43026: inst = 32'h10a00000;
      43027: inst = 32'hca0a817;
      43028: inst = 32'h13e00001;
      43029: inst = 32'hfe0d96a;
      43030: inst = 32'h5be00000;
      43031: inst = 32'h8c50000;
      43032: inst = 32'h24612800;
      43033: inst = 32'h10a0ffff;
      43034: inst = 32'hca0ffe5;
      43035: inst = 32'h24822800;
      43036: inst = 32'h10a00000;
      43037: inst = 32'hca00004;
      43038: inst = 32'h38632800;
      43039: inst = 32'h38842800;
      43040: inst = 32'h10a00000;
      43041: inst = 32'hca0a825;
      43042: inst = 32'h13e00001;
      43043: inst = 32'hfe0d96a;
      43044: inst = 32'h5be00000;
      43045: inst = 32'h8c50000;
      43046: inst = 32'h24612800;
      43047: inst = 32'h10a0ffff;
      43048: inst = 32'hca0ffe5;
      43049: inst = 32'h24822800;
      43050: inst = 32'h10a00000;
      43051: inst = 32'hca00004;
      43052: inst = 32'h38632800;
      43053: inst = 32'h38842800;
      43054: inst = 32'h10a00000;
      43055: inst = 32'hca0a833;
      43056: inst = 32'h13e00001;
      43057: inst = 32'hfe0d96a;
      43058: inst = 32'h5be00000;
      43059: inst = 32'h8c50000;
      43060: inst = 32'h24612800;
      43061: inst = 32'h10a0ffff;
      43062: inst = 32'hca0ffe5;
      43063: inst = 32'h24822800;
      43064: inst = 32'h10a00000;
      43065: inst = 32'hca00004;
      43066: inst = 32'h38632800;
      43067: inst = 32'h38842800;
      43068: inst = 32'h10a00000;
      43069: inst = 32'hca0a841;
      43070: inst = 32'h13e00001;
      43071: inst = 32'hfe0d96a;
      43072: inst = 32'h5be00000;
      43073: inst = 32'h8c50000;
      43074: inst = 32'h24612800;
      43075: inst = 32'h10a0ffff;
      43076: inst = 32'hca0ffe5;
      43077: inst = 32'h24822800;
      43078: inst = 32'h10a00000;
      43079: inst = 32'hca00004;
      43080: inst = 32'h38632800;
      43081: inst = 32'h38842800;
      43082: inst = 32'h10a00000;
      43083: inst = 32'hca0a84f;
      43084: inst = 32'h13e00001;
      43085: inst = 32'hfe0d96a;
      43086: inst = 32'h5be00000;
      43087: inst = 32'h8c50000;
      43088: inst = 32'h24612800;
      43089: inst = 32'h10a0ffff;
      43090: inst = 32'hca0ffe5;
      43091: inst = 32'h24822800;
      43092: inst = 32'h10a00000;
      43093: inst = 32'hca00004;
      43094: inst = 32'h38632800;
      43095: inst = 32'h38842800;
      43096: inst = 32'h10a00000;
      43097: inst = 32'hca0a85d;
      43098: inst = 32'h13e00001;
      43099: inst = 32'hfe0d96a;
      43100: inst = 32'h5be00000;
      43101: inst = 32'h8c50000;
      43102: inst = 32'h24612800;
      43103: inst = 32'h10a0ffff;
      43104: inst = 32'hca0ffe5;
      43105: inst = 32'h24822800;
      43106: inst = 32'h10a00000;
      43107: inst = 32'hca00004;
      43108: inst = 32'h38632800;
      43109: inst = 32'h38842800;
      43110: inst = 32'h10a00000;
      43111: inst = 32'hca0a86b;
      43112: inst = 32'h13e00001;
      43113: inst = 32'hfe0d96a;
      43114: inst = 32'h5be00000;
      43115: inst = 32'h8c50000;
      43116: inst = 32'h24612800;
      43117: inst = 32'h10a0ffff;
      43118: inst = 32'hca0ffe5;
      43119: inst = 32'h24822800;
      43120: inst = 32'h10a00000;
      43121: inst = 32'hca00004;
      43122: inst = 32'h38632800;
      43123: inst = 32'h38842800;
      43124: inst = 32'h10a00000;
      43125: inst = 32'hca0a879;
      43126: inst = 32'h13e00001;
      43127: inst = 32'hfe0d96a;
      43128: inst = 32'h5be00000;
      43129: inst = 32'h8c50000;
      43130: inst = 32'h24612800;
      43131: inst = 32'h10a0ffff;
      43132: inst = 32'hca0ffe5;
      43133: inst = 32'h24822800;
      43134: inst = 32'h10a00000;
      43135: inst = 32'hca00004;
      43136: inst = 32'h38632800;
      43137: inst = 32'h38842800;
      43138: inst = 32'h10a00000;
      43139: inst = 32'hca0a887;
      43140: inst = 32'h13e00001;
      43141: inst = 32'hfe0d96a;
      43142: inst = 32'h5be00000;
      43143: inst = 32'h8c50000;
      43144: inst = 32'h24612800;
      43145: inst = 32'h10a0ffff;
      43146: inst = 32'hca0ffe5;
      43147: inst = 32'h24822800;
      43148: inst = 32'h10a00000;
      43149: inst = 32'hca00004;
      43150: inst = 32'h38632800;
      43151: inst = 32'h38842800;
      43152: inst = 32'h10a00000;
      43153: inst = 32'hca0a895;
      43154: inst = 32'h13e00001;
      43155: inst = 32'hfe0d96a;
      43156: inst = 32'h5be00000;
      43157: inst = 32'h8c50000;
      43158: inst = 32'h24612800;
      43159: inst = 32'h10a0ffff;
      43160: inst = 32'hca0ffe5;
      43161: inst = 32'h24822800;
      43162: inst = 32'h10a00000;
      43163: inst = 32'hca00004;
      43164: inst = 32'h38632800;
      43165: inst = 32'h38842800;
      43166: inst = 32'h10a00000;
      43167: inst = 32'hca0a8a3;
      43168: inst = 32'h13e00001;
      43169: inst = 32'hfe0d96a;
      43170: inst = 32'h5be00000;
      43171: inst = 32'h8c50000;
      43172: inst = 32'h24612800;
      43173: inst = 32'h10a0ffff;
      43174: inst = 32'hca0ffe5;
      43175: inst = 32'h24822800;
      43176: inst = 32'h10a00000;
      43177: inst = 32'hca00004;
      43178: inst = 32'h38632800;
      43179: inst = 32'h38842800;
      43180: inst = 32'h10a00000;
      43181: inst = 32'hca0a8b1;
      43182: inst = 32'h13e00001;
      43183: inst = 32'hfe0d96a;
      43184: inst = 32'h5be00000;
      43185: inst = 32'h8c50000;
      43186: inst = 32'h24612800;
      43187: inst = 32'h10a0ffff;
      43188: inst = 32'hca0ffe5;
      43189: inst = 32'h24822800;
      43190: inst = 32'h10a00000;
      43191: inst = 32'hca00004;
      43192: inst = 32'h38632800;
      43193: inst = 32'h38842800;
      43194: inst = 32'h10a00000;
      43195: inst = 32'hca0a8bf;
      43196: inst = 32'h13e00001;
      43197: inst = 32'hfe0d96a;
      43198: inst = 32'h5be00000;
      43199: inst = 32'h8c50000;
      43200: inst = 32'h24612800;
      43201: inst = 32'h10a0ffff;
      43202: inst = 32'hca0ffe5;
      43203: inst = 32'h24822800;
      43204: inst = 32'h10a00000;
      43205: inst = 32'hca00004;
      43206: inst = 32'h38632800;
      43207: inst = 32'h38842800;
      43208: inst = 32'h10a00000;
      43209: inst = 32'hca0a8cd;
      43210: inst = 32'h13e00001;
      43211: inst = 32'hfe0d96a;
      43212: inst = 32'h5be00000;
      43213: inst = 32'h8c50000;
      43214: inst = 32'h24612800;
      43215: inst = 32'h10a0ffff;
      43216: inst = 32'hca0ffe5;
      43217: inst = 32'h24822800;
      43218: inst = 32'h10a00000;
      43219: inst = 32'hca00004;
      43220: inst = 32'h38632800;
      43221: inst = 32'h38842800;
      43222: inst = 32'h10a00000;
      43223: inst = 32'hca0a8db;
      43224: inst = 32'h13e00001;
      43225: inst = 32'hfe0d96a;
      43226: inst = 32'h5be00000;
      43227: inst = 32'h8c50000;
      43228: inst = 32'h24612800;
      43229: inst = 32'h10a0ffff;
      43230: inst = 32'hca0ffe5;
      43231: inst = 32'h24822800;
      43232: inst = 32'h10a00000;
      43233: inst = 32'hca00004;
      43234: inst = 32'h38632800;
      43235: inst = 32'h38842800;
      43236: inst = 32'h10a00000;
      43237: inst = 32'hca0a8e9;
      43238: inst = 32'h13e00001;
      43239: inst = 32'hfe0d96a;
      43240: inst = 32'h5be00000;
      43241: inst = 32'h8c50000;
      43242: inst = 32'h24612800;
      43243: inst = 32'h10a0ffff;
      43244: inst = 32'hca0ffe6;
      43245: inst = 32'h24822800;
      43246: inst = 32'h10a00000;
      43247: inst = 32'hca00004;
      43248: inst = 32'h38632800;
      43249: inst = 32'h38842800;
      43250: inst = 32'h10a00000;
      43251: inst = 32'hca0a8f7;
      43252: inst = 32'h13e00001;
      43253: inst = 32'hfe0d96a;
      43254: inst = 32'h5be00000;
      43255: inst = 32'h8c50000;
      43256: inst = 32'h24612800;
      43257: inst = 32'h10a0ffff;
      43258: inst = 32'hca0ffe6;
      43259: inst = 32'h24822800;
      43260: inst = 32'h10a00000;
      43261: inst = 32'hca00004;
      43262: inst = 32'h38632800;
      43263: inst = 32'h38842800;
      43264: inst = 32'h10a00000;
      43265: inst = 32'hca0a905;
      43266: inst = 32'h13e00001;
      43267: inst = 32'hfe0d96a;
      43268: inst = 32'h5be00000;
      43269: inst = 32'h8c50000;
      43270: inst = 32'h24612800;
      43271: inst = 32'h10a0ffff;
      43272: inst = 32'hca0ffe6;
      43273: inst = 32'h24822800;
      43274: inst = 32'h10a00000;
      43275: inst = 32'hca00004;
      43276: inst = 32'h38632800;
      43277: inst = 32'h38842800;
      43278: inst = 32'h10a00000;
      43279: inst = 32'hca0a913;
      43280: inst = 32'h13e00001;
      43281: inst = 32'hfe0d96a;
      43282: inst = 32'h5be00000;
      43283: inst = 32'h8c50000;
      43284: inst = 32'h24612800;
      43285: inst = 32'h10a0ffff;
      43286: inst = 32'hca0ffe6;
      43287: inst = 32'h24822800;
      43288: inst = 32'h10a00000;
      43289: inst = 32'hca00004;
      43290: inst = 32'h38632800;
      43291: inst = 32'h38842800;
      43292: inst = 32'h10a00000;
      43293: inst = 32'hca0a921;
      43294: inst = 32'h13e00001;
      43295: inst = 32'hfe0d96a;
      43296: inst = 32'h5be00000;
      43297: inst = 32'h8c50000;
      43298: inst = 32'h24612800;
      43299: inst = 32'h10a0ffff;
      43300: inst = 32'hca0ffe6;
      43301: inst = 32'h24822800;
      43302: inst = 32'h10a00000;
      43303: inst = 32'hca00004;
      43304: inst = 32'h38632800;
      43305: inst = 32'h38842800;
      43306: inst = 32'h10a00000;
      43307: inst = 32'hca0a92f;
      43308: inst = 32'h13e00001;
      43309: inst = 32'hfe0d96a;
      43310: inst = 32'h5be00000;
      43311: inst = 32'h8c50000;
      43312: inst = 32'h24612800;
      43313: inst = 32'h10a0ffff;
      43314: inst = 32'hca0ffe6;
      43315: inst = 32'h24822800;
      43316: inst = 32'h10a00000;
      43317: inst = 32'hca00004;
      43318: inst = 32'h38632800;
      43319: inst = 32'h38842800;
      43320: inst = 32'h10a00000;
      43321: inst = 32'hca0a93d;
      43322: inst = 32'h13e00001;
      43323: inst = 32'hfe0d96a;
      43324: inst = 32'h5be00000;
      43325: inst = 32'h8c50000;
      43326: inst = 32'h24612800;
      43327: inst = 32'h10a0ffff;
      43328: inst = 32'hca0ffe6;
      43329: inst = 32'h24822800;
      43330: inst = 32'h10a00000;
      43331: inst = 32'hca00004;
      43332: inst = 32'h38632800;
      43333: inst = 32'h38842800;
      43334: inst = 32'h10a00000;
      43335: inst = 32'hca0a94b;
      43336: inst = 32'h13e00001;
      43337: inst = 32'hfe0d96a;
      43338: inst = 32'h5be00000;
      43339: inst = 32'h8c50000;
      43340: inst = 32'h24612800;
      43341: inst = 32'h10a0ffff;
      43342: inst = 32'hca0ffe6;
      43343: inst = 32'h24822800;
      43344: inst = 32'h10a00000;
      43345: inst = 32'hca00004;
      43346: inst = 32'h38632800;
      43347: inst = 32'h38842800;
      43348: inst = 32'h10a00000;
      43349: inst = 32'hca0a959;
      43350: inst = 32'h13e00001;
      43351: inst = 32'hfe0d96a;
      43352: inst = 32'h5be00000;
      43353: inst = 32'h8c50000;
      43354: inst = 32'h24612800;
      43355: inst = 32'h10a0ffff;
      43356: inst = 32'hca0ffe6;
      43357: inst = 32'h24822800;
      43358: inst = 32'h10a00000;
      43359: inst = 32'hca00004;
      43360: inst = 32'h38632800;
      43361: inst = 32'h38842800;
      43362: inst = 32'h10a00000;
      43363: inst = 32'hca0a967;
      43364: inst = 32'h13e00001;
      43365: inst = 32'hfe0d96a;
      43366: inst = 32'h5be00000;
      43367: inst = 32'h8c50000;
      43368: inst = 32'h24612800;
      43369: inst = 32'h10a0ffff;
      43370: inst = 32'hca0ffe6;
      43371: inst = 32'h24822800;
      43372: inst = 32'h10a00000;
      43373: inst = 32'hca00004;
      43374: inst = 32'h38632800;
      43375: inst = 32'h38842800;
      43376: inst = 32'h10a00000;
      43377: inst = 32'hca0a975;
      43378: inst = 32'h13e00001;
      43379: inst = 32'hfe0d96a;
      43380: inst = 32'h5be00000;
      43381: inst = 32'h8c50000;
      43382: inst = 32'h24612800;
      43383: inst = 32'h10a0ffff;
      43384: inst = 32'hca0ffe6;
      43385: inst = 32'h24822800;
      43386: inst = 32'h10a00000;
      43387: inst = 32'hca00004;
      43388: inst = 32'h38632800;
      43389: inst = 32'h38842800;
      43390: inst = 32'h10a00000;
      43391: inst = 32'hca0a983;
      43392: inst = 32'h13e00001;
      43393: inst = 32'hfe0d96a;
      43394: inst = 32'h5be00000;
      43395: inst = 32'h8c50000;
      43396: inst = 32'h24612800;
      43397: inst = 32'h10a0ffff;
      43398: inst = 32'hca0ffe6;
      43399: inst = 32'h24822800;
      43400: inst = 32'h10a00000;
      43401: inst = 32'hca00004;
      43402: inst = 32'h38632800;
      43403: inst = 32'h38842800;
      43404: inst = 32'h10a00000;
      43405: inst = 32'hca0a991;
      43406: inst = 32'h13e00001;
      43407: inst = 32'hfe0d96a;
      43408: inst = 32'h5be00000;
      43409: inst = 32'h8c50000;
      43410: inst = 32'h24612800;
      43411: inst = 32'h10a0ffff;
      43412: inst = 32'hca0ffe6;
      43413: inst = 32'h24822800;
      43414: inst = 32'h10a00000;
      43415: inst = 32'hca00004;
      43416: inst = 32'h38632800;
      43417: inst = 32'h38842800;
      43418: inst = 32'h10a00000;
      43419: inst = 32'hca0a99f;
      43420: inst = 32'h13e00001;
      43421: inst = 32'hfe0d96a;
      43422: inst = 32'h5be00000;
      43423: inst = 32'h8c50000;
      43424: inst = 32'h24612800;
      43425: inst = 32'h10a0ffff;
      43426: inst = 32'hca0ffe6;
      43427: inst = 32'h24822800;
      43428: inst = 32'h10a00000;
      43429: inst = 32'hca00004;
      43430: inst = 32'h38632800;
      43431: inst = 32'h38842800;
      43432: inst = 32'h10a00000;
      43433: inst = 32'hca0a9ad;
      43434: inst = 32'h13e00001;
      43435: inst = 32'hfe0d96a;
      43436: inst = 32'h5be00000;
      43437: inst = 32'h8c50000;
      43438: inst = 32'h24612800;
      43439: inst = 32'h10a0ffff;
      43440: inst = 32'hca0ffe6;
      43441: inst = 32'h24822800;
      43442: inst = 32'h10a00000;
      43443: inst = 32'hca00004;
      43444: inst = 32'h38632800;
      43445: inst = 32'h38842800;
      43446: inst = 32'h10a00000;
      43447: inst = 32'hca0a9bb;
      43448: inst = 32'h13e00001;
      43449: inst = 32'hfe0d96a;
      43450: inst = 32'h5be00000;
      43451: inst = 32'h8c50000;
      43452: inst = 32'h24612800;
      43453: inst = 32'h10a0ffff;
      43454: inst = 32'hca0ffe6;
      43455: inst = 32'h24822800;
      43456: inst = 32'h10a00000;
      43457: inst = 32'hca00004;
      43458: inst = 32'h38632800;
      43459: inst = 32'h38842800;
      43460: inst = 32'h10a00000;
      43461: inst = 32'hca0a9c9;
      43462: inst = 32'h13e00001;
      43463: inst = 32'hfe0d96a;
      43464: inst = 32'h5be00000;
      43465: inst = 32'h8c50000;
      43466: inst = 32'h24612800;
      43467: inst = 32'h10a0ffff;
      43468: inst = 32'hca0ffe6;
      43469: inst = 32'h24822800;
      43470: inst = 32'h10a00000;
      43471: inst = 32'hca00004;
      43472: inst = 32'h38632800;
      43473: inst = 32'h38842800;
      43474: inst = 32'h10a00000;
      43475: inst = 32'hca0a9d7;
      43476: inst = 32'h13e00001;
      43477: inst = 32'hfe0d96a;
      43478: inst = 32'h5be00000;
      43479: inst = 32'h8c50000;
      43480: inst = 32'h24612800;
      43481: inst = 32'h10a0ffff;
      43482: inst = 32'hca0ffe6;
      43483: inst = 32'h24822800;
      43484: inst = 32'h10a00000;
      43485: inst = 32'hca00004;
      43486: inst = 32'h38632800;
      43487: inst = 32'h38842800;
      43488: inst = 32'h10a00000;
      43489: inst = 32'hca0a9e5;
      43490: inst = 32'h13e00001;
      43491: inst = 32'hfe0d96a;
      43492: inst = 32'h5be00000;
      43493: inst = 32'h8c50000;
      43494: inst = 32'h24612800;
      43495: inst = 32'h10a0ffff;
      43496: inst = 32'hca0ffe6;
      43497: inst = 32'h24822800;
      43498: inst = 32'h10a00000;
      43499: inst = 32'hca00004;
      43500: inst = 32'h38632800;
      43501: inst = 32'h38842800;
      43502: inst = 32'h10a00000;
      43503: inst = 32'hca0a9f3;
      43504: inst = 32'h13e00001;
      43505: inst = 32'hfe0d96a;
      43506: inst = 32'h5be00000;
      43507: inst = 32'h8c50000;
      43508: inst = 32'h24612800;
      43509: inst = 32'h10a0ffff;
      43510: inst = 32'hca0ffe6;
      43511: inst = 32'h24822800;
      43512: inst = 32'h10a00000;
      43513: inst = 32'hca00004;
      43514: inst = 32'h38632800;
      43515: inst = 32'h38842800;
      43516: inst = 32'h10a00000;
      43517: inst = 32'hca0aa01;
      43518: inst = 32'h13e00001;
      43519: inst = 32'hfe0d96a;
      43520: inst = 32'h5be00000;
      43521: inst = 32'h8c50000;
      43522: inst = 32'h24612800;
      43523: inst = 32'h10a0ffff;
      43524: inst = 32'hca0ffe6;
      43525: inst = 32'h24822800;
      43526: inst = 32'h10a00000;
      43527: inst = 32'hca00004;
      43528: inst = 32'h38632800;
      43529: inst = 32'h38842800;
      43530: inst = 32'h10a00000;
      43531: inst = 32'hca0aa0f;
      43532: inst = 32'h13e00001;
      43533: inst = 32'hfe0d96a;
      43534: inst = 32'h5be00000;
      43535: inst = 32'h8c50000;
      43536: inst = 32'h24612800;
      43537: inst = 32'h10a0ffff;
      43538: inst = 32'hca0ffe6;
      43539: inst = 32'h24822800;
      43540: inst = 32'h10a00000;
      43541: inst = 32'hca00004;
      43542: inst = 32'h38632800;
      43543: inst = 32'h38842800;
      43544: inst = 32'h10a00000;
      43545: inst = 32'hca0aa1d;
      43546: inst = 32'h13e00001;
      43547: inst = 32'hfe0d96a;
      43548: inst = 32'h5be00000;
      43549: inst = 32'h8c50000;
      43550: inst = 32'h24612800;
      43551: inst = 32'h10a0ffff;
      43552: inst = 32'hca0ffe6;
      43553: inst = 32'h24822800;
      43554: inst = 32'h10a00000;
      43555: inst = 32'hca00004;
      43556: inst = 32'h38632800;
      43557: inst = 32'h38842800;
      43558: inst = 32'h10a00000;
      43559: inst = 32'hca0aa2b;
      43560: inst = 32'h13e00001;
      43561: inst = 32'hfe0d96a;
      43562: inst = 32'h5be00000;
      43563: inst = 32'h8c50000;
      43564: inst = 32'h24612800;
      43565: inst = 32'h10a0ffff;
      43566: inst = 32'hca0ffe6;
      43567: inst = 32'h24822800;
      43568: inst = 32'h10a00000;
      43569: inst = 32'hca00004;
      43570: inst = 32'h38632800;
      43571: inst = 32'h38842800;
      43572: inst = 32'h10a00000;
      43573: inst = 32'hca0aa39;
      43574: inst = 32'h13e00001;
      43575: inst = 32'hfe0d96a;
      43576: inst = 32'h5be00000;
      43577: inst = 32'h8c50000;
      43578: inst = 32'h24612800;
      43579: inst = 32'h10a0ffff;
      43580: inst = 32'hca0ffe6;
      43581: inst = 32'h24822800;
      43582: inst = 32'h10a00000;
      43583: inst = 32'hca00004;
      43584: inst = 32'h38632800;
      43585: inst = 32'h38842800;
      43586: inst = 32'h10a00000;
      43587: inst = 32'hca0aa47;
      43588: inst = 32'h13e00001;
      43589: inst = 32'hfe0d96a;
      43590: inst = 32'h5be00000;
      43591: inst = 32'h8c50000;
      43592: inst = 32'h24612800;
      43593: inst = 32'h10a0ffff;
      43594: inst = 32'hca0ffe6;
      43595: inst = 32'h24822800;
      43596: inst = 32'h10a00000;
      43597: inst = 32'hca00004;
      43598: inst = 32'h38632800;
      43599: inst = 32'h38842800;
      43600: inst = 32'h10a00000;
      43601: inst = 32'hca0aa55;
      43602: inst = 32'h13e00001;
      43603: inst = 32'hfe0d96a;
      43604: inst = 32'h5be00000;
      43605: inst = 32'h8c50000;
      43606: inst = 32'h24612800;
      43607: inst = 32'h10a0ffff;
      43608: inst = 32'hca0ffe6;
      43609: inst = 32'h24822800;
      43610: inst = 32'h10a00000;
      43611: inst = 32'hca00004;
      43612: inst = 32'h38632800;
      43613: inst = 32'h38842800;
      43614: inst = 32'h10a00000;
      43615: inst = 32'hca0aa63;
      43616: inst = 32'h13e00001;
      43617: inst = 32'hfe0d96a;
      43618: inst = 32'h5be00000;
      43619: inst = 32'h8c50000;
      43620: inst = 32'h24612800;
      43621: inst = 32'h10a0ffff;
      43622: inst = 32'hca0ffe6;
      43623: inst = 32'h24822800;
      43624: inst = 32'h10a00000;
      43625: inst = 32'hca00004;
      43626: inst = 32'h38632800;
      43627: inst = 32'h38842800;
      43628: inst = 32'h10a00000;
      43629: inst = 32'hca0aa71;
      43630: inst = 32'h13e00001;
      43631: inst = 32'hfe0d96a;
      43632: inst = 32'h5be00000;
      43633: inst = 32'h8c50000;
      43634: inst = 32'h24612800;
      43635: inst = 32'h10a0ffff;
      43636: inst = 32'hca0ffe6;
      43637: inst = 32'h24822800;
      43638: inst = 32'h10a00000;
      43639: inst = 32'hca00004;
      43640: inst = 32'h38632800;
      43641: inst = 32'h38842800;
      43642: inst = 32'h10a00000;
      43643: inst = 32'hca0aa7f;
      43644: inst = 32'h13e00001;
      43645: inst = 32'hfe0d96a;
      43646: inst = 32'h5be00000;
      43647: inst = 32'h8c50000;
      43648: inst = 32'h24612800;
      43649: inst = 32'h10a0ffff;
      43650: inst = 32'hca0ffe6;
      43651: inst = 32'h24822800;
      43652: inst = 32'h10a00000;
      43653: inst = 32'hca00004;
      43654: inst = 32'h38632800;
      43655: inst = 32'h38842800;
      43656: inst = 32'h10a00000;
      43657: inst = 32'hca0aa8d;
      43658: inst = 32'h13e00001;
      43659: inst = 32'hfe0d96a;
      43660: inst = 32'h5be00000;
      43661: inst = 32'h8c50000;
      43662: inst = 32'h24612800;
      43663: inst = 32'h10a0ffff;
      43664: inst = 32'hca0ffe6;
      43665: inst = 32'h24822800;
      43666: inst = 32'h10a00000;
      43667: inst = 32'hca00004;
      43668: inst = 32'h38632800;
      43669: inst = 32'h38842800;
      43670: inst = 32'h10a00000;
      43671: inst = 32'hca0aa9b;
      43672: inst = 32'h13e00001;
      43673: inst = 32'hfe0d96a;
      43674: inst = 32'h5be00000;
      43675: inst = 32'h8c50000;
      43676: inst = 32'h24612800;
      43677: inst = 32'h10a0ffff;
      43678: inst = 32'hca0ffe6;
      43679: inst = 32'h24822800;
      43680: inst = 32'h10a00000;
      43681: inst = 32'hca00004;
      43682: inst = 32'h38632800;
      43683: inst = 32'h38842800;
      43684: inst = 32'h10a00000;
      43685: inst = 32'hca0aaa9;
      43686: inst = 32'h13e00001;
      43687: inst = 32'hfe0d96a;
      43688: inst = 32'h5be00000;
      43689: inst = 32'h8c50000;
      43690: inst = 32'h24612800;
      43691: inst = 32'h10a0ffff;
      43692: inst = 32'hca0ffe6;
      43693: inst = 32'h24822800;
      43694: inst = 32'h10a00000;
      43695: inst = 32'hca00004;
      43696: inst = 32'h38632800;
      43697: inst = 32'h38842800;
      43698: inst = 32'h10a00000;
      43699: inst = 32'hca0aab7;
      43700: inst = 32'h13e00001;
      43701: inst = 32'hfe0d96a;
      43702: inst = 32'h5be00000;
      43703: inst = 32'h8c50000;
      43704: inst = 32'h24612800;
      43705: inst = 32'h10a0ffff;
      43706: inst = 32'hca0ffe6;
      43707: inst = 32'h24822800;
      43708: inst = 32'h10a00000;
      43709: inst = 32'hca00004;
      43710: inst = 32'h38632800;
      43711: inst = 32'h38842800;
      43712: inst = 32'h10a00000;
      43713: inst = 32'hca0aac5;
      43714: inst = 32'h13e00001;
      43715: inst = 32'hfe0d96a;
      43716: inst = 32'h5be00000;
      43717: inst = 32'h8c50000;
      43718: inst = 32'h24612800;
      43719: inst = 32'h10a0ffff;
      43720: inst = 32'hca0ffe6;
      43721: inst = 32'h24822800;
      43722: inst = 32'h10a00000;
      43723: inst = 32'hca00004;
      43724: inst = 32'h38632800;
      43725: inst = 32'h38842800;
      43726: inst = 32'h10a00000;
      43727: inst = 32'hca0aad3;
      43728: inst = 32'h13e00001;
      43729: inst = 32'hfe0d96a;
      43730: inst = 32'h5be00000;
      43731: inst = 32'h8c50000;
      43732: inst = 32'h24612800;
      43733: inst = 32'h10a0ffff;
      43734: inst = 32'hca0ffe6;
      43735: inst = 32'h24822800;
      43736: inst = 32'h10a00000;
      43737: inst = 32'hca00004;
      43738: inst = 32'h38632800;
      43739: inst = 32'h38842800;
      43740: inst = 32'h10a00000;
      43741: inst = 32'hca0aae1;
      43742: inst = 32'h13e00001;
      43743: inst = 32'hfe0d96a;
      43744: inst = 32'h5be00000;
      43745: inst = 32'h8c50000;
      43746: inst = 32'h24612800;
      43747: inst = 32'h10a0ffff;
      43748: inst = 32'hca0ffe6;
      43749: inst = 32'h24822800;
      43750: inst = 32'h10a00000;
      43751: inst = 32'hca00004;
      43752: inst = 32'h38632800;
      43753: inst = 32'h38842800;
      43754: inst = 32'h10a00000;
      43755: inst = 32'hca0aaef;
      43756: inst = 32'h13e00001;
      43757: inst = 32'hfe0d96a;
      43758: inst = 32'h5be00000;
      43759: inst = 32'h8c50000;
      43760: inst = 32'h24612800;
      43761: inst = 32'h10a0ffff;
      43762: inst = 32'hca0ffe6;
      43763: inst = 32'h24822800;
      43764: inst = 32'h10a00000;
      43765: inst = 32'hca00004;
      43766: inst = 32'h38632800;
      43767: inst = 32'h38842800;
      43768: inst = 32'h10a00000;
      43769: inst = 32'hca0aafd;
      43770: inst = 32'h13e00001;
      43771: inst = 32'hfe0d96a;
      43772: inst = 32'h5be00000;
      43773: inst = 32'h8c50000;
      43774: inst = 32'h24612800;
      43775: inst = 32'h10a0ffff;
      43776: inst = 32'hca0ffe6;
      43777: inst = 32'h24822800;
      43778: inst = 32'h10a00000;
      43779: inst = 32'hca00004;
      43780: inst = 32'h38632800;
      43781: inst = 32'h38842800;
      43782: inst = 32'h10a00000;
      43783: inst = 32'hca0ab0b;
      43784: inst = 32'h13e00001;
      43785: inst = 32'hfe0d96a;
      43786: inst = 32'h5be00000;
      43787: inst = 32'h8c50000;
      43788: inst = 32'h24612800;
      43789: inst = 32'h10a0ffff;
      43790: inst = 32'hca0ffe6;
      43791: inst = 32'h24822800;
      43792: inst = 32'h10a00000;
      43793: inst = 32'hca00004;
      43794: inst = 32'h38632800;
      43795: inst = 32'h38842800;
      43796: inst = 32'h10a00000;
      43797: inst = 32'hca0ab19;
      43798: inst = 32'h13e00001;
      43799: inst = 32'hfe0d96a;
      43800: inst = 32'h5be00000;
      43801: inst = 32'h8c50000;
      43802: inst = 32'h24612800;
      43803: inst = 32'h10a0ffff;
      43804: inst = 32'hca0ffe6;
      43805: inst = 32'h24822800;
      43806: inst = 32'h10a00000;
      43807: inst = 32'hca00004;
      43808: inst = 32'h38632800;
      43809: inst = 32'h38842800;
      43810: inst = 32'h10a00000;
      43811: inst = 32'hca0ab27;
      43812: inst = 32'h13e00001;
      43813: inst = 32'hfe0d96a;
      43814: inst = 32'h5be00000;
      43815: inst = 32'h8c50000;
      43816: inst = 32'h24612800;
      43817: inst = 32'h10a0ffff;
      43818: inst = 32'hca0ffe6;
      43819: inst = 32'h24822800;
      43820: inst = 32'h10a00000;
      43821: inst = 32'hca00004;
      43822: inst = 32'h38632800;
      43823: inst = 32'h38842800;
      43824: inst = 32'h10a00000;
      43825: inst = 32'hca0ab35;
      43826: inst = 32'h13e00001;
      43827: inst = 32'hfe0d96a;
      43828: inst = 32'h5be00000;
      43829: inst = 32'h8c50000;
      43830: inst = 32'h24612800;
      43831: inst = 32'h10a0ffff;
      43832: inst = 32'hca0ffe6;
      43833: inst = 32'h24822800;
      43834: inst = 32'h10a00000;
      43835: inst = 32'hca00004;
      43836: inst = 32'h38632800;
      43837: inst = 32'h38842800;
      43838: inst = 32'h10a00000;
      43839: inst = 32'hca0ab43;
      43840: inst = 32'h13e00001;
      43841: inst = 32'hfe0d96a;
      43842: inst = 32'h5be00000;
      43843: inst = 32'h8c50000;
      43844: inst = 32'h24612800;
      43845: inst = 32'h10a0ffff;
      43846: inst = 32'hca0ffe6;
      43847: inst = 32'h24822800;
      43848: inst = 32'h10a00000;
      43849: inst = 32'hca00004;
      43850: inst = 32'h38632800;
      43851: inst = 32'h38842800;
      43852: inst = 32'h10a00000;
      43853: inst = 32'hca0ab51;
      43854: inst = 32'h13e00001;
      43855: inst = 32'hfe0d96a;
      43856: inst = 32'h5be00000;
      43857: inst = 32'h8c50000;
      43858: inst = 32'h24612800;
      43859: inst = 32'h10a0ffff;
      43860: inst = 32'hca0ffe6;
      43861: inst = 32'h24822800;
      43862: inst = 32'h10a00000;
      43863: inst = 32'hca00004;
      43864: inst = 32'h38632800;
      43865: inst = 32'h38842800;
      43866: inst = 32'h10a00000;
      43867: inst = 32'hca0ab5f;
      43868: inst = 32'h13e00001;
      43869: inst = 32'hfe0d96a;
      43870: inst = 32'h5be00000;
      43871: inst = 32'h8c50000;
      43872: inst = 32'h24612800;
      43873: inst = 32'h10a0ffff;
      43874: inst = 32'hca0ffe6;
      43875: inst = 32'h24822800;
      43876: inst = 32'h10a00000;
      43877: inst = 32'hca00004;
      43878: inst = 32'h38632800;
      43879: inst = 32'h38842800;
      43880: inst = 32'h10a00000;
      43881: inst = 32'hca0ab6d;
      43882: inst = 32'h13e00001;
      43883: inst = 32'hfe0d96a;
      43884: inst = 32'h5be00000;
      43885: inst = 32'h8c50000;
      43886: inst = 32'h24612800;
      43887: inst = 32'h10a0ffff;
      43888: inst = 32'hca0ffe6;
      43889: inst = 32'h24822800;
      43890: inst = 32'h10a00000;
      43891: inst = 32'hca00004;
      43892: inst = 32'h38632800;
      43893: inst = 32'h38842800;
      43894: inst = 32'h10a00000;
      43895: inst = 32'hca0ab7b;
      43896: inst = 32'h13e00001;
      43897: inst = 32'hfe0d96a;
      43898: inst = 32'h5be00000;
      43899: inst = 32'h8c50000;
      43900: inst = 32'h24612800;
      43901: inst = 32'h10a0ffff;
      43902: inst = 32'hca0ffe6;
      43903: inst = 32'h24822800;
      43904: inst = 32'h10a00000;
      43905: inst = 32'hca00004;
      43906: inst = 32'h38632800;
      43907: inst = 32'h38842800;
      43908: inst = 32'h10a00000;
      43909: inst = 32'hca0ab89;
      43910: inst = 32'h13e00001;
      43911: inst = 32'hfe0d96a;
      43912: inst = 32'h5be00000;
      43913: inst = 32'h8c50000;
      43914: inst = 32'h24612800;
      43915: inst = 32'h10a0ffff;
      43916: inst = 32'hca0ffe6;
      43917: inst = 32'h24822800;
      43918: inst = 32'h10a00000;
      43919: inst = 32'hca00004;
      43920: inst = 32'h38632800;
      43921: inst = 32'h38842800;
      43922: inst = 32'h10a00000;
      43923: inst = 32'hca0ab97;
      43924: inst = 32'h13e00001;
      43925: inst = 32'hfe0d96a;
      43926: inst = 32'h5be00000;
      43927: inst = 32'h8c50000;
      43928: inst = 32'h24612800;
      43929: inst = 32'h10a0ffff;
      43930: inst = 32'hca0ffe6;
      43931: inst = 32'h24822800;
      43932: inst = 32'h10a00000;
      43933: inst = 32'hca00004;
      43934: inst = 32'h38632800;
      43935: inst = 32'h38842800;
      43936: inst = 32'h10a00000;
      43937: inst = 32'hca0aba5;
      43938: inst = 32'h13e00001;
      43939: inst = 32'hfe0d96a;
      43940: inst = 32'h5be00000;
      43941: inst = 32'h8c50000;
      43942: inst = 32'h24612800;
      43943: inst = 32'h10a0ffff;
      43944: inst = 32'hca0ffe6;
      43945: inst = 32'h24822800;
      43946: inst = 32'h10a00000;
      43947: inst = 32'hca00004;
      43948: inst = 32'h38632800;
      43949: inst = 32'h38842800;
      43950: inst = 32'h10a00000;
      43951: inst = 32'hca0abb3;
      43952: inst = 32'h13e00001;
      43953: inst = 32'hfe0d96a;
      43954: inst = 32'h5be00000;
      43955: inst = 32'h8c50000;
      43956: inst = 32'h24612800;
      43957: inst = 32'h10a0ffff;
      43958: inst = 32'hca0ffe6;
      43959: inst = 32'h24822800;
      43960: inst = 32'h10a00000;
      43961: inst = 32'hca00004;
      43962: inst = 32'h38632800;
      43963: inst = 32'h38842800;
      43964: inst = 32'h10a00000;
      43965: inst = 32'hca0abc1;
      43966: inst = 32'h13e00001;
      43967: inst = 32'hfe0d96a;
      43968: inst = 32'h5be00000;
      43969: inst = 32'h8c50000;
      43970: inst = 32'h24612800;
      43971: inst = 32'h10a0ffff;
      43972: inst = 32'hca0ffe6;
      43973: inst = 32'h24822800;
      43974: inst = 32'h10a00000;
      43975: inst = 32'hca00004;
      43976: inst = 32'h38632800;
      43977: inst = 32'h38842800;
      43978: inst = 32'h10a00000;
      43979: inst = 32'hca0abcf;
      43980: inst = 32'h13e00001;
      43981: inst = 32'hfe0d96a;
      43982: inst = 32'h5be00000;
      43983: inst = 32'h8c50000;
      43984: inst = 32'h24612800;
      43985: inst = 32'h10a0ffff;
      43986: inst = 32'hca0ffe6;
      43987: inst = 32'h24822800;
      43988: inst = 32'h10a00000;
      43989: inst = 32'hca00004;
      43990: inst = 32'h38632800;
      43991: inst = 32'h38842800;
      43992: inst = 32'h10a00000;
      43993: inst = 32'hca0abdd;
      43994: inst = 32'h13e00001;
      43995: inst = 32'hfe0d96a;
      43996: inst = 32'h5be00000;
      43997: inst = 32'h8c50000;
      43998: inst = 32'h24612800;
      43999: inst = 32'h10a0ffff;
      44000: inst = 32'hca0ffe6;
      44001: inst = 32'h24822800;
      44002: inst = 32'h10a00000;
      44003: inst = 32'hca00004;
      44004: inst = 32'h38632800;
      44005: inst = 32'h38842800;
      44006: inst = 32'h10a00000;
      44007: inst = 32'hca0abeb;
      44008: inst = 32'h13e00001;
      44009: inst = 32'hfe0d96a;
      44010: inst = 32'h5be00000;
      44011: inst = 32'h8c50000;
      44012: inst = 32'h24612800;
      44013: inst = 32'h10a0ffff;
      44014: inst = 32'hca0ffe6;
      44015: inst = 32'h24822800;
      44016: inst = 32'h10a00000;
      44017: inst = 32'hca00004;
      44018: inst = 32'h38632800;
      44019: inst = 32'h38842800;
      44020: inst = 32'h10a00000;
      44021: inst = 32'hca0abf9;
      44022: inst = 32'h13e00001;
      44023: inst = 32'hfe0d96a;
      44024: inst = 32'h5be00000;
      44025: inst = 32'h8c50000;
      44026: inst = 32'h24612800;
      44027: inst = 32'h10a0ffff;
      44028: inst = 32'hca0ffe6;
      44029: inst = 32'h24822800;
      44030: inst = 32'h10a00000;
      44031: inst = 32'hca00004;
      44032: inst = 32'h38632800;
      44033: inst = 32'h38842800;
      44034: inst = 32'h10a00000;
      44035: inst = 32'hca0ac07;
      44036: inst = 32'h13e00001;
      44037: inst = 32'hfe0d96a;
      44038: inst = 32'h5be00000;
      44039: inst = 32'h8c50000;
      44040: inst = 32'h24612800;
      44041: inst = 32'h10a0ffff;
      44042: inst = 32'hca0ffe6;
      44043: inst = 32'h24822800;
      44044: inst = 32'h10a00000;
      44045: inst = 32'hca00004;
      44046: inst = 32'h38632800;
      44047: inst = 32'h38842800;
      44048: inst = 32'h10a00000;
      44049: inst = 32'hca0ac15;
      44050: inst = 32'h13e00001;
      44051: inst = 32'hfe0d96a;
      44052: inst = 32'h5be00000;
      44053: inst = 32'h8c50000;
      44054: inst = 32'h24612800;
      44055: inst = 32'h10a0ffff;
      44056: inst = 32'hca0ffe6;
      44057: inst = 32'h24822800;
      44058: inst = 32'h10a00000;
      44059: inst = 32'hca00004;
      44060: inst = 32'h38632800;
      44061: inst = 32'h38842800;
      44062: inst = 32'h10a00000;
      44063: inst = 32'hca0ac23;
      44064: inst = 32'h13e00001;
      44065: inst = 32'hfe0d96a;
      44066: inst = 32'h5be00000;
      44067: inst = 32'h8c50000;
      44068: inst = 32'h24612800;
      44069: inst = 32'h10a0ffff;
      44070: inst = 32'hca0ffe6;
      44071: inst = 32'h24822800;
      44072: inst = 32'h10a00000;
      44073: inst = 32'hca00004;
      44074: inst = 32'h38632800;
      44075: inst = 32'h38842800;
      44076: inst = 32'h10a00000;
      44077: inst = 32'hca0ac31;
      44078: inst = 32'h13e00001;
      44079: inst = 32'hfe0d96a;
      44080: inst = 32'h5be00000;
      44081: inst = 32'h8c50000;
      44082: inst = 32'h24612800;
      44083: inst = 32'h10a0ffff;
      44084: inst = 32'hca0ffe6;
      44085: inst = 32'h24822800;
      44086: inst = 32'h10a00000;
      44087: inst = 32'hca00004;
      44088: inst = 32'h38632800;
      44089: inst = 32'h38842800;
      44090: inst = 32'h10a00000;
      44091: inst = 32'hca0ac3f;
      44092: inst = 32'h13e00001;
      44093: inst = 32'hfe0d96a;
      44094: inst = 32'h5be00000;
      44095: inst = 32'h8c50000;
      44096: inst = 32'h24612800;
      44097: inst = 32'h10a0ffff;
      44098: inst = 32'hca0ffe6;
      44099: inst = 32'h24822800;
      44100: inst = 32'h10a00000;
      44101: inst = 32'hca00004;
      44102: inst = 32'h38632800;
      44103: inst = 32'h38842800;
      44104: inst = 32'h10a00000;
      44105: inst = 32'hca0ac4d;
      44106: inst = 32'h13e00001;
      44107: inst = 32'hfe0d96a;
      44108: inst = 32'h5be00000;
      44109: inst = 32'h8c50000;
      44110: inst = 32'h24612800;
      44111: inst = 32'h10a0ffff;
      44112: inst = 32'hca0ffe6;
      44113: inst = 32'h24822800;
      44114: inst = 32'h10a00000;
      44115: inst = 32'hca00004;
      44116: inst = 32'h38632800;
      44117: inst = 32'h38842800;
      44118: inst = 32'h10a00000;
      44119: inst = 32'hca0ac5b;
      44120: inst = 32'h13e00001;
      44121: inst = 32'hfe0d96a;
      44122: inst = 32'h5be00000;
      44123: inst = 32'h8c50000;
      44124: inst = 32'h24612800;
      44125: inst = 32'h10a0ffff;
      44126: inst = 32'hca0ffe6;
      44127: inst = 32'h24822800;
      44128: inst = 32'h10a00000;
      44129: inst = 32'hca00004;
      44130: inst = 32'h38632800;
      44131: inst = 32'h38842800;
      44132: inst = 32'h10a00000;
      44133: inst = 32'hca0ac69;
      44134: inst = 32'h13e00001;
      44135: inst = 32'hfe0d96a;
      44136: inst = 32'h5be00000;
      44137: inst = 32'h8c50000;
      44138: inst = 32'h24612800;
      44139: inst = 32'h10a0ffff;
      44140: inst = 32'hca0ffe6;
      44141: inst = 32'h24822800;
      44142: inst = 32'h10a00000;
      44143: inst = 32'hca00004;
      44144: inst = 32'h38632800;
      44145: inst = 32'h38842800;
      44146: inst = 32'h10a00000;
      44147: inst = 32'hca0ac77;
      44148: inst = 32'h13e00001;
      44149: inst = 32'hfe0d96a;
      44150: inst = 32'h5be00000;
      44151: inst = 32'h8c50000;
      44152: inst = 32'h24612800;
      44153: inst = 32'h10a0ffff;
      44154: inst = 32'hca0ffe6;
      44155: inst = 32'h24822800;
      44156: inst = 32'h10a00000;
      44157: inst = 32'hca00004;
      44158: inst = 32'h38632800;
      44159: inst = 32'h38842800;
      44160: inst = 32'h10a00000;
      44161: inst = 32'hca0ac85;
      44162: inst = 32'h13e00001;
      44163: inst = 32'hfe0d96a;
      44164: inst = 32'h5be00000;
      44165: inst = 32'h8c50000;
      44166: inst = 32'h24612800;
      44167: inst = 32'h10a0ffff;
      44168: inst = 32'hca0ffe6;
      44169: inst = 32'h24822800;
      44170: inst = 32'h10a00000;
      44171: inst = 32'hca00004;
      44172: inst = 32'h38632800;
      44173: inst = 32'h38842800;
      44174: inst = 32'h10a00000;
      44175: inst = 32'hca0ac93;
      44176: inst = 32'h13e00001;
      44177: inst = 32'hfe0d96a;
      44178: inst = 32'h5be00000;
      44179: inst = 32'h8c50000;
      44180: inst = 32'h24612800;
      44181: inst = 32'h10a0ffff;
      44182: inst = 32'hca0ffe6;
      44183: inst = 32'h24822800;
      44184: inst = 32'h10a00000;
      44185: inst = 32'hca00004;
      44186: inst = 32'h38632800;
      44187: inst = 32'h38842800;
      44188: inst = 32'h10a00000;
      44189: inst = 32'hca0aca1;
      44190: inst = 32'h13e00001;
      44191: inst = 32'hfe0d96a;
      44192: inst = 32'h5be00000;
      44193: inst = 32'h8c50000;
      44194: inst = 32'h24612800;
      44195: inst = 32'h10a0ffff;
      44196: inst = 32'hca0ffe6;
      44197: inst = 32'h24822800;
      44198: inst = 32'h10a00000;
      44199: inst = 32'hca00004;
      44200: inst = 32'h38632800;
      44201: inst = 32'h38842800;
      44202: inst = 32'h10a00000;
      44203: inst = 32'hca0acaf;
      44204: inst = 32'h13e00001;
      44205: inst = 32'hfe0d96a;
      44206: inst = 32'h5be00000;
      44207: inst = 32'h8c50000;
      44208: inst = 32'h24612800;
      44209: inst = 32'h10a0ffff;
      44210: inst = 32'hca0ffe6;
      44211: inst = 32'h24822800;
      44212: inst = 32'h10a00000;
      44213: inst = 32'hca00004;
      44214: inst = 32'h38632800;
      44215: inst = 32'h38842800;
      44216: inst = 32'h10a00000;
      44217: inst = 32'hca0acbd;
      44218: inst = 32'h13e00001;
      44219: inst = 32'hfe0d96a;
      44220: inst = 32'h5be00000;
      44221: inst = 32'h8c50000;
      44222: inst = 32'h24612800;
      44223: inst = 32'h10a0ffff;
      44224: inst = 32'hca0ffe6;
      44225: inst = 32'h24822800;
      44226: inst = 32'h10a00000;
      44227: inst = 32'hca00004;
      44228: inst = 32'h38632800;
      44229: inst = 32'h38842800;
      44230: inst = 32'h10a00000;
      44231: inst = 32'hca0accb;
      44232: inst = 32'h13e00001;
      44233: inst = 32'hfe0d96a;
      44234: inst = 32'h5be00000;
      44235: inst = 32'h8c50000;
      44236: inst = 32'h24612800;
      44237: inst = 32'h10a0ffff;
      44238: inst = 32'hca0ffe6;
      44239: inst = 32'h24822800;
      44240: inst = 32'h10a00000;
      44241: inst = 32'hca00004;
      44242: inst = 32'h38632800;
      44243: inst = 32'h38842800;
      44244: inst = 32'h10a00000;
      44245: inst = 32'hca0acd9;
      44246: inst = 32'h13e00001;
      44247: inst = 32'hfe0d96a;
      44248: inst = 32'h5be00000;
      44249: inst = 32'h8c50000;
      44250: inst = 32'h24612800;
      44251: inst = 32'h10a0ffff;
      44252: inst = 32'hca0ffe6;
      44253: inst = 32'h24822800;
      44254: inst = 32'h10a00000;
      44255: inst = 32'hca00004;
      44256: inst = 32'h38632800;
      44257: inst = 32'h38842800;
      44258: inst = 32'h10a00000;
      44259: inst = 32'hca0ace7;
      44260: inst = 32'h13e00001;
      44261: inst = 32'hfe0d96a;
      44262: inst = 32'h5be00000;
      44263: inst = 32'h8c50000;
      44264: inst = 32'h24612800;
      44265: inst = 32'h10a0ffff;
      44266: inst = 32'hca0ffe6;
      44267: inst = 32'h24822800;
      44268: inst = 32'h10a00000;
      44269: inst = 32'hca00004;
      44270: inst = 32'h38632800;
      44271: inst = 32'h38842800;
      44272: inst = 32'h10a00000;
      44273: inst = 32'hca0acf5;
      44274: inst = 32'h13e00001;
      44275: inst = 32'hfe0d96a;
      44276: inst = 32'h5be00000;
      44277: inst = 32'h8c50000;
      44278: inst = 32'h24612800;
      44279: inst = 32'h10a0ffff;
      44280: inst = 32'hca0ffe6;
      44281: inst = 32'h24822800;
      44282: inst = 32'h10a00000;
      44283: inst = 32'hca00004;
      44284: inst = 32'h38632800;
      44285: inst = 32'h38842800;
      44286: inst = 32'h10a00000;
      44287: inst = 32'hca0ad03;
      44288: inst = 32'h13e00001;
      44289: inst = 32'hfe0d96a;
      44290: inst = 32'h5be00000;
      44291: inst = 32'h8c50000;
      44292: inst = 32'h24612800;
      44293: inst = 32'h10a0ffff;
      44294: inst = 32'hca0ffe6;
      44295: inst = 32'h24822800;
      44296: inst = 32'h10a00000;
      44297: inst = 32'hca00004;
      44298: inst = 32'h38632800;
      44299: inst = 32'h38842800;
      44300: inst = 32'h10a00000;
      44301: inst = 32'hca0ad11;
      44302: inst = 32'h13e00001;
      44303: inst = 32'hfe0d96a;
      44304: inst = 32'h5be00000;
      44305: inst = 32'h8c50000;
      44306: inst = 32'h24612800;
      44307: inst = 32'h10a0ffff;
      44308: inst = 32'hca0ffe6;
      44309: inst = 32'h24822800;
      44310: inst = 32'h10a00000;
      44311: inst = 32'hca00004;
      44312: inst = 32'h38632800;
      44313: inst = 32'h38842800;
      44314: inst = 32'h10a00000;
      44315: inst = 32'hca0ad1f;
      44316: inst = 32'h13e00001;
      44317: inst = 32'hfe0d96a;
      44318: inst = 32'h5be00000;
      44319: inst = 32'h8c50000;
      44320: inst = 32'h24612800;
      44321: inst = 32'h10a0ffff;
      44322: inst = 32'hca0ffe6;
      44323: inst = 32'h24822800;
      44324: inst = 32'h10a00000;
      44325: inst = 32'hca00004;
      44326: inst = 32'h38632800;
      44327: inst = 32'h38842800;
      44328: inst = 32'h10a00000;
      44329: inst = 32'hca0ad2d;
      44330: inst = 32'h13e00001;
      44331: inst = 32'hfe0d96a;
      44332: inst = 32'h5be00000;
      44333: inst = 32'h8c50000;
      44334: inst = 32'h24612800;
      44335: inst = 32'h10a0ffff;
      44336: inst = 32'hca0ffe6;
      44337: inst = 32'h24822800;
      44338: inst = 32'h10a00000;
      44339: inst = 32'hca00004;
      44340: inst = 32'h38632800;
      44341: inst = 32'h38842800;
      44342: inst = 32'h10a00000;
      44343: inst = 32'hca0ad3b;
      44344: inst = 32'h13e00001;
      44345: inst = 32'hfe0d96a;
      44346: inst = 32'h5be00000;
      44347: inst = 32'h8c50000;
      44348: inst = 32'h24612800;
      44349: inst = 32'h10a0ffff;
      44350: inst = 32'hca0ffe6;
      44351: inst = 32'h24822800;
      44352: inst = 32'h10a00000;
      44353: inst = 32'hca00004;
      44354: inst = 32'h38632800;
      44355: inst = 32'h38842800;
      44356: inst = 32'h10a00000;
      44357: inst = 32'hca0ad49;
      44358: inst = 32'h13e00001;
      44359: inst = 32'hfe0d96a;
      44360: inst = 32'h5be00000;
      44361: inst = 32'h8c50000;
      44362: inst = 32'h24612800;
      44363: inst = 32'h10a0ffff;
      44364: inst = 32'hca0ffe6;
      44365: inst = 32'h24822800;
      44366: inst = 32'h10a00000;
      44367: inst = 32'hca00004;
      44368: inst = 32'h38632800;
      44369: inst = 32'h38842800;
      44370: inst = 32'h10a00000;
      44371: inst = 32'hca0ad57;
      44372: inst = 32'h13e00001;
      44373: inst = 32'hfe0d96a;
      44374: inst = 32'h5be00000;
      44375: inst = 32'h8c50000;
      44376: inst = 32'h24612800;
      44377: inst = 32'h10a0ffff;
      44378: inst = 32'hca0ffe6;
      44379: inst = 32'h24822800;
      44380: inst = 32'h10a00000;
      44381: inst = 32'hca00004;
      44382: inst = 32'h38632800;
      44383: inst = 32'h38842800;
      44384: inst = 32'h10a00000;
      44385: inst = 32'hca0ad65;
      44386: inst = 32'h13e00001;
      44387: inst = 32'hfe0d96a;
      44388: inst = 32'h5be00000;
      44389: inst = 32'h8c50000;
      44390: inst = 32'h24612800;
      44391: inst = 32'h10a0ffff;
      44392: inst = 32'hca0ffe6;
      44393: inst = 32'h24822800;
      44394: inst = 32'h10a00000;
      44395: inst = 32'hca00004;
      44396: inst = 32'h38632800;
      44397: inst = 32'h38842800;
      44398: inst = 32'h10a00000;
      44399: inst = 32'hca0ad73;
      44400: inst = 32'h13e00001;
      44401: inst = 32'hfe0d96a;
      44402: inst = 32'h5be00000;
      44403: inst = 32'h8c50000;
      44404: inst = 32'h24612800;
      44405: inst = 32'h10a0ffff;
      44406: inst = 32'hca0ffe6;
      44407: inst = 32'h24822800;
      44408: inst = 32'h10a00000;
      44409: inst = 32'hca00004;
      44410: inst = 32'h38632800;
      44411: inst = 32'h38842800;
      44412: inst = 32'h10a00000;
      44413: inst = 32'hca0ad81;
      44414: inst = 32'h13e00001;
      44415: inst = 32'hfe0d96a;
      44416: inst = 32'h5be00000;
      44417: inst = 32'h8c50000;
      44418: inst = 32'h24612800;
      44419: inst = 32'h10a0ffff;
      44420: inst = 32'hca0ffe6;
      44421: inst = 32'h24822800;
      44422: inst = 32'h10a00000;
      44423: inst = 32'hca00004;
      44424: inst = 32'h38632800;
      44425: inst = 32'h38842800;
      44426: inst = 32'h10a00000;
      44427: inst = 32'hca0ad8f;
      44428: inst = 32'h13e00001;
      44429: inst = 32'hfe0d96a;
      44430: inst = 32'h5be00000;
      44431: inst = 32'h8c50000;
      44432: inst = 32'h24612800;
      44433: inst = 32'h10a0ffff;
      44434: inst = 32'hca0ffe6;
      44435: inst = 32'h24822800;
      44436: inst = 32'h10a00000;
      44437: inst = 32'hca00004;
      44438: inst = 32'h38632800;
      44439: inst = 32'h38842800;
      44440: inst = 32'h10a00000;
      44441: inst = 32'hca0ad9d;
      44442: inst = 32'h13e00001;
      44443: inst = 32'hfe0d96a;
      44444: inst = 32'h5be00000;
      44445: inst = 32'h8c50000;
      44446: inst = 32'h24612800;
      44447: inst = 32'h10a0ffff;
      44448: inst = 32'hca0ffe6;
      44449: inst = 32'h24822800;
      44450: inst = 32'h10a00000;
      44451: inst = 32'hca00004;
      44452: inst = 32'h38632800;
      44453: inst = 32'h38842800;
      44454: inst = 32'h10a00000;
      44455: inst = 32'hca0adab;
      44456: inst = 32'h13e00001;
      44457: inst = 32'hfe0d96a;
      44458: inst = 32'h5be00000;
      44459: inst = 32'h8c50000;
      44460: inst = 32'h24612800;
      44461: inst = 32'h10a0ffff;
      44462: inst = 32'hca0ffe6;
      44463: inst = 32'h24822800;
      44464: inst = 32'h10a00000;
      44465: inst = 32'hca00004;
      44466: inst = 32'h38632800;
      44467: inst = 32'h38842800;
      44468: inst = 32'h10a00000;
      44469: inst = 32'hca0adb9;
      44470: inst = 32'h13e00001;
      44471: inst = 32'hfe0d96a;
      44472: inst = 32'h5be00000;
      44473: inst = 32'h8c50000;
      44474: inst = 32'h24612800;
      44475: inst = 32'h10a0ffff;
      44476: inst = 32'hca0ffe6;
      44477: inst = 32'h24822800;
      44478: inst = 32'h10a00000;
      44479: inst = 32'hca00004;
      44480: inst = 32'h38632800;
      44481: inst = 32'h38842800;
      44482: inst = 32'h10a00000;
      44483: inst = 32'hca0adc7;
      44484: inst = 32'h13e00001;
      44485: inst = 32'hfe0d96a;
      44486: inst = 32'h5be00000;
      44487: inst = 32'h8c50000;
      44488: inst = 32'h24612800;
      44489: inst = 32'h10a0ffff;
      44490: inst = 32'hca0ffe6;
      44491: inst = 32'h24822800;
      44492: inst = 32'h10a00000;
      44493: inst = 32'hca00004;
      44494: inst = 32'h38632800;
      44495: inst = 32'h38842800;
      44496: inst = 32'h10a00000;
      44497: inst = 32'hca0add5;
      44498: inst = 32'h13e00001;
      44499: inst = 32'hfe0d96a;
      44500: inst = 32'h5be00000;
      44501: inst = 32'h8c50000;
      44502: inst = 32'h24612800;
      44503: inst = 32'h10a0ffff;
      44504: inst = 32'hca0ffe6;
      44505: inst = 32'h24822800;
      44506: inst = 32'h10a00000;
      44507: inst = 32'hca00004;
      44508: inst = 32'h38632800;
      44509: inst = 32'h38842800;
      44510: inst = 32'h10a00000;
      44511: inst = 32'hca0ade3;
      44512: inst = 32'h13e00001;
      44513: inst = 32'hfe0d96a;
      44514: inst = 32'h5be00000;
      44515: inst = 32'h8c50000;
      44516: inst = 32'h24612800;
      44517: inst = 32'h10a0ffff;
      44518: inst = 32'hca0ffe6;
      44519: inst = 32'h24822800;
      44520: inst = 32'h10a00000;
      44521: inst = 32'hca00004;
      44522: inst = 32'h38632800;
      44523: inst = 32'h38842800;
      44524: inst = 32'h10a00000;
      44525: inst = 32'hca0adf1;
      44526: inst = 32'h13e00001;
      44527: inst = 32'hfe0d96a;
      44528: inst = 32'h5be00000;
      44529: inst = 32'h8c50000;
      44530: inst = 32'h24612800;
      44531: inst = 32'h10a0ffff;
      44532: inst = 32'hca0ffe6;
      44533: inst = 32'h24822800;
      44534: inst = 32'h10a00000;
      44535: inst = 32'hca00004;
      44536: inst = 32'h38632800;
      44537: inst = 32'h38842800;
      44538: inst = 32'h10a00000;
      44539: inst = 32'hca0adff;
      44540: inst = 32'h13e00001;
      44541: inst = 32'hfe0d96a;
      44542: inst = 32'h5be00000;
      44543: inst = 32'h8c50000;
      44544: inst = 32'h24612800;
      44545: inst = 32'h10a0ffff;
      44546: inst = 32'hca0ffe6;
      44547: inst = 32'h24822800;
      44548: inst = 32'h10a00000;
      44549: inst = 32'hca00004;
      44550: inst = 32'h38632800;
      44551: inst = 32'h38842800;
      44552: inst = 32'h10a00000;
      44553: inst = 32'hca0ae0d;
      44554: inst = 32'h13e00001;
      44555: inst = 32'hfe0d96a;
      44556: inst = 32'h5be00000;
      44557: inst = 32'h8c50000;
      44558: inst = 32'h24612800;
      44559: inst = 32'h10a0ffff;
      44560: inst = 32'hca0ffe6;
      44561: inst = 32'h24822800;
      44562: inst = 32'h10a00000;
      44563: inst = 32'hca00004;
      44564: inst = 32'h38632800;
      44565: inst = 32'h38842800;
      44566: inst = 32'h10a00000;
      44567: inst = 32'hca0ae1b;
      44568: inst = 32'h13e00001;
      44569: inst = 32'hfe0d96a;
      44570: inst = 32'h5be00000;
      44571: inst = 32'h8c50000;
      44572: inst = 32'h24612800;
      44573: inst = 32'h10a0ffff;
      44574: inst = 32'hca0ffe6;
      44575: inst = 32'h24822800;
      44576: inst = 32'h10a00000;
      44577: inst = 32'hca00004;
      44578: inst = 32'h38632800;
      44579: inst = 32'h38842800;
      44580: inst = 32'h10a00000;
      44581: inst = 32'hca0ae29;
      44582: inst = 32'h13e00001;
      44583: inst = 32'hfe0d96a;
      44584: inst = 32'h5be00000;
      44585: inst = 32'h8c50000;
      44586: inst = 32'h24612800;
      44587: inst = 32'h10a0ffff;
      44588: inst = 32'hca0ffe7;
      44589: inst = 32'h24822800;
      44590: inst = 32'h10a00000;
      44591: inst = 32'hca00004;
      44592: inst = 32'h38632800;
      44593: inst = 32'h38842800;
      44594: inst = 32'h10a00000;
      44595: inst = 32'hca0ae37;
      44596: inst = 32'h13e00001;
      44597: inst = 32'hfe0d96a;
      44598: inst = 32'h5be00000;
      44599: inst = 32'h8c50000;
      44600: inst = 32'h24612800;
      44601: inst = 32'h10a0ffff;
      44602: inst = 32'hca0ffe7;
      44603: inst = 32'h24822800;
      44604: inst = 32'h10a00000;
      44605: inst = 32'hca00004;
      44606: inst = 32'h38632800;
      44607: inst = 32'h38842800;
      44608: inst = 32'h10a00000;
      44609: inst = 32'hca0ae45;
      44610: inst = 32'h13e00001;
      44611: inst = 32'hfe0d96a;
      44612: inst = 32'h5be00000;
      44613: inst = 32'h8c50000;
      44614: inst = 32'h24612800;
      44615: inst = 32'h10a0ffff;
      44616: inst = 32'hca0ffe7;
      44617: inst = 32'h24822800;
      44618: inst = 32'h10a00000;
      44619: inst = 32'hca00004;
      44620: inst = 32'h38632800;
      44621: inst = 32'h38842800;
      44622: inst = 32'h10a00000;
      44623: inst = 32'hca0ae53;
      44624: inst = 32'h13e00001;
      44625: inst = 32'hfe0d96a;
      44626: inst = 32'h5be00000;
      44627: inst = 32'h8c50000;
      44628: inst = 32'h24612800;
      44629: inst = 32'h10a0ffff;
      44630: inst = 32'hca0ffe7;
      44631: inst = 32'h24822800;
      44632: inst = 32'h10a00000;
      44633: inst = 32'hca00004;
      44634: inst = 32'h38632800;
      44635: inst = 32'h38842800;
      44636: inst = 32'h10a00000;
      44637: inst = 32'hca0ae61;
      44638: inst = 32'h13e00001;
      44639: inst = 32'hfe0d96a;
      44640: inst = 32'h5be00000;
      44641: inst = 32'h8c50000;
      44642: inst = 32'h24612800;
      44643: inst = 32'h10a0ffff;
      44644: inst = 32'hca0ffe7;
      44645: inst = 32'h24822800;
      44646: inst = 32'h10a00000;
      44647: inst = 32'hca00004;
      44648: inst = 32'h38632800;
      44649: inst = 32'h38842800;
      44650: inst = 32'h10a00000;
      44651: inst = 32'hca0ae6f;
      44652: inst = 32'h13e00001;
      44653: inst = 32'hfe0d96a;
      44654: inst = 32'h5be00000;
      44655: inst = 32'h8c50000;
      44656: inst = 32'h24612800;
      44657: inst = 32'h10a0ffff;
      44658: inst = 32'hca0ffe7;
      44659: inst = 32'h24822800;
      44660: inst = 32'h10a00000;
      44661: inst = 32'hca00004;
      44662: inst = 32'h38632800;
      44663: inst = 32'h38842800;
      44664: inst = 32'h10a00000;
      44665: inst = 32'hca0ae7d;
      44666: inst = 32'h13e00001;
      44667: inst = 32'hfe0d96a;
      44668: inst = 32'h5be00000;
      44669: inst = 32'h8c50000;
      44670: inst = 32'h24612800;
      44671: inst = 32'h10a0ffff;
      44672: inst = 32'hca0ffe7;
      44673: inst = 32'h24822800;
      44674: inst = 32'h10a00000;
      44675: inst = 32'hca00004;
      44676: inst = 32'h38632800;
      44677: inst = 32'h38842800;
      44678: inst = 32'h10a00000;
      44679: inst = 32'hca0ae8b;
      44680: inst = 32'h13e00001;
      44681: inst = 32'hfe0d96a;
      44682: inst = 32'h5be00000;
      44683: inst = 32'h8c50000;
      44684: inst = 32'h24612800;
      44685: inst = 32'h10a0ffff;
      44686: inst = 32'hca0ffe7;
      44687: inst = 32'h24822800;
      44688: inst = 32'h10a00000;
      44689: inst = 32'hca00004;
      44690: inst = 32'h38632800;
      44691: inst = 32'h38842800;
      44692: inst = 32'h10a00000;
      44693: inst = 32'hca0ae99;
      44694: inst = 32'h13e00001;
      44695: inst = 32'hfe0d96a;
      44696: inst = 32'h5be00000;
      44697: inst = 32'h8c50000;
      44698: inst = 32'h24612800;
      44699: inst = 32'h10a0ffff;
      44700: inst = 32'hca0ffe7;
      44701: inst = 32'h24822800;
      44702: inst = 32'h10a00000;
      44703: inst = 32'hca00004;
      44704: inst = 32'h38632800;
      44705: inst = 32'h38842800;
      44706: inst = 32'h10a00000;
      44707: inst = 32'hca0aea7;
      44708: inst = 32'h13e00001;
      44709: inst = 32'hfe0d96a;
      44710: inst = 32'h5be00000;
      44711: inst = 32'h8c50000;
      44712: inst = 32'h24612800;
      44713: inst = 32'h10a0ffff;
      44714: inst = 32'hca0ffe7;
      44715: inst = 32'h24822800;
      44716: inst = 32'h10a00000;
      44717: inst = 32'hca00004;
      44718: inst = 32'h38632800;
      44719: inst = 32'h38842800;
      44720: inst = 32'h10a00000;
      44721: inst = 32'hca0aeb5;
      44722: inst = 32'h13e00001;
      44723: inst = 32'hfe0d96a;
      44724: inst = 32'h5be00000;
      44725: inst = 32'h8c50000;
      44726: inst = 32'h24612800;
      44727: inst = 32'h10a0ffff;
      44728: inst = 32'hca0ffe7;
      44729: inst = 32'h24822800;
      44730: inst = 32'h10a00000;
      44731: inst = 32'hca00004;
      44732: inst = 32'h38632800;
      44733: inst = 32'h38842800;
      44734: inst = 32'h10a00000;
      44735: inst = 32'hca0aec3;
      44736: inst = 32'h13e00001;
      44737: inst = 32'hfe0d96a;
      44738: inst = 32'h5be00000;
      44739: inst = 32'h8c50000;
      44740: inst = 32'h24612800;
      44741: inst = 32'h10a0ffff;
      44742: inst = 32'hca0ffe7;
      44743: inst = 32'h24822800;
      44744: inst = 32'h10a00000;
      44745: inst = 32'hca00004;
      44746: inst = 32'h38632800;
      44747: inst = 32'h38842800;
      44748: inst = 32'h10a00000;
      44749: inst = 32'hca0aed1;
      44750: inst = 32'h13e00001;
      44751: inst = 32'hfe0d96a;
      44752: inst = 32'h5be00000;
      44753: inst = 32'h8c50000;
      44754: inst = 32'h24612800;
      44755: inst = 32'h10a0ffff;
      44756: inst = 32'hca0ffe7;
      44757: inst = 32'h24822800;
      44758: inst = 32'h10a00000;
      44759: inst = 32'hca00004;
      44760: inst = 32'h38632800;
      44761: inst = 32'h38842800;
      44762: inst = 32'h10a00000;
      44763: inst = 32'hca0aedf;
      44764: inst = 32'h13e00001;
      44765: inst = 32'hfe0d96a;
      44766: inst = 32'h5be00000;
      44767: inst = 32'h8c50000;
      44768: inst = 32'h24612800;
      44769: inst = 32'h10a0ffff;
      44770: inst = 32'hca0ffe7;
      44771: inst = 32'h24822800;
      44772: inst = 32'h10a00000;
      44773: inst = 32'hca00004;
      44774: inst = 32'h38632800;
      44775: inst = 32'h38842800;
      44776: inst = 32'h10a00000;
      44777: inst = 32'hca0aeed;
      44778: inst = 32'h13e00001;
      44779: inst = 32'hfe0d96a;
      44780: inst = 32'h5be00000;
      44781: inst = 32'h8c50000;
      44782: inst = 32'h24612800;
      44783: inst = 32'h10a0ffff;
      44784: inst = 32'hca0ffe7;
      44785: inst = 32'h24822800;
      44786: inst = 32'h10a00000;
      44787: inst = 32'hca00004;
      44788: inst = 32'h38632800;
      44789: inst = 32'h38842800;
      44790: inst = 32'h10a00000;
      44791: inst = 32'hca0aefb;
      44792: inst = 32'h13e00001;
      44793: inst = 32'hfe0d96a;
      44794: inst = 32'h5be00000;
      44795: inst = 32'h8c50000;
      44796: inst = 32'h24612800;
      44797: inst = 32'h10a0ffff;
      44798: inst = 32'hca0ffe7;
      44799: inst = 32'h24822800;
      44800: inst = 32'h10a00000;
      44801: inst = 32'hca00004;
      44802: inst = 32'h38632800;
      44803: inst = 32'h38842800;
      44804: inst = 32'h10a00000;
      44805: inst = 32'hca0af09;
      44806: inst = 32'h13e00001;
      44807: inst = 32'hfe0d96a;
      44808: inst = 32'h5be00000;
      44809: inst = 32'h8c50000;
      44810: inst = 32'h24612800;
      44811: inst = 32'h10a0ffff;
      44812: inst = 32'hca0ffe7;
      44813: inst = 32'h24822800;
      44814: inst = 32'h10a00000;
      44815: inst = 32'hca00004;
      44816: inst = 32'h38632800;
      44817: inst = 32'h38842800;
      44818: inst = 32'h10a00000;
      44819: inst = 32'hca0af17;
      44820: inst = 32'h13e00001;
      44821: inst = 32'hfe0d96a;
      44822: inst = 32'h5be00000;
      44823: inst = 32'h8c50000;
      44824: inst = 32'h24612800;
      44825: inst = 32'h10a0ffff;
      44826: inst = 32'hca0ffe7;
      44827: inst = 32'h24822800;
      44828: inst = 32'h10a00000;
      44829: inst = 32'hca00004;
      44830: inst = 32'h38632800;
      44831: inst = 32'h38842800;
      44832: inst = 32'h10a00000;
      44833: inst = 32'hca0af25;
      44834: inst = 32'h13e00001;
      44835: inst = 32'hfe0d96a;
      44836: inst = 32'h5be00000;
      44837: inst = 32'h8c50000;
      44838: inst = 32'h24612800;
      44839: inst = 32'h10a0ffff;
      44840: inst = 32'hca0ffe7;
      44841: inst = 32'h24822800;
      44842: inst = 32'h10a00000;
      44843: inst = 32'hca00004;
      44844: inst = 32'h38632800;
      44845: inst = 32'h38842800;
      44846: inst = 32'h10a00000;
      44847: inst = 32'hca0af33;
      44848: inst = 32'h13e00001;
      44849: inst = 32'hfe0d96a;
      44850: inst = 32'h5be00000;
      44851: inst = 32'h8c50000;
      44852: inst = 32'h24612800;
      44853: inst = 32'h10a0ffff;
      44854: inst = 32'hca0ffe7;
      44855: inst = 32'h24822800;
      44856: inst = 32'h10a00000;
      44857: inst = 32'hca00004;
      44858: inst = 32'h38632800;
      44859: inst = 32'h38842800;
      44860: inst = 32'h10a00000;
      44861: inst = 32'hca0af41;
      44862: inst = 32'h13e00001;
      44863: inst = 32'hfe0d96a;
      44864: inst = 32'h5be00000;
      44865: inst = 32'h8c50000;
      44866: inst = 32'h24612800;
      44867: inst = 32'h10a0ffff;
      44868: inst = 32'hca0ffe7;
      44869: inst = 32'h24822800;
      44870: inst = 32'h10a00000;
      44871: inst = 32'hca00004;
      44872: inst = 32'h38632800;
      44873: inst = 32'h38842800;
      44874: inst = 32'h10a00000;
      44875: inst = 32'hca0af4f;
      44876: inst = 32'h13e00001;
      44877: inst = 32'hfe0d96a;
      44878: inst = 32'h5be00000;
      44879: inst = 32'h8c50000;
      44880: inst = 32'h24612800;
      44881: inst = 32'h10a0ffff;
      44882: inst = 32'hca0ffe7;
      44883: inst = 32'h24822800;
      44884: inst = 32'h10a00000;
      44885: inst = 32'hca00004;
      44886: inst = 32'h38632800;
      44887: inst = 32'h38842800;
      44888: inst = 32'h10a00000;
      44889: inst = 32'hca0af5d;
      44890: inst = 32'h13e00001;
      44891: inst = 32'hfe0d96a;
      44892: inst = 32'h5be00000;
      44893: inst = 32'h8c50000;
      44894: inst = 32'h24612800;
      44895: inst = 32'h10a0ffff;
      44896: inst = 32'hca0ffe7;
      44897: inst = 32'h24822800;
      44898: inst = 32'h10a00000;
      44899: inst = 32'hca00004;
      44900: inst = 32'h38632800;
      44901: inst = 32'h38842800;
      44902: inst = 32'h10a00000;
      44903: inst = 32'hca0af6b;
      44904: inst = 32'h13e00001;
      44905: inst = 32'hfe0d96a;
      44906: inst = 32'h5be00000;
      44907: inst = 32'h8c50000;
      44908: inst = 32'h24612800;
      44909: inst = 32'h10a0ffff;
      44910: inst = 32'hca0ffe7;
      44911: inst = 32'h24822800;
      44912: inst = 32'h10a00000;
      44913: inst = 32'hca00004;
      44914: inst = 32'h38632800;
      44915: inst = 32'h38842800;
      44916: inst = 32'h10a00000;
      44917: inst = 32'hca0af79;
      44918: inst = 32'h13e00001;
      44919: inst = 32'hfe0d96a;
      44920: inst = 32'h5be00000;
      44921: inst = 32'h8c50000;
      44922: inst = 32'h24612800;
      44923: inst = 32'h10a0ffff;
      44924: inst = 32'hca0ffe7;
      44925: inst = 32'h24822800;
      44926: inst = 32'h10a00000;
      44927: inst = 32'hca00004;
      44928: inst = 32'h38632800;
      44929: inst = 32'h38842800;
      44930: inst = 32'h10a00000;
      44931: inst = 32'hca0af87;
      44932: inst = 32'h13e00001;
      44933: inst = 32'hfe0d96a;
      44934: inst = 32'h5be00000;
      44935: inst = 32'h8c50000;
      44936: inst = 32'h24612800;
      44937: inst = 32'h10a0ffff;
      44938: inst = 32'hca0ffe7;
      44939: inst = 32'h24822800;
      44940: inst = 32'h10a00000;
      44941: inst = 32'hca00004;
      44942: inst = 32'h38632800;
      44943: inst = 32'h38842800;
      44944: inst = 32'h10a00000;
      44945: inst = 32'hca0af95;
      44946: inst = 32'h13e00001;
      44947: inst = 32'hfe0d96a;
      44948: inst = 32'h5be00000;
      44949: inst = 32'h8c50000;
      44950: inst = 32'h24612800;
      44951: inst = 32'h10a0ffff;
      44952: inst = 32'hca0ffe7;
      44953: inst = 32'h24822800;
      44954: inst = 32'h10a00000;
      44955: inst = 32'hca00004;
      44956: inst = 32'h38632800;
      44957: inst = 32'h38842800;
      44958: inst = 32'h10a00000;
      44959: inst = 32'hca0afa3;
      44960: inst = 32'h13e00001;
      44961: inst = 32'hfe0d96a;
      44962: inst = 32'h5be00000;
      44963: inst = 32'h8c50000;
      44964: inst = 32'h24612800;
      44965: inst = 32'h10a0ffff;
      44966: inst = 32'hca0ffe7;
      44967: inst = 32'h24822800;
      44968: inst = 32'h10a00000;
      44969: inst = 32'hca00004;
      44970: inst = 32'h38632800;
      44971: inst = 32'h38842800;
      44972: inst = 32'h10a00000;
      44973: inst = 32'hca0afb1;
      44974: inst = 32'h13e00001;
      44975: inst = 32'hfe0d96a;
      44976: inst = 32'h5be00000;
      44977: inst = 32'h8c50000;
      44978: inst = 32'h24612800;
      44979: inst = 32'h10a0ffff;
      44980: inst = 32'hca0ffe7;
      44981: inst = 32'h24822800;
      44982: inst = 32'h10a00000;
      44983: inst = 32'hca00004;
      44984: inst = 32'h38632800;
      44985: inst = 32'h38842800;
      44986: inst = 32'h10a00000;
      44987: inst = 32'hca0afbf;
      44988: inst = 32'h13e00001;
      44989: inst = 32'hfe0d96a;
      44990: inst = 32'h5be00000;
      44991: inst = 32'h8c50000;
      44992: inst = 32'h24612800;
      44993: inst = 32'h10a0ffff;
      44994: inst = 32'hca0ffe7;
      44995: inst = 32'h24822800;
      44996: inst = 32'h10a00000;
      44997: inst = 32'hca00004;
      44998: inst = 32'h38632800;
      44999: inst = 32'h38842800;
      45000: inst = 32'h10a00000;
      45001: inst = 32'hca0afcd;
      45002: inst = 32'h13e00001;
      45003: inst = 32'hfe0d96a;
      45004: inst = 32'h5be00000;
      45005: inst = 32'h8c50000;
      45006: inst = 32'h24612800;
      45007: inst = 32'h10a0ffff;
      45008: inst = 32'hca0ffe7;
      45009: inst = 32'h24822800;
      45010: inst = 32'h10a00000;
      45011: inst = 32'hca00004;
      45012: inst = 32'h38632800;
      45013: inst = 32'h38842800;
      45014: inst = 32'h10a00000;
      45015: inst = 32'hca0afdb;
      45016: inst = 32'h13e00001;
      45017: inst = 32'hfe0d96a;
      45018: inst = 32'h5be00000;
      45019: inst = 32'h8c50000;
      45020: inst = 32'h24612800;
      45021: inst = 32'h10a0ffff;
      45022: inst = 32'hca0ffe7;
      45023: inst = 32'h24822800;
      45024: inst = 32'h10a00000;
      45025: inst = 32'hca00004;
      45026: inst = 32'h38632800;
      45027: inst = 32'h38842800;
      45028: inst = 32'h10a00000;
      45029: inst = 32'hca0afe9;
      45030: inst = 32'h13e00001;
      45031: inst = 32'hfe0d96a;
      45032: inst = 32'h5be00000;
      45033: inst = 32'h8c50000;
      45034: inst = 32'h24612800;
      45035: inst = 32'h10a0ffff;
      45036: inst = 32'hca0ffe7;
      45037: inst = 32'h24822800;
      45038: inst = 32'h10a00000;
      45039: inst = 32'hca00004;
      45040: inst = 32'h38632800;
      45041: inst = 32'h38842800;
      45042: inst = 32'h10a00000;
      45043: inst = 32'hca0aff7;
      45044: inst = 32'h13e00001;
      45045: inst = 32'hfe0d96a;
      45046: inst = 32'h5be00000;
      45047: inst = 32'h8c50000;
      45048: inst = 32'h24612800;
      45049: inst = 32'h10a0ffff;
      45050: inst = 32'hca0ffe7;
      45051: inst = 32'h24822800;
      45052: inst = 32'h10a00000;
      45053: inst = 32'hca00004;
      45054: inst = 32'h38632800;
      45055: inst = 32'h38842800;
      45056: inst = 32'h10a00000;
      45057: inst = 32'hca0b005;
      45058: inst = 32'h13e00001;
      45059: inst = 32'hfe0d96a;
      45060: inst = 32'h5be00000;
      45061: inst = 32'h8c50000;
      45062: inst = 32'h24612800;
      45063: inst = 32'h10a0ffff;
      45064: inst = 32'hca0ffe7;
      45065: inst = 32'h24822800;
      45066: inst = 32'h10a00000;
      45067: inst = 32'hca00004;
      45068: inst = 32'h38632800;
      45069: inst = 32'h38842800;
      45070: inst = 32'h10a00000;
      45071: inst = 32'hca0b013;
      45072: inst = 32'h13e00001;
      45073: inst = 32'hfe0d96a;
      45074: inst = 32'h5be00000;
      45075: inst = 32'h8c50000;
      45076: inst = 32'h24612800;
      45077: inst = 32'h10a0ffff;
      45078: inst = 32'hca0ffe7;
      45079: inst = 32'h24822800;
      45080: inst = 32'h10a00000;
      45081: inst = 32'hca00004;
      45082: inst = 32'h38632800;
      45083: inst = 32'h38842800;
      45084: inst = 32'h10a00000;
      45085: inst = 32'hca0b021;
      45086: inst = 32'h13e00001;
      45087: inst = 32'hfe0d96a;
      45088: inst = 32'h5be00000;
      45089: inst = 32'h8c50000;
      45090: inst = 32'h24612800;
      45091: inst = 32'h10a0ffff;
      45092: inst = 32'hca0ffe7;
      45093: inst = 32'h24822800;
      45094: inst = 32'h10a00000;
      45095: inst = 32'hca00004;
      45096: inst = 32'h38632800;
      45097: inst = 32'h38842800;
      45098: inst = 32'h10a00000;
      45099: inst = 32'hca0b02f;
      45100: inst = 32'h13e00001;
      45101: inst = 32'hfe0d96a;
      45102: inst = 32'h5be00000;
      45103: inst = 32'h8c50000;
      45104: inst = 32'h24612800;
      45105: inst = 32'h10a0ffff;
      45106: inst = 32'hca0ffe7;
      45107: inst = 32'h24822800;
      45108: inst = 32'h10a00000;
      45109: inst = 32'hca00004;
      45110: inst = 32'h38632800;
      45111: inst = 32'h38842800;
      45112: inst = 32'h10a00000;
      45113: inst = 32'hca0b03d;
      45114: inst = 32'h13e00001;
      45115: inst = 32'hfe0d96a;
      45116: inst = 32'h5be00000;
      45117: inst = 32'h8c50000;
      45118: inst = 32'h24612800;
      45119: inst = 32'h10a0ffff;
      45120: inst = 32'hca0ffe7;
      45121: inst = 32'h24822800;
      45122: inst = 32'h10a00000;
      45123: inst = 32'hca00004;
      45124: inst = 32'h38632800;
      45125: inst = 32'h38842800;
      45126: inst = 32'h10a00000;
      45127: inst = 32'hca0b04b;
      45128: inst = 32'h13e00001;
      45129: inst = 32'hfe0d96a;
      45130: inst = 32'h5be00000;
      45131: inst = 32'h8c50000;
      45132: inst = 32'h24612800;
      45133: inst = 32'h10a0ffff;
      45134: inst = 32'hca0ffe7;
      45135: inst = 32'h24822800;
      45136: inst = 32'h10a00000;
      45137: inst = 32'hca00004;
      45138: inst = 32'h38632800;
      45139: inst = 32'h38842800;
      45140: inst = 32'h10a00000;
      45141: inst = 32'hca0b059;
      45142: inst = 32'h13e00001;
      45143: inst = 32'hfe0d96a;
      45144: inst = 32'h5be00000;
      45145: inst = 32'h8c50000;
      45146: inst = 32'h24612800;
      45147: inst = 32'h10a0ffff;
      45148: inst = 32'hca0ffe7;
      45149: inst = 32'h24822800;
      45150: inst = 32'h10a00000;
      45151: inst = 32'hca00004;
      45152: inst = 32'h38632800;
      45153: inst = 32'h38842800;
      45154: inst = 32'h10a00000;
      45155: inst = 32'hca0b067;
      45156: inst = 32'h13e00001;
      45157: inst = 32'hfe0d96a;
      45158: inst = 32'h5be00000;
      45159: inst = 32'h8c50000;
      45160: inst = 32'h24612800;
      45161: inst = 32'h10a0ffff;
      45162: inst = 32'hca0ffe7;
      45163: inst = 32'h24822800;
      45164: inst = 32'h10a00000;
      45165: inst = 32'hca00004;
      45166: inst = 32'h38632800;
      45167: inst = 32'h38842800;
      45168: inst = 32'h10a00000;
      45169: inst = 32'hca0b075;
      45170: inst = 32'h13e00001;
      45171: inst = 32'hfe0d96a;
      45172: inst = 32'h5be00000;
      45173: inst = 32'h8c50000;
      45174: inst = 32'h24612800;
      45175: inst = 32'h10a0ffff;
      45176: inst = 32'hca0ffe7;
      45177: inst = 32'h24822800;
      45178: inst = 32'h10a00000;
      45179: inst = 32'hca00004;
      45180: inst = 32'h38632800;
      45181: inst = 32'h38842800;
      45182: inst = 32'h10a00000;
      45183: inst = 32'hca0b083;
      45184: inst = 32'h13e00001;
      45185: inst = 32'hfe0d96a;
      45186: inst = 32'h5be00000;
      45187: inst = 32'h8c50000;
      45188: inst = 32'h24612800;
      45189: inst = 32'h10a0ffff;
      45190: inst = 32'hca0ffe7;
      45191: inst = 32'h24822800;
      45192: inst = 32'h10a00000;
      45193: inst = 32'hca00004;
      45194: inst = 32'h38632800;
      45195: inst = 32'h38842800;
      45196: inst = 32'h10a00000;
      45197: inst = 32'hca0b091;
      45198: inst = 32'h13e00001;
      45199: inst = 32'hfe0d96a;
      45200: inst = 32'h5be00000;
      45201: inst = 32'h8c50000;
      45202: inst = 32'h24612800;
      45203: inst = 32'h10a0ffff;
      45204: inst = 32'hca0ffe7;
      45205: inst = 32'h24822800;
      45206: inst = 32'h10a00000;
      45207: inst = 32'hca00004;
      45208: inst = 32'h38632800;
      45209: inst = 32'h38842800;
      45210: inst = 32'h10a00000;
      45211: inst = 32'hca0b09f;
      45212: inst = 32'h13e00001;
      45213: inst = 32'hfe0d96a;
      45214: inst = 32'h5be00000;
      45215: inst = 32'h8c50000;
      45216: inst = 32'h24612800;
      45217: inst = 32'h10a0ffff;
      45218: inst = 32'hca0ffe7;
      45219: inst = 32'h24822800;
      45220: inst = 32'h10a00000;
      45221: inst = 32'hca00004;
      45222: inst = 32'h38632800;
      45223: inst = 32'h38842800;
      45224: inst = 32'h10a00000;
      45225: inst = 32'hca0b0ad;
      45226: inst = 32'h13e00001;
      45227: inst = 32'hfe0d96a;
      45228: inst = 32'h5be00000;
      45229: inst = 32'h8c50000;
      45230: inst = 32'h24612800;
      45231: inst = 32'h10a0ffff;
      45232: inst = 32'hca0ffe7;
      45233: inst = 32'h24822800;
      45234: inst = 32'h10a00000;
      45235: inst = 32'hca00004;
      45236: inst = 32'h38632800;
      45237: inst = 32'h38842800;
      45238: inst = 32'h10a00000;
      45239: inst = 32'hca0b0bb;
      45240: inst = 32'h13e00001;
      45241: inst = 32'hfe0d96a;
      45242: inst = 32'h5be00000;
      45243: inst = 32'h8c50000;
      45244: inst = 32'h24612800;
      45245: inst = 32'h10a0ffff;
      45246: inst = 32'hca0ffe7;
      45247: inst = 32'h24822800;
      45248: inst = 32'h10a00000;
      45249: inst = 32'hca00004;
      45250: inst = 32'h38632800;
      45251: inst = 32'h38842800;
      45252: inst = 32'h10a00000;
      45253: inst = 32'hca0b0c9;
      45254: inst = 32'h13e00001;
      45255: inst = 32'hfe0d96a;
      45256: inst = 32'h5be00000;
      45257: inst = 32'h8c50000;
      45258: inst = 32'h24612800;
      45259: inst = 32'h10a0ffff;
      45260: inst = 32'hca0ffe7;
      45261: inst = 32'h24822800;
      45262: inst = 32'h10a00000;
      45263: inst = 32'hca00004;
      45264: inst = 32'h38632800;
      45265: inst = 32'h38842800;
      45266: inst = 32'h10a00000;
      45267: inst = 32'hca0b0d7;
      45268: inst = 32'h13e00001;
      45269: inst = 32'hfe0d96a;
      45270: inst = 32'h5be00000;
      45271: inst = 32'h8c50000;
      45272: inst = 32'h24612800;
      45273: inst = 32'h10a0ffff;
      45274: inst = 32'hca0ffe7;
      45275: inst = 32'h24822800;
      45276: inst = 32'h10a00000;
      45277: inst = 32'hca00004;
      45278: inst = 32'h38632800;
      45279: inst = 32'h38842800;
      45280: inst = 32'h10a00000;
      45281: inst = 32'hca0b0e5;
      45282: inst = 32'h13e00001;
      45283: inst = 32'hfe0d96a;
      45284: inst = 32'h5be00000;
      45285: inst = 32'h8c50000;
      45286: inst = 32'h24612800;
      45287: inst = 32'h10a0ffff;
      45288: inst = 32'hca0ffe7;
      45289: inst = 32'h24822800;
      45290: inst = 32'h10a00000;
      45291: inst = 32'hca00004;
      45292: inst = 32'h38632800;
      45293: inst = 32'h38842800;
      45294: inst = 32'h10a00000;
      45295: inst = 32'hca0b0f3;
      45296: inst = 32'h13e00001;
      45297: inst = 32'hfe0d96a;
      45298: inst = 32'h5be00000;
      45299: inst = 32'h8c50000;
      45300: inst = 32'h24612800;
      45301: inst = 32'h10a0ffff;
      45302: inst = 32'hca0ffe7;
      45303: inst = 32'h24822800;
      45304: inst = 32'h10a00000;
      45305: inst = 32'hca00004;
      45306: inst = 32'h38632800;
      45307: inst = 32'h38842800;
      45308: inst = 32'h10a00000;
      45309: inst = 32'hca0b101;
      45310: inst = 32'h13e00001;
      45311: inst = 32'hfe0d96a;
      45312: inst = 32'h5be00000;
      45313: inst = 32'h8c50000;
      45314: inst = 32'h24612800;
      45315: inst = 32'h10a0ffff;
      45316: inst = 32'hca0ffe7;
      45317: inst = 32'h24822800;
      45318: inst = 32'h10a00000;
      45319: inst = 32'hca00004;
      45320: inst = 32'h38632800;
      45321: inst = 32'h38842800;
      45322: inst = 32'h10a00000;
      45323: inst = 32'hca0b10f;
      45324: inst = 32'h13e00001;
      45325: inst = 32'hfe0d96a;
      45326: inst = 32'h5be00000;
      45327: inst = 32'h8c50000;
      45328: inst = 32'h24612800;
      45329: inst = 32'h10a0ffff;
      45330: inst = 32'hca0ffe7;
      45331: inst = 32'h24822800;
      45332: inst = 32'h10a00000;
      45333: inst = 32'hca00004;
      45334: inst = 32'h38632800;
      45335: inst = 32'h38842800;
      45336: inst = 32'h10a00000;
      45337: inst = 32'hca0b11d;
      45338: inst = 32'h13e00001;
      45339: inst = 32'hfe0d96a;
      45340: inst = 32'h5be00000;
      45341: inst = 32'h8c50000;
      45342: inst = 32'h24612800;
      45343: inst = 32'h10a0ffff;
      45344: inst = 32'hca0ffe7;
      45345: inst = 32'h24822800;
      45346: inst = 32'h10a00000;
      45347: inst = 32'hca00004;
      45348: inst = 32'h38632800;
      45349: inst = 32'h38842800;
      45350: inst = 32'h10a00000;
      45351: inst = 32'hca0b12b;
      45352: inst = 32'h13e00001;
      45353: inst = 32'hfe0d96a;
      45354: inst = 32'h5be00000;
      45355: inst = 32'h8c50000;
      45356: inst = 32'h24612800;
      45357: inst = 32'h10a0ffff;
      45358: inst = 32'hca0ffe7;
      45359: inst = 32'h24822800;
      45360: inst = 32'h10a00000;
      45361: inst = 32'hca00004;
      45362: inst = 32'h38632800;
      45363: inst = 32'h38842800;
      45364: inst = 32'h10a00000;
      45365: inst = 32'hca0b139;
      45366: inst = 32'h13e00001;
      45367: inst = 32'hfe0d96a;
      45368: inst = 32'h5be00000;
      45369: inst = 32'h8c50000;
      45370: inst = 32'h24612800;
      45371: inst = 32'h10a0ffff;
      45372: inst = 32'hca0ffe7;
      45373: inst = 32'h24822800;
      45374: inst = 32'h10a00000;
      45375: inst = 32'hca00004;
      45376: inst = 32'h38632800;
      45377: inst = 32'h38842800;
      45378: inst = 32'h10a00000;
      45379: inst = 32'hca0b147;
      45380: inst = 32'h13e00001;
      45381: inst = 32'hfe0d96a;
      45382: inst = 32'h5be00000;
      45383: inst = 32'h8c50000;
      45384: inst = 32'h24612800;
      45385: inst = 32'h10a0ffff;
      45386: inst = 32'hca0ffe7;
      45387: inst = 32'h24822800;
      45388: inst = 32'h10a00000;
      45389: inst = 32'hca00004;
      45390: inst = 32'h38632800;
      45391: inst = 32'h38842800;
      45392: inst = 32'h10a00000;
      45393: inst = 32'hca0b155;
      45394: inst = 32'h13e00001;
      45395: inst = 32'hfe0d96a;
      45396: inst = 32'h5be00000;
      45397: inst = 32'h8c50000;
      45398: inst = 32'h24612800;
      45399: inst = 32'h10a0ffff;
      45400: inst = 32'hca0ffe7;
      45401: inst = 32'h24822800;
      45402: inst = 32'h10a00000;
      45403: inst = 32'hca00004;
      45404: inst = 32'h38632800;
      45405: inst = 32'h38842800;
      45406: inst = 32'h10a00000;
      45407: inst = 32'hca0b163;
      45408: inst = 32'h13e00001;
      45409: inst = 32'hfe0d96a;
      45410: inst = 32'h5be00000;
      45411: inst = 32'h8c50000;
      45412: inst = 32'h24612800;
      45413: inst = 32'h10a0ffff;
      45414: inst = 32'hca0ffe7;
      45415: inst = 32'h24822800;
      45416: inst = 32'h10a00000;
      45417: inst = 32'hca00004;
      45418: inst = 32'h38632800;
      45419: inst = 32'h38842800;
      45420: inst = 32'h10a00000;
      45421: inst = 32'hca0b171;
      45422: inst = 32'h13e00001;
      45423: inst = 32'hfe0d96a;
      45424: inst = 32'h5be00000;
      45425: inst = 32'h8c50000;
      45426: inst = 32'h24612800;
      45427: inst = 32'h10a0ffff;
      45428: inst = 32'hca0ffe7;
      45429: inst = 32'h24822800;
      45430: inst = 32'h10a00000;
      45431: inst = 32'hca00004;
      45432: inst = 32'h38632800;
      45433: inst = 32'h38842800;
      45434: inst = 32'h10a00000;
      45435: inst = 32'hca0b17f;
      45436: inst = 32'h13e00001;
      45437: inst = 32'hfe0d96a;
      45438: inst = 32'h5be00000;
      45439: inst = 32'h8c50000;
      45440: inst = 32'h24612800;
      45441: inst = 32'h10a0ffff;
      45442: inst = 32'hca0ffe7;
      45443: inst = 32'h24822800;
      45444: inst = 32'h10a00000;
      45445: inst = 32'hca00004;
      45446: inst = 32'h38632800;
      45447: inst = 32'h38842800;
      45448: inst = 32'h10a00000;
      45449: inst = 32'hca0b18d;
      45450: inst = 32'h13e00001;
      45451: inst = 32'hfe0d96a;
      45452: inst = 32'h5be00000;
      45453: inst = 32'h8c50000;
      45454: inst = 32'h24612800;
      45455: inst = 32'h10a0ffff;
      45456: inst = 32'hca0ffe7;
      45457: inst = 32'h24822800;
      45458: inst = 32'h10a00000;
      45459: inst = 32'hca00004;
      45460: inst = 32'h38632800;
      45461: inst = 32'h38842800;
      45462: inst = 32'h10a00000;
      45463: inst = 32'hca0b19b;
      45464: inst = 32'h13e00001;
      45465: inst = 32'hfe0d96a;
      45466: inst = 32'h5be00000;
      45467: inst = 32'h8c50000;
      45468: inst = 32'h24612800;
      45469: inst = 32'h10a0ffff;
      45470: inst = 32'hca0ffe7;
      45471: inst = 32'h24822800;
      45472: inst = 32'h10a00000;
      45473: inst = 32'hca00004;
      45474: inst = 32'h38632800;
      45475: inst = 32'h38842800;
      45476: inst = 32'h10a00000;
      45477: inst = 32'hca0b1a9;
      45478: inst = 32'h13e00001;
      45479: inst = 32'hfe0d96a;
      45480: inst = 32'h5be00000;
      45481: inst = 32'h8c50000;
      45482: inst = 32'h24612800;
      45483: inst = 32'h10a0ffff;
      45484: inst = 32'hca0ffe7;
      45485: inst = 32'h24822800;
      45486: inst = 32'h10a00000;
      45487: inst = 32'hca00004;
      45488: inst = 32'h38632800;
      45489: inst = 32'h38842800;
      45490: inst = 32'h10a00000;
      45491: inst = 32'hca0b1b7;
      45492: inst = 32'h13e00001;
      45493: inst = 32'hfe0d96a;
      45494: inst = 32'h5be00000;
      45495: inst = 32'h8c50000;
      45496: inst = 32'h24612800;
      45497: inst = 32'h10a0ffff;
      45498: inst = 32'hca0ffe7;
      45499: inst = 32'h24822800;
      45500: inst = 32'h10a00000;
      45501: inst = 32'hca00004;
      45502: inst = 32'h38632800;
      45503: inst = 32'h38842800;
      45504: inst = 32'h10a00000;
      45505: inst = 32'hca0b1c5;
      45506: inst = 32'h13e00001;
      45507: inst = 32'hfe0d96a;
      45508: inst = 32'h5be00000;
      45509: inst = 32'h8c50000;
      45510: inst = 32'h24612800;
      45511: inst = 32'h10a0ffff;
      45512: inst = 32'hca0ffe7;
      45513: inst = 32'h24822800;
      45514: inst = 32'h10a00000;
      45515: inst = 32'hca00004;
      45516: inst = 32'h38632800;
      45517: inst = 32'h38842800;
      45518: inst = 32'h10a00000;
      45519: inst = 32'hca0b1d3;
      45520: inst = 32'h13e00001;
      45521: inst = 32'hfe0d96a;
      45522: inst = 32'h5be00000;
      45523: inst = 32'h8c50000;
      45524: inst = 32'h24612800;
      45525: inst = 32'h10a0ffff;
      45526: inst = 32'hca0ffe7;
      45527: inst = 32'h24822800;
      45528: inst = 32'h10a00000;
      45529: inst = 32'hca00004;
      45530: inst = 32'h38632800;
      45531: inst = 32'h38842800;
      45532: inst = 32'h10a00000;
      45533: inst = 32'hca0b1e1;
      45534: inst = 32'h13e00001;
      45535: inst = 32'hfe0d96a;
      45536: inst = 32'h5be00000;
      45537: inst = 32'h8c50000;
      45538: inst = 32'h24612800;
      45539: inst = 32'h10a0ffff;
      45540: inst = 32'hca0ffe7;
      45541: inst = 32'h24822800;
      45542: inst = 32'h10a00000;
      45543: inst = 32'hca00004;
      45544: inst = 32'h38632800;
      45545: inst = 32'h38842800;
      45546: inst = 32'h10a00000;
      45547: inst = 32'hca0b1ef;
      45548: inst = 32'h13e00001;
      45549: inst = 32'hfe0d96a;
      45550: inst = 32'h5be00000;
      45551: inst = 32'h8c50000;
      45552: inst = 32'h24612800;
      45553: inst = 32'h10a0ffff;
      45554: inst = 32'hca0ffe7;
      45555: inst = 32'h24822800;
      45556: inst = 32'h10a00000;
      45557: inst = 32'hca00004;
      45558: inst = 32'h38632800;
      45559: inst = 32'h38842800;
      45560: inst = 32'h10a00000;
      45561: inst = 32'hca0b1fd;
      45562: inst = 32'h13e00001;
      45563: inst = 32'hfe0d96a;
      45564: inst = 32'h5be00000;
      45565: inst = 32'h8c50000;
      45566: inst = 32'h24612800;
      45567: inst = 32'h10a0ffff;
      45568: inst = 32'hca0ffe7;
      45569: inst = 32'h24822800;
      45570: inst = 32'h10a00000;
      45571: inst = 32'hca00004;
      45572: inst = 32'h38632800;
      45573: inst = 32'h38842800;
      45574: inst = 32'h10a00000;
      45575: inst = 32'hca0b20b;
      45576: inst = 32'h13e00001;
      45577: inst = 32'hfe0d96a;
      45578: inst = 32'h5be00000;
      45579: inst = 32'h8c50000;
      45580: inst = 32'h24612800;
      45581: inst = 32'h10a0ffff;
      45582: inst = 32'hca0ffe7;
      45583: inst = 32'h24822800;
      45584: inst = 32'h10a00000;
      45585: inst = 32'hca00004;
      45586: inst = 32'h38632800;
      45587: inst = 32'h38842800;
      45588: inst = 32'h10a00000;
      45589: inst = 32'hca0b219;
      45590: inst = 32'h13e00001;
      45591: inst = 32'hfe0d96a;
      45592: inst = 32'h5be00000;
      45593: inst = 32'h8c50000;
      45594: inst = 32'h24612800;
      45595: inst = 32'h10a0ffff;
      45596: inst = 32'hca0ffe7;
      45597: inst = 32'h24822800;
      45598: inst = 32'h10a00000;
      45599: inst = 32'hca00004;
      45600: inst = 32'h38632800;
      45601: inst = 32'h38842800;
      45602: inst = 32'h10a00000;
      45603: inst = 32'hca0b227;
      45604: inst = 32'h13e00001;
      45605: inst = 32'hfe0d96a;
      45606: inst = 32'h5be00000;
      45607: inst = 32'h8c50000;
      45608: inst = 32'h24612800;
      45609: inst = 32'h10a0ffff;
      45610: inst = 32'hca0ffe7;
      45611: inst = 32'h24822800;
      45612: inst = 32'h10a00000;
      45613: inst = 32'hca00004;
      45614: inst = 32'h38632800;
      45615: inst = 32'h38842800;
      45616: inst = 32'h10a00000;
      45617: inst = 32'hca0b235;
      45618: inst = 32'h13e00001;
      45619: inst = 32'hfe0d96a;
      45620: inst = 32'h5be00000;
      45621: inst = 32'h8c50000;
      45622: inst = 32'h24612800;
      45623: inst = 32'h10a0ffff;
      45624: inst = 32'hca0ffe7;
      45625: inst = 32'h24822800;
      45626: inst = 32'h10a00000;
      45627: inst = 32'hca00004;
      45628: inst = 32'h38632800;
      45629: inst = 32'h38842800;
      45630: inst = 32'h10a00000;
      45631: inst = 32'hca0b243;
      45632: inst = 32'h13e00001;
      45633: inst = 32'hfe0d96a;
      45634: inst = 32'h5be00000;
      45635: inst = 32'h8c50000;
      45636: inst = 32'h24612800;
      45637: inst = 32'h10a0ffff;
      45638: inst = 32'hca0ffe7;
      45639: inst = 32'h24822800;
      45640: inst = 32'h10a00000;
      45641: inst = 32'hca00004;
      45642: inst = 32'h38632800;
      45643: inst = 32'h38842800;
      45644: inst = 32'h10a00000;
      45645: inst = 32'hca0b251;
      45646: inst = 32'h13e00001;
      45647: inst = 32'hfe0d96a;
      45648: inst = 32'h5be00000;
      45649: inst = 32'h8c50000;
      45650: inst = 32'h24612800;
      45651: inst = 32'h10a0ffff;
      45652: inst = 32'hca0ffe7;
      45653: inst = 32'h24822800;
      45654: inst = 32'h10a00000;
      45655: inst = 32'hca00004;
      45656: inst = 32'h38632800;
      45657: inst = 32'h38842800;
      45658: inst = 32'h10a00000;
      45659: inst = 32'hca0b25f;
      45660: inst = 32'h13e00001;
      45661: inst = 32'hfe0d96a;
      45662: inst = 32'h5be00000;
      45663: inst = 32'h8c50000;
      45664: inst = 32'h24612800;
      45665: inst = 32'h10a0ffff;
      45666: inst = 32'hca0ffe7;
      45667: inst = 32'h24822800;
      45668: inst = 32'h10a00000;
      45669: inst = 32'hca00004;
      45670: inst = 32'h38632800;
      45671: inst = 32'h38842800;
      45672: inst = 32'h10a00000;
      45673: inst = 32'hca0b26d;
      45674: inst = 32'h13e00001;
      45675: inst = 32'hfe0d96a;
      45676: inst = 32'h5be00000;
      45677: inst = 32'h8c50000;
      45678: inst = 32'h24612800;
      45679: inst = 32'h10a0ffff;
      45680: inst = 32'hca0ffe7;
      45681: inst = 32'h24822800;
      45682: inst = 32'h10a00000;
      45683: inst = 32'hca00004;
      45684: inst = 32'h38632800;
      45685: inst = 32'h38842800;
      45686: inst = 32'h10a00000;
      45687: inst = 32'hca0b27b;
      45688: inst = 32'h13e00001;
      45689: inst = 32'hfe0d96a;
      45690: inst = 32'h5be00000;
      45691: inst = 32'h8c50000;
      45692: inst = 32'h24612800;
      45693: inst = 32'h10a0ffff;
      45694: inst = 32'hca0ffe7;
      45695: inst = 32'h24822800;
      45696: inst = 32'h10a00000;
      45697: inst = 32'hca00004;
      45698: inst = 32'h38632800;
      45699: inst = 32'h38842800;
      45700: inst = 32'h10a00000;
      45701: inst = 32'hca0b289;
      45702: inst = 32'h13e00001;
      45703: inst = 32'hfe0d96a;
      45704: inst = 32'h5be00000;
      45705: inst = 32'h8c50000;
      45706: inst = 32'h24612800;
      45707: inst = 32'h10a0ffff;
      45708: inst = 32'hca0ffe7;
      45709: inst = 32'h24822800;
      45710: inst = 32'h10a00000;
      45711: inst = 32'hca00004;
      45712: inst = 32'h38632800;
      45713: inst = 32'h38842800;
      45714: inst = 32'h10a00000;
      45715: inst = 32'hca0b297;
      45716: inst = 32'h13e00001;
      45717: inst = 32'hfe0d96a;
      45718: inst = 32'h5be00000;
      45719: inst = 32'h8c50000;
      45720: inst = 32'h24612800;
      45721: inst = 32'h10a0ffff;
      45722: inst = 32'hca0ffe7;
      45723: inst = 32'h24822800;
      45724: inst = 32'h10a00000;
      45725: inst = 32'hca00004;
      45726: inst = 32'h38632800;
      45727: inst = 32'h38842800;
      45728: inst = 32'h10a00000;
      45729: inst = 32'hca0b2a5;
      45730: inst = 32'h13e00001;
      45731: inst = 32'hfe0d96a;
      45732: inst = 32'h5be00000;
      45733: inst = 32'h8c50000;
      45734: inst = 32'h24612800;
      45735: inst = 32'h10a0ffff;
      45736: inst = 32'hca0ffe7;
      45737: inst = 32'h24822800;
      45738: inst = 32'h10a00000;
      45739: inst = 32'hca00004;
      45740: inst = 32'h38632800;
      45741: inst = 32'h38842800;
      45742: inst = 32'h10a00000;
      45743: inst = 32'hca0b2b3;
      45744: inst = 32'h13e00001;
      45745: inst = 32'hfe0d96a;
      45746: inst = 32'h5be00000;
      45747: inst = 32'h8c50000;
      45748: inst = 32'h24612800;
      45749: inst = 32'h10a0ffff;
      45750: inst = 32'hca0ffe7;
      45751: inst = 32'h24822800;
      45752: inst = 32'h10a00000;
      45753: inst = 32'hca00004;
      45754: inst = 32'h38632800;
      45755: inst = 32'h38842800;
      45756: inst = 32'h10a00000;
      45757: inst = 32'hca0b2c1;
      45758: inst = 32'h13e00001;
      45759: inst = 32'hfe0d96a;
      45760: inst = 32'h5be00000;
      45761: inst = 32'h8c50000;
      45762: inst = 32'h24612800;
      45763: inst = 32'h10a0ffff;
      45764: inst = 32'hca0ffe7;
      45765: inst = 32'h24822800;
      45766: inst = 32'h10a00000;
      45767: inst = 32'hca00004;
      45768: inst = 32'h38632800;
      45769: inst = 32'h38842800;
      45770: inst = 32'h10a00000;
      45771: inst = 32'hca0b2cf;
      45772: inst = 32'h13e00001;
      45773: inst = 32'hfe0d96a;
      45774: inst = 32'h5be00000;
      45775: inst = 32'h8c50000;
      45776: inst = 32'h24612800;
      45777: inst = 32'h10a0ffff;
      45778: inst = 32'hca0ffe7;
      45779: inst = 32'h24822800;
      45780: inst = 32'h10a00000;
      45781: inst = 32'hca00004;
      45782: inst = 32'h38632800;
      45783: inst = 32'h38842800;
      45784: inst = 32'h10a00000;
      45785: inst = 32'hca0b2dd;
      45786: inst = 32'h13e00001;
      45787: inst = 32'hfe0d96a;
      45788: inst = 32'h5be00000;
      45789: inst = 32'h8c50000;
      45790: inst = 32'h24612800;
      45791: inst = 32'h10a0ffff;
      45792: inst = 32'hca0ffe7;
      45793: inst = 32'h24822800;
      45794: inst = 32'h10a00000;
      45795: inst = 32'hca00004;
      45796: inst = 32'h38632800;
      45797: inst = 32'h38842800;
      45798: inst = 32'h10a00000;
      45799: inst = 32'hca0b2eb;
      45800: inst = 32'h13e00001;
      45801: inst = 32'hfe0d96a;
      45802: inst = 32'h5be00000;
      45803: inst = 32'h8c50000;
      45804: inst = 32'h24612800;
      45805: inst = 32'h10a0ffff;
      45806: inst = 32'hca0ffe7;
      45807: inst = 32'h24822800;
      45808: inst = 32'h10a00000;
      45809: inst = 32'hca00004;
      45810: inst = 32'h38632800;
      45811: inst = 32'h38842800;
      45812: inst = 32'h10a00000;
      45813: inst = 32'hca0b2f9;
      45814: inst = 32'h13e00001;
      45815: inst = 32'hfe0d96a;
      45816: inst = 32'h5be00000;
      45817: inst = 32'h8c50000;
      45818: inst = 32'h24612800;
      45819: inst = 32'h10a0ffff;
      45820: inst = 32'hca0ffe7;
      45821: inst = 32'h24822800;
      45822: inst = 32'h10a00000;
      45823: inst = 32'hca00004;
      45824: inst = 32'h38632800;
      45825: inst = 32'h38842800;
      45826: inst = 32'h10a00000;
      45827: inst = 32'hca0b307;
      45828: inst = 32'h13e00001;
      45829: inst = 32'hfe0d96a;
      45830: inst = 32'h5be00000;
      45831: inst = 32'h8c50000;
      45832: inst = 32'h24612800;
      45833: inst = 32'h10a0ffff;
      45834: inst = 32'hca0ffe7;
      45835: inst = 32'h24822800;
      45836: inst = 32'h10a00000;
      45837: inst = 32'hca00004;
      45838: inst = 32'h38632800;
      45839: inst = 32'h38842800;
      45840: inst = 32'h10a00000;
      45841: inst = 32'hca0b315;
      45842: inst = 32'h13e00001;
      45843: inst = 32'hfe0d96a;
      45844: inst = 32'h5be00000;
      45845: inst = 32'h8c50000;
      45846: inst = 32'h24612800;
      45847: inst = 32'h10a0ffff;
      45848: inst = 32'hca0ffe7;
      45849: inst = 32'h24822800;
      45850: inst = 32'h10a00000;
      45851: inst = 32'hca00004;
      45852: inst = 32'h38632800;
      45853: inst = 32'h38842800;
      45854: inst = 32'h10a00000;
      45855: inst = 32'hca0b323;
      45856: inst = 32'h13e00001;
      45857: inst = 32'hfe0d96a;
      45858: inst = 32'h5be00000;
      45859: inst = 32'h8c50000;
      45860: inst = 32'h24612800;
      45861: inst = 32'h10a0ffff;
      45862: inst = 32'hca0ffe7;
      45863: inst = 32'h24822800;
      45864: inst = 32'h10a00000;
      45865: inst = 32'hca00004;
      45866: inst = 32'h38632800;
      45867: inst = 32'h38842800;
      45868: inst = 32'h10a00000;
      45869: inst = 32'hca0b331;
      45870: inst = 32'h13e00001;
      45871: inst = 32'hfe0d96a;
      45872: inst = 32'h5be00000;
      45873: inst = 32'h8c50000;
      45874: inst = 32'h24612800;
      45875: inst = 32'h10a0ffff;
      45876: inst = 32'hca0ffe7;
      45877: inst = 32'h24822800;
      45878: inst = 32'h10a00000;
      45879: inst = 32'hca00004;
      45880: inst = 32'h38632800;
      45881: inst = 32'h38842800;
      45882: inst = 32'h10a00000;
      45883: inst = 32'hca0b33f;
      45884: inst = 32'h13e00001;
      45885: inst = 32'hfe0d96a;
      45886: inst = 32'h5be00000;
      45887: inst = 32'h8c50000;
      45888: inst = 32'h24612800;
      45889: inst = 32'h10a0ffff;
      45890: inst = 32'hca0ffe7;
      45891: inst = 32'h24822800;
      45892: inst = 32'h10a00000;
      45893: inst = 32'hca00004;
      45894: inst = 32'h38632800;
      45895: inst = 32'h38842800;
      45896: inst = 32'h10a00000;
      45897: inst = 32'hca0b34d;
      45898: inst = 32'h13e00001;
      45899: inst = 32'hfe0d96a;
      45900: inst = 32'h5be00000;
      45901: inst = 32'h8c50000;
      45902: inst = 32'h24612800;
      45903: inst = 32'h10a0ffff;
      45904: inst = 32'hca0ffe7;
      45905: inst = 32'h24822800;
      45906: inst = 32'h10a00000;
      45907: inst = 32'hca00004;
      45908: inst = 32'h38632800;
      45909: inst = 32'h38842800;
      45910: inst = 32'h10a00000;
      45911: inst = 32'hca0b35b;
      45912: inst = 32'h13e00001;
      45913: inst = 32'hfe0d96a;
      45914: inst = 32'h5be00000;
      45915: inst = 32'h8c50000;
      45916: inst = 32'h24612800;
      45917: inst = 32'h10a0ffff;
      45918: inst = 32'hca0ffe7;
      45919: inst = 32'h24822800;
      45920: inst = 32'h10a00000;
      45921: inst = 32'hca00004;
      45922: inst = 32'h38632800;
      45923: inst = 32'h38842800;
      45924: inst = 32'h10a00000;
      45925: inst = 32'hca0b369;
      45926: inst = 32'h13e00001;
      45927: inst = 32'hfe0d96a;
      45928: inst = 32'h5be00000;
      45929: inst = 32'h8c50000;
      45930: inst = 32'h24612800;
      45931: inst = 32'h10a0ffff;
      45932: inst = 32'hca0ffe8;
      45933: inst = 32'h24822800;
      45934: inst = 32'h10a00000;
      45935: inst = 32'hca00004;
      45936: inst = 32'h38632800;
      45937: inst = 32'h38842800;
      45938: inst = 32'h10a00000;
      45939: inst = 32'hca0b377;
      45940: inst = 32'h13e00001;
      45941: inst = 32'hfe0d96a;
      45942: inst = 32'h5be00000;
      45943: inst = 32'h8c50000;
      45944: inst = 32'h24612800;
      45945: inst = 32'h10a0ffff;
      45946: inst = 32'hca0ffe8;
      45947: inst = 32'h24822800;
      45948: inst = 32'h10a00000;
      45949: inst = 32'hca00004;
      45950: inst = 32'h38632800;
      45951: inst = 32'h38842800;
      45952: inst = 32'h10a00000;
      45953: inst = 32'hca0b385;
      45954: inst = 32'h13e00001;
      45955: inst = 32'hfe0d96a;
      45956: inst = 32'h5be00000;
      45957: inst = 32'h8c50000;
      45958: inst = 32'h24612800;
      45959: inst = 32'h10a0ffff;
      45960: inst = 32'hca0ffe8;
      45961: inst = 32'h24822800;
      45962: inst = 32'h10a00000;
      45963: inst = 32'hca00004;
      45964: inst = 32'h38632800;
      45965: inst = 32'h38842800;
      45966: inst = 32'h10a00000;
      45967: inst = 32'hca0b393;
      45968: inst = 32'h13e00001;
      45969: inst = 32'hfe0d96a;
      45970: inst = 32'h5be00000;
      45971: inst = 32'h8c50000;
      45972: inst = 32'h24612800;
      45973: inst = 32'h10a0ffff;
      45974: inst = 32'hca0ffe8;
      45975: inst = 32'h24822800;
      45976: inst = 32'h10a00000;
      45977: inst = 32'hca00004;
      45978: inst = 32'h38632800;
      45979: inst = 32'h38842800;
      45980: inst = 32'h10a00000;
      45981: inst = 32'hca0b3a1;
      45982: inst = 32'h13e00001;
      45983: inst = 32'hfe0d96a;
      45984: inst = 32'h5be00000;
      45985: inst = 32'h8c50000;
      45986: inst = 32'h24612800;
      45987: inst = 32'h10a0ffff;
      45988: inst = 32'hca0ffe8;
      45989: inst = 32'h24822800;
      45990: inst = 32'h10a00000;
      45991: inst = 32'hca00004;
      45992: inst = 32'h38632800;
      45993: inst = 32'h38842800;
      45994: inst = 32'h10a00000;
      45995: inst = 32'hca0b3af;
      45996: inst = 32'h13e00001;
      45997: inst = 32'hfe0d96a;
      45998: inst = 32'h5be00000;
      45999: inst = 32'h8c50000;
      46000: inst = 32'h24612800;
      46001: inst = 32'h10a0ffff;
      46002: inst = 32'hca0ffe8;
      46003: inst = 32'h24822800;
      46004: inst = 32'h10a00000;
      46005: inst = 32'hca00004;
      46006: inst = 32'h38632800;
      46007: inst = 32'h38842800;
      46008: inst = 32'h10a00000;
      46009: inst = 32'hca0b3bd;
      46010: inst = 32'h13e00001;
      46011: inst = 32'hfe0d96a;
      46012: inst = 32'h5be00000;
      46013: inst = 32'h8c50000;
      46014: inst = 32'h24612800;
      46015: inst = 32'h10a0ffff;
      46016: inst = 32'hca0ffe8;
      46017: inst = 32'h24822800;
      46018: inst = 32'h10a00000;
      46019: inst = 32'hca00004;
      46020: inst = 32'h38632800;
      46021: inst = 32'h38842800;
      46022: inst = 32'h10a00000;
      46023: inst = 32'hca0b3cb;
      46024: inst = 32'h13e00001;
      46025: inst = 32'hfe0d96a;
      46026: inst = 32'h5be00000;
      46027: inst = 32'h8c50000;
      46028: inst = 32'h24612800;
      46029: inst = 32'h10a0ffff;
      46030: inst = 32'hca0ffe8;
      46031: inst = 32'h24822800;
      46032: inst = 32'h10a00000;
      46033: inst = 32'hca00004;
      46034: inst = 32'h38632800;
      46035: inst = 32'h38842800;
      46036: inst = 32'h10a00000;
      46037: inst = 32'hca0b3d9;
      46038: inst = 32'h13e00001;
      46039: inst = 32'hfe0d96a;
      46040: inst = 32'h5be00000;
      46041: inst = 32'h8c50000;
      46042: inst = 32'h24612800;
      46043: inst = 32'h10a0ffff;
      46044: inst = 32'hca0ffe8;
      46045: inst = 32'h24822800;
      46046: inst = 32'h10a00000;
      46047: inst = 32'hca00004;
      46048: inst = 32'h38632800;
      46049: inst = 32'h38842800;
      46050: inst = 32'h10a00000;
      46051: inst = 32'hca0b3e7;
      46052: inst = 32'h13e00001;
      46053: inst = 32'hfe0d96a;
      46054: inst = 32'h5be00000;
      46055: inst = 32'h8c50000;
      46056: inst = 32'h24612800;
      46057: inst = 32'h10a0ffff;
      46058: inst = 32'hca0ffe8;
      46059: inst = 32'h24822800;
      46060: inst = 32'h10a00000;
      46061: inst = 32'hca00004;
      46062: inst = 32'h38632800;
      46063: inst = 32'h38842800;
      46064: inst = 32'h10a00000;
      46065: inst = 32'hca0b3f5;
      46066: inst = 32'h13e00001;
      46067: inst = 32'hfe0d96a;
      46068: inst = 32'h5be00000;
      46069: inst = 32'h8c50000;
      46070: inst = 32'h24612800;
      46071: inst = 32'h10a0ffff;
      46072: inst = 32'hca0ffe8;
      46073: inst = 32'h24822800;
      46074: inst = 32'h10a00000;
      46075: inst = 32'hca00004;
      46076: inst = 32'h38632800;
      46077: inst = 32'h38842800;
      46078: inst = 32'h10a00000;
      46079: inst = 32'hca0b403;
      46080: inst = 32'h13e00001;
      46081: inst = 32'hfe0d96a;
      46082: inst = 32'h5be00000;
      46083: inst = 32'h8c50000;
      46084: inst = 32'h24612800;
      46085: inst = 32'h10a0ffff;
      46086: inst = 32'hca0ffe8;
      46087: inst = 32'h24822800;
      46088: inst = 32'h10a00000;
      46089: inst = 32'hca00004;
      46090: inst = 32'h38632800;
      46091: inst = 32'h38842800;
      46092: inst = 32'h10a00000;
      46093: inst = 32'hca0b411;
      46094: inst = 32'h13e00001;
      46095: inst = 32'hfe0d96a;
      46096: inst = 32'h5be00000;
      46097: inst = 32'h8c50000;
      46098: inst = 32'h24612800;
      46099: inst = 32'h10a0ffff;
      46100: inst = 32'hca0ffe8;
      46101: inst = 32'h24822800;
      46102: inst = 32'h10a00000;
      46103: inst = 32'hca00004;
      46104: inst = 32'h38632800;
      46105: inst = 32'h38842800;
      46106: inst = 32'h10a00000;
      46107: inst = 32'hca0b41f;
      46108: inst = 32'h13e00001;
      46109: inst = 32'hfe0d96a;
      46110: inst = 32'h5be00000;
      46111: inst = 32'h8c50000;
      46112: inst = 32'h24612800;
      46113: inst = 32'h10a0ffff;
      46114: inst = 32'hca0ffe8;
      46115: inst = 32'h24822800;
      46116: inst = 32'h10a00000;
      46117: inst = 32'hca00004;
      46118: inst = 32'h38632800;
      46119: inst = 32'h38842800;
      46120: inst = 32'h10a00000;
      46121: inst = 32'hca0b42d;
      46122: inst = 32'h13e00001;
      46123: inst = 32'hfe0d96a;
      46124: inst = 32'h5be00000;
      46125: inst = 32'h8c50000;
      46126: inst = 32'h24612800;
      46127: inst = 32'h10a0ffff;
      46128: inst = 32'hca0ffe8;
      46129: inst = 32'h24822800;
      46130: inst = 32'h10a00000;
      46131: inst = 32'hca00004;
      46132: inst = 32'h38632800;
      46133: inst = 32'h38842800;
      46134: inst = 32'h10a00000;
      46135: inst = 32'hca0b43b;
      46136: inst = 32'h13e00001;
      46137: inst = 32'hfe0d96a;
      46138: inst = 32'h5be00000;
      46139: inst = 32'h8c50000;
      46140: inst = 32'h24612800;
      46141: inst = 32'h10a0ffff;
      46142: inst = 32'hca0ffe8;
      46143: inst = 32'h24822800;
      46144: inst = 32'h10a00000;
      46145: inst = 32'hca00004;
      46146: inst = 32'h38632800;
      46147: inst = 32'h38842800;
      46148: inst = 32'h10a00000;
      46149: inst = 32'hca0b449;
      46150: inst = 32'h13e00001;
      46151: inst = 32'hfe0d96a;
      46152: inst = 32'h5be00000;
      46153: inst = 32'h8c50000;
      46154: inst = 32'h24612800;
      46155: inst = 32'h10a0ffff;
      46156: inst = 32'hca0ffe8;
      46157: inst = 32'h24822800;
      46158: inst = 32'h10a00000;
      46159: inst = 32'hca00004;
      46160: inst = 32'h38632800;
      46161: inst = 32'h38842800;
      46162: inst = 32'h10a00000;
      46163: inst = 32'hca0b457;
      46164: inst = 32'h13e00001;
      46165: inst = 32'hfe0d96a;
      46166: inst = 32'h5be00000;
      46167: inst = 32'h8c50000;
      46168: inst = 32'h24612800;
      46169: inst = 32'h10a0ffff;
      46170: inst = 32'hca0ffe8;
      46171: inst = 32'h24822800;
      46172: inst = 32'h10a00000;
      46173: inst = 32'hca00004;
      46174: inst = 32'h38632800;
      46175: inst = 32'h38842800;
      46176: inst = 32'h10a00000;
      46177: inst = 32'hca0b465;
      46178: inst = 32'h13e00001;
      46179: inst = 32'hfe0d96a;
      46180: inst = 32'h5be00000;
      46181: inst = 32'h8c50000;
      46182: inst = 32'h24612800;
      46183: inst = 32'h10a0ffff;
      46184: inst = 32'hca0ffe8;
      46185: inst = 32'h24822800;
      46186: inst = 32'h10a00000;
      46187: inst = 32'hca00004;
      46188: inst = 32'h38632800;
      46189: inst = 32'h38842800;
      46190: inst = 32'h10a00000;
      46191: inst = 32'hca0b473;
      46192: inst = 32'h13e00001;
      46193: inst = 32'hfe0d96a;
      46194: inst = 32'h5be00000;
      46195: inst = 32'h8c50000;
      46196: inst = 32'h24612800;
      46197: inst = 32'h10a0ffff;
      46198: inst = 32'hca0ffe8;
      46199: inst = 32'h24822800;
      46200: inst = 32'h10a00000;
      46201: inst = 32'hca00004;
      46202: inst = 32'h38632800;
      46203: inst = 32'h38842800;
      46204: inst = 32'h10a00000;
      46205: inst = 32'hca0b481;
      46206: inst = 32'h13e00001;
      46207: inst = 32'hfe0d96a;
      46208: inst = 32'h5be00000;
      46209: inst = 32'h8c50000;
      46210: inst = 32'h24612800;
      46211: inst = 32'h10a0ffff;
      46212: inst = 32'hca0ffe8;
      46213: inst = 32'h24822800;
      46214: inst = 32'h10a00000;
      46215: inst = 32'hca00004;
      46216: inst = 32'h38632800;
      46217: inst = 32'h38842800;
      46218: inst = 32'h10a00000;
      46219: inst = 32'hca0b48f;
      46220: inst = 32'h13e00001;
      46221: inst = 32'hfe0d96a;
      46222: inst = 32'h5be00000;
      46223: inst = 32'h8c50000;
      46224: inst = 32'h24612800;
      46225: inst = 32'h10a0ffff;
      46226: inst = 32'hca0ffe8;
      46227: inst = 32'h24822800;
      46228: inst = 32'h10a00000;
      46229: inst = 32'hca00004;
      46230: inst = 32'h38632800;
      46231: inst = 32'h38842800;
      46232: inst = 32'h10a00000;
      46233: inst = 32'hca0b49d;
      46234: inst = 32'h13e00001;
      46235: inst = 32'hfe0d96a;
      46236: inst = 32'h5be00000;
      46237: inst = 32'h8c50000;
      46238: inst = 32'h24612800;
      46239: inst = 32'h10a0ffff;
      46240: inst = 32'hca0ffe8;
      46241: inst = 32'h24822800;
      46242: inst = 32'h10a00000;
      46243: inst = 32'hca00004;
      46244: inst = 32'h38632800;
      46245: inst = 32'h38842800;
      46246: inst = 32'h10a00000;
      46247: inst = 32'hca0b4ab;
      46248: inst = 32'h13e00001;
      46249: inst = 32'hfe0d96a;
      46250: inst = 32'h5be00000;
      46251: inst = 32'h8c50000;
      46252: inst = 32'h24612800;
      46253: inst = 32'h10a0ffff;
      46254: inst = 32'hca0ffe8;
      46255: inst = 32'h24822800;
      46256: inst = 32'h10a00000;
      46257: inst = 32'hca00004;
      46258: inst = 32'h38632800;
      46259: inst = 32'h38842800;
      46260: inst = 32'h10a00000;
      46261: inst = 32'hca0b4b9;
      46262: inst = 32'h13e00001;
      46263: inst = 32'hfe0d96a;
      46264: inst = 32'h5be00000;
      46265: inst = 32'h8c50000;
      46266: inst = 32'h24612800;
      46267: inst = 32'h10a0ffff;
      46268: inst = 32'hca0ffe8;
      46269: inst = 32'h24822800;
      46270: inst = 32'h10a00000;
      46271: inst = 32'hca00004;
      46272: inst = 32'h38632800;
      46273: inst = 32'h38842800;
      46274: inst = 32'h10a00000;
      46275: inst = 32'hca0b4c7;
      46276: inst = 32'h13e00001;
      46277: inst = 32'hfe0d96a;
      46278: inst = 32'h5be00000;
      46279: inst = 32'h8c50000;
      46280: inst = 32'h24612800;
      46281: inst = 32'h10a0ffff;
      46282: inst = 32'hca0ffe8;
      46283: inst = 32'h24822800;
      46284: inst = 32'h10a00000;
      46285: inst = 32'hca00004;
      46286: inst = 32'h38632800;
      46287: inst = 32'h38842800;
      46288: inst = 32'h10a00000;
      46289: inst = 32'hca0b4d5;
      46290: inst = 32'h13e00001;
      46291: inst = 32'hfe0d96a;
      46292: inst = 32'h5be00000;
      46293: inst = 32'h8c50000;
      46294: inst = 32'h24612800;
      46295: inst = 32'h10a0ffff;
      46296: inst = 32'hca0ffe8;
      46297: inst = 32'h24822800;
      46298: inst = 32'h10a00000;
      46299: inst = 32'hca00004;
      46300: inst = 32'h38632800;
      46301: inst = 32'h38842800;
      46302: inst = 32'h10a00000;
      46303: inst = 32'hca0b4e3;
      46304: inst = 32'h13e00001;
      46305: inst = 32'hfe0d96a;
      46306: inst = 32'h5be00000;
      46307: inst = 32'h8c50000;
      46308: inst = 32'h24612800;
      46309: inst = 32'h10a0ffff;
      46310: inst = 32'hca0ffe8;
      46311: inst = 32'h24822800;
      46312: inst = 32'h10a00000;
      46313: inst = 32'hca00004;
      46314: inst = 32'h38632800;
      46315: inst = 32'h38842800;
      46316: inst = 32'h10a00000;
      46317: inst = 32'hca0b4f1;
      46318: inst = 32'h13e00001;
      46319: inst = 32'hfe0d96a;
      46320: inst = 32'h5be00000;
      46321: inst = 32'h8c50000;
      46322: inst = 32'h24612800;
      46323: inst = 32'h10a0ffff;
      46324: inst = 32'hca0ffe8;
      46325: inst = 32'h24822800;
      46326: inst = 32'h10a00000;
      46327: inst = 32'hca00004;
      46328: inst = 32'h38632800;
      46329: inst = 32'h38842800;
      46330: inst = 32'h10a00000;
      46331: inst = 32'hca0b4ff;
      46332: inst = 32'h13e00001;
      46333: inst = 32'hfe0d96a;
      46334: inst = 32'h5be00000;
      46335: inst = 32'h8c50000;
      46336: inst = 32'h24612800;
      46337: inst = 32'h10a0ffff;
      46338: inst = 32'hca0ffe8;
      46339: inst = 32'h24822800;
      46340: inst = 32'h10a00000;
      46341: inst = 32'hca00004;
      46342: inst = 32'h38632800;
      46343: inst = 32'h38842800;
      46344: inst = 32'h10a00000;
      46345: inst = 32'hca0b50d;
      46346: inst = 32'h13e00001;
      46347: inst = 32'hfe0d96a;
      46348: inst = 32'h5be00000;
      46349: inst = 32'h8c50000;
      46350: inst = 32'h24612800;
      46351: inst = 32'h10a0ffff;
      46352: inst = 32'hca0ffe8;
      46353: inst = 32'h24822800;
      46354: inst = 32'h10a00000;
      46355: inst = 32'hca00004;
      46356: inst = 32'h38632800;
      46357: inst = 32'h38842800;
      46358: inst = 32'h10a00000;
      46359: inst = 32'hca0b51b;
      46360: inst = 32'h13e00001;
      46361: inst = 32'hfe0d96a;
      46362: inst = 32'h5be00000;
      46363: inst = 32'h8c50000;
      46364: inst = 32'h24612800;
      46365: inst = 32'h10a0ffff;
      46366: inst = 32'hca0ffe8;
      46367: inst = 32'h24822800;
      46368: inst = 32'h10a00000;
      46369: inst = 32'hca00004;
      46370: inst = 32'h38632800;
      46371: inst = 32'h38842800;
      46372: inst = 32'h10a00000;
      46373: inst = 32'hca0b529;
      46374: inst = 32'h13e00001;
      46375: inst = 32'hfe0d96a;
      46376: inst = 32'h5be00000;
      46377: inst = 32'h8c50000;
      46378: inst = 32'h24612800;
      46379: inst = 32'h10a0ffff;
      46380: inst = 32'hca0ffe8;
      46381: inst = 32'h24822800;
      46382: inst = 32'h10a00000;
      46383: inst = 32'hca00004;
      46384: inst = 32'h38632800;
      46385: inst = 32'h38842800;
      46386: inst = 32'h10a00000;
      46387: inst = 32'hca0b537;
      46388: inst = 32'h13e00001;
      46389: inst = 32'hfe0d96a;
      46390: inst = 32'h5be00000;
      46391: inst = 32'h8c50000;
      46392: inst = 32'h24612800;
      46393: inst = 32'h10a0ffff;
      46394: inst = 32'hca0ffe8;
      46395: inst = 32'h24822800;
      46396: inst = 32'h10a00000;
      46397: inst = 32'hca00004;
      46398: inst = 32'h38632800;
      46399: inst = 32'h38842800;
      46400: inst = 32'h10a00000;
      46401: inst = 32'hca0b545;
      46402: inst = 32'h13e00001;
      46403: inst = 32'hfe0d96a;
      46404: inst = 32'h5be00000;
      46405: inst = 32'h8c50000;
      46406: inst = 32'h24612800;
      46407: inst = 32'h10a0ffff;
      46408: inst = 32'hca0ffe8;
      46409: inst = 32'h24822800;
      46410: inst = 32'h10a00000;
      46411: inst = 32'hca00004;
      46412: inst = 32'h38632800;
      46413: inst = 32'h38842800;
      46414: inst = 32'h10a00000;
      46415: inst = 32'hca0b553;
      46416: inst = 32'h13e00001;
      46417: inst = 32'hfe0d96a;
      46418: inst = 32'h5be00000;
      46419: inst = 32'h8c50000;
      46420: inst = 32'h24612800;
      46421: inst = 32'h10a0ffff;
      46422: inst = 32'hca0ffe8;
      46423: inst = 32'h24822800;
      46424: inst = 32'h10a00000;
      46425: inst = 32'hca00004;
      46426: inst = 32'h38632800;
      46427: inst = 32'h38842800;
      46428: inst = 32'h10a00000;
      46429: inst = 32'hca0b561;
      46430: inst = 32'h13e00001;
      46431: inst = 32'hfe0d96a;
      46432: inst = 32'h5be00000;
      46433: inst = 32'h8c50000;
      46434: inst = 32'h24612800;
      46435: inst = 32'h10a0ffff;
      46436: inst = 32'hca0ffe8;
      46437: inst = 32'h24822800;
      46438: inst = 32'h10a00000;
      46439: inst = 32'hca00004;
      46440: inst = 32'h38632800;
      46441: inst = 32'h38842800;
      46442: inst = 32'h10a00000;
      46443: inst = 32'hca0b56f;
      46444: inst = 32'h13e00001;
      46445: inst = 32'hfe0d96a;
      46446: inst = 32'h5be00000;
      46447: inst = 32'h8c50000;
      46448: inst = 32'h24612800;
      46449: inst = 32'h10a0ffff;
      46450: inst = 32'hca0ffe8;
      46451: inst = 32'h24822800;
      46452: inst = 32'h10a00000;
      46453: inst = 32'hca00004;
      46454: inst = 32'h38632800;
      46455: inst = 32'h38842800;
      46456: inst = 32'h10a00000;
      46457: inst = 32'hca0b57d;
      46458: inst = 32'h13e00001;
      46459: inst = 32'hfe0d96a;
      46460: inst = 32'h5be00000;
      46461: inst = 32'h8c50000;
      46462: inst = 32'h24612800;
      46463: inst = 32'h10a0ffff;
      46464: inst = 32'hca0ffe8;
      46465: inst = 32'h24822800;
      46466: inst = 32'h10a00000;
      46467: inst = 32'hca00004;
      46468: inst = 32'h38632800;
      46469: inst = 32'h38842800;
      46470: inst = 32'h10a00000;
      46471: inst = 32'hca0b58b;
      46472: inst = 32'h13e00001;
      46473: inst = 32'hfe0d96a;
      46474: inst = 32'h5be00000;
      46475: inst = 32'h8c50000;
      46476: inst = 32'h24612800;
      46477: inst = 32'h10a0ffff;
      46478: inst = 32'hca0ffe8;
      46479: inst = 32'h24822800;
      46480: inst = 32'h10a00000;
      46481: inst = 32'hca00004;
      46482: inst = 32'h38632800;
      46483: inst = 32'h38842800;
      46484: inst = 32'h10a00000;
      46485: inst = 32'hca0b599;
      46486: inst = 32'h13e00001;
      46487: inst = 32'hfe0d96a;
      46488: inst = 32'h5be00000;
      46489: inst = 32'h8c50000;
      46490: inst = 32'h24612800;
      46491: inst = 32'h10a0ffff;
      46492: inst = 32'hca0ffe8;
      46493: inst = 32'h24822800;
      46494: inst = 32'h10a00000;
      46495: inst = 32'hca00004;
      46496: inst = 32'h38632800;
      46497: inst = 32'h38842800;
      46498: inst = 32'h10a00000;
      46499: inst = 32'hca0b5a7;
      46500: inst = 32'h13e00001;
      46501: inst = 32'hfe0d96a;
      46502: inst = 32'h5be00000;
      46503: inst = 32'h8c50000;
      46504: inst = 32'h24612800;
      46505: inst = 32'h10a0ffff;
      46506: inst = 32'hca0ffe8;
      46507: inst = 32'h24822800;
      46508: inst = 32'h10a00000;
      46509: inst = 32'hca00004;
      46510: inst = 32'h38632800;
      46511: inst = 32'h38842800;
      46512: inst = 32'h10a00000;
      46513: inst = 32'hca0b5b5;
      46514: inst = 32'h13e00001;
      46515: inst = 32'hfe0d96a;
      46516: inst = 32'h5be00000;
      46517: inst = 32'h8c50000;
      46518: inst = 32'h24612800;
      46519: inst = 32'h10a0ffff;
      46520: inst = 32'hca0ffe8;
      46521: inst = 32'h24822800;
      46522: inst = 32'h10a00000;
      46523: inst = 32'hca00004;
      46524: inst = 32'h38632800;
      46525: inst = 32'h38842800;
      46526: inst = 32'h10a00000;
      46527: inst = 32'hca0b5c3;
      46528: inst = 32'h13e00001;
      46529: inst = 32'hfe0d96a;
      46530: inst = 32'h5be00000;
      46531: inst = 32'h8c50000;
      46532: inst = 32'h24612800;
      46533: inst = 32'h10a0ffff;
      46534: inst = 32'hca0ffe8;
      46535: inst = 32'h24822800;
      46536: inst = 32'h10a00000;
      46537: inst = 32'hca00004;
      46538: inst = 32'h38632800;
      46539: inst = 32'h38842800;
      46540: inst = 32'h10a00000;
      46541: inst = 32'hca0b5d1;
      46542: inst = 32'h13e00001;
      46543: inst = 32'hfe0d96a;
      46544: inst = 32'h5be00000;
      46545: inst = 32'h8c50000;
      46546: inst = 32'h24612800;
      46547: inst = 32'h10a0ffff;
      46548: inst = 32'hca0ffe8;
      46549: inst = 32'h24822800;
      46550: inst = 32'h10a00000;
      46551: inst = 32'hca00004;
      46552: inst = 32'h38632800;
      46553: inst = 32'h38842800;
      46554: inst = 32'h10a00000;
      46555: inst = 32'hca0b5df;
      46556: inst = 32'h13e00001;
      46557: inst = 32'hfe0d96a;
      46558: inst = 32'h5be00000;
      46559: inst = 32'h8c50000;
      46560: inst = 32'h24612800;
      46561: inst = 32'h10a0ffff;
      46562: inst = 32'hca0ffe8;
      46563: inst = 32'h24822800;
      46564: inst = 32'h10a00000;
      46565: inst = 32'hca00004;
      46566: inst = 32'h38632800;
      46567: inst = 32'h38842800;
      46568: inst = 32'h10a00000;
      46569: inst = 32'hca0b5ed;
      46570: inst = 32'h13e00001;
      46571: inst = 32'hfe0d96a;
      46572: inst = 32'h5be00000;
      46573: inst = 32'h8c50000;
      46574: inst = 32'h24612800;
      46575: inst = 32'h10a0ffff;
      46576: inst = 32'hca0ffe8;
      46577: inst = 32'h24822800;
      46578: inst = 32'h10a00000;
      46579: inst = 32'hca00004;
      46580: inst = 32'h38632800;
      46581: inst = 32'h38842800;
      46582: inst = 32'h10a00000;
      46583: inst = 32'hca0b5fb;
      46584: inst = 32'h13e00001;
      46585: inst = 32'hfe0d96a;
      46586: inst = 32'h5be00000;
      46587: inst = 32'h8c50000;
      46588: inst = 32'h24612800;
      46589: inst = 32'h10a0ffff;
      46590: inst = 32'hca0ffe8;
      46591: inst = 32'h24822800;
      46592: inst = 32'h10a00000;
      46593: inst = 32'hca00004;
      46594: inst = 32'h38632800;
      46595: inst = 32'h38842800;
      46596: inst = 32'h10a00000;
      46597: inst = 32'hca0b609;
      46598: inst = 32'h13e00001;
      46599: inst = 32'hfe0d96a;
      46600: inst = 32'h5be00000;
      46601: inst = 32'h8c50000;
      46602: inst = 32'h24612800;
      46603: inst = 32'h10a0ffff;
      46604: inst = 32'hca0ffe8;
      46605: inst = 32'h24822800;
      46606: inst = 32'h10a00000;
      46607: inst = 32'hca00004;
      46608: inst = 32'h38632800;
      46609: inst = 32'h38842800;
      46610: inst = 32'h10a00000;
      46611: inst = 32'hca0b617;
      46612: inst = 32'h13e00001;
      46613: inst = 32'hfe0d96a;
      46614: inst = 32'h5be00000;
      46615: inst = 32'h8c50000;
      46616: inst = 32'h24612800;
      46617: inst = 32'h10a0ffff;
      46618: inst = 32'hca0ffe8;
      46619: inst = 32'h24822800;
      46620: inst = 32'h10a00000;
      46621: inst = 32'hca00004;
      46622: inst = 32'h38632800;
      46623: inst = 32'h38842800;
      46624: inst = 32'h10a00000;
      46625: inst = 32'hca0b625;
      46626: inst = 32'h13e00001;
      46627: inst = 32'hfe0d96a;
      46628: inst = 32'h5be00000;
      46629: inst = 32'h8c50000;
      46630: inst = 32'h24612800;
      46631: inst = 32'h10a0ffff;
      46632: inst = 32'hca0ffe8;
      46633: inst = 32'h24822800;
      46634: inst = 32'h10a00000;
      46635: inst = 32'hca00004;
      46636: inst = 32'h38632800;
      46637: inst = 32'h38842800;
      46638: inst = 32'h10a00000;
      46639: inst = 32'hca0b633;
      46640: inst = 32'h13e00001;
      46641: inst = 32'hfe0d96a;
      46642: inst = 32'h5be00000;
      46643: inst = 32'h8c50000;
      46644: inst = 32'h24612800;
      46645: inst = 32'h10a0ffff;
      46646: inst = 32'hca0ffe8;
      46647: inst = 32'h24822800;
      46648: inst = 32'h10a00000;
      46649: inst = 32'hca00004;
      46650: inst = 32'h38632800;
      46651: inst = 32'h38842800;
      46652: inst = 32'h10a00000;
      46653: inst = 32'hca0b641;
      46654: inst = 32'h13e00001;
      46655: inst = 32'hfe0d96a;
      46656: inst = 32'h5be00000;
      46657: inst = 32'h8c50000;
      46658: inst = 32'h24612800;
      46659: inst = 32'h10a0ffff;
      46660: inst = 32'hca0ffe8;
      46661: inst = 32'h24822800;
      46662: inst = 32'h10a00000;
      46663: inst = 32'hca00004;
      46664: inst = 32'h38632800;
      46665: inst = 32'h38842800;
      46666: inst = 32'h10a00000;
      46667: inst = 32'hca0b64f;
      46668: inst = 32'h13e00001;
      46669: inst = 32'hfe0d96a;
      46670: inst = 32'h5be00000;
      46671: inst = 32'h8c50000;
      46672: inst = 32'h24612800;
      46673: inst = 32'h10a0ffff;
      46674: inst = 32'hca0ffe8;
      46675: inst = 32'h24822800;
      46676: inst = 32'h10a00000;
      46677: inst = 32'hca00004;
      46678: inst = 32'h38632800;
      46679: inst = 32'h38842800;
      46680: inst = 32'h10a00000;
      46681: inst = 32'hca0b65d;
      46682: inst = 32'h13e00001;
      46683: inst = 32'hfe0d96a;
      46684: inst = 32'h5be00000;
      46685: inst = 32'h8c50000;
      46686: inst = 32'h24612800;
      46687: inst = 32'h10a0ffff;
      46688: inst = 32'hca0ffe8;
      46689: inst = 32'h24822800;
      46690: inst = 32'h10a00000;
      46691: inst = 32'hca00004;
      46692: inst = 32'h38632800;
      46693: inst = 32'h38842800;
      46694: inst = 32'h10a00000;
      46695: inst = 32'hca0b66b;
      46696: inst = 32'h13e00001;
      46697: inst = 32'hfe0d96a;
      46698: inst = 32'h5be00000;
      46699: inst = 32'h8c50000;
      46700: inst = 32'h24612800;
      46701: inst = 32'h10a0ffff;
      46702: inst = 32'hca0ffe8;
      46703: inst = 32'h24822800;
      46704: inst = 32'h10a00000;
      46705: inst = 32'hca00004;
      46706: inst = 32'h38632800;
      46707: inst = 32'h38842800;
      46708: inst = 32'h10a00000;
      46709: inst = 32'hca0b679;
      46710: inst = 32'h13e00001;
      46711: inst = 32'hfe0d96a;
      46712: inst = 32'h5be00000;
      46713: inst = 32'h8c50000;
      46714: inst = 32'h24612800;
      46715: inst = 32'h10a0ffff;
      46716: inst = 32'hca0ffe8;
      46717: inst = 32'h24822800;
      46718: inst = 32'h10a00000;
      46719: inst = 32'hca00004;
      46720: inst = 32'h38632800;
      46721: inst = 32'h38842800;
      46722: inst = 32'h10a00000;
      46723: inst = 32'hca0b687;
      46724: inst = 32'h13e00001;
      46725: inst = 32'hfe0d96a;
      46726: inst = 32'h5be00000;
      46727: inst = 32'h8c50000;
      46728: inst = 32'h24612800;
      46729: inst = 32'h10a0ffff;
      46730: inst = 32'hca0ffe8;
      46731: inst = 32'h24822800;
      46732: inst = 32'h10a00000;
      46733: inst = 32'hca00004;
      46734: inst = 32'h38632800;
      46735: inst = 32'h38842800;
      46736: inst = 32'h10a00000;
      46737: inst = 32'hca0b695;
      46738: inst = 32'h13e00001;
      46739: inst = 32'hfe0d96a;
      46740: inst = 32'h5be00000;
      46741: inst = 32'h8c50000;
      46742: inst = 32'h24612800;
      46743: inst = 32'h10a0ffff;
      46744: inst = 32'hca0ffe8;
      46745: inst = 32'h24822800;
      46746: inst = 32'h10a00000;
      46747: inst = 32'hca00004;
      46748: inst = 32'h38632800;
      46749: inst = 32'h38842800;
      46750: inst = 32'h10a00000;
      46751: inst = 32'hca0b6a3;
      46752: inst = 32'h13e00001;
      46753: inst = 32'hfe0d96a;
      46754: inst = 32'h5be00000;
      46755: inst = 32'h8c50000;
      46756: inst = 32'h24612800;
      46757: inst = 32'h10a0ffff;
      46758: inst = 32'hca0ffe8;
      46759: inst = 32'h24822800;
      46760: inst = 32'h10a00000;
      46761: inst = 32'hca00004;
      46762: inst = 32'h38632800;
      46763: inst = 32'h38842800;
      46764: inst = 32'h10a00000;
      46765: inst = 32'hca0b6b1;
      46766: inst = 32'h13e00001;
      46767: inst = 32'hfe0d96a;
      46768: inst = 32'h5be00000;
      46769: inst = 32'h8c50000;
      46770: inst = 32'h24612800;
      46771: inst = 32'h10a0ffff;
      46772: inst = 32'hca0ffe8;
      46773: inst = 32'h24822800;
      46774: inst = 32'h10a00000;
      46775: inst = 32'hca00004;
      46776: inst = 32'h38632800;
      46777: inst = 32'h38842800;
      46778: inst = 32'h10a00000;
      46779: inst = 32'hca0b6bf;
      46780: inst = 32'h13e00001;
      46781: inst = 32'hfe0d96a;
      46782: inst = 32'h5be00000;
      46783: inst = 32'h8c50000;
      46784: inst = 32'h24612800;
      46785: inst = 32'h10a0ffff;
      46786: inst = 32'hca0ffe8;
      46787: inst = 32'h24822800;
      46788: inst = 32'h10a00000;
      46789: inst = 32'hca00004;
      46790: inst = 32'h38632800;
      46791: inst = 32'h38842800;
      46792: inst = 32'h10a00000;
      46793: inst = 32'hca0b6cd;
      46794: inst = 32'h13e00001;
      46795: inst = 32'hfe0d96a;
      46796: inst = 32'h5be00000;
      46797: inst = 32'h8c50000;
      46798: inst = 32'h24612800;
      46799: inst = 32'h10a0ffff;
      46800: inst = 32'hca0ffe8;
      46801: inst = 32'h24822800;
      46802: inst = 32'h10a00000;
      46803: inst = 32'hca00004;
      46804: inst = 32'h38632800;
      46805: inst = 32'h38842800;
      46806: inst = 32'h10a00000;
      46807: inst = 32'hca0b6db;
      46808: inst = 32'h13e00001;
      46809: inst = 32'hfe0d96a;
      46810: inst = 32'h5be00000;
      46811: inst = 32'h8c50000;
      46812: inst = 32'h24612800;
      46813: inst = 32'h10a0ffff;
      46814: inst = 32'hca0ffe8;
      46815: inst = 32'h24822800;
      46816: inst = 32'h10a00000;
      46817: inst = 32'hca00004;
      46818: inst = 32'h38632800;
      46819: inst = 32'h38842800;
      46820: inst = 32'h10a00000;
      46821: inst = 32'hca0b6e9;
      46822: inst = 32'h13e00001;
      46823: inst = 32'hfe0d96a;
      46824: inst = 32'h5be00000;
      46825: inst = 32'h8c50000;
      46826: inst = 32'h24612800;
      46827: inst = 32'h10a0ffff;
      46828: inst = 32'hca0ffe8;
      46829: inst = 32'h24822800;
      46830: inst = 32'h10a00000;
      46831: inst = 32'hca00004;
      46832: inst = 32'h38632800;
      46833: inst = 32'h38842800;
      46834: inst = 32'h10a00000;
      46835: inst = 32'hca0b6f7;
      46836: inst = 32'h13e00001;
      46837: inst = 32'hfe0d96a;
      46838: inst = 32'h5be00000;
      46839: inst = 32'h8c50000;
      46840: inst = 32'h24612800;
      46841: inst = 32'h10a0ffff;
      46842: inst = 32'hca0ffe8;
      46843: inst = 32'h24822800;
      46844: inst = 32'h10a00000;
      46845: inst = 32'hca00004;
      46846: inst = 32'h38632800;
      46847: inst = 32'h38842800;
      46848: inst = 32'h10a00000;
      46849: inst = 32'hca0b705;
      46850: inst = 32'h13e00001;
      46851: inst = 32'hfe0d96a;
      46852: inst = 32'h5be00000;
      46853: inst = 32'h8c50000;
      46854: inst = 32'h24612800;
      46855: inst = 32'h10a0ffff;
      46856: inst = 32'hca0ffe8;
      46857: inst = 32'h24822800;
      46858: inst = 32'h10a00000;
      46859: inst = 32'hca00004;
      46860: inst = 32'h38632800;
      46861: inst = 32'h38842800;
      46862: inst = 32'h10a00000;
      46863: inst = 32'hca0b713;
      46864: inst = 32'h13e00001;
      46865: inst = 32'hfe0d96a;
      46866: inst = 32'h5be00000;
      46867: inst = 32'h8c50000;
      46868: inst = 32'h24612800;
      46869: inst = 32'h10a0ffff;
      46870: inst = 32'hca0ffe8;
      46871: inst = 32'h24822800;
      46872: inst = 32'h10a00000;
      46873: inst = 32'hca00004;
      46874: inst = 32'h38632800;
      46875: inst = 32'h38842800;
      46876: inst = 32'h10a00000;
      46877: inst = 32'hca0b721;
      46878: inst = 32'h13e00001;
      46879: inst = 32'hfe0d96a;
      46880: inst = 32'h5be00000;
      46881: inst = 32'h8c50000;
      46882: inst = 32'h24612800;
      46883: inst = 32'h10a0ffff;
      46884: inst = 32'hca0ffe8;
      46885: inst = 32'h24822800;
      46886: inst = 32'h10a00000;
      46887: inst = 32'hca00004;
      46888: inst = 32'h38632800;
      46889: inst = 32'h38842800;
      46890: inst = 32'h10a00000;
      46891: inst = 32'hca0b72f;
      46892: inst = 32'h13e00001;
      46893: inst = 32'hfe0d96a;
      46894: inst = 32'h5be00000;
      46895: inst = 32'h8c50000;
      46896: inst = 32'h24612800;
      46897: inst = 32'h10a0ffff;
      46898: inst = 32'hca0ffe8;
      46899: inst = 32'h24822800;
      46900: inst = 32'h10a00000;
      46901: inst = 32'hca00004;
      46902: inst = 32'h38632800;
      46903: inst = 32'h38842800;
      46904: inst = 32'h10a00000;
      46905: inst = 32'hca0b73d;
      46906: inst = 32'h13e00001;
      46907: inst = 32'hfe0d96a;
      46908: inst = 32'h5be00000;
      46909: inst = 32'h8c50000;
      46910: inst = 32'h24612800;
      46911: inst = 32'h10a0ffff;
      46912: inst = 32'hca0ffe8;
      46913: inst = 32'h24822800;
      46914: inst = 32'h10a00000;
      46915: inst = 32'hca00004;
      46916: inst = 32'h38632800;
      46917: inst = 32'h38842800;
      46918: inst = 32'h10a00000;
      46919: inst = 32'hca0b74b;
      46920: inst = 32'h13e00001;
      46921: inst = 32'hfe0d96a;
      46922: inst = 32'h5be00000;
      46923: inst = 32'h8c50000;
      46924: inst = 32'h24612800;
      46925: inst = 32'h10a0ffff;
      46926: inst = 32'hca0ffe8;
      46927: inst = 32'h24822800;
      46928: inst = 32'h10a00000;
      46929: inst = 32'hca00004;
      46930: inst = 32'h38632800;
      46931: inst = 32'h38842800;
      46932: inst = 32'h10a00000;
      46933: inst = 32'hca0b759;
      46934: inst = 32'h13e00001;
      46935: inst = 32'hfe0d96a;
      46936: inst = 32'h5be00000;
      46937: inst = 32'h8c50000;
      46938: inst = 32'h24612800;
      46939: inst = 32'h10a0ffff;
      46940: inst = 32'hca0ffe8;
      46941: inst = 32'h24822800;
      46942: inst = 32'h10a00000;
      46943: inst = 32'hca00004;
      46944: inst = 32'h38632800;
      46945: inst = 32'h38842800;
      46946: inst = 32'h10a00000;
      46947: inst = 32'hca0b767;
      46948: inst = 32'h13e00001;
      46949: inst = 32'hfe0d96a;
      46950: inst = 32'h5be00000;
      46951: inst = 32'h8c50000;
      46952: inst = 32'h24612800;
      46953: inst = 32'h10a0ffff;
      46954: inst = 32'hca0ffe8;
      46955: inst = 32'h24822800;
      46956: inst = 32'h10a00000;
      46957: inst = 32'hca00004;
      46958: inst = 32'h38632800;
      46959: inst = 32'h38842800;
      46960: inst = 32'h10a00000;
      46961: inst = 32'hca0b775;
      46962: inst = 32'h13e00001;
      46963: inst = 32'hfe0d96a;
      46964: inst = 32'h5be00000;
      46965: inst = 32'h8c50000;
      46966: inst = 32'h24612800;
      46967: inst = 32'h10a0ffff;
      46968: inst = 32'hca0ffe8;
      46969: inst = 32'h24822800;
      46970: inst = 32'h10a00000;
      46971: inst = 32'hca00004;
      46972: inst = 32'h38632800;
      46973: inst = 32'h38842800;
      46974: inst = 32'h10a00000;
      46975: inst = 32'hca0b783;
      46976: inst = 32'h13e00001;
      46977: inst = 32'hfe0d96a;
      46978: inst = 32'h5be00000;
      46979: inst = 32'h8c50000;
      46980: inst = 32'h24612800;
      46981: inst = 32'h10a0ffff;
      46982: inst = 32'hca0ffe8;
      46983: inst = 32'h24822800;
      46984: inst = 32'h10a00000;
      46985: inst = 32'hca00004;
      46986: inst = 32'h38632800;
      46987: inst = 32'h38842800;
      46988: inst = 32'h10a00000;
      46989: inst = 32'hca0b791;
      46990: inst = 32'h13e00001;
      46991: inst = 32'hfe0d96a;
      46992: inst = 32'h5be00000;
      46993: inst = 32'h8c50000;
      46994: inst = 32'h24612800;
      46995: inst = 32'h10a0ffff;
      46996: inst = 32'hca0ffe8;
      46997: inst = 32'h24822800;
      46998: inst = 32'h10a00000;
      46999: inst = 32'hca00004;
      47000: inst = 32'h38632800;
      47001: inst = 32'h38842800;
      47002: inst = 32'h10a00000;
      47003: inst = 32'hca0b79f;
      47004: inst = 32'h13e00001;
      47005: inst = 32'hfe0d96a;
      47006: inst = 32'h5be00000;
      47007: inst = 32'h8c50000;
      47008: inst = 32'h24612800;
      47009: inst = 32'h10a0ffff;
      47010: inst = 32'hca0ffe8;
      47011: inst = 32'h24822800;
      47012: inst = 32'h10a00000;
      47013: inst = 32'hca00004;
      47014: inst = 32'h38632800;
      47015: inst = 32'h38842800;
      47016: inst = 32'h10a00000;
      47017: inst = 32'hca0b7ad;
      47018: inst = 32'h13e00001;
      47019: inst = 32'hfe0d96a;
      47020: inst = 32'h5be00000;
      47021: inst = 32'h8c50000;
      47022: inst = 32'h24612800;
      47023: inst = 32'h10a0ffff;
      47024: inst = 32'hca0ffe8;
      47025: inst = 32'h24822800;
      47026: inst = 32'h10a00000;
      47027: inst = 32'hca00004;
      47028: inst = 32'h38632800;
      47029: inst = 32'h38842800;
      47030: inst = 32'h10a00000;
      47031: inst = 32'hca0b7bb;
      47032: inst = 32'h13e00001;
      47033: inst = 32'hfe0d96a;
      47034: inst = 32'h5be00000;
      47035: inst = 32'h8c50000;
      47036: inst = 32'h24612800;
      47037: inst = 32'h10a0ffff;
      47038: inst = 32'hca0ffe8;
      47039: inst = 32'h24822800;
      47040: inst = 32'h10a00000;
      47041: inst = 32'hca00004;
      47042: inst = 32'h38632800;
      47043: inst = 32'h38842800;
      47044: inst = 32'h10a00000;
      47045: inst = 32'hca0b7c9;
      47046: inst = 32'h13e00001;
      47047: inst = 32'hfe0d96a;
      47048: inst = 32'h5be00000;
      47049: inst = 32'h8c50000;
      47050: inst = 32'h24612800;
      47051: inst = 32'h10a0ffff;
      47052: inst = 32'hca0ffe8;
      47053: inst = 32'h24822800;
      47054: inst = 32'h10a00000;
      47055: inst = 32'hca00004;
      47056: inst = 32'h38632800;
      47057: inst = 32'h38842800;
      47058: inst = 32'h10a00000;
      47059: inst = 32'hca0b7d7;
      47060: inst = 32'h13e00001;
      47061: inst = 32'hfe0d96a;
      47062: inst = 32'h5be00000;
      47063: inst = 32'h8c50000;
      47064: inst = 32'h24612800;
      47065: inst = 32'h10a0ffff;
      47066: inst = 32'hca0ffe8;
      47067: inst = 32'h24822800;
      47068: inst = 32'h10a00000;
      47069: inst = 32'hca00004;
      47070: inst = 32'h38632800;
      47071: inst = 32'h38842800;
      47072: inst = 32'h10a00000;
      47073: inst = 32'hca0b7e5;
      47074: inst = 32'h13e00001;
      47075: inst = 32'hfe0d96a;
      47076: inst = 32'h5be00000;
      47077: inst = 32'h8c50000;
      47078: inst = 32'h24612800;
      47079: inst = 32'h10a0ffff;
      47080: inst = 32'hca0ffe8;
      47081: inst = 32'h24822800;
      47082: inst = 32'h10a00000;
      47083: inst = 32'hca00004;
      47084: inst = 32'h38632800;
      47085: inst = 32'h38842800;
      47086: inst = 32'h10a00000;
      47087: inst = 32'hca0b7f3;
      47088: inst = 32'h13e00001;
      47089: inst = 32'hfe0d96a;
      47090: inst = 32'h5be00000;
      47091: inst = 32'h8c50000;
      47092: inst = 32'h24612800;
      47093: inst = 32'h10a0ffff;
      47094: inst = 32'hca0ffe8;
      47095: inst = 32'h24822800;
      47096: inst = 32'h10a00000;
      47097: inst = 32'hca00004;
      47098: inst = 32'h38632800;
      47099: inst = 32'h38842800;
      47100: inst = 32'h10a00000;
      47101: inst = 32'hca0b801;
      47102: inst = 32'h13e00001;
      47103: inst = 32'hfe0d96a;
      47104: inst = 32'h5be00000;
      47105: inst = 32'h8c50000;
      47106: inst = 32'h24612800;
      47107: inst = 32'h10a0ffff;
      47108: inst = 32'hca0ffe8;
      47109: inst = 32'h24822800;
      47110: inst = 32'h10a00000;
      47111: inst = 32'hca00004;
      47112: inst = 32'h38632800;
      47113: inst = 32'h38842800;
      47114: inst = 32'h10a00000;
      47115: inst = 32'hca0b80f;
      47116: inst = 32'h13e00001;
      47117: inst = 32'hfe0d96a;
      47118: inst = 32'h5be00000;
      47119: inst = 32'h8c50000;
      47120: inst = 32'h24612800;
      47121: inst = 32'h10a0ffff;
      47122: inst = 32'hca0ffe8;
      47123: inst = 32'h24822800;
      47124: inst = 32'h10a00000;
      47125: inst = 32'hca00004;
      47126: inst = 32'h38632800;
      47127: inst = 32'h38842800;
      47128: inst = 32'h10a00000;
      47129: inst = 32'hca0b81d;
      47130: inst = 32'h13e00001;
      47131: inst = 32'hfe0d96a;
      47132: inst = 32'h5be00000;
      47133: inst = 32'h8c50000;
      47134: inst = 32'h24612800;
      47135: inst = 32'h10a0ffff;
      47136: inst = 32'hca0ffe8;
      47137: inst = 32'h24822800;
      47138: inst = 32'h10a00000;
      47139: inst = 32'hca00004;
      47140: inst = 32'h38632800;
      47141: inst = 32'h38842800;
      47142: inst = 32'h10a00000;
      47143: inst = 32'hca0b82b;
      47144: inst = 32'h13e00001;
      47145: inst = 32'hfe0d96a;
      47146: inst = 32'h5be00000;
      47147: inst = 32'h8c50000;
      47148: inst = 32'h24612800;
      47149: inst = 32'h10a0ffff;
      47150: inst = 32'hca0ffe8;
      47151: inst = 32'h24822800;
      47152: inst = 32'h10a00000;
      47153: inst = 32'hca00004;
      47154: inst = 32'h38632800;
      47155: inst = 32'h38842800;
      47156: inst = 32'h10a00000;
      47157: inst = 32'hca0b839;
      47158: inst = 32'h13e00001;
      47159: inst = 32'hfe0d96a;
      47160: inst = 32'h5be00000;
      47161: inst = 32'h8c50000;
      47162: inst = 32'h24612800;
      47163: inst = 32'h10a0ffff;
      47164: inst = 32'hca0ffe8;
      47165: inst = 32'h24822800;
      47166: inst = 32'h10a00000;
      47167: inst = 32'hca00004;
      47168: inst = 32'h38632800;
      47169: inst = 32'h38842800;
      47170: inst = 32'h10a00000;
      47171: inst = 32'hca0b847;
      47172: inst = 32'h13e00001;
      47173: inst = 32'hfe0d96a;
      47174: inst = 32'h5be00000;
      47175: inst = 32'h8c50000;
      47176: inst = 32'h24612800;
      47177: inst = 32'h10a0ffff;
      47178: inst = 32'hca0ffe8;
      47179: inst = 32'h24822800;
      47180: inst = 32'h10a00000;
      47181: inst = 32'hca00004;
      47182: inst = 32'h38632800;
      47183: inst = 32'h38842800;
      47184: inst = 32'h10a00000;
      47185: inst = 32'hca0b855;
      47186: inst = 32'h13e00001;
      47187: inst = 32'hfe0d96a;
      47188: inst = 32'h5be00000;
      47189: inst = 32'h8c50000;
      47190: inst = 32'h24612800;
      47191: inst = 32'h10a0ffff;
      47192: inst = 32'hca0ffe8;
      47193: inst = 32'h24822800;
      47194: inst = 32'h10a00000;
      47195: inst = 32'hca00004;
      47196: inst = 32'h38632800;
      47197: inst = 32'h38842800;
      47198: inst = 32'h10a00000;
      47199: inst = 32'hca0b863;
      47200: inst = 32'h13e00001;
      47201: inst = 32'hfe0d96a;
      47202: inst = 32'h5be00000;
      47203: inst = 32'h8c50000;
      47204: inst = 32'h24612800;
      47205: inst = 32'h10a0ffff;
      47206: inst = 32'hca0ffe8;
      47207: inst = 32'h24822800;
      47208: inst = 32'h10a00000;
      47209: inst = 32'hca00004;
      47210: inst = 32'h38632800;
      47211: inst = 32'h38842800;
      47212: inst = 32'h10a00000;
      47213: inst = 32'hca0b871;
      47214: inst = 32'h13e00001;
      47215: inst = 32'hfe0d96a;
      47216: inst = 32'h5be00000;
      47217: inst = 32'h8c50000;
      47218: inst = 32'h24612800;
      47219: inst = 32'h10a0ffff;
      47220: inst = 32'hca0ffe8;
      47221: inst = 32'h24822800;
      47222: inst = 32'h10a00000;
      47223: inst = 32'hca00004;
      47224: inst = 32'h38632800;
      47225: inst = 32'h38842800;
      47226: inst = 32'h10a00000;
      47227: inst = 32'hca0b87f;
      47228: inst = 32'h13e00001;
      47229: inst = 32'hfe0d96a;
      47230: inst = 32'h5be00000;
      47231: inst = 32'h8c50000;
      47232: inst = 32'h24612800;
      47233: inst = 32'h10a0ffff;
      47234: inst = 32'hca0ffe8;
      47235: inst = 32'h24822800;
      47236: inst = 32'h10a00000;
      47237: inst = 32'hca00004;
      47238: inst = 32'h38632800;
      47239: inst = 32'h38842800;
      47240: inst = 32'h10a00000;
      47241: inst = 32'hca0b88d;
      47242: inst = 32'h13e00001;
      47243: inst = 32'hfe0d96a;
      47244: inst = 32'h5be00000;
      47245: inst = 32'h8c50000;
      47246: inst = 32'h24612800;
      47247: inst = 32'h10a0ffff;
      47248: inst = 32'hca0ffe8;
      47249: inst = 32'h24822800;
      47250: inst = 32'h10a00000;
      47251: inst = 32'hca00004;
      47252: inst = 32'h38632800;
      47253: inst = 32'h38842800;
      47254: inst = 32'h10a00000;
      47255: inst = 32'hca0b89b;
      47256: inst = 32'h13e00001;
      47257: inst = 32'hfe0d96a;
      47258: inst = 32'h5be00000;
      47259: inst = 32'h8c50000;
      47260: inst = 32'h24612800;
      47261: inst = 32'h10a0ffff;
      47262: inst = 32'hca0ffe8;
      47263: inst = 32'h24822800;
      47264: inst = 32'h10a00000;
      47265: inst = 32'hca00004;
      47266: inst = 32'h38632800;
      47267: inst = 32'h38842800;
      47268: inst = 32'h10a00000;
      47269: inst = 32'hca0b8a9;
      47270: inst = 32'h13e00001;
      47271: inst = 32'hfe0d96a;
      47272: inst = 32'h5be00000;
      47273: inst = 32'h8c50000;
      47274: inst = 32'h24612800;
      47275: inst = 32'h10a0ffff;
      47276: inst = 32'hca0ffe9;
      47277: inst = 32'h24822800;
      47278: inst = 32'h10a00000;
      47279: inst = 32'hca00004;
      47280: inst = 32'h38632800;
      47281: inst = 32'h38842800;
      47282: inst = 32'h10a00000;
      47283: inst = 32'hca0b8b7;
      47284: inst = 32'h13e00001;
      47285: inst = 32'hfe0d96a;
      47286: inst = 32'h5be00000;
      47287: inst = 32'h8c50000;
      47288: inst = 32'h24612800;
      47289: inst = 32'h10a0ffff;
      47290: inst = 32'hca0ffe9;
      47291: inst = 32'h24822800;
      47292: inst = 32'h10a00000;
      47293: inst = 32'hca00004;
      47294: inst = 32'h38632800;
      47295: inst = 32'h38842800;
      47296: inst = 32'h10a00000;
      47297: inst = 32'hca0b8c5;
      47298: inst = 32'h13e00001;
      47299: inst = 32'hfe0d96a;
      47300: inst = 32'h5be00000;
      47301: inst = 32'h8c50000;
      47302: inst = 32'h24612800;
      47303: inst = 32'h10a0ffff;
      47304: inst = 32'hca0ffe9;
      47305: inst = 32'h24822800;
      47306: inst = 32'h10a00000;
      47307: inst = 32'hca00004;
      47308: inst = 32'h38632800;
      47309: inst = 32'h38842800;
      47310: inst = 32'h10a00000;
      47311: inst = 32'hca0b8d3;
      47312: inst = 32'h13e00001;
      47313: inst = 32'hfe0d96a;
      47314: inst = 32'h5be00000;
      47315: inst = 32'h8c50000;
      47316: inst = 32'h24612800;
      47317: inst = 32'h10a0ffff;
      47318: inst = 32'hca0ffe9;
      47319: inst = 32'h24822800;
      47320: inst = 32'h10a00000;
      47321: inst = 32'hca00004;
      47322: inst = 32'h38632800;
      47323: inst = 32'h38842800;
      47324: inst = 32'h10a00000;
      47325: inst = 32'hca0b8e1;
      47326: inst = 32'h13e00001;
      47327: inst = 32'hfe0d96a;
      47328: inst = 32'h5be00000;
      47329: inst = 32'h8c50000;
      47330: inst = 32'h24612800;
      47331: inst = 32'h10a0ffff;
      47332: inst = 32'hca0ffe9;
      47333: inst = 32'h24822800;
      47334: inst = 32'h10a00000;
      47335: inst = 32'hca00004;
      47336: inst = 32'h38632800;
      47337: inst = 32'h38842800;
      47338: inst = 32'h10a00000;
      47339: inst = 32'hca0b8ef;
      47340: inst = 32'h13e00001;
      47341: inst = 32'hfe0d96a;
      47342: inst = 32'h5be00000;
      47343: inst = 32'h8c50000;
      47344: inst = 32'h24612800;
      47345: inst = 32'h10a0ffff;
      47346: inst = 32'hca0ffe9;
      47347: inst = 32'h24822800;
      47348: inst = 32'h10a00000;
      47349: inst = 32'hca00004;
      47350: inst = 32'h38632800;
      47351: inst = 32'h38842800;
      47352: inst = 32'h10a00000;
      47353: inst = 32'hca0b8fd;
      47354: inst = 32'h13e00001;
      47355: inst = 32'hfe0d96a;
      47356: inst = 32'h5be00000;
      47357: inst = 32'h8c50000;
      47358: inst = 32'h24612800;
      47359: inst = 32'h10a0ffff;
      47360: inst = 32'hca0ffe9;
      47361: inst = 32'h24822800;
      47362: inst = 32'h10a00000;
      47363: inst = 32'hca00004;
      47364: inst = 32'h38632800;
      47365: inst = 32'h38842800;
      47366: inst = 32'h10a00000;
      47367: inst = 32'hca0b90b;
      47368: inst = 32'h13e00001;
      47369: inst = 32'hfe0d96a;
      47370: inst = 32'h5be00000;
      47371: inst = 32'h8c50000;
      47372: inst = 32'h24612800;
      47373: inst = 32'h10a0ffff;
      47374: inst = 32'hca0ffe9;
      47375: inst = 32'h24822800;
      47376: inst = 32'h10a00000;
      47377: inst = 32'hca00004;
      47378: inst = 32'h38632800;
      47379: inst = 32'h38842800;
      47380: inst = 32'h10a00000;
      47381: inst = 32'hca0b919;
      47382: inst = 32'h13e00001;
      47383: inst = 32'hfe0d96a;
      47384: inst = 32'h5be00000;
      47385: inst = 32'h8c50000;
      47386: inst = 32'h24612800;
      47387: inst = 32'h10a0ffff;
      47388: inst = 32'hca0ffe9;
      47389: inst = 32'h24822800;
      47390: inst = 32'h10a00000;
      47391: inst = 32'hca00004;
      47392: inst = 32'h38632800;
      47393: inst = 32'h38842800;
      47394: inst = 32'h10a00000;
      47395: inst = 32'hca0b927;
      47396: inst = 32'h13e00001;
      47397: inst = 32'hfe0d96a;
      47398: inst = 32'h5be00000;
      47399: inst = 32'h8c50000;
      47400: inst = 32'h24612800;
      47401: inst = 32'h10a0ffff;
      47402: inst = 32'hca0ffe9;
      47403: inst = 32'h24822800;
      47404: inst = 32'h10a00000;
      47405: inst = 32'hca00004;
      47406: inst = 32'h38632800;
      47407: inst = 32'h38842800;
      47408: inst = 32'h10a00000;
      47409: inst = 32'hca0b935;
      47410: inst = 32'h13e00001;
      47411: inst = 32'hfe0d96a;
      47412: inst = 32'h5be00000;
      47413: inst = 32'h8c50000;
      47414: inst = 32'h24612800;
      47415: inst = 32'h10a0ffff;
      47416: inst = 32'hca0ffe9;
      47417: inst = 32'h24822800;
      47418: inst = 32'h10a00000;
      47419: inst = 32'hca00004;
      47420: inst = 32'h38632800;
      47421: inst = 32'h38842800;
      47422: inst = 32'h10a00000;
      47423: inst = 32'hca0b943;
      47424: inst = 32'h13e00001;
      47425: inst = 32'hfe0d96a;
      47426: inst = 32'h5be00000;
      47427: inst = 32'h8c50000;
      47428: inst = 32'h24612800;
      47429: inst = 32'h10a0ffff;
      47430: inst = 32'hca0ffe9;
      47431: inst = 32'h24822800;
      47432: inst = 32'h10a00000;
      47433: inst = 32'hca00004;
      47434: inst = 32'h38632800;
      47435: inst = 32'h38842800;
      47436: inst = 32'h10a00000;
      47437: inst = 32'hca0b951;
      47438: inst = 32'h13e00001;
      47439: inst = 32'hfe0d96a;
      47440: inst = 32'h5be00000;
      47441: inst = 32'h8c50000;
      47442: inst = 32'h24612800;
      47443: inst = 32'h10a0ffff;
      47444: inst = 32'hca0ffe9;
      47445: inst = 32'h24822800;
      47446: inst = 32'h10a00000;
      47447: inst = 32'hca00004;
      47448: inst = 32'h38632800;
      47449: inst = 32'h38842800;
      47450: inst = 32'h10a00000;
      47451: inst = 32'hca0b95f;
      47452: inst = 32'h13e00001;
      47453: inst = 32'hfe0d96a;
      47454: inst = 32'h5be00000;
      47455: inst = 32'h8c50000;
      47456: inst = 32'h24612800;
      47457: inst = 32'h10a0ffff;
      47458: inst = 32'hca0ffe9;
      47459: inst = 32'h24822800;
      47460: inst = 32'h10a00000;
      47461: inst = 32'hca00004;
      47462: inst = 32'h38632800;
      47463: inst = 32'h38842800;
      47464: inst = 32'h10a00000;
      47465: inst = 32'hca0b96d;
      47466: inst = 32'h13e00001;
      47467: inst = 32'hfe0d96a;
      47468: inst = 32'h5be00000;
      47469: inst = 32'h8c50000;
      47470: inst = 32'h24612800;
      47471: inst = 32'h10a0ffff;
      47472: inst = 32'hca0ffe9;
      47473: inst = 32'h24822800;
      47474: inst = 32'h10a00000;
      47475: inst = 32'hca00004;
      47476: inst = 32'h38632800;
      47477: inst = 32'h38842800;
      47478: inst = 32'h10a00000;
      47479: inst = 32'hca0b97b;
      47480: inst = 32'h13e00001;
      47481: inst = 32'hfe0d96a;
      47482: inst = 32'h5be00000;
      47483: inst = 32'h8c50000;
      47484: inst = 32'h24612800;
      47485: inst = 32'h10a0ffff;
      47486: inst = 32'hca0ffe9;
      47487: inst = 32'h24822800;
      47488: inst = 32'h10a00000;
      47489: inst = 32'hca00004;
      47490: inst = 32'h38632800;
      47491: inst = 32'h38842800;
      47492: inst = 32'h10a00000;
      47493: inst = 32'hca0b989;
      47494: inst = 32'h13e00001;
      47495: inst = 32'hfe0d96a;
      47496: inst = 32'h5be00000;
      47497: inst = 32'h8c50000;
      47498: inst = 32'h24612800;
      47499: inst = 32'h10a0ffff;
      47500: inst = 32'hca0ffe9;
      47501: inst = 32'h24822800;
      47502: inst = 32'h10a00000;
      47503: inst = 32'hca00004;
      47504: inst = 32'h38632800;
      47505: inst = 32'h38842800;
      47506: inst = 32'h10a00000;
      47507: inst = 32'hca0b997;
      47508: inst = 32'h13e00001;
      47509: inst = 32'hfe0d96a;
      47510: inst = 32'h5be00000;
      47511: inst = 32'h8c50000;
      47512: inst = 32'h24612800;
      47513: inst = 32'h10a0ffff;
      47514: inst = 32'hca0ffe9;
      47515: inst = 32'h24822800;
      47516: inst = 32'h10a00000;
      47517: inst = 32'hca00004;
      47518: inst = 32'h38632800;
      47519: inst = 32'h38842800;
      47520: inst = 32'h10a00000;
      47521: inst = 32'hca0b9a5;
      47522: inst = 32'h13e00001;
      47523: inst = 32'hfe0d96a;
      47524: inst = 32'h5be00000;
      47525: inst = 32'h8c50000;
      47526: inst = 32'h24612800;
      47527: inst = 32'h10a0ffff;
      47528: inst = 32'hca0ffe9;
      47529: inst = 32'h24822800;
      47530: inst = 32'h10a00000;
      47531: inst = 32'hca00004;
      47532: inst = 32'h38632800;
      47533: inst = 32'h38842800;
      47534: inst = 32'h10a00000;
      47535: inst = 32'hca0b9b3;
      47536: inst = 32'h13e00001;
      47537: inst = 32'hfe0d96a;
      47538: inst = 32'h5be00000;
      47539: inst = 32'h8c50000;
      47540: inst = 32'h24612800;
      47541: inst = 32'h10a0ffff;
      47542: inst = 32'hca0ffe9;
      47543: inst = 32'h24822800;
      47544: inst = 32'h10a00000;
      47545: inst = 32'hca00004;
      47546: inst = 32'h38632800;
      47547: inst = 32'h38842800;
      47548: inst = 32'h10a00000;
      47549: inst = 32'hca0b9c1;
      47550: inst = 32'h13e00001;
      47551: inst = 32'hfe0d96a;
      47552: inst = 32'h5be00000;
      47553: inst = 32'h8c50000;
      47554: inst = 32'h24612800;
      47555: inst = 32'h10a0ffff;
      47556: inst = 32'hca0ffe9;
      47557: inst = 32'h24822800;
      47558: inst = 32'h10a00000;
      47559: inst = 32'hca00004;
      47560: inst = 32'h38632800;
      47561: inst = 32'h38842800;
      47562: inst = 32'h10a00000;
      47563: inst = 32'hca0b9cf;
      47564: inst = 32'h13e00001;
      47565: inst = 32'hfe0d96a;
      47566: inst = 32'h5be00000;
      47567: inst = 32'h8c50000;
      47568: inst = 32'h24612800;
      47569: inst = 32'h10a0ffff;
      47570: inst = 32'hca0ffe9;
      47571: inst = 32'h24822800;
      47572: inst = 32'h10a00000;
      47573: inst = 32'hca00004;
      47574: inst = 32'h38632800;
      47575: inst = 32'h38842800;
      47576: inst = 32'h10a00000;
      47577: inst = 32'hca0b9dd;
      47578: inst = 32'h13e00001;
      47579: inst = 32'hfe0d96a;
      47580: inst = 32'h5be00000;
      47581: inst = 32'h8c50000;
      47582: inst = 32'h24612800;
      47583: inst = 32'h10a0ffff;
      47584: inst = 32'hca0ffe9;
      47585: inst = 32'h24822800;
      47586: inst = 32'h10a00000;
      47587: inst = 32'hca00004;
      47588: inst = 32'h38632800;
      47589: inst = 32'h38842800;
      47590: inst = 32'h10a00000;
      47591: inst = 32'hca0b9eb;
      47592: inst = 32'h13e00001;
      47593: inst = 32'hfe0d96a;
      47594: inst = 32'h5be00000;
      47595: inst = 32'h8c50000;
      47596: inst = 32'h24612800;
      47597: inst = 32'h10a0ffff;
      47598: inst = 32'hca0ffe9;
      47599: inst = 32'h24822800;
      47600: inst = 32'h10a00000;
      47601: inst = 32'hca00004;
      47602: inst = 32'h38632800;
      47603: inst = 32'h38842800;
      47604: inst = 32'h10a00000;
      47605: inst = 32'hca0b9f9;
      47606: inst = 32'h13e00001;
      47607: inst = 32'hfe0d96a;
      47608: inst = 32'h5be00000;
      47609: inst = 32'h8c50000;
      47610: inst = 32'h24612800;
      47611: inst = 32'h10a0ffff;
      47612: inst = 32'hca0ffe9;
      47613: inst = 32'h24822800;
      47614: inst = 32'h10a00000;
      47615: inst = 32'hca00004;
      47616: inst = 32'h38632800;
      47617: inst = 32'h38842800;
      47618: inst = 32'h10a00000;
      47619: inst = 32'hca0ba07;
      47620: inst = 32'h13e00001;
      47621: inst = 32'hfe0d96a;
      47622: inst = 32'h5be00000;
      47623: inst = 32'h8c50000;
      47624: inst = 32'h24612800;
      47625: inst = 32'h10a0ffff;
      47626: inst = 32'hca0ffe9;
      47627: inst = 32'h24822800;
      47628: inst = 32'h10a00000;
      47629: inst = 32'hca00004;
      47630: inst = 32'h38632800;
      47631: inst = 32'h38842800;
      47632: inst = 32'h10a00000;
      47633: inst = 32'hca0ba15;
      47634: inst = 32'h13e00001;
      47635: inst = 32'hfe0d96a;
      47636: inst = 32'h5be00000;
      47637: inst = 32'h8c50000;
      47638: inst = 32'h24612800;
      47639: inst = 32'h10a0ffff;
      47640: inst = 32'hca0ffe9;
      47641: inst = 32'h24822800;
      47642: inst = 32'h10a00000;
      47643: inst = 32'hca00004;
      47644: inst = 32'h38632800;
      47645: inst = 32'h38842800;
      47646: inst = 32'h10a00000;
      47647: inst = 32'hca0ba23;
      47648: inst = 32'h13e00001;
      47649: inst = 32'hfe0d96a;
      47650: inst = 32'h5be00000;
      47651: inst = 32'h8c50000;
      47652: inst = 32'h24612800;
      47653: inst = 32'h10a0ffff;
      47654: inst = 32'hca0ffe9;
      47655: inst = 32'h24822800;
      47656: inst = 32'h10a00000;
      47657: inst = 32'hca00004;
      47658: inst = 32'h38632800;
      47659: inst = 32'h38842800;
      47660: inst = 32'h10a00000;
      47661: inst = 32'hca0ba31;
      47662: inst = 32'h13e00001;
      47663: inst = 32'hfe0d96a;
      47664: inst = 32'h5be00000;
      47665: inst = 32'h8c50000;
      47666: inst = 32'h24612800;
      47667: inst = 32'h10a0ffff;
      47668: inst = 32'hca0ffe9;
      47669: inst = 32'h24822800;
      47670: inst = 32'h10a00000;
      47671: inst = 32'hca00004;
      47672: inst = 32'h38632800;
      47673: inst = 32'h38842800;
      47674: inst = 32'h10a00000;
      47675: inst = 32'hca0ba3f;
      47676: inst = 32'h13e00001;
      47677: inst = 32'hfe0d96a;
      47678: inst = 32'h5be00000;
      47679: inst = 32'h8c50000;
      47680: inst = 32'h24612800;
      47681: inst = 32'h10a0ffff;
      47682: inst = 32'hca0ffe9;
      47683: inst = 32'h24822800;
      47684: inst = 32'h10a00000;
      47685: inst = 32'hca00004;
      47686: inst = 32'h38632800;
      47687: inst = 32'h38842800;
      47688: inst = 32'h10a00000;
      47689: inst = 32'hca0ba4d;
      47690: inst = 32'h13e00001;
      47691: inst = 32'hfe0d96a;
      47692: inst = 32'h5be00000;
      47693: inst = 32'h8c50000;
      47694: inst = 32'h24612800;
      47695: inst = 32'h10a0ffff;
      47696: inst = 32'hca0ffe9;
      47697: inst = 32'h24822800;
      47698: inst = 32'h10a00000;
      47699: inst = 32'hca00004;
      47700: inst = 32'h38632800;
      47701: inst = 32'h38842800;
      47702: inst = 32'h10a00000;
      47703: inst = 32'hca0ba5b;
      47704: inst = 32'h13e00001;
      47705: inst = 32'hfe0d96a;
      47706: inst = 32'h5be00000;
      47707: inst = 32'h8c50000;
      47708: inst = 32'h24612800;
      47709: inst = 32'h10a0ffff;
      47710: inst = 32'hca0ffe9;
      47711: inst = 32'h24822800;
      47712: inst = 32'h10a00000;
      47713: inst = 32'hca00004;
      47714: inst = 32'h38632800;
      47715: inst = 32'h38842800;
      47716: inst = 32'h10a00000;
      47717: inst = 32'hca0ba69;
      47718: inst = 32'h13e00001;
      47719: inst = 32'hfe0d96a;
      47720: inst = 32'h5be00000;
      47721: inst = 32'h8c50000;
      47722: inst = 32'h24612800;
      47723: inst = 32'h10a0ffff;
      47724: inst = 32'hca0ffe9;
      47725: inst = 32'h24822800;
      47726: inst = 32'h10a00000;
      47727: inst = 32'hca00004;
      47728: inst = 32'h38632800;
      47729: inst = 32'h38842800;
      47730: inst = 32'h10a00000;
      47731: inst = 32'hca0ba77;
      47732: inst = 32'h13e00001;
      47733: inst = 32'hfe0d96a;
      47734: inst = 32'h5be00000;
      47735: inst = 32'h8c50000;
      47736: inst = 32'h24612800;
      47737: inst = 32'h10a0ffff;
      47738: inst = 32'hca0ffe9;
      47739: inst = 32'h24822800;
      47740: inst = 32'h10a00000;
      47741: inst = 32'hca00004;
      47742: inst = 32'h38632800;
      47743: inst = 32'h38842800;
      47744: inst = 32'h10a00000;
      47745: inst = 32'hca0ba85;
      47746: inst = 32'h13e00001;
      47747: inst = 32'hfe0d96a;
      47748: inst = 32'h5be00000;
      47749: inst = 32'h8c50000;
      47750: inst = 32'h24612800;
      47751: inst = 32'h10a0ffff;
      47752: inst = 32'hca0ffe9;
      47753: inst = 32'h24822800;
      47754: inst = 32'h10a00000;
      47755: inst = 32'hca00004;
      47756: inst = 32'h38632800;
      47757: inst = 32'h38842800;
      47758: inst = 32'h10a00000;
      47759: inst = 32'hca0ba93;
      47760: inst = 32'h13e00001;
      47761: inst = 32'hfe0d96a;
      47762: inst = 32'h5be00000;
      47763: inst = 32'h8c50000;
      47764: inst = 32'h24612800;
      47765: inst = 32'h10a0ffff;
      47766: inst = 32'hca0ffe9;
      47767: inst = 32'h24822800;
      47768: inst = 32'h10a00000;
      47769: inst = 32'hca00004;
      47770: inst = 32'h38632800;
      47771: inst = 32'h38842800;
      47772: inst = 32'h10a00000;
      47773: inst = 32'hca0baa1;
      47774: inst = 32'h13e00001;
      47775: inst = 32'hfe0d96a;
      47776: inst = 32'h5be00000;
      47777: inst = 32'h8c50000;
      47778: inst = 32'h24612800;
      47779: inst = 32'h10a0ffff;
      47780: inst = 32'hca0ffe9;
      47781: inst = 32'h24822800;
      47782: inst = 32'h10a00000;
      47783: inst = 32'hca00004;
      47784: inst = 32'h38632800;
      47785: inst = 32'h38842800;
      47786: inst = 32'h10a00000;
      47787: inst = 32'hca0baaf;
      47788: inst = 32'h13e00001;
      47789: inst = 32'hfe0d96a;
      47790: inst = 32'h5be00000;
      47791: inst = 32'h8c50000;
      47792: inst = 32'h24612800;
      47793: inst = 32'h10a0ffff;
      47794: inst = 32'hca0ffe9;
      47795: inst = 32'h24822800;
      47796: inst = 32'h10a00000;
      47797: inst = 32'hca00004;
      47798: inst = 32'h38632800;
      47799: inst = 32'h38842800;
      47800: inst = 32'h10a00000;
      47801: inst = 32'hca0babd;
      47802: inst = 32'h13e00001;
      47803: inst = 32'hfe0d96a;
      47804: inst = 32'h5be00000;
      47805: inst = 32'h8c50000;
      47806: inst = 32'h24612800;
      47807: inst = 32'h10a0ffff;
      47808: inst = 32'hca0ffe9;
      47809: inst = 32'h24822800;
      47810: inst = 32'h10a00000;
      47811: inst = 32'hca00004;
      47812: inst = 32'h38632800;
      47813: inst = 32'h38842800;
      47814: inst = 32'h10a00000;
      47815: inst = 32'hca0bacb;
      47816: inst = 32'h13e00001;
      47817: inst = 32'hfe0d96a;
      47818: inst = 32'h5be00000;
      47819: inst = 32'h8c50000;
      47820: inst = 32'h24612800;
      47821: inst = 32'h10a0ffff;
      47822: inst = 32'hca0ffe9;
      47823: inst = 32'h24822800;
      47824: inst = 32'h10a00000;
      47825: inst = 32'hca00004;
      47826: inst = 32'h38632800;
      47827: inst = 32'h38842800;
      47828: inst = 32'h10a00000;
      47829: inst = 32'hca0bad9;
      47830: inst = 32'h13e00001;
      47831: inst = 32'hfe0d96a;
      47832: inst = 32'h5be00000;
      47833: inst = 32'h8c50000;
      47834: inst = 32'h24612800;
      47835: inst = 32'h10a0ffff;
      47836: inst = 32'hca0ffe9;
      47837: inst = 32'h24822800;
      47838: inst = 32'h10a00000;
      47839: inst = 32'hca00004;
      47840: inst = 32'h38632800;
      47841: inst = 32'h38842800;
      47842: inst = 32'h10a00000;
      47843: inst = 32'hca0bae7;
      47844: inst = 32'h13e00001;
      47845: inst = 32'hfe0d96a;
      47846: inst = 32'h5be00000;
      47847: inst = 32'h8c50000;
      47848: inst = 32'h24612800;
      47849: inst = 32'h10a0ffff;
      47850: inst = 32'hca0ffe9;
      47851: inst = 32'h24822800;
      47852: inst = 32'h10a00000;
      47853: inst = 32'hca00004;
      47854: inst = 32'h38632800;
      47855: inst = 32'h38842800;
      47856: inst = 32'h10a00000;
      47857: inst = 32'hca0baf5;
      47858: inst = 32'h13e00001;
      47859: inst = 32'hfe0d96a;
      47860: inst = 32'h5be00000;
      47861: inst = 32'h8c50000;
      47862: inst = 32'h24612800;
      47863: inst = 32'h10a0ffff;
      47864: inst = 32'hca0ffe9;
      47865: inst = 32'h24822800;
      47866: inst = 32'h10a00000;
      47867: inst = 32'hca00004;
      47868: inst = 32'h38632800;
      47869: inst = 32'h38842800;
      47870: inst = 32'h10a00000;
      47871: inst = 32'hca0bb03;
      47872: inst = 32'h13e00001;
      47873: inst = 32'hfe0d96a;
      47874: inst = 32'h5be00000;
      47875: inst = 32'h8c50000;
      47876: inst = 32'h24612800;
      47877: inst = 32'h10a0ffff;
      47878: inst = 32'hca0ffe9;
      47879: inst = 32'h24822800;
      47880: inst = 32'h10a00000;
      47881: inst = 32'hca00004;
      47882: inst = 32'h38632800;
      47883: inst = 32'h38842800;
      47884: inst = 32'h10a00000;
      47885: inst = 32'hca0bb11;
      47886: inst = 32'h13e00001;
      47887: inst = 32'hfe0d96a;
      47888: inst = 32'h5be00000;
      47889: inst = 32'h8c50000;
      47890: inst = 32'h24612800;
      47891: inst = 32'h10a0ffff;
      47892: inst = 32'hca0ffe9;
      47893: inst = 32'h24822800;
      47894: inst = 32'h10a00000;
      47895: inst = 32'hca00004;
      47896: inst = 32'h38632800;
      47897: inst = 32'h38842800;
      47898: inst = 32'h10a00000;
      47899: inst = 32'hca0bb1f;
      47900: inst = 32'h13e00001;
      47901: inst = 32'hfe0d96a;
      47902: inst = 32'h5be00000;
      47903: inst = 32'h8c50000;
      47904: inst = 32'h24612800;
      47905: inst = 32'h10a0ffff;
      47906: inst = 32'hca0ffe9;
      47907: inst = 32'h24822800;
      47908: inst = 32'h10a00000;
      47909: inst = 32'hca00004;
      47910: inst = 32'h38632800;
      47911: inst = 32'h38842800;
      47912: inst = 32'h10a00000;
      47913: inst = 32'hca0bb2d;
      47914: inst = 32'h13e00001;
      47915: inst = 32'hfe0d96a;
      47916: inst = 32'h5be00000;
      47917: inst = 32'h8c50000;
      47918: inst = 32'h24612800;
      47919: inst = 32'h10a0ffff;
      47920: inst = 32'hca0ffe9;
      47921: inst = 32'h24822800;
      47922: inst = 32'h10a00000;
      47923: inst = 32'hca00004;
      47924: inst = 32'h38632800;
      47925: inst = 32'h38842800;
      47926: inst = 32'h10a00000;
      47927: inst = 32'hca0bb3b;
      47928: inst = 32'h13e00001;
      47929: inst = 32'hfe0d96a;
      47930: inst = 32'h5be00000;
      47931: inst = 32'h8c50000;
      47932: inst = 32'h24612800;
      47933: inst = 32'h10a0ffff;
      47934: inst = 32'hca0ffe9;
      47935: inst = 32'h24822800;
      47936: inst = 32'h10a00000;
      47937: inst = 32'hca00004;
      47938: inst = 32'h38632800;
      47939: inst = 32'h38842800;
      47940: inst = 32'h10a00000;
      47941: inst = 32'hca0bb49;
      47942: inst = 32'h13e00001;
      47943: inst = 32'hfe0d96a;
      47944: inst = 32'h5be00000;
      47945: inst = 32'h8c50000;
      47946: inst = 32'h24612800;
      47947: inst = 32'h10a0ffff;
      47948: inst = 32'hca0ffe9;
      47949: inst = 32'h24822800;
      47950: inst = 32'h10a00000;
      47951: inst = 32'hca00004;
      47952: inst = 32'h38632800;
      47953: inst = 32'h38842800;
      47954: inst = 32'h10a00000;
      47955: inst = 32'hca0bb57;
      47956: inst = 32'h13e00001;
      47957: inst = 32'hfe0d96a;
      47958: inst = 32'h5be00000;
      47959: inst = 32'h8c50000;
      47960: inst = 32'h24612800;
      47961: inst = 32'h10a0ffff;
      47962: inst = 32'hca0ffe9;
      47963: inst = 32'h24822800;
      47964: inst = 32'h10a00000;
      47965: inst = 32'hca00004;
      47966: inst = 32'h38632800;
      47967: inst = 32'h38842800;
      47968: inst = 32'h10a00000;
      47969: inst = 32'hca0bb65;
      47970: inst = 32'h13e00001;
      47971: inst = 32'hfe0d96a;
      47972: inst = 32'h5be00000;
      47973: inst = 32'h8c50000;
      47974: inst = 32'h24612800;
      47975: inst = 32'h10a0ffff;
      47976: inst = 32'hca0ffe9;
      47977: inst = 32'h24822800;
      47978: inst = 32'h10a00000;
      47979: inst = 32'hca00004;
      47980: inst = 32'h38632800;
      47981: inst = 32'h38842800;
      47982: inst = 32'h10a00000;
      47983: inst = 32'hca0bb73;
      47984: inst = 32'h13e00001;
      47985: inst = 32'hfe0d96a;
      47986: inst = 32'h5be00000;
      47987: inst = 32'h8c50000;
      47988: inst = 32'h24612800;
      47989: inst = 32'h10a0ffff;
      47990: inst = 32'hca0ffe9;
      47991: inst = 32'h24822800;
      47992: inst = 32'h10a00000;
      47993: inst = 32'hca00004;
      47994: inst = 32'h38632800;
      47995: inst = 32'h38842800;
      47996: inst = 32'h10a00000;
      47997: inst = 32'hca0bb81;
      47998: inst = 32'h13e00001;
      47999: inst = 32'hfe0d96a;
      48000: inst = 32'h5be00000;
      48001: inst = 32'h8c50000;
      48002: inst = 32'h24612800;
      48003: inst = 32'h10a0ffff;
      48004: inst = 32'hca0ffe9;
      48005: inst = 32'h24822800;
      48006: inst = 32'h10a00000;
      48007: inst = 32'hca00004;
      48008: inst = 32'h38632800;
      48009: inst = 32'h38842800;
      48010: inst = 32'h10a00000;
      48011: inst = 32'hca0bb8f;
      48012: inst = 32'h13e00001;
      48013: inst = 32'hfe0d96a;
      48014: inst = 32'h5be00000;
      48015: inst = 32'h8c50000;
      48016: inst = 32'h24612800;
      48017: inst = 32'h10a0ffff;
      48018: inst = 32'hca0ffe9;
      48019: inst = 32'h24822800;
      48020: inst = 32'h10a00000;
      48021: inst = 32'hca00004;
      48022: inst = 32'h38632800;
      48023: inst = 32'h38842800;
      48024: inst = 32'h10a00000;
      48025: inst = 32'hca0bb9d;
      48026: inst = 32'h13e00001;
      48027: inst = 32'hfe0d96a;
      48028: inst = 32'h5be00000;
      48029: inst = 32'h8c50000;
      48030: inst = 32'h24612800;
      48031: inst = 32'h10a0ffff;
      48032: inst = 32'hca0ffe9;
      48033: inst = 32'h24822800;
      48034: inst = 32'h10a00000;
      48035: inst = 32'hca00004;
      48036: inst = 32'h38632800;
      48037: inst = 32'h38842800;
      48038: inst = 32'h10a00000;
      48039: inst = 32'hca0bbab;
      48040: inst = 32'h13e00001;
      48041: inst = 32'hfe0d96a;
      48042: inst = 32'h5be00000;
      48043: inst = 32'h8c50000;
      48044: inst = 32'h24612800;
      48045: inst = 32'h10a0ffff;
      48046: inst = 32'hca0ffe9;
      48047: inst = 32'h24822800;
      48048: inst = 32'h10a00000;
      48049: inst = 32'hca00004;
      48050: inst = 32'h38632800;
      48051: inst = 32'h38842800;
      48052: inst = 32'h10a00000;
      48053: inst = 32'hca0bbb9;
      48054: inst = 32'h13e00001;
      48055: inst = 32'hfe0d96a;
      48056: inst = 32'h5be00000;
      48057: inst = 32'h8c50000;
      48058: inst = 32'h24612800;
      48059: inst = 32'h10a0ffff;
      48060: inst = 32'hca0ffe9;
      48061: inst = 32'h24822800;
      48062: inst = 32'h10a00000;
      48063: inst = 32'hca00004;
      48064: inst = 32'h38632800;
      48065: inst = 32'h38842800;
      48066: inst = 32'h10a00000;
      48067: inst = 32'hca0bbc7;
      48068: inst = 32'h13e00001;
      48069: inst = 32'hfe0d96a;
      48070: inst = 32'h5be00000;
      48071: inst = 32'h8c50000;
      48072: inst = 32'h24612800;
      48073: inst = 32'h10a0ffff;
      48074: inst = 32'hca0ffe9;
      48075: inst = 32'h24822800;
      48076: inst = 32'h10a00000;
      48077: inst = 32'hca00004;
      48078: inst = 32'h38632800;
      48079: inst = 32'h38842800;
      48080: inst = 32'h10a00000;
      48081: inst = 32'hca0bbd5;
      48082: inst = 32'h13e00001;
      48083: inst = 32'hfe0d96a;
      48084: inst = 32'h5be00000;
      48085: inst = 32'h8c50000;
      48086: inst = 32'h24612800;
      48087: inst = 32'h10a0ffff;
      48088: inst = 32'hca0ffe9;
      48089: inst = 32'h24822800;
      48090: inst = 32'h10a00000;
      48091: inst = 32'hca00004;
      48092: inst = 32'h38632800;
      48093: inst = 32'h38842800;
      48094: inst = 32'h10a00000;
      48095: inst = 32'hca0bbe3;
      48096: inst = 32'h13e00001;
      48097: inst = 32'hfe0d96a;
      48098: inst = 32'h5be00000;
      48099: inst = 32'h8c50000;
      48100: inst = 32'h24612800;
      48101: inst = 32'h10a0ffff;
      48102: inst = 32'hca0ffe9;
      48103: inst = 32'h24822800;
      48104: inst = 32'h10a00000;
      48105: inst = 32'hca00004;
      48106: inst = 32'h38632800;
      48107: inst = 32'h38842800;
      48108: inst = 32'h10a00000;
      48109: inst = 32'hca0bbf1;
      48110: inst = 32'h13e00001;
      48111: inst = 32'hfe0d96a;
      48112: inst = 32'h5be00000;
      48113: inst = 32'h8c50000;
      48114: inst = 32'h24612800;
      48115: inst = 32'h10a0ffff;
      48116: inst = 32'hca0ffe9;
      48117: inst = 32'h24822800;
      48118: inst = 32'h10a00000;
      48119: inst = 32'hca00004;
      48120: inst = 32'h38632800;
      48121: inst = 32'h38842800;
      48122: inst = 32'h10a00000;
      48123: inst = 32'hca0bbff;
      48124: inst = 32'h13e00001;
      48125: inst = 32'hfe0d96a;
      48126: inst = 32'h5be00000;
      48127: inst = 32'h8c50000;
      48128: inst = 32'h24612800;
      48129: inst = 32'h10a0ffff;
      48130: inst = 32'hca0ffe9;
      48131: inst = 32'h24822800;
      48132: inst = 32'h10a00000;
      48133: inst = 32'hca00004;
      48134: inst = 32'h38632800;
      48135: inst = 32'h38842800;
      48136: inst = 32'h10a00000;
      48137: inst = 32'hca0bc0d;
      48138: inst = 32'h13e00001;
      48139: inst = 32'hfe0d96a;
      48140: inst = 32'h5be00000;
      48141: inst = 32'h8c50000;
      48142: inst = 32'h24612800;
      48143: inst = 32'h10a0ffff;
      48144: inst = 32'hca0ffe9;
      48145: inst = 32'h24822800;
      48146: inst = 32'h10a00000;
      48147: inst = 32'hca00004;
      48148: inst = 32'h38632800;
      48149: inst = 32'h38842800;
      48150: inst = 32'h10a00000;
      48151: inst = 32'hca0bc1b;
      48152: inst = 32'h13e00001;
      48153: inst = 32'hfe0d96a;
      48154: inst = 32'h5be00000;
      48155: inst = 32'h8c50000;
      48156: inst = 32'h24612800;
      48157: inst = 32'h10a0ffff;
      48158: inst = 32'hca0ffe9;
      48159: inst = 32'h24822800;
      48160: inst = 32'h10a00000;
      48161: inst = 32'hca00004;
      48162: inst = 32'h38632800;
      48163: inst = 32'h38842800;
      48164: inst = 32'h10a00000;
      48165: inst = 32'hca0bc29;
      48166: inst = 32'h13e00001;
      48167: inst = 32'hfe0d96a;
      48168: inst = 32'h5be00000;
      48169: inst = 32'h8c50000;
      48170: inst = 32'h24612800;
      48171: inst = 32'h10a0ffff;
      48172: inst = 32'hca0ffe9;
      48173: inst = 32'h24822800;
      48174: inst = 32'h10a00000;
      48175: inst = 32'hca00004;
      48176: inst = 32'h38632800;
      48177: inst = 32'h38842800;
      48178: inst = 32'h10a00000;
      48179: inst = 32'hca0bc37;
      48180: inst = 32'h13e00001;
      48181: inst = 32'hfe0d96a;
      48182: inst = 32'h5be00000;
      48183: inst = 32'h8c50000;
      48184: inst = 32'h24612800;
      48185: inst = 32'h10a0ffff;
      48186: inst = 32'hca0ffe9;
      48187: inst = 32'h24822800;
      48188: inst = 32'h10a00000;
      48189: inst = 32'hca00004;
      48190: inst = 32'h38632800;
      48191: inst = 32'h38842800;
      48192: inst = 32'h10a00000;
      48193: inst = 32'hca0bc45;
      48194: inst = 32'h13e00001;
      48195: inst = 32'hfe0d96a;
      48196: inst = 32'h5be00000;
      48197: inst = 32'h8c50000;
      48198: inst = 32'h24612800;
      48199: inst = 32'h10a0ffff;
      48200: inst = 32'hca0ffe9;
      48201: inst = 32'h24822800;
      48202: inst = 32'h10a00000;
      48203: inst = 32'hca00004;
      48204: inst = 32'h38632800;
      48205: inst = 32'h38842800;
      48206: inst = 32'h10a00000;
      48207: inst = 32'hca0bc53;
      48208: inst = 32'h13e00001;
      48209: inst = 32'hfe0d96a;
      48210: inst = 32'h5be00000;
      48211: inst = 32'h8c50000;
      48212: inst = 32'h24612800;
      48213: inst = 32'h10a0ffff;
      48214: inst = 32'hca0ffe9;
      48215: inst = 32'h24822800;
      48216: inst = 32'h10a00000;
      48217: inst = 32'hca00004;
      48218: inst = 32'h38632800;
      48219: inst = 32'h38842800;
      48220: inst = 32'h10a00000;
      48221: inst = 32'hca0bc61;
      48222: inst = 32'h13e00001;
      48223: inst = 32'hfe0d96a;
      48224: inst = 32'h5be00000;
      48225: inst = 32'h8c50000;
      48226: inst = 32'h24612800;
      48227: inst = 32'h10a0ffff;
      48228: inst = 32'hca0ffe9;
      48229: inst = 32'h24822800;
      48230: inst = 32'h10a00000;
      48231: inst = 32'hca00004;
      48232: inst = 32'h38632800;
      48233: inst = 32'h38842800;
      48234: inst = 32'h10a00000;
      48235: inst = 32'hca0bc6f;
      48236: inst = 32'h13e00001;
      48237: inst = 32'hfe0d96a;
      48238: inst = 32'h5be00000;
      48239: inst = 32'h8c50000;
      48240: inst = 32'h24612800;
      48241: inst = 32'h10a0ffff;
      48242: inst = 32'hca0ffe9;
      48243: inst = 32'h24822800;
      48244: inst = 32'h10a00000;
      48245: inst = 32'hca00004;
      48246: inst = 32'h38632800;
      48247: inst = 32'h38842800;
      48248: inst = 32'h10a00000;
      48249: inst = 32'hca0bc7d;
      48250: inst = 32'h13e00001;
      48251: inst = 32'hfe0d96a;
      48252: inst = 32'h5be00000;
      48253: inst = 32'h8c50000;
      48254: inst = 32'h24612800;
      48255: inst = 32'h10a0ffff;
      48256: inst = 32'hca0ffe9;
      48257: inst = 32'h24822800;
      48258: inst = 32'h10a00000;
      48259: inst = 32'hca00004;
      48260: inst = 32'h38632800;
      48261: inst = 32'h38842800;
      48262: inst = 32'h10a00000;
      48263: inst = 32'hca0bc8b;
      48264: inst = 32'h13e00001;
      48265: inst = 32'hfe0d96a;
      48266: inst = 32'h5be00000;
      48267: inst = 32'h8c50000;
      48268: inst = 32'h24612800;
      48269: inst = 32'h10a0ffff;
      48270: inst = 32'hca0ffe9;
      48271: inst = 32'h24822800;
      48272: inst = 32'h10a00000;
      48273: inst = 32'hca00004;
      48274: inst = 32'h38632800;
      48275: inst = 32'h38842800;
      48276: inst = 32'h10a00000;
      48277: inst = 32'hca0bc99;
      48278: inst = 32'h13e00001;
      48279: inst = 32'hfe0d96a;
      48280: inst = 32'h5be00000;
      48281: inst = 32'h8c50000;
      48282: inst = 32'h24612800;
      48283: inst = 32'h10a0ffff;
      48284: inst = 32'hca0ffe9;
      48285: inst = 32'h24822800;
      48286: inst = 32'h10a00000;
      48287: inst = 32'hca00004;
      48288: inst = 32'h38632800;
      48289: inst = 32'h38842800;
      48290: inst = 32'h10a00000;
      48291: inst = 32'hca0bca7;
      48292: inst = 32'h13e00001;
      48293: inst = 32'hfe0d96a;
      48294: inst = 32'h5be00000;
      48295: inst = 32'h8c50000;
      48296: inst = 32'h24612800;
      48297: inst = 32'h10a0ffff;
      48298: inst = 32'hca0ffe9;
      48299: inst = 32'h24822800;
      48300: inst = 32'h10a00000;
      48301: inst = 32'hca00004;
      48302: inst = 32'h38632800;
      48303: inst = 32'h38842800;
      48304: inst = 32'h10a00000;
      48305: inst = 32'hca0bcb5;
      48306: inst = 32'h13e00001;
      48307: inst = 32'hfe0d96a;
      48308: inst = 32'h5be00000;
      48309: inst = 32'h8c50000;
      48310: inst = 32'h24612800;
      48311: inst = 32'h10a0ffff;
      48312: inst = 32'hca0ffe9;
      48313: inst = 32'h24822800;
      48314: inst = 32'h10a00000;
      48315: inst = 32'hca00004;
      48316: inst = 32'h38632800;
      48317: inst = 32'h38842800;
      48318: inst = 32'h10a00000;
      48319: inst = 32'hca0bcc3;
      48320: inst = 32'h13e00001;
      48321: inst = 32'hfe0d96a;
      48322: inst = 32'h5be00000;
      48323: inst = 32'h8c50000;
      48324: inst = 32'h24612800;
      48325: inst = 32'h10a0ffff;
      48326: inst = 32'hca0ffe9;
      48327: inst = 32'h24822800;
      48328: inst = 32'h10a00000;
      48329: inst = 32'hca00004;
      48330: inst = 32'h38632800;
      48331: inst = 32'h38842800;
      48332: inst = 32'h10a00000;
      48333: inst = 32'hca0bcd1;
      48334: inst = 32'h13e00001;
      48335: inst = 32'hfe0d96a;
      48336: inst = 32'h5be00000;
      48337: inst = 32'h8c50000;
      48338: inst = 32'h24612800;
      48339: inst = 32'h10a0ffff;
      48340: inst = 32'hca0ffe9;
      48341: inst = 32'h24822800;
      48342: inst = 32'h10a00000;
      48343: inst = 32'hca00004;
      48344: inst = 32'h38632800;
      48345: inst = 32'h38842800;
      48346: inst = 32'h10a00000;
      48347: inst = 32'hca0bcdf;
      48348: inst = 32'h13e00001;
      48349: inst = 32'hfe0d96a;
      48350: inst = 32'h5be00000;
      48351: inst = 32'h8c50000;
      48352: inst = 32'h24612800;
      48353: inst = 32'h10a0ffff;
      48354: inst = 32'hca0ffe9;
      48355: inst = 32'h24822800;
      48356: inst = 32'h10a00000;
      48357: inst = 32'hca00004;
      48358: inst = 32'h38632800;
      48359: inst = 32'h38842800;
      48360: inst = 32'h10a00000;
      48361: inst = 32'hca0bced;
      48362: inst = 32'h13e00001;
      48363: inst = 32'hfe0d96a;
      48364: inst = 32'h5be00000;
      48365: inst = 32'h8c50000;
      48366: inst = 32'h24612800;
      48367: inst = 32'h10a0ffff;
      48368: inst = 32'hca0ffe9;
      48369: inst = 32'h24822800;
      48370: inst = 32'h10a00000;
      48371: inst = 32'hca00004;
      48372: inst = 32'h38632800;
      48373: inst = 32'h38842800;
      48374: inst = 32'h10a00000;
      48375: inst = 32'hca0bcfb;
      48376: inst = 32'h13e00001;
      48377: inst = 32'hfe0d96a;
      48378: inst = 32'h5be00000;
      48379: inst = 32'h8c50000;
      48380: inst = 32'h24612800;
      48381: inst = 32'h10a0ffff;
      48382: inst = 32'hca0ffe9;
      48383: inst = 32'h24822800;
      48384: inst = 32'h10a00000;
      48385: inst = 32'hca00004;
      48386: inst = 32'h38632800;
      48387: inst = 32'h38842800;
      48388: inst = 32'h10a00000;
      48389: inst = 32'hca0bd09;
      48390: inst = 32'h13e00001;
      48391: inst = 32'hfe0d96a;
      48392: inst = 32'h5be00000;
      48393: inst = 32'h8c50000;
      48394: inst = 32'h24612800;
      48395: inst = 32'h10a0ffff;
      48396: inst = 32'hca0ffe9;
      48397: inst = 32'h24822800;
      48398: inst = 32'h10a00000;
      48399: inst = 32'hca00004;
      48400: inst = 32'h38632800;
      48401: inst = 32'h38842800;
      48402: inst = 32'h10a00000;
      48403: inst = 32'hca0bd17;
      48404: inst = 32'h13e00001;
      48405: inst = 32'hfe0d96a;
      48406: inst = 32'h5be00000;
      48407: inst = 32'h8c50000;
      48408: inst = 32'h24612800;
      48409: inst = 32'h10a0ffff;
      48410: inst = 32'hca0ffe9;
      48411: inst = 32'h24822800;
      48412: inst = 32'h10a00000;
      48413: inst = 32'hca00004;
      48414: inst = 32'h38632800;
      48415: inst = 32'h38842800;
      48416: inst = 32'h10a00000;
      48417: inst = 32'hca0bd25;
      48418: inst = 32'h13e00001;
      48419: inst = 32'hfe0d96a;
      48420: inst = 32'h5be00000;
      48421: inst = 32'h8c50000;
      48422: inst = 32'h24612800;
      48423: inst = 32'h10a0ffff;
      48424: inst = 32'hca0ffe9;
      48425: inst = 32'h24822800;
      48426: inst = 32'h10a00000;
      48427: inst = 32'hca00004;
      48428: inst = 32'h38632800;
      48429: inst = 32'h38842800;
      48430: inst = 32'h10a00000;
      48431: inst = 32'hca0bd33;
      48432: inst = 32'h13e00001;
      48433: inst = 32'hfe0d96a;
      48434: inst = 32'h5be00000;
      48435: inst = 32'h8c50000;
      48436: inst = 32'h24612800;
      48437: inst = 32'h10a0ffff;
      48438: inst = 32'hca0ffe9;
      48439: inst = 32'h24822800;
      48440: inst = 32'h10a00000;
      48441: inst = 32'hca00004;
      48442: inst = 32'h38632800;
      48443: inst = 32'h38842800;
      48444: inst = 32'h10a00000;
      48445: inst = 32'hca0bd41;
      48446: inst = 32'h13e00001;
      48447: inst = 32'hfe0d96a;
      48448: inst = 32'h5be00000;
      48449: inst = 32'h8c50000;
      48450: inst = 32'h24612800;
      48451: inst = 32'h10a0ffff;
      48452: inst = 32'hca0ffe9;
      48453: inst = 32'h24822800;
      48454: inst = 32'h10a00000;
      48455: inst = 32'hca00004;
      48456: inst = 32'h38632800;
      48457: inst = 32'h38842800;
      48458: inst = 32'h10a00000;
      48459: inst = 32'hca0bd4f;
      48460: inst = 32'h13e00001;
      48461: inst = 32'hfe0d96a;
      48462: inst = 32'h5be00000;
      48463: inst = 32'h8c50000;
      48464: inst = 32'h24612800;
      48465: inst = 32'h10a0ffff;
      48466: inst = 32'hca0ffe9;
      48467: inst = 32'h24822800;
      48468: inst = 32'h10a00000;
      48469: inst = 32'hca00004;
      48470: inst = 32'h38632800;
      48471: inst = 32'h38842800;
      48472: inst = 32'h10a00000;
      48473: inst = 32'hca0bd5d;
      48474: inst = 32'h13e00001;
      48475: inst = 32'hfe0d96a;
      48476: inst = 32'h5be00000;
      48477: inst = 32'h8c50000;
      48478: inst = 32'h24612800;
      48479: inst = 32'h10a0ffff;
      48480: inst = 32'hca0ffe9;
      48481: inst = 32'h24822800;
      48482: inst = 32'h10a00000;
      48483: inst = 32'hca00004;
      48484: inst = 32'h38632800;
      48485: inst = 32'h38842800;
      48486: inst = 32'h10a00000;
      48487: inst = 32'hca0bd6b;
      48488: inst = 32'h13e00001;
      48489: inst = 32'hfe0d96a;
      48490: inst = 32'h5be00000;
      48491: inst = 32'h8c50000;
      48492: inst = 32'h24612800;
      48493: inst = 32'h10a0ffff;
      48494: inst = 32'hca0ffe9;
      48495: inst = 32'h24822800;
      48496: inst = 32'h10a00000;
      48497: inst = 32'hca00004;
      48498: inst = 32'h38632800;
      48499: inst = 32'h38842800;
      48500: inst = 32'h10a00000;
      48501: inst = 32'hca0bd79;
      48502: inst = 32'h13e00001;
      48503: inst = 32'hfe0d96a;
      48504: inst = 32'h5be00000;
      48505: inst = 32'h8c50000;
      48506: inst = 32'h24612800;
      48507: inst = 32'h10a0ffff;
      48508: inst = 32'hca0ffe9;
      48509: inst = 32'h24822800;
      48510: inst = 32'h10a00000;
      48511: inst = 32'hca00004;
      48512: inst = 32'h38632800;
      48513: inst = 32'h38842800;
      48514: inst = 32'h10a00000;
      48515: inst = 32'hca0bd87;
      48516: inst = 32'h13e00001;
      48517: inst = 32'hfe0d96a;
      48518: inst = 32'h5be00000;
      48519: inst = 32'h8c50000;
      48520: inst = 32'h24612800;
      48521: inst = 32'h10a0ffff;
      48522: inst = 32'hca0ffe9;
      48523: inst = 32'h24822800;
      48524: inst = 32'h10a00000;
      48525: inst = 32'hca00004;
      48526: inst = 32'h38632800;
      48527: inst = 32'h38842800;
      48528: inst = 32'h10a00000;
      48529: inst = 32'hca0bd95;
      48530: inst = 32'h13e00001;
      48531: inst = 32'hfe0d96a;
      48532: inst = 32'h5be00000;
      48533: inst = 32'h8c50000;
      48534: inst = 32'h24612800;
      48535: inst = 32'h10a0ffff;
      48536: inst = 32'hca0ffe9;
      48537: inst = 32'h24822800;
      48538: inst = 32'h10a00000;
      48539: inst = 32'hca00004;
      48540: inst = 32'h38632800;
      48541: inst = 32'h38842800;
      48542: inst = 32'h10a00000;
      48543: inst = 32'hca0bda3;
      48544: inst = 32'h13e00001;
      48545: inst = 32'hfe0d96a;
      48546: inst = 32'h5be00000;
      48547: inst = 32'h8c50000;
      48548: inst = 32'h24612800;
      48549: inst = 32'h10a0ffff;
      48550: inst = 32'hca0ffe9;
      48551: inst = 32'h24822800;
      48552: inst = 32'h10a00000;
      48553: inst = 32'hca00004;
      48554: inst = 32'h38632800;
      48555: inst = 32'h38842800;
      48556: inst = 32'h10a00000;
      48557: inst = 32'hca0bdb1;
      48558: inst = 32'h13e00001;
      48559: inst = 32'hfe0d96a;
      48560: inst = 32'h5be00000;
      48561: inst = 32'h8c50000;
      48562: inst = 32'h24612800;
      48563: inst = 32'h10a0ffff;
      48564: inst = 32'hca0ffe9;
      48565: inst = 32'h24822800;
      48566: inst = 32'h10a00000;
      48567: inst = 32'hca00004;
      48568: inst = 32'h38632800;
      48569: inst = 32'h38842800;
      48570: inst = 32'h10a00000;
      48571: inst = 32'hca0bdbf;
      48572: inst = 32'h13e00001;
      48573: inst = 32'hfe0d96a;
      48574: inst = 32'h5be00000;
      48575: inst = 32'h8c50000;
      48576: inst = 32'h24612800;
      48577: inst = 32'h10a0ffff;
      48578: inst = 32'hca0ffe9;
      48579: inst = 32'h24822800;
      48580: inst = 32'h10a00000;
      48581: inst = 32'hca00004;
      48582: inst = 32'h38632800;
      48583: inst = 32'h38842800;
      48584: inst = 32'h10a00000;
      48585: inst = 32'hca0bdcd;
      48586: inst = 32'h13e00001;
      48587: inst = 32'hfe0d96a;
      48588: inst = 32'h5be00000;
      48589: inst = 32'h8c50000;
      48590: inst = 32'h24612800;
      48591: inst = 32'h10a0ffff;
      48592: inst = 32'hca0ffe9;
      48593: inst = 32'h24822800;
      48594: inst = 32'h10a00000;
      48595: inst = 32'hca00004;
      48596: inst = 32'h38632800;
      48597: inst = 32'h38842800;
      48598: inst = 32'h10a00000;
      48599: inst = 32'hca0bddb;
      48600: inst = 32'h13e00001;
      48601: inst = 32'hfe0d96a;
      48602: inst = 32'h5be00000;
      48603: inst = 32'h8c50000;
      48604: inst = 32'h24612800;
      48605: inst = 32'h10a0ffff;
      48606: inst = 32'hca0ffe9;
      48607: inst = 32'h24822800;
      48608: inst = 32'h10a00000;
      48609: inst = 32'hca00004;
      48610: inst = 32'h38632800;
      48611: inst = 32'h38842800;
      48612: inst = 32'h10a00000;
      48613: inst = 32'hca0bde9;
      48614: inst = 32'h13e00001;
      48615: inst = 32'hfe0d96a;
      48616: inst = 32'h5be00000;
      48617: inst = 32'h8c50000;
      48618: inst = 32'h24612800;
      48619: inst = 32'h10a0ffff;
      48620: inst = 32'hca0ffea;
      48621: inst = 32'h24822800;
      48622: inst = 32'h10a00000;
      48623: inst = 32'hca00004;
      48624: inst = 32'h38632800;
      48625: inst = 32'h38842800;
      48626: inst = 32'h10a00000;
      48627: inst = 32'hca0bdf7;
      48628: inst = 32'h13e00001;
      48629: inst = 32'hfe0d96a;
      48630: inst = 32'h5be00000;
      48631: inst = 32'h8c50000;
      48632: inst = 32'h24612800;
      48633: inst = 32'h10a0ffff;
      48634: inst = 32'hca0ffea;
      48635: inst = 32'h24822800;
      48636: inst = 32'h10a00000;
      48637: inst = 32'hca00004;
      48638: inst = 32'h38632800;
      48639: inst = 32'h38842800;
      48640: inst = 32'h10a00000;
      48641: inst = 32'hca0be05;
      48642: inst = 32'h13e00001;
      48643: inst = 32'hfe0d96a;
      48644: inst = 32'h5be00000;
      48645: inst = 32'h8c50000;
      48646: inst = 32'h24612800;
      48647: inst = 32'h10a0ffff;
      48648: inst = 32'hca0ffea;
      48649: inst = 32'h24822800;
      48650: inst = 32'h10a00000;
      48651: inst = 32'hca00004;
      48652: inst = 32'h38632800;
      48653: inst = 32'h38842800;
      48654: inst = 32'h10a00000;
      48655: inst = 32'hca0be13;
      48656: inst = 32'h13e00001;
      48657: inst = 32'hfe0d96a;
      48658: inst = 32'h5be00000;
      48659: inst = 32'h8c50000;
      48660: inst = 32'h24612800;
      48661: inst = 32'h10a0ffff;
      48662: inst = 32'hca0ffea;
      48663: inst = 32'h24822800;
      48664: inst = 32'h10a00000;
      48665: inst = 32'hca00004;
      48666: inst = 32'h38632800;
      48667: inst = 32'h38842800;
      48668: inst = 32'h10a00000;
      48669: inst = 32'hca0be21;
      48670: inst = 32'h13e00001;
      48671: inst = 32'hfe0d96a;
      48672: inst = 32'h5be00000;
      48673: inst = 32'h8c50000;
      48674: inst = 32'h24612800;
      48675: inst = 32'h10a0ffff;
      48676: inst = 32'hca0ffea;
      48677: inst = 32'h24822800;
      48678: inst = 32'h10a00000;
      48679: inst = 32'hca00004;
      48680: inst = 32'h38632800;
      48681: inst = 32'h38842800;
      48682: inst = 32'h10a00000;
      48683: inst = 32'hca0be2f;
      48684: inst = 32'h13e00001;
      48685: inst = 32'hfe0d96a;
      48686: inst = 32'h5be00000;
      48687: inst = 32'h8c50000;
      48688: inst = 32'h24612800;
      48689: inst = 32'h10a0ffff;
      48690: inst = 32'hca0ffea;
      48691: inst = 32'h24822800;
      48692: inst = 32'h10a00000;
      48693: inst = 32'hca00004;
      48694: inst = 32'h38632800;
      48695: inst = 32'h38842800;
      48696: inst = 32'h10a00000;
      48697: inst = 32'hca0be3d;
      48698: inst = 32'h13e00001;
      48699: inst = 32'hfe0d96a;
      48700: inst = 32'h5be00000;
      48701: inst = 32'h8c50000;
      48702: inst = 32'h24612800;
      48703: inst = 32'h10a0ffff;
      48704: inst = 32'hca0ffea;
      48705: inst = 32'h24822800;
      48706: inst = 32'h10a00000;
      48707: inst = 32'hca00004;
      48708: inst = 32'h38632800;
      48709: inst = 32'h38842800;
      48710: inst = 32'h10a00000;
      48711: inst = 32'hca0be4b;
      48712: inst = 32'h13e00001;
      48713: inst = 32'hfe0d96a;
      48714: inst = 32'h5be00000;
      48715: inst = 32'h8c50000;
      48716: inst = 32'h24612800;
      48717: inst = 32'h10a0ffff;
      48718: inst = 32'hca0ffea;
      48719: inst = 32'h24822800;
      48720: inst = 32'h10a00000;
      48721: inst = 32'hca00004;
      48722: inst = 32'h38632800;
      48723: inst = 32'h38842800;
      48724: inst = 32'h10a00000;
      48725: inst = 32'hca0be59;
      48726: inst = 32'h13e00001;
      48727: inst = 32'hfe0d96a;
      48728: inst = 32'h5be00000;
      48729: inst = 32'h8c50000;
      48730: inst = 32'h24612800;
      48731: inst = 32'h10a0ffff;
      48732: inst = 32'hca0ffea;
      48733: inst = 32'h24822800;
      48734: inst = 32'h10a00000;
      48735: inst = 32'hca00004;
      48736: inst = 32'h38632800;
      48737: inst = 32'h38842800;
      48738: inst = 32'h10a00000;
      48739: inst = 32'hca0be67;
      48740: inst = 32'h13e00001;
      48741: inst = 32'hfe0d96a;
      48742: inst = 32'h5be00000;
      48743: inst = 32'h8c50000;
      48744: inst = 32'h24612800;
      48745: inst = 32'h10a0ffff;
      48746: inst = 32'hca0ffea;
      48747: inst = 32'h24822800;
      48748: inst = 32'h10a00000;
      48749: inst = 32'hca00004;
      48750: inst = 32'h38632800;
      48751: inst = 32'h38842800;
      48752: inst = 32'h10a00000;
      48753: inst = 32'hca0be75;
      48754: inst = 32'h13e00001;
      48755: inst = 32'hfe0d96a;
      48756: inst = 32'h5be00000;
      48757: inst = 32'h8c50000;
      48758: inst = 32'h24612800;
      48759: inst = 32'h10a0ffff;
      48760: inst = 32'hca0ffea;
      48761: inst = 32'h24822800;
      48762: inst = 32'h10a00000;
      48763: inst = 32'hca00004;
      48764: inst = 32'h38632800;
      48765: inst = 32'h38842800;
      48766: inst = 32'h10a00000;
      48767: inst = 32'hca0be83;
      48768: inst = 32'h13e00001;
      48769: inst = 32'hfe0d96a;
      48770: inst = 32'h5be00000;
      48771: inst = 32'h8c50000;
      48772: inst = 32'h24612800;
      48773: inst = 32'h10a0ffff;
      48774: inst = 32'hca0ffea;
      48775: inst = 32'h24822800;
      48776: inst = 32'h10a00000;
      48777: inst = 32'hca00004;
      48778: inst = 32'h38632800;
      48779: inst = 32'h38842800;
      48780: inst = 32'h10a00000;
      48781: inst = 32'hca0be91;
      48782: inst = 32'h13e00001;
      48783: inst = 32'hfe0d96a;
      48784: inst = 32'h5be00000;
      48785: inst = 32'h8c50000;
      48786: inst = 32'h24612800;
      48787: inst = 32'h10a0ffff;
      48788: inst = 32'hca0ffea;
      48789: inst = 32'h24822800;
      48790: inst = 32'h10a00000;
      48791: inst = 32'hca00004;
      48792: inst = 32'h38632800;
      48793: inst = 32'h38842800;
      48794: inst = 32'h10a00000;
      48795: inst = 32'hca0be9f;
      48796: inst = 32'h13e00001;
      48797: inst = 32'hfe0d96a;
      48798: inst = 32'h5be00000;
      48799: inst = 32'h8c50000;
      48800: inst = 32'h24612800;
      48801: inst = 32'h10a0ffff;
      48802: inst = 32'hca0ffea;
      48803: inst = 32'h24822800;
      48804: inst = 32'h10a00000;
      48805: inst = 32'hca00004;
      48806: inst = 32'h38632800;
      48807: inst = 32'h38842800;
      48808: inst = 32'h10a00000;
      48809: inst = 32'hca0bead;
      48810: inst = 32'h13e00001;
      48811: inst = 32'hfe0d96a;
      48812: inst = 32'h5be00000;
      48813: inst = 32'h8c50000;
      48814: inst = 32'h24612800;
      48815: inst = 32'h10a0ffff;
      48816: inst = 32'hca0ffea;
      48817: inst = 32'h24822800;
      48818: inst = 32'h10a00000;
      48819: inst = 32'hca00004;
      48820: inst = 32'h38632800;
      48821: inst = 32'h38842800;
      48822: inst = 32'h10a00000;
      48823: inst = 32'hca0bebb;
      48824: inst = 32'h13e00001;
      48825: inst = 32'hfe0d96a;
      48826: inst = 32'h5be00000;
      48827: inst = 32'h8c50000;
      48828: inst = 32'h24612800;
      48829: inst = 32'h10a0ffff;
      48830: inst = 32'hca0ffea;
      48831: inst = 32'h24822800;
      48832: inst = 32'h10a00000;
      48833: inst = 32'hca00004;
      48834: inst = 32'h38632800;
      48835: inst = 32'h38842800;
      48836: inst = 32'h10a00000;
      48837: inst = 32'hca0bec9;
      48838: inst = 32'h13e00001;
      48839: inst = 32'hfe0d96a;
      48840: inst = 32'h5be00000;
      48841: inst = 32'h8c50000;
      48842: inst = 32'h24612800;
      48843: inst = 32'h10a0ffff;
      48844: inst = 32'hca0ffea;
      48845: inst = 32'h24822800;
      48846: inst = 32'h10a00000;
      48847: inst = 32'hca00004;
      48848: inst = 32'h38632800;
      48849: inst = 32'h38842800;
      48850: inst = 32'h10a00000;
      48851: inst = 32'hca0bed7;
      48852: inst = 32'h13e00001;
      48853: inst = 32'hfe0d96a;
      48854: inst = 32'h5be00000;
      48855: inst = 32'h8c50000;
      48856: inst = 32'h24612800;
      48857: inst = 32'h10a0ffff;
      48858: inst = 32'hca0ffea;
      48859: inst = 32'h24822800;
      48860: inst = 32'h10a00000;
      48861: inst = 32'hca00004;
      48862: inst = 32'h38632800;
      48863: inst = 32'h38842800;
      48864: inst = 32'h10a00000;
      48865: inst = 32'hca0bee5;
      48866: inst = 32'h13e00001;
      48867: inst = 32'hfe0d96a;
      48868: inst = 32'h5be00000;
      48869: inst = 32'h8c50000;
      48870: inst = 32'h24612800;
      48871: inst = 32'h10a0ffff;
      48872: inst = 32'hca0ffea;
      48873: inst = 32'h24822800;
      48874: inst = 32'h10a00000;
      48875: inst = 32'hca00004;
      48876: inst = 32'h38632800;
      48877: inst = 32'h38842800;
      48878: inst = 32'h10a00000;
      48879: inst = 32'hca0bef3;
      48880: inst = 32'h13e00001;
      48881: inst = 32'hfe0d96a;
      48882: inst = 32'h5be00000;
      48883: inst = 32'h8c50000;
      48884: inst = 32'h24612800;
      48885: inst = 32'h10a0ffff;
      48886: inst = 32'hca0ffea;
      48887: inst = 32'h24822800;
      48888: inst = 32'h10a00000;
      48889: inst = 32'hca00004;
      48890: inst = 32'h38632800;
      48891: inst = 32'h38842800;
      48892: inst = 32'h10a00000;
      48893: inst = 32'hca0bf01;
      48894: inst = 32'h13e00001;
      48895: inst = 32'hfe0d96a;
      48896: inst = 32'h5be00000;
      48897: inst = 32'h8c50000;
      48898: inst = 32'h24612800;
      48899: inst = 32'h10a0ffff;
      48900: inst = 32'hca0ffea;
      48901: inst = 32'h24822800;
      48902: inst = 32'h10a00000;
      48903: inst = 32'hca00004;
      48904: inst = 32'h38632800;
      48905: inst = 32'h38842800;
      48906: inst = 32'h10a00000;
      48907: inst = 32'hca0bf0f;
      48908: inst = 32'h13e00001;
      48909: inst = 32'hfe0d96a;
      48910: inst = 32'h5be00000;
      48911: inst = 32'h8c50000;
      48912: inst = 32'h24612800;
      48913: inst = 32'h10a0ffff;
      48914: inst = 32'hca0ffea;
      48915: inst = 32'h24822800;
      48916: inst = 32'h10a00000;
      48917: inst = 32'hca00004;
      48918: inst = 32'h38632800;
      48919: inst = 32'h38842800;
      48920: inst = 32'h10a00000;
      48921: inst = 32'hca0bf1d;
      48922: inst = 32'h13e00001;
      48923: inst = 32'hfe0d96a;
      48924: inst = 32'h5be00000;
      48925: inst = 32'h8c50000;
      48926: inst = 32'h24612800;
      48927: inst = 32'h10a0ffff;
      48928: inst = 32'hca0ffea;
      48929: inst = 32'h24822800;
      48930: inst = 32'h10a00000;
      48931: inst = 32'hca00004;
      48932: inst = 32'h38632800;
      48933: inst = 32'h38842800;
      48934: inst = 32'h10a00000;
      48935: inst = 32'hca0bf2b;
      48936: inst = 32'h13e00001;
      48937: inst = 32'hfe0d96a;
      48938: inst = 32'h5be00000;
      48939: inst = 32'h8c50000;
      48940: inst = 32'h24612800;
      48941: inst = 32'h10a0ffff;
      48942: inst = 32'hca0ffea;
      48943: inst = 32'h24822800;
      48944: inst = 32'h10a00000;
      48945: inst = 32'hca00004;
      48946: inst = 32'h38632800;
      48947: inst = 32'h38842800;
      48948: inst = 32'h10a00000;
      48949: inst = 32'hca0bf39;
      48950: inst = 32'h13e00001;
      48951: inst = 32'hfe0d96a;
      48952: inst = 32'h5be00000;
      48953: inst = 32'h8c50000;
      48954: inst = 32'h24612800;
      48955: inst = 32'h10a0ffff;
      48956: inst = 32'hca0ffea;
      48957: inst = 32'h24822800;
      48958: inst = 32'h10a00000;
      48959: inst = 32'hca00004;
      48960: inst = 32'h38632800;
      48961: inst = 32'h38842800;
      48962: inst = 32'h10a00000;
      48963: inst = 32'hca0bf47;
      48964: inst = 32'h13e00001;
      48965: inst = 32'hfe0d96a;
      48966: inst = 32'h5be00000;
      48967: inst = 32'h8c50000;
      48968: inst = 32'h24612800;
      48969: inst = 32'h10a0ffff;
      48970: inst = 32'hca0ffea;
      48971: inst = 32'h24822800;
      48972: inst = 32'h10a00000;
      48973: inst = 32'hca00004;
      48974: inst = 32'h38632800;
      48975: inst = 32'h38842800;
      48976: inst = 32'h10a00000;
      48977: inst = 32'hca0bf55;
      48978: inst = 32'h13e00001;
      48979: inst = 32'hfe0d96a;
      48980: inst = 32'h5be00000;
      48981: inst = 32'h8c50000;
      48982: inst = 32'h24612800;
      48983: inst = 32'h10a0ffff;
      48984: inst = 32'hca0ffea;
      48985: inst = 32'h24822800;
      48986: inst = 32'h10a00000;
      48987: inst = 32'hca00004;
      48988: inst = 32'h38632800;
      48989: inst = 32'h38842800;
      48990: inst = 32'h10a00000;
      48991: inst = 32'hca0bf63;
      48992: inst = 32'h13e00001;
      48993: inst = 32'hfe0d96a;
      48994: inst = 32'h5be00000;
      48995: inst = 32'h8c50000;
      48996: inst = 32'h24612800;
      48997: inst = 32'h10a0ffff;
      48998: inst = 32'hca0ffea;
      48999: inst = 32'h24822800;
      49000: inst = 32'h10a00000;
      49001: inst = 32'hca00004;
      49002: inst = 32'h38632800;
      49003: inst = 32'h38842800;
      49004: inst = 32'h10a00000;
      49005: inst = 32'hca0bf71;
      49006: inst = 32'h13e00001;
      49007: inst = 32'hfe0d96a;
      49008: inst = 32'h5be00000;
      49009: inst = 32'h8c50000;
      49010: inst = 32'h24612800;
      49011: inst = 32'h10a0ffff;
      49012: inst = 32'hca0ffea;
      49013: inst = 32'h24822800;
      49014: inst = 32'h10a00000;
      49015: inst = 32'hca00004;
      49016: inst = 32'h38632800;
      49017: inst = 32'h38842800;
      49018: inst = 32'h10a00000;
      49019: inst = 32'hca0bf7f;
      49020: inst = 32'h13e00001;
      49021: inst = 32'hfe0d96a;
      49022: inst = 32'h5be00000;
      49023: inst = 32'h8c50000;
      49024: inst = 32'h24612800;
      49025: inst = 32'h10a0ffff;
      49026: inst = 32'hca0ffea;
      49027: inst = 32'h24822800;
      49028: inst = 32'h10a00000;
      49029: inst = 32'hca00004;
      49030: inst = 32'h38632800;
      49031: inst = 32'h38842800;
      49032: inst = 32'h10a00000;
      49033: inst = 32'hca0bf8d;
      49034: inst = 32'h13e00001;
      49035: inst = 32'hfe0d96a;
      49036: inst = 32'h5be00000;
      49037: inst = 32'h8c50000;
      49038: inst = 32'h24612800;
      49039: inst = 32'h10a0ffff;
      49040: inst = 32'hca0ffea;
      49041: inst = 32'h24822800;
      49042: inst = 32'h10a00000;
      49043: inst = 32'hca00004;
      49044: inst = 32'h38632800;
      49045: inst = 32'h38842800;
      49046: inst = 32'h10a00000;
      49047: inst = 32'hca0bf9b;
      49048: inst = 32'h13e00001;
      49049: inst = 32'hfe0d96a;
      49050: inst = 32'h5be00000;
      49051: inst = 32'h8c50000;
      49052: inst = 32'h24612800;
      49053: inst = 32'h10a0ffff;
      49054: inst = 32'hca0ffea;
      49055: inst = 32'h24822800;
      49056: inst = 32'h10a00000;
      49057: inst = 32'hca00004;
      49058: inst = 32'h38632800;
      49059: inst = 32'h38842800;
      49060: inst = 32'h10a00000;
      49061: inst = 32'hca0bfa9;
      49062: inst = 32'h13e00001;
      49063: inst = 32'hfe0d96a;
      49064: inst = 32'h5be00000;
      49065: inst = 32'h8c50000;
      49066: inst = 32'h24612800;
      49067: inst = 32'h10a0ffff;
      49068: inst = 32'hca0ffea;
      49069: inst = 32'h24822800;
      49070: inst = 32'h10a00000;
      49071: inst = 32'hca00004;
      49072: inst = 32'h38632800;
      49073: inst = 32'h38842800;
      49074: inst = 32'h10a00000;
      49075: inst = 32'hca0bfb7;
      49076: inst = 32'h13e00001;
      49077: inst = 32'hfe0d96a;
      49078: inst = 32'h5be00000;
      49079: inst = 32'h8c50000;
      49080: inst = 32'h24612800;
      49081: inst = 32'h10a0ffff;
      49082: inst = 32'hca0ffea;
      49083: inst = 32'h24822800;
      49084: inst = 32'h10a00000;
      49085: inst = 32'hca00004;
      49086: inst = 32'h38632800;
      49087: inst = 32'h38842800;
      49088: inst = 32'h10a00000;
      49089: inst = 32'hca0bfc5;
      49090: inst = 32'h13e00001;
      49091: inst = 32'hfe0d96a;
      49092: inst = 32'h5be00000;
      49093: inst = 32'h8c50000;
      49094: inst = 32'h24612800;
      49095: inst = 32'h10a0ffff;
      49096: inst = 32'hca0ffea;
      49097: inst = 32'h24822800;
      49098: inst = 32'h10a00000;
      49099: inst = 32'hca00004;
      49100: inst = 32'h38632800;
      49101: inst = 32'h38842800;
      49102: inst = 32'h10a00000;
      49103: inst = 32'hca0bfd3;
      49104: inst = 32'h13e00001;
      49105: inst = 32'hfe0d96a;
      49106: inst = 32'h5be00000;
      49107: inst = 32'h8c50000;
      49108: inst = 32'h24612800;
      49109: inst = 32'h10a0ffff;
      49110: inst = 32'hca0ffea;
      49111: inst = 32'h24822800;
      49112: inst = 32'h10a00000;
      49113: inst = 32'hca00004;
      49114: inst = 32'h38632800;
      49115: inst = 32'h38842800;
      49116: inst = 32'h10a00000;
      49117: inst = 32'hca0bfe1;
      49118: inst = 32'h13e00001;
      49119: inst = 32'hfe0d96a;
      49120: inst = 32'h5be00000;
      49121: inst = 32'h8c50000;
      49122: inst = 32'h24612800;
      49123: inst = 32'h10a0ffff;
      49124: inst = 32'hca0ffea;
      49125: inst = 32'h24822800;
      49126: inst = 32'h10a00000;
      49127: inst = 32'hca00004;
      49128: inst = 32'h38632800;
      49129: inst = 32'h38842800;
      49130: inst = 32'h10a00000;
      49131: inst = 32'hca0bfef;
      49132: inst = 32'h13e00001;
      49133: inst = 32'hfe0d96a;
      49134: inst = 32'h5be00000;
      49135: inst = 32'h8c50000;
      49136: inst = 32'h24612800;
      49137: inst = 32'h10a0ffff;
      49138: inst = 32'hca0ffea;
      49139: inst = 32'h24822800;
      49140: inst = 32'h10a00000;
      49141: inst = 32'hca00004;
      49142: inst = 32'h38632800;
      49143: inst = 32'h38842800;
      49144: inst = 32'h10a00000;
      49145: inst = 32'hca0bffd;
      49146: inst = 32'h13e00001;
      49147: inst = 32'hfe0d96a;
      49148: inst = 32'h5be00000;
      49149: inst = 32'h8c50000;
      49150: inst = 32'h24612800;
      49151: inst = 32'h10a0ffff;
      49152: inst = 32'hca0ffea;
      49153: inst = 32'h24822800;
      49154: inst = 32'h10a00000;
      49155: inst = 32'hca00004;
      49156: inst = 32'h38632800;
      49157: inst = 32'h38842800;
      49158: inst = 32'h10a00000;
      49159: inst = 32'hca0c00b;
      49160: inst = 32'h13e00001;
      49161: inst = 32'hfe0d96a;
      49162: inst = 32'h5be00000;
      49163: inst = 32'h8c50000;
      49164: inst = 32'h24612800;
      49165: inst = 32'h10a0ffff;
      49166: inst = 32'hca0ffea;
      49167: inst = 32'h24822800;
      49168: inst = 32'h10a00000;
      49169: inst = 32'hca00004;
      49170: inst = 32'h38632800;
      49171: inst = 32'h38842800;
      49172: inst = 32'h10a00000;
      49173: inst = 32'hca0c019;
      49174: inst = 32'h13e00001;
      49175: inst = 32'hfe0d96a;
      49176: inst = 32'h5be00000;
      49177: inst = 32'h8c50000;
      49178: inst = 32'h24612800;
      49179: inst = 32'h10a0ffff;
      49180: inst = 32'hca0ffea;
      49181: inst = 32'h24822800;
      49182: inst = 32'h10a00000;
      49183: inst = 32'hca00004;
      49184: inst = 32'h38632800;
      49185: inst = 32'h38842800;
      49186: inst = 32'h10a00000;
      49187: inst = 32'hca0c027;
      49188: inst = 32'h13e00001;
      49189: inst = 32'hfe0d96a;
      49190: inst = 32'h5be00000;
      49191: inst = 32'h8c50000;
      49192: inst = 32'h24612800;
      49193: inst = 32'h10a0ffff;
      49194: inst = 32'hca0ffea;
      49195: inst = 32'h24822800;
      49196: inst = 32'h10a00000;
      49197: inst = 32'hca00004;
      49198: inst = 32'h38632800;
      49199: inst = 32'h38842800;
      49200: inst = 32'h10a00000;
      49201: inst = 32'hca0c035;
      49202: inst = 32'h13e00001;
      49203: inst = 32'hfe0d96a;
      49204: inst = 32'h5be00000;
      49205: inst = 32'h8c50000;
      49206: inst = 32'h24612800;
      49207: inst = 32'h10a0ffff;
      49208: inst = 32'hca0ffea;
      49209: inst = 32'h24822800;
      49210: inst = 32'h10a00000;
      49211: inst = 32'hca00004;
      49212: inst = 32'h38632800;
      49213: inst = 32'h38842800;
      49214: inst = 32'h10a00000;
      49215: inst = 32'hca0c043;
      49216: inst = 32'h13e00001;
      49217: inst = 32'hfe0d96a;
      49218: inst = 32'h5be00000;
      49219: inst = 32'h8c50000;
      49220: inst = 32'h24612800;
      49221: inst = 32'h10a0ffff;
      49222: inst = 32'hca0ffea;
      49223: inst = 32'h24822800;
      49224: inst = 32'h10a00000;
      49225: inst = 32'hca00004;
      49226: inst = 32'h38632800;
      49227: inst = 32'h38842800;
      49228: inst = 32'h10a00000;
      49229: inst = 32'hca0c051;
      49230: inst = 32'h13e00001;
      49231: inst = 32'hfe0d96a;
      49232: inst = 32'h5be00000;
      49233: inst = 32'h8c50000;
      49234: inst = 32'h24612800;
      49235: inst = 32'h10a0ffff;
      49236: inst = 32'hca0ffea;
      49237: inst = 32'h24822800;
      49238: inst = 32'h10a00000;
      49239: inst = 32'hca00004;
      49240: inst = 32'h38632800;
      49241: inst = 32'h38842800;
      49242: inst = 32'h10a00000;
      49243: inst = 32'hca0c05f;
      49244: inst = 32'h13e00001;
      49245: inst = 32'hfe0d96a;
      49246: inst = 32'h5be00000;
      49247: inst = 32'h8c50000;
      49248: inst = 32'h24612800;
      49249: inst = 32'h10a0ffff;
      49250: inst = 32'hca0ffea;
      49251: inst = 32'h24822800;
      49252: inst = 32'h10a00000;
      49253: inst = 32'hca00004;
      49254: inst = 32'h38632800;
      49255: inst = 32'h38842800;
      49256: inst = 32'h10a00000;
      49257: inst = 32'hca0c06d;
      49258: inst = 32'h13e00001;
      49259: inst = 32'hfe0d96a;
      49260: inst = 32'h5be00000;
      49261: inst = 32'h8c50000;
      49262: inst = 32'h24612800;
      49263: inst = 32'h10a0ffff;
      49264: inst = 32'hca0ffea;
      49265: inst = 32'h24822800;
      49266: inst = 32'h10a00000;
      49267: inst = 32'hca00004;
      49268: inst = 32'h38632800;
      49269: inst = 32'h38842800;
      49270: inst = 32'h10a00000;
      49271: inst = 32'hca0c07b;
      49272: inst = 32'h13e00001;
      49273: inst = 32'hfe0d96a;
      49274: inst = 32'h5be00000;
      49275: inst = 32'h8c50000;
      49276: inst = 32'h24612800;
      49277: inst = 32'h10a0ffff;
      49278: inst = 32'hca0ffea;
      49279: inst = 32'h24822800;
      49280: inst = 32'h10a00000;
      49281: inst = 32'hca00004;
      49282: inst = 32'h38632800;
      49283: inst = 32'h38842800;
      49284: inst = 32'h10a00000;
      49285: inst = 32'hca0c089;
      49286: inst = 32'h13e00001;
      49287: inst = 32'hfe0d96a;
      49288: inst = 32'h5be00000;
      49289: inst = 32'h8c50000;
      49290: inst = 32'h24612800;
      49291: inst = 32'h10a0ffff;
      49292: inst = 32'hca0ffea;
      49293: inst = 32'h24822800;
      49294: inst = 32'h10a00000;
      49295: inst = 32'hca00004;
      49296: inst = 32'h38632800;
      49297: inst = 32'h38842800;
      49298: inst = 32'h10a00000;
      49299: inst = 32'hca0c097;
      49300: inst = 32'h13e00001;
      49301: inst = 32'hfe0d96a;
      49302: inst = 32'h5be00000;
      49303: inst = 32'h8c50000;
      49304: inst = 32'h24612800;
      49305: inst = 32'h10a0ffff;
      49306: inst = 32'hca0ffea;
      49307: inst = 32'h24822800;
      49308: inst = 32'h10a00000;
      49309: inst = 32'hca00004;
      49310: inst = 32'h38632800;
      49311: inst = 32'h38842800;
      49312: inst = 32'h10a00000;
      49313: inst = 32'hca0c0a5;
      49314: inst = 32'h13e00001;
      49315: inst = 32'hfe0d96a;
      49316: inst = 32'h5be00000;
      49317: inst = 32'h8c50000;
      49318: inst = 32'h24612800;
      49319: inst = 32'h10a0ffff;
      49320: inst = 32'hca0ffea;
      49321: inst = 32'h24822800;
      49322: inst = 32'h10a00000;
      49323: inst = 32'hca00004;
      49324: inst = 32'h38632800;
      49325: inst = 32'h38842800;
      49326: inst = 32'h10a00000;
      49327: inst = 32'hca0c0b3;
      49328: inst = 32'h13e00001;
      49329: inst = 32'hfe0d96a;
      49330: inst = 32'h5be00000;
      49331: inst = 32'h8c50000;
      49332: inst = 32'h24612800;
      49333: inst = 32'h10a0ffff;
      49334: inst = 32'hca0ffea;
      49335: inst = 32'h24822800;
      49336: inst = 32'h10a00000;
      49337: inst = 32'hca00004;
      49338: inst = 32'h38632800;
      49339: inst = 32'h38842800;
      49340: inst = 32'h10a00000;
      49341: inst = 32'hca0c0c1;
      49342: inst = 32'h13e00001;
      49343: inst = 32'hfe0d96a;
      49344: inst = 32'h5be00000;
      49345: inst = 32'h8c50000;
      49346: inst = 32'h24612800;
      49347: inst = 32'h10a0ffff;
      49348: inst = 32'hca0ffea;
      49349: inst = 32'h24822800;
      49350: inst = 32'h10a00000;
      49351: inst = 32'hca00004;
      49352: inst = 32'h38632800;
      49353: inst = 32'h38842800;
      49354: inst = 32'h10a00000;
      49355: inst = 32'hca0c0cf;
      49356: inst = 32'h13e00001;
      49357: inst = 32'hfe0d96a;
      49358: inst = 32'h5be00000;
      49359: inst = 32'h8c50000;
      49360: inst = 32'h24612800;
      49361: inst = 32'h10a0ffff;
      49362: inst = 32'hca0ffea;
      49363: inst = 32'h24822800;
      49364: inst = 32'h10a00000;
      49365: inst = 32'hca00004;
      49366: inst = 32'h38632800;
      49367: inst = 32'h38842800;
      49368: inst = 32'h10a00000;
      49369: inst = 32'hca0c0dd;
      49370: inst = 32'h13e00001;
      49371: inst = 32'hfe0d96a;
      49372: inst = 32'h5be00000;
      49373: inst = 32'h8c50000;
      49374: inst = 32'h24612800;
      49375: inst = 32'h10a0ffff;
      49376: inst = 32'hca0ffea;
      49377: inst = 32'h24822800;
      49378: inst = 32'h10a00000;
      49379: inst = 32'hca00004;
      49380: inst = 32'h38632800;
      49381: inst = 32'h38842800;
      49382: inst = 32'h10a00000;
      49383: inst = 32'hca0c0eb;
      49384: inst = 32'h13e00001;
      49385: inst = 32'hfe0d96a;
      49386: inst = 32'h5be00000;
      49387: inst = 32'h8c50000;
      49388: inst = 32'h24612800;
      49389: inst = 32'h10a0ffff;
      49390: inst = 32'hca0ffea;
      49391: inst = 32'h24822800;
      49392: inst = 32'h10a00000;
      49393: inst = 32'hca00004;
      49394: inst = 32'h38632800;
      49395: inst = 32'h38842800;
      49396: inst = 32'h10a00000;
      49397: inst = 32'hca0c0f9;
      49398: inst = 32'h13e00001;
      49399: inst = 32'hfe0d96a;
      49400: inst = 32'h5be00000;
      49401: inst = 32'h8c50000;
      49402: inst = 32'h24612800;
      49403: inst = 32'h10a0ffff;
      49404: inst = 32'hca0ffea;
      49405: inst = 32'h24822800;
      49406: inst = 32'h10a00000;
      49407: inst = 32'hca00004;
      49408: inst = 32'h38632800;
      49409: inst = 32'h38842800;
      49410: inst = 32'h10a00000;
      49411: inst = 32'hca0c107;
      49412: inst = 32'h13e00001;
      49413: inst = 32'hfe0d96a;
      49414: inst = 32'h5be00000;
      49415: inst = 32'h8c50000;
      49416: inst = 32'h24612800;
      49417: inst = 32'h10a0ffff;
      49418: inst = 32'hca0ffea;
      49419: inst = 32'h24822800;
      49420: inst = 32'h10a00000;
      49421: inst = 32'hca00004;
      49422: inst = 32'h38632800;
      49423: inst = 32'h38842800;
      49424: inst = 32'h10a00000;
      49425: inst = 32'hca0c115;
      49426: inst = 32'h13e00001;
      49427: inst = 32'hfe0d96a;
      49428: inst = 32'h5be00000;
      49429: inst = 32'h8c50000;
      49430: inst = 32'h24612800;
      49431: inst = 32'h10a0ffff;
      49432: inst = 32'hca0ffea;
      49433: inst = 32'h24822800;
      49434: inst = 32'h10a00000;
      49435: inst = 32'hca00004;
      49436: inst = 32'h38632800;
      49437: inst = 32'h38842800;
      49438: inst = 32'h10a00000;
      49439: inst = 32'hca0c123;
      49440: inst = 32'h13e00001;
      49441: inst = 32'hfe0d96a;
      49442: inst = 32'h5be00000;
      49443: inst = 32'h8c50000;
      49444: inst = 32'h24612800;
      49445: inst = 32'h10a0ffff;
      49446: inst = 32'hca0ffea;
      49447: inst = 32'h24822800;
      49448: inst = 32'h10a00000;
      49449: inst = 32'hca00004;
      49450: inst = 32'h38632800;
      49451: inst = 32'h38842800;
      49452: inst = 32'h10a00000;
      49453: inst = 32'hca0c131;
      49454: inst = 32'h13e00001;
      49455: inst = 32'hfe0d96a;
      49456: inst = 32'h5be00000;
      49457: inst = 32'h8c50000;
      49458: inst = 32'h24612800;
      49459: inst = 32'h10a0ffff;
      49460: inst = 32'hca0ffea;
      49461: inst = 32'h24822800;
      49462: inst = 32'h10a00000;
      49463: inst = 32'hca00004;
      49464: inst = 32'h38632800;
      49465: inst = 32'h38842800;
      49466: inst = 32'h10a00000;
      49467: inst = 32'hca0c13f;
      49468: inst = 32'h13e00001;
      49469: inst = 32'hfe0d96a;
      49470: inst = 32'h5be00000;
      49471: inst = 32'h8c50000;
      49472: inst = 32'h24612800;
      49473: inst = 32'h10a0ffff;
      49474: inst = 32'hca0ffea;
      49475: inst = 32'h24822800;
      49476: inst = 32'h10a00000;
      49477: inst = 32'hca00004;
      49478: inst = 32'h38632800;
      49479: inst = 32'h38842800;
      49480: inst = 32'h10a00000;
      49481: inst = 32'hca0c14d;
      49482: inst = 32'h13e00001;
      49483: inst = 32'hfe0d96a;
      49484: inst = 32'h5be00000;
      49485: inst = 32'h8c50000;
      49486: inst = 32'h24612800;
      49487: inst = 32'h10a0ffff;
      49488: inst = 32'hca0ffea;
      49489: inst = 32'h24822800;
      49490: inst = 32'h10a00000;
      49491: inst = 32'hca00004;
      49492: inst = 32'h38632800;
      49493: inst = 32'h38842800;
      49494: inst = 32'h10a00000;
      49495: inst = 32'hca0c15b;
      49496: inst = 32'h13e00001;
      49497: inst = 32'hfe0d96a;
      49498: inst = 32'h5be00000;
      49499: inst = 32'h8c50000;
      49500: inst = 32'h24612800;
      49501: inst = 32'h10a0ffff;
      49502: inst = 32'hca0ffea;
      49503: inst = 32'h24822800;
      49504: inst = 32'h10a00000;
      49505: inst = 32'hca00004;
      49506: inst = 32'h38632800;
      49507: inst = 32'h38842800;
      49508: inst = 32'h10a00000;
      49509: inst = 32'hca0c169;
      49510: inst = 32'h13e00001;
      49511: inst = 32'hfe0d96a;
      49512: inst = 32'h5be00000;
      49513: inst = 32'h8c50000;
      49514: inst = 32'h24612800;
      49515: inst = 32'h10a0ffff;
      49516: inst = 32'hca0ffea;
      49517: inst = 32'h24822800;
      49518: inst = 32'h10a00000;
      49519: inst = 32'hca00004;
      49520: inst = 32'h38632800;
      49521: inst = 32'h38842800;
      49522: inst = 32'h10a00000;
      49523: inst = 32'hca0c177;
      49524: inst = 32'h13e00001;
      49525: inst = 32'hfe0d96a;
      49526: inst = 32'h5be00000;
      49527: inst = 32'h8c50000;
      49528: inst = 32'h24612800;
      49529: inst = 32'h10a0ffff;
      49530: inst = 32'hca0ffea;
      49531: inst = 32'h24822800;
      49532: inst = 32'h10a00000;
      49533: inst = 32'hca00004;
      49534: inst = 32'h38632800;
      49535: inst = 32'h38842800;
      49536: inst = 32'h10a00000;
      49537: inst = 32'hca0c185;
      49538: inst = 32'h13e00001;
      49539: inst = 32'hfe0d96a;
      49540: inst = 32'h5be00000;
      49541: inst = 32'h8c50000;
      49542: inst = 32'h24612800;
      49543: inst = 32'h10a0ffff;
      49544: inst = 32'hca0ffea;
      49545: inst = 32'h24822800;
      49546: inst = 32'h10a00000;
      49547: inst = 32'hca00004;
      49548: inst = 32'h38632800;
      49549: inst = 32'h38842800;
      49550: inst = 32'h10a00000;
      49551: inst = 32'hca0c193;
      49552: inst = 32'h13e00001;
      49553: inst = 32'hfe0d96a;
      49554: inst = 32'h5be00000;
      49555: inst = 32'h8c50000;
      49556: inst = 32'h24612800;
      49557: inst = 32'h10a0ffff;
      49558: inst = 32'hca0ffea;
      49559: inst = 32'h24822800;
      49560: inst = 32'h10a00000;
      49561: inst = 32'hca00004;
      49562: inst = 32'h38632800;
      49563: inst = 32'h38842800;
      49564: inst = 32'h10a00000;
      49565: inst = 32'hca0c1a1;
      49566: inst = 32'h13e00001;
      49567: inst = 32'hfe0d96a;
      49568: inst = 32'h5be00000;
      49569: inst = 32'h8c50000;
      49570: inst = 32'h24612800;
      49571: inst = 32'h10a0ffff;
      49572: inst = 32'hca0ffea;
      49573: inst = 32'h24822800;
      49574: inst = 32'h10a00000;
      49575: inst = 32'hca00004;
      49576: inst = 32'h38632800;
      49577: inst = 32'h38842800;
      49578: inst = 32'h10a00000;
      49579: inst = 32'hca0c1af;
      49580: inst = 32'h13e00001;
      49581: inst = 32'hfe0d96a;
      49582: inst = 32'h5be00000;
      49583: inst = 32'h8c50000;
      49584: inst = 32'h24612800;
      49585: inst = 32'h10a0ffff;
      49586: inst = 32'hca0ffea;
      49587: inst = 32'h24822800;
      49588: inst = 32'h10a00000;
      49589: inst = 32'hca00004;
      49590: inst = 32'h38632800;
      49591: inst = 32'h38842800;
      49592: inst = 32'h10a00000;
      49593: inst = 32'hca0c1bd;
      49594: inst = 32'h13e00001;
      49595: inst = 32'hfe0d96a;
      49596: inst = 32'h5be00000;
      49597: inst = 32'h8c50000;
      49598: inst = 32'h24612800;
      49599: inst = 32'h10a0ffff;
      49600: inst = 32'hca0ffea;
      49601: inst = 32'h24822800;
      49602: inst = 32'h10a00000;
      49603: inst = 32'hca00004;
      49604: inst = 32'h38632800;
      49605: inst = 32'h38842800;
      49606: inst = 32'h10a00000;
      49607: inst = 32'hca0c1cb;
      49608: inst = 32'h13e00001;
      49609: inst = 32'hfe0d96a;
      49610: inst = 32'h5be00000;
      49611: inst = 32'h8c50000;
      49612: inst = 32'h24612800;
      49613: inst = 32'h10a0ffff;
      49614: inst = 32'hca0ffea;
      49615: inst = 32'h24822800;
      49616: inst = 32'h10a00000;
      49617: inst = 32'hca00004;
      49618: inst = 32'h38632800;
      49619: inst = 32'h38842800;
      49620: inst = 32'h10a00000;
      49621: inst = 32'hca0c1d9;
      49622: inst = 32'h13e00001;
      49623: inst = 32'hfe0d96a;
      49624: inst = 32'h5be00000;
      49625: inst = 32'h8c50000;
      49626: inst = 32'h24612800;
      49627: inst = 32'h10a0ffff;
      49628: inst = 32'hca0ffea;
      49629: inst = 32'h24822800;
      49630: inst = 32'h10a00000;
      49631: inst = 32'hca00004;
      49632: inst = 32'h38632800;
      49633: inst = 32'h38842800;
      49634: inst = 32'h10a00000;
      49635: inst = 32'hca0c1e7;
      49636: inst = 32'h13e00001;
      49637: inst = 32'hfe0d96a;
      49638: inst = 32'h5be00000;
      49639: inst = 32'h8c50000;
      49640: inst = 32'h24612800;
      49641: inst = 32'h10a0ffff;
      49642: inst = 32'hca0ffea;
      49643: inst = 32'h24822800;
      49644: inst = 32'h10a00000;
      49645: inst = 32'hca00004;
      49646: inst = 32'h38632800;
      49647: inst = 32'h38842800;
      49648: inst = 32'h10a00000;
      49649: inst = 32'hca0c1f5;
      49650: inst = 32'h13e00001;
      49651: inst = 32'hfe0d96a;
      49652: inst = 32'h5be00000;
      49653: inst = 32'h8c50000;
      49654: inst = 32'h24612800;
      49655: inst = 32'h10a0ffff;
      49656: inst = 32'hca0ffea;
      49657: inst = 32'h24822800;
      49658: inst = 32'h10a00000;
      49659: inst = 32'hca00004;
      49660: inst = 32'h38632800;
      49661: inst = 32'h38842800;
      49662: inst = 32'h10a00000;
      49663: inst = 32'hca0c203;
      49664: inst = 32'h13e00001;
      49665: inst = 32'hfe0d96a;
      49666: inst = 32'h5be00000;
      49667: inst = 32'h8c50000;
      49668: inst = 32'h24612800;
      49669: inst = 32'h10a0ffff;
      49670: inst = 32'hca0ffea;
      49671: inst = 32'h24822800;
      49672: inst = 32'h10a00000;
      49673: inst = 32'hca00004;
      49674: inst = 32'h38632800;
      49675: inst = 32'h38842800;
      49676: inst = 32'h10a00000;
      49677: inst = 32'hca0c211;
      49678: inst = 32'h13e00001;
      49679: inst = 32'hfe0d96a;
      49680: inst = 32'h5be00000;
      49681: inst = 32'h8c50000;
      49682: inst = 32'h24612800;
      49683: inst = 32'h10a0ffff;
      49684: inst = 32'hca0ffea;
      49685: inst = 32'h24822800;
      49686: inst = 32'h10a00000;
      49687: inst = 32'hca00004;
      49688: inst = 32'h38632800;
      49689: inst = 32'h38842800;
      49690: inst = 32'h10a00000;
      49691: inst = 32'hca0c21f;
      49692: inst = 32'h13e00001;
      49693: inst = 32'hfe0d96a;
      49694: inst = 32'h5be00000;
      49695: inst = 32'h8c50000;
      49696: inst = 32'h24612800;
      49697: inst = 32'h10a0ffff;
      49698: inst = 32'hca0ffea;
      49699: inst = 32'h24822800;
      49700: inst = 32'h10a00000;
      49701: inst = 32'hca00004;
      49702: inst = 32'h38632800;
      49703: inst = 32'h38842800;
      49704: inst = 32'h10a00000;
      49705: inst = 32'hca0c22d;
      49706: inst = 32'h13e00001;
      49707: inst = 32'hfe0d96a;
      49708: inst = 32'h5be00000;
      49709: inst = 32'h8c50000;
      49710: inst = 32'h24612800;
      49711: inst = 32'h10a0ffff;
      49712: inst = 32'hca0ffea;
      49713: inst = 32'h24822800;
      49714: inst = 32'h10a00000;
      49715: inst = 32'hca00004;
      49716: inst = 32'h38632800;
      49717: inst = 32'h38842800;
      49718: inst = 32'h10a00000;
      49719: inst = 32'hca0c23b;
      49720: inst = 32'h13e00001;
      49721: inst = 32'hfe0d96a;
      49722: inst = 32'h5be00000;
      49723: inst = 32'h8c50000;
      49724: inst = 32'h24612800;
      49725: inst = 32'h10a0ffff;
      49726: inst = 32'hca0ffea;
      49727: inst = 32'h24822800;
      49728: inst = 32'h10a00000;
      49729: inst = 32'hca00004;
      49730: inst = 32'h38632800;
      49731: inst = 32'h38842800;
      49732: inst = 32'h10a00000;
      49733: inst = 32'hca0c249;
      49734: inst = 32'h13e00001;
      49735: inst = 32'hfe0d96a;
      49736: inst = 32'h5be00000;
      49737: inst = 32'h8c50000;
      49738: inst = 32'h24612800;
      49739: inst = 32'h10a0ffff;
      49740: inst = 32'hca0ffea;
      49741: inst = 32'h24822800;
      49742: inst = 32'h10a00000;
      49743: inst = 32'hca00004;
      49744: inst = 32'h38632800;
      49745: inst = 32'h38842800;
      49746: inst = 32'h10a00000;
      49747: inst = 32'hca0c257;
      49748: inst = 32'h13e00001;
      49749: inst = 32'hfe0d96a;
      49750: inst = 32'h5be00000;
      49751: inst = 32'h8c50000;
      49752: inst = 32'h24612800;
      49753: inst = 32'h10a0ffff;
      49754: inst = 32'hca0ffea;
      49755: inst = 32'h24822800;
      49756: inst = 32'h10a00000;
      49757: inst = 32'hca00004;
      49758: inst = 32'h38632800;
      49759: inst = 32'h38842800;
      49760: inst = 32'h10a00000;
      49761: inst = 32'hca0c265;
      49762: inst = 32'h13e00001;
      49763: inst = 32'hfe0d96a;
      49764: inst = 32'h5be00000;
      49765: inst = 32'h8c50000;
      49766: inst = 32'h24612800;
      49767: inst = 32'h10a0ffff;
      49768: inst = 32'hca0ffea;
      49769: inst = 32'h24822800;
      49770: inst = 32'h10a00000;
      49771: inst = 32'hca00004;
      49772: inst = 32'h38632800;
      49773: inst = 32'h38842800;
      49774: inst = 32'h10a00000;
      49775: inst = 32'hca0c273;
      49776: inst = 32'h13e00001;
      49777: inst = 32'hfe0d96a;
      49778: inst = 32'h5be00000;
      49779: inst = 32'h8c50000;
      49780: inst = 32'h24612800;
      49781: inst = 32'h10a0ffff;
      49782: inst = 32'hca0ffea;
      49783: inst = 32'h24822800;
      49784: inst = 32'h10a00000;
      49785: inst = 32'hca00004;
      49786: inst = 32'h38632800;
      49787: inst = 32'h38842800;
      49788: inst = 32'h10a00000;
      49789: inst = 32'hca0c281;
      49790: inst = 32'h13e00001;
      49791: inst = 32'hfe0d96a;
      49792: inst = 32'h5be00000;
      49793: inst = 32'h8c50000;
      49794: inst = 32'h24612800;
      49795: inst = 32'h10a0ffff;
      49796: inst = 32'hca0ffea;
      49797: inst = 32'h24822800;
      49798: inst = 32'h10a00000;
      49799: inst = 32'hca00004;
      49800: inst = 32'h38632800;
      49801: inst = 32'h38842800;
      49802: inst = 32'h10a00000;
      49803: inst = 32'hca0c28f;
      49804: inst = 32'h13e00001;
      49805: inst = 32'hfe0d96a;
      49806: inst = 32'h5be00000;
      49807: inst = 32'h8c50000;
      49808: inst = 32'h24612800;
      49809: inst = 32'h10a0ffff;
      49810: inst = 32'hca0ffea;
      49811: inst = 32'h24822800;
      49812: inst = 32'h10a00000;
      49813: inst = 32'hca00004;
      49814: inst = 32'h38632800;
      49815: inst = 32'h38842800;
      49816: inst = 32'h10a00000;
      49817: inst = 32'hca0c29d;
      49818: inst = 32'h13e00001;
      49819: inst = 32'hfe0d96a;
      49820: inst = 32'h5be00000;
      49821: inst = 32'h8c50000;
      49822: inst = 32'h24612800;
      49823: inst = 32'h10a0ffff;
      49824: inst = 32'hca0ffea;
      49825: inst = 32'h24822800;
      49826: inst = 32'h10a00000;
      49827: inst = 32'hca00004;
      49828: inst = 32'h38632800;
      49829: inst = 32'h38842800;
      49830: inst = 32'h10a00000;
      49831: inst = 32'hca0c2ab;
      49832: inst = 32'h13e00001;
      49833: inst = 32'hfe0d96a;
      49834: inst = 32'h5be00000;
      49835: inst = 32'h8c50000;
      49836: inst = 32'h24612800;
      49837: inst = 32'h10a0ffff;
      49838: inst = 32'hca0ffea;
      49839: inst = 32'h24822800;
      49840: inst = 32'h10a00000;
      49841: inst = 32'hca00004;
      49842: inst = 32'h38632800;
      49843: inst = 32'h38842800;
      49844: inst = 32'h10a00000;
      49845: inst = 32'hca0c2b9;
      49846: inst = 32'h13e00001;
      49847: inst = 32'hfe0d96a;
      49848: inst = 32'h5be00000;
      49849: inst = 32'h8c50000;
      49850: inst = 32'h24612800;
      49851: inst = 32'h10a0ffff;
      49852: inst = 32'hca0ffea;
      49853: inst = 32'h24822800;
      49854: inst = 32'h10a00000;
      49855: inst = 32'hca00004;
      49856: inst = 32'h38632800;
      49857: inst = 32'h38842800;
      49858: inst = 32'h10a00000;
      49859: inst = 32'hca0c2c7;
      49860: inst = 32'h13e00001;
      49861: inst = 32'hfe0d96a;
      49862: inst = 32'h5be00000;
      49863: inst = 32'h8c50000;
      49864: inst = 32'h24612800;
      49865: inst = 32'h10a0ffff;
      49866: inst = 32'hca0ffea;
      49867: inst = 32'h24822800;
      49868: inst = 32'h10a00000;
      49869: inst = 32'hca00004;
      49870: inst = 32'h38632800;
      49871: inst = 32'h38842800;
      49872: inst = 32'h10a00000;
      49873: inst = 32'hca0c2d5;
      49874: inst = 32'h13e00001;
      49875: inst = 32'hfe0d96a;
      49876: inst = 32'h5be00000;
      49877: inst = 32'h8c50000;
      49878: inst = 32'h24612800;
      49879: inst = 32'h10a0ffff;
      49880: inst = 32'hca0ffea;
      49881: inst = 32'h24822800;
      49882: inst = 32'h10a00000;
      49883: inst = 32'hca00004;
      49884: inst = 32'h38632800;
      49885: inst = 32'h38842800;
      49886: inst = 32'h10a00000;
      49887: inst = 32'hca0c2e3;
      49888: inst = 32'h13e00001;
      49889: inst = 32'hfe0d96a;
      49890: inst = 32'h5be00000;
      49891: inst = 32'h8c50000;
      49892: inst = 32'h24612800;
      49893: inst = 32'h10a0ffff;
      49894: inst = 32'hca0ffea;
      49895: inst = 32'h24822800;
      49896: inst = 32'h10a00000;
      49897: inst = 32'hca00004;
      49898: inst = 32'h38632800;
      49899: inst = 32'h38842800;
      49900: inst = 32'h10a00000;
      49901: inst = 32'hca0c2f1;
      49902: inst = 32'h13e00001;
      49903: inst = 32'hfe0d96a;
      49904: inst = 32'h5be00000;
      49905: inst = 32'h8c50000;
      49906: inst = 32'h24612800;
      49907: inst = 32'h10a0ffff;
      49908: inst = 32'hca0ffea;
      49909: inst = 32'h24822800;
      49910: inst = 32'h10a00000;
      49911: inst = 32'hca00004;
      49912: inst = 32'h38632800;
      49913: inst = 32'h38842800;
      49914: inst = 32'h10a00000;
      49915: inst = 32'hca0c2ff;
      49916: inst = 32'h13e00001;
      49917: inst = 32'hfe0d96a;
      49918: inst = 32'h5be00000;
      49919: inst = 32'h8c50000;
      49920: inst = 32'h24612800;
      49921: inst = 32'h10a0ffff;
      49922: inst = 32'hca0ffea;
      49923: inst = 32'h24822800;
      49924: inst = 32'h10a00000;
      49925: inst = 32'hca00004;
      49926: inst = 32'h38632800;
      49927: inst = 32'h38842800;
      49928: inst = 32'h10a00000;
      49929: inst = 32'hca0c30d;
      49930: inst = 32'h13e00001;
      49931: inst = 32'hfe0d96a;
      49932: inst = 32'h5be00000;
      49933: inst = 32'h8c50000;
      49934: inst = 32'h24612800;
      49935: inst = 32'h10a0ffff;
      49936: inst = 32'hca0ffea;
      49937: inst = 32'h24822800;
      49938: inst = 32'h10a00000;
      49939: inst = 32'hca00004;
      49940: inst = 32'h38632800;
      49941: inst = 32'h38842800;
      49942: inst = 32'h10a00000;
      49943: inst = 32'hca0c31b;
      49944: inst = 32'h13e00001;
      49945: inst = 32'hfe0d96a;
      49946: inst = 32'h5be00000;
      49947: inst = 32'h8c50000;
      49948: inst = 32'h24612800;
      49949: inst = 32'h10a0ffff;
      49950: inst = 32'hca0ffea;
      49951: inst = 32'h24822800;
      49952: inst = 32'h10a00000;
      49953: inst = 32'hca00004;
      49954: inst = 32'h38632800;
      49955: inst = 32'h38842800;
      49956: inst = 32'h10a00000;
      49957: inst = 32'hca0c329;
      49958: inst = 32'h13e00001;
      49959: inst = 32'hfe0d96a;
      49960: inst = 32'h5be00000;
      49961: inst = 32'h8c50000;
      49962: inst = 32'h24612800;
      49963: inst = 32'h10a0ffff;
      49964: inst = 32'hca0ffeb;
      49965: inst = 32'h24822800;
      49966: inst = 32'h10a00000;
      49967: inst = 32'hca00004;
      49968: inst = 32'h38632800;
      49969: inst = 32'h38842800;
      49970: inst = 32'h10a00000;
      49971: inst = 32'hca0c337;
      49972: inst = 32'h13e00001;
      49973: inst = 32'hfe0d96a;
      49974: inst = 32'h5be00000;
      49975: inst = 32'h8c50000;
      49976: inst = 32'h24612800;
      49977: inst = 32'h10a0ffff;
      49978: inst = 32'hca0ffeb;
      49979: inst = 32'h24822800;
      49980: inst = 32'h10a00000;
      49981: inst = 32'hca00004;
      49982: inst = 32'h38632800;
      49983: inst = 32'h38842800;
      49984: inst = 32'h10a00000;
      49985: inst = 32'hca0c345;
      49986: inst = 32'h13e00001;
      49987: inst = 32'hfe0d96a;
      49988: inst = 32'h5be00000;
      49989: inst = 32'h8c50000;
      49990: inst = 32'h24612800;
      49991: inst = 32'h10a0ffff;
      49992: inst = 32'hca0ffeb;
      49993: inst = 32'h24822800;
      49994: inst = 32'h10a00000;
      49995: inst = 32'hca00004;
      49996: inst = 32'h38632800;
      49997: inst = 32'h38842800;
      49998: inst = 32'h10a00000;
      49999: inst = 32'hca0c353;
      50000: inst = 32'h13e00001;
      50001: inst = 32'hfe0d96a;
      50002: inst = 32'h5be00000;
      50003: inst = 32'h8c50000;
      50004: inst = 32'h24612800;
      50005: inst = 32'h10a0ffff;
      50006: inst = 32'hca0ffeb;
      50007: inst = 32'h24822800;
      50008: inst = 32'h10a00000;
      50009: inst = 32'hca00004;
      50010: inst = 32'h38632800;
      50011: inst = 32'h38842800;
      50012: inst = 32'h10a00000;
      50013: inst = 32'hca0c361;
      50014: inst = 32'h13e00001;
      50015: inst = 32'hfe0d96a;
      50016: inst = 32'h5be00000;
      50017: inst = 32'h8c50000;
      50018: inst = 32'h24612800;
      50019: inst = 32'h10a0ffff;
      50020: inst = 32'hca0ffeb;
      50021: inst = 32'h24822800;
      50022: inst = 32'h10a00000;
      50023: inst = 32'hca00004;
      50024: inst = 32'h38632800;
      50025: inst = 32'h38842800;
      50026: inst = 32'h10a00000;
      50027: inst = 32'hca0c36f;
      50028: inst = 32'h13e00001;
      50029: inst = 32'hfe0d96a;
      50030: inst = 32'h5be00000;
      50031: inst = 32'h8c50000;
      50032: inst = 32'h24612800;
      50033: inst = 32'h10a0ffff;
      50034: inst = 32'hca0ffeb;
      50035: inst = 32'h24822800;
      50036: inst = 32'h10a00000;
      50037: inst = 32'hca00004;
      50038: inst = 32'h38632800;
      50039: inst = 32'h38842800;
      50040: inst = 32'h10a00000;
      50041: inst = 32'hca0c37d;
      50042: inst = 32'h13e00001;
      50043: inst = 32'hfe0d96a;
      50044: inst = 32'h5be00000;
      50045: inst = 32'h8c50000;
      50046: inst = 32'h24612800;
      50047: inst = 32'h10a0ffff;
      50048: inst = 32'hca0ffeb;
      50049: inst = 32'h24822800;
      50050: inst = 32'h10a00000;
      50051: inst = 32'hca00004;
      50052: inst = 32'h38632800;
      50053: inst = 32'h38842800;
      50054: inst = 32'h10a00000;
      50055: inst = 32'hca0c38b;
      50056: inst = 32'h13e00001;
      50057: inst = 32'hfe0d96a;
      50058: inst = 32'h5be00000;
      50059: inst = 32'h8c50000;
      50060: inst = 32'h24612800;
      50061: inst = 32'h10a0ffff;
      50062: inst = 32'hca0ffeb;
      50063: inst = 32'h24822800;
      50064: inst = 32'h10a00000;
      50065: inst = 32'hca00004;
      50066: inst = 32'h38632800;
      50067: inst = 32'h38842800;
      50068: inst = 32'h10a00000;
      50069: inst = 32'hca0c399;
      50070: inst = 32'h13e00001;
      50071: inst = 32'hfe0d96a;
      50072: inst = 32'h5be00000;
      50073: inst = 32'h8c50000;
      50074: inst = 32'h24612800;
      50075: inst = 32'h10a0ffff;
      50076: inst = 32'hca0ffeb;
      50077: inst = 32'h24822800;
      50078: inst = 32'h10a00000;
      50079: inst = 32'hca00004;
      50080: inst = 32'h38632800;
      50081: inst = 32'h38842800;
      50082: inst = 32'h10a00000;
      50083: inst = 32'hca0c3a7;
      50084: inst = 32'h13e00001;
      50085: inst = 32'hfe0d96a;
      50086: inst = 32'h5be00000;
      50087: inst = 32'h8c50000;
      50088: inst = 32'h24612800;
      50089: inst = 32'h10a0ffff;
      50090: inst = 32'hca0ffeb;
      50091: inst = 32'h24822800;
      50092: inst = 32'h10a00000;
      50093: inst = 32'hca00004;
      50094: inst = 32'h38632800;
      50095: inst = 32'h38842800;
      50096: inst = 32'h10a00000;
      50097: inst = 32'hca0c3b5;
      50098: inst = 32'h13e00001;
      50099: inst = 32'hfe0d96a;
      50100: inst = 32'h5be00000;
      50101: inst = 32'h8c50000;
      50102: inst = 32'h24612800;
      50103: inst = 32'h10a0ffff;
      50104: inst = 32'hca0ffeb;
      50105: inst = 32'h24822800;
      50106: inst = 32'h10a00000;
      50107: inst = 32'hca00004;
      50108: inst = 32'h38632800;
      50109: inst = 32'h38842800;
      50110: inst = 32'h10a00000;
      50111: inst = 32'hca0c3c3;
      50112: inst = 32'h13e00001;
      50113: inst = 32'hfe0d96a;
      50114: inst = 32'h5be00000;
      50115: inst = 32'h8c50000;
      50116: inst = 32'h24612800;
      50117: inst = 32'h10a0ffff;
      50118: inst = 32'hca0ffeb;
      50119: inst = 32'h24822800;
      50120: inst = 32'h10a00000;
      50121: inst = 32'hca00004;
      50122: inst = 32'h38632800;
      50123: inst = 32'h38842800;
      50124: inst = 32'h10a00000;
      50125: inst = 32'hca0c3d1;
      50126: inst = 32'h13e00001;
      50127: inst = 32'hfe0d96a;
      50128: inst = 32'h5be00000;
      50129: inst = 32'h8c50000;
      50130: inst = 32'h24612800;
      50131: inst = 32'h10a0ffff;
      50132: inst = 32'hca0ffeb;
      50133: inst = 32'h24822800;
      50134: inst = 32'h10a00000;
      50135: inst = 32'hca00004;
      50136: inst = 32'h38632800;
      50137: inst = 32'h38842800;
      50138: inst = 32'h10a00000;
      50139: inst = 32'hca0c3df;
      50140: inst = 32'h13e00001;
      50141: inst = 32'hfe0d96a;
      50142: inst = 32'h5be00000;
      50143: inst = 32'h8c50000;
      50144: inst = 32'h24612800;
      50145: inst = 32'h10a0ffff;
      50146: inst = 32'hca0ffeb;
      50147: inst = 32'h24822800;
      50148: inst = 32'h10a00000;
      50149: inst = 32'hca00004;
      50150: inst = 32'h38632800;
      50151: inst = 32'h38842800;
      50152: inst = 32'h10a00000;
      50153: inst = 32'hca0c3ed;
      50154: inst = 32'h13e00001;
      50155: inst = 32'hfe0d96a;
      50156: inst = 32'h5be00000;
      50157: inst = 32'h8c50000;
      50158: inst = 32'h24612800;
      50159: inst = 32'h10a0ffff;
      50160: inst = 32'hca0ffeb;
      50161: inst = 32'h24822800;
      50162: inst = 32'h10a00000;
      50163: inst = 32'hca00004;
      50164: inst = 32'h38632800;
      50165: inst = 32'h38842800;
      50166: inst = 32'h10a00000;
      50167: inst = 32'hca0c3fb;
      50168: inst = 32'h13e00001;
      50169: inst = 32'hfe0d96a;
      50170: inst = 32'h5be00000;
      50171: inst = 32'h8c50000;
      50172: inst = 32'h24612800;
      50173: inst = 32'h10a0ffff;
      50174: inst = 32'hca0ffeb;
      50175: inst = 32'h24822800;
      50176: inst = 32'h10a00000;
      50177: inst = 32'hca00004;
      50178: inst = 32'h38632800;
      50179: inst = 32'h38842800;
      50180: inst = 32'h10a00000;
      50181: inst = 32'hca0c409;
      50182: inst = 32'h13e00001;
      50183: inst = 32'hfe0d96a;
      50184: inst = 32'h5be00000;
      50185: inst = 32'h8c50000;
      50186: inst = 32'h24612800;
      50187: inst = 32'h10a0ffff;
      50188: inst = 32'hca0ffeb;
      50189: inst = 32'h24822800;
      50190: inst = 32'h10a00000;
      50191: inst = 32'hca00004;
      50192: inst = 32'h38632800;
      50193: inst = 32'h38842800;
      50194: inst = 32'h10a00000;
      50195: inst = 32'hca0c417;
      50196: inst = 32'h13e00001;
      50197: inst = 32'hfe0d96a;
      50198: inst = 32'h5be00000;
      50199: inst = 32'h8c50000;
      50200: inst = 32'h24612800;
      50201: inst = 32'h10a0ffff;
      50202: inst = 32'hca0ffeb;
      50203: inst = 32'h24822800;
      50204: inst = 32'h10a00000;
      50205: inst = 32'hca00004;
      50206: inst = 32'h38632800;
      50207: inst = 32'h38842800;
      50208: inst = 32'h10a00000;
      50209: inst = 32'hca0c425;
      50210: inst = 32'h13e00001;
      50211: inst = 32'hfe0d96a;
      50212: inst = 32'h5be00000;
      50213: inst = 32'h8c50000;
      50214: inst = 32'h24612800;
      50215: inst = 32'h10a0ffff;
      50216: inst = 32'hca0ffeb;
      50217: inst = 32'h24822800;
      50218: inst = 32'h10a00000;
      50219: inst = 32'hca00004;
      50220: inst = 32'h38632800;
      50221: inst = 32'h38842800;
      50222: inst = 32'h10a00000;
      50223: inst = 32'hca0c433;
      50224: inst = 32'h13e00001;
      50225: inst = 32'hfe0d96a;
      50226: inst = 32'h5be00000;
      50227: inst = 32'h8c50000;
      50228: inst = 32'h24612800;
      50229: inst = 32'h10a0ffff;
      50230: inst = 32'hca0ffeb;
      50231: inst = 32'h24822800;
      50232: inst = 32'h10a00000;
      50233: inst = 32'hca00004;
      50234: inst = 32'h38632800;
      50235: inst = 32'h38842800;
      50236: inst = 32'h10a00000;
      50237: inst = 32'hca0c441;
      50238: inst = 32'h13e00001;
      50239: inst = 32'hfe0d96a;
      50240: inst = 32'h5be00000;
      50241: inst = 32'h8c50000;
      50242: inst = 32'h24612800;
      50243: inst = 32'h10a0ffff;
      50244: inst = 32'hca0ffeb;
      50245: inst = 32'h24822800;
      50246: inst = 32'h10a00000;
      50247: inst = 32'hca00004;
      50248: inst = 32'h38632800;
      50249: inst = 32'h38842800;
      50250: inst = 32'h10a00000;
      50251: inst = 32'hca0c44f;
      50252: inst = 32'h13e00001;
      50253: inst = 32'hfe0d96a;
      50254: inst = 32'h5be00000;
      50255: inst = 32'h8c50000;
      50256: inst = 32'h24612800;
      50257: inst = 32'h10a0ffff;
      50258: inst = 32'hca0ffeb;
      50259: inst = 32'h24822800;
      50260: inst = 32'h10a00000;
      50261: inst = 32'hca00004;
      50262: inst = 32'h38632800;
      50263: inst = 32'h38842800;
      50264: inst = 32'h10a00000;
      50265: inst = 32'hca0c45d;
      50266: inst = 32'h13e00001;
      50267: inst = 32'hfe0d96a;
      50268: inst = 32'h5be00000;
      50269: inst = 32'h8c50000;
      50270: inst = 32'h24612800;
      50271: inst = 32'h10a0ffff;
      50272: inst = 32'hca0ffeb;
      50273: inst = 32'h24822800;
      50274: inst = 32'h10a00000;
      50275: inst = 32'hca00004;
      50276: inst = 32'h38632800;
      50277: inst = 32'h38842800;
      50278: inst = 32'h10a00000;
      50279: inst = 32'hca0c46b;
      50280: inst = 32'h13e00001;
      50281: inst = 32'hfe0d96a;
      50282: inst = 32'h5be00000;
      50283: inst = 32'h8c50000;
      50284: inst = 32'h24612800;
      50285: inst = 32'h10a0ffff;
      50286: inst = 32'hca0ffeb;
      50287: inst = 32'h24822800;
      50288: inst = 32'h10a00000;
      50289: inst = 32'hca00004;
      50290: inst = 32'h38632800;
      50291: inst = 32'h38842800;
      50292: inst = 32'h10a00000;
      50293: inst = 32'hca0c479;
      50294: inst = 32'h13e00001;
      50295: inst = 32'hfe0d96a;
      50296: inst = 32'h5be00000;
      50297: inst = 32'h8c50000;
      50298: inst = 32'h24612800;
      50299: inst = 32'h10a0ffff;
      50300: inst = 32'hca0ffeb;
      50301: inst = 32'h24822800;
      50302: inst = 32'h10a00000;
      50303: inst = 32'hca00004;
      50304: inst = 32'h38632800;
      50305: inst = 32'h38842800;
      50306: inst = 32'h10a00000;
      50307: inst = 32'hca0c487;
      50308: inst = 32'h13e00001;
      50309: inst = 32'hfe0d96a;
      50310: inst = 32'h5be00000;
      50311: inst = 32'h8c50000;
      50312: inst = 32'h24612800;
      50313: inst = 32'h10a0ffff;
      50314: inst = 32'hca0ffeb;
      50315: inst = 32'h24822800;
      50316: inst = 32'h10a00000;
      50317: inst = 32'hca00004;
      50318: inst = 32'h38632800;
      50319: inst = 32'h38842800;
      50320: inst = 32'h10a00000;
      50321: inst = 32'hca0c495;
      50322: inst = 32'h13e00001;
      50323: inst = 32'hfe0d96a;
      50324: inst = 32'h5be00000;
      50325: inst = 32'h8c50000;
      50326: inst = 32'h24612800;
      50327: inst = 32'h10a0ffff;
      50328: inst = 32'hca0ffeb;
      50329: inst = 32'h24822800;
      50330: inst = 32'h10a00000;
      50331: inst = 32'hca00004;
      50332: inst = 32'h38632800;
      50333: inst = 32'h38842800;
      50334: inst = 32'h10a00000;
      50335: inst = 32'hca0c4a3;
      50336: inst = 32'h13e00001;
      50337: inst = 32'hfe0d96a;
      50338: inst = 32'h5be00000;
      50339: inst = 32'h8c50000;
      50340: inst = 32'h24612800;
      50341: inst = 32'h10a0ffff;
      50342: inst = 32'hca0ffeb;
      50343: inst = 32'h24822800;
      50344: inst = 32'h10a00000;
      50345: inst = 32'hca00004;
      50346: inst = 32'h38632800;
      50347: inst = 32'h38842800;
      50348: inst = 32'h10a00000;
      50349: inst = 32'hca0c4b1;
      50350: inst = 32'h13e00001;
      50351: inst = 32'hfe0d96a;
      50352: inst = 32'h5be00000;
      50353: inst = 32'h8c50000;
      50354: inst = 32'h24612800;
      50355: inst = 32'h10a0ffff;
      50356: inst = 32'hca0ffeb;
      50357: inst = 32'h24822800;
      50358: inst = 32'h10a00000;
      50359: inst = 32'hca00004;
      50360: inst = 32'h38632800;
      50361: inst = 32'h38842800;
      50362: inst = 32'h10a00000;
      50363: inst = 32'hca0c4bf;
      50364: inst = 32'h13e00001;
      50365: inst = 32'hfe0d96a;
      50366: inst = 32'h5be00000;
      50367: inst = 32'h8c50000;
      50368: inst = 32'h24612800;
      50369: inst = 32'h10a0ffff;
      50370: inst = 32'hca0ffeb;
      50371: inst = 32'h24822800;
      50372: inst = 32'h10a00000;
      50373: inst = 32'hca00004;
      50374: inst = 32'h38632800;
      50375: inst = 32'h38842800;
      50376: inst = 32'h10a00000;
      50377: inst = 32'hca0c4cd;
      50378: inst = 32'h13e00001;
      50379: inst = 32'hfe0d96a;
      50380: inst = 32'h5be00000;
      50381: inst = 32'h8c50000;
      50382: inst = 32'h24612800;
      50383: inst = 32'h10a0ffff;
      50384: inst = 32'hca0ffeb;
      50385: inst = 32'h24822800;
      50386: inst = 32'h10a00000;
      50387: inst = 32'hca00004;
      50388: inst = 32'h38632800;
      50389: inst = 32'h38842800;
      50390: inst = 32'h10a00000;
      50391: inst = 32'hca0c4db;
      50392: inst = 32'h13e00001;
      50393: inst = 32'hfe0d96a;
      50394: inst = 32'h5be00000;
      50395: inst = 32'h8c50000;
      50396: inst = 32'h24612800;
      50397: inst = 32'h10a0ffff;
      50398: inst = 32'hca0ffeb;
      50399: inst = 32'h24822800;
      50400: inst = 32'h10a00000;
      50401: inst = 32'hca00004;
      50402: inst = 32'h38632800;
      50403: inst = 32'h38842800;
      50404: inst = 32'h10a00000;
      50405: inst = 32'hca0c4e9;
      50406: inst = 32'h13e00001;
      50407: inst = 32'hfe0d96a;
      50408: inst = 32'h5be00000;
      50409: inst = 32'h8c50000;
      50410: inst = 32'h24612800;
      50411: inst = 32'h10a0ffff;
      50412: inst = 32'hca0ffeb;
      50413: inst = 32'h24822800;
      50414: inst = 32'h10a00000;
      50415: inst = 32'hca00004;
      50416: inst = 32'h38632800;
      50417: inst = 32'h38842800;
      50418: inst = 32'h10a00000;
      50419: inst = 32'hca0c4f7;
      50420: inst = 32'h13e00001;
      50421: inst = 32'hfe0d96a;
      50422: inst = 32'h5be00000;
      50423: inst = 32'h8c50000;
      50424: inst = 32'h24612800;
      50425: inst = 32'h10a0ffff;
      50426: inst = 32'hca0ffeb;
      50427: inst = 32'h24822800;
      50428: inst = 32'h10a00000;
      50429: inst = 32'hca00004;
      50430: inst = 32'h38632800;
      50431: inst = 32'h38842800;
      50432: inst = 32'h10a00000;
      50433: inst = 32'hca0c505;
      50434: inst = 32'h13e00001;
      50435: inst = 32'hfe0d96a;
      50436: inst = 32'h5be00000;
      50437: inst = 32'h8c50000;
      50438: inst = 32'h24612800;
      50439: inst = 32'h10a0ffff;
      50440: inst = 32'hca0ffeb;
      50441: inst = 32'h24822800;
      50442: inst = 32'h10a00000;
      50443: inst = 32'hca00004;
      50444: inst = 32'h38632800;
      50445: inst = 32'h38842800;
      50446: inst = 32'h10a00000;
      50447: inst = 32'hca0c513;
      50448: inst = 32'h13e00001;
      50449: inst = 32'hfe0d96a;
      50450: inst = 32'h5be00000;
      50451: inst = 32'h8c50000;
      50452: inst = 32'h24612800;
      50453: inst = 32'h10a0ffff;
      50454: inst = 32'hca0ffeb;
      50455: inst = 32'h24822800;
      50456: inst = 32'h10a00000;
      50457: inst = 32'hca00004;
      50458: inst = 32'h38632800;
      50459: inst = 32'h38842800;
      50460: inst = 32'h10a00000;
      50461: inst = 32'hca0c521;
      50462: inst = 32'h13e00001;
      50463: inst = 32'hfe0d96a;
      50464: inst = 32'h5be00000;
      50465: inst = 32'h8c50000;
      50466: inst = 32'h24612800;
      50467: inst = 32'h10a0ffff;
      50468: inst = 32'hca0ffeb;
      50469: inst = 32'h24822800;
      50470: inst = 32'h10a00000;
      50471: inst = 32'hca00004;
      50472: inst = 32'h38632800;
      50473: inst = 32'h38842800;
      50474: inst = 32'h10a00000;
      50475: inst = 32'hca0c52f;
      50476: inst = 32'h13e00001;
      50477: inst = 32'hfe0d96a;
      50478: inst = 32'h5be00000;
      50479: inst = 32'h8c50000;
      50480: inst = 32'h24612800;
      50481: inst = 32'h10a0ffff;
      50482: inst = 32'hca0ffeb;
      50483: inst = 32'h24822800;
      50484: inst = 32'h10a00000;
      50485: inst = 32'hca00004;
      50486: inst = 32'h38632800;
      50487: inst = 32'h38842800;
      50488: inst = 32'h10a00000;
      50489: inst = 32'hca0c53d;
      50490: inst = 32'h13e00001;
      50491: inst = 32'hfe0d96a;
      50492: inst = 32'h5be00000;
      50493: inst = 32'h8c50000;
      50494: inst = 32'h24612800;
      50495: inst = 32'h10a0ffff;
      50496: inst = 32'hca0ffeb;
      50497: inst = 32'h24822800;
      50498: inst = 32'h10a00000;
      50499: inst = 32'hca00004;
      50500: inst = 32'h38632800;
      50501: inst = 32'h38842800;
      50502: inst = 32'h10a00000;
      50503: inst = 32'hca0c54b;
      50504: inst = 32'h13e00001;
      50505: inst = 32'hfe0d96a;
      50506: inst = 32'h5be00000;
      50507: inst = 32'h8c50000;
      50508: inst = 32'h24612800;
      50509: inst = 32'h10a0ffff;
      50510: inst = 32'hca0ffeb;
      50511: inst = 32'h24822800;
      50512: inst = 32'h10a00000;
      50513: inst = 32'hca00004;
      50514: inst = 32'h38632800;
      50515: inst = 32'h38842800;
      50516: inst = 32'h10a00000;
      50517: inst = 32'hca0c559;
      50518: inst = 32'h13e00001;
      50519: inst = 32'hfe0d96a;
      50520: inst = 32'h5be00000;
      50521: inst = 32'h8c50000;
      50522: inst = 32'h24612800;
      50523: inst = 32'h10a0ffff;
      50524: inst = 32'hca0ffeb;
      50525: inst = 32'h24822800;
      50526: inst = 32'h10a00000;
      50527: inst = 32'hca00004;
      50528: inst = 32'h38632800;
      50529: inst = 32'h38842800;
      50530: inst = 32'h10a00000;
      50531: inst = 32'hca0c567;
      50532: inst = 32'h13e00001;
      50533: inst = 32'hfe0d96a;
      50534: inst = 32'h5be00000;
      50535: inst = 32'h8c50000;
      50536: inst = 32'h24612800;
      50537: inst = 32'h10a0ffff;
      50538: inst = 32'hca0ffeb;
      50539: inst = 32'h24822800;
      50540: inst = 32'h10a00000;
      50541: inst = 32'hca00004;
      50542: inst = 32'h38632800;
      50543: inst = 32'h38842800;
      50544: inst = 32'h10a00000;
      50545: inst = 32'hca0c575;
      50546: inst = 32'h13e00001;
      50547: inst = 32'hfe0d96a;
      50548: inst = 32'h5be00000;
      50549: inst = 32'h8c50000;
      50550: inst = 32'h24612800;
      50551: inst = 32'h10a0ffff;
      50552: inst = 32'hca0ffeb;
      50553: inst = 32'h24822800;
      50554: inst = 32'h10a00000;
      50555: inst = 32'hca00004;
      50556: inst = 32'h38632800;
      50557: inst = 32'h38842800;
      50558: inst = 32'h10a00000;
      50559: inst = 32'hca0c583;
      50560: inst = 32'h13e00001;
      50561: inst = 32'hfe0d96a;
      50562: inst = 32'h5be00000;
      50563: inst = 32'h8c50000;
      50564: inst = 32'h24612800;
      50565: inst = 32'h10a0ffff;
      50566: inst = 32'hca0ffeb;
      50567: inst = 32'h24822800;
      50568: inst = 32'h10a00000;
      50569: inst = 32'hca00004;
      50570: inst = 32'h38632800;
      50571: inst = 32'h38842800;
      50572: inst = 32'h10a00000;
      50573: inst = 32'hca0c591;
      50574: inst = 32'h13e00001;
      50575: inst = 32'hfe0d96a;
      50576: inst = 32'h5be00000;
      50577: inst = 32'h8c50000;
      50578: inst = 32'h24612800;
      50579: inst = 32'h10a0ffff;
      50580: inst = 32'hca0ffeb;
      50581: inst = 32'h24822800;
      50582: inst = 32'h10a00000;
      50583: inst = 32'hca00004;
      50584: inst = 32'h38632800;
      50585: inst = 32'h38842800;
      50586: inst = 32'h10a00000;
      50587: inst = 32'hca0c59f;
      50588: inst = 32'h13e00001;
      50589: inst = 32'hfe0d96a;
      50590: inst = 32'h5be00000;
      50591: inst = 32'h8c50000;
      50592: inst = 32'h24612800;
      50593: inst = 32'h10a0ffff;
      50594: inst = 32'hca0ffeb;
      50595: inst = 32'h24822800;
      50596: inst = 32'h10a00000;
      50597: inst = 32'hca00004;
      50598: inst = 32'h38632800;
      50599: inst = 32'h38842800;
      50600: inst = 32'h10a00000;
      50601: inst = 32'hca0c5ad;
      50602: inst = 32'h13e00001;
      50603: inst = 32'hfe0d96a;
      50604: inst = 32'h5be00000;
      50605: inst = 32'h8c50000;
      50606: inst = 32'h24612800;
      50607: inst = 32'h10a0ffff;
      50608: inst = 32'hca0ffeb;
      50609: inst = 32'h24822800;
      50610: inst = 32'h10a00000;
      50611: inst = 32'hca00004;
      50612: inst = 32'h38632800;
      50613: inst = 32'h38842800;
      50614: inst = 32'h10a00000;
      50615: inst = 32'hca0c5bb;
      50616: inst = 32'h13e00001;
      50617: inst = 32'hfe0d96a;
      50618: inst = 32'h5be00000;
      50619: inst = 32'h8c50000;
      50620: inst = 32'h24612800;
      50621: inst = 32'h10a0ffff;
      50622: inst = 32'hca0ffeb;
      50623: inst = 32'h24822800;
      50624: inst = 32'h10a00000;
      50625: inst = 32'hca00004;
      50626: inst = 32'h38632800;
      50627: inst = 32'h38842800;
      50628: inst = 32'h10a00000;
      50629: inst = 32'hca0c5c9;
      50630: inst = 32'h13e00001;
      50631: inst = 32'hfe0d96a;
      50632: inst = 32'h5be00000;
      50633: inst = 32'h8c50000;
      50634: inst = 32'h24612800;
      50635: inst = 32'h10a0ffff;
      50636: inst = 32'hca0ffeb;
      50637: inst = 32'h24822800;
      50638: inst = 32'h10a00000;
      50639: inst = 32'hca00004;
      50640: inst = 32'h38632800;
      50641: inst = 32'h38842800;
      50642: inst = 32'h10a00000;
      50643: inst = 32'hca0c5d7;
      50644: inst = 32'h13e00001;
      50645: inst = 32'hfe0d96a;
      50646: inst = 32'h5be00000;
      50647: inst = 32'h8c50000;
      50648: inst = 32'h24612800;
      50649: inst = 32'h10a0ffff;
      50650: inst = 32'hca0ffeb;
      50651: inst = 32'h24822800;
      50652: inst = 32'h10a00000;
      50653: inst = 32'hca00004;
      50654: inst = 32'h38632800;
      50655: inst = 32'h38842800;
      50656: inst = 32'h10a00000;
      50657: inst = 32'hca0c5e5;
      50658: inst = 32'h13e00001;
      50659: inst = 32'hfe0d96a;
      50660: inst = 32'h5be00000;
      50661: inst = 32'h8c50000;
      50662: inst = 32'h24612800;
      50663: inst = 32'h10a0ffff;
      50664: inst = 32'hca0ffeb;
      50665: inst = 32'h24822800;
      50666: inst = 32'h10a00000;
      50667: inst = 32'hca00004;
      50668: inst = 32'h38632800;
      50669: inst = 32'h38842800;
      50670: inst = 32'h10a00000;
      50671: inst = 32'hca0c5f3;
      50672: inst = 32'h13e00001;
      50673: inst = 32'hfe0d96a;
      50674: inst = 32'h5be00000;
      50675: inst = 32'h8c50000;
      50676: inst = 32'h24612800;
      50677: inst = 32'h10a0ffff;
      50678: inst = 32'hca0ffeb;
      50679: inst = 32'h24822800;
      50680: inst = 32'h10a00000;
      50681: inst = 32'hca00004;
      50682: inst = 32'h38632800;
      50683: inst = 32'h38842800;
      50684: inst = 32'h10a00000;
      50685: inst = 32'hca0c601;
      50686: inst = 32'h13e00001;
      50687: inst = 32'hfe0d96a;
      50688: inst = 32'h5be00000;
      50689: inst = 32'h8c50000;
      50690: inst = 32'h24612800;
      50691: inst = 32'h10a0ffff;
      50692: inst = 32'hca0ffeb;
      50693: inst = 32'h24822800;
      50694: inst = 32'h10a00000;
      50695: inst = 32'hca00004;
      50696: inst = 32'h38632800;
      50697: inst = 32'h38842800;
      50698: inst = 32'h10a00000;
      50699: inst = 32'hca0c60f;
      50700: inst = 32'h13e00001;
      50701: inst = 32'hfe0d96a;
      50702: inst = 32'h5be00000;
      50703: inst = 32'h8c50000;
      50704: inst = 32'h24612800;
      50705: inst = 32'h10a0ffff;
      50706: inst = 32'hca0ffeb;
      50707: inst = 32'h24822800;
      50708: inst = 32'h10a00000;
      50709: inst = 32'hca00004;
      50710: inst = 32'h38632800;
      50711: inst = 32'h38842800;
      50712: inst = 32'h10a00000;
      50713: inst = 32'hca0c61d;
      50714: inst = 32'h13e00001;
      50715: inst = 32'hfe0d96a;
      50716: inst = 32'h5be00000;
      50717: inst = 32'h8c50000;
      50718: inst = 32'h24612800;
      50719: inst = 32'h10a0ffff;
      50720: inst = 32'hca0ffeb;
      50721: inst = 32'h24822800;
      50722: inst = 32'h10a00000;
      50723: inst = 32'hca00004;
      50724: inst = 32'h38632800;
      50725: inst = 32'h38842800;
      50726: inst = 32'h10a00000;
      50727: inst = 32'hca0c62b;
      50728: inst = 32'h13e00001;
      50729: inst = 32'hfe0d96a;
      50730: inst = 32'h5be00000;
      50731: inst = 32'h8c50000;
      50732: inst = 32'h24612800;
      50733: inst = 32'h10a0ffff;
      50734: inst = 32'hca0ffeb;
      50735: inst = 32'h24822800;
      50736: inst = 32'h10a00000;
      50737: inst = 32'hca00004;
      50738: inst = 32'h38632800;
      50739: inst = 32'h38842800;
      50740: inst = 32'h10a00000;
      50741: inst = 32'hca0c639;
      50742: inst = 32'h13e00001;
      50743: inst = 32'hfe0d96a;
      50744: inst = 32'h5be00000;
      50745: inst = 32'h8c50000;
      50746: inst = 32'h24612800;
      50747: inst = 32'h10a0ffff;
      50748: inst = 32'hca0ffeb;
      50749: inst = 32'h24822800;
      50750: inst = 32'h10a00000;
      50751: inst = 32'hca00004;
      50752: inst = 32'h38632800;
      50753: inst = 32'h38842800;
      50754: inst = 32'h10a00000;
      50755: inst = 32'hca0c647;
      50756: inst = 32'h13e00001;
      50757: inst = 32'hfe0d96a;
      50758: inst = 32'h5be00000;
      50759: inst = 32'h8c50000;
      50760: inst = 32'h24612800;
      50761: inst = 32'h10a0ffff;
      50762: inst = 32'hca0ffeb;
      50763: inst = 32'h24822800;
      50764: inst = 32'h10a00000;
      50765: inst = 32'hca00004;
      50766: inst = 32'h38632800;
      50767: inst = 32'h38842800;
      50768: inst = 32'h10a00000;
      50769: inst = 32'hca0c655;
      50770: inst = 32'h13e00001;
      50771: inst = 32'hfe0d96a;
      50772: inst = 32'h5be00000;
      50773: inst = 32'h8c50000;
      50774: inst = 32'h24612800;
      50775: inst = 32'h10a0ffff;
      50776: inst = 32'hca0ffeb;
      50777: inst = 32'h24822800;
      50778: inst = 32'h10a00000;
      50779: inst = 32'hca00004;
      50780: inst = 32'h38632800;
      50781: inst = 32'h38842800;
      50782: inst = 32'h10a00000;
      50783: inst = 32'hca0c663;
      50784: inst = 32'h13e00001;
      50785: inst = 32'hfe0d96a;
      50786: inst = 32'h5be00000;
      50787: inst = 32'h8c50000;
      50788: inst = 32'h24612800;
      50789: inst = 32'h10a0ffff;
      50790: inst = 32'hca0ffeb;
      50791: inst = 32'h24822800;
      50792: inst = 32'h10a00000;
      50793: inst = 32'hca00004;
      50794: inst = 32'h38632800;
      50795: inst = 32'h38842800;
      50796: inst = 32'h10a00000;
      50797: inst = 32'hca0c671;
      50798: inst = 32'h13e00001;
      50799: inst = 32'hfe0d96a;
      50800: inst = 32'h5be00000;
      50801: inst = 32'h8c50000;
      50802: inst = 32'h24612800;
      50803: inst = 32'h10a0ffff;
      50804: inst = 32'hca0ffeb;
      50805: inst = 32'h24822800;
      50806: inst = 32'h10a00000;
      50807: inst = 32'hca00004;
      50808: inst = 32'h38632800;
      50809: inst = 32'h38842800;
      50810: inst = 32'h10a00000;
      50811: inst = 32'hca0c67f;
      50812: inst = 32'h13e00001;
      50813: inst = 32'hfe0d96a;
      50814: inst = 32'h5be00000;
      50815: inst = 32'h8c50000;
      50816: inst = 32'h24612800;
      50817: inst = 32'h10a0ffff;
      50818: inst = 32'hca0ffeb;
      50819: inst = 32'h24822800;
      50820: inst = 32'h10a00000;
      50821: inst = 32'hca00004;
      50822: inst = 32'h38632800;
      50823: inst = 32'h38842800;
      50824: inst = 32'h10a00000;
      50825: inst = 32'hca0c68d;
      50826: inst = 32'h13e00001;
      50827: inst = 32'hfe0d96a;
      50828: inst = 32'h5be00000;
      50829: inst = 32'h8c50000;
      50830: inst = 32'h24612800;
      50831: inst = 32'h10a0ffff;
      50832: inst = 32'hca0ffeb;
      50833: inst = 32'h24822800;
      50834: inst = 32'h10a00000;
      50835: inst = 32'hca00004;
      50836: inst = 32'h38632800;
      50837: inst = 32'h38842800;
      50838: inst = 32'h10a00000;
      50839: inst = 32'hca0c69b;
      50840: inst = 32'h13e00001;
      50841: inst = 32'hfe0d96a;
      50842: inst = 32'h5be00000;
      50843: inst = 32'h8c50000;
      50844: inst = 32'h24612800;
      50845: inst = 32'h10a0ffff;
      50846: inst = 32'hca0ffeb;
      50847: inst = 32'h24822800;
      50848: inst = 32'h10a00000;
      50849: inst = 32'hca00004;
      50850: inst = 32'h38632800;
      50851: inst = 32'h38842800;
      50852: inst = 32'h10a00000;
      50853: inst = 32'hca0c6a9;
      50854: inst = 32'h13e00001;
      50855: inst = 32'hfe0d96a;
      50856: inst = 32'h5be00000;
      50857: inst = 32'h8c50000;
      50858: inst = 32'h24612800;
      50859: inst = 32'h10a0ffff;
      50860: inst = 32'hca0ffeb;
      50861: inst = 32'h24822800;
      50862: inst = 32'h10a00000;
      50863: inst = 32'hca00004;
      50864: inst = 32'h38632800;
      50865: inst = 32'h38842800;
      50866: inst = 32'h10a00000;
      50867: inst = 32'hca0c6b7;
      50868: inst = 32'h13e00001;
      50869: inst = 32'hfe0d96a;
      50870: inst = 32'h5be00000;
      50871: inst = 32'h8c50000;
      50872: inst = 32'h24612800;
      50873: inst = 32'h10a0ffff;
      50874: inst = 32'hca0ffeb;
      50875: inst = 32'h24822800;
      50876: inst = 32'h10a00000;
      50877: inst = 32'hca00004;
      50878: inst = 32'h38632800;
      50879: inst = 32'h38842800;
      50880: inst = 32'h10a00000;
      50881: inst = 32'hca0c6c5;
      50882: inst = 32'h13e00001;
      50883: inst = 32'hfe0d96a;
      50884: inst = 32'h5be00000;
      50885: inst = 32'h8c50000;
      50886: inst = 32'h24612800;
      50887: inst = 32'h10a0ffff;
      50888: inst = 32'hca0ffeb;
      50889: inst = 32'h24822800;
      50890: inst = 32'h10a00000;
      50891: inst = 32'hca00004;
      50892: inst = 32'h38632800;
      50893: inst = 32'h38842800;
      50894: inst = 32'h10a00000;
      50895: inst = 32'hca0c6d3;
      50896: inst = 32'h13e00001;
      50897: inst = 32'hfe0d96a;
      50898: inst = 32'h5be00000;
      50899: inst = 32'h8c50000;
      50900: inst = 32'h24612800;
      50901: inst = 32'h10a0ffff;
      50902: inst = 32'hca0ffeb;
      50903: inst = 32'h24822800;
      50904: inst = 32'h10a00000;
      50905: inst = 32'hca00004;
      50906: inst = 32'h38632800;
      50907: inst = 32'h38842800;
      50908: inst = 32'h10a00000;
      50909: inst = 32'hca0c6e1;
      50910: inst = 32'h13e00001;
      50911: inst = 32'hfe0d96a;
      50912: inst = 32'h5be00000;
      50913: inst = 32'h8c50000;
      50914: inst = 32'h24612800;
      50915: inst = 32'h10a0ffff;
      50916: inst = 32'hca0ffeb;
      50917: inst = 32'h24822800;
      50918: inst = 32'h10a00000;
      50919: inst = 32'hca00004;
      50920: inst = 32'h38632800;
      50921: inst = 32'h38842800;
      50922: inst = 32'h10a00000;
      50923: inst = 32'hca0c6ef;
      50924: inst = 32'h13e00001;
      50925: inst = 32'hfe0d96a;
      50926: inst = 32'h5be00000;
      50927: inst = 32'h8c50000;
      50928: inst = 32'h24612800;
      50929: inst = 32'h10a0ffff;
      50930: inst = 32'hca0ffeb;
      50931: inst = 32'h24822800;
      50932: inst = 32'h10a00000;
      50933: inst = 32'hca00004;
      50934: inst = 32'h38632800;
      50935: inst = 32'h38842800;
      50936: inst = 32'h10a00000;
      50937: inst = 32'hca0c6fd;
      50938: inst = 32'h13e00001;
      50939: inst = 32'hfe0d96a;
      50940: inst = 32'h5be00000;
      50941: inst = 32'h8c50000;
      50942: inst = 32'h24612800;
      50943: inst = 32'h10a0ffff;
      50944: inst = 32'hca0ffeb;
      50945: inst = 32'h24822800;
      50946: inst = 32'h10a00000;
      50947: inst = 32'hca00004;
      50948: inst = 32'h38632800;
      50949: inst = 32'h38842800;
      50950: inst = 32'h10a00000;
      50951: inst = 32'hca0c70b;
      50952: inst = 32'h13e00001;
      50953: inst = 32'hfe0d96a;
      50954: inst = 32'h5be00000;
      50955: inst = 32'h8c50000;
      50956: inst = 32'h24612800;
      50957: inst = 32'h10a0ffff;
      50958: inst = 32'hca0ffeb;
      50959: inst = 32'h24822800;
      50960: inst = 32'h10a00000;
      50961: inst = 32'hca00004;
      50962: inst = 32'h38632800;
      50963: inst = 32'h38842800;
      50964: inst = 32'h10a00000;
      50965: inst = 32'hca0c719;
      50966: inst = 32'h13e00001;
      50967: inst = 32'hfe0d96a;
      50968: inst = 32'h5be00000;
      50969: inst = 32'h8c50000;
      50970: inst = 32'h24612800;
      50971: inst = 32'h10a0ffff;
      50972: inst = 32'hca0ffeb;
      50973: inst = 32'h24822800;
      50974: inst = 32'h10a00000;
      50975: inst = 32'hca00004;
      50976: inst = 32'h38632800;
      50977: inst = 32'h38842800;
      50978: inst = 32'h10a00000;
      50979: inst = 32'hca0c727;
      50980: inst = 32'h13e00001;
      50981: inst = 32'hfe0d96a;
      50982: inst = 32'h5be00000;
      50983: inst = 32'h8c50000;
      50984: inst = 32'h24612800;
      50985: inst = 32'h10a0ffff;
      50986: inst = 32'hca0ffeb;
      50987: inst = 32'h24822800;
      50988: inst = 32'h10a00000;
      50989: inst = 32'hca00004;
      50990: inst = 32'h38632800;
      50991: inst = 32'h38842800;
      50992: inst = 32'h10a00000;
      50993: inst = 32'hca0c735;
      50994: inst = 32'h13e00001;
      50995: inst = 32'hfe0d96a;
      50996: inst = 32'h5be00000;
      50997: inst = 32'h8c50000;
      50998: inst = 32'h24612800;
      50999: inst = 32'h10a0ffff;
      51000: inst = 32'hca0ffeb;
      51001: inst = 32'h24822800;
      51002: inst = 32'h10a00000;
      51003: inst = 32'hca00004;
      51004: inst = 32'h38632800;
      51005: inst = 32'h38842800;
      51006: inst = 32'h10a00000;
      51007: inst = 32'hca0c743;
      51008: inst = 32'h13e00001;
      51009: inst = 32'hfe0d96a;
      51010: inst = 32'h5be00000;
      51011: inst = 32'h8c50000;
      51012: inst = 32'h24612800;
      51013: inst = 32'h10a0ffff;
      51014: inst = 32'hca0ffeb;
      51015: inst = 32'h24822800;
      51016: inst = 32'h10a00000;
      51017: inst = 32'hca00004;
      51018: inst = 32'h38632800;
      51019: inst = 32'h38842800;
      51020: inst = 32'h10a00000;
      51021: inst = 32'hca0c751;
      51022: inst = 32'h13e00001;
      51023: inst = 32'hfe0d96a;
      51024: inst = 32'h5be00000;
      51025: inst = 32'h8c50000;
      51026: inst = 32'h24612800;
      51027: inst = 32'h10a0ffff;
      51028: inst = 32'hca0ffeb;
      51029: inst = 32'h24822800;
      51030: inst = 32'h10a00000;
      51031: inst = 32'hca00004;
      51032: inst = 32'h38632800;
      51033: inst = 32'h38842800;
      51034: inst = 32'h10a00000;
      51035: inst = 32'hca0c75f;
      51036: inst = 32'h13e00001;
      51037: inst = 32'hfe0d96a;
      51038: inst = 32'h5be00000;
      51039: inst = 32'h8c50000;
      51040: inst = 32'h24612800;
      51041: inst = 32'h10a0ffff;
      51042: inst = 32'hca0ffeb;
      51043: inst = 32'h24822800;
      51044: inst = 32'h10a00000;
      51045: inst = 32'hca00004;
      51046: inst = 32'h38632800;
      51047: inst = 32'h38842800;
      51048: inst = 32'h10a00000;
      51049: inst = 32'hca0c76d;
      51050: inst = 32'h13e00001;
      51051: inst = 32'hfe0d96a;
      51052: inst = 32'h5be00000;
      51053: inst = 32'h8c50000;
      51054: inst = 32'h24612800;
      51055: inst = 32'h10a0ffff;
      51056: inst = 32'hca0ffeb;
      51057: inst = 32'h24822800;
      51058: inst = 32'h10a00000;
      51059: inst = 32'hca00004;
      51060: inst = 32'h38632800;
      51061: inst = 32'h38842800;
      51062: inst = 32'h10a00000;
      51063: inst = 32'hca0c77b;
      51064: inst = 32'h13e00001;
      51065: inst = 32'hfe0d96a;
      51066: inst = 32'h5be00000;
      51067: inst = 32'h8c50000;
      51068: inst = 32'h24612800;
      51069: inst = 32'h10a0ffff;
      51070: inst = 32'hca0ffeb;
      51071: inst = 32'h24822800;
      51072: inst = 32'h10a00000;
      51073: inst = 32'hca00004;
      51074: inst = 32'h38632800;
      51075: inst = 32'h38842800;
      51076: inst = 32'h10a00000;
      51077: inst = 32'hca0c789;
      51078: inst = 32'h13e00001;
      51079: inst = 32'hfe0d96a;
      51080: inst = 32'h5be00000;
      51081: inst = 32'h8c50000;
      51082: inst = 32'h24612800;
      51083: inst = 32'h10a0ffff;
      51084: inst = 32'hca0ffeb;
      51085: inst = 32'h24822800;
      51086: inst = 32'h10a00000;
      51087: inst = 32'hca00004;
      51088: inst = 32'h38632800;
      51089: inst = 32'h38842800;
      51090: inst = 32'h10a00000;
      51091: inst = 32'hca0c797;
      51092: inst = 32'h13e00001;
      51093: inst = 32'hfe0d96a;
      51094: inst = 32'h5be00000;
      51095: inst = 32'h8c50000;
      51096: inst = 32'h24612800;
      51097: inst = 32'h10a0ffff;
      51098: inst = 32'hca0ffeb;
      51099: inst = 32'h24822800;
      51100: inst = 32'h10a00000;
      51101: inst = 32'hca00004;
      51102: inst = 32'h38632800;
      51103: inst = 32'h38842800;
      51104: inst = 32'h10a00000;
      51105: inst = 32'hca0c7a5;
      51106: inst = 32'h13e00001;
      51107: inst = 32'hfe0d96a;
      51108: inst = 32'h5be00000;
      51109: inst = 32'h8c50000;
      51110: inst = 32'h24612800;
      51111: inst = 32'h10a0ffff;
      51112: inst = 32'hca0ffeb;
      51113: inst = 32'h24822800;
      51114: inst = 32'h10a00000;
      51115: inst = 32'hca00004;
      51116: inst = 32'h38632800;
      51117: inst = 32'h38842800;
      51118: inst = 32'h10a00000;
      51119: inst = 32'hca0c7b3;
      51120: inst = 32'h13e00001;
      51121: inst = 32'hfe0d96a;
      51122: inst = 32'h5be00000;
      51123: inst = 32'h8c50000;
      51124: inst = 32'h24612800;
      51125: inst = 32'h10a0ffff;
      51126: inst = 32'hca0ffeb;
      51127: inst = 32'h24822800;
      51128: inst = 32'h10a00000;
      51129: inst = 32'hca00004;
      51130: inst = 32'h38632800;
      51131: inst = 32'h38842800;
      51132: inst = 32'h10a00000;
      51133: inst = 32'hca0c7c1;
      51134: inst = 32'h13e00001;
      51135: inst = 32'hfe0d96a;
      51136: inst = 32'h5be00000;
      51137: inst = 32'h8c50000;
      51138: inst = 32'h24612800;
      51139: inst = 32'h10a0ffff;
      51140: inst = 32'hca0ffeb;
      51141: inst = 32'h24822800;
      51142: inst = 32'h10a00000;
      51143: inst = 32'hca00004;
      51144: inst = 32'h38632800;
      51145: inst = 32'h38842800;
      51146: inst = 32'h10a00000;
      51147: inst = 32'hca0c7cf;
      51148: inst = 32'h13e00001;
      51149: inst = 32'hfe0d96a;
      51150: inst = 32'h5be00000;
      51151: inst = 32'h8c50000;
      51152: inst = 32'h24612800;
      51153: inst = 32'h10a0ffff;
      51154: inst = 32'hca0ffeb;
      51155: inst = 32'h24822800;
      51156: inst = 32'h10a00000;
      51157: inst = 32'hca00004;
      51158: inst = 32'h38632800;
      51159: inst = 32'h38842800;
      51160: inst = 32'h10a00000;
      51161: inst = 32'hca0c7dd;
      51162: inst = 32'h13e00001;
      51163: inst = 32'hfe0d96a;
      51164: inst = 32'h5be00000;
      51165: inst = 32'h8c50000;
      51166: inst = 32'h24612800;
      51167: inst = 32'h10a0ffff;
      51168: inst = 32'hca0ffeb;
      51169: inst = 32'h24822800;
      51170: inst = 32'h10a00000;
      51171: inst = 32'hca00004;
      51172: inst = 32'h38632800;
      51173: inst = 32'h38842800;
      51174: inst = 32'h10a00000;
      51175: inst = 32'hca0c7eb;
      51176: inst = 32'h13e00001;
      51177: inst = 32'hfe0d96a;
      51178: inst = 32'h5be00000;
      51179: inst = 32'h8c50000;
      51180: inst = 32'h24612800;
      51181: inst = 32'h10a0ffff;
      51182: inst = 32'hca0ffeb;
      51183: inst = 32'h24822800;
      51184: inst = 32'h10a00000;
      51185: inst = 32'hca00004;
      51186: inst = 32'h38632800;
      51187: inst = 32'h38842800;
      51188: inst = 32'h10a00000;
      51189: inst = 32'hca0c7f9;
      51190: inst = 32'h13e00001;
      51191: inst = 32'hfe0d96a;
      51192: inst = 32'h5be00000;
      51193: inst = 32'h8c50000;
      51194: inst = 32'h24612800;
      51195: inst = 32'h10a0ffff;
      51196: inst = 32'hca0ffeb;
      51197: inst = 32'h24822800;
      51198: inst = 32'h10a00000;
      51199: inst = 32'hca00004;
      51200: inst = 32'h38632800;
      51201: inst = 32'h38842800;
      51202: inst = 32'h10a00000;
      51203: inst = 32'hca0c807;
      51204: inst = 32'h13e00001;
      51205: inst = 32'hfe0d96a;
      51206: inst = 32'h5be00000;
      51207: inst = 32'h8c50000;
      51208: inst = 32'h24612800;
      51209: inst = 32'h10a0ffff;
      51210: inst = 32'hca0ffeb;
      51211: inst = 32'h24822800;
      51212: inst = 32'h10a00000;
      51213: inst = 32'hca00004;
      51214: inst = 32'h38632800;
      51215: inst = 32'h38842800;
      51216: inst = 32'h10a00000;
      51217: inst = 32'hca0c815;
      51218: inst = 32'h13e00001;
      51219: inst = 32'hfe0d96a;
      51220: inst = 32'h5be00000;
      51221: inst = 32'h8c50000;
      51222: inst = 32'h24612800;
      51223: inst = 32'h10a0ffff;
      51224: inst = 32'hca0ffeb;
      51225: inst = 32'h24822800;
      51226: inst = 32'h10a00000;
      51227: inst = 32'hca00004;
      51228: inst = 32'h38632800;
      51229: inst = 32'h38842800;
      51230: inst = 32'h10a00000;
      51231: inst = 32'hca0c823;
      51232: inst = 32'h13e00001;
      51233: inst = 32'hfe0d96a;
      51234: inst = 32'h5be00000;
      51235: inst = 32'h8c50000;
      51236: inst = 32'h24612800;
      51237: inst = 32'h10a0ffff;
      51238: inst = 32'hca0ffeb;
      51239: inst = 32'h24822800;
      51240: inst = 32'h10a00000;
      51241: inst = 32'hca00004;
      51242: inst = 32'h38632800;
      51243: inst = 32'h38842800;
      51244: inst = 32'h10a00000;
      51245: inst = 32'hca0c831;
      51246: inst = 32'h13e00001;
      51247: inst = 32'hfe0d96a;
      51248: inst = 32'h5be00000;
      51249: inst = 32'h8c50000;
      51250: inst = 32'h24612800;
      51251: inst = 32'h10a0ffff;
      51252: inst = 32'hca0ffeb;
      51253: inst = 32'h24822800;
      51254: inst = 32'h10a00000;
      51255: inst = 32'hca00004;
      51256: inst = 32'h38632800;
      51257: inst = 32'h38842800;
      51258: inst = 32'h10a00000;
      51259: inst = 32'hca0c83f;
      51260: inst = 32'h13e00001;
      51261: inst = 32'hfe0d96a;
      51262: inst = 32'h5be00000;
      51263: inst = 32'h8c50000;
      51264: inst = 32'h24612800;
      51265: inst = 32'h10a0ffff;
      51266: inst = 32'hca0ffeb;
      51267: inst = 32'h24822800;
      51268: inst = 32'h10a00000;
      51269: inst = 32'hca00004;
      51270: inst = 32'h38632800;
      51271: inst = 32'h38842800;
      51272: inst = 32'h10a00000;
      51273: inst = 32'hca0c84d;
      51274: inst = 32'h13e00001;
      51275: inst = 32'hfe0d96a;
      51276: inst = 32'h5be00000;
      51277: inst = 32'h8c50000;
      51278: inst = 32'h24612800;
      51279: inst = 32'h10a0ffff;
      51280: inst = 32'hca0ffeb;
      51281: inst = 32'h24822800;
      51282: inst = 32'h10a00000;
      51283: inst = 32'hca00004;
      51284: inst = 32'h38632800;
      51285: inst = 32'h38842800;
      51286: inst = 32'h10a00000;
      51287: inst = 32'hca0c85b;
      51288: inst = 32'h13e00001;
      51289: inst = 32'hfe0d96a;
      51290: inst = 32'h5be00000;
      51291: inst = 32'h8c50000;
      51292: inst = 32'h24612800;
      51293: inst = 32'h10a0ffff;
      51294: inst = 32'hca0ffeb;
      51295: inst = 32'h24822800;
      51296: inst = 32'h10a00000;
      51297: inst = 32'hca00004;
      51298: inst = 32'h38632800;
      51299: inst = 32'h38842800;
      51300: inst = 32'h10a00000;
      51301: inst = 32'hca0c869;
      51302: inst = 32'h13e00001;
      51303: inst = 32'hfe0d96a;
      51304: inst = 32'h5be00000;
      51305: inst = 32'h8c50000;
      51306: inst = 32'h24612800;
      51307: inst = 32'h10a0ffff;
      51308: inst = 32'hca0ffec;
      51309: inst = 32'h24822800;
      51310: inst = 32'h10a00000;
      51311: inst = 32'hca00004;
      51312: inst = 32'h38632800;
      51313: inst = 32'h38842800;
      51314: inst = 32'h10a00000;
      51315: inst = 32'hca0c877;
      51316: inst = 32'h13e00001;
      51317: inst = 32'hfe0d96a;
      51318: inst = 32'h5be00000;
      51319: inst = 32'h8c50000;
      51320: inst = 32'h24612800;
      51321: inst = 32'h10a0ffff;
      51322: inst = 32'hca0ffec;
      51323: inst = 32'h24822800;
      51324: inst = 32'h10a00000;
      51325: inst = 32'hca00004;
      51326: inst = 32'h38632800;
      51327: inst = 32'h38842800;
      51328: inst = 32'h10a00000;
      51329: inst = 32'hca0c885;
      51330: inst = 32'h13e00001;
      51331: inst = 32'hfe0d96a;
      51332: inst = 32'h5be00000;
      51333: inst = 32'h8c50000;
      51334: inst = 32'h24612800;
      51335: inst = 32'h10a0ffff;
      51336: inst = 32'hca0ffec;
      51337: inst = 32'h24822800;
      51338: inst = 32'h10a00000;
      51339: inst = 32'hca00004;
      51340: inst = 32'h38632800;
      51341: inst = 32'h38842800;
      51342: inst = 32'h10a00000;
      51343: inst = 32'hca0c893;
      51344: inst = 32'h13e00001;
      51345: inst = 32'hfe0d96a;
      51346: inst = 32'h5be00000;
      51347: inst = 32'h8c50000;
      51348: inst = 32'h24612800;
      51349: inst = 32'h10a0ffff;
      51350: inst = 32'hca0ffec;
      51351: inst = 32'h24822800;
      51352: inst = 32'h10a00000;
      51353: inst = 32'hca00004;
      51354: inst = 32'h38632800;
      51355: inst = 32'h38842800;
      51356: inst = 32'h10a00000;
      51357: inst = 32'hca0c8a1;
      51358: inst = 32'h13e00001;
      51359: inst = 32'hfe0d96a;
      51360: inst = 32'h5be00000;
      51361: inst = 32'h8c50000;
      51362: inst = 32'h24612800;
      51363: inst = 32'h10a0ffff;
      51364: inst = 32'hca0ffec;
      51365: inst = 32'h24822800;
      51366: inst = 32'h10a00000;
      51367: inst = 32'hca00004;
      51368: inst = 32'h38632800;
      51369: inst = 32'h38842800;
      51370: inst = 32'h10a00000;
      51371: inst = 32'hca0c8af;
      51372: inst = 32'h13e00001;
      51373: inst = 32'hfe0d96a;
      51374: inst = 32'h5be00000;
      51375: inst = 32'h8c50000;
      51376: inst = 32'h24612800;
      51377: inst = 32'h10a0ffff;
      51378: inst = 32'hca0ffec;
      51379: inst = 32'h24822800;
      51380: inst = 32'h10a00000;
      51381: inst = 32'hca00004;
      51382: inst = 32'h38632800;
      51383: inst = 32'h38842800;
      51384: inst = 32'h10a00000;
      51385: inst = 32'hca0c8bd;
      51386: inst = 32'h13e00001;
      51387: inst = 32'hfe0d96a;
      51388: inst = 32'h5be00000;
      51389: inst = 32'h8c50000;
      51390: inst = 32'h24612800;
      51391: inst = 32'h10a0ffff;
      51392: inst = 32'hca0ffec;
      51393: inst = 32'h24822800;
      51394: inst = 32'h10a00000;
      51395: inst = 32'hca00004;
      51396: inst = 32'h38632800;
      51397: inst = 32'h38842800;
      51398: inst = 32'h10a00000;
      51399: inst = 32'hca0c8cb;
      51400: inst = 32'h13e00001;
      51401: inst = 32'hfe0d96a;
      51402: inst = 32'h5be00000;
      51403: inst = 32'h8c50000;
      51404: inst = 32'h24612800;
      51405: inst = 32'h10a0ffff;
      51406: inst = 32'hca0ffec;
      51407: inst = 32'h24822800;
      51408: inst = 32'h10a00000;
      51409: inst = 32'hca00004;
      51410: inst = 32'h38632800;
      51411: inst = 32'h38842800;
      51412: inst = 32'h10a00000;
      51413: inst = 32'hca0c8d9;
      51414: inst = 32'h13e00001;
      51415: inst = 32'hfe0d96a;
      51416: inst = 32'h5be00000;
      51417: inst = 32'h8c50000;
      51418: inst = 32'h24612800;
      51419: inst = 32'h10a0ffff;
      51420: inst = 32'hca0ffec;
      51421: inst = 32'h24822800;
      51422: inst = 32'h10a00000;
      51423: inst = 32'hca00004;
      51424: inst = 32'h38632800;
      51425: inst = 32'h38842800;
      51426: inst = 32'h10a00000;
      51427: inst = 32'hca0c8e7;
      51428: inst = 32'h13e00001;
      51429: inst = 32'hfe0d96a;
      51430: inst = 32'h5be00000;
      51431: inst = 32'h8c50000;
      51432: inst = 32'h24612800;
      51433: inst = 32'h10a0ffff;
      51434: inst = 32'hca0ffec;
      51435: inst = 32'h24822800;
      51436: inst = 32'h10a00000;
      51437: inst = 32'hca00004;
      51438: inst = 32'h38632800;
      51439: inst = 32'h38842800;
      51440: inst = 32'h10a00000;
      51441: inst = 32'hca0c8f5;
      51442: inst = 32'h13e00001;
      51443: inst = 32'hfe0d96a;
      51444: inst = 32'h5be00000;
      51445: inst = 32'h8c50000;
      51446: inst = 32'h24612800;
      51447: inst = 32'h10a0ffff;
      51448: inst = 32'hca0ffec;
      51449: inst = 32'h24822800;
      51450: inst = 32'h10a00000;
      51451: inst = 32'hca00004;
      51452: inst = 32'h38632800;
      51453: inst = 32'h38842800;
      51454: inst = 32'h10a00000;
      51455: inst = 32'hca0c903;
      51456: inst = 32'h13e00001;
      51457: inst = 32'hfe0d96a;
      51458: inst = 32'h5be00000;
      51459: inst = 32'h8c50000;
      51460: inst = 32'h24612800;
      51461: inst = 32'h10a0ffff;
      51462: inst = 32'hca0ffec;
      51463: inst = 32'h24822800;
      51464: inst = 32'h10a00000;
      51465: inst = 32'hca00004;
      51466: inst = 32'h38632800;
      51467: inst = 32'h38842800;
      51468: inst = 32'h10a00000;
      51469: inst = 32'hca0c911;
      51470: inst = 32'h13e00001;
      51471: inst = 32'hfe0d96a;
      51472: inst = 32'h5be00000;
      51473: inst = 32'h8c50000;
      51474: inst = 32'h24612800;
      51475: inst = 32'h10a0ffff;
      51476: inst = 32'hca0ffec;
      51477: inst = 32'h24822800;
      51478: inst = 32'h10a00000;
      51479: inst = 32'hca00004;
      51480: inst = 32'h38632800;
      51481: inst = 32'h38842800;
      51482: inst = 32'h10a00000;
      51483: inst = 32'hca0c91f;
      51484: inst = 32'h13e00001;
      51485: inst = 32'hfe0d96a;
      51486: inst = 32'h5be00000;
      51487: inst = 32'h8c50000;
      51488: inst = 32'h24612800;
      51489: inst = 32'h10a0ffff;
      51490: inst = 32'hca0ffec;
      51491: inst = 32'h24822800;
      51492: inst = 32'h10a00000;
      51493: inst = 32'hca00004;
      51494: inst = 32'h38632800;
      51495: inst = 32'h38842800;
      51496: inst = 32'h10a00000;
      51497: inst = 32'hca0c92d;
      51498: inst = 32'h13e00001;
      51499: inst = 32'hfe0d96a;
      51500: inst = 32'h5be00000;
      51501: inst = 32'h8c50000;
      51502: inst = 32'h24612800;
      51503: inst = 32'h10a0ffff;
      51504: inst = 32'hca0ffec;
      51505: inst = 32'h24822800;
      51506: inst = 32'h10a00000;
      51507: inst = 32'hca00004;
      51508: inst = 32'h38632800;
      51509: inst = 32'h38842800;
      51510: inst = 32'h10a00000;
      51511: inst = 32'hca0c93b;
      51512: inst = 32'h13e00001;
      51513: inst = 32'hfe0d96a;
      51514: inst = 32'h5be00000;
      51515: inst = 32'h8c50000;
      51516: inst = 32'h24612800;
      51517: inst = 32'h10a0ffff;
      51518: inst = 32'hca0ffec;
      51519: inst = 32'h24822800;
      51520: inst = 32'h10a00000;
      51521: inst = 32'hca00004;
      51522: inst = 32'h38632800;
      51523: inst = 32'h38842800;
      51524: inst = 32'h10a00000;
      51525: inst = 32'hca0c949;
      51526: inst = 32'h13e00001;
      51527: inst = 32'hfe0d96a;
      51528: inst = 32'h5be00000;
      51529: inst = 32'h8c50000;
      51530: inst = 32'h24612800;
      51531: inst = 32'h10a0ffff;
      51532: inst = 32'hca0ffec;
      51533: inst = 32'h24822800;
      51534: inst = 32'h10a00000;
      51535: inst = 32'hca00004;
      51536: inst = 32'h38632800;
      51537: inst = 32'h38842800;
      51538: inst = 32'h10a00000;
      51539: inst = 32'hca0c957;
      51540: inst = 32'h13e00001;
      51541: inst = 32'hfe0d96a;
      51542: inst = 32'h5be00000;
      51543: inst = 32'h8c50000;
      51544: inst = 32'h24612800;
      51545: inst = 32'h10a0ffff;
      51546: inst = 32'hca0ffec;
      51547: inst = 32'h24822800;
      51548: inst = 32'h10a00000;
      51549: inst = 32'hca00004;
      51550: inst = 32'h38632800;
      51551: inst = 32'h38842800;
      51552: inst = 32'h10a00000;
      51553: inst = 32'hca0c965;
      51554: inst = 32'h13e00001;
      51555: inst = 32'hfe0d96a;
      51556: inst = 32'h5be00000;
      51557: inst = 32'h8c50000;
      51558: inst = 32'h24612800;
      51559: inst = 32'h10a0ffff;
      51560: inst = 32'hca0ffec;
      51561: inst = 32'h24822800;
      51562: inst = 32'h10a00000;
      51563: inst = 32'hca00004;
      51564: inst = 32'h38632800;
      51565: inst = 32'h38842800;
      51566: inst = 32'h10a00000;
      51567: inst = 32'hca0c973;
      51568: inst = 32'h13e00001;
      51569: inst = 32'hfe0d96a;
      51570: inst = 32'h5be00000;
      51571: inst = 32'h8c50000;
      51572: inst = 32'h24612800;
      51573: inst = 32'h10a0ffff;
      51574: inst = 32'hca0ffec;
      51575: inst = 32'h24822800;
      51576: inst = 32'h10a00000;
      51577: inst = 32'hca00004;
      51578: inst = 32'h38632800;
      51579: inst = 32'h38842800;
      51580: inst = 32'h10a00000;
      51581: inst = 32'hca0c981;
      51582: inst = 32'h13e00001;
      51583: inst = 32'hfe0d96a;
      51584: inst = 32'h5be00000;
      51585: inst = 32'h8c50000;
      51586: inst = 32'h24612800;
      51587: inst = 32'h10a0ffff;
      51588: inst = 32'hca0ffec;
      51589: inst = 32'h24822800;
      51590: inst = 32'h10a00000;
      51591: inst = 32'hca00004;
      51592: inst = 32'h38632800;
      51593: inst = 32'h38842800;
      51594: inst = 32'h10a00000;
      51595: inst = 32'hca0c98f;
      51596: inst = 32'h13e00001;
      51597: inst = 32'hfe0d96a;
      51598: inst = 32'h5be00000;
      51599: inst = 32'h8c50000;
      51600: inst = 32'h24612800;
      51601: inst = 32'h10a0ffff;
      51602: inst = 32'hca0ffec;
      51603: inst = 32'h24822800;
      51604: inst = 32'h10a00000;
      51605: inst = 32'hca00004;
      51606: inst = 32'h38632800;
      51607: inst = 32'h38842800;
      51608: inst = 32'h10a00000;
      51609: inst = 32'hca0c99d;
      51610: inst = 32'h13e00001;
      51611: inst = 32'hfe0d96a;
      51612: inst = 32'h5be00000;
      51613: inst = 32'h8c50000;
      51614: inst = 32'h24612800;
      51615: inst = 32'h10a0ffff;
      51616: inst = 32'hca0ffec;
      51617: inst = 32'h24822800;
      51618: inst = 32'h10a00000;
      51619: inst = 32'hca00004;
      51620: inst = 32'h38632800;
      51621: inst = 32'h38842800;
      51622: inst = 32'h10a00000;
      51623: inst = 32'hca0c9ab;
      51624: inst = 32'h13e00001;
      51625: inst = 32'hfe0d96a;
      51626: inst = 32'h5be00000;
      51627: inst = 32'h8c50000;
      51628: inst = 32'h24612800;
      51629: inst = 32'h10a0ffff;
      51630: inst = 32'hca0ffec;
      51631: inst = 32'h24822800;
      51632: inst = 32'h10a00000;
      51633: inst = 32'hca00004;
      51634: inst = 32'h38632800;
      51635: inst = 32'h38842800;
      51636: inst = 32'h10a00000;
      51637: inst = 32'hca0c9b9;
      51638: inst = 32'h13e00001;
      51639: inst = 32'hfe0d96a;
      51640: inst = 32'h5be00000;
      51641: inst = 32'h8c50000;
      51642: inst = 32'h24612800;
      51643: inst = 32'h10a0ffff;
      51644: inst = 32'hca0ffec;
      51645: inst = 32'h24822800;
      51646: inst = 32'h10a00000;
      51647: inst = 32'hca00004;
      51648: inst = 32'h38632800;
      51649: inst = 32'h38842800;
      51650: inst = 32'h10a00000;
      51651: inst = 32'hca0c9c7;
      51652: inst = 32'h13e00001;
      51653: inst = 32'hfe0d96a;
      51654: inst = 32'h5be00000;
      51655: inst = 32'h8c50000;
      51656: inst = 32'h24612800;
      51657: inst = 32'h10a0ffff;
      51658: inst = 32'hca0ffec;
      51659: inst = 32'h24822800;
      51660: inst = 32'h10a00000;
      51661: inst = 32'hca00004;
      51662: inst = 32'h38632800;
      51663: inst = 32'h38842800;
      51664: inst = 32'h10a00000;
      51665: inst = 32'hca0c9d5;
      51666: inst = 32'h13e00001;
      51667: inst = 32'hfe0d96a;
      51668: inst = 32'h5be00000;
      51669: inst = 32'h8c50000;
      51670: inst = 32'h24612800;
      51671: inst = 32'h10a0ffff;
      51672: inst = 32'hca0ffec;
      51673: inst = 32'h24822800;
      51674: inst = 32'h10a00000;
      51675: inst = 32'hca00004;
      51676: inst = 32'h38632800;
      51677: inst = 32'h38842800;
      51678: inst = 32'h10a00000;
      51679: inst = 32'hca0c9e3;
      51680: inst = 32'h13e00001;
      51681: inst = 32'hfe0d96a;
      51682: inst = 32'h5be00000;
      51683: inst = 32'h8c50000;
      51684: inst = 32'h24612800;
      51685: inst = 32'h10a0ffff;
      51686: inst = 32'hca0ffec;
      51687: inst = 32'h24822800;
      51688: inst = 32'h10a00000;
      51689: inst = 32'hca00004;
      51690: inst = 32'h38632800;
      51691: inst = 32'h38842800;
      51692: inst = 32'h10a00000;
      51693: inst = 32'hca0c9f1;
      51694: inst = 32'h13e00001;
      51695: inst = 32'hfe0d96a;
      51696: inst = 32'h5be00000;
      51697: inst = 32'h8c50000;
      51698: inst = 32'h24612800;
      51699: inst = 32'h10a0ffff;
      51700: inst = 32'hca0ffec;
      51701: inst = 32'h24822800;
      51702: inst = 32'h10a00000;
      51703: inst = 32'hca00004;
      51704: inst = 32'h38632800;
      51705: inst = 32'h38842800;
      51706: inst = 32'h10a00000;
      51707: inst = 32'hca0c9ff;
      51708: inst = 32'h13e00001;
      51709: inst = 32'hfe0d96a;
      51710: inst = 32'h5be00000;
      51711: inst = 32'h8c50000;
      51712: inst = 32'h24612800;
      51713: inst = 32'h10a0ffff;
      51714: inst = 32'hca0ffec;
      51715: inst = 32'h24822800;
      51716: inst = 32'h10a00000;
      51717: inst = 32'hca00004;
      51718: inst = 32'h38632800;
      51719: inst = 32'h38842800;
      51720: inst = 32'h10a00000;
      51721: inst = 32'hca0ca0d;
      51722: inst = 32'h13e00001;
      51723: inst = 32'hfe0d96a;
      51724: inst = 32'h5be00000;
      51725: inst = 32'h8c50000;
      51726: inst = 32'h24612800;
      51727: inst = 32'h10a0ffff;
      51728: inst = 32'hca0ffec;
      51729: inst = 32'h24822800;
      51730: inst = 32'h10a00000;
      51731: inst = 32'hca00004;
      51732: inst = 32'h38632800;
      51733: inst = 32'h38842800;
      51734: inst = 32'h10a00000;
      51735: inst = 32'hca0ca1b;
      51736: inst = 32'h13e00001;
      51737: inst = 32'hfe0d96a;
      51738: inst = 32'h5be00000;
      51739: inst = 32'h8c50000;
      51740: inst = 32'h24612800;
      51741: inst = 32'h10a0ffff;
      51742: inst = 32'hca0ffec;
      51743: inst = 32'h24822800;
      51744: inst = 32'h10a00000;
      51745: inst = 32'hca00004;
      51746: inst = 32'h38632800;
      51747: inst = 32'h38842800;
      51748: inst = 32'h10a00000;
      51749: inst = 32'hca0ca29;
      51750: inst = 32'h13e00001;
      51751: inst = 32'hfe0d96a;
      51752: inst = 32'h5be00000;
      51753: inst = 32'h8c50000;
      51754: inst = 32'h24612800;
      51755: inst = 32'h10a0ffff;
      51756: inst = 32'hca0ffec;
      51757: inst = 32'h24822800;
      51758: inst = 32'h10a00000;
      51759: inst = 32'hca00004;
      51760: inst = 32'h38632800;
      51761: inst = 32'h38842800;
      51762: inst = 32'h10a00000;
      51763: inst = 32'hca0ca37;
      51764: inst = 32'h13e00001;
      51765: inst = 32'hfe0d96a;
      51766: inst = 32'h5be00000;
      51767: inst = 32'h8c50000;
      51768: inst = 32'h24612800;
      51769: inst = 32'h10a0ffff;
      51770: inst = 32'hca0ffec;
      51771: inst = 32'h24822800;
      51772: inst = 32'h10a00000;
      51773: inst = 32'hca00004;
      51774: inst = 32'h38632800;
      51775: inst = 32'h38842800;
      51776: inst = 32'h10a00000;
      51777: inst = 32'hca0ca45;
      51778: inst = 32'h13e00001;
      51779: inst = 32'hfe0d96a;
      51780: inst = 32'h5be00000;
      51781: inst = 32'h8c50000;
      51782: inst = 32'h24612800;
      51783: inst = 32'h10a0ffff;
      51784: inst = 32'hca0ffec;
      51785: inst = 32'h24822800;
      51786: inst = 32'h10a00000;
      51787: inst = 32'hca00004;
      51788: inst = 32'h38632800;
      51789: inst = 32'h38842800;
      51790: inst = 32'h10a00000;
      51791: inst = 32'hca0ca53;
      51792: inst = 32'h13e00001;
      51793: inst = 32'hfe0d96a;
      51794: inst = 32'h5be00000;
      51795: inst = 32'h8c50000;
      51796: inst = 32'h24612800;
      51797: inst = 32'h10a0ffff;
      51798: inst = 32'hca0ffec;
      51799: inst = 32'h24822800;
      51800: inst = 32'h10a00000;
      51801: inst = 32'hca00004;
      51802: inst = 32'h38632800;
      51803: inst = 32'h38842800;
      51804: inst = 32'h10a00000;
      51805: inst = 32'hca0ca61;
      51806: inst = 32'h13e00001;
      51807: inst = 32'hfe0d96a;
      51808: inst = 32'h5be00000;
      51809: inst = 32'h8c50000;
      51810: inst = 32'h24612800;
      51811: inst = 32'h10a0ffff;
      51812: inst = 32'hca0ffec;
      51813: inst = 32'h24822800;
      51814: inst = 32'h10a00000;
      51815: inst = 32'hca00004;
      51816: inst = 32'h38632800;
      51817: inst = 32'h38842800;
      51818: inst = 32'h10a00000;
      51819: inst = 32'hca0ca6f;
      51820: inst = 32'h13e00001;
      51821: inst = 32'hfe0d96a;
      51822: inst = 32'h5be00000;
      51823: inst = 32'h8c50000;
      51824: inst = 32'h24612800;
      51825: inst = 32'h10a0ffff;
      51826: inst = 32'hca0ffec;
      51827: inst = 32'h24822800;
      51828: inst = 32'h10a00000;
      51829: inst = 32'hca00004;
      51830: inst = 32'h38632800;
      51831: inst = 32'h38842800;
      51832: inst = 32'h10a00000;
      51833: inst = 32'hca0ca7d;
      51834: inst = 32'h13e00001;
      51835: inst = 32'hfe0d96a;
      51836: inst = 32'h5be00000;
      51837: inst = 32'h8c50000;
      51838: inst = 32'h24612800;
      51839: inst = 32'h10a0ffff;
      51840: inst = 32'hca0ffec;
      51841: inst = 32'h24822800;
      51842: inst = 32'h10a00000;
      51843: inst = 32'hca00004;
      51844: inst = 32'h38632800;
      51845: inst = 32'h38842800;
      51846: inst = 32'h10a00000;
      51847: inst = 32'hca0ca8b;
      51848: inst = 32'h13e00001;
      51849: inst = 32'hfe0d96a;
      51850: inst = 32'h5be00000;
      51851: inst = 32'h8c50000;
      51852: inst = 32'h24612800;
      51853: inst = 32'h10a0ffff;
      51854: inst = 32'hca0ffec;
      51855: inst = 32'h24822800;
      51856: inst = 32'h10a00000;
      51857: inst = 32'hca00004;
      51858: inst = 32'h38632800;
      51859: inst = 32'h38842800;
      51860: inst = 32'h10a00000;
      51861: inst = 32'hca0ca99;
      51862: inst = 32'h13e00001;
      51863: inst = 32'hfe0d96a;
      51864: inst = 32'h5be00000;
      51865: inst = 32'h8c50000;
      51866: inst = 32'h24612800;
      51867: inst = 32'h10a0ffff;
      51868: inst = 32'hca0ffec;
      51869: inst = 32'h24822800;
      51870: inst = 32'h10a00000;
      51871: inst = 32'hca00004;
      51872: inst = 32'h38632800;
      51873: inst = 32'h38842800;
      51874: inst = 32'h10a00000;
      51875: inst = 32'hca0caa7;
      51876: inst = 32'h13e00001;
      51877: inst = 32'hfe0d96a;
      51878: inst = 32'h5be00000;
      51879: inst = 32'h8c50000;
      51880: inst = 32'h24612800;
      51881: inst = 32'h10a0ffff;
      51882: inst = 32'hca0ffec;
      51883: inst = 32'h24822800;
      51884: inst = 32'h10a00000;
      51885: inst = 32'hca00004;
      51886: inst = 32'h38632800;
      51887: inst = 32'h38842800;
      51888: inst = 32'h10a00000;
      51889: inst = 32'hca0cab5;
      51890: inst = 32'h13e00001;
      51891: inst = 32'hfe0d96a;
      51892: inst = 32'h5be00000;
      51893: inst = 32'h8c50000;
      51894: inst = 32'h24612800;
      51895: inst = 32'h10a0ffff;
      51896: inst = 32'hca0ffec;
      51897: inst = 32'h24822800;
      51898: inst = 32'h10a00000;
      51899: inst = 32'hca00004;
      51900: inst = 32'h38632800;
      51901: inst = 32'h38842800;
      51902: inst = 32'h10a00000;
      51903: inst = 32'hca0cac3;
      51904: inst = 32'h13e00001;
      51905: inst = 32'hfe0d96a;
      51906: inst = 32'h5be00000;
      51907: inst = 32'h8c50000;
      51908: inst = 32'h24612800;
      51909: inst = 32'h10a0ffff;
      51910: inst = 32'hca0ffec;
      51911: inst = 32'h24822800;
      51912: inst = 32'h10a00000;
      51913: inst = 32'hca00004;
      51914: inst = 32'h38632800;
      51915: inst = 32'h38842800;
      51916: inst = 32'h10a00000;
      51917: inst = 32'hca0cad1;
      51918: inst = 32'h13e00001;
      51919: inst = 32'hfe0d96a;
      51920: inst = 32'h5be00000;
      51921: inst = 32'h8c50000;
      51922: inst = 32'h24612800;
      51923: inst = 32'h10a0ffff;
      51924: inst = 32'hca0ffec;
      51925: inst = 32'h24822800;
      51926: inst = 32'h10a00000;
      51927: inst = 32'hca00004;
      51928: inst = 32'h38632800;
      51929: inst = 32'h38842800;
      51930: inst = 32'h10a00000;
      51931: inst = 32'hca0cadf;
      51932: inst = 32'h13e00001;
      51933: inst = 32'hfe0d96a;
      51934: inst = 32'h5be00000;
      51935: inst = 32'h8c50000;
      51936: inst = 32'h24612800;
      51937: inst = 32'h10a0ffff;
      51938: inst = 32'hca0ffec;
      51939: inst = 32'h24822800;
      51940: inst = 32'h10a00000;
      51941: inst = 32'hca00004;
      51942: inst = 32'h38632800;
      51943: inst = 32'h38842800;
      51944: inst = 32'h10a00000;
      51945: inst = 32'hca0caed;
      51946: inst = 32'h13e00001;
      51947: inst = 32'hfe0d96a;
      51948: inst = 32'h5be00000;
      51949: inst = 32'h8c50000;
      51950: inst = 32'h24612800;
      51951: inst = 32'h10a0ffff;
      51952: inst = 32'hca0ffec;
      51953: inst = 32'h24822800;
      51954: inst = 32'h10a00000;
      51955: inst = 32'hca00004;
      51956: inst = 32'h38632800;
      51957: inst = 32'h38842800;
      51958: inst = 32'h10a00000;
      51959: inst = 32'hca0cafb;
      51960: inst = 32'h13e00001;
      51961: inst = 32'hfe0d96a;
      51962: inst = 32'h5be00000;
      51963: inst = 32'h8c50000;
      51964: inst = 32'h24612800;
      51965: inst = 32'h10a0ffff;
      51966: inst = 32'hca0ffec;
      51967: inst = 32'h24822800;
      51968: inst = 32'h10a00000;
      51969: inst = 32'hca00004;
      51970: inst = 32'h38632800;
      51971: inst = 32'h38842800;
      51972: inst = 32'h10a00000;
      51973: inst = 32'hca0cb09;
      51974: inst = 32'h13e00001;
      51975: inst = 32'hfe0d96a;
      51976: inst = 32'h5be00000;
      51977: inst = 32'h8c50000;
      51978: inst = 32'h24612800;
      51979: inst = 32'h10a0ffff;
      51980: inst = 32'hca0ffec;
      51981: inst = 32'h24822800;
      51982: inst = 32'h10a00000;
      51983: inst = 32'hca00004;
      51984: inst = 32'h38632800;
      51985: inst = 32'h38842800;
      51986: inst = 32'h10a00000;
      51987: inst = 32'hca0cb17;
      51988: inst = 32'h13e00001;
      51989: inst = 32'hfe0d96a;
      51990: inst = 32'h5be00000;
      51991: inst = 32'h8c50000;
      51992: inst = 32'h24612800;
      51993: inst = 32'h10a0ffff;
      51994: inst = 32'hca0ffec;
      51995: inst = 32'h24822800;
      51996: inst = 32'h10a00000;
      51997: inst = 32'hca00004;
      51998: inst = 32'h38632800;
      51999: inst = 32'h38842800;
      52000: inst = 32'h10a00000;
      52001: inst = 32'hca0cb25;
      52002: inst = 32'h13e00001;
      52003: inst = 32'hfe0d96a;
      52004: inst = 32'h5be00000;
      52005: inst = 32'h8c50000;
      52006: inst = 32'h24612800;
      52007: inst = 32'h10a0ffff;
      52008: inst = 32'hca0ffec;
      52009: inst = 32'h24822800;
      52010: inst = 32'h10a00000;
      52011: inst = 32'hca00004;
      52012: inst = 32'h38632800;
      52013: inst = 32'h38842800;
      52014: inst = 32'h10a00000;
      52015: inst = 32'hca0cb33;
      52016: inst = 32'h13e00001;
      52017: inst = 32'hfe0d96a;
      52018: inst = 32'h5be00000;
      52019: inst = 32'h8c50000;
      52020: inst = 32'h24612800;
      52021: inst = 32'h10a0ffff;
      52022: inst = 32'hca0ffec;
      52023: inst = 32'h24822800;
      52024: inst = 32'h10a00000;
      52025: inst = 32'hca00004;
      52026: inst = 32'h38632800;
      52027: inst = 32'h38842800;
      52028: inst = 32'h10a00000;
      52029: inst = 32'hca0cb41;
      52030: inst = 32'h13e00001;
      52031: inst = 32'hfe0d96a;
      52032: inst = 32'h5be00000;
      52033: inst = 32'h8c50000;
      52034: inst = 32'h24612800;
      52035: inst = 32'h10a0ffff;
      52036: inst = 32'hca0ffec;
      52037: inst = 32'h24822800;
      52038: inst = 32'h10a00000;
      52039: inst = 32'hca00004;
      52040: inst = 32'h38632800;
      52041: inst = 32'h38842800;
      52042: inst = 32'h10a00000;
      52043: inst = 32'hca0cb4f;
      52044: inst = 32'h13e00001;
      52045: inst = 32'hfe0d96a;
      52046: inst = 32'h5be00000;
      52047: inst = 32'h8c50000;
      52048: inst = 32'h24612800;
      52049: inst = 32'h10a0ffff;
      52050: inst = 32'hca0ffec;
      52051: inst = 32'h24822800;
      52052: inst = 32'h10a00000;
      52053: inst = 32'hca00004;
      52054: inst = 32'h38632800;
      52055: inst = 32'h38842800;
      52056: inst = 32'h10a00000;
      52057: inst = 32'hca0cb5d;
      52058: inst = 32'h13e00001;
      52059: inst = 32'hfe0d96a;
      52060: inst = 32'h5be00000;
      52061: inst = 32'h8c50000;
      52062: inst = 32'h24612800;
      52063: inst = 32'h10a0ffff;
      52064: inst = 32'hca0ffec;
      52065: inst = 32'h24822800;
      52066: inst = 32'h10a00000;
      52067: inst = 32'hca00004;
      52068: inst = 32'h38632800;
      52069: inst = 32'h38842800;
      52070: inst = 32'h10a00000;
      52071: inst = 32'hca0cb6b;
      52072: inst = 32'h13e00001;
      52073: inst = 32'hfe0d96a;
      52074: inst = 32'h5be00000;
      52075: inst = 32'h8c50000;
      52076: inst = 32'h24612800;
      52077: inst = 32'h10a0ffff;
      52078: inst = 32'hca0ffec;
      52079: inst = 32'h24822800;
      52080: inst = 32'h10a00000;
      52081: inst = 32'hca00004;
      52082: inst = 32'h38632800;
      52083: inst = 32'h38842800;
      52084: inst = 32'h10a00000;
      52085: inst = 32'hca0cb79;
      52086: inst = 32'h13e00001;
      52087: inst = 32'hfe0d96a;
      52088: inst = 32'h5be00000;
      52089: inst = 32'h8c50000;
      52090: inst = 32'h24612800;
      52091: inst = 32'h10a0ffff;
      52092: inst = 32'hca0ffec;
      52093: inst = 32'h24822800;
      52094: inst = 32'h10a00000;
      52095: inst = 32'hca00004;
      52096: inst = 32'h38632800;
      52097: inst = 32'h38842800;
      52098: inst = 32'h10a00000;
      52099: inst = 32'hca0cb87;
      52100: inst = 32'h13e00001;
      52101: inst = 32'hfe0d96a;
      52102: inst = 32'h5be00000;
      52103: inst = 32'h8c50000;
      52104: inst = 32'h24612800;
      52105: inst = 32'h10a0ffff;
      52106: inst = 32'hca0ffec;
      52107: inst = 32'h24822800;
      52108: inst = 32'h10a00000;
      52109: inst = 32'hca00004;
      52110: inst = 32'h38632800;
      52111: inst = 32'h38842800;
      52112: inst = 32'h10a00000;
      52113: inst = 32'hca0cb95;
      52114: inst = 32'h13e00001;
      52115: inst = 32'hfe0d96a;
      52116: inst = 32'h5be00000;
      52117: inst = 32'h8c50000;
      52118: inst = 32'h24612800;
      52119: inst = 32'h10a0ffff;
      52120: inst = 32'hca0ffec;
      52121: inst = 32'h24822800;
      52122: inst = 32'h10a00000;
      52123: inst = 32'hca00004;
      52124: inst = 32'h38632800;
      52125: inst = 32'h38842800;
      52126: inst = 32'h10a00000;
      52127: inst = 32'hca0cba3;
      52128: inst = 32'h13e00001;
      52129: inst = 32'hfe0d96a;
      52130: inst = 32'h5be00000;
      52131: inst = 32'h8c50000;
      52132: inst = 32'h24612800;
      52133: inst = 32'h10a0ffff;
      52134: inst = 32'hca0ffec;
      52135: inst = 32'h24822800;
      52136: inst = 32'h10a00000;
      52137: inst = 32'hca00004;
      52138: inst = 32'h38632800;
      52139: inst = 32'h38842800;
      52140: inst = 32'h10a00000;
      52141: inst = 32'hca0cbb1;
      52142: inst = 32'h13e00001;
      52143: inst = 32'hfe0d96a;
      52144: inst = 32'h5be00000;
      52145: inst = 32'h8c50000;
      52146: inst = 32'h24612800;
      52147: inst = 32'h10a0ffff;
      52148: inst = 32'hca0ffec;
      52149: inst = 32'h24822800;
      52150: inst = 32'h10a00000;
      52151: inst = 32'hca00004;
      52152: inst = 32'h38632800;
      52153: inst = 32'h38842800;
      52154: inst = 32'h10a00000;
      52155: inst = 32'hca0cbbf;
      52156: inst = 32'h13e00001;
      52157: inst = 32'hfe0d96a;
      52158: inst = 32'h5be00000;
      52159: inst = 32'h8c50000;
      52160: inst = 32'h24612800;
      52161: inst = 32'h10a0ffff;
      52162: inst = 32'hca0ffec;
      52163: inst = 32'h24822800;
      52164: inst = 32'h10a00000;
      52165: inst = 32'hca00004;
      52166: inst = 32'h38632800;
      52167: inst = 32'h38842800;
      52168: inst = 32'h10a00000;
      52169: inst = 32'hca0cbcd;
      52170: inst = 32'h13e00001;
      52171: inst = 32'hfe0d96a;
      52172: inst = 32'h5be00000;
      52173: inst = 32'h8c50000;
      52174: inst = 32'h24612800;
      52175: inst = 32'h10a0ffff;
      52176: inst = 32'hca0ffec;
      52177: inst = 32'h24822800;
      52178: inst = 32'h10a00000;
      52179: inst = 32'hca00004;
      52180: inst = 32'h38632800;
      52181: inst = 32'h38842800;
      52182: inst = 32'h10a00000;
      52183: inst = 32'hca0cbdb;
      52184: inst = 32'h13e00001;
      52185: inst = 32'hfe0d96a;
      52186: inst = 32'h5be00000;
      52187: inst = 32'h8c50000;
      52188: inst = 32'h24612800;
      52189: inst = 32'h10a0ffff;
      52190: inst = 32'hca0ffec;
      52191: inst = 32'h24822800;
      52192: inst = 32'h10a00000;
      52193: inst = 32'hca00004;
      52194: inst = 32'h38632800;
      52195: inst = 32'h38842800;
      52196: inst = 32'h10a00000;
      52197: inst = 32'hca0cbe9;
      52198: inst = 32'h13e00001;
      52199: inst = 32'hfe0d96a;
      52200: inst = 32'h5be00000;
      52201: inst = 32'h8c50000;
      52202: inst = 32'h24612800;
      52203: inst = 32'h10a0ffff;
      52204: inst = 32'hca0ffec;
      52205: inst = 32'h24822800;
      52206: inst = 32'h10a00000;
      52207: inst = 32'hca00004;
      52208: inst = 32'h38632800;
      52209: inst = 32'h38842800;
      52210: inst = 32'h10a00000;
      52211: inst = 32'hca0cbf7;
      52212: inst = 32'h13e00001;
      52213: inst = 32'hfe0d96a;
      52214: inst = 32'h5be00000;
      52215: inst = 32'h8c50000;
      52216: inst = 32'h24612800;
      52217: inst = 32'h10a0ffff;
      52218: inst = 32'hca0ffec;
      52219: inst = 32'h24822800;
      52220: inst = 32'h10a00000;
      52221: inst = 32'hca00004;
      52222: inst = 32'h38632800;
      52223: inst = 32'h38842800;
      52224: inst = 32'h10a00000;
      52225: inst = 32'hca0cc05;
      52226: inst = 32'h13e00001;
      52227: inst = 32'hfe0d96a;
      52228: inst = 32'h5be00000;
      52229: inst = 32'h8c50000;
      52230: inst = 32'h24612800;
      52231: inst = 32'h10a0ffff;
      52232: inst = 32'hca0ffec;
      52233: inst = 32'h24822800;
      52234: inst = 32'h10a00000;
      52235: inst = 32'hca00004;
      52236: inst = 32'h38632800;
      52237: inst = 32'h38842800;
      52238: inst = 32'h10a00000;
      52239: inst = 32'hca0cc13;
      52240: inst = 32'h13e00001;
      52241: inst = 32'hfe0d96a;
      52242: inst = 32'h5be00000;
      52243: inst = 32'h8c50000;
      52244: inst = 32'h24612800;
      52245: inst = 32'h10a0ffff;
      52246: inst = 32'hca0ffec;
      52247: inst = 32'h24822800;
      52248: inst = 32'h10a00000;
      52249: inst = 32'hca00004;
      52250: inst = 32'h38632800;
      52251: inst = 32'h38842800;
      52252: inst = 32'h10a00000;
      52253: inst = 32'hca0cc21;
      52254: inst = 32'h13e00001;
      52255: inst = 32'hfe0d96a;
      52256: inst = 32'h5be00000;
      52257: inst = 32'h8c50000;
      52258: inst = 32'h24612800;
      52259: inst = 32'h10a0ffff;
      52260: inst = 32'hca0ffec;
      52261: inst = 32'h24822800;
      52262: inst = 32'h10a00000;
      52263: inst = 32'hca00004;
      52264: inst = 32'h38632800;
      52265: inst = 32'h38842800;
      52266: inst = 32'h10a00000;
      52267: inst = 32'hca0cc2f;
      52268: inst = 32'h13e00001;
      52269: inst = 32'hfe0d96a;
      52270: inst = 32'h5be00000;
      52271: inst = 32'h8c50000;
      52272: inst = 32'h24612800;
      52273: inst = 32'h10a0ffff;
      52274: inst = 32'hca0ffec;
      52275: inst = 32'h24822800;
      52276: inst = 32'h10a00000;
      52277: inst = 32'hca00004;
      52278: inst = 32'h38632800;
      52279: inst = 32'h38842800;
      52280: inst = 32'h10a00000;
      52281: inst = 32'hca0cc3d;
      52282: inst = 32'h13e00001;
      52283: inst = 32'hfe0d96a;
      52284: inst = 32'h5be00000;
      52285: inst = 32'h8c50000;
      52286: inst = 32'h24612800;
      52287: inst = 32'h10a0ffff;
      52288: inst = 32'hca0ffec;
      52289: inst = 32'h24822800;
      52290: inst = 32'h10a00000;
      52291: inst = 32'hca00004;
      52292: inst = 32'h38632800;
      52293: inst = 32'h38842800;
      52294: inst = 32'h10a00000;
      52295: inst = 32'hca0cc4b;
      52296: inst = 32'h13e00001;
      52297: inst = 32'hfe0d96a;
      52298: inst = 32'h5be00000;
      52299: inst = 32'h8c50000;
      52300: inst = 32'h24612800;
      52301: inst = 32'h10a0ffff;
      52302: inst = 32'hca0ffec;
      52303: inst = 32'h24822800;
      52304: inst = 32'h10a00000;
      52305: inst = 32'hca00004;
      52306: inst = 32'h38632800;
      52307: inst = 32'h38842800;
      52308: inst = 32'h10a00000;
      52309: inst = 32'hca0cc59;
      52310: inst = 32'h13e00001;
      52311: inst = 32'hfe0d96a;
      52312: inst = 32'h5be00000;
      52313: inst = 32'h8c50000;
      52314: inst = 32'h24612800;
      52315: inst = 32'h10a0ffff;
      52316: inst = 32'hca0ffec;
      52317: inst = 32'h24822800;
      52318: inst = 32'h10a00000;
      52319: inst = 32'hca00004;
      52320: inst = 32'h38632800;
      52321: inst = 32'h38842800;
      52322: inst = 32'h10a00000;
      52323: inst = 32'hca0cc67;
      52324: inst = 32'h13e00001;
      52325: inst = 32'hfe0d96a;
      52326: inst = 32'h5be00000;
      52327: inst = 32'h8c50000;
      52328: inst = 32'h24612800;
      52329: inst = 32'h10a0ffff;
      52330: inst = 32'hca0ffec;
      52331: inst = 32'h24822800;
      52332: inst = 32'h10a00000;
      52333: inst = 32'hca00004;
      52334: inst = 32'h38632800;
      52335: inst = 32'h38842800;
      52336: inst = 32'h10a00000;
      52337: inst = 32'hca0cc75;
      52338: inst = 32'h13e00001;
      52339: inst = 32'hfe0d96a;
      52340: inst = 32'h5be00000;
      52341: inst = 32'h8c50000;
      52342: inst = 32'h24612800;
      52343: inst = 32'h10a0ffff;
      52344: inst = 32'hca0ffec;
      52345: inst = 32'h24822800;
      52346: inst = 32'h10a00000;
      52347: inst = 32'hca00004;
      52348: inst = 32'h38632800;
      52349: inst = 32'h38842800;
      52350: inst = 32'h10a00000;
      52351: inst = 32'hca0cc83;
      52352: inst = 32'h13e00001;
      52353: inst = 32'hfe0d96a;
      52354: inst = 32'h5be00000;
      52355: inst = 32'h8c50000;
      52356: inst = 32'h24612800;
      52357: inst = 32'h10a0ffff;
      52358: inst = 32'hca0ffec;
      52359: inst = 32'h24822800;
      52360: inst = 32'h10a00000;
      52361: inst = 32'hca00004;
      52362: inst = 32'h38632800;
      52363: inst = 32'h38842800;
      52364: inst = 32'h10a00000;
      52365: inst = 32'hca0cc91;
      52366: inst = 32'h13e00001;
      52367: inst = 32'hfe0d96a;
      52368: inst = 32'h5be00000;
      52369: inst = 32'h8c50000;
      52370: inst = 32'h24612800;
      52371: inst = 32'h10a0ffff;
      52372: inst = 32'hca0ffec;
      52373: inst = 32'h24822800;
      52374: inst = 32'h10a00000;
      52375: inst = 32'hca00004;
      52376: inst = 32'h38632800;
      52377: inst = 32'h38842800;
      52378: inst = 32'h10a00000;
      52379: inst = 32'hca0cc9f;
      52380: inst = 32'h13e00001;
      52381: inst = 32'hfe0d96a;
      52382: inst = 32'h5be00000;
      52383: inst = 32'h8c50000;
      52384: inst = 32'h24612800;
      52385: inst = 32'h10a0ffff;
      52386: inst = 32'hca0ffec;
      52387: inst = 32'h24822800;
      52388: inst = 32'h10a00000;
      52389: inst = 32'hca00004;
      52390: inst = 32'h38632800;
      52391: inst = 32'h38842800;
      52392: inst = 32'h10a00000;
      52393: inst = 32'hca0ccad;
      52394: inst = 32'h13e00001;
      52395: inst = 32'hfe0d96a;
      52396: inst = 32'h5be00000;
      52397: inst = 32'h8c50000;
      52398: inst = 32'h24612800;
      52399: inst = 32'h10a0ffff;
      52400: inst = 32'hca0ffec;
      52401: inst = 32'h24822800;
      52402: inst = 32'h10a00000;
      52403: inst = 32'hca00004;
      52404: inst = 32'h38632800;
      52405: inst = 32'h38842800;
      52406: inst = 32'h10a00000;
      52407: inst = 32'hca0ccbb;
      52408: inst = 32'h13e00001;
      52409: inst = 32'hfe0d96a;
      52410: inst = 32'h5be00000;
      52411: inst = 32'h8c50000;
      52412: inst = 32'h24612800;
      52413: inst = 32'h10a0ffff;
      52414: inst = 32'hca0ffec;
      52415: inst = 32'h24822800;
      52416: inst = 32'h10a00000;
      52417: inst = 32'hca00004;
      52418: inst = 32'h38632800;
      52419: inst = 32'h38842800;
      52420: inst = 32'h10a00000;
      52421: inst = 32'hca0ccc9;
      52422: inst = 32'h13e00001;
      52423: inst = 32'hfe0d96a;
      52424: inst = 32'h5be00000;
      52425: inst = 32'h8c50000;
      52426: inst = 32'h24612800;
      52427: inst = 32'h10a0ffff;
      52428: inst = 32'hca0ffec;
      52429: inst = 32'h24822800;
      52430: inst = 32'h10a00000;
      52431: inst = 32'hca00004;
      52432: inst = 32'h38632800;
      52433: inst = 32'h38842800;
      52434: inst = 32'h10a00000;
      52435: inst = 32'hca0ccd7;
      52436: inst = 32'h13e00001;
      52437: inst = 32'hfe0d96a;
      52438: inst = 32'h5be00000;
      52439: inst = 32'h8c50000;
      52440: inst = 32'h24612800;
      52441: inst = 32'h10a0ffff;
      52442: inst = 32'hca0ffec;
      52443: inst = 32'h24822800;
      52444: inst = 32'h10a00000;
      52445: inst = 32'hca00004;
      52446: inst = 32'h38632800;
      52447: inst = 32'h38842800;
      52448: inst = 32'h10a00000;
      52449: inst = 32'hca0cce5;
      52450: inst = 32'h13e00001;
      52451: inst = 32'hfe0d96a;
      52452: inst = 32'h5be00000;
      52453: inst = 32'h8c50000;
      52454: inst = 32'h24612800;
      52455: inst = 32'h10a0ffff;
      52456: inst = 32'hca0ffec;
      52457: inst = 32'h24822800;
      52458: inst = 32'h10a00000;
      52459: inst = 32'hca00004;
      52460: inst = 32'h38632800;
      52461: inst = 32'h38842800;
      52462: inst = 32'h10a00000;
      52463: inst = 32'hca0ccf3;
      52464: inst = 32'h13e00001;
      52465: inst = 32'hfe0d96a;
      52466: inst = 32'h5be00000;
      52467: inst = 32'h8c50000;
      52468: inst = 32'h24612800;
      52469: inst = 32'h10a0ffff;
      52470: inst = 32'hca0ffec;
      52471: inst = 32'h24822800;
      52472: inst = 32'h10a00000;
      52473: inst = 32'hca00004;
      52474: inst = 32'h38632800;
      52475: inst = 32'h38842800;
      52476: inst = 32'h10a00000;
      52477: inst = 32'hca0cd01;
      52478: inst = 32'h13e00001;
      52479: inst = 32'hfe0d96a;
      52480: inst = 32'h5be00000;
      52481: inst = 32'h8c50000;
      52482: inst = 32'h24612800;
      52483: inst = 32'h10a0ffff;
      52484: inst = 32'hca0ffec;
      52485: inst = 32'h24822800;
      52486: inst = 32'h10a00000;
      52487: inst = 32'hca00004;
      52488: inst = 32'h38632800;
      52489: inst = 32'h38842800;
      52490: inst = 32'h10a00000;
      52491: inst = 32'hca0cd0f;
      52492: inst = 32'h13e00001;
      52493: inst = 32'hfe0d96a;
      52494: inst = 32'h5be00000;
      52495: inst = 32'h8c50000;
      52496: inst = 32'h24612800;
      52497: inst = 32'h10a0ffff;
      52498: inst = 32'hca0ffec;
      52499: inst = 32'h24822800;
      52500: inst = 32'h10a00000;
      52501: inst = 32'hca00004;
      52502: inst = 32'h38632800;
      52503: inst = 32'h38842800;
      52504: inst = 32'h10a00000;
      52505: inst = 32'hca0cd1d;
      52506: inst = 32'h13e00001;
      52507: inst = 32'hfe0d96a;
      52508: inst = 32'h5be00000;
      52509: inst = 32'h8c50000;
      52510: inst = 32'h24612800;
      52511: inst = 32'h10a0ffff;
      52512: inst = 32'hca0ffec;
      52513: inst = 32'h24822800;
      52514: inst = 32'h10a00000;
      52515: inst = 32'hca00004;
      52516: inst = 32'h38632800;
      52517: inst = 32'h38842800;
      52518: inst = 32'h10a00000;
      52519: inst = 32'hca0cd2b;
      52520: inst = 32'h13e00001;
      52521: inst = 32'hfe0d96a;
      52522: inst = 32'h5be00000;
      52523: inst = 32'h8c50000;
      52524: inst = 32'h24612800;
      52525: inst = 32'h10a0ffff;
      52526: inst = 32'hca0ffec;
      52527: inst = 32'h24822800;
      52528: inst = 32'h10a00000;
      52529: inst = 32'hca00004;
      52530: inst = 32'h38632800;
      52531: inst = 32'h38842800;
      52532: inst = 32'h10a00000;
      52533: inst = 32'hca0cd39;
      52534: inst = 32'h13e00001;
      52535: inst = 32'hfe0d96a;
      52536: inst = 32'h5be00000;
      52537: inst = 32'h8c50000;
      52538: inst = 32'h24612800;
      52539: inst = 32'h10a0ffff;
      52540: inst = 32'hca0ffec;
      52541: inst = 32'h24822800;
      52542: inst = 32'h10a00000;
      52543: inst = 32'hca00004;
      52544: inst = 32'h38632800;
      52545: inst = 32'h38842800;
      52546: inst = 32'h10a00000;
      52547: inst = 32'hca0cd47;
      52548: inst = 32'h13e00001;
      52549: inst = 32'hfe0d96a;
      52550: inst = 32'h5be00000;
      52551: inst = 32'h8c50000;
      52552: inst = 32'h24612800;
      52553: inst = 32'h10a0ffff;
      52554: inst = 32'hca0ffec;
      52555: inst = 32'h24822800;
      52556: inst = 32'h10a00000;
      52557: inst = 32'hca00004;
      52558: inst = 32'h38632800;
      52559: inst = 32'h38842800;
      52560: inst = 32'h10a00000;
      52561: inst = 32'hca0cd55;
      52562: inst = 32'h13e00001;
      52563: inst = 32'hfe0d96a;
      52564: inst = 32'h5be00000;
      52565: inst = 32'h8c50000;
      52566: inst = 32'h24612800;
      52567: inst = 32'h10a0ffff;
      52568: inst = 32'hca0ffec;
      52569: inst = 32'h24822800;
      52570: inst = 32'h10a00000;
      52571: inst = 32'hca00004;
      52572: inst = 32'h38632800;
      52573: inst = 32'h38842800;
      52574: inst = 32'h10a00000;
      52575: inst = 32'hca0cd63;
      52576: inst = 32'h13e00001;
      52577: inst = 32'hfe0d96a;
      52578: inst = 32'h5be00000;
      52579: inst = 32'h8c50000;
      52580: inst = 32'h24612800;
      52581: inst = 32'h10a0ffff;
      52582: inst = 32'hca0ffec;
      52583: inst = 32'h24822800;
      52584: inst = 32'h10a00000;
      52585: inst = 32'hca00004;
      52586: inst = 32'h38632800;
      52587: inst = 32'h38842800;
      52588: inst = 32'h10a00000;
      52589: inst = 32'hca0cd71;
      52590: inst = 32'h13e00001;
      52591: inst = 32'hfe0d96a;
      52592: inst = 32'h5be00000;
      52593: inst = 32'h8c50000;
      52594: inst = 32'h24612800;
      52595: inst = 32'h10a0ffff;
      52596: inst = 32'hca0ffec;
      52597: inst = 32'h24822800;
      52598: inst = 32'h10a00000;
      52599: inst = 32'hca00004;
      52600: inst = 32'h38632800;
      52601: inst = 32'h38842800;
      52602: inst = 32'h10a00000;
      52603: inst = 32'hca0cd7f;
      52604: inst = 32'h13e00001;
      52605: inst = 32'hfe0d96a;
      52606: inst = 32'h5be00000;
      52607: inst = 32'h8c50000;
      52608: inst = 32'h24612800;
      52609: inst = 32'h10a0ffff;
      52610: inst = 32'hca0ffec;
      52611: inst = 32'h24822800;
      52612: inst = 32'h10a00000;
      52613: inst = 32'hca00004;
      52614: inst = 32'h38632800;
      52615: inst = 32'h38842800;
      52616: inst = 32'h10a00000;
      52617: inst = 32'hca0cd8d;
      52618: inst = 32'h13e00001;
      52619: inst = 32'hfe0d96a;
      52620: inst = 32'h5be00000;
      52621: inst = 32'h8c50000;
      52622: inst = 32'h24612800;
      52623: inst = 32'h10a0ffff;
      52624: inst = 32'hca0ffec;
      52625: inst = 32'h24822800;
      52626: inst = 32'h10a00000;
      52627: inst = 32'hca00004;
      52628: inst = 32'h38632800;
      52629: inst = 32'h38842800;
      52630: inst = 32'h10a00000;
      52631: inst = 32'hca0cd9b;
      52632: inst = 32'h13e00001;
      52633: inst = 32'hfe0d96a;
      52634: inst = 32'h5be00000;
      52635: inst = 32'h8c50000;
      52636: inst = 32'h24612800;
      52637: inst = 32'h10a0ffff;
      52638: inst = 32'hca0ffec;
      52639: inst = 32'h24822800;
      52640: inst = 32'h10a00000;
      52641: inst = 32'hca00004;
      52642: inst = 32'h38632800;
      52643: inst = 32'h38842800;
      52644: inst = 32'h10a00000;
      52645: inst = 32'hca0cda9;
      52646: inst = 32'h13e00001;
      52647: inst = 32'hfe0d96a;
      52648: inst = 32'h5be00000;
      52649: inst = 32'h8c50000;
      52650: inst = 32'h24612800;
      52651: inst = 32'h10a0ffff;
      52652: inst = 32'hca0ffed;
      52653: inst = 32'h24822800;
      52654: inst = 32'h10a00000;
      52655: inst = 32'hca00004;
      52656: inst = 32'h38632800;
      52657: inst = 32'h38842800;
      52658: inst = 32'h10a00000;
      52659: inst = 32'hca0cdb7;
      52660: inst = 32'h13e00001;
      52661: inst = 32'hfe0d96a;
      52662: inst = 32'h5be00000;
      52663: inst = 32'h8c50000;
      52664: inst = 32'h24612800;
      52665: inst = 32'h10a0ffff;
      52666: inst = 32'hca0ffed;
      52667: inst = 32'h24822800;
      52668: inst = 32'h10a00000;
      52669: inst = 32'hca00004;
      52670: inst = 32'h38632800;
      52671: inst = 32'h38842800;
      52672: inst = 32'h10a00000;
      52673: inst = 32'hca0cdc5;
      52674: inst = 32'h13e00001;
      52675: inst = 32'hfe0d96a;
      52676: inst = 32'h5be00000;
      52677: inst = 32'h8c50000;
      52678: inst = 32'h24612800;
      52679: inst = 32'h10a0ffff;
      52680: inst = 32'hca0ffed;
      52681: inst = 32'h24822800;
      52682: inst = 32'h10a00000;
      52683: inst = 32'hca00004;
      52684: inst = 32'h38632800;
      52685: inst = 32'h38842800;
      52686: inst = 32'h10a00000;
      52687: inst = 32'hca0cdd3;
      52688: inst = 32'h13e00001;
      52689: inst = 32'hfe0d96a;
      52690: inst = 32'h5be00000;
      52691: inst = 32'h8c50000;
      52692: inst = 32'h24612800;
      52693: inst = 32'h10a0ffff;
      52694: inst = 32'hca0ffed;
      52695: inst = 32'h24822800;
      52696: inst = 32'h10a00000;
      52697: inst = 32'hca00004;
      52698: inst = 32'h38632800;
      52699: inst = 32'h38842800;
      52700: inst = 32'h10a00000;
      52701: inst = 32'hca0cde1;
      52702: inst = 32'h13e00001;
      52703: inst = 32'hfe0d96a;
      52704: inst = 32'h5be00000;
      52705: inst = 32'h8c50000;
      52706: inst = 32'h24612800;
      52707: inst = 32'h10a0ffff;
      52708: inst = 32'hca0ffed;
      52709: inst = 32'h24822800;
      52710: inst = 32'h10a00000;
      52711: inst = 32'hca00004;
      52712: inst = 32'h38632800;
      52713: inst = 32'h38842800;
      52714: inst = 32'h10a00000;
      52715: inst = 32'hca0cdef;
      52716: inst = 32'h13e00001;
      52717: inst = 32'hfe0d96a;
      52718: inst = 32'h5be00000;
      52719: inst = 32'h8c50000;
      52720: inst = 32'h24612800;
      52721: inst = 32'h10a0ffff;
      52722: inst = 32'hca0ffed;
      52723: inst = 32'h24822800;
      52724: inst = 32'h10a00000;
      52725: inst = 32'hca00004;
      52726: inst = 32'h38632800;
      52727: inst = 32'h38842800;
      52728: inst = 32'h10a00000;
      52729: inst = 32'hca0cdfd;
      52730: inst = 32'h13e00001;
      52731: inst = 32'hfe0d96a;
      52732: inst = 32'h5be00000;
      52733: inst = 32'h8c50000;
      52734: inst = 32'h24612800;
      52735: inst = 32'h10a0ffff;
      52736: inst = 32'hca0ffed;
      52737: inst = 32'h24822800;
      52738: inst = 32'h10a00000;
      52739: inst = 32'hca00004;
      52740: inst = 32'h38632800;
      52741: inst = 32'h38842800;
      52742: inst = 32'h10a00000;
      52743: inst = 32'hca0ce0b;
      52744: inst = 32'h13e00001;
      52745: inst = 32'hfe0d96a;
      52746: inst = 32'h5be00000;
      52747: inst = 32'h8c50000;
      52748: inst = 32'h24612800;
      52749: inst = 32'h10a0ffff;
      52750: inst = 32'hca0ffed;
      52751: inst = 32'h24822800;
      52752: inst = 32'h10a00000;
      52753: inst = 32'hca00004;
      52754: inst = 32'h38632800;
      52755: inst = 32'h38842800;
      52756: inst = 32'h10a00000;
      52757: inst = 32'hca0ce19;
      52758: inst = 32'h13e00001;
      52759: inst = 32'hfe0d96a;
      52760: inst = 32'h5be00000;
      52761: inst = 32'h8c50000;
      52762: inst = 32'h24612800;
      52763: inst = 32'h10a0ffff;
      52764: inst = 32'hca0ffed;
      52765: inst = 32'h24822800;
      52766: inst = 32'h10a00000;
      52767: inst = 32'hca00004;
      52768: inst = 32'h38632800;
      52769: inst = 32'h38842800;
      52770: inst = 32'h10a00000;
      52771: inst = 32'hca0ce27;
      52772: inst = 32'h13e00001;
      52773: inst = 32'hfe0d96a;
      52774: inst = 32'h5be00000;
      52775: inst = 32'h8c50000;
      52776: inst = 32'h24612800;
      52777: inst = 32'h10a0ffff;
      52778: inst = 32'hca0ffed;
      52779: inst = 32'h24822800;
      52780: inst = 32'h10a00000;
      52781: inst = 32'hca00004;
      52782: inst = 32'h38632800;
      52783: inst = 32'h38842800;
      52784: inst = 32'h10a00000;
      52785: inst = 32'hca0ce35;
      52786: inst = 32'h13e00001;
      52787: inst = 32'hfe0d96a;
      52788: inst = 32'h5be00000;
      52789: inst = 32'h8c50000;
      52790: inst = 32'h24612800;
      52791: inst = 32'h10a0ffff;
      52792: inst = 32'hca0ffed;
      52793: inst = 32'h24822800;
      52794: inst = 32'h10a00000;
      52795: inst = 32'hca00004;
      52796: inst = 32'h38632800;
      52797: inst = 32'h38842800;
      52798: inst = 32'h10a00000;
      52799: inst = 32'hca0ce43;
      52800: inst = 32'h13e00001;
      52801: inst = 32'hfe0d96a;
      52802: inst = 32'h5be00000;
      52803: inst = 32'h8c50000;
      52804: inst = 32'h24612800;
      52805: inst = 32'h10a0ffff;
      52806: inst = 32'hca0ffed;
      52807: inst = 32'h24822800;
      52808: inst = 32'h10a00000;
      52809: inst = 32'hca00004;
      52810: inst = 32'h38632800;
      52811: inst = 32'h38842800;
      52812: inst = 32'h10a00000;
      52813: inst = 32'hca0ce51;
      52814: inst = 32'h13e00001;
      52815: inst = 32'hfe0d96a;
      52816: inst = 32'h5be00000;
      52817: inst = 32'h8c50000;
      52818: inst = 32'h24612800;
      52819: inst = 32'h10a0ffff;
      52820: inst = 32'hca0ffed;
      52821: inst = 32'h24822800;
      52822: inst = 32'h10a00000;
      52823: inst = 32'hca00004;
      52824: inst = 32'h38632800;
      52825: inst = 32'h38842800;
      52826: inst = 32'h10a00000;
      52827: inst = 32'hca0ce5f;
      52828: inst = 32'h13e00001;
      52829: inst = 32'hfe0d96a;
      52830: inst = 32'h5be00000;
      52831: inst = 32'h8c50000;
      52832: inst = 32'h24612800;
      52833: inst = 32'h10a0ffff;
      52834: inst = 32'hca0ffed;
      52835: inst = 32'h24822800;
      52836: inst = 32'h10a00000;
      52837: inst = 32'hca00004;
      52838: inst = 32'h38632800;
      52839: inst = 32'h38842800;
      52840: inst = 32'h10a00000;
      52841: inst = 32'hca0ce6d;
      52842: inst = 32'h13e00001;
      52843: inst = 32'hfe0d96a;
      52844: inst = 32'h5be00000;
      52845: inst = 32'h8c50000;
      52846: inst = 32'h24612800;
      52847: inst = 32'h10a0ffff;
      52848: inst = 32'hca0ffed;
      52849: inst = 32'h24822800;
      52850: inst = 32'h10a00000;
      52851: inst = 32'hca00004;
      52852: inst = 32'h38632800;
      52853: inst = 32'h38842800;
      52854: inst = 32'h10a00000;
      52855: inst = 32'hca0ce7b;
      52856: inst = 32'h13e00001;
      52857: inst = 32'hfe0d96a;
      52858: inst = 32'h5be00000;
      52859: inst = 32'h8c50000;
      52860: inst = 32'h24612800;
      52861: inst = 32'h10a0ffff;
      52862: inst = 32'hca0ffed;
      52863: inst = 32'h24822800;
      52864: inst = 32'h10a00000;
      52865: inst = 32'hca00004;
      52866: inst = 32'h38632800;
      52867: inst = 32'h38842800;
      52868: inst = 32'h10a00000;
      52869: inst = 32'hca0ce89;
      52870: inst = 32'h13e00001;
      52871: inst = 32'hfe0d96a;
      52872: inst = 32'h5be00000;
      52873: inst = 32'h8c50000;
      52874: inst = 32'h24612800;
      52875: inst = 32'h10a0ffff;
      52876: inst = 32'hca0ffed;
      52877: inst = 32'h24822800;
      52878: inst = 32'h10a00000;
      52879: inst = 32'hca00004;
      52880: inst = 32'h38632800;
      52881: inst = 32'h38842800;
      52882: inst = 32'h10a00000;
      52883: inst = 32'hca0ce97;
      52884: inst = 32'h13e00001;
      52885: inst = 32'hfe0d96a;
      52886: inst = 32'h5be00000;
      52887: inst = 32'h8c50000;
      52888: inst = 32'h24612800;
      52889: inst = 32'h10a0ffff;
      52890: inst = 32'hca0ffed;
      52891: inst = 32'h24822800;
      52892: inst = 32'h10a00000;
      52893: inst = 32'hca00004;
      52894: inst = 32'h38632800;
      52895: inst = 32'h38842800;
      52896: inst = 32'h10a00000;
      52897: inst = 32'hca0cea5;
      52898: inst = 32'h13e00001;
      52899: inst = 32'hfe0d96a;
      52900: inst = 32'h5be00000;
      52901: inst = 32'h8c50000;
      52902: inst = 32'h24612800;
      52903: inst = 32'h10a0ffff;
      52904: inst = 32'hca0ffed;
      52905: inst = 32'h24822800;
      52906: inst = 32'h10a00000;
      52907: inst = 32'hca00004;
      52908: inst = 32'h38632800;
      52909: inst = 32'h38842800;
      52910: inst = 32'h10a00000;
      52911: inst = 32'hca0ceb3;
      52912: inst = 32'h13e00001;
      52913: inst = 32'hfe0d96a;
      52914: inst = 32'h5be00000;
      52915: inst = 32'h8c50000;
      52916: inst = 32'h24612800;
      52917: inst = 32'h10a0ffff;
      52918: inst = 32'hca0ffed;
      52919: inst = 32'h24822800;
      52920: inst = 32'h10a00000;
      52921: inst = 32'hca00004;
      52922: inst = 32'h38632800;
      52923: inst = 32'h38842800;
      52924: inst = 32'h10a00000;
      52925: inst = 32'hca0cec1;
      52926: inst = 32'h13e00001;
      52927: inst = 32'hfe0d96a;
      52928: inst = 32'h5be00000;
      52929: inst = 32'h8c50000;
      52930: inst = 32'h24612800;
      52931: inst = 32'h10a0ffff;
      52932: inst = 32'hca0ffed;
      52933: inst = 32'h24822800;
      52934: inst = 32'h10a00000;
      52935: inst = 32'hca00004;
      52936: inst = 32'h38632800;
      52937: inst = 32'h38842800;
      52938: inst = 32'h10a00000;
      52939: inst = 32'hca0cecf;
      52940: inst = 32'h13e00001;
      52941: inst = 32'hfe0d96a;
      52942: inst = 32'h5be00000;
      52943: inst = 32'h8c50000;
      52944: inst = 32'h24612800;
      52945: inst = 32'h10a0ffff;
      52946: inst = 32'hca0ffed;
      52947: inst = 32'h24822800;
      52948: inst = 32'h10a00000;
      52949: inst = 32'hca00004;
      52950: inst = 32'h38632800;
      52951: inst = 32'h38842800;
      52952: inst = 32'h10a00000;
      52953: inst = 32'hca0cedd;
      52954: inst = 32'h13e00001;
      52955: inst = 32'hfe0d96a;
      52956: inst = 32'h5be00000;
      52957: inst = 32'h8c50000;
      52958: inst = 32'h24612800;
      52959: inst = 32'h10a0ffff;
      52960: inst = 32'hca0ffed;
      52961: inst = 32'h24822800;
      52962: inst = 32'h10a00000;
      52963: inst = 32'hca00004;
      52964: inst = 32'h38632800;
      52965: inst = 32'h38842800;
      52966: inst = 32'h10a00000;
      52967: inst = 32'hca0ceeb;
      52968: inst = 32'h13e00001;
      52969: inst = 32'hfe0d96a;
      52970: inst = 32'h5be00000;
      52971: inst = 32'h8c50000;
      52972: inst = 32'h24612800;
      52973: inst = 32'h10a0ffff;
      52974: inst = 32'hca0ffed;
      52975: inst = 32'h24822800;
      52976: inst = 32'h10a00000;
      52977: inst = 32'hca00004;
      52978: inst = 32'h38632800;
      52979: inst = 32'h38842800;
      52980: inst = 32'h10a00000;
      52981: inst = 32'hca0cef9;
      52982: inst = 32'h13e00001;
      52983: inst = 32'hfe0d96a;
      52984: inst = 32'h5be00000;
      52985: inst = 32'h8c50000;
      52986: inst = 32'h24612800;
      52987: inst = 32'h10a0ffff;
      52988: inst = 32'hca0ffed;
      52989: inst = 32'h24822800;
      52990: inst = 32'h10a00000;
      52991: inst = 32'hca00004;
      52992: inst = 32'h38632800;
      52993: inst = 32'h38842800;
      52994: inst = 32'h10a00000;
      52995: inst = 32'hca0cf07;
      52996: inst = 32'h13e00001;
      52997: inst = 32'hfe0d96a;
      52998: inst = 32'h5be00000;
      52999: inst = 32'h8c50000;
      53000: inst = 32'h24612800;
      53001: inst = 32'h10a0ffff;
      53002: inst = 32'hca0ffed;
      53003: inst = 32'h24822800;
      53004: inst = 32'h10a00000;
      53005: inst = 32'hca00004;
      53006: inst = 32'h38632800;
      53007: inst = 32'h38842800;
      53008: inst = 32'h10a00000;
      53009: inst = 32'hca0cf15;
      53010: inst = 32'h13e00001;
      53011: inst = 32'hfe0d96a;
      53012: inst = 32'h5be00000;
      53013: inst = 32'h8c50000;
      53014: inst = 32'h24612800;
      53015: inst = 32'h10a0ffff;
      53016: inst = 32'hca0ffed;
      53017: inst = 32'h24822800;
      53018: inst = 32'h10a00000;
      53019: inst = 32'hca00004;
      53020: inst = 32'h38632800;
      53021: inst = 32'h38842800;
      53022: inst = 32'h10a00000;
      53023: inst = 32'hca0cf23;
      53024: inst = 32'h13e00001;
      53025: inst = 32'hfe0d96a;
      53026: inst = 32'h5be00000;
      53027: inst = 32'h8c50000;
      53028: inst = 32'h24612800;
      53029: inst = 32'h10a0ffff;
      53030: inst = 32'hca0ffed;
      53031: inst = 32'h24822800;
      53032: inst = 32'h10a00000;
      53033: inst = 32'hca00004;
      53034: inst = 32'h38632800;
      53035: inst = 32'h38842800;
      53036: inst = 32'h10a00000;
      53037: inst = 32'hca0cf31;
      53038: inst = 32'h13e00001;
      53039: inst = 32'hfe0d96a;
      53040: inst = 32'h5be00000;
      53041: inst = 32'h8c50000;
      53042: inst = 32'h24612800;
      53043: inst = 32'h10a0ffff;
      53044: inst = 32'hca0ffed;
      53045: inst = 32'h24822800;
      53046: inst = 32'h10a00000;
      53047: inst = 32'hca00004;
      53048: inst = 32'h38632800;
      53049: inst = 32'h38842800;
      53050: inst = 32'h10a00000;
      53051: inst = 32'hca0cf3f;
      53052: inst = 32'h13e00001;
      53053: inst = 32'hfe0d96a;
      53054: inst = 32'h5be00000;
      53055: inst = 32'h8c50000;
      53056: inst = 32'h24612800;
      53057: inst = 32'h10a0ffff;
      53058: inst = 32'hca0ffed;
      53059: inst = 32'h24822800;
      53060: inst = 32'h10a00000;
      53061: inst = 32'hca00004;
      53062: inst = 32'h38632800;
      53063: inst = 32'h38842800;
      53064: inst = 32'h10a00000;
      53065: inst = 32'hca0cf4d;
      53066: inst = 32'h13e00001;
      53067: inst = 32'hfe0d96a;
      53068: inst = 32'h5be00000;
      53069: inst = 32'h8c50000;
      53070: inst = 32'h24612800;
      53071: inst = 32'h10a0ffff;
      53072: inst = 32'hca0ffed;
      53073: inst = 32'h24822800;
      53074: inst = 32'h10a00000;
      53075: inst = 32'hca00004;
      53076: inst = 32'h38632800;
      53077: inst = 32'h38842800;
      53078: inst = 32'h10a00000;
      53079: inst = 32'hca0cf5b;
      53080: inst = 32'h13e00001;
      53081: inst = 32'hfe0d96a;
      53082: inst = 32'h5be00000;
      53083: inst = 32'h8c50000;
      53084: inst = 32'h24612800;
      53085: inst = 32'h10a0ffff;
      53086: inst = 32'hca0ffed;
      53087: inst = 32'h24822800;
      53088: inst = 32'h10a00000;
      53089: inst = 32'hca00004;
      53090: inst = 32'h38632800;
      53091: inst = 32'h38842800;
      53092: inst = 32'h10a00000;
      53093: inst = 32'hca0cf69;
      53094: inst = 32'h13e00001;
      53095: inst = 32'hfe0d96a;
      53096: inst = 32'h5be00000;
      53097: inst = 32'h8c50000;
      53098: inst = 32'h24612800;
      53099: inst = 32'h10a0ffff;
      53100: inst = 32'hca0ffed;
      53101: inst = 32'h24822800;
      53102: inst = 32'h10a00000;
      53103: inst = 32'hca00004;
      53104: inst = 32'h38632800;
      53105: inst = 32'h38842800;
      53106: inst = 32'h10a00000;
      53107: inst = 32'hca0cf77;
      53108: inst = 32'h13e00001;
      53109: inst = 32'hfe0d96a;
      53110: inst = 32'h5be00000;
      53111: inst = 32'h8c50000;
      53112: inst = 32'h24612800;
      53113: inst = 32'h10a0ffff;
      53114: inst = 32'hca0ffed;
      53115: inst = 32'h24822800;
      53116: inst = 32'h10a00000;
      53117: inst = 32'hca00004;
      53118: inst = 32'h38632800;
      53119: inst = 32'h38842800;
      53120: inst = 32'h10a00000;
      53121: inst = 32'hca0cf85;
      53122: inst = 32'h13e00001;
      53123: inst = 32'hfe0d96a;
      53124: inst = 32'h5be00000;
      53125: inst = 32'h8c50000;
      53126: inst = 32'h24612800;
      53127: inst = 32'h10a0ffff;
      53128: inst = 32'hca0ffed;
      53129: inst = 32'h24822800;
      53130: inst = 32'h10a00000;
      53131: inst = 32'hca00004;
      53132: inst = 32'h38632800;
      53133: inst = 32'h38842800;
      53134: inst = 32'h10a00000;
      53135: inst = 32'hca0cf93;
      53136: inst = 32'h13e00001;
      53137: inst = 32'hfe0d96a;
      53138: inst = 32'h5be00000;
      53139: inst = 32'h8c50000;
      53140: inst = 32'h24612800;
      53141: inst = 32'h10a0ffff;
      53142: inst = 32'hca0ffed;
      53143: inst = 32'h24822800;
      53144: inst = 32'h10a00000;
      53145: inst = 32'hca00004;
      53146: inst = 32'h38632800;
      53147: inst = 32'h38842800;
      53148: inst = 32'h10a00000;
      53149: inst = 32'hca0cfa1;
      53150: inst = 32'h13e00001;
      53151: inst = 32'hfe0d96a;
      53152: inst = 32'h5be00000;
      53153: inst = 32'h8c50000;
      53154: inst = 32'h24612800;
      53155: inst = 32'h10a0ffff;
      53156: inst = 32'hca0ffed;
      53157: inst = 32'h24822800;
      53158: inst = 32'h10a00000;
      53159: inst = 32'hca00004;
      53160: inst = 32'h38632800;
      53161: inst = 32'h38842800;
      53162: inst = 32'h10a00000;
      53163: inst = 32'hca0cfaf;
      53164: inst = 32'h13e00001;
      53165: inst = 32'hfe0d96a;
      53166: inst = 32'h5be00000;
      53167: inst = 32'h8c50000;
      53168: inst = 32'h24612800;
      53169: inst = 32'h10a0ffff;
      53170: inst = 32'hca0ffed;
      53171: inst = 32'h24822800;
      53172: inst = 32'h10a00000;
      53173: inst = 32'hca00004;
      53174: inst = 32'h38632800;
      53175: inst = 32'h38842800;
      53176: inst = 32'h10a00000;
      53177: inst = 32'hca0cfbd;
      53178: inst = 32'h13e00001;
      53179: inst = 32'hfe0d96a;
      53180: inst = 32'h5be00000;
      53181: inst = 32'h8c50000;
      53182: inst = 32'h24612800;
      53183: inst = 32'h10a0ffff;
      53184: inst = 32'hca0ffed;
      53185: inst = 32'h24822800;
      53186: inst = 32'h10a00000;
      53187: inst = 32'hca00004;
      53188: inst = 32'h38632800;
      53189: inst = 32'h38842800;
      53190: inst = 32'h10a00000;
      53191: inst = 32'hca0cfcb;
      53192: inst = 32'h13e00001;
      53193: inst = 32'hfe0d96a;
      53194: inst = 32'h5be00000;
      53195: inst = 32'h8c50000;
      53196: inst = 32'h24612800;
      53197: inst = 32'h10a0ffff;
      53198: inst = 32'hca0ffed;
      53199: inst = 32'h24822800;
      53200: inst = 32'h10a00000;
      53201: inst = 32'hca00004;
      53202: inst = 32'h38632800;
      53203: inst = 32'h38842800;
      53204: inst = 32'h10a00000;
      53205: inst = 32'hca0cfd9;
      53206: inst = 32'h13e00001;
      53207: inst = 32'hfe0d96a;
      53208: inst = 32'h5be00000;
      53209: inst = 32'h8c50000;
      53210: inst = 32'h24612800;
      53211: inst = 32'h10a0ffff;
      53212: inst = 32'hca0ffed;
      53213: inst = 32'h24822800;
      53214: inst = 32'h10a00000;
      53215: inst = 32'hca00004;
      53216: inst = 32'h38632800;
      53217: inst = 32'h38842800;
      53218: inst = 32'h10a00000;
      53219: inst = 32'hca0cfe7;
      53220: inst = 32'h13e00001;
      53221: inst = 32'hfe0d96a;
      53222: inst = 32'h5be00000;
      53223: inst = 32'h8c50000;
      53224: inst = 32'h24612800;
      53225: inst = 32'h10a0ffff;
      53226: inst = 32'hca0ffed;
      53227: inst = 32'h24822800;
      53228: inst = 32'h10a00000;
      53229: inst = 32'hca00004;
      53230: inst = 32'h38632800;
      53231: inst = 32'h38842800;
      53232: inst = 32'h10a00000;
      53233: inst = 32'hca0cff5;
      53234: inst = 32'h13e00001;
      53235: inst = 32'hfe0d96a;
      53236: inst = 32'h5be00000;
      53237: inst = 32'h8c50000;
      53238: inst = 32'h24612800;
      53239: inst = 32'h10a0ffff;
      53240: inst = 32'hca0ffed;
      53241: inst = 32'h24822800;
      53242: inst = 32'h10a00000;
      53243: inst = 32'hca00004;
      53244: inst = 32'h38632800;
      53245: inst = 32'h38842800;
      53246: inst = 32'h10a00000;
      53247: inst = 32'hca0d003;
      53248: inst = 32'h13e00001;
      53249: inst = 32'hfe0d96a;
      53250: inst = 32'h5be00000;
      53251: inst = 32'h8c50000;
      53252: inst = 32'h24612800;
      53253: inst = 32'h10a0ffff;
      53254: inst = 32'hca0ffed;
      53255: inst = 32'h24822800;
      53256: inst = 32'h10a00000;
      53257: inst = 32'hca00004;
      53258: inst = 32'h38632800;
      53259: inst = 32'h38842800;
      53260: inst = 32'h10a00000;
      53261: inst = 32'hca0d011;
      53262: inst = 32'h13e00001;
      53263: inst = 32'hfe0d96a;
      53264: inst = 32'h5be00000;
      53265: inst = 32'h8c50000;
      53266: inst = 32'h24612800;
      53267: inst = 32'h10a0ffff;
      53268: inst = 32'hca0ffed;
      53269: inst = 32'h24822800;
      53270: inst = 32'h10a00000;
      53271: inst = 32'hca00004;
      53272: inst = 32'h38632800;
      53273: inst = 32'h38842800;
      53274: inst = 32'h10a00000;
      53275: inst = 32'hca0d01f;
      53276: inst = 32'h13e00001;
      53277: inst = 32'hfe0d96a;
      53278: inst = 32'h5be00000;
      53279: inst = 32'h8c50000;
      53280: inst = 32'h24612800;
      53281: inst = 32'h10a0ffff;
      53282: inst = 32'hca0ffed;
      53283: inst = 32'h24822800;
      53284: inst = 32'h10a00000;
      53285: inst = 32'hca00004;
      53286: inst = 32'h38632800;
      53287: inst = 32'h38842800;
      53288: inst = 32'h10a00000;
      53289: inst = 32'hca0d02d;
      53290: inst = 32'h13e00001;
      53291: inst = 32'hfe0d96a;
      53292: inst = 32'h5be00000;
      53293: inst = 32'h8c50000;
      53294: inst = 32'h24612800;
      53295: inst = 32'h10a0ffff;
      53296: inst = 32'hca0ffed;
      53297: inst = 32'h24822800;
      53298: inst = 32'h10a00000;
      53299: inst = 32'hca00004;
      53300: inst = 32'h38632800;
      53301: inst = 32'h38842800;
      53302: inst = 32'h10a00000;
      53303: inst = 32'hca0d03b;
      53304: inst = 32'h13e00001;
      53305: inst = 32'hfe0d96a;
      53306: inst = 32'h5be00000;
      53307: inst = 32'h8c50000;
      53308: inst = 32'h24612800;
      53309: inst = 32'h10a0ffff;
      53310: inst = 32'hca0ffed;
      53311: inst = 32'h24822800;
      53312: inst = 32'h10a00000;
      53313: inst = 32'hca00004;
      53314: inst = 32'h38632800;
      53315: inst = 32'h38842800;
      53316: inst = 32'h10a00000;
      53317: inst = 32'hca0d049;
      53318: inst = 32'h13e00001;
      53319: inst = 32'hfe0d96a;
      53320: inst = 32'h5be00000;
      53321: inst = 32'h8c50000;
      53322: inst = 32'h24612800;
      53323: inst = 32'h10a0ffff;
      53324: inst = 32'hca0ffed;
      53325: inst = 32'h24822800;
      53326: inst = 32'h10a00000;
      53327: inst = 32'hca00004;
      53328: inst = 32'h38632800;
      53329: inst = 32'h38842800;
      53330: inst = 32'h10a00000;
      53331: inst = 32'hca0d057;
      53332: inst = 32'h13e00001;
      53333: inst = 32'hfe0d96a;
      53334: inst = 32'h5be00000;
      53335: inst = 32'h8c50000;
      53336: inst = 32'h24612800;
      53337: inst = 32'h10a0ffff;
      53338: inst = 32'hca0ffed;
      53339: inst = 32'h24822800;
      53340: inst = 32'h10a00000;
      53341: inst = 32'hca00004;
      53342: inst = 32'h38632800;
      53343: inst = 32'h38842800;
      53344: inst = 32'h10a00000;
      53345: inst = 32'hca0d065;
      53346: inst = 32'h13e00001;
      53347: inst = 32'hfe0d96a;
      53348: inst = 32'h5be00000;
      53349: inst = 32'h8c50000;
      53350: inst = 32'h24612800;
      53351: inst = 32'h10a0ffff;
      53352: inst = 32'hca0ffed;
      53353: inst = 32'h24822800;
      53354: inst = 32'h10a00000;
      53355: inst = 32'hca00004;
      53356: inst = 32'h38632800;
      53357: inst = 32'h38842800;
      53358: inst = 32'h10a00000;
      53359: inst = 32'hca0d073;
      53360: inst = 32'h13e00001;
      53361: inst = 32'hfe0d96a;
      53362: inst = 32'h5be00000;
      53363: inst = 32'h8c50000;
      53364: inst = 32'h24612800;
      53365: inst = 32'h10a0ffff;
      53366: inst = 32'hca0ffed;
      53367: inst = 32'h24822800;
      53368: inst = 32'h10a00000;
      53369: inst = 32'hca00004;
      53370: inst = 32'h38632800;
      53371: inst = 32'h38842800;
      53372: inst = 32'h10a00000;
      53373: inst = 32'hca0d081;
      53374: inst = 32'h13e00001;
      53375: inst = 32'hfe0d96a;
      53376: inst = 32'h5be00000;
      53377: inst = 32'h8c50000;
      53378: inst = 32'h24612800;
      53379: inst = 32'h10a0ffff;
      53380: inst = 32'hca0ffed;
      53381: inst = 32'h24822800;
      53382: inst = 32'h10a00000;
      53383: inst = 32'hca00004;
      53384: inst = 32'h38632800;
      53385: inst = 32'h38842800;
      53386: inst = 32'h10a00000;
      53387: inst = 32'hca0d08f;
      53388: inst = 32'h13e00001;
      53389: inst = 32'hfe0d96a;
      53390: inst = 32'h5be00000;
      53391: inst = 32'h8c50000;
      53392: inst = 32'h24612800;
      53393: inst = 32'h10a0ffff;
      53394: inst = 32'hca0ffed;
      53395: inst = 32'h24822800;
      53396: inst = 32'h10a00000;
      53397: inst = 32'hca00004;
      53398: inst = 32'h38632800;
      53399: inst = 32'h38842800;
      53400: inst = 32'h10a00000;
      53401: inst = 32'hca0d09d;
      53402: inst = 32'h13e00001;
      53403: inst = 32'hfe0d96a;
      53404: inst = 32'h5be00000;
      53405: inst = 32'h8c50000;
      53406: inst = 32'h24612800;
      53407: inst = 32'h10a0ffff;
      53408: inst = 32'hca0ffed;
      53409: inst = 32'h24822800;
      53410: inst = 32'h10a00000;
      53411: inst = 32'hca00004;
      53412: inst = 32'h38632800;
      53413: inst = 32'h38842800;
      53414: inst = 32'h10a00000;
      53415: inst = 32'hca0d0ab;
      53416: inst = 32'h13e00001;
      53417: inst = 32'hfe0d96a;
      53418: inst = 32'h5be00000;
      53419: inst = 32'h8c50000;
      53420: inst = 32'h24612800;
      53421: inst = 32'h10a0ffff;
      53422: inst = 32'hca0ffed;
      53423: inst = 32'h24822800;
      53424: inst = 32'h10a00000;
      53425: inst = 32'hca00004;
      53426: inst = 32'h38632800;
      53427: inst = 32'h38842800;
      53428: inst = 32'h10a00000;
      53429: inst = 32'hca0d0b9;
      53430: inst = 32'h13e00001;
      53431: inst = 32'hfe0d96a;
      53432: inst = 32'h5be00000;
      53433: inst = 32'h8c50000;
      53434: inst = 32'h24612800;
      53435: inst = 32'h10a0ffff;
      53436: inst = 32'hca0ffed;
      53437: inst = 32'h24822800;
      53438: inst = 32'h10a00000;
      53439: inst = 32'hca00004;
      53440: inst = 32'h38632800;
      53441: inst = 32'h38842800;
      53442: inst = 32'h10a00000;
      53443: inst = 32'hca0d0c7;
      53444: inst = 32'h13e00001;
      53445: inst = 32'hfe0d96a;
      53446: inst = 32'h5be00000;
      53447: inst = 32'h8c50000;
      53448: inst = 32'h24612800;
      53449: inst = 32'h10a0ffff;
      53450: inst = 32'hca0ffed;
      53451: inst = 32'h24822800;
      53452: inst = 32'h10a00000;
      53453: inst = 32'hca00004;
      53454: inst = 32'h38632800;
      53455: inst = 32'h38842800;
      53456: inst = 32'h10a00000;
      53457: inst = 32'hca0d0d5;
      53458: inst = 32'h13e00001;
      53459: inst = 32'hfe0d96a;
      53460: inst = 32'h5be00000;
      53461: inst = 32'h8c50000;
      53462: inst = 32'h24612800;
      53463: inst = 32'h10a0ffff;
      53464: inst = 32'hca0ffed;
      53465: inst = 32'h24822800;
      53466: inst = 32'h10a00000;
      53467: inst = 32'hca00004;
      53468: inst = 32'h38632800;
      53469: inst = 32'h38842800;
      53470: inst = 32'h10a00000;
      53471: inst = 32'hca0d0e3;
      53472: inst = 32'h13e00001;
      53473: inst = 32'hfe0d96a;
      53474: inst = 32'h5be00000;
      53475: inst = 32'h8c50000;
      53476: inst = 32'h24612800;
      53477: inst = 32'h10a0ffff;
      53478: inst = 32'hca0ffed;
      53479: inst = 32'h24822800;
      53480: inst = 32'h10a00000;
      53481: inst = 32'hca00004;
      53482: inst = 32'h38632800;
      53483: inst = 32'h38842800;
      53484: inst = 32'h10a00000;
      53485: inst = 32'hca0d0f1;
      53486: inst = 32'h13e00001;
      53487: inst = 32'hfe0d96a;
      53488: inst = 32'h5be00000;
      53489: inst = 32'h8c50000;
      53490: inst = 32'h24612800;
      53491: inst = 32'h10a0ffff;
      53492: inst = 32'hca0ffed;
      53493: inst = 32'h24822800;
      53494: inst = 32'h10a00000;
      53495: inst = 32'hca00004;
      53496: inst = 32'h38632800;
      53497: inst = 32'h38842800;
      53498: inst = 32'h10a00000;
      53499: inst = 32'hca0d0ff;
      53500: inst = 32'h13e00001;
      53501: inst = 32'hfe0d96a;
      53502: inst = 32'h5be00000;
      53503: inst = 32'h8c50000;
      53504: inst = 32'h24612800;
      53505: inst = 32'h10a0ffff;
      53506: inst = 32'hca0ffed;
      53507: inst = 32'h24822800;
      53508: inst = 32'h10a00000;
      53509: inst = 32'hca00004;
      53510: inst = 32'h38632800;
      53511: inst = 32'h38842800;
      53512: inst = 32'h10a00000;
      53513: inst = 32'hca0d10d;
      53514: inst = 32'h13e00001;
      53515: inst = 32'hfe0d96a;
      53516: inst = 32'h5be00000;
      53517: inst = 32'h8c50000;
      53518: inst = 32'h24612800;
      53519: inst = 32'h10a0ffff;
      53520: inst = 32'hca0ffed;
      53521: inst = 32'h24822800;
      53522: inst = 32'h10a00000;
      53523: inst = 32'hca00004;
      53524: inst = 32'h38632800;
      53525: inst = 32'h38842800;
      53526: inst = 32'h10a00000;
      53527: inst = 32'hca0d11b;
      53528: inst = 32'h13e00001;
      53529: inst = 32'hfe0d96a;
      53530: inst = 32'h5be00000;
      53531: inst = 32'h8c50000;
      53532: inst = 32'h24612800;
      53533: inst = 32'h10a0ffff;
      53534: inst = 32'hca0ffed;
      53535: inst = 32'h24822800;
      53536: inst = 32'h10a00000;
      53537: inst = 32'hca00004;
      53538: inst = 32'h38632800;
      53539: inst = 32'h38842800;
      53540: inst = 32'h10a00000;
      53541: inst = 32'hca0d129;
      53542: inst = 32'h13e00001;
      53543: inst = 32'hfe0d96a;
      53544: inst = 32'h5be00000;
      53545: inst = 32'h8c50000;
      53546: inst = 32'h24612800;
      53547: inst = 32'h10a0ffff;
      53548: inst = 32'hca0ffed;
      53549: inst = 32'h24822800;
      53550: inst = 32'h10a00000;
      53551: inst = 32'hca00004;
      53552: inst = 32'h38632800;
      53553: inst = 32'h38842800;
      53554: inst = 32'h10a00000;
      53555: inst = 32'hca0d137;
      53556: inst = 32'h13e00001;
      53557: inst = 32'hfe0d96a;
      53558: inst = 32'h5be00000;
      53559: inst = 32'h8c50000;
      53560: inst = 32'h24612800;
      53561: inst = 32'h10a0ffff;
      53562: inst = 32'hca0ffed;
      53563: inst = 32'h24822800;
      53564: inst = 32'h10a00000;
      53565: inst = 32'hca00004;
      53566: inst = 32'h38632800;
      53567: inst = 32'h38842800;
      53568: inst = 32'h10a00000;
      53569: inst = 32'hca0d145;
      53570: inst = 32'h13e00001;
      53571: inst = 32'hfe0d96a;
      53572: inst = 32'h5be00000;
      53573: inst = 32'h8c50000;
      53574: inst = 32'h24612800;
      53575: inst = 32'h10a0ffff;
      53576: inst = 32'hca0ffed;
      53577: inst = 32'h24822800;
      53578: inst = 32'h10a00000;
      53579: inst = 32'hca00004;
      53580: inst = 32'h38632800;
      53581: inst = 32'h38842800;
      53582: inst = 32'h10a00000;
      53583: inst = 32'hca0d153;
      53584: inst = 32'h13e00001;
      53585: inst = 32'hfe0d96a;
      53586: inst = 32'h5be00000;
      53587: inst = 32'h8c50000;
      53588: inst = 32'h24612800;
      53589: inst = 32'h10a0ffff;
      53590: inst = 32'hca0ffed;
      53591: inst = 32'h24822800;
      53592: inst = 32'h10a00000;
      53593: inst = 32'hca00004;
      53594: inst = 32'h38632800;
      53595: inst = 32'h38842800;
      53596: inst = 32'h10a00000;
      53597: inst = 32'hca0d161;
      53598: inst = 32'h13e00001;
      53599: inst = 32'hfe0d96a;
      53600: inst = 32'h5be00000;
      53601: inst = 32'h8c50000;
      53602: inst = 32'h24612800;
      53603: inst = 32'h10a0ffff;
      53604: inst = 32'hca0ffed;
      53605: inst = 32'h24822800;
      53606: inst = 32'h10a00000;
      53607: inst = 32'hca00004;
      53608: inst = 32'h38632800;
      53609: inst = 32'h38842800;
      53610: inst = 32'h10a00000;
      53611: inst = 32'hca0d16f;
      53612: inst = 32'h13e00001;
      53613: inst = 32'hfe0d96a;
      53614: inst = 32'h5be00000;
      53615: inst = 32'h8c50000;
      53616: inst = 32'h24612800;
      53617: inst = 32'h10a0ffff;
      53618: inst = 32'hca0ffed;
      53619: inst = 32'h24822800;
      53620: inst = 32'h10a00000;
      53621: inst = 32'hca00004;
      53622: inst = 32'h38632800;
      53623: inst = 32'h38842800;
      53624: inst = 32'h10a00000;
      53625: inst = 32'hca0d17d;
      53626: inst = 32'h13e00001;
      53627: inst = 32'hfe0d96a;
      53628: inst = 32'h5be00000;
      53629: inst = 32'h8c50000;
      53630: inst = 32'h24612800;
      53631: inst = 32'h10a0ffff;
      53632: inst = 32'hca0ffed;
      53633: inst = 32'h24822800;
      53634: inst = 32'h10a00000;
      53635: inst = 32'hca00004;
      53636: inst = 32'h38632800;
      53637: inst = 32'h38842800;
      53638: inst = 32'h10a00000;
      53639: inst = 32'hca0d18b;
      53640: inst = 32'h13e00001;
      53641: inst = 32'hfe0d96a;
      53642: inst = 32'h5be00000;
      53643: inst = 32'h8c50000;
      53644: inst = 32'h24612800;
      53645: inst = 32'h10a0ffff;
      53646: inst = 32'hca0ffed;
      53647: inst = 32'h24822800;
      53648: inst = 32'h10a00000;
      53649: inst = 32'hca00004;
      53650: inst = 32'h38632800;
      53651: inst = 32'h38842800;
      53652: inst = 32'h10a00000;
      53653: inst = 32'hca0d199;
      53654: inst = 32'h13e00001;
      53655: inst = 32'hfe0d96a;
      53656: inst = 32'h5be00000;
      53657: inst = 32'h8c50000;
      53658: inst = 32'h24612800;
      53659: inst = 32'h10a0ffff;
      53660: inst = 32'hca0ffed;
      53661: inst = 32'h24822800;
      53662: inst = 32'h10a00000;
      53663: inst = 32'hca00004;
      53664: inst = 32'h38632800;
      53665: inst = 32'h38842800;
      53666: inst = 32'h10a00000;
      53667: inst = 32'hca0d1a7;
      53668: inst = 32'h13e00001;
      53669: inst = 32'hfe0d96a;
      53670: inst = 32'h5be00000;
      53671: inst = 32'h8c50000;
      53672: inst = 32'h24612800;
      53673: inst = 32'h10a0ffff;
      53674: inst = 32'hca0ffed;
      53675: inst = 32'h24822800;
      53676: inst = 32'h10a00000;
      53677: inst = 32'hca00004;
      53678: inst = 32'h38632800;
      53679: inst = 32'h38842800;
      53680: inst = 32'h10a00000;
      53681: inst = 32'hca0d1b5;
      53682: inst = 32'h13e00001;
      53683: inst = 32'hfe0d96a;
      53684: inst = 32'h5be00000;
      53685: inst = 32'h8c50000;
      53686: inst = 32'h24612800;
      53687: inst = 32'h10a0ffff;
      53688: inst = 32'hca0ffed;
      53689: inst = 32'h24822800;
      53690: inst = 32'h10a00000;
      53691: inst = 32'hca00004;
      53692: inst = 32'h38632800;
      53693: inst = 32'h38842800;
      53694: inst = 32'h10a00000;
      53695: inst = 32'hca0d1c3;
      53696: inst = 32'h13e00001;
      53697: inst = 32'hfe0d96a;
      53698: inst = 32'h5be00000;
      53699: inst = 32'h8c50000;
      53700: inst = 32'h24612800;
      53701: inst = 32'h10a0ffff;
      53702: inst = 32'hca0ffed;
      53703: inst = 32'h24822800;
      53704: inst = 32'h10a00000;
      53705: inst = 32'hca00004;
      53706: inst = 32'h38632800;
      53707: inst = 32'h38842800;
      53708: inst = 32'h10a00000;
      53709: inst = 32'hca0d1d1;
      53710: inst = 32'h13e00001;
      53711: inst = 32'hfe0d96a;
      53712: inst = 32'h5be00000;
      53713: inst = 32'h8c50000;
      53714: inst = 32'h24612800;
      53715: inst = 32'h10a0ffff;
      53716: inst = 32'hca0ffed;
      53717: inst = 32'h24822800;
      53718: inst = 32'h10a00000;
      53719: inst = 32'hca00004;
      53720: inst = 32'h38632800;
      53721: inst = 32'h38842800;
      53722: inst = 32'h10a00000;
      53723: inst = 32'hca0d1df;
      53724: inst = 32'h13e00001;
      53725: inst = 32'hfe0d96a;
      53726: inst = 32'h5be00000;
      53727: inst = 32'h8c50000;
      53728: inst = 32'h24612800;
      53729: inst = 32'h10a0ffff;
      53730: inst = 32'hca0ffed;
      53731: inst = 32'h24822800;
      53732: inst = 32'h10a00000;
      53733: inst = 32'hca00004;
      53734: inst = 32'h38632800;
      53735: inst = 32'h38842800;
      53736: inst = 32'h10a00000;
      53737: inst = 32'hca0d1ed;
      53738: inst = 32'h13e00001;
      53739: inst = 32'hfe0d96a;
      53740: inst = 32'h5be00000;
      53741: inst = 32'h8c50000;
      53742: inst = 32'h24612800;
      53743: inst = 32'h10a0ffff;
      53744: inst = 32'hca0ffed;
      53745: inst = 32'h24822800;
      53746: inst = 32'h10a00000;
      53747: inst = 32'hca00004;
      53748: inst = 32'h38632800;
      53749: inst = 32'h38842800;
      53750: inst = 32'h10a00000;
      53751: inst = 32'hca0d1fb;
      53752: inst = 32'h13e00001;
      53753: inst = 32'hfe0d96a;
      53754: inst = 32'h5be00000;
      53755: inst = 32'h8c50000;
      53756: inst = 32'h24612800;
      53757: inst = 32'h10a0ffff;
      53758: inst = 32'hca0ffed;
      53759: inst = 32'h24822800;
      53760: inst = 32'h10a00000;
      53761: inst = 32'hca00004;
      53762: inst = 32'h38632800;
      53763: inst = 32'h38842800;
      53764: inst = 32'h10a00000;
      53765: inst = 32'hca0d209;
      53766: inst = 32'h13e00001;
      53767: inst = 32'hfe0d96a;
      53768: inst = 32'h5be00000;
      53769: inst = 32'h8c50000;
      53770: inst = 32'h24612800;
      53771: inst = 32'h10a0ffff;
      53772: inst = 32'hca0ffed;
      53773: inst = 32'h24822800;
      53774: inst = 32'h10a00000;
      53775: inst = 32'hca00004;
      53776: inst = 32'h38632800;
      53777: inst = 32'h38842800;
      53778: inst = 32'h10a00000;
      53779: inst = 32'hca0d217;
      53780: inst = 32'h13e00001;
      53781: inst = 32'hfe0d96a;
      53782: inst = 32'h5be00000;
      53783: inst = 32'h8c50000;
      53784: inst = 32'h24612800;
      53785: inst = 32'h10a0ffff;
      53786: inst = 32'hca0ffed;
      53787: inst = 32'h24822800;
      53788: inst = 32'h10a00000;
      53789: inst = 32'hca00004;
      53790: inst = 32'h38632800;
      53791: inst = 32'h38842800;
      53792: inst = 32'h10a00000;
      53793: inst = 32'hca0d225;
      53794: inst = 32'h13e00001;
      53795: inst = 32'hfe0d96a;
      53796: inst = 32'h5be00000;
      53797: inst = 32'h8c50000;
      53798: inst = 32'h24612800;
      53799: inst = 32'h10a0ffff;
      53800: inst = 32'hca0ffed;
      53801: inst = 32'h24822800;
      53802: inst = 32'h10a00000;
      53803: inst = 32'hca00004;
      53804: inst = 32'h38632800;
      53805: inst = 32'h38842800;
      53806: inst = 32'h10a00000;
      53807: inst = 32'hca0d233;
      53808: inst = 32'h13e00001;
      53809: inst = 32'hfe0d96a;
      53810: inst = 32'h5be00000;
      53811: inst = 32'h8c50000;
      53812: inst = 32'h24612800;
      53813: inst = 32'h10a0ffff;
      53814: inst = 32'hca0ffed;
      53815: inst = 32'h24822800;
      53816: inst = 32'h10a00000;
      53817: inst = 32'hca00004;
      53818: inst = 32'h38632800;
      53819: inst = 32'h38842800;
      53820: inst = 32'h10a00000;
      53821: inst = 32'hca0d241;
      53822: inst = 32'h13e00001;
      53823: inst = 32'hfe0d96a;
      53824: inst = 32'h5be00000;
      53825: inst = 32'h8c50000;
      53826: inst = 32'h24612800;
      53827: inst = 32'h10a0ffff;
      53828: inst = 32'hca0ffed;
      53829: inst = 32'h24822800;
      53830: inst = 32'h10a00000;
      53831: inst = 32'hca00004;
      53832: inst = 32'h38632800;
      53833: inst = 32'h38842800;
      53834: inst = 32'h10a00000;
      53835: inst = 32'hca0d24f;
      53836: inst = 32'h13e00001;
      53837: inst = 32'hfe0d96a;
      53838: inst = 32'h5be00000;
      53839: inst = 32'h8c50000;
      53840: inst = 32'h24612800;
      53841: inst = 32'h10a0ffff;
      53842: inst = 32'hca0ffed;
      53843: inst = 32'h24822800;
      53844: inst = 32'h10a00000;
      53845: inst = 32'hca00004;
      53846: inst = 32'h38632800;
      53847: inst = 32'h38842800;
      53848: inst = 32'h10a00000;
      53849: inst = 32'hca0d25d;
      53850: inst = 32'h13e00001;
      53851: inst = 32'hfe0d96a;
      53852: inst = 32'h5be00000;
      53853: inst = 32'h8c50000;
      53854: inst = 32'h24612800;
      53855: inst = 32'h10a0ffff;
      53856: inst = 32'hca0ffed;
      53857: inst = 32'h24822800;
      53858: inst = 32'h10a00000;
      53859: inst = 32'hca00004;
      53860: inst = 32'h38632800;
      53861: inst = 32'h38842800;
      53862: inst = 32'h10a00000;
      53863: inst = 32'hca0d26b;
      53864: inst = 32'h13e00001;
      53865: inst = 32'hfe0d96a;
      53866: inst = 32'h5be00000;
      53867: inst = 32'h8c50000;
      53868: inst = 32'h24612800;
      53869: inst = 32'h10a0ffff;
      53870: inst = 32'hca0ffed;
      53871: inst = 32'h24822800;
      53872: inst = 32'h10a00000;
      53873: inst = 32'hca00004;
      53874: inst = 32'h38632800;
      53875: inst = 32'h38842800;
      53876: inst = 32'h10a00000;
      53877: inst = 32'hca0d279;
      53878: inst = 32'h13e00001;
      53879: inst = 32'hfe0d96a;
      53880: inst = 32'h5be00000;
      53881: inst = 32'h8c50000;
      53882: inst = 32'h24612800;
      53883: inst = 32'h10a0ffff;
      53884: inst = 32'hca0ffed;
      53885: inst = 32'h24822800;
      53886: inst = 32'h10a00000;
      53887: inst = 32'hca00004;
      53888: inst = 32'h38632800;
      53889: inst = 32'h38842800;
      53890: inst = 32'h10a00000;
      53891: inst = 32'hca0d287;
      53892: inst = 32'h13e00001;
      53893: inst = 32'hfe0d96a;
      53894: inst = 32'h5be00000;
      53895: inst = 32'h8c50000;
      53896: inst = 32'h24612800;
      53897: inst = 32'h10a0ffff;
      53898: inst = 32'hca0ffed;
      53899: inst = 32'h24822800;
      53900: inst = 32'h10a00000;
      53901: inst = 32'hca00004;
      53902: inst = 32'h38632800;
      53903: inst = 32'h38842800;
      53904: inst = 32'h10a00000;
      53905: inst = 32'hca0d295;
      53906: inst = 32'h13e00001;
      53907: inst = 32'hfe0d96a;
      53908: inst = 32'h5be00000;
      53909: inst = 32'h8c50000;
      53910: inst = 32'h24612800;
      53911: inst = 32'h10a0ffff;
      53912: inst = 32'hca0ffed;
      53913: inst = 32'h24822800;
      53914: inst = 32'h10a00000;
      53915: inst = 32'hca00004;
      53916: inst = 32'h38632800;
      53917: inst = 32'h38842800;
      53918: inst = 32'h10a00000;
      53919: inst = 32'hca0d2a3;
      53920: inst = 32'h13e00001;
      53921: inst = 32'hfe0d96a;
      53922: inst = 32'h5be00000;
      53923: inst = 32'h8c50000;
      53924: inst = 32'h24612800;
      53925: inst = 32'h10a0ffff;
      53926: inst = 32'hca0ffed;
      53927: inst = 32'h24822800;
      53928: inst = 32'h10a00000;
      53929: inst = 32'hca00004;
      53930: inst = 32'h38632800;
      53931: inst = 32'h38842800;
      53932: inst = 32'h10a00000;
      53933: inst = 32'hca0d2b1;
      53934: inst = 32'h13e00001;
      53935: inst = 32'hfe0d96a;
      53936: inst = 32'h5be00000;
      53937: inst = 32'h8c50000;
      53938: inst = 32'h24612800;
      53939: inst = 32'h10a0ffff;
      53940: inst = 32'hca0ffed;
      53941: inst = 32'h24822800;
      53942: inst = 32'h10a00000;
      53943: inst = 32'hca00004;
      53944: inst = 32'h38632800;
      53945: inst = 32'h38842800;
      53946: inst = 32'h10a00000;
      53947: inst = 32'hca0d2bf;
      53948: inst = 32'h13e00001;
      53949: inst = 32'hfe0d96a;
      53950: inst = 32'h5be00000;
      53951: inst = 32'h8c50000;
      53952: inst = 32'h24612800;
      53953: inst = 32'h10a0ffff;
      53954: inst = 32'hca0ffed;
      53955: inst = 32'h24822800;
      53956: inst = 32'h10a00000;
      53957: inst = 32'hca00004;
      53958: inst = 32'h38632800;
      53959: inst = 32'h38842800;
      53960: inst = 32'h10a00000;
      53961: inst = 32'hca0d2cd;
      53962: inst = 32'h13e00001;
      53963: inst = 32'hfe0d96a;
      53964: inst = 32'h5be00000;
      53965: inst = 32'h8c50000;
      53966: inst = 32'h24612800;
      53967: inst = 32'h10a0ffff;
      53968: inst = 32'hca0ffed;
      53969: inst = 32'h24822800;
      53970: inst = 32'h10a00000;
      53971: inst = 32'hca00004;
      53972: inst = 32'h38632800;
      53973: inst = 32'h38842800;
      53974: inst = 32'h10a00000;
      53975: inst = 32'hca0d2db;
      53976: inst = 32'h13e00001;
      53977: inst = 32'hfe0d96a;
      53978: inst = 32'h5be00000;
      53979: inst = 32'h8c50000;
      53980: inst = 32'h24612800;
      53981: inst = 32'h10a0ffff;
      53982: inst = 32'hca0ffed;
      53983: inst = 32'h24822800;
      53984: inst = 32'h10a00000;
      53985: inst = 32'hca00004;
      53986: inst = 32'h38632800;
      53987: inst = 32'h38842800;
      53988: inst = 32'h10a00000;
      53989: inst = 32'hca0d2e9;
      53990: inst = 32'h13e00001;
      53991: inst = 32'hfe0d96a;
      53992: inst = 32'h5be00000;
      53993: inst = 32'h8c50000;
      53994: inst = 32'h24612800;
      53995: inst = 32'h10a0ffff;
      53996: inst = 32'hca0ffee;
      53997: inst = 32'h24822800;
      53998: inst = 32'h10a00000;
      53999: inst = 32'hca00004;
      54000: inst = 32'h38632800;
      54001: inst = 32'h38842800;
      54002: inst = 32'h10a00000;
      54003: inst = 32'hca0d2f7;
      54004: inst = 32'h13e00001;
      54005: inst = 32'hfe0d96a;
      54006: inst = 32'h5be00000;
      54007: inst = 32'h8c50000;
      54008: inst = 32'h24612800;
      54009: inst = 32'h10a0ffff;
      54010: inst = 32'hca0ffee;
      54011: inst = 32'h24822800;
      54012: inst = 32'h10a00000;
      54013: inst = 32'hca00004;
      54014: inst = 32'h38632800;
      54015: inst = 32'h38842800;
      54016: inst = 32'h10a00000;
      54017: inst = 32'hca0d305;
      54018: inst = 32'h13e00001;
      54019: inst = 32'hfe0d96a;
      54020: inst = 32'h5be00000;
      54021: inst = 32'h8c50000;
      54022: inst = 32'h24612800;
      54023: inst = 32'h10a0ffff;
      54024: inst = 32'hca0ffee;
      54025: inst = 32'h24822800;
      54026: inst = 32'h10a00000;
      54027: inst = 32'hca00004;
      54028: inst = 32'h38632800;
      54029: inst = 32'h38842800;
      54030: inst = 32'h10a00000;
      54031: inst = 32'hca0d313;
      54032: inst = 32'h13e00001;
      54033: inst = 32'hfe0d96a;
      54034: inst = 32'h5be00000;
      54035: inst = 32'h8c50000;
      54036: inst = 32'h24612800;
      54037: inst = 32'h10a0ffff;
      54038: inst = 32'hca0ffee;
      54039: inst = 32'h24822800;
      54040: inst = 32'h10a00000;
      54041: inst = 32'hca00004;
      54042: inst = 32'h38632800;
      54043: inst = 32'h38842800;
      54044: inst = 32'h10a00000;
      54045: inst = 32'hca0d321;
      54046: inst = 32'h13e00001;
      54047: inst = 32'hfe0d96a;
      54048: inst = 32'h5be00000;
      54049: inst = 32'h8c50000;
      54050: inst = 32'h24612800;
      54051: inst = 32'h10a0ffff;
      54052: inst = 32'hca0ffee;
      54053: inst = 32'h24822800;
      54054: inst = 32'h10a00000;
      54055: inst = 32'hca00004;
      54056: inst = 32'h38632800;
      54057: inst = 32'h38842800;
      54058: inst = 32'h10a00000;
      54059: inst = 32'hca0d32f;
      54060: inst = 32'h13e00001;
      54061: inst = 32'hfe0d96a;
      54062: inst = 32'h5be00000;
      54063: inst = 32'h8c50000;
      54064: inst = 32'h24612800;
      54065: inst = 32'h10a0ffff;
      54066: inst = 32'hca0ffee;
      54067: inst = 32'h24822800;
      54068: inst = 32'h10a00000;
      54069: inst = 32'hca00004;
      54070: inst = 32'h38632800;
      54071: inst = 32'h38842800;
      54072: inst = 32'h10a00000;
      54073: inst = 32'hca0d33d;
      54074: inst = 32'h13e00001;
      54075: inst = 32'hfe0d96a;
      54076: inst = 32'h5be00000;
      54077: inst = 32'h8c50000;
      54078: inst = 32'h24612800;
      54079: inst = 32'h10a0ffff;
      54080: inst = 32'hca0ffee;
      54081: inst = 32'h24822800;
      54082: inst = 32'h10a00000;
      54083: inst = 32'hca00004;
      54084: inst = 32'h38632800;
      54085: inst = 32'h38842800;
      54086: inst = 32'h10a00000;
      54087: inst = 32'hca0d34b;
      54088: inst = 32'h13e00001;
      54089: inst = 32'hfe0d96a;
      54090: inst = 32'h5be00000;
      54091: inst = 32'h8c50000;
      54092: inst = 32'h24612800;
      54093: inst = 32'h10a0ffff;
      54094: inst = 32'hca0ffee;
      54095: inst = 32'h24822800;
      54096: inst = 32'h10a00000;
      54097: inst = 32'hca00004;
      54098: inst = 32'h38632800;
      54099: inst = 32'h38842800;
      54100: inst = 32'h10a00000;
      54101: inst = 32'hca0d359;
      54102: inst = 32'h13e00001;
      54103: inst = 32'hfe0d96a;
      54104: inst = 32'h5be00000;
      54105: inst = 32'h8c50000;
      54106: inst = 32'h24612800;
      54107: inst = 32'h10a0ffff;
      54108: inst = 32'hca0ffee;
      54109: inst = 32'h24822800;
      54110: inst = 32'h10a00000;
      54111: inst = 32'hca00004;
      54112: inst = 32'h38632800;
      54113: inst = 32'h38842800;
      54114: inst = 32'h10a00000;
      54115: inst = 32'hca0d367;
      54116: inst = 32'h13e00001;
      54117: inst = 32'hfe0d96a;
      54118: inst = 32'h5be00000;
      54119: inst = 32'h8c50000;
      54120: inst = 32'h24612800;
      54121: inst = 32'h10a0ffff;
      54122: inst = 32'hca0ffee;
      54123: inst = 32'h24822800;
      54124: inst = 32'h10a00000;
      54125: inst = 32'hca00004;
      54126: inst = 32'h38632800;
      54127: inst = 32'h38842800;
      54128: inst = 32'h10a00000;
      54129: inst = 32'hca0d375;
      54130: inst = 32'h13e00001;
      54131: inst = 32'hfe0d96a;
      54132: inst = 32'h5be00000;
      54133: inst = 32'h8c50000;
      54134: inst = 32'h24612800;
      54135: inst = 32'h10a0ffff;
      54136: inst = 32'hca0ffee;
      54137: inst = 32'h24822800;
      54138: inst = 32'h10a00000;
      54139: inst = 32'hca00004;
      54140: inst = 32'h38632800;
      54141: inst = 32'h38842800;
      54142: inst = 32'h10a00000;
      54143: inst = 32'hca0d383;
      54144: inst = 32'h13e00001;
      54145: inst = 32'hfe0d96a;
      54146: inst = 32'h5be00000;
      54147: inst = 32'h8c50000;
      54148: inst = 32'h24612800;
      54149: inst = 32'h10a0ffff;
      54150: inst = 32'hca0ffee;
      54151: inst = 32'h24822800;
      54152: inst = 32'h10a00000;
      54153: inst = 32'hca00004;
      54154: inst = 32'h38632800;
      54155: inst = 32'h38842800;
      54156: inst = 32'h10a00000;
      54157: inst = 32'hca0d391;
      54158: inst = 32'h13e00001;
      54159: inst = 32'hfe0d96a;
      54160: inst = 32'h5be00000;
      54161: inst = 32'h8c50000;
      54162: inst = 32'h24612800;
      54163: inst = 32'h10a0ffff;
      54164: inst = 32'hca0ffee;
      54165: inst = 32'h24822800;
      54166: inst = 32'h10a00000;
      54167: inst = 32'hca00004;
      54168: inst = 32'h38632800;
      54169: inst = 32'h38842800;
      54170: inst = 32'h10a00000;
      54171: inst = 32'hca0d39f;
      54172: inst = 32'h13e00001;
      54173: inst = 32'hfe0d96a;
      54174: inst = 32'h5be00000;
      54175: inst = 32'h8c50000;
      54176: inst = 32'h24612800;
      54177: inst = 32'h10a0ffff;
      54178: inst = 32'hca0ffee;
      54179: inst = 32'h24822800;
      54180: inst = 32'h10a00000;
      54181: inst = 32'hca00004;
      54182: inst = 32'h38632800;
      54183: inst = 32'h38842800;
      54184: inst = 32'h10a00000;
      54185: inst = 32'hca0d3ad;
      54186: inst = 32'h13e00001;
      54187: inst = 32'hfe0d96a;
      54188: inst = 32'h5be00000;
      54189: inst = 32'h8c50000;
      54190: inst = 32'h24612800;
      54191: inst = 32'h10a0ffff;
      54192: inst = 32'hca0ffee;
      54193: inst = 32'h24822800;
      54194: inst = 32'h10a00000;
      54195: inst = 32'hca00004;
      54196: inst = 32'h38632800;
      54197: inst = 32'h38842800;
      54198: inst = 32'h10a00000;
      54199: inst = 32'hca0d3bb;
      54200: inst = 32'h13e00001;
      54201: inst = 32'hfe0d96a;
      54202: inst = 32'h5be00000;
      54203: inst = 32'h8c50000;
      54204: inst = 32'h24612800;
      54205: inst = 32'h10a0ffff;
      54206: inst = 32'hca0ffee;
      54207: inst = 32'h24822800;
      54208: inst = 32'h10a00000;
      54209: inst = 32'hca00004;
      54210: inst = 32'h38632800;
      54211: inst = 32'h38842800;
      54212: inst = 32'h10a00000;
      54213: inst = 32'hca0d3c9;
      54214: inst = 32'h13e00001;
      54215: inst = 32'hfe0d96a;
      54216: inst = 32'h5be00000;
      54217: inst = 32'h8c50000;
      54218: inst = 32'h24612800;
      54219: inst = 32'h10a0ffff;
      54220: inst = 32'hca0ffee;
      54221: inst = 32'h24822800;
      54222: inst = 32'h10a00000;
      54223: inst = 32'hca00004;
      54224: inst = 32'h38632800;
      54225: inst = 32'h38842800;
      54226: inst = 32'h10a00000;
      54227: inst = 32'hca0d3d7;
      54228: inst = 32'h13e00001;
      54229: inst = 32'hfe0d96a;
      54230: inst = 32'h5be00000;
      54231: inst = 32'h8c50000;
      54232: inst = 32'h24612800;
      54233: inst = 32'h10a0ffff;
      54234: inst = 32'hca0ffee;
      54235: inst = 32'h24822800;
      54236: inst = 32'h10a00000;
      54237: inst = 32'hca00004;
      54238: inst = 32'h38632800;
      54239: inst = 32'h38842800;
      54240: inst = 32'h10a00000;
      54241: inst = 32'hca0d3e5;
      54242: inst = 32'h13e00001;
      54243: inst = 32'hfe0d96a;
      54244: inst = 32'h5be00000;
      54245: inst = 32'h8c50000;
      54246: inst = 32'h24612800;
      54247: inst = 32'h10a0ffff;
      54248: inst = 32'hca0ffee;
      54249: inst = 32'h24822800;
      54250: inst = 32'h10a00000;
      54251: inst = 32'hca00004;
      54252: inst = 32'h38632800;
      54253: inst = 32'h38842800;
      54254: inst = 32'h10a00000;
      54255: inst = 32'hca0d3f3;
      54256: inst = 32'h13e00001;
      54257: inst = 32'hfe0d96a;
      54258: inst = 32'h5be00000;
      54259: inst = 32'h8c50000;
      54260: inst = 32'h24612800;
      54261: inst = 32'h10a0ffff;
      54262: inst = 32'hca0ffee;
      54263: inst = 32'h24822800;
      54264: inst = 32'h10a00000;
      54265: inst = 32'hca00004;
      54266: inst = 32'h38632800;
      54267: inst = 32'h38842800;
      54268: inst = 32'h10a00000;
      54269: inst = 32'hca0d401;
      54270: inst = 32'h13e00001;
      54271: inst = 32'hfe0d96a;
      54272: inst = 32'h5be00000;
      54273: inst = 32'h8c50000;
      54274: inst = 32'h24612800;
      54275: inst = 32'h10a0ffff;
      54276: inst = 32'hca0ffee;
      54277: inst = 32'h24822800;
      54278: inst = 32'h10a00000;
      54279: inst = 32'hca00004;
      54280: inst = 32'h38632800;
      54281: inst = 32'h38842800;
      54282: inst = 32'h10a00000;
      54283: inst = 32'hca0d40f;
      54284: inst = 32'h13e00001;
      54285: inst = 32'hfe0d96a;
      54286: inst = 32'h5be00000;
      54287: inst = 32'h8c50000;
      54288: inst = 32'h24612800;
      54289: inst = 32'h10a0ffff;
      54290: inst = 32'hca0ffee;
      54291: inst = 32'h24822800;
      54292: inst = 32'h10a00000;
      54293: inst = 32'hca00004;
      54294: inst = 32'h38632800;
      54295: inst = 32'h38842800;
      54296: inst = 32'h10a00000;
      54297: inst = 32'hca0d41d;
      54298: inst = 32'h13e00001;
      54299: inst = 32'hfe0d96a;
      54300: inst = 32'h5be00000;
      54301: inst = 32'h8c50000;
      54302: inst = 32'h24612800;
      54303: inst = 32'h10a0ffff;
      54304: inst = 32'hca0ffee;
      54305: inst = 32'h24822800;
      54306: inst = 32'h10a00000;
      54307: inst = 32'hca00004;
      54308: inst = 32'h38632800;
      54309: inst = 32'h38842800;
      54310: inst = 32'h10a00000;
      54311: inst = 32'hca0d42b;
      54312: inst = 32'h13e00001;
      54313: inst = 32'hfe0d96a;
      54314: inst = 32'h5be00000;
      54315: inst = 32'h8c50000;
      54316: inst = 32'h24612800;
      54317: inst = 32'h10a0ffff;
      54318: inst = 32'hca0ffee;
      54319: inst = 32'h24822800;
      54320: inst = 32'h10a00000;
      54321: inst = 32'hca00004;
      54322: inst = 32'h38632800;
      54323: inst = 32'h38842800;
      54324: inst = 32'h10a00000;
      54325: inst = 32'hca0d439;
      54326: inst = 32'h13e00001;
      54327: inst = 32'hfe0d96a;
      54328: inst = 32'h5be00000;
      54329: inst = 32'h8c50000;
      54330: inst = 32'h24612800;
      54331: inst = 32'h10a0ffff;
      54332: inst = 32'hca0ffee;
      54333: inst = 32'h24822800;
      54334: inst = 32'h10a00000;
      54335: inst = 32'hca00004;
      54336: inst = 32'h38632800;
      54337: inst = 32'h38842800;
      54338: inst = 32'h10a00000;
      54339: inst = 32'hca0d447;
      54340: inst = 32'h13e00001;
      54341: inst = 32'hfe0d96a;
      54342: inst = 32'h5be00000;
      54343: inst = 32'h8c50000;
      54344: inst = 32'h24612800;
      54345: inst = 32'h10a0ffff;
      54346: inst = 32'hca0ffee;
      54347: inst = 32'h24822800;
      54348: inst = 32'h10a00000;
      54349: inst = 32'hca00004;
      54350: inst = 32'h38632800;
      54351: inst = 32'h38842800;
      54352: inst = 32'h10a00000;
      54353: inst = 32'hca0d455;
      54354: inst = 32'h13e00001;
      54355: inst = 32'hfe0d96a;
      54356: inst = 32'h5be00000;
      54357: inst = 32'h8c50000;
      54358: inst = 32'h24612800;
      54359: inst = 32'h10a0ffff;
      54360: inst = 32'hca0ffee;
      54361: inst = 32'h24822800;
      54362: inst = 32'h10a00000;
      54363: inst = 32'hca00004;
      54364: inst = 32'h38632800;
      54365: inst = 32'h38842800;
      54366: inst = 32'h10a00000;
      54367: inst = 32'hca0d463;
      54368: inst = 32'h13e00001;
      54369: inst = 32'hfe0d96a;
      54370: inst = 32'h5be00000;
      54371: inst = 32'h8c50000;
      54372: inst = 32'h24612800;
      54373: inst = 32'h10a0ffff;
      54374: inst = 32'hca0ffee;
      54375: inst = 32'h24822800;
      54376: inst = 32'h10a00000;
      54377: inst = 32'hca00004;
      54378: inst = 32'h38632800;
      54379: inst = 32'h38842800;
      54380: inst = 32'h10a00000;
      54381: inst = 32'hca0d471;
      54382: inst = 32'h13e00001;
      54383: inst = 32'hfe0d96a;
      54384: inst = 32'h5be00000;
      54385: inst = 32'h8c50000;
      54386: inst = 32'h24612800;
      54387: inst = 32'h10a0ffff;
      54388: inst = 32'hca0ffee;
      54389: inst = 32'h24822800;
      54390: inst = 32'h10a00000;
      54391: inst = 32'hca00004;
      54392: inst = 32'h38632800;
      54393: inst = 32'h38842800;
      54394: inst = 32'h10a00000;
      54395: inst = 32'hca0d47f;
      54396: inst = 32'h13e00001;
      54397: inst = 32'hfe0d96a;
      54398: inst = 32'h5be00000;
      54399: inst = 32'h8c50000;
      54400: inst = 32'h24612800;
      54401: inst = 32'h10a0ffff;
      54402: inst = 32'hca0ffee;
      54403: inst = 32'h24822800;
      54404: inst = 32'h10a00000;
      54405: inst = 32'hca00004;
      54406: inst = 32'h38632800;
      54407: inst = 32'h38842800;
      54408: inst = 32'h10a00000;
      54409: inst = 32'hca0d48d;
      54410: inst = 32'h13e00001;
      54411: inst = 32'hfe0d96a;
      54412: inst = 32'h5be00000;
      54413: inst = 32'h8c50000;
      54414: inst = 32'h24612800;
      54415: inst = 32'h10a0ffff;
      54416: inst = 32'hca0ffee;
      54417: inst = 32'h24822800;
      54418: inst = 32'h10a00000;
      54419: inst = 32'hca00004;
      54420: inst = 32'h38632800;
      54421: inst = 32'h38842800;
      54422: inst = 32'h10a00000;
      54423: inst = 32'hca0d49b;
      54424: inst = 32'h13e00001;
      54425: inst = 32'hfe0d96a;
      54426: inst = 32'h5be00000;
      54427: inst = 32'h8c50000;
      54428: inst = 32'h24612800;
      54429: inst = 32'h10a0ffff;
      54430: inst = 32'hca0ffee;
      54431: inst = 32'h24822800;
      54432: inst = 32'h10a00000;
      54433: inst = 32'hca00004;
      54434: inst = 32'h38632800;
      54435: inst = 32'h38842800;
      54436: inst = 32'h10a00000;
      54437: inst = 32'hca0d4a9;
      54438: inst = 32'h13e00001;
      54439: inst = 32'hfe0d96a;
      54440: inst = 32'h5be00000;
      54441: inst = 32'h8c50000;
      54442: inst = 32'h24612800;
      54443: inst = 32'h10a0ffff;
      54444: inst = 32'hca0ffee;
      54445: inst = 32'h24822800;
      54446: inst = 32'h10a00000;
      54447: inst = 32'hca00004;
      54448: inst = 32'h38632800;
      54449: inst = 32'h38842800;
      54450: inst = 32'h10a00000;
      54451: inst = 32'hca0d4b7;
      54452: inst = 32'h13e00001;
      54453: inst = 32'hfe0d96a;
      54454: inst = 32'h5be00000;
      54455: inst = 32'h8c50000;
      54456: inst = 32'h24612800;
      54457: inst = 32'h10a0ffff;
      54458: inst = 32'hca0ffee;
      54459: inst = 32'h24822800;
      54460: inst = 32'h10a00000;
      54461: inst = 32'hca00004;
      54462: inst = 32'h38632800;
      54463: inst = 32'h38842800;
      54464: inst = 32'h10a00000;
      54465: inst = 32'hca0d4c5;
      54466: inst = 32'h13e00001;
      54467: inst = 32'hfe0d96a;
      54468: inst = 32'h5be00000;
      54469: inst = 32'h8c50000;
      54470: inst = 32'h24612800;
      54471: inst = 32'h10a0ffff;
      54472: inst = 32'hca0ffee;
      54473: inst = 32'h24822800;
      54474: inst = 32'h10a00000;
      54475: inst = 32'hca00004;
      54476: inst = 32'h38632800;
      54477: inst = 32'h38842800;
      54478: inst = 32'h10a00000;
      54479: inst = 32'hca0d4d3;
      54480: inst = 32'h13e00001;
      54481: inst = 32'hfe0d96a;
      54482: inst = 32'h5be00000;
      54483: inst = 32'h8c50000;
      54484: inst = 32'h24612800;
      54485: inst = 32'h10a0ffff;
      54486: inst = 32'hca0ffee;
      54487: inst = 32'h24822800;
      54488: inst = 32'h10a00000;
      54489: inst = 32'hca00004;
      54490: inst = 32'h38632800;
      54491: inst = 32'h38842800;
      54492: inst = 32'h10a00000;
      54493: inst = 32'hca0d4e1;
      54494: inst = 32'h13e00001;
      54495: inst = 32'hfe0d96a;
      54496: inst = 32'h5be00000;
      54497: inst = 32'h8c50000;
      54498: inst = 32'h24612800;
      54499: inst = 32'h10a0ffff;
      54500: inst = 32'hca0ffee;
      54501: inst = 32'h24822800;
      54502: inst = 32'h10a00000;
      54503: inst = 32'hca00004;
      54504: inst = 32'h38632800;
      54505: inst = 32'h38842800;
      54506: inst = 32'h10a00000;
      54507: inst = 32'hca0d4ef;
      54508: inst = 32'h13e00001;
      54509: inst = 32'hfe0d96a;
      54510: inst = 32'h5be00000;
      54511: inst = 32'h8c50000;
      54512: inst = 32'h24612800;
      54513: inst = 32'h10a0ffff;
      54514: inst = 32'hca0ffee;
      54515: inst = 32'h24822800;
      54516: inst = 32'h10a00000;
      54517: inst = 32'hca00004;
      54518: inst = 32'h38632800;
      54519: inst = 32'h38842800;
      54520: inst = 32'h10a00000;
      54521: inst = 32'hca0d4fd;
      54522: inst = 32'h13e00001;
      54523: inst = 32'hfe0d96a;
      54524: inst = 32'h5be00000;
      54525: inst = 32'h8c50000;
      54526: inst = 32'h24612800;
      54527: inst = 32'h10a0ffff;
      54528: inst = 32'hca0ffee;
      54529: inst = 32'h24822800;
      54530: inst = 32'h10a00000;
      54531: inst = 32'hca00004;
      54532: inst = 32'h38632800;
      54533: inst = 32'h38842800;
      54534: inst = 32'h10a00000;
      54535: inst = 32'hca0d50b;
      54536: inst = 32'h13e00001;
      54537: inst = 32'hfe0d96a;
      54538: inst = 32'h5be00000;
      54539: inst = 32'h8c50000;
      54540: inst = 32'h24612800;
      54541: inst = 32'h10a0ffff;
      54542: inst = 32'hca0ffee;
      54543: inst = 32'h24822800;
      54544: inst = 32'h10a00000;
      54545: inst = 32'hca00004;
      54546: inst = 32'h38632800;
      54547: inst = 32'h38842800;
      54548: inst = 32'h10a00000;
      54549: inst = 32'hca0d519;
      54550: inst = 32'h13e00001;
      54551: inst = 32'hfe0d96a;
      54552: inst = 32'h5be00000;
      54553: inst = 32'h8c50000;
      54554: inst = 32'h24612800;
      54555: inst = 32'h10a0ffff;
      54556: inst = 32'hca0ffee;
      54557: inst = 32'h24822800;
      54558: inst = 32'h10a00000;
      54559: inst = 32'hca00004;
      54560: inst = 32'h38632800;
      54561: inst = 32'h38842800;
      54562: inst = 32'h10a00000;
      54563: inst = 32'hca0d527;
      54564: inst = 32'h13e00001;
      54565: inst = 32'hfe0d96a;
      54566: inst = 32'h5be00000;
      54567: inst = 32'h8c50000;
      54568: inst = 32'h24612800;
      54569: inst = 32'h10a0ffff;
      54570: inst = 32'hca0ffee;
      54571: inst = 32'h24822800;
      54572: inst = 32'h10a00000;
      54573: inst = 32'hca00004;
      54574: inst = 32'h38632800;
      54575: inst = 32'h38842800;
      54576: inst = 32'h10a00000;
      54577: inst = 32'hca0d535;
      54578: inst = 32'h13e00001;
      54579: inst = 32'hfe0d96a;
      54580: inst = 32'h5be00000;
      54581: inst = 32'h8c50000;
      54582: inst = 32'h24612800;
      54583: inst = 32'h10a0ffff;
      54584: inst = 32'hca0ffee;
      54585: inst = 32'h24822800;
      54586: inst = 32'h10a00000;
      54587: inst = 32'hca00004;
      54588: inst = 32'h38632800;
      54589: inst = 32'h38842800;
      54590: inst = 32'h10a00000;
      54591: inst = 32'hca0d543;
      54592: inst = 32'h13e00001;
      54593: inst = 32'hfe0d96a;
      54594: inst = 32'h5be00000;
      54595: inst = 32'h8c50000;
      54596: inst = 32'h24612800;
      54597: inst = 32'h10a0ffff;
      54598: inst = 32'hca0ffee;
      54599: inst = 32'h24822800;
      54600: inst = 32'h10a00000;
      54601: inst = 32'hca00004;
      54602: inst = 32'h38632800;
      54603: inst = 32'h38842800;
      54604: inst = 32'h10a00000;
      54605: inst = 32'hca0d551;
      54606: inst = 32'h13e00001;
      54607: inst = 32'hfe0d96a;
      54608: inst = 32'h5be00000;
      54609: inst = 32'h8c50000;
      54610: inst = 32'h24612800;
      54611: inst = 32'h10a0ffff;
      54612: inst = 32'hca0ffee;
      54613: inst = 32'h24822800;
      54614: inst = 32'h10a00000;
      54615: inst = 32'hca00004;
      54616: inst = 32'h38632800;
      54617: inst = 32'h38842800;
      54618: inst = 32'h10a00000;
      54619: inst = 32'hca0d55f;
      54620: inst = 32'h13e00001;
      54621: inst = 32'hfe0d96a;
      54622: inst = 32'h5be00000;
      54623: inst = 32'h8c50000;
      54624: inst = 32'h24612800;
      54625: inst = 32'h10a0ffff;
      54626: inst = 32'hca0ffee;
      54627: inst = 32'h24822800;
      54628: inst = 32'h10a00000;
      54629: inst = 32'hca00004;
      54630: inst = 32'h38632800;
      54631: inst = 32'h38842800;
      54632: inst = 32'h10a00000;
      54633: inst = 32'hca0d56d;
      54634: inst = 32'h13e00001;
      54635: inst = 32'hfe0d96a;
      54636: inst = 32'h5be00000;
      54637: inst = 32'h8c50000;
      54638: inst = 32'h24612800;
      54639: inst = 32'h10a0ffff;
      54640: inst = 32'hca0ffee;
      54641: inst = 32'h24822800;
      54642: inst = 32'h10a00000;
      54643: inst = 32'hca00004;
      54644: inst = 32'h38632800;
      54645: inst = 32'h38842800;
      54646: inst = 32'h10a00000;
      54647: inst = 32'hca0d57b;
      54648: inst = 32'h13e00001;
      54649: inst = 32'hfe0d96a;
      54650: inst = 32'h5be00000;
      54651: inst = 32'h8c50000;
      54652: inst = 32'h24612800;
      54653: inst = 32'h10a0ffff;
      54654: inst = 32'hca0ffee;
      54655: inst = 32'h24822800;
      54656: inst = 32'h10a00000;
      54657: inst = 32'hca00004;
      54658: inst = 32'h38632800;
      54659: inst = 32'h38842800;
      54660: inst = 32'h10a00000;
      54661: inst = 32'hca0d589;
      54662: inst = 32'h13e00001;
      54663: inst = 32'hfe0d96a;
      54664: inst = 32'h5be00000;
      54665: inst = 32'h8c50000;
      54666: inst = 32'h24612800;
      54667: inst = 32'h10a0ffff;
      54668: inst = 32'hca0ffee;
      54669: inst = 32'h24822800;
      54670: inst = 32'h10a00000;
      54671: inst = 32'hca00004;
      54672: inst = 32'h38632800;
      54673: inst = 32'h38842800;
      54674: inst = 32'h10a00000;
      54675: inst = 32'hca0d597;
      54676: inst = 32'h13e00001;
      54677: inst = 32'hfe0d96a;
      54678: inst = 32'h5be00000;
      54679: inst = 32'h8c50000;
      54680: inst = 32'h24612800;
      54681: inst = 32'h10a0ffff;
      54682: inst = 32'hca0ffee;
      54683: inst = 32'h24822800;
      54684: inst = 32'h10a00000;
      54685: inst = 32'hca00004;
      54686: inst = 32'h38632800;
      54687: inst = 32'h38842800;
      54688: inst = 32'h10a00000;
      54689: inst = 32'hca0d5a5;
      54690: inst = 32'h13e00001;
      54691: inst = 32'hfe0d96a;
      54692: inst = 32'h5be00000;
      54693: inst = 32'h8c50000;
      54694: inst = 32'h24612800;
      54695: inst = 32'h10a0ffff;
      54696: inst = 32'hca0ffee;
      54697: inst = 32'h24822800;
      54698: inst = 32'h10a00000;
      54699: inst = 32'hca00004;
      54700: inst = 32'h38632800;
      54701: inst = 32'h38842800;
      54702: inst = 32'h10a00000;
      54703: inst = 32'hca0d5b3;
      54704: inst = 32'h13e00001;
      54705: inst = 32'hfe0d96a;
      54706: inst = 32'h5be00000;
      54707: inst = 32'h8c50000;
      54708: inst = 32'h24612800;
      54709: inst = 32'h10a0ffff;
      54710: inst = 32'hca0ffee;
      54711: inst = 32'h24822800;
      54712: inst = 32'h10a00000;
      54713: inst = 32'hca00004;
      54714: inst = 32'h38632800;
      54715: inst = 32'h38842800;
      54716: inst = 32'h10a00000;
      54717: inst = 32'hca0d5c1;
      54718: inst = 32'h13e00001;
      54719: inst = 32'hfe0d96a;
      54720: inst = 32'h5be00000;
      54721: inst = 32'h8c50000;
      54722: inst = 32'h24612800;
      54723: inst = 32'h10a0ffff;
      54724: inst = 32'hca0ffee;
      54725: inst = 32'h24822800;
      54726: inst = 32'h10a00000;
      54727: inst = 32'hca00004;
      54728: inst = 32'h38632800;
      54729: inst = 32'h38842800;
      54730: inst = 32'h10a00000;
      54731: inst = 32'hca0d5cf;
      54732: inst = 32'h13e00001;
      54733: inst = 32'hfe0d96a;
      54734: inst = 32'h5be00000;
      54735: inst = 32'h8c50000;
      54736: inst = 32'h24612800;
      54737: inst = 32'h10a0ffff;
      54738: inst = 32'hca0ffee;
      54739: inst = 32'h24822800;
      54740: inst = 32'h10a00000;
      54741: inst = 32'hca00004;
      54742: inst = 32'h38632800;
      54743: inst = 32'h38842800;
      54744: inst = 32'h10a00000;
      54745: inst = 32'hca0d5dd;
      54746: inst = 32'h13e00001;
      54747: inst = 32'hfe0d96a;
      54748: inst = 32'h5be00000;
      54749: inst = 32'h8c50000;
      54750: inst = 32'h24612800;
      54751: inst = 32'h10a0ffff;
      54752: inst = 32'hca0ffee;
      54753: inst = 32'h24822800;
      54754: inst = 32'h10a00000;
      54755: inst = 32'hca00004;
      54756: inst = 32'h38632800;
      54757: inst = 32'h38842800;
      54758: inst = 32'h10a00000;
      54759: inst = 32'hca0d5eb;
      54760: inst = 32'h13e00001;
      54761: inst = 32'hfe0d96a;
      54762: inst = 32'h5be00000;
      54763: inst = 32'h8c50000;
      54764: inst = 32'h24612800;
      54765: inst = 32'h10a0ffff;
      54766: inst = 32'hca0ffee;
      54767: inst = 32'h24822800;
      54768: inst = 32'h10a00000;
      54769: inst = 32'hca00004;
      54770: inst = 32'h38632800;
      54771: inst = 32'h38842800;
      54772: inst = 32'h10a00000;
      54773: inst = 32'hca0d5f9;
      54774: inst = 32'h13e00001;
      54775: inst = 32'hfe0d96a;
      54776: inst = 32'h5be00000;
      54777: inst = 32'h8c50000;
      54778: inst = 32'h24612800;
      54779: inst = 32'h10a0ffff;
      54780: inst = 32'hca0ffee;
      54781: inst = 32'h24822800;
      54782: inst = 32'h10a00000;
      54783: inst = 32'hca00004;
      54784: inst = 32'h38632800;
      54785: inst = 32'h38842800;
      54786: inst = 32'h10a00000;
      54787: inst = 32'hca0d607;
      54788: inst = 32'h13e00001;
      54789: inst = 32'hfe0d96a;
      54790: inst = 32'h5be00000;
      54791: inst = 32'h8c50000;
      54792: inst = 32'h24612800;
      54793: inst = 32'h10a0ffff;
      54794: inst = 32'hca0ffee;
      54795: inst = 32'h24822800;
      54796: inst = 32'h10a00000;
      54797: inst = 32'hca00004;
      54798: inst = 32'h38632800;
      54799: inst = 32'h38842800;
      54800: inst = 32'h10a00000;
      54801: inst = 32'hca0d615;
      54802: inst = 32'h13e00001;
      54803: inst = 32'hfe0d96a;
      54804: inst = 32'h5be00000;
      54805: inst = 32'h8c50000;
      54806: inst = 32'h24612800;
      54807: inst = 32'h10a0ffff;
      54808: inst = 32'hca0ffee;
      54809: inst = 32'h24822800;
      54810: inst = 32'h10a00000;
      54811: inst = 32'hca00004;
      54812: inst = 32'h38632800;
      54813: inst = 32'h38842800;
      54814: inst = 32'h10a00000;
      54815: inst = 32'hca0d623;
      54816: inst = 32'h13e00001;
      54817: inst = 32'hfe0d96a;
      54818: inst = 32'h5be00000;
      54819: inst = 32'h8c50000;
      54820: inst = 32'h24612800;
      54821: inst = 32'h10a0ffff;
      54822: inst = 32'hca0ffee;
      54823: inst = 32'h24822800;
      54824: inst = 32'h10a00000;
      54825: inst = 32'hca00004;
      54826: inst = 32'h38632800;
      54827: inst = 32'h38842800;
      54828: inst = 32'h10a00000;
      54829: inst = 32'hca0d631;
      54830: inst = 32'h13e00001;
      54831: inst = 32'hfe0d96a;
      54832: inst = 32'h5be00000;
      54833: inst = 32'h8c50000;
      54834: inst = 32'h24612800;
      54835: inst = 32'h10a0ffff;
      54836: inst = 32'hca0ffee;
      54837: inst = 32'h24822800;
      54838: inst = 32'h10a00000;
      54839: inst = 32'hca00004;
      54840: inst = 32'h38632800;
      54841: inst = 32'h38842800;
      54842: inst = 32'h10a00000;
      54843: inst = 32'hca0d63f;
      54844: inst = 32'h13e00001;
      54845: inst = 32'hfe0d96a;
      54846: inst = 32'h5be00000;
      54847: inst = 32'h8c50000;
      54848: inst = 32'h24612800;
      54849: inst = 32'h10a0ffff;
      54850: inst = 32'hca0ffee;
      54851: inst = 32'h24822800;
      54852: inst = 32'h10a00000;
      54853: inst = 32'hca00004;
      54854: inst = 32'h38632800;
      54855: inst = 32'h38842800;
      54856: inst = 32'h10a00000;
      54857: inst = 32'hca0d64d;
      54858: inst = 32'h13e00001;
      54859: inst = 32'hfe0d96a;
      54860: inst = 32'h5be00000;
      54861: inst = 32'h8c50000;
      54862: inst = 32'h24612800;
      54863: inst = 32'h10a0ffff;
      54864: inst = 32'hca0ffee;
      54865: inst = 32'h24822800;
      54866: inst = 32'h10a00000;
      54867: inst = 32'hca00004;
      54868: inst = 32'h38632800;
      54869: inst = 32'h38842800;
      54870: inst = 32'h10a00000;
      54871: inst = 32'hca0d65b;
      54872: inst = 32'h13e00001;
      54873: inst = 32'hfe0d96a;
      54874: inst = 32'h5be00000;
      54875: inst = 32'h8c50000;
      54876: inst = 32'h24612800;
      54877: inst = 32'h10a0ffff;
      54878: inst = 32'hca0ffee;
      54879: inst = 32'h24822800;
      54880: inst = 32'h10a00000;
      54881: inst = 32'hca00004;
      54882: inst = 32'h38632800;
      54883: inst = 32'h38842800;
      54884: inst = 32'h10a00000;
      54885: inst = 32'hca0d669;
      54886: inst = 32'h13e00001;
      54887: inst = 32'hfe0d96a;
      54888: inst = 32'h5be00000;
      54889: inst = 32'h8c50000;
      54890: inst = 32'h24612800;
      54891: inst = 32'h10a0ffff;
      54892: inst = 32'hca0ffee;
      54893: inst = 32'h24822800;
      54894: inst = 32'h10a00000;
      54895: inst = 32'hca00004;
      54896: inst = 32'h38632800;
      54897: inst = 32'h38842800;
      54898: inst = 32'h10a00000;
      54899: inst = 32'hca0d677;
      54900: inst = 32'h13e00001;
      54901: inst = 32'hfe0d96a;
      54902: inst = 32'h5be00000;
      54903: inst = 32'h8c50000;
      54904: inst = 32'h24612800;
      54905: inst = 32'h10a0ffff;
      54906: inst = 32'hca0ffee;
      54907: inst = 32'h24822800;
      54908: inst = 32'h10a00000;
      54909: inst = 32'hca00004;
      54910: inst = 32'h38632800;
      54911: inst = 32'h38842800;
      54912: inst = 32'h10a00000;
      54913: inst = 32'hca0d685;
      54914: inst = 32'h13e00001;
      54915: inst = 32'hfe0d96a;
      54916: inst = 32'h5be00000;
      54917: inst = 32'h8c50000;
      54918: inst = 32'h24612800;
      54919: inst = 32'h10a0ffff;
      54920: inst = 32'hca0ffee;
      54921: inst = 32'h24822800;
      54922: inst = 32'h10a00000;
      54923: inst = 32'hca00004;
      54924: inst = 32'h38632800;
      54925: inst = 32'h38842800;
      54926: inst = 32'h10a00000;
      54927: inst = 32'hca0d693;
      54928: inst = 32'h13e00001;
      54929: inst = 32'hfe0d96a;
      54930: inst = 32'h5be00000;
      54931: inst = 32'h8c50000;
      54932: inst = 32'h24612800;
      54933: inst = 32'h10a0ffff;
      54934: inst = 32'hca0ffee;
      54935: inst = 32'h24822800;
      54936: inst = 32'h10a00000;
      54937: inst = 32'hca00004;
      54938: inst = 32'h38632800;
      54939: inst = 32'h38842800;
      54940: inst = 32'h10a00000;
      54941: inst = 32'hca0d6a1;
      54942: inst = 32'h13e00001;
      54943: inst = 32'hfe0d96a;
      54944: inst = 32'h5be00000;
      54945: inst = 32'h8c50000;
      54946: inst = 32'h24612800;
      54947: inst = 32'h10a0ffff;
      54948: inst = 32'hca0ffee;
      54949: inst = 32'h24822800;
      54950: inst = 32'h10a00000;
      54951: inst = 32'hca00004;
      54952: inst = 32'h38632800;
      54953: inst = 32'h38842800;
      54954: inst = 32'h10a00000;
      54955: inst = 32'hca0d6af;
      54956: inst = 32'h13e00001;
      54957: inst = 32'hfe0d96a;
      54958: inst = 32'h5be00000;
      54959: inst = 32'h8c50000;
      54960: inst = 32'h24612800;
      54961: inst = 32'h10a0ffff;
      54962: inst = 32'hca0ffee;
      54963: inst = 32'h24822800;
      54964: inst = 32'h10a00000;
      54965: inst = 32'hca00004;
      54966: inst = 32'h38632800;
      54967: inst = 32'h38842800;
      54968: inst = 32'h10a00000;
      54969: inst = 32'hca0d6bd;
      54970: inst = 32'h13e00001;
      54971: inst = 32'hfe0d96a;
      54972: inst = 32'h5be00000;
      54973: inst = 32'h8c50000;
      54974: inst = 32'h24612800;
      54975: inst = 32'h10a0ffff;
      54976: inst = 32'hca0ffee;
      54977: inst = 32'h24822800;
      54978: inst = 32'h10a00000;
      54979: inst = 32'hca00004;
      54980: inst = 32'h38632800;
      54981: inst = 32'h38842800;
      54982: inst = 32'h10a00000;
      54983: inst = 32'hca0d6cb;
      54984: inst = 32'h13e00001;
      54985: inst = 32'hfe0d96a;
      54986: inst = 32'h5be00000;
      54987: inst = 32'h8c50000;
      54988: inst = 32'h24612800;
      54989: inst = 32'h10a0ffff;
      54990: inst = 32'hca0ffee;
      54991: inst = 32'h24822800;
      54992: inst = 32'h10a00000;
      54993: inst = 32'hca00004;
      54994: inst = 32'h38632800;
      54995: inst = 32'h38842800;
      54996: inst = 32'h10a00000;
      54997: inst = 32'hca0d6d9;
      54998: inst = 32'h13e00001;
      54999: inst = 32'hfe0d96a;
      55000: inst = 32'h5be00000;
      55001: inst = 32'h8c50000;
      55002: inst = 32'h24612800;
      55003: inst = 32'h10a0ffff;
      55004: inst = 32'hca0ffee;
      55005: inst = 32'h24822800;
      55006: inst = 32'h10a00000;
      55007: inst = 32'hca00004;
      55008: inst = 32'h38632800;
      55009: inst = 32'h38842800;
      55010: inst = 32'h10a00000;
      55011: inst = 32'hca0d6e7;
      55012: inst = 32'h13e00001;
      55013: inst = 32'hfe0d96a;
      55014: inst = 32'h5be00000;
      55015: inst = 32'h8c50000;
      55016: inst = 32'h24612800;
      55017: inst = 32'h10a0ffff;
      55018: inst = 32'hca0ffee;
      55019: inst = 32'h24822800;
      55020: inst = 32'h10a00000;
      55021: inst = 32'hca00004;
      55022: inst = 32'h38632800;
      55023: inst = 32'h38842800;
      55024: inst = 32'h10a00000;
      55025: inst = 32'hca0d6f5;
      55026: inst = 32'h13e00001;
      55027: inst = 32'hfe0d96a;
      55028: inst = 32'h5be00000;
      55029: inst = 32'h8c50000;
      55030: inst = 32'h24612800;
      55031: inst = 32'h10a0ffff;
      55032: inst = 32'hca0ffee;
      55033: inst = 32'h24822800;
      55034: inst = 32'h10a00000;
      55035: inst = 32'hca00004;
      55036: inst = 32'h38632800;
      55037: inst = 32'h38842800;
      55038: inst = 32'h10a00000;
      55039: inst = 32'hca0d703;
      55040: inst = 32'h13e00001;
      55041: inst = 32'hfe0d96a;
      55042: inst = 32'h5be00000;
      55043: inst = 32'h8c50000;
      55044: inst = 32'h24612800;
      55045: inst = 32'h10a0ffff;
      55046: inst = 32'hca0ffee;
      55047: inst = 32'h24822800;
      55048: inst = 32'h10a00000;
      55049: inst = 32'hca00004;
      55050: inst = 32'h38632800;
      55051: inst = 32'h38842800;
      55052: inst = 32'h10a00000;
      55053: inst = 32'hca0d711;
      55054: inst = 32'h13e00001;
      55055: inst = 32'hfe0d96a;
      55056: inst = 32'h5be00000;
      55057: inst = 32'h8c50000;
      55058: inst = 32'h24612800;
      55059: inst = 32'h10a0ffff;
      55060: inst = 32'hca0ffee;
      55061: inst = 32'h24822800;
      55062: inst = 32'h10a00000;
      55063: inst = 32'hca00004;
      55064: inst = 32'h38632800;
      55065: inst = 32'h38842800;
      55066: inst = 32'h10a00000;
      55067: inst = 32'hca0d71f;
      55068: inst = 32'h13e00001;
      55069: inst = 32'hfe0d96a;
      55070: inst = 32'h5be00000;
      55071: inst = 32'h8c50000;
      55072: inst = 32'h24612800;
      55073: inst = 32'h10a0ffff;
      55074: inst = 32'hca0ffee;
      55075: inst = 32'h24822800;
      55076: inst = 32'h10a00000;
      55077: inst = 32'hca00004;
      55078: inst = 32'h38632800;
      55079: inst = 32'h38842800;
      55080: inst = 32'h10a00000;
      55081: inst = 32'hca0d72d;
      55082: inst = 32'h13e00001;
      55083: inst = 32'hfe0d96a;
      55084: inst = 32'h5be00000;
      55085: inst = 32'h8c50000;
      55086: inst = 32'h24612800;
      55087: inst = 32'h10a0ffff;
      55088: inst = 32'hca0ffee;
      55089: inst = 32'h24822800;
      55090: inst = 32'h10a00000;
      55091: inst = 32'hca00004;
      55092: inst = 32'h38632800;
      55093: inst = 32'h38842800;
      55094: inst = 32'h10a00000;
      55095: inst = 32'hca0d73b;
      55096: inst = 32'h13e00001;
      55097: inst = 32'hfe0d96a;
      55098: inst = 32'h5be00000;
      55099: inst = 32'h8c50000;
      55100: inst = 32'h24612800;
      55101: inst = 32'h10a0ffff;
      55102: inst = 32'hca0ffee;
      55103: inst = 32'h24822800;
      55104: inst = 32'h10a00000;
      55105: inst = 32'hca00004;
      55106: inst = 32'h38632800;
      55107: inst = 32'h38842800;
      55108: inst = 32'h10a00000;
      55109: inst = 32'hca0d749;
      55110: inst = 32'h13e00001;
      55111: inst = 32'hfe0d96a;
      55112: inst = 32'h5be00000;
      55113: inst = 32'h8c50000;
      55114: inst = 32'h24612800;
      55115: inst = 32'h10a0ffff;
      55116: inst = 32'hca0ffee;
      55117: inst = 32'h24822800;
      55118: inst = 32'h10a00000;
      55119: inst = 32'hca00004;
      55120: inst = 32'h38632800;
      55121: inst = 32'h38842800;
      55122: inst = 32'h10a00000;
      55123: inst = 32'hca0d757;
      55124: inst = 32'h13e00001;
      55125: inst = 32'hfe0d96a;
      55126: inst = 32'h5be00000;
      55127: inst = 32'h8c50000;
      55128: inst = 32'h24612800;
      55129: inst = 32'h10a0ffff;
      55130: inst = 32'hca0ffee;
      55131: inst = 32'h24822800;
      55132: inst = 32'h10a00000;
      55133: inst = 32'hca00004;
      55134: inst = 32'h38632800;
      55135: inst = 32'h38842800;
      55136: inst = 32'h10a00000;
      55137: inst = 32'hca0d765;
      55138: inst = 32'h13e00001;
      55139: inst = 32'hfe0d96a;
      55140: inst = 32'h5be00000;
      55141: inst = 32'h8c50000;
      55142: inst = 32'h24612800;
      55143: inst = 32'h10a0ffff;
      55144: inst = 32'hca0ffee;
      55145: inst = 32'h24822800;
      55146: inst = 32'h10a00000;
      55147: inst = 32'hca00004;
      55148: inst = 32'h38632800;
      55149: inst = 32'h38842800;
      55150: inst = 32'h10a00000;
      55151: inst = 32'hca0d773;
      55152: inst = 32'h13e00001;
      55153: inst = 32'hfe0d96a;
      55154: inst = 32'h5be00000;
      55155: inst = 32'h8c50000;
      55156: inst = 32'h24612800;
      55157: inst = 32'h10a0ffff;
      55158: inst = 32'hca0ffee;
      55159: inst = 32'h24822800;
      55160: inst = 32'h10a00000;
      55161: inst = 32'hca00004;
      55162: inst = 32'h38632800;
      55163: inst = 32'h38842800;
      55164: inst = 32'h10a00000;
      55165: inst = 32'hca0d781;
      55166: inst = 32'h13e00001;
      55167: inst = 32'hfe0d96a;
      55168: inst = 32'h5be00000;
      55169: inst = 32'h8c50000;
      55170: inst = 32'h24612800;
      55171: inst = 32'h10a0ffff;
      55172: inst = 32'hca0ffee;
      55173: inst = 32'h24822800;
      55174: inst = 32'h10a00000;
      55175: inst = 32'hca00004;
      55176: inst = 32'h38632800;
      55177: inst = 32'h38842800;
      55178: inst = 32'h10a00000;
      55179: inst = 32'hca0d78f;
      55180: inst = 32'h13e00001;
      55181: inst = 32'hfe0d96a;
      55182: inst = 32'h5be00000;
      55183: inst = 32'h8c50000;
      55184: inst = 32'h24612800;
      55185: inst = 32'h10a0ffff;
      55186: inst = 32'hca0ffee;
      55187: inst = 32'h24822800;
      55188: inst = 32'h10a00000;
      55189: inst = 32'hca00004;
      55190: inst = 32'h38632800;
      55191: inst = 32'h38842800;
      55192: inst = 32'h10a00000;
      55193: inst = 32'hca0d79d;
      55194: inst = 32'h13e00001;
      55195: inst = 32'hfe0d96a;
      55196: inst = 32'h5be00000;
      55197: inst = 32'h8c50000;
      55198: inst = 32'h24612800;
      55199: inst = 32'h10a0ffff;
      55200: inst = 32'hca0ffee;
      55201: inst = 32'h24822800;
      55202: inst = 32'h10a00000;
      55203: inst = 32'hca00004;
      55204: inst = 32'h38632800;
      55205: inst = 32'h38842800;
      55206: inst = 32'h10a00000;
      55207: inst = 32'hca0d7ab;
      55208: inst = 32'h13e00001;
      55209: inst = 32'hfe0d96a;
      55210: inst = 32'h5be00000;
      55211: inst = 32'h8c50000;
      55212: inst = 32'h24612800;
      55213: inst = 32'h10a0ffff;
      55214: inst = 32'hca0ffee;
      55215: inst = 32'h24822800;
      55216: inst = 32'h10a00000;
      55217: inst = 32'hca00004;
      55218: inst = 32'h38632800;
      55219: inst = 32'h38842800;
      55220: inst = 32'h10a00000;
      55221: inst = 32'hca0d7b9;
      55222: inst = 32'h13e00001;
      55223: inst = 32'hfe0d96a;
      55224: inst = 32'h5be00000;
      55225: inst = 32'h8c50000;
      55226: inst = 32'h24612800;
      55227: inst = 32'h10a0ffff;
      55228: inst = 32'hca0ffee;
      55229: inst = 32'h24822800;
      55230: inst = 32'h10a00000;
      55231: inst = 32'hca00004;
      55232: inst = 32'h38632800;
      55233: inst = 32'h38842800;
      55234: inst = 32'h10a00000;
      55235: inst = 32'hca0d7c7;
      55236: inst = 32'h13e00001;
      55237: inst = 32'hfe0d96a;
      55238: inst = 32'h5be00000;
      55239: inst = 32'h8c50000;
      55240: inst = 32'h24612800;
      55241: inst = 32'h10a0ffff;
      55242: inst = 32'hca0ffee;
      55243: inst = 32'h24822800;
      55244: inst = 32'h10a00000;
      55245: inst = 32'hca00004;
      55246: inst = 32'h38632800;
      55247: inst = 32'h38842800;
      55248: inst = 32'h10a00000;
      55249: inst = 32'hca0d7d5;
      55250: inst = 32'h13e00001;
      55251: inst = 32'hfe0d96a;
      55252: inst = 32'h5be00000;
      55253: inst = 32'h8c50000;
      55254: inst = 32'h24612800;
      55255: inst = 32'h10a0ffff;
      55256: inst = 32'hca0ffee;
      55257: inst = 32'h24822800;
      55258: inst = 32'h10a00000;
      55259: inst = 32'hca00004;
      55260: inst = 32'h38632800;
      55261: inst = 32'h38842800;
      55262: inst = 32'h10a00000;
      55263: inst = 32'hca0d7e3;
      55264: inst = 32'h13e00001;
      55265: inst = 32'hfe0d96a;
      55266: inst = 32'h5be00000;
      55267: inst = 32'h8c50000;
      55268: inst = 32'h24612800;
      55269: inst = 32'h10a0ffff;
      55270: inst = 32'hca0ffee;
      55271: inst = 32'h24822800;
      55272: inst = 32'h10a00000;
      55273: inst = 32'hca00004;
      55274: inst = 32'h38632800;
      55275: inst = 32'h38842800;
      55276: inst = 32'h10a00000;
      55277: inst = 32'hca0d7f1;
      55278: inst = 32'h13e00001;
      55279: inst = 32'hfe0d96a;
      55280: inst = 32'h5be00000;
      55281: inst = 32'h8c50000;
      55282: inst = 32'h24612800;
      55283: inst = 32'h10a0ffff;
      55284: inst = 32'hca0ffee;
      55285: inst = 32'h24822800;
      55286: inst = 32'h10a00000;
      55287: inst = 32'hca00004;
      55288: inst = 32'h38632800;
      55289: inst = 32'h38842800;
      55290: inst = 32'h10a00000;
      55291: inst = 32'hca0d7ff;
      55292: inst = 32'h13e00001;
      55293: inst = 32'hfe0d96a;
      55294: inst = 32'h5be00000;
      55295: inst = 32'h8c50000;
      55296: inst = 32'h24612800;
      55297: inst = 32'h10a0ffff;
      55298: inst = 32'hca0ffee;
      55299: inst = 32'h24822800;
      55300: inst = 32'h10a00000;
      55301: inst = 32'hca00004;
      55302: inst = 32'h38632800;
      55303: inst = 32'h38842800;
      55304: inst = 32'h10a00000;
      55305: inst = 32'hca0d80d;
      55306: inst = 32'h13e00001;
      55307: inst = 32'hfe0d96a;
      55308: inst = 32'h5be00000;
      55309: inst = 32'h8c50000;
      55310: inst = 32'h24612800;
      55311: inst = 32'h10a0ffff;
      55312: inst = 32'hca0ffee;
      55313: inst = 32'h24822800;
      55314: inst = 32'h10a00000;
      55315: inst = 32'hca00004;
      55316: inst = 32'h38632800;
      55317: inst = 32'h38842800;
      55318: inst = 32'h10a00000;
      55319: inst = 32'hca0d81b;
      55320: inst = 32'h13e00001;
      55321: inst = 32'hfe0d96a;
      55322: inst = 32'h5be00000;
      55323: inst = 32'h8c50000;
      55324: inst = 32'h24612800;
      55325: inst = 32'h10a0ffff;
      55326: inst = 32'hca0ffee;
      55327: inst = 32'h24822800;
      55328: inst = 32'h10a00000;
      55329: inst = 32'hca00004;
      55330: inst = 32'h38632800;
      55331: inst = 32'h38842800;
      55332: inst = 32'h10a00000;
      55333: inst = 32'hca0d829;
      55334: inst = 32'h13e00001;
      55335: inst = 32'hfe0d96a;
      55336: inst = 32'h5be00000;
      55337: inst = 32'h8c50000;
      55338: inst = 32'h24612800;
      55339: inst = 32'h10a0ffff;
      55340: inst = 32'hca0ffef;
      55341: inst = 32'h24822800;
      55342: inst = 32'h10a00000;
      55343: inst = 32'hca00004;
      55344: inst = 32'h38632800;
      55345: inst = 32'h38842800;
      55346: inst = 32'h10a00000;
      55347: inst = 32'hca0d837;
      55348: inst = 32'h13e00001;
      55349: inst = 32'hfe0d96a;
      55350: inst = 32'h5be00000;
      55351: inst = 32'h8c50000;
      55352: inst = 32'h24612800;
      55353: inst = 32'h10a0ffff;
      55354: inst = 32'hca0ffef;
      55355: inst = 32'h24822800;
      55356: inst = 32'h10a00000;
      55357: inst = 32'hca00004;
      55358: inst = 32'h38632800;
      55359: inst = 32'h38842800;
      55360: inst = 32'h10a00000;
      55361: inst = 32'hca0d845;
      55362: inst = 32'h13e00001;
      55363: inst = 32'hfe0d96a;
      55364: inst = 32'h5be00000;
      55365: inst = 32'h8c50000;
      55366: inst = 32'h24612800;
      55367: inst = 32'h10a0ffff;
      55368: inst = 32'hca0ffef;
      55369: inst = 32'h24822800;
      55370: inst = 32'h10a00000;
      55371: inst = 32'hca00004;
      55372: inst = 32'h38632800;
      55373: inst = 32'h38842800;
      55374: inst = 32'h10a00000;
      55375: inst = 32'hca0d853;
      55376: inst = 32'h13e00001;
      55377: inst = 32'hfe0d96a;
      55378: inst = 32'h5be00000;
      55379: inst = 32'h8c50000;
      55380: inst = 32'h24612800;
      55381: inst = 32'h10a0ffff;
      55382: inst = 32'hca0ffef;
      55383: inst = 32'h24822800;
      55384: inst = 32'h10a00000;
      55385: inst = 32'hca00004;
      55386: inst = 32'h38632800;
      55387: inst = 32'h38842800;
      55388: inst = 32'h10a00000;
      55389: inst = 32'hca0d861;
      55390: inst = 32'h13e00001;
      55391: inst = 32'hfe0d96a;
      55392: inst = 32'h5be00000;
      55393: inst = 32'h8c50000;
      55394: inst = 32'h24612800;
      55395: inst = 32'h10a0ffff;
      55396: inst = 32'hca0ffef;
      55397: inst = 32'h24822800;
      55398: inst = 32'h10a00000;
      55399: inst = 32'hca00004;
      55400: inst = 32'h38632800;
      55401: inst = 32'h38842800;
      55402: inst = 32'h10a00000;
      55403: inst = 32'hca0d86f;
      55404: inst = 32'h13e00001;
      55405: inst = 32'hfe0d96a;
      55406: inst = 32'h5be00000;
      55407: inst = 32'h8c50000;
      55408: inst = 32'h24612800;
      55409: inst = 32'h10a0ffff;
      55410: inst = 32'hca0ffef;
      55411: inst = 32'h24822800;
      55412: inst = 32'h10a00000;
      55413: inst = 32'hca00004;
      55414: inst = 32'h38632800;
      55415: inst = 32'h38842800;
      55416: inst = 32'h10a00000;
      55417: inst = 32'hca0d87d;
      55418: inst = 32'h13e00001;
      55419: inst = 32'hfe0d96a;
      55420: inst = 32'h5be00000;
      55421: inst = 32'h8c50000;
      55422: inst = 32'h24612800;
      55423: inst = 32'h10a0ffff;
      55424: inst = 32'hca0ffef;
      55425: inst = 32'h24822800;
      55426: inst = 32'h10a00000;
      55427: inst = 32'hca00004;
      55428: inst = 32'h38632800;
      55429: inst = 32'h38842800;
      55430: inst = 32'h10a00000;
      55431: inst = 32'hca0d88b;
      55432: inst = 32'h13e00001;
      55433: inst = 32'hfe0d96a;
      55434: inst = 32'h5be00000;
      55435: inst = 32'h8c50000;
      55436: inst = 32'h24612800;
      55437: inst = 32'h10a0ffff;
      55438: inst = 32'hca0ffef;
      55439: inst = 32'h24822800;
      55440: inst = 32'h10a00000;
      55441: inst = 32'hca00004;
      55442: inst = 32'h38632800;
      55443: inst = 32'h38842800;
      55444: inst = 32'h10a00000;
      55445: inst = 32'hca0d899;
      55446: inst = 32'h13e00001;
      55447: inst = 32'hfe0d96a;
      55448: inst = 32'h5be00000;
      55449: inst = 32'h8c50000;
      55450: inst = 32'h24612800;
      55451: inst = 32'h10a0ffff;
      55452: inst = 32'hca0ffef;
      55453: inst = 32'h24822800;
      55454: inst = 32'h10a00000;
      55455: inst = 32'hca00004;
      55456: inst = 32'h38632800;
      55457: inst = 32'h38842800;
      55458: inst = 32'h10a00000;
      55459: inst = 32'hca0d8a7;
      55460: inst = 32'h13e00001;
      55461: inst = 32'hfe0d96a;
      55462: inst = 32'h5be00000;
      55463: inst = 32'h8c50000;
      55464: inst = 32'h24612800;
      55465: inst = 32'h10a0ffff;
      55466: inst = 32'hca0ffef;
      55467: inst = 32'h24822800;
      55468: inst = 32'h10a00000;
      55469: inst = 32'hca00004;
      55470: inst = 32'h38632800;
      55471: inst = 32'h38842800;
      55472: inst = 32'h10a00000;
      55473: inst = 32'hca0d8b5;
      55474: inst = 32'h13e00001;
      55475: inst = 32'hfe0d96a;
      55476: inst = 32'h5be00000;
      55477: inst = 32'h8c50000;
      55478: inst = 32'h24612800;
      55479: inst = 32'h10a0ffff;
      55480: inst = 32'hca0ffef;
      55481: inst = 32'h24822800;
      55482: inst = 32'h10a00000;
      55483: inst = 32'hca00004;
      55484: inst = 32'h38632800;
      55485: inst = 32'h38842800;
      55486: inst = 32'h10a00000;
      55487: inst = 32'hca0d8c3;
      55488: inst = 32'h13e00001;
      55489: inst = 32'hfe0d96a;
      55490: inst = 32'h5be00000;
      55491: inst = 32'h8c50000;
      55492: inst = 32'h24612800;
      55493: inst = 32'h10a0ffff;
      55494: inst = 32'hca0ffef;
      55495: inst = 32'h24822800;
      55496: inst = 32'h10a00000;
      55497: inst = 32'hca00004;
      55498: inst = 32'h38632800;
      55499: inst = 32'h38842800;
      55500: inst = 32'h10a00000;
      55501: inst = 32'hca0d8d1;
      55502: inst = 32'h13e00001;
      55503: inst = 32'hfe0d96a;
      55504: inst = 32'h5be00000;
      55505: inst = 32'h8c50000;
      55506: inst = 32'h24612800;
      55507: inst = 32'h10a0ffff;
      55508: inst = 32'hca0ffef;
      55509: inst = 32'h24822800;
      55510: inst = 32'h10a00000;
      55511: inst = 32'hca00004;
      55512: inst = 32'h38632800;
      55513: inst = 32'h38842800;
      55514: inst = 32'h10a00000;
      55515: inst = 32'hca0d8df;
      55516: inst = 32'h13e00001;
      55517: inst = 32'hfe0d96a;
      55518: inst = 32'h5be00000;
      55519: inst = 32'h8c50000;
      55520: inst = 32'h24612800;
      55521: inst = 32'h10a0ffff;
      55522: inst = 32'hca0ffef;
      55523: inst = 32'h24822800;
      55524: inst = 32'h10a00000;
      55525: inst = 32'hca00004;
      55526: inst = 32'h38632800;
      55527: inst = 32'h38842800;
      55528: inst = 32'h10a00000;
      55529: inst = 32'hca0d8ed;
      55530: inst = 32'h13e00001;
      55531: inst = 32'hfe0d96a;
      55532: inst = 32'h5be00000;
      55533: inst = 32'h8c50000;
      55534: inst = 32'h24612800;
      55535: inst = 32'h10a0ffff;
      55536: inst = 32'hca0ffef;
      55537: inst = 32'h24822800;
      55538: inst = 32'h10a00000;
      55539: inst = 32'hca00004;
      55540: inst = 32'h38632800;
      55541: inst = 32'h38842800;
      55542: inst = 32'h10a00000;
      55543: inst = 32'hca0d8fb;
      55544: inst = 32'h13e00001;
      55545: inst = 32'hfe0d96a;
      55546: inst = 32'h5be00000;
      55547: inst = 32'h8c50000;
      55548: inst = 32'h24612800;
      55549: inst = 32'h10a0ffff;
      55550: inst = 32'hca0ffef;
      55551: inst = 32'h24822800;
      55552: inst = 32'h10a00000;
      55553: inst = 32'hca00004;
      55554: inst = 32'h38632800;
      55555: inst = 32'h38842800;
      55556: inst = 32'h10a00000;
      55557: inst = 32'hca0d909;
      55558: inst = 32'h13e00001;
      55559: inst = 32'hfe0d96a;
      55560: inst = 32'h5be00000;
      55561: inst = 32'h8c50000;
      55562: inst = 32'h24612800;
      55563: inst = 32'h10a0ffff;
      55564: inst = 32'hca0ffef;
      55565: inst = 32'h24822800;
      55566: inst = 32'h10a00000;
      55567: inst = 32'hca00004;
      55568: inst = 32'h38632800;
      55569: inst = 32'h38842800;
      55570: inst = 32'h10a00000;
      55571: inst = 32'hca0d917;
      55572: inst = 32'h13e00001;
      55573: inst = 32'hfe0d96a;
      55574: inst = 32'h5be00000;
      55575: inst = 32'h8c50000;
      55576: inst = 32'h24612800;
      55577: inst = 32'h10a0ffff;
      55578: inst = 32'hca0ffef;
      55579: inst = 32'h24822800;
      55580: inst = 32'h10a00000;
      55581: inst = 32'hca00004;
      55582: inst = 32'h38632800;
      55583: inst = 32'h38842800;
      55584: inst = 32'h10a00000;
      55585: inst = 32'hca0d925;
      55586: inst = 32'h13e00001;
      55587: inst = 32'hfe0d96a;
      55588: inst = 32'h5be00000;
      55589: inst = 32'h8c50000;
      55590: inst = 32'h24612800;
      55591: inst = 32'h10a0ffff;
      55592: inst = 32'hca0ffef;
      55593: inst = 32'h24822800;
      55594: inst = 32'h10a00000;
      55595: inst = 32'hca00004;
      55596: inst = 32'h38632800;
      55597: inst = 32'h38842800;
      55598: inst = 32'h10a00000;
      55599: inst = 32'hca0d933;
      55600: inst = 32'h13e00001;
      55601: inst = 32'hfe0d96a;
      55602: inst = 32'h5be00000;
      55603: inst = 32'h8c50000;
      55604: inst = 32'h24612800;
      55605: inst = 32'h10a0ffff;
      55606: inst = 32'hca0ffef;
      55607: inst = 32'h24822800;
      55608: inst = 32'h10a00000;
      55609: inst = 32'hca00004;
      55610: inst = 32'h38632800;
      55611: inst = 32'h38842800;
      55612: inst = 32'h10a00000;
      55613: inst = 32'hca0d941;
      55614: inst = 32'h13e00001;
      55615: inst = 32'hfe0d96a;
      55616: inst = 32'h5be00000;
      55617: inst = 32'h8c50000;
      55618: inst = 32'h24612800;
      55619: inst = 32'h10a0ffff;
      55620: inst = 32'hca0ffef;
      55621: inst = 32'h24822800;
      55622: inst = 32'h10a00000;
      55623: inst = 32'hca00004;
      55624: inst = 32'h38632800;
      55625: inst = 32'h38842800;
      55626: inst = 32'h10a00000;
      55627: inst = 32'hca0d94f;
      55628: inst = 32'h13e00001;
      55629: inst = 32'hfe0d96a;
      55630: inst = 32'h5be00000;
      55631: inst = 32'h8c50000;
      55632: inst = 32'h24612800;
      55633: inst = 32'h10a0ffff;
      55634: inst = 32'hca0ffef;
      55635: inst = 32'h24822800;
      55636: inst = 32'h10a00000;
      55637: inst = 32'hca00004;
      55638: inst = 32'h38632800;
      55639: inst = 32'h38842800;
      55640: inst = 32'h10a00000;
      55641: inst = 32'hca0d95d;
      55642: inst = 32'h13e00001;
      55643: inst = 32'hfe0d96a;
      55644: inst = 32'h5be00000;
      55645: inst = 32'h8c50000;
      55646: inst = 32'h24612800;
      55647: inst = 32'h10a0ffff;
      55648: inst = 32'hca0ffef;
      55649: inst = 32'h24822800;
      55650: inst = 32'h10a00000;
      55651: inst = 32'hca00004;
      55652: inst = 32'h38632800;
      55653: inst = 32'h38842800;
      55654: inst = 32'h10a00000;
      55655: inst = 32'hca0d96b;
      55656: inst = 32'h13e00001;
      55657: inst = 32'hfe0d96a;
      55658: inst = 32'h5be00000;
      55659: inst = 32'h8c50000;
      55660: inst = 32'h24612800;
      55661: inst = 32'h10a0ffff;
      55662: inst = 32'hca0ffef;
      55663: inst = 32'h24822800;
      55664: inst = 32'h10a00000;
      55665: inst = 32'hca00004;
      55666: inst = 32'h38632800;
      55667: inst = 32'h38842800;
      55668: inst = 32'h10a00000;
      55669: inst = 32'hca0d979;
      55670: inst = 32'h13e00001;
      55671: inst = 32'hfe0d96a;
      55672: inst = 32'h5be00000;
      55673: inst = 32'h8c50000;
      55674: inst = 32'h24612800;
      55675: inst = 32'h10a0ffff;
      55676: inst = 32'hca0ffef;
      55677: inst = 32'h24822800;
      55678: inst = 32'h10a00000;
      55679: inst = 32'hca00004;
      55680: inst = 32'h38632800;
      55681: inst = 32'h38842800;
      55682: inst = 32'h10a00000;
      55683: inst = 32'hca0d987;
      55684: inst = 32'h13e00001;
      55685: inst = 32'hfe0d96a;
      55686: inst = 32'h5be00000;
      55687: inst = 32'h8c50000;
      55688: inst = 32'h24612800;
      55689: inst = 32'h10a0ffff;
      55690: inst = 32'hca0ffef;
      55691: inst = 32'h24822800;
      55692: inst = 32'h10a00000;
      55693: inst = 32'hca00004;
      55694: inst = 32'h38632800;
      55695: inst = 32'h38842800;
      55696: inst = 32'h10a00000;
      55697: inst = 32'hca0d995;
      55698: inst = 32'h13e00001;
      55699: inst = 32'hfe0d96a;
      55700: inst = 32'h5be00000;
      55701: inst = 32'h8c50000;
      55702: inst = 32'h24612800;
      55703: inst = 32'h10a0ffff;
      55704: inst = 32'hca0ffef;
      55705: inst = 32'h24822800;
      55706: inst = 32'h10a00000;
      55707: inst = 32'hca00004;
      55708: inst = 32'h38632800;
      55709: inst = 32'h38842800;
      55710: inst = 32'h10a00000;
      55711: inst = 32'hca0d9a3;
      55712: inst = 32'h13e00001;
      55713: inst = 32'hfe0d96a;
      55714: inst = 32'h5be00000;
      55715: inst = 32'h8c50000;
      55716: inst = 32'h24612800;
      55717: inst = 32'h10a0ffff;
      55718: inst = 32'hca0ffef;
      55719: inst = 32'h24822800;
      55720: inst = 32'h10a00000;
      55721: inst = 32'hca00004;
      55722: inst = 32'h38632800;
      55723: inst = 32'h38842800;
      55724: inst = 32'h10a00000;
      55725: inst = 32'hca0d9b1;
      55726: inst = 32'h13e00001;
      55727: inst = 32'hfe0d96a;
      55728: inst = 32'h5be00000;
      55729: inst = 32'h8c50000;
      55730: inst = 32'h24612800;
      55731: inst = 32'h10a0ffff;
      55732: inst = 32'hca0ffef;
      55733: inst = 32'h24822800;
      55734: inst = 32'h10a00000;
      55735: inst = 32'hca00004;
      55736: inst = 32'h38632800;
      55737: inst = 32'h38842800;
      55738: inst = 32'h10a00000;
      55739: inst = 32'hca0d9bf;
      55740: inst = 32'h13e00001;
      55741: inst = 32'hfe0d96a;
      55742: inst = 32'h5be00000;
      55743: inst = 32'h8c50000;
      55744: inst = 32'h24612800;
      55745: inst = 32'h10a0ffff;
      55746: inst = 32'hca0ffef;
      55747: inst = 32'h24822800;
      55748: inst = 32'h10a00000;
      55749: inst = 32'hca00004;
      55750: inst = 32'h38632800;
      55751: inst = 32'h38842800;
      55752: inst = 32'h10a00000;
      55753: inst = 32'hca0d9cd;
      55754: inst = 32'h13e00001;
      55755: inst = 32'hfe0d96a;
      55756: inst = 32'h5be00000;
      55757: inst = 32'h8c50000;
      55758: inst = 32'h24612800;
      55759: inst = 32'h10a0ffff;
      55760: inst = 32'hca0ffef;
      55761: inst = 32'h24822800;
      55762: inst = 32'h10a00000;
      55763: inst = 32'hca00004;
      55764: inst = 32'h38632800;
      55765: inst = 32'h38842800;
      55766: inst = 32'h10a00000;
      55767: inst = 32'hca0d9db;
      55768: inst = 32'h13e00001;
      55769: inst = 32'hfe0d96a;
      55770: inst = 32'h5be00000;
      55771: inst = 32'h8c50000;
      55772: inst = 32'h24612800;
      55773: inst = 32'h10a0ffff;
      55774: inst = 32'hca0ffef;
      55775: inst = 32'h24822800;
      55776: inst = 32'h10a00000;
      55777: inst = 32'hca00004;
      55778: inst = 32'h38632800;
      55779: inst = 32'h38842800;
      55780: inst = 32'h10a00000;
      55781: inst = 32'hca0d9e9;
      55782: inst = 32'h13e00001;
      55783: inst = 32'hfe0d96a;
      55784: inst = 32'h5be00000;
      55785: inst = 32'h8c50000;
      55786: inst = 32'h24612800;
      55787: inst = 32'h10a0ffff;
      55788: inst = 32'hca0ffef;
      55789: inst = 32'h24822800;
      55790: inst = 32'h10a00000;
      55791: inst = 32'hca00004;
      55792: inst = 32'h38632800;
      55793: inst = 32'h38842800;
      55794: inst = 32'h10a00000;
      55795: inst = 32'hca0d9f7;
      55796: inst = 32'h13e00001;
      55797: inst = 32'hfe0d96a;
      55798: inst = 32'h5be00000;
      55799: inst = 32'h8c50000;
      55800: inst = 32'h24612800;
      55801: inst = 32'h10a0ffff;
      55802: inst = 32'hca0ffef;
      55803: inst = 32'h24822800;
      55804: inst = 32'h10a00000;
      55805: inst = 32'hca00004;
      55806: inst = 32'h38632800;
      55807: inst = 32'h38842800;
      55808: inst = 32'h10a00000;
      55809: inst = 32'hca0da05;
      55810: inst = 32'h13e00001;
      55811: inst = 32'hfe0d96a;
      55812: inst = 32'h5be00000;
      55813: inst = 32'h8c50000;
      55814: inst = 32'h24612800;
      55815: inst = 32'h10a0ffff;
      55816: inst = 32'hca0ffef;
      55817: inst = 32'h24822800;
      55818: inst = 32'h10a00000;
      55819: inst = 32'hca00004;
      55820: inst = 32'h38632800;
      55821: inst = 32'h38842800;
      55822: inst = 32'h10a00000;
      55823: inst = 32'hca0da13;
      55824: inst = 32'h13e00001;
      55825: inst = 32'hfe0d96a;
      55826: inst = 32'h5be00000;
      55827: inst = 32'h8c50000;
      55828: inst = 32'h24612800;
      55829: inst = 32'h10a0ffff;
      55830: inst = 32'hca0ffef;
      55831: inst = 32'h24822800;
      55832: inst = 32'h10a00000;
      55833: inst = 32'hca00004;
      55834: inst = 32'h38632800;
      55835: inst = 32'h38842800;
      55836: inst = 32'h10a00000;
      55837: inst = 32'hca0da21;
      55838: inst = 32'h13e00001;
      55839: inst = 32'hfe0d96a;
      55840: inst = 32'h5be00000;
      55841: inst = 32'h8c50000;
      55842: inst = 32'h24612800;
      55843: inst = 32'h10a0ffff;
      55844: inst = 32'hca0ffef;
      55845: inst = 32'h24822800;
      55846: inst = 32'h10a00000;
      55847: inst = 32'hca00004;
      55848: inst = 32'h38632800;
      55849: inst = 32'h38842800;
      55850: inst = 32'h10a00000;
      55851: inst = 32'hca0da2f;
      55852: inst = 32'h13e00001;
      55853: inst = 32'hfe0d96a;
      55854: inst = 32'h5be00000;
      55855: inst = 32'h8c50000;
      55856: inst = 32'h24612800;
      55857: inst = 32'h10a0ffff;
      55858: inst = 32'hca0ffef;
      55859: inst = 32'h24822800;
      55860: inst = 32'h10a00000;
      55861: inst = 32'hca00004;
      55862: inst = 32'h38632800;
      55863: inst = 32'h38842800;
      55864: inst = 32'h10a00000;
      55865: inst = 32'hca0da3d;
      55866: inst = 32'h13e00001;
      55867: inst = 32'hfe0d96a;
      55868: inst = 32'h5be00000;
      55869: inst = 32'h8c50000;
      55870: inst = 32'h24612800;
      55871: inst = 32'h10a0ffff;
      55872: inst = 32'hca0ffef;
      55873: inst = 32'h24822800;
      55874: inst = 32'h10a00000;
      55875: inst = 32'hca00004;
      55876: inst = 32'h38632800;
      55877: inst = 32'h38842800;
      55878: inst = 32'h10a00000;
      55879: inst = 32'hca0da4b;
      55880: inst = 32'h13e00001;
      55881: inst = 32'hfe0d96a;
      55882: inst = 32'h5be00000;
      55883: inst = 32'h8c50000;
      55884: inst = 32'h24612800;
      55885: inst = 32'h10a0ffff;
      55886: inst = 32'hca0ffef;
      55887: inst = 32'h24822800;
      55888: inst = 32'h10a00000;
      55889: inst = 32'hca00004;
      55890: inst = 32'h38632800;
      55891: inst = 32'h38842800;
      55892: inst = 32'h10a00000;
      55893: inst = 32'hca0da59;
      55894: inst = 32'h13e00001;
      55895: inst = 32'hfe0d96a;
      55896: inst = 32'h5be00000;
      55897: inst = 32'h8c50000;
      55898: inst = 32'h24612800;
      55899: inst = 32'h10a0ffff;
      55900: inst = 32'hca0ffef;
      55901: inst = 32'h24822800;
      55902: inst = 32'h10a00000;
      55903: inst = 32'hca00004;
      55904: inst = 32'h38632800;
      55905: inst = 32'h38842800;
      55906: inst = 32'h10a00000;
      55907: inst = 32'hca0da67;
      55908: inst = 32'h13e00001;
      55909: inst = 32'hfe0d96a;
      55910: inst = 32'h5be00000;
      55911: inst = 32'h8c50000;
      55912: inst = 32'h24612800;
      55913: inst = 32'h10a0ffff;
      55914: inst = 32'hca0ffef;
      55915: inst = 32'h24822800;
      55916: inst = 32'h10a00000;
      55917: inst = 32'hca00004;
      55918: inst = 32'h38632800;
      55919: inst = 32'h38842800;
      55920: inst = 32'h10a00000;
      55921: inst = 32'hca0da75;
      55922: inst = 32'h13e00001;
      55923: inst = 32'hfe0d96a;
      55924: inst = 32'h5be00000;
      55925: inst = 32'h8c50000;
      55926: inst = 32'h24612800;
      55927: inst = 32'h10a0ffff;
      55928: inst = 32'hca0ffef;
      55929: inst = 32'h24822800;
      55930: inst = 32'h10a00000;
      55931: inst = 32'hca00004;
      55932: inst = 32'h38632800;
      55933: inst = 32'h38842800;
      55934: inst = 32'h10a00000;
      55935: inst = 32'hca0da83;
      55936: inst = 32'h13e00001;
      55937: inst = 32'hfe0d96a;
      55938: inst = 32'h5be00000;
      55939: inst = 32'h8c50000;
      55940: inst = 32'h24612800;
      55941: inst = 32'h10a0ffff;
      55942: inst = 32'hca0ffef;
      55943: inst = 32'h24822800;
      55944: inst = 32'h10a00000;
      55945: inst = 32'hca00004;
      55946: inst = 32'h38632800;
      55947: inst = 32'h38842800;
      55948: inst = 32'h10a00000;
      55949: inst = 32'hca0da91;
      55950: inst = 32'h13e00001;
      55951: inst = 32'hfe0d96a;
      55952: inst = 32'h5be00000;
      55953: inst = 32'h8c50000;
      55954: inst = 32'h24612800;
      55955: inst = 32'h10a0ffff;
      55956: inst = 32'hca0ffef;
      55957: inst = 32'h24822800;
      55958: inst = 32'h10a00000;
      55959: inst = 32'hca00004;
      55960: inst = 32'h38632800;
      55961: inst = 32'h38842800;
      55962: inst = 32'h10a00000;
      55963: inst = 32'hca0da9f;
      55964: inst = 32'h13e00001;
      55965: inst = 32'hfe0d96a;
      55966: inst = 32'h5be00000;
      55967: inst = 32'h8c50000;
      55968: inst = 32'h24612800;
      55969: inst = 32'h10a0ffff;
      55970: inst = 32'hca0ffef;
      55971: inst = 32'h24822800;
      55972: inst = 32'h10a00000;
      55973: inst = 32'hca00004;
      55974: inst = 32'h38632800;
      55975: inst = 32'h38842800;
      55976: inst = 32'h10a00000;
      55977: inst = 32'hca0daad;
      55978: inst = 32'h13e00001;
      55979: inst = 32'hfe0d96a;
      55980: inst = 32'h5be00000;
      55981: inst = 32'h8c50000;
      55982: inst = 32'h24612800;
      55983: inst = 32'h10a0ffff;
      55984: inst = 32'hca0ffef;
      55985: inst = 32'h24822800;
      55986: inst = 32'h10a00000;
      55987: inst = 32'hca00004;
      55988: inst = 32'h38632800;
      55989: inst = 32'h38842800;
      55990: inst = 32'h10a00000;
      55991: inst = 32'hca0dabb;
      55992: inst = 32'h13e00001;
      55993: inst = 32'hfe0d96a;
      55994: inst = 32'h5be00000;
      55995: inst = 32'h8c50000;
      55996: inst = 32'h24612800;
      55997: inst = 32'h10a0ffff;
      55998: inst = 32'hca0ffef;
      55999: inst = 32'h24822800;
      56000: inst = 32'h10a00000;
      56001: inst = 32'hca00004;
      56002: inst = 32'h38632800;
      56003: inst = 32'h38842800;
      56004: inst = 32'h10a00000;
      56005: inst = 32'hca0dac9;
      56006: inst = 32'h13e00001;
      56007: inst = 32'hfe0d96a;
      56008: inst = 32'h5be00000;
      56009: inst = 32'h8c50000;
      56010: inst = 32'h24612800;
      56011: inst = 32'h10a0ffff;
      56012: inst = 32'hca0ffef;
      56013: inst = 32'h24822800;
      56014: inst = 32'h10a00000;
      56015: inst = 32'hca00004;
      56016: inst = 32'h38632800;
      56017: inst = 32'h38842800;
      56018: inst = 32'h10a00000;
      56019: inst = 32'hca0dad7;
      56020: inst = 32'h13e00001;
      56021: inst = 32'hfe0d96a;
      56022: inst = 32'h5be00000;
      56023: inst = 32'h8c50000;
      56024: inst = 32'h24612800;
      56025: inst = 32'h10a0ffff;
      56026: inst = 32'hca0ffef;
      56027: inst = 32'h24822800;
      56028: inst = 32'h10a00000;
      56029: inst = 32'hca00004;
      56030: inst = 32'h38632800;
      56031: inst = 32'h38842800;
      56032: inst = 32'h10a00000;
      56033: inst = 32'hca0dae5;
      56034: inst = 32'h13e00001;
      56035: inst = 32'hfe0d96a;
      56036: inst = 32'h5be00000;
      56037: inst = 32'h8c50000;
      56038: inst = 32'h24612800;
      56039: inst = 32'h10a0ffff;
      56040: inst = 32'hca0ffef;
      56041: inst = 32'h24822800;
      56042: inst = 32'h10a00000;
      56043: inst = 32'hca00004;
      56044: inst = 32'h38632800;
      56045: inst = 32'h38842800;
      56046: inst = 32'h10a00000;
      56047: inst = 32'hca0daf3;
      56048: inst = 32'h13e00001;
      56049: inst = 32'hfe0d96a;
      56050: inst = 32'h5be00000;
      56051: inst = 32'h8c50000;
      56052: inst = 32'h24612800;
      56053: inst = 32'h10a0ffff;
      56054: inst = 32'hca0ffef;
      56055: inst = 32'h24822800;
      56056: inst = 32'h10a00000;
      56057: inst = 32'hca00004;
      56058: inst = 32'h38632800;
      56059: inst = 32'h38842800;
      56060: inst = 32'h10a00000;
      56061: inst = 32'hca0db01;
      56062: inst = 32'h13e00001;
      56063: inst = 32'hfe0d96a;
      56064: inst = 32'h5be00000;
      56065: inst = 32'h8c50000;
      56066: inst = 32'h24612800;
      56067: inst = 32'h10a0ffff;
      56068: inst = 32'hca0ffef;
      56069: inst = 32'h24822800;
      56070: inst = 32'h10a00000;
      56071: inst = 32'hca00004;
      56072: inst = 32'h38632800;
      56073: inst = 32'h38842800;
      56074: inst = 32'h10a00000;
      56075: inst = 32'hca0db0f;
      56076: inst = 32'h13e00001;
      56077: inst = 32'hfe0d96a;
      56078: inst = 32'h5be00000;
      56079: inst = 32'h8c50000;
      56080: inst = 32'h24612800;
      56081: inst = 32'h10a0ffff;
      56082: inst = 32'hca0ffef;
      56083: inst = 32'h24822800;
      56084: inst = 32'h10a00000;
      56085: inst = 32'hca00004;
      56086: inst = 32'h38632800;
      56087: inst = 32'h38842800;
      56088: inst = 32'h10a00000;
      56089: inst = 32'hca0db1d;
      56090: inst = 32'h13e00001;
      56091: inst = 32'hfe0d96a;
      56092: inst = 32'h5be00000;
      56093: inst = 32'h8c50000;
      56094: inst = 32'h24612800;
      56095: inst = 32'h10a0ffff;
      56096: inst = 32'hca0ffef;
      56097: inst = 32'h24822800;
      56098: inst = 32'h10a00000;
      56099: inst = 32'hca00004;
      56100: inst = 32'h38632800;
      56101: inst = 32'h38842800;
      56102: inst = 32'h10a00000;
      56103: inst = 32'hca0db2b;
      56104: inst = 32'h13e00001;
      56105: inst = 32'hfe0d96a;
      56106: inst = 32'h5be00000;
      56107: inst = 32'h8c50000;
      56108: inst = 32'h24612800;
      56109: inst = 32'h10a0ffff;
      56110: inst = 32'hca0ffef;
      56111: inst = 32'h24822800;
      56112: inst = 32'h10a00000;
      56113: inst = 32'hca00004;
      56114: inst = 32'h38632800;
      56115: inst = 32'h38842800;
      56116: inst = 32'h10a00000;
      56117: inst = 32'hca0db39;
      56118: inst = 32'h13e00001;
      56119: inst = 32'hfe0d96a;
      56120: inst = 32'h5be00000;
      56121: inst = 32'h8c50000;
      56122: inst = 32'h24612800;
      56123: inst = 32'h10a0ffff;
      56124: inst = 32'hca0ffef;
      56125: inst = 32'h24822800;
      56126: inst = 32'h10a00000;
      56127: inst = 32'hca00004;
      56128: inst = 32'h38632800;
      56129: inst = 32'h38842800;
      56130: inst = 32'h10a00000;
      56131: inst = 32'hca0db47;
      56132: inst = 32'h13e00001;
      56133: inst = 32'hfe0d96a;
      56134: inst = 32'h5be00000;
      56135: inst = 32'h8c50000;
      56136: inst = 32'h24612800;
      56137: inst = 32'h10a0ffff;
      56138: inst = 32'hca0ffef;
      56139: inst = 32'h24822800;
      56140: inst = 32'h10a00000;
      56141: inst = 32'hca00004;
      56142: inst = 32'h38632800;
      56143: inst = 32'h38842800;
      56144: inst = 32'h10a00000;
      56145: inst = 32'hca0db55;
      56146: inst = 32'h13e00001;
      56147: inst = 32'hfe0d96a;
      56148: inst = 32'h5be00000;
      56149: inst = 32'h8c50000;
      56150: inst = 32'h24612800;
      56151: inst = 32'h10a0ffff;
      56152: inst = 32'hca0ffef;
      56153: inst = 32'h24822800;
      56154: inst = 32'h10a00000;
      56155: inst = 32'hca00004;
      56156: inst = 32'h38632800;
      56157: inst = 32'h38842800;
      56158: inst = 32'h10a00000;
      56159: inst = 32'hca0db63;
      56160: inst = 32'h13e00001;
      56161: inst = 32'hfe0d96a;
      56162: inst = 32'h5be00000;
      56163: inst = 32'h8c50000;
      56164: inst = 32'h24612800;
      56165: inst = 32'h10a0ffff;
      56166: inst = 32'hca0ffef;
      56167: inst = 32'h24822800;
      56168: inst = 32'h10a00000;
      56169: inst = 32'hca00004;
      56170: inst = 32'h38632800;
      56171: inst = 32'h38842800;
      56172: inst = 32'h10a00000;
      56173: inst = 32'hca0db71;
      56174: inst = 32'h13e00001;
      56175: inst = 32'hfe0d96a;
      56176: inst = 32'h5be00000;
      56177: inst = 32'h8c50000;
      56178: inst = 32'h24612800;
      56179: inst = 32'h10a0ffff;
      56180: inst = 32'hca0ffef;
      56181: inst = 32'h24822800;
      56182: inst = 32'h10a00000;
      56183: inst = 32'hca00004;
      56184: inst = 32'h38632800;
      56185: inst = 32'h38842800;
      56186: inst = 32'h10a00000;
      56187: inst = 32'hca0db7f;
      56188: inst = 32'h13e00001;
      56189: inst = 32'hfe0d96a;
      56190: inst = 32'h5be00000;
      56191: inst = 32'h8c50000;
      56192: inst = 32'h24612800;
      56193: inst = 32'h10a0ffff;
      56194: inst = 32'hca0ffef;
      56195: inst = 32'h24822800;
      56196: inst = 32'h10a00000;
      56197: inst = 32'hca00004;
      56198: inst = 32'h38632800;
      56199: inst = 32'h38842800;
      56200: inst = 32'h10a00000;
      56201: inst = 32'hca0db8d;
      56202: inst = 32'h13e00001;
      56203: inst = 32'hfe0d96a;
      56204: inst = 32'h5be00000;
      56205: inst = 32'h8c50000;
      56206: inst = 32'h24612800;
      56207: inst = 32'h10a0ffff;
      56208: inst = 32'hca0ffef;
      56209: inst = 32'h24822800;
      56210: inst = 32'h10a00000;
      56211: inst = 32'hca00004;
      56212: inst = 32'h38632800;
      56213: inst = 32'h38842800;
      56214: inst = 32'h10a00000;
      56215: inst = 32'hca0db9b;
      56216: inst = 32'h13e00001;
      56217: inst = 32'hfe0d96a;
      56218: inst = 32'h5be00000;
      56219: inst = 32'h8c50000;
      56220: inst = 32'h24612800;
      56221: inst = 32'h10a0ffff;
      56222: inst = 32'hca0ffef;
      56223: inst = 32'h24822800;
      56224: inst = 32'h10a00000;
      56225: inst = 32'hca00004;
      56226: inst = 32'h38632800;
      56227: inst = 32'h38842800;
      56228: inst = 32'h10a00000;
      56229: inst = 32'hca0dba9;
      56230: inst = 32'h13e00001;
      56231: inst = 32'hfe0d96a;
      56232: inst = 32'h5be00000;
      56233: inst = 32'h8c50000;
      56234: inst = 32'h24612800;
      56235: inst = 32'h10a0ffff;
      56236: inst = 32'hca0ffef;
      56237: inst = 32'h24822800;
      56238: inst = 32'h10a00000;
      56239: inst = 32'hca00004;
      56240: inst = 32'h38632800;
      56241: inst = 32'h38842800;
      56242: inst = 32'h10a00000;
      56243: inst = 32'hca0dbb7;
      56244: inst = 32'h13e00001;
      56245: inst = 32'hfe0d96a;
      56246: inst = 32'h5be00000;
      56247: inst = 32'h8c50000;
      56248: inst = 32'h24612800;
      56249: inst = 32'h10a0ffff;
      56250: inst = 32'hca0ffef;
      56251: inst = 32'h24822800;
      56252: inst = 32'h10a00000;
      56253: inst = 32'hca00004;
      56254: inst = 32'h38632800;
      56255: inst = 32'h38842800;
      56256: inst = 32'h10a00000;
      56257: inst = 32'hca0dbc5;
      56258: inst = 32'h13e00001;
      56259: inst = 32'hfe0d96a;
      56260: inst = 32'h5be00000;
      56261: inst = 32'h8c50000;
      56262: inst = 32'h24612800;
      56263: inst = 32'h10a0ffff;
      56264: inst = 32'hca0ffef;
      56265: inst = 32'h24822800;
      56266: inst = 32'h10a00000;
      56267: inst = 32'hca00004;
      56268: inst = 32'h38632800;
      56269: inst = 32'h38842800;
      56270: inst = 32'h10a00000;
      56271: inst = 32'hca0dbd3;
      56272: inst = 32'h13e00001;
      56273: inst = 32'hfe0d96a;
      56274: inst = 32'h5be00000;
      56275: inst = 32'h8c50000;
      56276: inst = 32'h24612800;
      56277: inst = 32'h10a0ffff;
      56278: inst = 32'hca0ffef;
      56279: inst = 32'h24822800;
      56280: inst = 32'h10a00000;
      56281: inst = 32'hca00004;
      56282: inst = 32'h38632800;
      56283: inst = 32'h38842800;
      56284: inst = 32'h10a00000;
      56285: inst = 32'hca0dbe1;
      56286: inst = 32'h13e00001;
      56287: inst = 32'hfe0d96a;
      56288: inst = 32'h5be00000;
      56289: inst = 32'h8c50000;
      56290: inst = 32'h24612800;
      56291: inst = 32'h10a0ffff;
      56292: inst = 32'hca0ffef;
      56293: inst = 32'h24822800;
      56294: inst = 32'h10a00000;
      56295: inst = 32'hca00004;
      56296: inst = 32'h38632800;
      56297: inst = 32'h38842800;
      56298: inst = 32'h10a00000;
      56299: inst = 32'hca0dbef;
      56300: inst = 32'h13e00001;
      56301: inst = 32'hfe0d96a;
      56302: inst = 32'h5be00000;
      56303: inst = 32'h8c50000;
      56304: inst = 32'h24612800;
      56305: inst = 32'h10a0ffff;
      56306: inst = 32'hca0ffef;
      56307: inst = 32'h24822800;
      56308: inst = 32'h10a00000;
      56309: inst = 32'hca00004;
      56310: inst = 32'h38632800;
      56311: inst = 32'h38842800;
      56312: inst = 32'h10a00000;
      56313: inst = 32'hca0dbfd;
      56314: inst = 32'h13e00001;
      56315: inst = 32'hfe0d96a;
      56316: inst = 32'h5be00000;
      56317: inst = 32'h8c50000;
      56318: inst = 32'h24612800;
      56319: inst = 32'h10a0ffff;
      56320: inst = 32'hca0ffef;
      56321: inst = 32'h24822800;
      56322: inst = 32'h10a00000;
      56323: inst = 32'hca00004;
      56324: inst = 32'h38632800;
      56325: inst = 32'h38842800;
      56326: inst = 32'h10a00000;
      56327: inst = 32'hca0dc0b;
      56328: inst = 32'h13e00001;
      56329: inst = 32'hfe0d96a;
      56330: inst = 32'h5be00000;
      56331: inst = 32'h8c50000;
      56332: inst = 32'h24612800;
      56333: inst = 32'h10a0ffff;
      56334: inst = 32'hca0ffef;
      56335: inst = 32'h24822800;
      56336: inst = 32'h10a00000;
      56337: inst = 32'hca00004;
      56338: inst = 32'h38632800;
      56339: inst = 32'h38842800;
      56340: inst = 32'h10a00000;
      56341: inst = 32'hca0dc19;
      56342: inst = 32'h13e00001;
      56343: inst = 32'hfe0d96a;
      56344: inst = 32'h5be00000;
      56345: inst = 32'h8c50000;
      56346: inst = 32'h24612800;
      56347: inst = 32'h10a0ffff;
      56348: inst = 32'hca0ffef;
      56349: inst = 32'h24822800;
      56350: inst = 32'h10a00000;
      56351: inst = 32'hca00004;
      56352: inst = 32'h38632800;
      56353: inst = 32'h38842800;
      56354: inst = 32'h10a00000;
      56355: inst = 32'hca0dc27;
      56356: inst = 32'h13e00001;
      56357: inst = 32'hfe0d96a;
      56358: inst = 32'h5be00000;
      56359: inst = 32'h8c50000;
      56360: inst = 32'h24612800;
      56361: inst = 32'h10a0ffff;
      56362: inst = 32'hca0ffef;
      56363: inst = 32'h24822800;
      56364: inst = 32'h10a00000;
      56365: inst = 32'hca00004;
      56366: inst = 32'h38632800;
      56367: inst = 32'h38842800;
      56368: inst = 32'h10a00000;
      56369: inst = 32'hca0dc35;
      56370: inst = 32'h13e00001;
      56371: inst = 32'hfe0d96a;
      56372: inst = 32'h5be00000;
      56373: inst = 32'h8c50000;
      56374: inst = 32'h24612800;
      56375: inst = 32'h10a0ffff;
      56376: inst = 32'hca0ffef;
      56377: inst = 32'h24822800;
      56378: inst = 32'h10a00000;
      56379: inst = 32'hca00004;
      56380: inst = 32'h38632800;
      56381: inst = 32'h38842800;
      56382: inst = 32'h10a00000;
      56383: inst = 32'hca0dc43;
      56384: inst = 32'h13e00001;
      56385: inst = 32'hfe0d96a;
      56386: inst = 32'h5be00000;
      56387: inst = 32'h8c50000;
      56388: inst = 32'h24612800;
      56389: inst = 32'h10a0ffff;
      56390: inst = 32'hca0ffef;
      56391: inst = 32'h24822800;
      56392: inst = 32'h10a00000;
      56393: inst = 32'hca00004;
      56394: inst = 32'h38632800;
      56395: inst = 32'h38842800;
      56396: inst = 32'h10a00000;
      56397: inst = 32'hca0dc51;
      56398: inst = 32'h13e00001;
      56399: inst = 32'hfe0d96a;
      56400: inst = 32'h5be00000;
      56401: inst = 32'h8c50000;
      56402: inst = 32'h24612800;
      56403: inst = 32'h10a0ffff;
      56404: inst = 32'hca0ffef;
      56405: inst = 32'h24822800;
      56406: inst = 32'h10a00000;
      56407: inst = 32'hca00004;
      56408: inst = 32'h38632800;
      56409: inst = 32'h38842800;
      56410: inst = 32'h10a00000;
      56411: inst = 32'hca0dc5f;
      56412: inst = 32'h13e00001;
      56413: inst = 32'hfe0d96a;
      56414: inst = 32'h5be00000;
      56415: inst = 32'h8c50000;
      56416: inst = 32'h24612800;
      56417: inst = 32'h10a0ffff;
      56418: inst = 32'hca0ffef;
      56419: inst = 32'h24822800;
      56420: inst = 32'h10a00000;
      56421: inst = 32'hca00004;
      56422: inst = 32'h38632800;
      56423: inst = 32'h38842800;
      56424: inst = 32'h10a00000;
      56425: inst = 32'hca0dc6d;
      56426: inst = 32'h13e00001;
      56427: inst = 32'hfe0d96a;
      56428: inst = 32'h5be00000;
      56429: inst = 32'h8c50000;
      56430: inst = 32'h24612800;
      56431: inst = 32'h10a0ffff;
      56432: inst = 32'hca0ffef;
      56433: inst = 32'h24822800;
      56434: inst = 32'h10a00000;
      56435: inst = 32'hca00004;
      56436: inst = 32'h38632800;
      56437: inst = 32'h38842800;
      56438: inst = 32'h10a00000;
      56439: inst = 32'hca0dc7b;
      56440: inst = 32'h13e00001;
      56441: inst = 32'hfe0d96a;
      56442: inst = 32'h5be00000;
      56443: inst = 32'h8c50000;
      56444: inst = 32'h24612800;
      56445: inst = 32'h10a0ffff;
      56446: inst = 32'hca0ffef;
      56447: inst = 32'h24822800;
      56448: inst = 32'h10a00000;
      56449: inst = 32'hca00004;
      56450: inst = 32'h38632800;
      56451: inst = 32'h38842800;
      56452: inst = 32'h10a00000;
      56453: inst = 32'hca0dc89;
      56454: inst = 32'h13e00001;
      56455: inst = 32'hfe0d96a;
      56456: inst = 32'h5be00000;
      56457: inst = 32'h8c50000;
      56458: inst = 32'h24612800;
      56459: inst = 32'h10a0ffff;
      56460: inst = 32'hca0ffef;
      56461: inst = 32'h24822800;
      56462: inst = 32'h10a00000;
      56463: inst = 32'hca00004;
      56464: inst = 32'h38632800;
      56465: inst = 32'h38842800;
      56466: inst = 32'h10a00000;
      56467: inst = 32'hca0dc97;
      56468: inst = 32'h13e00001;
      56469: inst = 32'hfe0d96a;
      56470: inst = 32'h5be00000;
      56471: inst = 32'h8c50000;
      56472: inst = 32'h24612800;
      56473: inst = 32'h10a0ffff;
      56474: inst = 32'hca0ffef;
      56475: inst = 32'h24822800;
      56476: inst = 32'h10a00000;
      56477: inst = 32'hca00004;
      56478: inst = 32'h38632800;
      56479: inst = 32'h38842800;
      56480: inst = 32'h10a00000;
      56481: inst = 32'hca0dca5;
      56482: inst = 32'h13e00001;
      56483: inst = 32'hfe0d96a;
      56484: inst = 32'h5be00000;
      56485: inst = 32'h8c50000;
      56486: inst = 32'h24612800;
      56487: inst = 32'h10a0ffff;
      56488: inst = 32'hca0ffef;
      56489: inst = 32'h24822800;
      56490: inst = 32'h10a00000;
      56491: inst = 32'hca00004;
      56492: inst = 32'h38632800;
      56493: inst = 32'h38842800;
      56494: inst = 32'h10a00000;
      56495: inst = 32'hca0dcb3;
      56496: inst = 32'h13e00001;
      56497: inst = 32'hfe0d96a;
      56498: inst = 32'h5be00000;
      56499: inst = 32'h8c50000;
      56500: inst = 32'h24612800;
      56501: inst = 32'h10a0ffff;
      56502: inst = 32'hca0ffef;
      56503: inst = 32'h24822800;
      56504: inst = 32'h10a00000;
      56505: inst = 32'hca00004;
      56506: inst = 32'h38632800;
      56507: inst = 32'h38842800;
      56508: inst = 32'h10a00000;
      56509: inst = 32'hca0dcc1;
      56510: inst = 32'h13e00001;
      56511: inst = 32'hfe0d96a;
      56512: inst = 32'h5be00000;
      56513: inst = 32'h8c50000;
      56514: inst = 32'h24612800;
      56515: inst = 32'h10a0ffff;
      56516: inst = 32'hca0ffef;
      56517: inst = 32'h24822800;
      56518: inst = 32'h10a00000;
      56519: inst = 32'hca00004;
      56520: inst = 32'h38632800;
      56521: inst = 32'h38842800;
      56522: inst = 32'h10a00000;
      56523: inst = 32'hca0dccf;
      56524: inst = 32'h13e00001;
      56525: inst = 32'hfe0d96a;
      56526: inst = 32'h5be00000;
      56527: inst = 32'h8c50000;
      56528: inst = 32'h24612800;
      56529: inst = 32'h10a0ffff;
      56530: inst = 32'hca0ffef;
      56531: inst = 32'h24822800;
      56532: inst = 32'h10a00000;
      56533: inst = 32'hca00004;
      56534: inst = 32'h38632800;
      56535: inst = 32'h38842800;
      56536: inst = 32'h10a00000;
      56537: inst = 32'hca0dcdd;
      56538: inst = 32'h13e00001;
      56539: inst = 32'hfe0d96a;
      56540: inst = 32'h5be00000;
      56541: inst = 32'h8c50000;
      56542: inst = 32'h24612800;
      56543: inst = 32'h10a0ffff;
      56544: inst = 32'hca0ffef;
      56545: inst = 32'h24822800;
      56546: inst = 32'h10a00000;
      56547: inst = 32'hca00004;
      56548: inst = 32'h38632800;
      56549: inst = 32'h38842800;
      56550: inst = 32'h10a00000;
      56551: inst = 32'hca0dceb;
      56552: inst = 32'h13e00001;
      56553: inst = 32'hfe0d96a;
      56554: inst = 32'h5be00000;
      56555: inst = 32'h8c50000;
      56556: inst = 32'h24612800;
      56557: inst = 32'h10a0ffff;
      56558: inst = 32'hca0ffef;
      56559: inst = 32'h24822800;
      56560: inst = 32'h10a00000;
      56561: inst = 32'hca00004;
      56562: inst = 32'h38632800;
      56563: inst = 32'h38842800;
      56564: inst = 32'h10a00000;
      56565: inst = 32'hca0dcf9;
      56566: inst = 32'h13e00001;
      56567: inst = 32'hfe0d96a;
      56568: inst = 32'h5be00000;
      56569: inst = 32'h8c50000;
      56570: inst = 32'h24612800;
      56571: inst = 32'h10a0ffff;
      56572: inst = 32'hca0ffef;
      56573: inst = 32'h24822800;
      56574: inst = 32'h10a00000;
      56575: inst = 32'hca00004;
      56576: inst = 32'h38632800;
      56577: inst = 32'h38842800;
      56578: inst = 32'h10a00000;
      56579: inst = 32'hca0dd07;
      56580: inst = 32'h13e00001;
      56581: inst = 32'hfe0d96a;
      56582: inst = 32'h5be00000;
      56583: inst = 32'h8c50000;
      56584: inst = 32'h24612800;
      56585: inst = 32'h10a0ffff;
      56586: inst = 32'hca0ffef;
      56587: inst = 32'h24822800;
      56588: inst = 32'h10a00000;
      56589: inst = 32'hca00004;
      56590: inst = 32'h38632800;
      56591: inst = 32'h38842800;
      56592: inst = 32'h10a00000;
      56593: inst = 32'hca0dd15;
      56594: inst = 32'h13e00001;
      56595: inst = 32'hfe0d96a;
      56596: inst = 32'h5be00000;
      56597: inst = 32'h8c50000;
      56598: inst = 32'h24612800;
      56599: inst = 32'h10a0ffff;
      56600: inst = 32'hca0ffef;
      56601: inst = 32'h24822800;
      56602: inst = 32'h10a00000;
      56603: inst = 32'hca00004;
      56604: inst = 32'h38632800;
      56605: inst = 32'h38842800;
      56606: inst = 32'h10a00000;
      56607: inst = 32'hca0dd23;
      56608: inst = 32'h13e00001;
      56609: inst = 32'hfe0d96a;
      56610: inst = 32'h5be00000;
      56611: inst = 32'h8c50000;
      56612: inst = 32'h24612800;
      56613: inst = 32'h10a0ffff;
      56614: inst = 32'hca0ffef;
      56615: inst = 32'h24822800;
      56616: inst = 32'h10a00000;
      56617: inst = 32'hca00004;
      56618: inst = 32'h38632800;
      56619: inst = 32'h38842800;
      56620: inst = 32'h10a00000;
      56621: inst = 32'hca0dd31;
      56622: inst = 32'h13e00001;
      56623: inst = 32'hfe0d96a;
      56624: inst = 32'h5be00000;
      56625: inst = 32'h8c50000;
      56626: inst = 32'h24612800;
      56627: inst = 32'h10a0ffff;
      56628: inst = 32'hca0ffef;
      56629: inst = 32'h24822800;
      56630: inst = 32'h10a00000;
      56631: inst = 32'hca00004;
      56632: inst = 32'h38632800;
      56633: inst = 32'h38842800;
      56634: inst = 32'h10a00000;
      56635: inst = 32'hca0dd3f;
      56636: inst = 32'h13e00001;
      56637: inst = 32'hfe0d96a;
      56638: inst = 32'h5be00000;
      56639: inst = 32'h8c50000;
      56640: inst = 32'h24612800;
      56641: inst = 32'h10a0ffff;
      56642: inst = 32'hca0ffef;
      56643: inst = 32'h24822800;
      56644: inst = 32'h10a00000;
      56645: inst = 32'hca00004;
      56646: inst = 32'h38632800;
      56647: inst = 32'h38842800;
      56648: inst = 32'h10a00000;
      56649: inst = 32'hca0dd4d;
      56650: inst = 32'h13e00001;
      56651: inst = 32'hfe0d96a;
      56652: inst = 32'h5be00000;
      56653: inst = 32'h8c50000;
      56654: inst = 32'h24612800;
      56655: inst = 32'h10a0ffff;
      56656: inst = 32'hca0ffef;
      56657: inst = 32'h24822800;
      56658: inst = 32'h10a00000;
      56659: inst = 32'hca00004;
      56660: inst = 32'h38632800;
      56661: inst = 32'h38842800;
      56662: inst = 32'h10a00000;
      56663: inst = 32'hca0dd5b;
      56664: inst = 32'h13e00001;
      56665: inst = 32'hfe0d96a;
      56666: inst = 32'h5be00000;
      56667: inst = 32'h8c50000;
      56668: inst = 32'h24612800;
      56669: inst = 32'h10a0ffff;
      56670: inst = 32'hca0ffef;
      56671: inst = 32'h24822800;
      56672: inst = 32'h10a00000;
      56673: inst = 32'hca00004;
      56674: inst = 32'h38632800;
      56675: inst = 32'h38842800;
      56676: inst = 32'h10a00000;
      56677: inst = 32'hca0dd69;
      56678: inst = 32'h13e00001;
      56679: inst = 32'hfe0d96a;
      56680: inst = 32'h5be00000;
      56681: inst = 32'h8c50000;
      56682: inst = 32'h24612800;
      56683: inst = 32'h10a0ffff;
      56684: inst = 32'hca0fff0;
      56685: inst = 32'h24822800;
      56686: inst = 32'h10a00000;
      56687: inst = 32'hca00004;
      56688: inst = 32'h38632800;
      56689: inst = 32'h38842800;
      56690: inst = 32'h10a00000;
      56691: inst = 32'hca0dd77;
      56692: inst = 32'h13e00001;
      56693: inst = 32'hfe0d96a;
      56694: inst = 32'h5be00000;
      56695: inst = 32'h8c50000;
      56696: inst = 32'h24612800;
      56697: inst = 32'h10a0ffff;
      56698: inst = 32'hca0fff0;
      56699: inst = 32'h24822800;
      56700: inst = 32'h10a00000;
      56701: inst = 32'hca00004;
      56702: inst = 32'h38632800;
      56703: inst = 32'h38842800;
      56704: inst = 32'h10a00000;
      56705: inst = 32'hca0dd85;
      56706: inst = 32'h13e00001;
      56707: inst = 32'hfe0d96a;
      56708: inst = 32'h5be00000;
      56709: inst = 32'h8c50000;
      56710: inst = 32'h24612800;
      56711: inst = 32'h10a0ffff;
      56712: inst = 32'hca0fff0;
      56713: inst = 32'h24822800;
      56714: inst = 32'h10a00000;
      56715: inst = 32'hca00004;
      56716: inst = 32'h38632800;
      56717: inst = 32'h38842800;
      56718: inst = 32'h10a00000;
      56719: inst = 32'hca0dd93;
      56720: inst = 32'h13e00001;
      56721: inst = 32'hfe0d96a;
      56722: inst = 32'h5be00000;
      56723: inst = 32'h8c50000;
      56724: inst = 32'h24612800;
      56725: inst = 32'h10a0ffff;
      56726: inst = 32'hca0fff0;
      56727: inst = 32'h24822800;
      56728: inst = 32'h10a00000;
      56729: inst = 32'hca00004;
      56730: inst = 32'h38632800;
      56731: inst = 32'h38842800;
      56732: inst = 32'h10a00000;
      56733: inst = 32'hca0dda1;
      56734: inst = 32'h13e00001;
      56735: inst = 32'hfe0d96a;
      56736: inst = 32'h5be00000;
      56737: inst = 32'h8c50000;
      56738: inst = 32'h24612800;
      56739: inst = 32'h10a0ffff;
      56740: inst = 32'hca0fff0;
      56741: inst = 32'h24822800;
      56742: inst = 32'h10a00000;
      56743: inst = 32'hca00004;
      56744: inst = 32'h38632800;
      56745: inst = 32'h38842800;
      56746: inst = 32'h10a00000;
      56747: inst = 32'hca0ddaf;
      56748: inst = 32'h13e00001;
      56749: inst = 32'hfe0d96a;
      56750: inst = 32'h5be00000;
      56751: inst = 32'h8c50000;
      56752: inst = 32'h24612800;
      56753: inst = 32'h10a0ffff;
      56754: inst = 32'hca0fff0;
      56755: inst = 32'h24822800;
      56756: inst = 32'h10a00000;
      56757: inst = 32'hca00004;
      56758: inst = 32'h38632800;
      56759: inst = 32'h38842800;
      56760: inst = 32'h10a00000;
      56761: inst = 32'hca0ddbd;
      56762: inst = 32'h13e00001;
      56763: inst = 32'hfe0d96a;
      56764: inst = 32'h5be00000;
      56765: inst = 32'h8c50000;
      56766: inst = 32'h24612800;
      56767: inst = 32'h10a0ffff;
      56768: inst = 32'hca0fff0;
      56769: inst = 32'h24822800;
      56770: inst = 32'h10a00000;
      56771: inst = 32'hca00004;
      56772: inst = 32'h38632800;
      56773: inst = 32'h38842800;
      56774: inst = 32'h10a00000;
      56775: inst = 32'hca0ddcb;
      56776: inst = 32'h13e00001;
      56777: inst = 32'hfe0d96a;
      56778: inst = 32'h5be00000;
      56779: inst = 32'h8c50000;
      56780: inst = 32'h24612800;
      56781: inst = 32'h10a0ffff;
      56782: inst = 32'hca0fff0;
      56783: inst = 32'h24822800;
      56784: inst = 32'h10a00000;
      56785: inst = 32'hca00004;
      56786: inst = 32'h38632800;
      56787: inst = 32'h38842800;
      56788: inst = 32'h10a00000;
      56789: inst = 32'hca0ddd9;
      56790: inst = 32'h13e00001;
      56791: inst = 32'hfe0d96a;
      56792: inst = 32'h5be00000;
      56793: inst = 32'h8c50000;
      56794: inst = 32'h24612800;
      56795: inst = 32'h10a0ffff;
      56796: inst = 32'hca0fff0;
      56797: inst = 32'h24822800;
      56798: inst = 32'h10a00000;
      56799: inst = 32'hca00004;
      56800: inst = 32'h38632800;
      56801: inst = 32'h38842800;
      56802: inst = 32'h10a00000;
      56803: inst = 32'hca0dde7;
      56804: inst = 32'h13e00001;
      56805: inst = 32'hfe0d96a;
      56806: inst = 32'h5be00000;
      56807: inst = 32'h8c50000;
      56808: inst = 32'h24612800;
      56809: inst = 32'h10a0ffff;
      56810: inst = 32'hca0fff0;
      56811: inst = 32'h24822800;
      56812: inst = 32'h10a00000;
      56813: inst = 32'hca00004;
      56814: inst = 32'h38632800;
      56815: inst = 32'h38842800;
      56816: inst = 32'h10a00000;
      56817: inst = 32'hca0ddf5;
      56818: inst = 32'h13e00001;
      56819: inst = 32'hfe0d96a;
      56820: inst = 32'h5be00000;
      56821: inst = 32'h8c50000;
      56822: inst = 32'h24612800;
      56823: inst = 32'h10a0ffff;
      56824: inst = 32'hca0fff0;
      56825: inst = 32'h24822800;
      56826: inst = 32'h10a00000;
      56827: inst = 32'hca00004;
      56828: inst = 32'h38632800;
      56829: inst = 32'h38842800;
      56830: inst = 32'h10a00000;
      56831: inst = 32'hca0de03;
      56832: inst = 32'h13e00001;
      56833: inst = 32'hfe0d96a;
      56834: inst = 32'h5be00000;
      56835: inst = 32'h8c50000;
      56836: inst = 32'h24612800;
      56837: inst = 32'h10a0ffff;
      56838: inst = 32'hca0fff0;
      56839: inst = 32'h24822800;
      56840: inst = 32'h10a00000;
      56841: inst = 32'hca00004;
      56842: inst = 32'h38632800;
      56843: inst = 32'h38842800;
      56844: inst = 32'h10a00000;
      56845: inst = 32'hca0de11;
      56846: inst = 32'h13e00001;
      56847: inst = 32'hfe0d96a;
      56848: inst = 32'h5be00000;
      56849: inst = 32'h8c50000;
      56850: inst = 32'h24612800;
      56851: inst = 32'h10a0ffff;
      56852: inst = 32'hca0fff0;
      56853: inst = 32'h24822800;
      56854: inst = 32'h10a00000;
      56855: inst = 32'hca00004;
      56856: inst = 32'h38632800;
      56857: inst = 32'h38842800;
      56858: inst = 32'h10a00000;
      56859: inst = 32'hca0de1f;
      56860: inst = 32'h13e00001;
      56861: inst = 32'hfe0d96a;
      56862: inst = 32'h5be00000;
      56863: inst = 32'h8c50000;
      56864: inst = 32'h24612800;
      56865: inst = 32'h10a0ffff;
      56866: inst = 32'hca0fff0;
      56867: inst = 32'h24822800;
      56868: inst = 32'h10a00000;
      56869: inst = 32'hca00004;
      56870: inst = 32'h38632800;
      56871: inst = 32'h38842800;
      56872: inst = 32'h10a00000;
      56873: inst = 32'hca0de2d;
      56874: inst = 32'h13e00001;
      56875: inst = 32'hfe0d96a;
      56876: inst = 32'h5be00000;
      56877: inst = 32'h8c50000;
      56878: inst = 32'h24612800;
      56879: inst = 32'h10a0ffff;
      56880: inst = 32'hca0fff0;
      56881: inst = 32'h24822800;
      56882: inst = 32'h10a00000;
      56883: inst = 32'hca00004;
      56884: inst = 32'h38632800;
      56885: inst = 32'h38842800;
      56886: inst = 32'h10a00000;
      56887: inst = 32'hca0de3b;
      56888: inst = 32'h13e00001;
      56889: inst = 32'hfe0d96a;
      56890: inst = 32'h5be00000;
      56891: inst = 32'h8c50000;
      56892: inst = 32'h24612800;
      56893: inst = 32'h10a0ffff;
      56894: inst = 32'hca0fff0;
      56895: inst = 32'h24822800;
      56896: inst = 32'h10a00000;
      56897: inst = 32'hca00004;
      56898: inst = 32'h38632800;
      56899: inst = 32'h38842800;
      56900: inst = 32'h10a00000;
      56901: inst = 32'hca0de49;
      56902: inst = 32'h13e00001;
      56903: inst = 32'hfe0d96a;
      56904: inst = 32'h5be00000;
      56905: inst = 32'h8c50000;
      56906: inst = 32'h24612800;
      56907: inst = 32'h10a0ffff;
      56908: inst = 32'hca0fff0;
      56909: inst = 32'h24822800;
      56910: inst = 32'h10a00000;
      56911: inst = 32'hca00004;
      56912: inst = 32'h38632800;
      56913: inst = 32'h38842800;
      56914: inst = 32'h10a00000;
      56915: inst = 32'hca0de57;
      56916: inst = 32'h13e00001;
      56917: inst = 32'hfe0d96a;
      56918: inst = 32'h5be00000;
      56919: inst = 32'h8c50000;
      56920: inst = 32'h24612800;
      56921: inst = 32'h10a0ffff;
      56922: inst = 32'hca0fff0;
      56923: inst = 32'h24822800;
      56924: inst = 32'h10a00000;
      56925: inst = 32'hca00004;
      56926: inst = 32'h38632800;
      56927: inst = 32'h38842800;
      56928: inst = 32'h10a00000;
      56929: inst = 32'hca0de65;
      56930: inst = 32'h13e00001;
      56931: inst = 32'hfe0d96a;
      56932: inst = 32'h5be00000;
      56933: inst = 32'h8c50000;
      56934: inst = 32'h24612800;
      56935: inst = 32'h10a0ffff;
      56936: inst = 32'hca0fff0;
      56937: inst = 32'h24822800;
      56938: inst = 32'h10a00000;
      56939: inst = 32'hca00004;
      56940: inst = 32'h38632800;
      56941: inst = 32'h38842800;
      56942: inst = 32'h10a00000;
      56943: inst = 32'hca0de73;
      56944: inst = 32'h13e00001;
      56945: inst = 32'hfe0d96a;
      56946: inst = 32'h5be00000;
      56947: inst = 32'h8c50000;
      56948: inst = 32'h24612800;
      56949: inst = 32'h10a0ffff;
      56950: inst = 32'hca0fff0;
      56951: inst = 32'h24822800;
      56952: inst = 32'h10a00000;
      56953: inst = 32'hca00004;
      56954: inst = 32'h38632800;
      56955: inst = 32'h38842800;
      56956: inst = 32'h10a00000;
      56957: inst = 32'hca0de81;
      56958: inst = 32'h13e00001;
      56959: inst = 32'hfe0d96a;
      56960: inst = 32'h5be00000;
      56961: inst = 32'h8c50000;
      56962: inst = 32'h24612800;
      56963: inst = 32'h10a0ffff;
      56964: inst = 32'hca0fff0;
      56965: inst = 32'h24822800;
      56966: inst = 32'h10a00000;
      56967: inst = 32'hca00004;
      56968: inst = 32'h38632800;
      56969: inst = 32'h38842800;
      56970: inst = 32'h10a00000;
      56971: inst = 32'hca0de8f;
      56972: inst = 32'h13e00001;
      56973: inst = 32'hfe0d96a;
      56974: inst = 32'h5be00000;
      56975: inst = 32'h8c50000;
      56976: inst = 32'h24612800;
      56977: inst = 32'h10a0ffff;
      56978: inst = 32'hca0fff0;
      56979: inst = 32'h24822800;
      56980: inst = 32'h10a00000;
      56981: inst = 32'hca00004;
      56982: inst = 32'h38632800;
      56983: inst = 32'h38842800;
      56984: inst = 32'h10a00000;
      56985: inst = 32'hca0de9d;
      56986: inst = 32'h13e00001;
      56987: inst = 32'hfe0d96a;
      56988: inst = 32'h5be00000;
      56989: inst = 32'h8c50000;
      56990: inst = 32'h24612800;
      56991: inst = 32'h10a0ffff;
      56992: inst = 32'hca0fff0;
      56993: inst = 32'h24822800;
      56994: inst = 32'h10a00000;
      56995: inst = 32'hca00004;
      56996: inst = 32'h38632800;
      56997: inst = 32'h38842800;
      56998: inst = 32'h10a00000;
      56999: inst = 32'hca0deab;
      57000: inst = 32'h13e00001;
      57001: inst = 32'hfe0d96a;
      57002: inst = 32'h5be00000;
      57003: inst = 32'h8c50000;
      57004: inst = 32'h24612800;
      57005: inst = 32'h10a0ffff;
      57006: inst = 32'hca0fff0;
      57007: inst = 32'h24822800;
      57008: inst = 32'h10a00000;
      57009: inst = 32'hca00004;
      57010: inst = 32'h38632800;
      57011: inst = 32'h38842800;
      57012: inst = 32'h10a00000;
      57013: inst = 32'hca0deb9;
      57014: inst = 32'h13e00001;
      57015: inst = 32'hfe0d96a;
      57016: inst = 32'h5be00000;
      57017: inst = 32'h8c50000;
      57018: inst = 32'h24612800;
      57019: inst = 32'h10a0ffff;
      57020: inst = 32'hca0fff0;
      57021: inst = 32'h24822800;
      57022: inst = 32'h10a00000;
      57023: inst = 32'hca00004;
      57024: inst = 32'h38632800;
      57025: inst = 32'h38842800;
      57026: inst = 32'h10a00000;
      57027: inst = 32'hca0dec7;
      57028: inst = 32'h13e00001;
      57029: inst = 32'hfe0d96a;
      57030: inst = 32'h5be00000;
      57031: inst = 32'h8c50000;
      57032: inst = 32'h24612800;
      57033: inst = 32'h10a0ffff;
      57034: inst = 32'hca0fff0;
      57035: inst = 32'h24822800;
      57036: inst = 32'h10a00000;
      57037: inst = 32'hca00004;
      57038: inst = 32'h38632800;
      57039: inst = 32'h38842800;
      57040: inst = 32'h10a00000;
      57041: inst = 32'hca0ded5;
      57042: inst = 32'h13e00001;
      57043: inst = 32'hfe0d96a;
      57044: inst = 32'h5be00000;
      57045: inst = 32'h8c50000;
      57046: inst = 32'h24612800;
      57047: inst = 32'h10a0ffff;
      57048: inst = 32'hca0fff0;
      57049: inst = 32'h24822800;
      57050: inst = 32'h10a00000;
      57051: inst = 32'hca00004;
      57052: inst = 32'h38632800;
      57053: inst = 32'h38842800;
      57054: inst = 32'h10a00000;
      57055: inst = 32'hca0dee3;
      57056: inst = 32'h13e00001;
      57057: inst = 32'hfe0d96a;
      57058: inst = 32'h5be00000;
      57059: inst = 32'h8c50000;
      57060: inst = 32'h24612800;
      57061: inst = 32'h10a0ffff;
      57062: inst = 32'hca0fff0;
      57063: inst = 32'h24822800;
      57064: inst = 32'h10a00000;
      57065: inst = 32'hca00004;
      57066: inst = 32'h38632800;
      57067: inst = 32'h38842800;
      57068: inst = 32'h10a00000;
      57069: inst = 32'hca0def1;
      57070: inst = 32'h13e00001;
      57071: inst = 32'hfe0d96a;
      57072: inst = 32'h5be00000;
      57073: inst = 32'h8c50000;
      57074: inst = 32'h24612800;
      57075: inst = 32'h10a0ffff;
      57076: inst = 32'hca0fff0;
      57077: inst = 32'h24822800;
      57078: inst = 32'h10a00000;
      57079: inst = 32'hca00004;
      57080: inst = 32'h38632800;
      57081: inst = 32'h38842800;
      57082: inst = 32'h10a00000;
      57083: inst = 32'hca0deff;
      57084: inst = 32'h13e00001;
      57085: inst = 32'hfe0d96a;
      57086: inst = 32'h5be00000;
      57087: inst = 32'h8c50000;
      57088: inst = 32'h24612800;
      57089: inst = 32'h10a0ffff;
      57090: inst = 32'hca0fff0;
      57091: inst = 32'h24822800;
      57092: inst = 32'h10a00000;
      57093: inst = 32'hca00004;
      57094: inst = 32'h38632800;
      57095: inst = 32'h38842800;
      57096: inst = 32'h10a00000;
      57097: inst = 32'hca0df0d;
      57098: inst = 32'h13e00001;
      57099: inst = 32'hfe0d96a;
      57100: inst = 32'h5be00000;
      57101: inst = 32'h8c50000;
      57102: inst = 32'h24612800;
      57103: inst = 32'h10a0ffff;
      57104: inst = 32'hca0fff0;
      57105: inst = 32'h24822800;
      57106: inst = 32'h10a00000;
      57107: inst = 32'hca00004;
      57108: inst = 32'h38632800;
      57109: inst = 32'h38842800;
      57110: inst = 32'h10a00000;
      57111: inst = 32'hca0df1b;
      57112: inst = 32'h13e00001;
      57113: inst = 32'hfe0d96a;
      57114: inst = 32'h5be00000;
      57115: inst = 32'h8c50000;
      57116: inst = 32'h24612800;
      57117: inst = 32'h10a0ffff;
      57118: inst = 32'hca0fff0;
      57119: inst = 32'h24822800;
      57120: inst = 32'h10a00000;
      57121: inst = 32'hca00004;
      57122: inst = 32'h38632800;
      57123: inst = 32'h38842800;
      57124: inst = 32'h10a00000;
      57125: inst = 32'hca0df29;
      57126: inst = 32'h13e00001;
      57127: inst = 32'hfe0d96a;
      57128: inst = 32'h5be00000;
      57129: inst = 32'h8c50000;
      57130: inst = 32'h24612800;
      57131: inst = 32'h10a0ffff;
      57132: inst = 32'hca0fff0;
      57133: inst = 32'h24822800;
      57134: inst = 32'h10a00000;
      57135: inst = 32'hca00004;
      57136: inst = 32'h38632800;
      57137: inst = 32'h38842800;
      57138: inst = 32'h10a00000;
      57139: inst = 32'hca0df37;
      57140: inst = 32'h13e00001;
      57141: inst = 32'hfe0d96a;
      57142: inst = 32'h5be00000;
      57143: inst = 32'h8c50000;
      57144: inst = 32'h24612800;
      57145: inst = 32'h10a0ffff;
      57146: inst = 32'hca0fff0;
      57147: inst = 32'h24822800;
      57148: inst = 32'h10a00000;
      57149: inst = 32'hca00004;
      57150: inst = 32'h38632800;
      57151: inst = 32'h38842800;
      57152: inst = 32'h10a00000;
      57153: inst = 32'hca0df45;
      57154: inst = 32'h13e00001;
      57155: inst = 32'hfe0d96a;
      57156: inst = 32'h5be00000;
      57157: inst = 32'h8c50000;
      57158: inst = 32'h24612800;
      57159: inst = 32'h10a0ffff;
      57160: inst = 32'hca0fff0;
      57161: inst = 32'h24822800;
      57162: inst = 32'h10a00000;
      57163: inst = 32'hca00004;
      57164: inst = 32'h38632800;
      57165: inst = 32'h38842800;
      57166: inst = 32'h10a00000;
      57167: inst = 32'hca0df53;
      57168: inst = 32'h13e00001;
      57169: inst = 32'hfe0d96a;
      57170: inst = 32'h5be00000;
      57171: inst = 32'h8c50000;
      57172: inst = 32'h24612800;
      57173: inst = 32'h10a0ffff;
      57174: inst = 32'hca0fff0;
      57175: inst = 32'h24822800;
      57176: inst = 32'h10a00000;
      57177: inst = 32'hca00004;
      57178: inst = 32'h38632800;
      57179: inst = 32'h38842800;
      57180: inst = 32'h10a00000;
      57181: inst = 32'hca0df61;
      57182: inst = 32'h13e00001;
      57183: inst = 32'hfe0d96a;
      57184: inst = 32'h5be00000;
      57185: inst = 32'h8c50000;
      57186: inst = 32'h24612800;
      57187: inst = 32'h10a0ffff;
      57188: inst = 32'hca0fff0;
      57189: inst = 32'h24822800;
      57190: inst = 32'h10a00000;
      57191: inst = 32'hca00004;
      57192: inst = 32'h38632800;
      57193: inst = 32'h38842800;
      57194: inst = 32'h10a00000;
      57195: inst = 32'hca0df6f;
      57196: inst = 32'h13e00001;
      57197: inst = 32'hfe0d96a;
      57198: inst = 32'h5be00000;
      57199: inst = 32'h8c50000;
      57200: inst = 32'h24612800;
      57201: inst = 32'h10a0ffff;
      57202: inst = 32'hca0fff0;
      57203: inst = 32'h24822800;
      57204: inst = 32'h10a00000;
      57205: inst = 32'hca00004;
      57206: inst = 32'h38632800;
      57207: inst = 32'h38842800;
      57208: inst = 32'h10a00000;
      57209: inst = 32'hca0df7d;
      57210: inst = 32'h13e00001;
      57211: inst = 32'hfe0d96a;
      57212: inst = 32'h5be00000;
      57213: inst = 32'h8c50000;
      57214: inst = 32'h24612800;
      57215: inst = 32'h10a0ffff;
      57216: inst = 32'hca0fff0;
      57217: inst = 32'h24822800;
      57218: inst = 32'h10a00000;
      57219: inst = 32'hca00004;
      57220: inst = 32'h38632800;
      57221: inst = 32'h38842800;
      57222: inst = 32'h10a00000;
      57223: inst = 32'hca0df8b;
      57224: inst = 32'h13e00001;
      57225: inst = 32'hfe0d96a;
      57226: inst = 32'h5be00000;
      57227: inst = 32'h8c50000;
      57228: inst = 32'h24612800;
      57229: inst = 32'h10a0ffff;
      57230: inst = 32'hca0fff0;
      57231: inst = 32'h24822800;
      57232: inst = 32'h10a00000;
      57233: inst = 32'hca00004;
      57234: inst = 32'h38632800;
      57235: inst = 32'h38842800;
      57236: inst = 32'h10a00000;
      57237: inst = 32'hca0df99;
      57238: inst = 32'h13e00001;
      57239: inst = 32'hfe0d96a;
      57240: inst = 32'h5be00000;
      57241: inst = 32'h8c50000;
      57242: inst = 32'h24612800;
      57243: inst = 32'h10a0ffff;
      57244: inst = 32'hca0fff0;
      57245: inst = 32'h24822800;
      57246: inst = 32'h10a00000;
      57247: inst = 32'hca00004;
      57248: inst = 32'h38632800;
      57249: inst = 32'h38842800;
      57250: inst = 32'h10a00000;
      57251: inst = 32'hca0dfa7;
      57252: inst = 32'h13e00001;
      57253: inst = 32'hfe0d96a;
      57254: inst = 32'h5be00000;
      57255: inst = 32'h8c50000;
      57256: inst = 32'h24612800;
      57257: inst = 32'h10a0ffff;
      57258: inst = 32'hca0fff0;
      57259: inst = 32'h24822800;
      57260: inst = 32'h10a00000;
      57261: inst = 32'hca00004;
      57262: inst = 32'h38632800;
      57263: inst = 32'h38842800;
      57264: inst = 32'h10a00000;
      57265: inst = 32'hca0dfb5;
      57266: inst = 32'h13e00001;
      57267: inst = 32'hfe0d96a;
      57268: inst = 32'h5be00000;
      57269: inst = 32'h8c50000;
      57270: inst = 32'h24612800;
      57271: inst = 32'h10a0ffff;
      57272: inst = 32'hca0fff0;
      57273: inst = 32'h24822800;
      57274: inst = 32'h10a00000;
      57275: inst = 32'hca00004;
      57276: inst = 32'h38632800;
      57277: inst = 32'h38842800;
      57278: inst = 32'h10a00000;
      57279: inst = 32'hca0dfc3;
      57280: inst = 32'h13e00001;
      57281: inst = 32'hfe0d96a;
      57282: inst = 32'h5be00000;
      57283: inst = 32'h8c50000;
      57284: inst = 32'h24612800;
      57285: inst = 32'h10a0ffff;
      57286: inst = 32'hca0fff0;
      57287: inst = 32'h24822800;
      57288: inst = 32'h10a00000;
      57289: inst = 32'hca00004;
      57290: inst = 32'h38632800;
      57291: inst = 32'h38842800;
      57292: inst = 32'h10a00000;
      57293: inst = 32'hca0dfd1;
      57294: inst = 32'h13e00001;
      57295: inst = 32'hfe0d96a;
      57296: inst = 32'h5be00000;
      57297: inst = 32'h8c50000;
      57298: inst = 32'h24612800;
      57299: inst = 32'h10a0ffff;
      57300: inst = 32'hca0fff0;
      57301: inst = 32'h24822800;
      57302: inst = 32'h10a00000;
      57303: inst = 32'hca00004;
      57304: inst = 32'h38632800;
      57305: inst = 32'h38842800;
      57306: inst = 32'h10a00000;
      57307: inst = 32'hca0dfdf;
      57308: inst = 32'h13e00001;
      57309: inst = 32'hfe0d96a;
      57310: inst = 32'h5be00000;
      57311: inst = 32'h8c50000;
      57312: inst = 32'h24612800;
      57313: inst = 32'h10a0ffff;
      57314: inst = 32'hca0fff0;
      57315: inst = 32'h24822800;
      57316: inst = 32'h10a00000;
      57317: inst = 32'hca00004;
      57318: inst = 32'h38632800;
      57319: inst = 32'h38842800;
      57320: inst = 32'h10a00000;
      57321: inst = 32'hca0dfed;
      57322: inst = 32'h13e00001;
      57323: inst = 32'hfe0d96a;
      57324: inst = 32'h5be00000;
      57325: inst = 32'h8c50000;
      57326: inst = 32'h24612800;
      57327: inst = 32'h10a0ffff;
      57328: inst = 32'hca0fff0;
      57329: inst = 32'h24822800;
      57330: inst = 32'h10a00000;
      57331: inst = 32'hca00004;
      57332: inst = 32'h38632800;
      57333: inst = 32'h38842800;
      57334: inst = 32'h10a00000;
      57335: inst = 32'hca0dffb;
      57336: inst = 32'h13e00001;
      57337: inst = 32'hfe0d96a;
      57338: inst = 32'h5be00000;
      57339: inst = 32'h8c50000;
      57340: inst = 32'h24612800;
      57341: inst = 32'h10a0ffff;
      57342: inst = 32'hca0fff0;
      57343: inst = 32'h24822800;
      57344: inst = 32'h10a00000;
      57345: inst = 32'hca00004;
      57346: inst = 32'h38632800;
      57347: inst = 32'h38842800;
      57348: inst = 32'h10a00000;
      57349: inst = 32'hca0e009;
      57350: inst = 32'h13e00001;
      57351: inst = 32'hfe0d96a;
      57352: inst = 32'h5be00000;
      57353: inst = 32'h8c50000;
      57354: inst = 32'h24612800;
      57355: inst = 32'h10a0ffff;
      57356: inst = 32'hca0fff0;
      57357: inst = 32'h24822800;
      57358: inst = 32'h10a00000;
      57359: inst = 32'hca00004;
      57360: inst = 32'h38632800;
      57361: inst = 32'h38842800;
      57362: inst = 32'h10a00000;
      57363: inst = 32'hca0e017;
      57364: inst = 32'h13e00001;
      57365: inst = 32'hfe0d96a;
      57366: inst = 32'h5be00000;
      57367: inst = 32'h8c50000;
      57368: inst = 32'h24612800;
      57369: inst = 32'h10a0ffff;
      57370: inst = 32'hca0fff0;
      57371: inst = 32'h24822800;
      57372: inst = 32'h10a00000;
      57373: inst = 32'hca00004;
      57374: inst = 32'h38632800;
      57375: inst = 32'h38842800;
      57376: inst = 32'h10a00000;
      57377: inst = 32'hca0e025;
      57378: inst = 32'h13e00001;
      57379: inst = 32'hfe0d96a;
      57380: inst = 32'h5be00000;
      57381: inst = 32'h8c50000;
      57382: inst = 32'h24612800;
      57383: inst = 32'h10a0ffff;
      57384: inst = 32'hca0fff0;
      57385: inst = 32'h24822800;
      57386: inst = 32'h10a00000;
      57387: inst = 32'hca00004;
      57388: inst = 32'h38632800;
      57389: inst = 32'h38842800;
      57390: inst = 32'h10a00000;
      57391: inst = 32'hca0e033;
      57392: inst = 32'h13e00001;
      57393: inst = 32'hfe0d96a;
      57394: inst = 32'h5be00000;
      57395: inst = 32'h8c50000;
      57396: inst = 32'h24612800;
      57397: inst = 32'h10a0ffff;
      57398: inst = 32'hca0fff0;
      57399: inst = 32'h24822800;
      57400: inst = 32'h10a00000;
      57401: inst = 32'hca00004;
      57402: inst = 32'h38632800;
      57403: inst = 32'h38842800;
      57404: inst = 32'h10a00000;
      57405: inst = 32'hca0e041;
      57406: inst = 32'h13e00001;
      57407: inst = 32'hfe0d96a;
      57408: inst = 32'h5be00000;
      57409: inst = 32'h8c50000;
      57410: inst = 32'h24612800;
      57411: inst = 32'h10a0ffff;
      57412: inst = 32'hca0fff0;
      57413: inst = 32'h24822800;
      57414: inst = 32'h10a00000;
      57415: inst = 32'hca00004;
      57416: inst = 32'h38632800;
      57417: inst = 32'h38842800;
      57418: inst = 32'h10a00000;
      57419: inst = 32'hca0e04f;
      57420: inst = 32'h13e00001;
      57421: inst = 32'hfe0d96a;
      57422: inst = 32'h5be00000;
      57423: inst = 32'h8c50000;
      57424: inst = 32'h24612800;
      57425: inst = 32'h10a0ffff;
      57426: inst = 32'hca0fff0;
      57427: inst = 32'h24822800;
      57428: inst = 32'h10a00000;
      57429: inst = 32'hca00004;
      57430: inst = 32'h38632800;
      57431: inst = 32'h38842800;
      57432: inst = 32'h10a00000;
      57433: inst = 32'hca0e05d;
      57434: inst = 32'h13e00001;
      57435: inst = 32'hfe0d96a;
      57436: inst = 32'h5be00000;
      57437: inst = 32'h8c50000;
      57438: inst = 32'h24612800;
      57439: inst = 32'h10a0ffff;
      57440: inst = 32'hca0fff0;
      57441: inst = 32'h24822800;
      57442: inst = 32'h10a00000;
      57443: inst = 32'hca00004;
      57444: inst = 32'h38632800;
      57445: inst = 32'h38842800;
      57446: inst = 32'h10a00000;
      57447: inst = 32'hca0e06b;
      57448: inst = 32'h13e00001;
      57449: inst = 32'hfe0d96a;
      57450: inst = 32'h5be00000;
      57451: inst = 32'h8c50000;
      57452: inst = 32'h24612800;
      57453: inst = 32'h10a0ffff;
      57454: inst = 32'hca0fff0;
      57455: inst = 32'h24822800;
      57456: inst = 32'h10a00000;
      57457: inst = 32'hca00004;
      57458: inst = 32'h38632800;
      57459: inst = 32'h38842800;
      57460: inst = 32'h10a00000;
      57461: inst = 32'hca0e079;
      57462: inst = 32'h13e00001;
      57463: inst = 32'hfe0d96a;
      57464: inst = 32'h5be00000;
      57465: inst = 32'h8c50000;
      57466: inst = 32'h24612800;
      57467: inst = 32'h10a0ffff;
      57468: inst = 32'hca0fff0;
      57469: inst = 32'h24822800;
      57470: inst = 32'h10a00000;
      57471: inst = 32'hca00004;
      57472: inst = 32'h38632800;
      57473: inst = 32'h38842800;
      57474: inst = 32'h10a00000;
      57475: inst = 32'hca0e087;
      57476: inst = 32'h13e00001;
      57477: inst = 32'hfe0d96a;
      57478: inst = 32'h5be00000;
      57479: inst = 32'h8c50000;
      57480: inst = 32'h24612800;
      57481: inst = 32'h10a0ffff;
      57482: inst = 32'hca0fff0;
      57483: inst = 32'h24822800;
      57484: inst = 32'h10a00000;
      57485: inst = 32'hca00004;
      57486: inst = 32'h38632800;
      57487: inst = 32'h38842800;
      57488: inst = 32'h10a00000;
      57489: inst = 32'hca0e095;
      57490: inst = 32'h13e00001;
      57491: inst = 32'hfe0d96a;
      57492: inst = 32'h5be00000;
      57493: inst = 32'h8c50000;
      57494: inst = 32'h24612800;
      57495: inst = 32'h10a0ffff;
      57496: inst = 32'hca0fff0;
      57497: inst = 32'h24822800;
      57498: inst = 32'h10a00000;
      57499: inst = 32'hca00004;
      57500: inst = 32'h38632800;
      57501: inst = 32'h38842800;
      57502: inst = 32'h10a00000;
      57503: inst = 32'hca0e0a3;
      57504: inst = 32'h13e00001;
      57505: inst = 32'hfe0d96a;
      57506: inst = 32'h5be00000;
      57507: inst = 32'h8c50000;
      57508: inst = 32'h24612800;
      57509: inst = 32'h10a0ffff;
      57510: inst = 32'hca0fff0;
      57511: inst = 32'h24822800;
      57512: inst = 32'h10a00000;
      57513: inst = 32'hca00004;
      57514: inst = 32'h38632800;
      57515: inst = 32'h38842800;
      57516: inst = 32'h10a00000;
      57517: inst = 32'hca0e0b1;
      57518: inst = 32'h13e00001;
      57519: inst = 32'hfe0d96a;
      57520: inst = 32'h5be00000;
      57521: inst = 32'h8c50000;
      57522: inst = 32'h24612800;
      57523: inst = 32'h10a0ffff;
      57524: inst = 32'hca0fff0;
      57525: inst = 32'h24822800;
      57526: inst = 32'h10a00000;
      57527: inst = 32'hca00004;
      57528: inst = 32'h38632800;
      57529: inst = 32'h38842800;
      57530: inst = 32'h10a00000;
      57531: inst = 32'hca0e0bf;
      57532: inst = 32'h13e00001;
      57533: inst = 32'hfe0d96a;
      57534: inst = 32'h5be00000;
      57535: inst = 32'h8c50000;
      57536: inst = 32'h24612800;
      57537: inst = 32'h10a0ffff;
      57538: inst = 32'hca0fff0;
      57539: inst = 32'h24822800;
      57540: inst = 32'h10a00000;
      57541: inst = 32'hca00004;
      57542: inst = 32'h38632800;
      57543: inst = 32'h38842800;
      57544: inst = 32'h10a00000;
      57545: inst = 32'hca0e0cd;
      57546: inst = 32'h13e00001;
      57547: inst = 32'hfe0d96a;
      57548: inst = 32'h5be00000;
      57549: inst = 32'h8c50000;
      57550: inst = 32'h24612800;
      57551: inst = 32'h10a0ffff;
      57552: inst = 32'hca0fff0;
      57553: inst = 32'h24822800;
      57554: inst = 32'h10a00000;
      57555: inst = 32'hca00004;
      57556: inst = 32'h38632800;
      57557: inst = 32'h38842800;
      57558: inst = 32'h10a00000;
      57559: inst = 32'hca0e0db;
      57560: inst = 32'h13e00001;
      57561: inst = 32'hfe0d96a;
      57562: inst = 32'h5be00000;
      57563: inst = 32'h8c50000;
      57564: inst = 32'h24612800;
      57565: inst = 32'h10a0ffff;
      57566: inst = 32'hca0fff0;
      57567: inst = 32'h24822800;
      57568: inst = 32'h10a00000;
      57569: inst = 32'hca00004;
      57570: inst = 32'h38632800;
      57571: inst = 32'h38842800;
      57572: inst = 32'h10a00000;
      57573: inst = 32'hca0e0e9;
      57574: inst = 32'h13e00001;
      57575: inst = 32'hfe0d96a;
      57576: inst = 32'h5be00000;
      57577: inst = 32'h8c50000;
      57578: inst = 32'h24612800;
      57579: inst = 32'h10a0ffff;
      57580: inst = 32'hca0fff0;
      57581: inst = 32'h24822800;
      57582: inst = 32'h10a00000;
      57583: inst = 32'hca00004;
      57584: inst = 32'h38632800;
      57585: inst = 32'h38842800;
      57586: inst = 32'h10a00000;
      57587: inst = 32'hca0e0f7;
      57588: inst = 32'h13e00001;
      57589: inst = 32'hfe0d96a;
      57590: inst = 32'h5be00000;
      57591: inst = 32'h8c50000;
      57592: inst = 32'h24612800;
      57593: inst = 32'h10a0ffff;
      57594: inst = 32'hca0fff0;
      57595: inst = 32'h24822800;
      57596: inst = 32'h10a00000;
      57597: inst = 32'hca00004;
      57598: inst = 32'h38632800;
      57599: inst = 32'h38842800;
      57600: inst = 32'h10a00000;
      57601: inst = 32'hca0e105;
      57602: inst = 32'h13e00001;
      57603: inst = 32'hfe0d96a;
      57604: inst = 32'h5be00000;
      57605: inst = 32'h8c50000;
      57606: inst = 32'h24612800;
      57607: inst = 32'h10a0ffff;
      57608: inst = 32'hca0fff0;
      57609: inst = 32'h24822800;
      57610: inst = 32'h10a00000;
      57611: inst = 32'hca00004;
      57612: inst = 32'h38632800;
      57613: inst = 32'h38842800;
      57614: inst = 32'h10a00000;
      57615: inst = 32'hca0e113;
      57616: inst = 32'h13e00001;
      57617: inst = 32'hfe0d96a;
      57618: inst = 32'h5be00000;
      57619: inst = 32'h8c50000;
      57620: inst = 32'h24612800;
      57621: inst = 32'h10a0ffff;
      57622: inst = 32'hca0fff0;
      57623: inst = 32'h24822800;
      57624: inst = 32'h10a00000;
      57625: inst = 32'hca00004;
      57626: inst = 32'h38632800;
      57627: inst = 32'h38842800;
      57628: inst = 32'h10a00000;
      57629: inst = 32'hca0e121;
      57630: inst = 32'h13e00001;
      57631: inst = 32'hfe0d96a;
      57632: inst = 32'h5be00000;
      57633: inst = 32'h8c50000;
      57634: inst = 32'h24612800;
      57635: inst = 32'h10a0ffff;
      57636: inst = 32'hca0fff0;
      57637: inst = 32'h24822800;
      57638: inst = 32'h10a00000;
      57639: inst = 32'hca00004;
      57640: inst = 32'h38632800;
      57641: inst = 32'h38842800;
      57642: inst = 32'h10a00000;
      57643: inst = 32'hca0e12f;
      57644: inst = 32'h13e00001;
      57645: inst = 32'hfe0d96a;
      57646: inst = 32'h5be00000;
      57647: inst = 32'h8c50000;
      57648: inst = 32'h24612800;
      57649: inst = 32'h10a0ffff;
      57650: inst = 32'hca0fff0;
      57651: inst = 32'h24822800;
      57652: inst = 32'h10a00000;
      57653: inst = 32'hca00004;
      57654: inst = 32'h38632800;
      57655: inst = 32'h38842800;
      57656: inst = 32'h10a00000;
      57657: inst = 32'hca0e13d;
      57658: inst = 32'h13e00001;
      57659: inst = 32'hfe0d96a;
      57660: inst = 32'h5be00000;
      57661: inst = 32'h8c50000;
      57662: inst = 32'h24612800;
      57663: inst = 32'h10a0ffff;
      57664: inst = 32'hca0fff0;
      57665: inst = 32'h24822800;
      57666: inst = 32'h10a00000;
      57667: inst = 32'hca00004;
      57668: inst = 32'h38632800;
      57669: inst = 32'h38842800;
      57670: inst = 32'h10a00000;
      57671: inst = 32'hca0e14b;
      57672: inst = 32'h13e00001;
      57673: inst = 32'hfe0d96a;
      57674: inst = 32'h5be00000;
      57675: inst = 32'h8c50000;
      57676: inst = 32'h24612800;
      57677: inst = 32'h10a0ffff;
      57678: inst = 32'hca0fff0;
      57679: inst = 32'h24822800;
      57680: inst = 32'h10a00000;
      57681: inst = 32'hca00004;
      57682: inst = 32'h38632800;
      57683: inst = 32'h38842800;
      57684: inst = 32'h10a00000;
      57685: inst = 32'hca0e159;
      57686: inst = 32'h13e00001;
      57687: inst = 32'hfe0d96a;
      57688: inst = 32'h5be00000;
      57689: inst = 32'h8c50000;
      57690: inst = 32'h24612800;
      57691: inst = 32'h10a0ffff;
      57692: inst = 32'hca0fff0;
      57693: inst = 32'h24822800;
      57694: inst = 32'h10a00000;
      57695: inst = 32'hca00004;
      57696: inst = 32'h38632800;
      57697: inst = 32'h38842800;
      57698: inst = 32'h10a00000;
      57699: inst = 32'hca0e167;
      57700: inst = 32'h13e00001;
      57701: inst = 32'hfe0d96a;
      57702: inst = 32'h5be00000;
      57703: inst = 32'h8c50000;
      57704: inst = 32'h24612800;
      57705: inst = 32'h10a0ffff;
      57706: inst = 32'hca0fff0;
      57707: inst = 32'h24822800;
      57708: inst = 32'h10a00000;
      57709: inst = 32'hca00004;
      57710: inst = 32'h38632800;
      57711: inst = 32'h38842800;
      57712: inst = 32'h10a00000;
      57713: inst = 32'hca0e175;
      57714: inst = 32'h13e00001;
      57715: inst = 32'hfe0d96a;
      57716: inst = 32'h5be00000;
      57717: inst = 32'h8c50000;
      57718: inst = 32'h24612800;
      57719: inst = 32'h10a0ffff;
      57720: inst = 32'hca0fff0;
      57721: inst = 32'h24822800;
      57722: inst = 32'h10a00000;
      57723: inst = 32'hca00004;
      57724: inst = 32'h38632800;
      57725: inst = 32'h38842800;
      57726: inst = 32'h10a00000;
      57727: inst = 32'hca0e183;
      57728: inst = 32'h13e00001;
      57729: inst = 32'hfe0d96a;
      57730: inst = 32'h5be00000;
      57731: inst = 32'h8c50000;
      57732: inst = 32'h24612800;
      57733: inst = 32'h10a0ffff;
      57734: inst = 32'hca0fff0;
      57735: inst = 32'h24822800;
      57736: inst = 32'h10a00000;
      57737: inst = 32'hca00004;
      57738: inst = 32'h38632800;
      57739: inst = 32'h38842800;
      57740: inst = 32'h10a00000;
      57741: inst = 32'hca0e191;
      57742: inst = 32'h13e00001;
      57743: inst = 32'hfe0d96a;
      57744: inst = 32'h5be00000;
      57745: inst = 32'h8c50000;
      57746: inst = 32'h24612800;
      57747: inst = 32'h10a0ffff;
      57748: inst = 32'hca0fff0;
      57749: inst = 32'h24822800;
      57750: inst = 32'h10a00000;
      57751: inst = 32'hca00004;
      57752: inst = 32'h38632800;
      57753: inst = 32'h38842800;
      57754: inst = 32'h10a00000;
      57755: inst = 32'hca0e19f;
      57756: inst = 32'h13e00001;
      57757: inst = 32'hfe0d96a;
      57758: inst = 32'h5be00000;
      57759: inst = 32'h8c50000;
      57760: inst = 32'h24612800;
      57761: inst = 32'h10a0ffff;
      57762: inst = 32'hca0fff0;
      57763: inst = 32'h24822800;
      57764: inst = 32'h10a00000;
      57765: inst = 32'hca00004;
      57766: inst = 32'h38632800;
      57767: inst = 32'h38842800;
      57768: inst = 32'h10a00000;
      57769: inst = 32'hca0e1ad;
      57770: inst = 32'h13e00001;
      57771: inst = 32'hfe0d96a;
      57772: inst = 32'h5be00000;
      57773: inst = 32'h8c50000;
      57774: inst = 32'h24612800;
      57775: inst = 32'h10a0ffff;
      57776: inst = 32'hca0fff0;
      57777: inst = 32'h24822800;
      57778: inst = 32'h10a00000;
      57779: inst = 32'hca00004;
      57780: inst = 32'h38632800;
      57781: inst = 32'h38842800;
      57782: inst = 32'h10a00000;
      57783: inst = 32'hca0e1bb;
      57784: inst = 32'h13e00001;
      57785: inst = 32'hfe0d96a;
      57786: inst = 32'h5be00000;
      57787: inst = 32'h8c50000;
      57788: inst = 32'h24612800;
      57789: inst = 32'h10a0ffff;
      57790: inst = 32'hca0fff0;
      57791: inst = 32'h24822800;
      57792: inst = 32'h10a00000;
      57793: inst = 32'hca00004;
      57794: inst = 32'h38632800;
      57795: inst = 32'h38842800;
      57796: inst = 32'h10a00000;
      57797: inst = 32'hca0e1c9;
      57798: inst = 32'h13e00001;
      57799: inst = 32'hfe0d96a;
      57800: inst = 32'h5be00000;
      57801: inst = 32'h8c50000;
      57802: inst = 32'h24612800;
      57803: inst = 32'h10a0ffff;
      57804: inst = 32'hca0fff0;
      57805: inst = 32'h24822800;
      57806: inst = 32'h10a00000;
      57807: inst = 32'hca00004;
      57808: inst = 32'h38632800;
      57809: inst = 32'h38842800;
      57810: inst = 32'h10a00000;
      57811: inst = 32'hca0e1d7;
      57812: inst = 32'h13e00001;
      57813: inst = 32'hfe0d96a;
      57814: inst = 32'h5be00000;
      57815: inst = 32'h8c50000;
      57816: inst = 32'h24612800;
      57817: inst = 32'h10a0ffff;
      57818: inst = 32'hca0fff0;
      57819: inst = 32'h24822800;
      57820: inst = 32'h10a00000;
      57821: inst = 32'hca00004;
      57822: inst = 32'h38632800;
      57823: inst = 32'h38842800;
      57824: inst = 32'h10a00000;
      57825: inst = 32'hca0e1e5;
      57826: inst = 32'h13e00001;
      57827: inst = 32'hfe0d96a;
      57828: inst = 32'h5be00000;
      57829: inst = 32'h8c50000;
      57830: inst = 32'h24612800;
      57831: inst = 32'h10a0ffff;
      57832: inst = 32'hca0fff0;
      57833: inst = 32'h24822800;
      57834: inst = 32'h10a00000;
      57835: inst = 32'hca00004;
      57836: inst = 32'h38632800;
      57837: inst = 32'h38842800;
      57838: inst = 32'h10a00000;
      57839: inst = 32'hca0e1f3;
      57840: inst = 32'h13e00001;
      57841: inst = 32'hfe0d96a;
      57842: inst = 32'h5be00000;
      57843: inst = 32'h8c50000;
      57844: inst = 32'h24612800;
      57845: inst = 32'h10a0ffff;
      57846: inst = 32'hca0fff0;
      57847: inst = 32'h24822800;
      57848: inst = 32'h10a00000;
      57849: inst = 32'hca00004;
      57850: inst = 32'h38632800;
      57851: inst = 32'h38842800;
      57852: inst = 32'h10a00000;
      57853: inst = 32'hca0e201;
      57854: inst = 32'h13e00001;
      57855: inst = 32'hfe0d96a;
      57856: inst = 32'h5be00000;
      57857: inst = 32'h8c50000;
      57858: inst = 32'h24612800;
      57859: inst = 32'h10a0ffff;
      57860: inst = 32'hca0fff0;
      57861: inst = 32'h24822800;
      57862: inst = 32'h10a00000;
      57863: inst = 32'hca00004;
      57864: inst = 32'h38632800;
      57865: inst = 32'h38842800;
      57866: inst = 32'h10a00000;
      57867: inst = 32'hca0e20f;
      57868: inst = 32'h13e00001;
      57869: inst = 32'hfe0d96a;
      57870: inst = 32'h5be00000;
      57871: inst = 32'h8c50000;
      57872: inst = 32'h24612800;
      57873: inst = 32'h10a0ffff;
      57874: inst = 32'hca0fff0;
      57875: inst = 32'h24822800;
      57876: inst = 32'h10a00000;
      57877: inst = 32'hca00004;
      57878: inst = 32'h38632800;
      57879: inst = 32'h38842800;
      57880: inst = 32'h10a00000;
      57881: inst = 32'hca0e21d;
      57882: inst = 32'h13e00001;
      57883: inst = 32'hfe0d96a;
      57884: inst = 32'h5be00000;
      57885: inst = 32'h8c50000;
      57886: inst = 32'h24612800;
      57887: inst = 32'h10a0ffff;
      57888: inst = 32'hca0fff0;
      57889: inst = 32'h24822800;
      57890: inst = 32'h10a00000;
      57891: inst = 32'hca00004;
      57892: inst = 32'h38632800;
      57893: inst = 32'h38842800;
      57894: inst = 32'h10a00000;
      57895: inst = 32'hca0e22b;
      57896: inst = 32'h13e00001;
      57897: inst = 32'hfe0d96a;
      57898: inst = 32'h5be00000;
      57899: inst = 32'h8c50000;
      57900: inst = 32'h24612800;
      57901: inst = 32'h10a0ffff;
      57902: inst = 32'hca0fff0;
      57903: inst = 32'h24822800;
      57904: inst = 32'h10a00000;
      57905: inst = 32'hca00004;
      57906: inst = 32'h38632800;
      57907: inst = 32'h38842800;
      57908: inst = 32'h10a00000;
      57909: inst = 32'hca0e239;
      57910: inst = 32'h13e00001;
      57911: inst = 32'hfe0d96a;
      57912: inst = 32'h5be00000;
      57913: inst = 32'h8c50000;
      57914: inst = 32'h24612800;
      57915: inst = 32'h10a0ffff;
      57916: inst = 32'hca0fff0;
      57917: inst = 32'h24822800;
      57918: inst = 32'h10a00000;
      57919: inst = 32'hca00004;
      57920: inst = 32'h38632800;
      57921: inst = 32'h38842800;
      57922: inst = 32'h10a00000;
      57923: inst = 32'hca0e247;
      57924: inst = 32'h13e00001;
      57925: inst = 32'hfe0d96a;
      57926: inst = 32'h5be00000;
      57927: inst = 32'h8c50000;
      57928: inst = 32'h24612800;
      57929: inst = 32'h10a0ffff;
      57930: inst = 32'hca0fff0;
      57931: inst = 32'h24822800;
      57932: inst = 32'h10a00000;
      57933: inst = 32'hca00004;
      57934: inst = 32'h38632800;
      57935: inst = 32'h38842800;
      57936: inst = 32'h10a00000;
      57937: inst = 32'hca0e255;
      57938: inst = 32'h13e00001;
      57939: inst = 32'hfe0d96a;
      57940: inst = 32'h5be00000;
      57941: inst = 32'h8c50000;
      57942: inst = 32'h24612800;
      57943: inst = 32'h10a0ffff;
      57944: inst = 32'hca0fff0;
      57945: inst = 32'h24822800;
      57946: inst = 32'h10a00000;
      57947: inst = 32'hca00004;
      57948: inst = 32'h38632800;
      57949: inst = 32'h38842800;
      57950: inst = 32'h10a00000;
      57951: inst = 32'hca0e263;
      57952: inst = 32'h13e00001;
      57953: inst = 32'hfe0d96a;
      57954: inst = 32'h5be00000;
      57955: inst = 32'h8c50000;
      57956: inst = 32'h24612800;
      57957: inst = 32'h10a0ffff;
      57958: inst = 32'hca0fff0;
      57959: inst = 32'h24822800;
      57960: inst = 32'h10a00000;
      57961: inst = 32'hca00004;
      57962: inst = 32'h38632800;
      57963: inst = 32'h38842800;
      57964: inst = 32'h10a00000;
      57965: inst = 32'hca0e271;
      57966: inst = 32'h13e00001;
      57967: inst = 32'hfe0d96a;
      57968: inst = 32'h5be00000;
      57969: inst = 32'h8c50000;
      57970: inst = 32'h24612800;
      57971: inst = 32'h10a0ffff;
      57972: inst = 32'hca0fff0;
      57973: inst = 32'h24822800;
      57974: inst = 32'h10a00000;
      57975: inst = 32'hca00004;
      57976: inst = 32'h38632800;
      57977: inst = 32'h38842800;
      57978: inst = 32'h10a00000;
      57979: inst = 32'hca0e27f;
      57980: inst = 32'h13e00001;
      57981: inst = 32'hfe0d96a;
      57982: inst = 32'h5be00000;
      57983: inst = 32'h8c50000;
      57984: inst = 32'h24612800;
      57985: inst = 32'h10a0ffff;
      57986: inst = 32'hca0fff0;
      57987: inst = 32'h24822800;
      57988: inst = 32'h10a00000;
      57989: inst = 32'hca00004;
      57990: inst = 32'h38632800;
      57991: inst = 32'h38842800;
      57992: inst = 32'h10a00000;
      57993: inst = 32'hca0e28d;
      57994: inst = 32'h13e00001;
      57995: inst = 32'hfe0d96a;
      57996: inst = 32'h5be00000;
      57997: inst = 32'h8c50000;
      57998: inst = 32'h24612800;
      57999: inst = 32'h10a0ffff;
      58000: inst = 32'hca0fff0;
      58001: inst = 32'h24822800;
      58002: inst = 32'h10a00000;
      58003: inst = 32'hca00004;
      58004: inst = 32'h38632800;
      58005: inst = 32'h38842800;
      58006: inst = 32'h10a00000;
      58007: inst = 32'hca0e29b;
      58008: inst = 32'h13e00001;
      58009: inst = 32'hfe0d96a;
      58010: inst = 32'h5be00000;
      58011: inst = 32'h8c50000;
      58012: inst = 32'h24612800;
      58013: inst = 32'h10a0ffff;
      58014: inst = 32'hca0fff0;
      58015: inst = 32'h24822800;
      58016: inst = 32'h10a00000;
      58017: inst = 32'hca00004;
      58018: inst = 32'h38632800;
      58019: inst = 32'h38842800;
      58020: inst = 32'h10a00000;
      58021: inst = 32'hca0e2a9;
      58022: inst = 32'h13e00001;
      58023: inst = 32'hfe0d96a;
      58024: inst = 32'h5be00000;
      58025: inst = 32'h8c50000;
      58026: inst = 32'h24612800;
      58027: inst = 32'h10a0ffff;
      58028: inst = 32'hca0fff1;
      58029: inst = 32'h24822800;
      58030: inst = 32'h10a00000;
      58031: inst = 32'hca00004;
      58032: inst = 32'h38632800;
      58033: inst = 32'h38842800;
      58034: inst = 32'h10a00000;
      58035: inst = 32'hca0e2b7;
      58036: inst = 32'h13e00001;
      58037: inst = 32'hfe0d96a;
      58038: inst = 32'h5be00000;
      58039: inst = 32'h8c50000;
      58040: inst = 32'h24612800;
      58041: inst = 32'h10a0ffff;
      58042: inst = 32'hca0fff1;
      58043: inst = 32'h24822800;
      58044: inst = 32'h10a00000;
      58045: inst = 32'hca00004;
      58046: inst = 32'h38632800;
      58047: inst = 32'h38842800;
      58048: inst = 32'h10a00000;
      58049: inst = 32'hca0e2c5;
      58050: inst = 32'h13e00001;
      58051: inst = 32'hfe0d96a;
      58052: inst = 32'h5be00000;
      58053: inst = 32'h8c50000;
      58054: inst = 32'h24612800;
      58055: inst = 32'h10a0ffff;
      58056: inst = 32'hca0fff1;
      58057: inst = 32'h24822800;
      58058: inst = 32'h10a00000;
      58059: inst = 32'hca00004;
      58060: inst = 32'h38632800;
      58061: inst = 32'h38842800;
      58062: inst = 32'h10a00000;
      58063: inst = 32'hca0e2d3;
      58064: inst = 32'h13e00001;
      58065: inst = 32'hfe0d96a;
      58066: inst = 32'h5be00000;
      58067: inst = 32'h8c50000;
      58068: inst = 32'h24612800;
      58069: inst = 32'h10a0ffff;
      58070: inst = 32'hca0fff1;
      58071: inst = 32'h24822800;
      58072: inst = 32'h10a00000;
      58073: inst = 32'hca00004;
      58074: inst = 32'h38632800;
      58075: inst = 32'h38842800;
      58076: inst = 32'h10a00000;
      58077: inst = 32'hca0e2e1;
      58078: inst = 32'h13e00001;
      58079: inst = 32'hfe0d96a;
      58080: inst = 32'h5be00000;
      58081: inst = 32'h8c50000;
      58082: inst = 32'h24612800;
      58083: inst = 32'h10a0ffff;
      58084: inst = 32'hca0fff1;
      58085: inst = 32'h24822800;
      58086: inst = 32'h10a00000;
      58087: inst = 32'hca00004;
      58088: inst = 32'h38632800;
      58089: inst = 32'h38842800;
      58090: inst = 32'h10a00000;
      58091: inst = 32'hca0e2ef;
      58092: inst = 32'h13e00001;
      58093: inst = 32'hfe0d96a;
      58094: inst = 32'h5be00000;
      58095: inst = 32'h8c50000;
      58096: inst = 32'h24612800;
      58097: inst = 32'h10a0ffff;
      58098: inst = 32'hca0fff1;
      58099: inst = 32'h24822800;
      58100: inst = 32'h10a00000;
      58101: inst = 32'hca00004;
      58102: inst = 32'h38632800;
      58103: inst = 32'h38842800;
      58104: inst = 32'h10a00000;
      58105: inst = 32'hca0e2fd;
      58106: inst = 32'h13e00001;
      58107: inst = 32'hfe0d96a;
      58108: inst = 32'h5be00000;
      58109: inst = 32'h8c50000;
      58110: inst = 32'h24612800;
      58111: inst = 32'h10a0ffff;
      58112: inst = 32'hca0fff1;
      58113: inst = 32'h24822800;
      58114: inst = 32'h10a00000;
      58115: inst = 32'hca00004;
      58116: inst = 32'h38632800;
      58117: inst = 32'h38842800;
      58118: inst = 32'h10a00000;
      58119: inst = 32'hca0e30b;
      58120: inst = 32'h13e00001;
      58121: inst = 32'hfe0d96a;
      58122: inst = 32'h5be00000;
      58123: inst = 32'h8c50000;
      58124: inst = 32'h24612800;
      58125: inst = 32'h10a0ffff;
      58126: inst = 32'hca0fff1;
      58127: inst = 32'h24822800;
      58128: inst = 32'h10a00000;
      58129: inst = 32'hca00004;
      58130: inst = 32'h38632800;
      58131: inst = 32'h38842800;
      58132: inst = 32'h10a00000;
      58133: inst = 32'hca0e319;
      58134: inst = 32'h13e00001;
      58135: inst = 32'hfe0d96a;
      58136: inst = 32'h5be00000;
      58137: inst = 32'h8c50000;
      58138: inst = 32'h24612800;
      58139: inst = 32'h10a0ffff;
      58140: inst = 32'hca0fff1;
      58141: inst = 32'h24822800;
      58142: inst = 32'h10a00000;
      58143: inst = 32'hca00004;
      58144: inst = 32'h38632800;
      58145: inst = 32'h38842800;
      58146: inst = 32'h10a00000;
      58147: inst = 32'hca0e327;
      58148: inst = 32'h13e00001;
      58149: inst = 32'hfe0d96a;
      58150: inst = 32'h5be00000;
      58151: inst = 32'h8c50000;
      58152: inst = 32'h24612800;
      58153: inst = 32'h10a0ffff;
      58154: inst = 32'hca0fff1;
      58155: inst = 32'h24822800;
      58156: inst = 32'h10a00000;
      58157: inst = 32'hca00004;
      58158: inst = 32'h38632800;
      58159: inst = 32'h38842800;
      58160: inst = 32'h10a00000;
      58161: inst = 32'hca0e335;
      58162: inst = 32'h13e00001;
      58163: inst = 32'hfe0d96a;
      58164: inst = 32'h5be00000;
      58165: inst = 32'h8c50000;
      58166: inst = 32'h24612800;
      58167: inst = 32'h10a0ffff;
      58168: inst = 32'hca0fff1;
      58169: inst = 32'h24822800;
      58170: inst = 32'h10a00000;
      58171: inst = 32'hca00004;
      58172: inst = 32'h38632800;
      58173: inst = 32'h38842800;
      58174: inst = 32'h10a00000;
      58175: inst = 32'hca0e343;
      58176: inst = 32'h13e00001;
      58177: inst = 32'hfe0d96a;
      58178: inst = 32'h5be00000;
      58179: inst = 32'h8c50000;
      58180: inst = 32'h24612800;
      58181: inst = 32'h10a0ffff;
      58182: inst = 32'hca0fff1;
      58183: inst = 32'h24822800;
      58184: inst = 32'h10a00000;
      58185: inst = 32'hca00004;
      58186: inst = 32'h38632800;
      58187: inst = 32'h38842800;
      58188: inst = 32'h10a00000;
      58189: inst = 32'hca0e351;
      58190: inst = 32'h13e00001;
      58191: inst = 32'hfe0d96a;
      58192: inst = 32'h5be00000;
      58193: inst = 32'h8c50000;
      58194: inst = 32'h24612800;
      58195: inst = 32'h10a0ffff;
      58196: inst = 32'hca0fff1;
      58197: inst = 32'h24822800;
      58198: inst = 32'h10a00000;
      58199: inst = 32'hca00004;
      58200: inst = 32'h38632800;
      58201: inst = 32'h38842800;
      58202: inst = 32'h10a00000;
      58203: inst = 32'hca0e35f;
      58204: inst = 32'h13e00001;
      58205: inst = 32'hfe0d96a;
      58206: inst = 32'h5be00000;
      58207: inst = 32'h8c50000;
      58208: inst = 32'h24612800;
      58209: inst = 32'h10a0ffff;
      58210: inst = 32'hca0fff1;
      58211: inst = 32'h24822800;
      58212: inst = 32'h10a00000;
      58213: inst = 32'hca00004;
      58214: inst = 32'h38632800;
      58215: inst = 32'h38842800;
      58216: inst = 32'h10a00000;
      58217: inst = 32'hca0e36d;
      58218: inst = 32'h13e00001;
      58219: inst = 32'hfe0d96a;
      58220: inst = 32'h5be00000;
      58221: inst = 32'h8c50000;
      58222: inst = 32'h24612800;
      58223: inst = 32'h10a0ffff;
      58224: inst = 32'hca0fff1;
      58225: inst = 32'h24822800;
      58226: inst = 32'h10a00000;
      58227: inst = 32'hca00004;
      58228: inst = 32'h38632800;
      58229: inst = 32'h38842800;
      58230: inst = 32'h10a00000;
      58231: inst = 32'hca0e37b;
      58232: inst = 32'h13e00001;
      58233: inst = 32'hfe0d96a;
      58234: inst = 32'h5be00000;
      58235: inst = 32'h8c50000;
      58236: inst = 32'h24612800;
      58237: inst = 32'h10a0ffff;
      58238: inst = 32'hca0fff1;
      58239: inst = 32'h24822800;
      58240: inst = 32'h10a00000;
      58241: inst = 32'hca00004;
      58242: inst = 32'h38632800;
      58243: inst = 32'h38842800;
      58244: inst = 32'h10a00000;
      58245: inst = 32'hca0e389;
      58246: inst = 32'h13e00001;
      58247: inst = 32'hfe0d96a;
      58248: inst = 32'h5be00000;
      58249: inst = 32'h8c50000;
      58250: inst = 32'h24612800;
      58251: inst = 32'h10a0ffff;
      58252: inst = 32'hca0fff1;
      58253: inst = 32'h24822800;
      58254: inst = 32'h10a00000;
      58255: inst = 32'hca00004;
      58256: inst = 32'h38632800;
      58257: inst = 32'h38842800;
      58258: inst = 32'h10a00000;
      58259: inst = 32'hca0e397;
      58260: inst = 32'h13e00001;
      58261: inst = 32'hfe0d96a;
      58262: inst = 32'h5be00000;
      58263: inst = 32'h8c50000;
      58264: inst = 32'h24612800;
      58265: inst = 32'h10a0ffff;
      58266: inst = 32'hca0fff1;
      58267: inst = 32'h24822800;
      58268: inst = 32'h10a00000;
      58269: inst = 32'hca00004;
      58270: inst = 32'h38632800;
      58271: inst = 32'h38842800;
      58272: inst = 32'h10a00000;
      58273: inst = 32'hca0e3a5;
      58274: inst = 32'h13e00001;
      58275: inst = 32'hfe0d96a;
      58276: inst = 32'h5be00000;
      58277: inst = 32'h8c50000;
      58278: inst = 32'h24612800;
      58279: inst = 32'h10a0ffff;
      58280: inst = 32'hca0fff1;
      58281: inst = 32'h24822800;
      58282: inst = 32'h10a00000;
      58283: inst = 32'hca00004;
      58284: inst = 32'h38632800;
      58285: inst = 32'h38842800;
      58286: inst = 32'h10a00000;
      58287: inst = 32'hca0e3b3;
      58288: inst = 32'h13e00001;
      58289: inst = 32'hfe0d96a;
      58290: inst = 32'h5be00000;
      58291: inst = 32'h8c50000;
      58292: inst = 32'h24612800;
      58293: inst = 32'h10a0ffff;
      58294: inst = 32'hca0fff1;
      58295: inst = 32'h24822800;
      58296: inst = 32'h10a00000;
      58297: inst = 32'hca00004;
      58298: inst = 32'h38632800;
      58299: inst = 32'h38842800;
      58300: inst = 32'h10a00000;
      58301: inst = 32'hca0e3c1;
      58302: inst = 32'h13e00001;
      58303: inst = 32'hfe0d96a;
      58304: inst = 32'h5be00000;
      58305: inst = 32'h8c50000;
      58306: inst = 32'h24612800;
      58307: inst = 32'h10a0ffff;
      58308: inst = 32'hca0fff1;
      58309: inst = 32'h24822800;
      58310: inst = 32'h10a00000;
      58311: inst = 32'hca00004;
      58312: inst = 32'h38632800;
      58313: inst = 32'h38842800;
      58314: inst = 32'h10a00000;
      58315: inst = 32'hca0e3cf;
      58316: inst = 32'h13e00001;
      58317: inst = 32'hfe0d96a;
      58318: inst = 32'h5be00000;
      58319: inst = 32'h8c50000;
      58320: inst = 32'h24612800;
      58321: inst = 32'h10a0ffff;
      58322: inst = 32'hca0fff1;
      58323: inst = 32'h24822800;
      58324: inst = 32'h10a00000;
      58325: inst = 32'hca00004;
      58326: inst = 32'h38632800;
      58327: inst = 32'h38842800;
      58328: inst = 32'h10a00000;
      58329: inst = 32'hca0e3dd;
      58330: inst = 32'h13e00001;
      58331: inst = 32'hfe0d96a;
      58332: inst = 32'h5be00000;
      58333: inst = 32'h8c50000;
      58334: inst = 32'h24612800;
      58335: inst = 32'h10a0ffff;
      58336: inst = 32'hca0fff1;
      58337: inst = 32'h24822800;
      58338: inst = 32'h10a00000;
      58339: inst = 32'hca00004;
      58340: inst = 32'h38632800;
      58341: inst = 32'h38842800;
      58342: inst = 32'h10a00000;
      58343: inst = 32'hca0e3eb;
      58344: inst = 32'h13e00001;
      58345: inst = 32'hfe0d96a;
      58346: inst = 32'h5be00000;
      58347: inst = 32'h8c50000;
      58348: inst = 32'h24612800;
      58349: inst = 32'h10a0ffff;
      58350: inst = 32'hca0fff1;
      58351: inst = 32'h24822800;
      58352: inst = 32'h10a00000;
      58353: inst = 32'hca00004;
      58354: inst = 32'h38632800;
      58355: inst = 32'h38842800;
      58356: inst = 32'h10a00000;
      58357: inst = 32'hca0e3f9;
      58358: inst = 32'h13e00001;
      58359: inst = 32'hfe0d96a;
      58360: inst = 32'h5be00000;
      58361: inst = 32'h8c50000;
      58362: inst = 32'h24612800;
      58363: inst = 32'h10a0ffff;
      58364: inst = 32'hca0fff1;
      58365: inst = 32'h24822800;
      58366: inst = 32'h10a00000;
      58367: inst = 32'hca00004;
      58368: inst = 32'h38632800;
      58369: inst = 32'h38842800;
      58370: inst = 32'h10a00000;
      58371: inst = 32'hca0e407;
      58372: inst = 32'h13e00001;
      58373: inst = 32'hfe0d96a;
      58374: inst = 32'h5be00000;
      58375: inst = 32'h8c50000;
      58376: inst = 32'h24612800;
      58377: inst = 32'h10a0ffff;
      58378: inst = 32'hca0fff1;
      58379: inst = 32'h24822800;
      58380: inst = 32'h10a00000;
      58381: inst = 32'hca00004;
      58382: inst = 32'h38632800;
      58383: inst = 32'h38842800;
      58384: inst = 32'h10a00000;
      58385: inst = 32'hca0e415;
      58386: inst = 32'h13e00001;
      58387: inst = 32'hfe0d96a;
      58388: inst = 32'h5be00000;
      58389: inst = 32'h8c50000;
      58390: inst = 32'h24612800;
      58391: inst = 32'h10a0ffff;
      58392: inst = 32'hca0fff1;
      58393: inst = 32'h24822800;
      58394: inst = 32'h10a00000;
      58395: inst = 32'hca00004;
      58396: inst = 32'h38632800;
      58397: inst = 32'h38842800;
      58398: inst = 32'h10a00000;
      58399: inst = 32'hca0e423;
      58400: inst = 32'h13e00001;
      58401: inst = 32'hfe0d96a;
      58402: inst = 32'h5be00000;
      58403: inst = 32'h8c50000;
      58404: inst = 32'h24612800;
      58405: inst = 32'h10a0ffff;
      58406: inst = 32'hca0fff1;
      58407: inst = 32'h24822800;
      58408: inst = 32'h10a00000;
      58409: inst = 32'hca00004;
      58410: inst = 32'h38632800;
      58411: inst = 32'h38842800;
      58412: inst = 32'h10a00000;
      58413: inst = 32'hca0e431;
      58414: inst = 32'h13e00001;
      58415: inst = 32'hfe0d96a;
      58416: inst = 32'h5be00000;
      58417: inst = 32'h8c50000;
      58418: inst = 32'h24612800;
      58419: inst = 32'h10a0ffff;
      58420: inst = 32'hca0fff1;
      58421: inst = 32'h24822800;
      58422: inst = 32'h10a00000;
      58423: inst = 32'hca00004;
      58424: inst = 32'h38632800;
      58425: inst = 32'h38842800;
      58426: inst = 32'h10a00000;
      58427: inst = 32'hca0e43f;
      58428: inst = 32'h13e00001;
      58429: inst = 32'hfe0d96a;
      58430: inst = 32'h5be00000;
      58431: inst = 32'h8c50000;
      58432: inst = 32'h24612800;
      58433: inst = 32'h10a0ffff;
      58434: inst = 32'hca0fff1;
      58435: inst = 32'h24822800;
      58436: inst = 32'h10a00000;
      58437: inst = 32'hca00004;
      58438: inst = 32'h38632800;
      58439: inst = 32'h38842800;
      58440: inst = 32'h10a00000;
      58441: inst = 32'hca0e44d;
      58442: inst = 32'h13e00001;
      58443: inst = 32'hfe0d96a;
      58444: inst = 32'h5be00000;
      58445: inst = 32'h8c50000;
      58446: inst = 32'h24612800;
      58447: inst = 32'h10a0ffff;
      58448: inst = 32'hca0fff1;
      58449: inst = 32'h24822800;
      58450: inst = 32'h10a00000;
      58451: inst = 32'hca00004;
      58452: inst = 32'h38632800;
      58453: inst = 32'h38842800;
      58454: inst = 32'h10a00000;
      58455: inst = 32'hca0e45b;
      58456: inst = 32'h13e00001;
      58457: inst = 32'hfe0d96a;
      58458: inst = 32'h5be00000;
      58459: inst = 32'h8c50000;
      58460: inst = 32'h24612800;
      58461: inst = 32'h10a0ffff;
      58462: inst = 32'hca0fff1;
      58463: inst = 32'h24822800;
      58464: inst = 32'h10a00000;
      58465: inst = 32'hca00004;
      58466: inst = 32'h38632800;
      58467: inst = 32'h38842800;
      58468: inst = 32'h10a00000;
      58469: inst = 32'hca0e469;
      58470: inst = 32'h13e00001;
      58471: inst = 32'hfe0d96a;
      58472: inst = 32'h5be00000;
      58473: inst = 32'h8c50000;
      58474: inst = 32'h24612800;
      58475: inst = 32'h10a0ffff;
      58476: inst = 32'hca0fff1;
      58477: inst = 32'h24822800;
      58478: inst = 32'h10a00000;
      58479: inst = 32'hca00004;
      58480: inst = 32'h38632800;
      58481: inst = 32'h38842800;
      58482: inst = 32'h10a00000;
      58483: inst = 32'hca0e477;
      58484: inst = 32'h13e00001;
      58485: inst = 32'hfe0d96a;
      58486: inst = 32'h5be00000;
      58487: inst = 32'h8c50000;
      58488: inst = 32'h24612800;
      58489: inst = 32'h10a0ffff;
      58490: inst = 32'hca0fff1;
      58491: inst = 32'h24822800;
      58492: inst = 32'h10a00000;
      58493: inst = 32'hca00004;
      58494: inst = 32'h38632800;
      58495: inst = 32'h38842800;
      58496: inst = 32'h10a00000;
      58497: inst = 32'hca0e485;
      58498: inst = 32'h13e00001;
      58499: inst = 32'hfe0d96a;
      58500: inst = 32'h5be00000;
      58501: inst = 32'h8c50000;
      58502: inst = 32'h24612800;
      58503: inst = 32'h10a0ffff;
      58504: inst = 32'hca0fff1;
      58505: inst = 32'h24822800;
      58506: inst = 32'h10a00000;
      58507: inst = 32'hca00004;
      58508: inst = 32'h38632800;
      58509: inst = 32'h38842800;
      58510: inst = 32'h10a00000;
      58511: inst = 32'hca0e493;
      58512: inst = 32'h13e00001;
      58513: inst = 32'hfe0d96a;
      58514: inst = 32'h5be00000;
      58515: inst = 32'h8c50000;
      58516: inst = 32'h24612800;
      58517: inst = 32'h10a0ffff;
      58518: inst = 32'hca0fff1;
      58519: inst = 32'h24822800;
      58520: inst = 32'h10a00000;
      58521: inst = 32'hca00004;
      58522: inst = 32'h38632800;
      58523: inst = 32'h38842800;
      58524: inst = 32'h10a00000;
      58525: inst = 32'hca0e4a1;
      58526: inst = 32'h13e00001;
      58527: inst = 32'hfe0d96a;
      58528: inst = 32'h5be00000;
      58529: inst = 32'h8c50000;
      58530: inst = 32'h24612800;
      58531: inst = 32'h10a0ffff;
      58532: inst = 32'hca0fff1;
      58533: inst = 32'h24822800;
      58534: inst = 32'h10a00000;
      58535: inst = 32'hca00004;
      58536: inst = 32'h38632800;
      58537: inst = 32'h38842800;
      58538: inst = 32'h10a00000;
      58539: inst = 32'hca0e4af;
      58540: inst = 32'h13e00001;
      58541: inst = 32'hfe0d96a;
      58542: inst = 32'h5be00000;
      58543: inst = 32'h8c50000;
      58544: inst = 32'h24612800;
      58545: inst = 32'h10a0ffff;
      58546: inst = 32'hca0fff1;
      58547: inst = 32'h24822800;
      58548: inst = 32'h10a00000;
      58549: inst = 32'hca00004;
      58550: inst = 32'h38632800;
      58551: inst = 32'h38842800;
      58552: inst = 32'h10a00000;
      58553: inst = 32'hca0e4bd;
      58554: inst = 32'h13e00001;
      58555: inst = 32'hfe0d96a;
      58556: inst = 32'h5be00000;
      58557: inst = 32'h8c50000;
      58558: inst = 32'h24612800;
      58559: inst = 32'h10a0ffff;
      58560: inst = 32'hca0fff1;
      58561: inst = 32'h24822800;
      58562: inst = 32'h10a00000;
      58563: inst = 32'hca00004;
      58564: inst = 32'h38632800;
      58565: inst = 32'h38842800;
      58566: inst = 32'h10a00000;
      58567: inst = 32'hca0e4cb;
      58568: inst = 32'h13e00001;
      58569: inst = 32'hfe0d96a;
      58570: inst = 32'h5be00000;
      58571: inst = 32'h8c50000;
      58572: inst = 32'h24612800;
      58573: inst = 32'h10a0ffff;
      58574: inst = 32'hca0fff1;
      58575: inst = 32'h24822800;
      58576: inst = 32'h10a00000;
      58577: inst = 32'hca00004;
      58578: inst = 32'h38632800;
      58579: inst = 32'h38842800;
      58580: inst = 32'h10a00000;
      58581: inst = 32'hca0e4d9;
      58582: inst = 32'h13e00001;
      58583: inst = 32'hfe0d96a;
      58584: inst = 32'h5be00000;
      58585: inst = 32'h8c50000;
      58586: inst = 32'h24612800;
      58587: inst = 32'h10a0ffff;
      58588: inst = 32'hca0fff1;
      58589: inst = 32'h24822800;
      58590: inst = 32'h10a00000;
      58591: inst = 32'hca00004;
      58592: inst = 32'h38632800;
      58593: inst = 32'h38842800;
      58594: inst = 32'h10a00000;
      58595: inst = 32'hca0e4e7;
      58596: inst = 32'h13e00001;
      58597: inst = 32'hfe0d96a;
      58598: inst = 32'h5be00000;
      58599: inst = 32'h8c50000;
      58600: inst = 32'h24612800;
      58601: inst = 32'h10a0ffff;
      58602: inst = 32'hca0fff1;
      58603: inst = 32'h24822800;
      58604: inst = 32'h10a00000;
      58605: inst = 32'hca00004;
      58606: inst = 32'h38632800;
      58607: inst = 32'h38842800;
      58608: inst = 32'h10a00000;
      58609: inst = 32'hca0e4f5;
      58610: inst = 32'h13e00001;
      58611: inst = 32'hfe0d96a;
      58612: inst = 32'h5be00000;
      58613: inst = 32'h8c50000;
      58614: inst = 32'h24612800;
      58615: inst = 32'h10a0ffff;
      58616: inst = 32'hca0fff1;
      58617: inst = 32'h24822800;
      58618: inst = 32'h10a00000;
      58619: inst = 32'hca00004;
      58620: inst = 32'h38632800;
      58621: inst = 32'h38842800;
      58622: inst = 32'h10a00000;
      58623: inst = 32'hca0e503;
      58624: inst = 32'h13e00001;
      58625: inst = 32'hfe0d96a;
      58626: inst = 32'h5be00000;
      58627: inst = 32'h8c50000;
      58628: inst = 32'h24612800;
      58629: inst = 32'h10a0ffff;
      58630: inst = 32'hca0fff1;
      58631: inst = 32'h24822800;
      58632: inst = 32'h10a00000;
      58633: inst = 32'hca00004;
      58634: inst = 32'h38632800;
      58635: inst = 32'h38842800;
      58636: inst = 32'h10a00000;
      58637: inst = 32'hca0e511;
      58638: inst = 32'h13e00001;
      58639: inst = 32'hfe0d96a;
      58640: inst = 32'h5be00000;
      58641: inst = 32'h8c50000;
      58642: inst = 32'h24612800;
      58643: inst = 32'h10a0ffff;
      58644: inst = 32'hca0fff1;
      58645: inst = 32'h24822800;
      58646: inst = 32'h10a00000;
      58647: inst = 32'hca00004;
      58648: inst = 32'h38632800;
      58649: inst = 32'h38842800;
      58650: inst = 32'h10a00000;
      58651: inst = 32'hca0e51f;
      58652: inst = 32'h13e00001;
      58653: inst = 32'hfe0d96a;
      58654: inst = 32'h5be00000;
      58655: inst = 32'h8c50000;
      58656: inst = 32'h24612800;
      58657: inst = 32'h10a0ffff;
      58658: inst = 32'hca0fff1;
      58659: inst = 32'h24822800;
      58660: inst = 32'h10a00000;
      58661: inst = 32'hca00004;
      58662: inst = 32'h38632800;
      58663: inst = 32'h38842800;
      58664: inst = 32'h10a00000;
      58665: inst = 32'hca0e52d;
      58666: inst = 32'h13e00001;
      58667: inst = 32'hfe0d96a;
      58668: inst = 32'h5be00000;
      58669: inst = 32'h8c50000;
      58670: inst = 32'h24612800;
      58671: inst = 32'h10a0ffff;
      58672: inst = 32'hca0fff1;
      58673: inst = 32'h24822800;
      58674: inst = 32'h10a00000;
      58675: inst = 32'hca00004;
      58676: inst = 32'h38632800;
      58677: inst = 32'h38842800;
      58678: inst = 32'h10a00000;
      58679: inst = 32'hca0e53b;
      58680: inst = 32'h13e00001;
      58681: inst = 32'hfe0d96a;
      58682: inst = 32'h5be00000;
      58683: inst = 32'h8c50000;
      58684: inst = 32'h24612800;
      58685: inst = 32'h10a0ffff;
      58686: inst = 32'hca0fff1;
      58687: inst = 32'h24822800;
      58688: inst = 32'h10a00000;
      58689: inst = 32'hca00004;
      58690: inst = 32'h38632800;
      58691: inst = 32'h38842800;
      58692: inst = 32'h10a00000;
      58693: inst = 32'hca0e549;
      58694: inst = 32'h13e00001;
      58695: inst = 32'hfe0d96a;
      58696: inst = 32'h5be00000;
      58697: inst = 32'h8c50000;
      58698: inst = 32'h24612800;
      58699: inst = 32'h10a0ffff;
      58700: inst = 32'hca0fff1;
      58701: inst = 32'h24822800;
      58702: inst = 32'h10a00000;
      58703: inst = 32'hca00004;
      58704: inst = 32'h38632800;
      58705: inst = 32'h38842800;
      58706: inst = 32'h10a00000;
      58707: inst = 32'hca0e557;
      58708: inst = 32'h13e00001;
      58709: inst = 32'hfe0d96a;
      58710: inst = 32'h5be00000;
      58711: inst = 32'h8c50000;
      58712: inst = 32'h24612800;
      58713: inst = 32'h10a0ffff;
      58714: inst = 32'hca0fff1;
      58715: inst = 32'h24822800;
      58716: inst = 32'h10a00000;
      58717: inst = 32'hca00004;
      58718: inst = 32'h38632800;
      58719: inst = 32'h38842800;
      58720: inst = 32'h10a00000;
      58721: inst = 32'hca0e565;
      58722: inst = 32'h13e00001;
      58723: inst = 32'hfe0d96a;
      58724: inst = 32'h5be00000;
      58725: inst = 32'h8c50000;
      58726: inst = 32'h24612800;
      58727: inst = 32'h10a0ffff;
      58728: inst = 32'hca0fff1;
      58729: inst = 32'h24822800;
      58730: inst = 32'h10a00000;
      58731: inst = 32'hca00004;
      58732: inst = 32'h38632800;
      58733: inst = 32'h38842800;
      58734: inst = 32'h10a00000;
      58735: inst = 32'hca0e573;
      58736: inst = 32'h13e00001;
      58737: inst = 32'hfe0d96a;
      58738: inst = 32'h5be00000;
      58739: inst = 32'h8c50000;
      58740: inst = 32'h24612800;
      58741: inst = 32'h10a0ffff;
      58742: inst = 32'hca0fff1;
      58743: inst = 32'h24822800;
      58744: inst = 32'h10a00000;
      58745: inst = 32'hca00004;
      58746: inst = 32'h38632800;
      58747: inst = 32'h38842800;
      58748: inst = 32'h10a00000;
      58749: inst = 32'hca0e581;
      58750: inst = 32'h13e00001;
      58751: inst = 32'hfe0d96a;
      58752: inst = 32'h5be00000;
      58753: inst = 32'h8c50000;
      58754: inst = 32'h24612800;
      58755: inst = 32'h10a0ffff;
      58756: inst = 32'hca0fff1;
      58757: inst = 32'h24822800;
      58758: inst = 32'h10a00000;
      58759: inst = 32'hca00004;
      58760: inst = 32'h38632800;
      58761: inst = 32'h38842800;
      58762: inst = 32'h10a00000;
      58763: inst = 32'hca0e58f;
      58764: inst = 32'h13e00001;
      58765: inst = 32'hfe0d96a;
      58766: inst = 32'h5be00000;
      58767: inst = 32'h8c50000;
      58768: inst = 32'h24612800;
      58769: inst = 32'h10a0ffff;
      58770: inst = 32'hca0fff1;
      58771: inst = 32'h24822800;
      58772: inst = 32'h10a00000;
      58773: inst = 32'hca00004;
      58774: inst = 32'h38632800;
      58775: inst = 32'h38842800;
      58776: inst = 32'h10a00000;
      58777: inst = 32'hca0e59d;
      58778: inst = 32'h13e00001;
      58779: inst = 32'hfe0d96a;
      58780: inst = 32'h5be00000;
      58781: inst = 32'h8c50000;
      58782: inst = 32'h24612800;
      58783: inst = 32'h10a0ffff;
      58784: inst = 32'hca0fff1;
      58785: inst = 32'h24822800;
      58786: inst = 32'h10a00000;
      58787: inst = 32'hca00004;
      58788: inst = 32'h38632800;
      58789: inst = 32'h38842800;
      58790: inst = 32'h10a00000;
      58791: inst = 32'hca0e5ab;
      58792: inst = 32'h13e00001;
      58793: inst = 32'hfe0d96a;
      58794: inst = 32'h5be00000;
      58795: inst = 32'h8c50000;
      58796: inst = 32'h24612800;
      58797: inst = 32'h10a0ffff;
      58798: inst = 32'hca0fff1;
      58799: inst = 32'h24822800;
      58800: inst = 32'h10a00000;
      58801: inst = 32'hca00004;
      58802: inst = 32'h38632800;
      58803: inst = 32'h38842800;
      58804: inst = 32'h10a00000;
      58805: inst = 32'hca0e5b9;
      58806: inst = 32'h13e00001;
      58807: inst = 32'hfe0d96a;
      58808: inst = 32'h5be00000;
      58809: inst = 32'h8c50000;
      58810: inst = 32'h24612800;
      58811: inst = 32'h10a0ffff;
      58812: inst = 32'hca0fff1;
      58813: inst = 32'h24822800;
      58814: inst = 32'h10a00000;
      58815: inst = 32'hca00004;
      58816: inst = 32'h38632800;
      58817: inst = 32'h38842800;
      58818: inst = 32'h10a00000;
      58819: inst = 32'hca0e5c7;
      58820: inst = 32'h13e00001;
      58821: inst = 32'hfe0d96a;
      58822: inst = 32'h5be00000;
      58823: inst = 32'h8c50000;
      58824: inst = 32'h24612800;
      58825: inst = 32'h10a0ffff;
      58826: inst = 32'hca0fff1;
      58827: inst = 32'h24822800;
      58828: inst = 32'h10a00000;
      58829: inst = 32'hca00004;
      58830: inst = 32'h38632800;
      58831: inst = 32'h38842800;
      58832: inst = 32'h10a00000;
      58833: inst = 32'hca0e5d5;
      58834: inst = 32'h13e00001;
      58835: inst = 32'hfe0d96a;
      58836: inst = 32'h5be00000;
      58837: inst = 32'h8c50000;
      58838: inst = 32'h24612800;
      58839: inst = 32'h10a0ffff;
      58840: inst = 32'hca0fff1;
      58841: inst = 32'h24822800;
      58842: inst = 32'h10a00000;
      58843: inst = 32'hca00004;
      58844: inst = 32'h38632800;
      58845: inst = 32'h38842800;
      58846: inst = 32'h10a00000;
      58847: inst = 32'hca0e5e3;
      58848: inst = 32'h13e00001;
      58849: inst = 32'hfe0d96a;
      58850: inst = 32'h5be00000;
      58851: inst = 32'h8c50000;
      58852: inst = 32'h24612800;
      58853: inst = 32'h10a0ffff;
      58854: inst = 32'hca0fff1;
      58855: inst = 32'h24822800;
      58856: inst = 32'h10a00000;
      58857: inst = 32'hca00004;
      58858: inst = 32'h38632800;
      58859: inst = 32'h38842800;
      58860: inst = 32'h10a00000;
      58861: inst = 32'hca0e5f1;
      58862: inst = 32'h13e00001;
      58863: inst = 32'hfe0d96a;
      58864: inst = 32'h5be00000;
      58865: inst = 32'h8c50000;
      58866: inst = 32'h24612800;
      58867: inst = 32'h10a0ffff;
      58868: inst = 32'hca0fff1;
      58869: inst = 32'h24822800;
      58870: inst = 32'h10a00000;
      58871: inst = 32'hca00004;
      58872: inst = 32'h38632800;
      58873: inst = 32'h38842800;
      58874: inst = 32'h10a00000;
      58875: inst = 32'hca0e5ff;
      58876: inst = 32'h13e00001;
      58877: inst = 32'hfe0d96a;
      58878: inst = 32'h5be00000;
      58879: inst = 32'h8c50000;
      58880: inst = 32'h24612800;
      58881: inst = 32'h10a0ffff;
      58882: inst = 32'hca0fff1;
      58883: inst = 32'h24822800;
      58884: inst = 32'h10a00000;
      58885: inst = 32'hca00004;
      58886: inst = 32'h38632800;
      58887: inst = 32'h38842800;
      58888: inst = 32'h10a00000;
      58889: inst = 32'hca0e60d;
      58890: inst = 32'h13e00001;
      58891: inst = 32'hfe0d96a;
      58892: inst = 32'h5be00000;
      58893: inst = 32'h8c50000;
      58894: inst = 32'h24612800;
      58895: inst = 32'h10a0ffff;
      58896: inst = 32'hca0fff1;
      58897: inst = 32'h24822800;
      58898: inst = 32'h10a00000;
      58899: inst = 32'hca00004;
      58900: inst = 32'h38632800;
      58901: inst = 32'h38842800;
      58902: inst = 32'h10a00000;
      58903: inst = 32'hca0e61b;
      58904: inst = 32'h13e00001;
      58905: inst = 32'hfe0d96a;
      58906: inst = 32'h5be00000;
      58907: inst = 32'h8c50000;
      58908: inst = 32'h24612800;
      58909: inst = 32'h10a0ffff;
      58910: inst = 32'hca0fff1;
      58911: inst = 32'h24822800;
      58912: inst = 32'h10a00000;
      58913: inst = 32'hca00004;
      58914: inst = 32'h38632800;
      58915: inst = 32'h38842800;
      58916: inst = 32'h10a00000;
      58917: inst = 32'hca0e629;
      58918: inst = 32'h13e00001;
      58919: inst = 32'hfe0d96a;
      58920: inst = 32'h5be00000;
      58921: inst = 32'h8c50000;
      58922: inst = 32'h24612800;
      58923: inst = 32'h10a0ffff;
      58924: inst = 32'hca0fff1;
      58925: inst = 32'h24822800;
      58926: inst = 32'h10a00000;
      58927: inst = 32'hca00004;
      58928: inst = 32'h38632800;
      58929: inst = 32'h38842800;
      58930: inst = 32'h10a00000;
      58931: inst = 32'hca0e637;
      58932: inst = 32'h13e00001;
      58933: inst = 32'hfe0d96a;
      58934: inst = 32'h5be00000;
      58935: inst = 32'h8c50000;
      58936: inst = 32'h24612800;
      58937: inst = 32'h10a0ffff;
      58938: inst = 32'hca0fff1;
      58939: inst = 32'h24822800;
      58940: inst = 32'h10a00000;
      58941: inst = 32'hca00004;
      58942: inst = 32'h38632800;
      58943: inst = 32'h38842800;
      58944: inst = 32'h10a00000;
      58945: inst = 32'hca0e645;
      58946: inst = 32'h13e00001;
      58947: inst = 32'hfe0d96a;
      58948: inst = 32'h5be00000;
      58949: inst = 32'h8c50000;
      58950: inst = 32'h24612800;
      58951: inst = 32'h10a0ffff;
      58952: inst = 32'hca0fff1;
      58953: inst = 32'h24822800;
      58954: inst = 32'h10a00000;
      58955: inst = 32'hca00004;
      58956: inst = 32'h38632800;
      58957: inst = 32'h38842800;
      58958: inst = 32'h10a00000;
      58959: inst = 32'hca0e653;
      58960: inst = 32'h13e00001;
      58961: inst = 32'hfe0d96a;
      58962: inst = 32'h5be00000;
      58963: inst = 32'h8c50000;
      58964: inst = 32'h24612800;
      58965: inst = 32'h10a0ffff;
      58966: inst = 32'hca0fff1;
      58967: inst = 32'h24822800;
      58968: inst = 32'h10a00000;
      58969: inst = 32'hca00004;
      58970: inst = 32'h38632800;
      58971: inst = 32'h38842800;
      58972: inst = 32'h10a00000;
      58973: inst = 32'hca0e661;
      58974: inst = 32'h13e00001;
      58975: inst = 32'hfe0d96a;
      58976: inst = 32'h5be00000;
      58977: inst = 32'h8c50000;
      58978: inst = 32'h24612800;
      58979: inst = 32'h10a0ffff;
      58980: inst = 32'hca0fff1;
      58981: inst = 32'h24822800;
      58982: inst = 32'h10a00000;
      58983: inst = 32'hca00004;
      58984: inst = 32'h38632800;
      58985: inst = 32'h38842800;
      58986: inst = 32'h10a00000;
      58987: inst = 32'hca0e66f;
      58988: inst = 32'h13e00001;
      58989: inst = 32'hfe0d96a;
      58990: inst = 32'h5be00000;
      58991: inst = 32'h8c50000;
      58992: inst = 32'h24612800;
      58993: inst = 32'h10a0ffff;
      58994: inst = 32'hca0fff1;
      58995: inst = 32'h24822800;
      58996: inst = 32'h10a00000;
      58997: inst = 32'hca00004;
      58998: inst = 32'h38632800;
      58999: inst = 32'h38842800;
      59000: inst = 32'h10a00000;
      59001: inst = 32'hca0e67d;
      59002: inst = 32'h13e00001;
      59003: inst = 32'hfe0d96a;
      59004: inst = 32'h5be00000;
      59005: inst = 32'h8c50000;
      59006: inst = 32'h24612800;
      59007: inst = 32'h10a0ffff;
      59008: inst = 32'hca0fff1;
      59009: inst = 32'h24822800;
      59010: inst = 32'h10a00000;
      59011: inst = 32'hca00004;
      59012: inst = 32'h38632800;
      59013: inst = 32'h38842800;
      59014: inst = 32'h10a00000;
      59015: inst = 32'hca0e68b;
      59016: inst = 32'h13e00001;
      59017: inst = 32'hfe0d96a;
      59018: inst = 32'h5be00000;
      59019: inst = 32'h8c50000;
      59020: inst = 32'h24612800;
      59021: inst = 32'h10a0ffff;
      59022: inst = 32'hca0fff1;
      59023: inst = 32'h24822800;
      59024: inst = 32'h10a00000;
      59025: inst = 32'hca00004;
      59026: inst = 32'h38632800;
      59027: inst = 32'h38842800;
      59028: inst = 32'h10a00000;
      59029: inst = 32'hca0e699;
      59030: inst = 32'h13e00001;
      59031: inst = 32'hfe0d96a;
      59032: inst = 32'h5be00000;
      59033: inst = 32'h8c50000;
      59034: inst = 32'h24612800;
      59035: inst = 32'h10a0ffff;
      59036: inst = 32'hca0fff1;
      59037: inst = 32'h24822800;
      59038: inst = 32'h10a00000;
      59039: inst = 32'hca00004;
      59040: inst = 32'h38632800;
      59041: inst = 32'h38842800;
      59042: inst = 32'h10a00000;
      59043: inst = 32'hca0e6a7;
      59044: inst = 32'h13e00001;
      59045: inst = 32'hfe0d96a;
      59046: inst = 32'h5be00000;
      59047: inst = 32'h8c50000;
      59048: inst = 32'h24612800;
      59049: inst = 32'h10a0ffff;
      59050: inst = 32'hca0fff1;
      59051: inst = 32'h24822800;
      59052: inst = 32'h10a00000;
      59053: inst = 32'hca00004;
      59054: inst = 32'h38632800;
      59055: inst = 32'h38842800;
      59056: inst = 32'h10a00000;
      59057: inst = 32'hca0e6b5;
      59058: inst = 32'h13e00001;
      59059: inst = 32'hfe0d96a;
      59060: inst = 32'h5be00000;
      59061: inst = 32'h8c50000;
      59062: inst = 32'h24612800;
      59063: inst = 32'h10a0ffff;
      59064: inst = 32'hca0fff1;
      59065: inst = 32'h24822800;
      59066: inst = 32'h10a00000;
      59067: inst = 32'hca00004;
      59068: inst = 32'h38632800;
      59069: inst = 32'h38842800;
      59070: inst = 32'h10a00000;
      59071: inst = 32'hca0e6c3;
      59072: inst = 32'h13e00001;
      59073: inst = 32'hfe0d96a;
      59074: inst = 32'h5be00000;
      59075: inst = 32'h8c50000;
      59076: inst = 32'h24612800;
      59077: inst = 32'h10a0ffff;
      59078: inst = 32'hca0fff1;
      59079: inst = 32'h24822800;
      59080: inst = 32'h10a00000;
      59081: inst = 32'hca00004;
      59082: inst = 32'h38632800;
      59083: inst = 32'h38842800;
      59084: inst = 32'h10a00000;
      59085: inst = 32'hca0e6d1;
      59086: inst = 32'h13e00001;
      59087: inst = 32'hfe0d96a;
      59088: inst = 32'h5be00000;
      59089: inst = 32'h8c50000;
      59090: inst = 32'h24612800;
      59091: inst = 32'h10a0ffff;
      59092: inst = 32'hca0fff1;
      59093: inst = 32'h24822800;
      59094: inst = 32'h10a00000;
      59095: inst = 32'hca00004;
      59096: inst = 32'h38632800;
      59097: inst = 32'h38842800;
      59098: inst = 32'h10a00000;
      59099: inst = 32'hca0e6df;
      59100: inst = 32'h13e00001;
      59101: inst = 32'hfe0d96a;
      59102: inst = 32'h5be00000;
      59103: inst = 32'h8c50000;
      59104: inst = 32'h24612800;
      59105: inst = 32'h10a0ffff;
      59106: inst = 32'hca0fff1;
      59107: inst = 32'h24822800;
      59108: inst = 32'h10a00000;
      59109: inst = 32'hca00004;
      59110: inst = 32'h38632800;
      59111: inst = 32'h38842800;
      59112: inst = 32'h10a00000;
      59113: inst = 32'hca0e6ed;
      59114: inst = 32'h13e00001;
      59115: inst = 32'hfe0d96a;
      59116: inst = 32'h5be00000;
      59117: inst = 32'h8c50000;
      59118: inst = 32'h24612800;
      59119: inst = 32'h10a0ffff;
      59120: inst = 32'hca0fff1;
      59121: inst = 32'h24822800;
      59122: inst = 32'h10a00000;
      59123: inst = 32'hca00004;
      59124: inst = 32'h38632800;
      59125: inst = 32'h38842800;
      59126: inst = 32'h10a00000;
      59127: inst = 32'hca0e6fb;
      59128: inst = 32'h13e00001;
      59129: inst = 32'hfe0d96a;
      59130: inst = 32'h5be00000;
      59131: inst = 32'h8c50000;
      59132: inst = 32'h24612800;
      59133: inst = 32'h10a0ffff;
      59134: inst = 32'hca0fff1;
      59135: inst = 32'h24822800;
      59136: inst = 32'h10a00000;
      59137: inst = 32'hca00004;
      59138: inst = 32'h38632800;
      59139: inst = 32'h38842800;
      59140: inst = 32'h10a00000;
      59141: inst = 32'hca0e709;
      59142: inst = 32'h13e00001;
      59143: inst = 32'hfe0d96a;
      59144: inst = 32'h5be00000;
      59145: inst = 32'h8c50000;
      59146: inst = 32'h24612800;
      59147: inst = 32'h10a0ffff;
      59148: inst = 32'hca0fff1;
      59149: inst = 32'h24822800;
      59150: inst = 32'h10a00000;
      59151: inst = 32'hca00004;
      59152: inst = 32'h38632800;
      59153: inst = 32'h38842800;
      59154: inst = 32'h10a00000;
      59155: inst = 32'hca0e717;
      59156: inst = 32'h13e00001;
      59157: inst = 32'hfe0d96a;
      59158: inst = 32'h5be00000;
      59159: inst = 32'h8c50000;
      59160: inst = 32'h24612800;
      59161: inst = 32'h10a0ffff;
      59162: inst = 32'hca0fff1;
      59163: inst = 32'h24822800;
      59164: inst = 32'h10a00000;
      59165: inst = 32'hca00004;
      59166: inst = 32'h38632800;
      59167: inst = 32'h38842800;
      59168: inst = 32'h10a00000;
      59169: inst = 32'hca0e725;
      59170: inst = 32'h13e00001;
      59171: inst = 32'hfe0d96a;
      59172: inst = 32'h5be00000;
      59173: inst = 32'h8c50000;
      59174: inst = 32'h24612800;
      59175: inst = 32'h10a0ffff;
      59176: inst = 32'hca0fff1;
      59177: inst = 32'h24822800;
      59178: inst = 32'h10a00000;
      59179: inst = 32'hca00004;
      59180: inst = 32'h38632800;
      59181: inst = 32'h38842800;
      59182: inst = 32'h10a00000;
      59183: inst = 32'hca0e733;
      59184: inst = 32'h13e00001;
      59185: inst = 32'hfe0d96a;
      59186: inst = 32'h5be00000;
      59187: inst = 32'h8c50000;
      59188: inst = 32'h24612800;
      59189: inst = 32'h10a0ffff;
      59190: inst = 32'hca0fff1;
      59191: inst = 32'h24822800;
      59192: inst = 32'h10a00000;
      59193: inst = 32'hca00004;
      59194: inst = 32'h38632800;
      59195: inst = 32'h38842800;
      59196: inst = 32'h10a00000;
      59197: inst = 32'hca0e741;
      59198: inst = 32'h13e00001;
      59199: inst = 32'hfe0d96a;
      59200: inst = 32'h5be00000;
      59201: inst = 32'h8c50000;
      59202: inst = 32'h24612800;
      59203: inst = 32'h10a0ffff;
      59204: inst = 32'hca0fff1;
      59205: inst = 32'h24822800;
      59206: inst = 32'h10a00000;
      59207: inst = 32'hca00004;
      59208: inst = 32'h38632800;
      59209: inst = 32'h38842800;
      59210: inst = 32'h10a00000;
      59211: inst = 32'hca0e74f;
      59212: inst = 32'h13e00001;
      59213: inst = 32'hfe0d96a;
      59214: inst = 32'h5be00000;
      59215: inst = 32'h8c50000;
      59216: inst = 32'h24612800;
      59217: inst = 32'h10a0ffff;
      59218: inst = 32'hca0fff1;
      59219: inst = 32'h24822800;
      59220: inst = 32'h10a00000;
      59221: inst = 32'hca00004;
      59222: inst = 32'h38632800;
      59223: inst = 32'h38842800;
      59224: inst = 32'h10a00000;
      59225: inst = 32'hca0e75d;
      59226: inst = 32'h13e00001;
      59227: inst = 32'hfe0d96a;
      59228: inst = 32'h5be00000;
      59229: inst = 32'h8c50000;
      59230: inst = 32'h24612800;
      59231: inst = 32'h10a0ffff;
      59232: inst = 32'hca0fff1;
      59233: inst = 32'h24822800;
      59234: inst = 32'h10a00000;
      59235: inst = 32'hca00004;
      59236: inst = 32'h38632800;
      59237: inst = 32'h38842800;
      59238: inst = 32'h10a00000;
      59239: inst = 32'hca0e76b;
      59240: inst = 32'h13e00001;
      59241: inst = 32'hfe0d96a;
      59242: inst = 32'h5be00000;
      59243: inst = 32'h8c50000;
      59244: inst = 32'h24612800;
      59245: inst = 32'h10a0ffff;
      59246: inst = 32'hca0fff1;
      59247: inst = 32'h24822800;
      59248: inst = 32'h10a00000;
      59249: inst = 32'hca00004;
      59250: inst = 32'h38632800;
      59251: inst = 32'h38842800;
      59252: inst = 32'h10a00000;
      59253: inst = 32'hca0e779;
      59254: inst = 32'h13e00001;
      59255: inst = 32'hfe0d96a;
      59256: inst = 32'h5be00000;
      59257: inst = 32'h8c50000;
      59258: inst = 32'h24612800;
      59259: inst = 32'h10a0ffff;
      59260: inst = 32'hca0fff1;
      59261: inst = 32'h24822800;
      59262: inst = 32'h10a00000;
      59263: inst = 32'hca00004;
      59264: inst = 32'h38632800;
      59265: inst = 32'h38842800;
      59266: inst = 32'h10a00000;
      59267: inst = 32'hca0e787;
      59268: inst = 32'h13e00001;
      59269: inst = 32'hfe0d96a;
      59270: inst = 32'h5be00000;
      59271: inst = 32'h8c50000;
      59272: inst = 32'h24612800;
      59273: inst = 32'h10a0ffff;
      59274: inst = 32'hca0fff1;
      59275: inst = 32'h24822800;
      59276: inst = 32'h10a00000;
      59277: inst = 32'hca00004;
      59278: inst = 32'h38632800;
      59279: inst = 32'h38842800;
      59280: inst = 32'h10a00000;
      59281: inst = 32'hca0e795;
      59282: inst = 32'h13e00001;
      59283: inst = 32'hfe0d96a;
      59284: inst = 32'h5be00000;
      59285: inst = 32'h8c50000;
      59286: inst = 32'h24612800;
      59287: inst = 32'h10a0ffff;
      59288: inst = 32'hca0fff1;
      59289: inst = 32'h24822800;
      59290: inst = 32'h10a00000;
      59291: inst = 32'hca00004;
      59292: inst = 32'h38632800;
      59293: inst = 32'h38842800;
      59294: inst = 32'h10a00000;
      59295: inst = 32'hca0e7a3;
      59296: inst = 32'h13e00001;
      59297: inst = 32'hfe0d96a;
      59298: inst = 32'h5be00000;
      59299: inst = 32'h8c50000;
      59300: inst = 32'h24612800;
      59301: inst = 32'h10a0ffff;
      59302: inst = 32'hca0fff1;
      59303: inst = 32'h24822800;
      59304: inst = 32'h10a00000;
      59305: inst = 32'hca00004;
      59306: inst = 32'h38632800;
      59307: inst = 32'h38842800;
      59308: inst = 32'h10a00000;
      59309: inst = 32'hca0e7b1;
      59310: inst = 32'h13e00001;
      59311: inst = 32'hfe0d96a;
      59312: inst = 32'h5be00000;
      59313: inst = 32'h8c50000;
      59314: inst = 32'h24612800;
      59315: inst = 32'h10a0ffff;
      59316: inst = 32'hca0fff1;
      59317: inst = 32'h24822800;
      59318: inst = 32'h10a00000;
      59319: inst = 32'hca00004;
      59320: inst = 32'h38632800;
      59321: inst = 32'h38842800;
      59322: inst = 32'h10a00000;
      59323: inst = 32'hca0e7bf;
      59324: inst = 32'h13e00001;
      59325: inst = 32'hfe0d96a;
      59326: inst = 32'h5be00000;
      59327: inst = 32'h8c50000;
      59328: inst = 32'h24612800;
      59329: inst = 32'h10a0ffff;
      59330: inst = 32'hca0fff1;
      59331: inst = 32'h24822800;
      59332: inst = 32'h10a00000;
      59333: inst = 32'hca00004;
      59334: inst = 32'h38632800;
      59335: inst = 32'h38842800;
      59336: inst = 32'h10a00000;
      59337: inst = 32'hca0e7cd;
      59338: inst = 32'h13e00001;
      59339: inst = 32'hfe0d96a;
      59340: inst = 32'h5be00000;
      59341: inst = 32'h8c50000;
      59342: inst = 32'h24612800;
      59343: inst = 32'h10a0ffff;
      59344: inst = 32'hca0fff1;
      59345: inst = 32'h24822800;
      59346: inst = 32'h10a00000;
      59347: inst = 32'hca00004;
      59348: inst = 32'h38632800;
      59349: inst = 32'h38842800;
      59350: inst = 32'h10a00000;
      59351: inst = 32'hca0e7db;
      59352: inst = 32'h13e00001;
      59353: inst = 32'hfe0d96a;
      59354: inst = 32'h5be00000;
      59355: inst = 32'h8c50000;
      59356: inst = 32'h24612800;
      59357: inst = 32'h10a0ffff;
      59358: inst = 32'hca0fff1;
      59359: inst = 32'h24822800;
      59360: inst = 32'h10a00000;
      59361: inst = 32'hca00004;
      59362: inst = 32'h38632800;
      59363: inst = 32'h38842800;
      59364: inst = 32'h10a00000;
      59365: inst = 32'hca0e7e9;
      59366: inst = 32'h13e00001;
      59367: inst = 32'hfe0d96a;
      59368: inst = 32'h5be00000;
      59369: inst = 32'h8c50000;
      59370: inst = 32'h24612800;
      59371: inst = 32'h10a0ffff;
      59372: inst = 32'hca0fff2;
      59373: inst = 32'h24822800;
      59374: inst = 32'h10a00000;
      59375: inst = 32'hca00004;
      59376: inst = 32'h38632800;
      59377: inst = 32'h38842800;
      59378: inst = 32'h10a00000;
      59379: inst = 32'hca0e7f7;
      59380: inst = 32'h13e00001;
      59381: inst = 32'hfe0d96a;
      59382: inst = 32'h5be00000;
      59383: inst = 32'h8c50000;
      59384: inst = 32'h24612800;
      59385: inst = 32'h10a0ffff;
      59386: inst = 32'hca0fff2;
      59387: inst = 32'h24822800;
      59388: inst = 32'h10a00000;
      59389: inst = 32'hca00004;
      59390: inst = 32'h38632800;
      59391: inst = 32'h38842800;
      59392: inst = 32'h10a00000;
      59393: inst = 32'hca0e805;
      59394: inst = 32'h13e00001;
      59395: inst = 32'hfe0d96a;
      59396: inst = 32'h5be00000;
      59397: inst = 32'h8c50000;
      59398: inst = 32'h24612800;
      59399: inst = 32'h10a0ffff;
      59400: inst = 32'hca0fff2;
      59401: inst = 32'h24822800;
      59402: inst = 32'h10a00000;
      59403: inst = 32'hca00004;
      59404: inst = 32'h38632800;
      59405: inst = 32'h38842800;
      59406: inst = 32'h10a00000;
      59407: inst = 32'hca0e813;
      59408: inst = 32'h13e00001;
      59409: inst = 32'hfe0d96a;
      59410: inst = 32'h5be00000;
      59411: inst = 32'h8c50000;
      59412: inst = 32'h24612800;
      59413: inst = 32'h10a0ffff;
      59414: inst = 32'hca0fff2;
      59415: inst = 32'h24822800;
      59416: inst = 32'h10a00000;
      59417: inst = 32'hca00004;
      59418: inst = 32'h38632800;
      59419: inst = 32'h38842800;
      59420: inst = 32'h10a00000;
      59421: inst = 32'hca0e821;
      59422: inst = 32'h13e00001;
      59423: inst = 32'hfe0d96a;
      59424: inst = 32'h5be00000;
      59425: inst = 32'h8c50000;
      59426: inst = 32'h24612800;
      59427: inst = 32'h10a0ffff;
      59428: inst = 32'hca0fff2;
      59429: inst = 32'h24822800;
      59430: inst = 32'h10a00000;
      59431: inst = 32'hca00004;
      59432: inst = 32'h38632800;
      59433: inst = 32'h38842800;
      59434: inst = 32'h10a00000;
      59435: inst = 32'hca0e82f;
      59436: inst = 32'h13e00001;
      59437: inst = 32'hfe0d96a;
      59438: inst = 32'h5be00000;
      59439: inst = 32'h8c50000;
      59440: inst = 32'h24612800;
      59441: inst = 32'h10a0ffff;
      59442: inst = 32'hca0fff2;
      59443: inst = 32'h24822800;
      59444: inst = 32'h10a00000;
      59445: inst = 32'hca00004;
      59446: inst = 32'h38632800;
      59447: inst = 32'h38842800;
      59448: inst = 32'h10a00000;
      59449: inst = 32'hca0e83d;
      59450: inst = 32'h13e00001;
      59451: inst = 32'hfe0d96a;
      59452: inst = 32'h5be00000;
      59453: inst = 32'h8c50000;
      59454: inst = 32'h24612800;
      59455: inst = 32'h10a0ffff;
      59456: inst = 32'hca0fff2;
      59457: inst = 32'h24822800;
      59458: inst = 32'h10a00000;
      59459: inst = 32'hca00004;
      59460: inst = 32'h38632800;
      59461: inst = 32'h38842800;
      59462: inst = 32'h10a00000;
      59463: inst = 32'hca0e84b;
      59464: inst = 32'h13e00001;
      59465: inst = 32'hfe0d96a;
      59466: inst = 32'h5be00000;
      59467: inst = 32'h8c50000;
      59468: inst = 32'h24612800;
      59469: inst = 32'h10a0ffff;
      59470: inst = 32'hca0fff2;
      59471: inst = 32'h24822800;
      59472: inst = 32'h10a00000;
      59473: inst = 32'hca00004;
      59474: inst = 32'h38632800;
      59475: inst = 32'h38842800;
      59476: inst = 32'h10a00000;
      59477: inst = 32'hca0e859;
      59478: inst = 32'h13e00001;
      59479: inst = 32'hfe0d96a;
      59480: inst = 32'h5be00000;
      59481: inst = 32'h8c50000;
      59482: inst = 32'h24612800;
      59483: inst = 32'h10a0ffff;
      59484: inst = 32'hca0fff2;
      59485: inst = 32'h24822800;
      59486: inst = 32'h10a00000;
      59487: inst = 32'hca00004;
      59488: inst = 32'h38632800;
      59489: inst = 32'h38842800;
      59490: inst = 32'h10a00000;
      59491: inst = 32'hca0e867;
      59492: inst = 32'h13e00001;
      59493: inst = 32'hfe0d96a;
      59494: inst = 32'h5be00000;
      59495: inst = 32'h8c50000;
      59496: inst = 32'h24612800;
      59497: inst = 32'h10a0ffff;
      59498: inst = 32'hca0fff2;
      59499: inst = 32'h24822800;
      59500: inst = 32'h10a00000;
      59501: inst = 32'hca00004;
      59502: inst = 32'h38632800;
      59503: inst = 32'h38842800;
      59504: inst = 32'h10a00000;
      59505: inst = 32'hca0e875;
      59506: inst = 32'h13e00001;
      59507: inst = 32'hfe0d96a;
      59508: inst = 32'h5be00000;
      59509: inst = 32'h8c50000;
      59510: inst = 32'h24612800;
      59511: inst = 32'h10a0ffff;
      59512: inst = 32'hca0fff2;
      59513: inst = 32'h24822800;
      59514: inst = 32'h10a00000;
      59515: inst = 32'hca00004;
      59516: inst = 32'h38632800;
      59517: inst = 32'h38842800;
      59518: inst = 32'h10a00000;
      59519: inst = 32'hca0e883;
      59520: inst = 32'h13e00001;
      59521: inst = 32'hfe0d96a;
      59522: inst = 32'h5be00000;
      59523: inst = 32'h8c50000;
      59524: inst = 32'h24612800;
      59525: inst = 32'h10a0ffff;
      59526: inst = 32'hca0fff2;
      59527: inst = 32'h24822800;
      59528: inst = 32'h10a00000;
      59529: inst = 32'hca00004;
      59530: inst = 32'h38632800;
      59531: inst = 32'h38842800;
      59532: inst = 32'h10a00000;
      59533: inst = 32'hca0e891;
      59534: inst = 32'h13e00001;
      59535: inst = 32'hfe0d96a;
      59536: inst = 32'h5be00000;
      59537: inst = 32'h8c50000;
      59538: inst = 32'h24612800;
      59539: inst = 32'h10a0ffff;
      59540: inst = 32'hca0fff2;
      59541: inst = 32'h24822800;
      59542: inst = 32'h10a00000;
      59543: inst = 32'hca00004;
      59544: inst = 32'h38632800;
      59545: inst = 32'h38842800;
      59546: inst = 32'h10a00000;
      59547: inst = 32'hca0e89f;
      59548: inst = 32'h13e00001;
      59549: inst = 32'hfe0d96a;
      59550: inst = 32'h5be00000;
      59551: inst = 32'h8c50000;
      59552: inst = 32'h24612800;
      59553: inst = 32'h10a0ffff;
      59554: inst = 32'hca0fff2;
      59555: inst = 32'h24822800;
      59556: inst = 32'h10a00000;
      59557: inst = 32'hca00004;
      59558: inst = 32'h38632800;
      59559: inst = 32'h38842800;
      59560: inst = 32'h10a00000;
      59561: inst = 32'hca0e8ad;
      59562: inst = 32'h13e00001;
      59563: inst = 32'hfe0d96a;
      59564: inst = 32'h5be00000;
      59565: inst = 32'h8c50000;
      59566: inst = 32'h24612800;
      59567: inst = 32'h10a0ffff;
      59568: inst = 32'hca0fff2;
      59569: inst = 32'h24822800;
      59570: inst = 32'h10a00000;
      59571: inst = 32'hca00004;
      59572: inst = 32'h38632800;
      59573: inst = 32'h38842800;
      59574: inst = 32'h10a00000;
      59575: inst = 32'hca0e8bb;
      59576: inst = 32'h13e00001;
      59577: inst = 32'hfe0d96a;
      59578: inst = 32'h5be00000;
      59579: inst = 32'h8c50000;
      59580: inst = 32'h24612800;
      59581: inst = 32'h10a0ffff;
      59582: inst = 32'hca0fff2;
      59583: inst = 32'h24822800;
      59584: inst = 32'h10a00000;
      59585: inst = 32'hca00004;
      59586: inst = 32'h38632800;
      59587: inst = 32'h38842800;
      59588: inst = 32'h10a00000;
      59589: inst = 32'hca0e8c9;
      59590: inst = 32'h13e00001;
      59591: inst = 32'hfe0d96a;
      59592: inst = 32'h5be00000;
      59593: inst = 32'h8c50000;
      59594: inst = 32'h24612800;
      59595: inst = 32'h10a0ffff;
      59596: inst = 32'hca0fff2;
      59597: inst = 32'h24822800;
      59598: inst = 32'h10a00000;
      59599: inst = 32'hca00004;
      59600: inst = 32'h38632800;
      59601: inst = 32'h38842800;
      59602: inst = 32'h10a00000;
      59603: inst = 32'hca0e8d7;
      59604: inst = 32'h13e00001;
      59605: inst = 32'hfe0d96a;
      59606: inst = 32'h5be00000;
      59607: inst = 32'h8c50000;
      59608: inst = 32'h24612800;
      59609: inst = 32'h10a0ffff;
      59610: inst = 32'hca0fff2;
      59611: inst = 32'h24822800;
      59612: inst = 32'h10a00000;
      59613: inst = 32'hca00004;
      59614: inst = 32'h38632800;
      59615: inst = 32'h38842800;
      59616: inst = 32'h10a00000;
      59617: inst = 32'hca0e8e5;
      59618: inst = 32'h13e00001;
      59619: inst = 32'hfe0d96a;
      59620: inst = 32'h5be00000;
      59621: inst = 32'h8c50000;
      59622: inst = 32'h24612800;
      59623: inst = 32'h10a0ffff;
      59624: inst = 32'hca0fff2;
      59625: inst = 32'h24822800;
      59626: inst = 32'h10a00000;
      59627: inst = 32'hca00004;
      59628: inst = 32'h38632800;
      59629: inst = 32'h38842800;
      59630: inst = 32'h10a00000;
      59631: inst = 32'hca0e8f3;
      59632: inst = 32'h13e00001;
      59633: inst = 32'hfe0d96a;
      59634: inst = 32'h5be00000;
      59635: inst = 32'h8c50000;
      59636: inst = 32'h24612800;
      59637: inst = 32'h10a0ffff;
      59638: inst = 32'hca0fff2;
      59639: inst = 32'h24822800;
      59640: inst = 32'h10a00000;
      59641: inst = 32'hca00004;
      59642: inst = 32'h38632800;
      59643: inst = 32'h38842800;
      59644: inst = 32'h10a00000;
      59645: inst = 32'hca0e901;
      59646: inst = 32'h13e00001;
      59647: inst = 32'hfe0d96a;
      59648: inst = 32'h5be00000;
      59649: inst = 32'h8c50000;
      59650: inst = 32'h24612800;
      59651: inst = 32'h10a0ffff;
      59652: inst = 32'hca0fff2;
      59653: inst = 32'h24822800;
      59654: inst = 32'h10a00000;
      59655: inst = 32'hca00004;
      59656: inst = 32'h38632800;
      59657: inst = 32'h38842800;
      59658: inst = 32'h10a00000;
      59659: inst = 32'hca0e90f;
      59660: inst = 32'h13e00001;
      59661: inst = 32'hfe0d96a;
      59662: inst = 32'h5be00000;
      59663: inst = 32'h8c50000;
      59664: inst = 32'h24612800;
      59665: inst = 32'h10a0ffff;
      59666: inst = 32'hca0fff2;
      59667: inst = 32'h24822800;
      59668: inst = 32'h10a00000;
      59669: inst = 32'hca00004;
      59670: inst = 32'h38632800;
      59671: inst = 32'h38842800;
      59672: inst = 32'h10a00000;
      59673: inst = 32'hca0e91d;
      59674: inst = 32'h13e00001;
      59675: inst = 32'hfe0d96a;
      59676: inst = 32'h5be00000;
      59677: inst = 32'h8c50000;
      59678: inst = 32'h24612800;
      59679: inst = 32'h10a0ffff;
      59680: inst = 32'hca0fff2;
      59681: inst = 32'h24822800;
      59682: inst = 32'h10a00000;
      59683: inst = 32'hca00004;
      59684: inst = 32'h38632800;
      59685: inst = 32'h38842800;
      59686: inst = 32'h10a00000;
      59687: inst = 32'hca0e92b;
      59688: inst = 32'h13e00001;
      59689: inst = 32'hfe0d96a;
      59690: inst = 32'h5be00000;
      59691: inst = 32'h8c50000;
      59692: inst = 32'h24612800;
      59693: inst = 32'h10a0ffff;
      59694: inst = 32'hca0fff2;
      59695: inst = 32'h24822800;
      59696: inst = 32'h10a00000;
      59697: inst = 32'hca00004;
      59698: inst = 32'h38632800;
      59699: inst = 32'h38842800;
      59700: inst = 32'h10a00000;
      59701: inst = 32'hca0e939;
      59702: inst = 32'h13e00001;
      59703: inst = 32'hfe0d96a;
      59704: inst = 32'h5be00000;
      59705: inst = 32'h8c50000;
      59706: inst = 32'h24612800;
      59707: inst = 32'h10a0ffff;
      59708: inst = 32'hca0fff2;
      59709: inst = 32'h24822800;
      59710: inst = 32'h10a00000;
      59711: inst = 32'hca00004;
      59712: inst = 32'h38632800;
      59713: inst = 32'h38842800;
      59714: inst = 32'h10a00000;
      59715: inst = 32'hca0e947;
      59716: inst = 32'h13e00001;
      59717: inst = 32'hfe0d96a;
      59718: inst = 32'h5be00000;
      59719: inst = 32'h8c50000;
      59720: inst = 32'h24612800;
      59721: inst = 32'h10a0ffff;
      59722: inst = 32'hca0fff2;
      59723: inst = 32'h24822800;
      59724: inst = 32'h10a00000;
      59725: inst = 32'hca00004;
      59726: inst = 32'h38632800;
      59727: inst = 32'h38842800;
      59728: inst = 32'h10a00000;
      59729: inst = 32'hca0e955;
      59730: inst = 32'h13e00001;
      59731: inst = 32'hfe0d96a;
      59732: inst = 32'h5be00000;
      59733: inst = 32'h8c50000;
      59734: inst = 32'h24612800;
      59735: inst = 32'h10a0ffff;
      59736: inst = 32'hca0fff2;
      59737: inst = 32'h24822800;
      59738: inst = 32'h10a00000;
      59739: inst = 32'hca00004;
      59740: inst = 32'h38632800;
      59741: inst = 32'h38842800;
      59742: inst = 32'h10a00000;
      59743: inst = 32'hca0e963;
      59744: inst = 32'h13e00001;
      59745: inst = 32'hfe0d96a;
      59746: inst = 32'h5be00000;
      59747: inst = 32'h8c50000;
      59748: inst = 32'h24612800;
      59749: inst = 32'h10a0ffff;
      59750: inst = 32'hca0fff2;
      59751: inst = 32'h24822800;
      59752: inst = 32'h10a00000;
      59753: inst = 32'hca00004;
      59754: inst = 32'h38632800;
      59755: inst = 32'h38842800;
      59756: inst = 32'h10a00000;
      59757: inst = 32'hca0e971;
      59758: inst = 32'h13e00001;
      59759: inst = 32'hfe0d96a;
      59760: inst = 32'h5be00000;
      59761: inst = 32'h8c50000;
      59762: inst = 32'h24612800;
      59763: inst = 32'h10a0ffff;
      59764: inst = 32'hca0fff2;
      59765: inst = 32'h24822800;
      59766: inst = 32'h10a00000;
      59767: inst = 32'hca00004;
      59768: inst = 32'h38632800;
      59769: inst = 32'h38842800;
      59770: inst = 32'h10a00000;
      59771: inst = 32'hca0e97f;
      59772: inst = 32'h13e00001;
      59773: inst = 32'hfe0d96a;
      59774: inst = 32'h5be00000;
      59775: inst = 32'h8c50000;
      59776: inst = 32'h24612800;
      59777: inst = 32'h10a0ffff;
      59778: inst = 32'hca0fff2;
      59779: inst = 32'h24822800;
      59780: inst = 32'h10a00000;
      59781: inst = 32'hca00004;
      59782: inst = 32'h38632800;
      59783: inst = 32'h38842800;
      59784: inst = 32'h10a00000;
      59785: inst = 32'hca0e98d;
      59786: inst = 32'h13e00001;
      59787: inst = 32'hfe0d96a;
      59788: inst = 32'h5be00000;
      59789: inst = 32'h8c50000;
      59790: inst = 32'h24612800;
      59791: inst = 32'h10a0ffff;
      59792: inst = 32'hca0fff2;
      59793: inst = 32'h24822800;
      59794: inst = 32'h10a00000;
      59795: inst = 32'hca00004;
      59796: inst = 32'h38632800;
      59797: inst = 32'h38842800;
      59798: inst = 32'h10a00000;
      59799: inst = 32'hca0e99b;
      59800: inst = 32'h13e00001;
      59801: inst = 32'hfe0d96a;
      59802: inst = 32'h5be00000;
      59803: inst = 32'h8c50000;
      59804: inst = 32'h24612800;
      59805: inst = 32'h10a0ffff;
      59806: inst = 32'hca0fff2;
      59807: inst = 32'h24822800;
      59808: inst = 32'h10a00000;
      59809: inst = 32'hca00004;
      59810: inst = 32'h38632800;
      59811: inst = 32'h38842800;
      59812: inst = 32'h10a00000;
      59813: inst = 32'hca0e9a9;
      59814: inst = 32'h13e00001;
      59815: inst = 32'hfe0d96a;
      59816: inst = 32'h5be00000;
      59817: inst = 32'h8c50000;
      59818: inst = 32'h24612800;
      59819: inst = 32'h10a0ffff;
      59820: inst = 32'hca0fff2;
      59821: inst = 32'h24822800;
      59822: inst = 32'h10a00000;
      59823: inst = 32'hca00004;
      59824: inst = 32'h38632800;
      59825: inst = 32'h38842800;
      59826: inst = 32'h10a00000;
      59827: inst = 32'hca0e9b7;
      59828: inst = 32'h13e00001;
      59829: inst = 32'hfe0d96a;
      59830: inst = 32'h5be00000;
      59831: inst = 32'h8c50000;
      59832: inst = 32'h24612800;
      59833: inst = 32'h10a0ffff;
      59834: inst = 32'hca0fff2;
      59835: inst = 32'h24822800;
      59836: inst = 32'h10a00000;
      59837: inst = 32'hca00004;
      59838: inst = 32'h38632800;
      59839: inst = 32'h38842800;
      59840: inst = 32'h10a00000;
      59841: inst = 32'hca0e9c5;
      59842: inst = 32'h13e00001;
      59843: inst = 32'hfe0d96a;
      59844: inst = 32'h5be00000;
      59845: inst = 32'h8c50000;
      59846: inst = 32'h24612800;
      59847: inst = 32'h10a0ffff;
      59848: inst = 32'hca0fff2;
      59849: inst = 32'h24822800;
      59850: inst = 32'h10a00000;
      59851: inst = 32'hca00004;
      59852: inst = 32'h38632800;
      59853: inst = 32'h38842800;
      59854: inst = 32'h10a00000;
      59855: inst = 32'hca0e9d3;
      59856: inst = 32'h13e00001;
      59857: inst = 32'hfe0d96a;
      59858: inst = 32'h5be00000;
      59859: inst = 32'h8c50000;
      59860: inst = 32'h24612800;
      59861: inst = 32'h10a0ffff;
      59862: inst = 32'hca0fff2;
      59863: inst = 32'h24822800;
      59864: inst = 32'h10a00000;
      59865: inst = 32'hca00004;
      59866: inst = 32'h38632800;
      59867: inst = 32'h38842800;
      59868: inst = 32'h10a00000;
      59869: inst = 32'hca0e9e1;
      59870: inst = 32'h13e00001;
      59871: inst = 32'hfe0d96a;
      59872: inst = 32'h5be00000;
      59873: inst = 32'h8c50000;
      59874: inst = 32'h24612800;
      59875: inst = 32'h10a0ffff;
      59876: inst = 32'hca0fff2;
      59877: inst = 32'h24822800;
      59878: inst = 32'h10a00000;
      59879: inst = 32'hca00004;
      59880: inst = 32'h38632800;
      59881: inst = 32'h38842800;
      59882: inst = 32'h10a00000;
      59883: inst = 32'hca0e9ef;
      59884: inst = 32'h13e00001;
      59885: inst = 32'hfe0d96a;
      59886: inst = 32'h5be00000;
      59887: inst = 32'h8c50000;
      59888: inst = 32'h24612800;
      59889: inst = 32'h10a0ffff;
      59890: inst = 32'hca0fff2;
      59891: inst = 32'h24822800;
      59892: inst = 32'h10a00000;
      59893: inst = 32'hca00004;
      59894: inst = 32'h38632800;
      59895: inst = 32'h38842800;
      59896: inst = 32'h10a00000;
      59897: inst = 32'hca0e9fd;
      59898: inst = 32'h13e00001;
      59899: inst = 32'hfe0d96a;
      59900: inst = 32'h5be00000;
      59901: inst = 32'h8c50000;
      59902: inst = 32'h24612800;
      59903: inst = 32'h10a0ffff;
      59904: inst = 32'hca0fff2;
      59905: inst = 32'h24822800;
      59906: inst = 32'h10a00000;
      59907: inst = 32'hca00004;
      59908: inst = 32'h38632800;
      59909: inst = 32'h38842800;
      59910: inst = 32'h10a00000;
      59911: inst = 32'hca0ea0b;
      59912: inst = 32'h13e00001;
      59913: inst = 32'hfe0d96a;
      59914: inst = 32'h5be00000;
      59915: inst = 32'h8c50000;
      59916: inst = 32'h24612800;
      59917: inst = 32'h10a0ffff;
      59918: inst = 32'hca0fff2;
      59919: inst = 32'h24822800;
      59920: inst = 32'h10a00000;
      59921: inst = 32'hca00004;
      59922: inst = 32'h38632800;
      59923: inst = 32'h38842800;
      59924: inst = 32'h10a00000;
      59925: inst = 32'hca0ea19;
      59926: inst = 32'h13e00001;
      59927: inst = 32'hfe0d96a;
      59928: inst = 32'h5be00000;
      59929: inst = 32'h8c50000;
      59930: inst = 32'h24612800;
      59931: inst = 32'h10a0ffff;
      59932: inst = 32'hca0fff2;
      59933: inst = 32'h24822800;
      59934: inst = 32'h10a00000;
      59935: inst = 32'hca00004;
      59936: inst = 32'h38632800;
      59937: inst = 32'h38842800;
      59938: inst = 32'h10a00000;
      59939: inst = 32'hca0ea27;
      59940: inst = 32'h13e00001;
      59941: inst = 32'hfe0d96a;
      59942: inst = 32'h5be00000;
      59943: inst = 32'h8c50000;
      59944: inst = 32'h24612800;
      59945: inst = 32'h10a0ffff;
      59946: inst = 32'hca0fff2;
      59947: inst = 32'h24822800;
      59948: inst = 32'h10a00000;
      59949: inst = 32'hca00004;
      59950: inst = 32'h38632800;
      59951: inst = 32'h38842800;
      59952: inst = 32'h10a00000;
      59953: inst = 32'hca0ea35;
      59954: inst = 32'h13e00001;
      59955: inst = 32'hfe0d96a;
      59956: inst = 32'h5be00000;
      59957: inst = 32'h8c50000;
      59958: inst = 32'h24612800;
      59959: inst = 32'h10a0ffff;
      59960: inst = 32'hca0fff2;
      59961: inst = 32'h24822800;
      59962: inst = 32'h10a00000;
      59963: inst = 32'hca00004;
      59964: inst = 32'h38632800;
      59965: inst = 32'h38842800;
      59966: inst = 32'h10a00000;
      59967: inst = 32'hca0ea43;
      59968: inst = 32'h13e00001;
      59969: inst = 32'hfe0d96a;
      59970: inst = 32'h5be00000;
      59971: inst = 32'h8c50000;
      59972: inst = 32'h24612800;
      59973: inst = 32'h10a0ffff;
      59974: inst = 32'hca0fff2;
      59975: inst = 32'h24822800;
      59976: inst = 32'h10a00000;
      59977: inst = 32'hca00004;
      59978: inst = 32'h38632800;
      59979: inst = 32'h38842800;
      59980: inst = 32'h10a00000;
      59981: inst = 32'hca0ea51;
      59982: inst = 32'h13e00001;
      59983: inst = 32'hfe0d96a;
      59984: inst = 32'h5be00000;
      59985: inst = 32'h8c50000;
      59986: inst = 32'h24612800;
      59987: inst = 32'h10a0ffff;
      59988: inst = 32'hca0fff2;
      59989: inst = 32'h24822800;
      59990: inst = 32'h10a00000;
      59991: inst = 32'hca00004;
      59992: inst = 32'h38632800;
      59993: inst = 32'h38842800;
      59994: inst = 32'h10a00000;
      59995: inst = 32'hca0ea5f;
      59996: inst = 32'h13e00001;
      59997: inst = 32'hfe0d96a;
      59998: inst = 32'h5be00000;
      59999: inst = 32'h8c50000;
      60000: inst = 32'h24612800;
      60001: inst = 32'h10a0ffff;
      60002: inst = 32'hca0fff2;
      60003: inst = 32'h24822800;
      60004: inst = 32'h10a00000;
      60005: inst = 32'hca00004;
      60006: inst = 32'h38632800;
      60007: inst = 32'h38842800;
      60008: inst = 32'h10a00000;
      60009: inst = 32'hca0ea6d;
      60010: inst = 32'h13e00001;
      60011: inst = 32'hfe0d96a;
      60012: inst = 32'h5be00000;
      60013: inst = 32'h8c50000;
      60014: inst = 32'h24612800;
      60015: inst = 32'h10a0ffff;
      60016: inst = 32'hca0fff2;
      60017: inst = 32'h24822800;
      60018: inst = 32'h10a00000;
      60019: inst = 32'hca00004;
      60020: inst = 32'h38632800;
      60021: inst = 32'h38842800;
      60022: inst = 32'h10a00000;
      60023: inst = 32'hca0ea7b;
      60024: inst = 32'h13e00001;
      60025: inst = 32'hfe0d96a;
      60026: inst = 32'h5be00000;
      60027: inst = 32'h8c50000;
      60028: inst = 32'h24612800;
      60029: inst = 32'h10a0ffff;
      60030: inst = 32'hca0fff2;
      60031: inst = 32'h24822800;
      60032: inst = 32'h10a00000;
      60033: inst = 32'hca00004;
      60034: inst = 32'h38632800;
      60035: inst = 32'h38842800;
      60036: inst = 32'h10a00000;
      60037: inst = 32'hca0ea89;
      60038: inst = 32'h13e00001;
      60039: inst = 32'hfe0d96a;
      60040: inst = 32'h5be00000;
      60041: inst = 32'h8c50000;
      60042: inst = 32'h24612800;
      60043: inst = 32'h10a0ffff;
      60044: inst = 32'hca0fff2;
      60045: inst = 32'h24822800;
      60046: inst = 32'h10a00000;
      60047: inst = 32'hca00004;
      60048: inst = 32'h38632800;
      60049: inst = 32'h38842800;
      60050: inst = 32'h10a00000;
      60051: inst = 32'hca0ea97;
      60052: inst = 32'h13e00001;
      60053: inst = 32'hfe0d96a;
      60054: inst = 32'h5be00000;
      60055: inst = 32'h8c50000;
      60056: inst = 32'h24612800;
      60057: inst = 32'h10a0ffff;
      60058: inst = 32'hca0fff2;
      60059: inst = 32'h24822800;
      60060: inst = 32'h10a00000;
      60061: inst = 32'hca00004;
      60062: inst = 32'h38632800;
      60063: inst = 32'h38842800;
      60064: inst = 32'h10a00000;
      60065: inst = 32'hca0eaa5;
      60066: inst = 32'h13e00001;
      60067: inst = 32'hfe0d96a;
      60068: inst = 32'h5be00000;
      60069: inst = 32'h8c50000;
      60070: inst = 32'h24612800;
      60071: inst = 32'h10a0ffff;
      60072: inst = 32'hca0fff2;
      60073: inst = 32'h24822800;
      60074: inst = 32'h10a00000;
      60075: inst = 32'hca00004;
      60076: inst = 32'h38632800;
      60077: inst = 32'h38842800;
      60078: inst = 32'h10a00000;
      60079: inst = 32'hca0eab3;
      60080: inst = 32'h13e00001;
      60081: inst = 32'hfe0d96a;
      60082: inst = 32'h5be00000;
      60083: inst = 32'h8c50000;
      60084: inst = 32'h24612800;
      60085: inst = 32'h10a0ffff;
      60086: inst = 32'hca0fff2;
      60087: inst = 32'h24822800;
      60088: inst = 32'h10a00000;
      60089: inst = 32'hca00004;
      60090: inst = 32'h38632800;
      60091: inst = 32'h38842800;
      60092: inst = 32'h10a00000;
      60093: inst = 32'hca0eac1;
      60094: inst = 32'h13e00001;
      60095: inst = 32'hfe0d96a;
      60096: inst = 32'h5be00000;
      60097: inst = 32'h8c50000;
      60098: inst = 32'h24612800;
      60099: inst = 32'h10a0ffff;
      60100: inst = 32'hca0fff2;
      60101: inst = 32'h24822800;
      60102: inst = 32'h10a00000;
      60103: inst = 32'hca00004;
      60104: inst = 32'h38632800;
      60105: inst = 32'h38842800;
      60106: inst = 32'h10a00000;
      60107: inst = 32'hca0eacf;
      60108: inst = 32'h13e00001;
      60109: inst = 32'hfe0d96a;
      60110: inst = 32'h5be00000;
      60111: inst = 32'h8c50000;
      60112: inst = 32'h24612800;
      60113: inst = 32'h10a0ffff;
      60114: inst = 32'hca0fff2;
      60115: inst = 32'h24822800;
      60116: inst = 32'h10a00000;
      60117: inst = 32'hca00004;
      60118: inst = 32'h38632800;
      60119: inst = 32'h38842800;
      60120: inst = 32'h10a00000;
      60121: inst = 32'hca0eadd;
      60122: inst = 32'h13e00001;
      60123: inst = 32'hfe0d96a;
      60124: inst = 32'h5be00000;
      60125: inst = 32'h8c50000;
      60126: inst = 32'h24612800;
      60127: inst = 32'h10a0ffff;
      60128: inst = 32'hca0fff2;
      60129: inst = 32'h24822800;
      60130: inst = 32'h10a00000;
      60131: inst = 32'hca00004;
      60132: inst = 32'h38632800;
      60133: inst = 32'h38842800;
      60134: inst = 32'h10a00000;
      60135: inst = 32'hca0eaeb;
      60136: inst = 32'h13e00001;
      60137: inst = 32'hfe0d96a;
      60138: inst = 32'h5be00000;
      60139: inst = 32'h8c50000;
      60140: inst = 32'h24612800;
      60141: inst = 32'h10a0ffff;
      60142: inst = 32'hca0fff2;
      60143: inst = 32'h24822800;
      60144: inst = 32'h10a00000;
      60145: inst = 32'hca00004;
      60146: inst = 32'h38632800;
      60147: inst = 32'h38842800;
      60148: inst = 32'h10a00000;
      60149: inst = 32'hca0eaf9;
      60150: inst = 32'h13e00001;
      60151: inst = 32'hfe0d96a;
      60152: inst = 32'h5be00000;
      60153: inst = 32'h8c50000;
      60154: inst = 32'h24612800;
      60155: inst = 32'h10a0ffff;
      60156: inst = 32'hca0fff2;
      60157: inst = 32'h24822800;
      60158: inst = 32'h10a00000;
      60159: inst = 32'hca00004;
      60160: inst = 32'h38632800;
      60161: inst = 32'h38842800;
      60162: inst = 32'h10a00000;
      60163: inst = 32'hca0eb07;
      60164: inst = 32'h13e00001;
      60165: inst = 32'hfe0d96a;
      60166: inst = 32'h5be00000;
      60167: inst = 32'h8c50000;
      60168: inst = 32'h24612800;
      60169: inst = 32'h10a0ffff;
      60170: inst = 32'hca0fff2;
      60171: inst = 32'h24822800;
      60172: inst = 32'h10a00000;
      60173: inst = 32'hca00004;
      60174: inst = 32'h38632800;
      60175: inst = 32'h38842800;
      60176: inst = 32'h10a00000;
      60177: inst = 32'hca0eb15;
      60178: inst = 32'h13e00001;
      60179: inst = 32'hfe0d96a;
      60180: inst = 32'h5be00000;
      60181: inst = 32'h8c50000;
      60182: inst = 32'h24612800;
      60183: inst = 32'h10a0ffff;
      60184: inst = 32'hca0fff2;
      60185: inst = 32'h24822800;
      60186: inst = 32'h10a00000;
      60187: inst = 32'hca00004;
      60188: inst = 32'h38632800;
      60189: inst = 32'h38842800;
      60190: inst = 32'h10a00000;
      60191: inst = 32'hca0eb23;
      60192: inst = 32'h13e00001;
      60193: inst = 32'hfe0d96a;
      60194: inst = 32'h5be00000;
      60195: inst = 32'h8c50000;
      60196: inst = 32'h24612800;
      60197: inst = 32'h10a0ffff;
      60198: inst = 32'hca0fff2;
      60199: inst = 32'h24822800;
      60200: inst = 32'h10a00000;
      60201: inst = 32'hca00004;
      60202: inst = 32'h38632800;
      60203: inst = 32'h38842800;
      60204: inst = 32'h10a00000;
      60205: inst = 32'hca0eb31;
      60206: inst = 32'h13e00001;
      60207: inst = 32'hfe0d96a;
      60208: inst = 32'h5be00000;
      60209: inst = 32'h8c50000;
      60210: inst = 32'h24612800;
      60211: inst = 32'h10a0ffff;
      60212: inst = 32'hca0fff2;
      60213: inst = 32'h24822800;
      60214: inst = 32'h10a00000;
      60215: inst = 32'hca00004;
      60216: inst = 32'h38632800;
      60217: inst = 32'h38842800;
      60218: inst = 32'h10a00000;
      60219: inst = 32'hca0eb3f;
      60220: inst = 32'h13e00001;
      60221: inst = 32'hfe0d96a;
      60222: inst = 32'h5be00000;
      60223: inst = 32'h8c50000;
      60224: inst = 32'h24612800;
      60225: inst = 32'h10a0ffff;
      60226: inst = 32'hca0fff2;
      60227: inst = 32'h24822800;
      60228: inst = 32'h10a00000;
      60229: inst = 32'hca00004;
      60230: inst = 32'h38632800;
      60231: inst = 32'h38842800;
      60232: inst = 32'h10a00000;
      60233: inst = 32'hca0eb4d;
      60234: inst = 32'h13e00001;
      60235: inst = 32'hfe0d96a;
      60236: inst = 32'h5be00000;
      60237: inst = 32'h8c50000;
      60238: inst = 32'h24612800;
      60239: inst = 32'h10a0ffff;
      60240: inst = 32'hca0fff2;
      60241: inst = 32'h24822800;
      60242: inst = 32'h10a00000;
      60243: inst = 32'hca00004;
      60244: inst = 32'h38632800;
      60245: inst = 32'h38842800;
      60246: inst = 32'h10a00000;
      60247: inst = 32'hca0eb5b;
      60248: inst = 32'h13e00001;
      60249: inst = 32'hfe0d96a;
      60250: inst = 32'h5be00000;
      60251: inst = 32'h8c50000;
      60252: inst = 32'h24612800;
      60253: inst = 32'h10a0ffff;
      60254: inst = 32'hca0fff2;
      60255: inst = 32'h24822800;
      60256: inst = 32'h10a00000;
      60257: inst = 32'hca00004;
      60258: inst = 32'h38632800;
      60259: inst = 32'h38842800;
      60260: inst = 32'h10a00000;
      60261: inst = 32'hca0eb69;
      60262: inst = 32'h13e00001;
      60263: inst = 32'hfe0d96a;
      60264: inst = 32'h5be00000;
      60265: inst = 32'h8c50000;
      60266: inst = 32'h24612800;
      60267: inst = 32'h10a0ffff;
      60268: inst = 32'hca0fff2;
      60269: inst = 32'h24822800;
      60270: inst = 32'h10a00000;
      60271: inst = 32'hca00004;
      60272: inst = 32'h38632800;
      60273: inst = 32'h38842800;
      60274: inst = 32'h10a00000;
      60275: inst = 32'hca0eb77;
      60276: inst = 32'h13e00001;
      60277: inst = 32'hfe0d96a;
      60278: inst = 32'h5be00000;
      60279: inst = 32'h8c50000;
      60280: inst = 32'h24612800;
      60281: inst = 32'h10a0ffff;
      60282: inst = 32'hca0fff2;
      60283: inst = 32'h24822800;
      60284: inst = 32'h10a00000;
      60285: inst = 32'hca00004;
      60286: inst = 32'h38632800;
      60287: inst = 32'h38842800;
      60288: inst = 32'h10a00000;
      60289: inst = 32'hca0eb85;
      60290: inst = 32'h13e00001;
      60291: inst = 32'hfe0d96a;
      60292: inst = 32'h5be00000;
      60293: inst = 32'h8c50000;
      60294: inst = 32'h24612800;
      60295: inst = 32'h10a0ffff;
      60296: inst = 32'hca0fff2;
      60297: inst = 32'h24822800;
      60298: inst = 32'h10a00000;
      60299: inst = 32'hca00004;
      60300: inst = 32'h38632800;
      60301: inst = 32'h38842800;
      60302: inst = 32'h10a00000;
      60303: inst = 32'hca0eb93;
      60304: inst = 32'h13e00001;
      60305: inst = 32'hfe0d96a;
      60306: inst = 32'h5be00000;
      60307: inst = 32'h8c50000;
      60308: inst = 32'h24612800;
      60309: inst = 32'h10a0ffff;
      60310: inst = 32'hca0fff2;
      60311: inst = 32'h24822800;
      60312: inst = 32'h10a00000;
      60313: inst = 32'hca00004;
      60314: inst = 32'h38632800;
      60315: inst = 32'h38842800;
      60316: inst = 32'h10a00000;
      60317: inst = 32'hca0eba1;
      60318: inst = 32'h13e00001;
      60319: inst = 32'hfe0d96a;
      60320: inst = 32'h5be00000;
      60321: inst = 32'h8c50000;
      60322: inst = 32'h24612800;
      60323: inst = 32'h10a0ffff;
      60324: inst = 32'hca0fff2;
      60325: inst = 32'h24822800;
      60326: inst = 32'h10a00000;
      60327: inst = 32'hca00004;
      60328: inst = 32'h38632800;
      60329: inst = 32'h38842800;
      60330: inst = 32'h10a00000;
      60331: inst = 32'hca0ebaf;
      60332: inst = 32'h13e00001;
      60333: inst = 32'hfe0d96a;
      60334: inst = 32'h5be00000;
      60335: inst = 32'h8c50000;
      60336: inst = 32'h24612800;
      60337: inst = 32'h10a0ffff;
      60338: inst = 32'hca0fff2;
      60339: inst = 32'h24822800;
      60340: inst = 32'h10a00000;
      60341: inst = 32'hca00004;
      60342: inst = 32'h38632800;
      60343: inst = 32'h38842800;
      60344: inst = 32'h10a00000;
      60345: inst = 32'hca0ebbd;
      60346: inst = 32'h13e00001;
      60347: inst = 32'hfe0d96a;
      60348: inst = 32'h5be00000;
      60349: inst = 32'h8c50000;
      60350: inst = 32'h24612800;
      60351: inst = 32'h10a0ffff;
      60352: inst = 32'hca0fff2;
      60353: inst = 32'h24822800;
      60354: inst = 32'h10a00000;
      60355: inst = 32'hca00004;
      60356: inst = 32'h38632800;
      60357: inst = 32'h38842800;
      60358: inst = 32'h10a00000;
      60359: inst = 32'hca0ebcb;
      60360: inst = 32'h13e00001;
      60361: inst = 32'hfe0d96a;
      60362: inst = 32'h5be00000;
      60363: inst = 32'h8c50000;
      60364: inst = 32'h24612800;
      60365: inst = 32'h10a0ffff;
      60366: inst = 32'hca0fff2;
      60367: inst = 32'h24822800;
      60368: inst = 32'h10a00000;
      60369: inst = 32'hca00004;
      60370: inst = 32'h38632800;
      60371: inst = 32'h38842800;
      60372: inst = 32'h10a00000;
      60373: inst = 32'hca0ebd9;
      60374: inst = 32'h13e00001;
      60375: inst = 32'hfe0d96a;
      60376: inst = 32'h5be00000;
      60377: inst = 32'h8c50000;
      60378: inst = 32'h24612800;
      60379: inst = 32'h10a0ffff;
      60380: inst = 32'hca0fff2;
      60381: inst = 32'h24822800;
      60382: inst = 32'h10a00000;
      60383: inst = 32'hca00004;
      60384: inst = 32'h38632800;
      60385: inst = 32'h38842800;
      60386: inst = 32'h10a00000;
      60387: inst = 32'hca0ebe7;
      60388: inst = 32'h13e00001;
      60389: inst = 32'hfe0d96a;
      60390: inst = 32'h5be00000;
      60391: inst = 32'h8c50000;
      60392: inst = 32'h24612800;
      60393: inst = 32'h10a0ffff;
      60394: inst = 32'hca0fff2;
      60395: inst = 32'h24822800;
      60396: inst = 32'h10a00000;
      60397: inst = 32'hca00004;
      60398: inst = 32'h38632800;
      60399: inst = 32'h38842800;
      60400: inst = 32'h10a00000;
      60401: inst = 32'hca0ebf5;
      60402: inst = 32'h13e00001;
      60403: inst = 32'hfe0d96a;
      60404: inst = 32'h5be00000;
      60405: inst = 32'h8c50000;
      60406: inst = 32'h24612800;
      60407: inst = 32'h10a0ffff;
      60408: inst = 32'hca0fff2;
      60409: inst = 32'h24822800;
      60410: inst = 32'h10a00000;
      60411: inst = 32'hca00004;
      60412: inst = 32'h38632800;
      60413: inst = 32'h38842800;
      60414: inst = 32'h10a00000;
      60415: inst = 32'hca0ec03;
      60416: inst = 32'h13e00001;
      60417: inst = 32'hfe0d96a;
      60418: inst = 32'h5be00000;
      60419: inst = 32'h8c50000;
      60420: inst = 32'h24612800;
      60421: inst = 32'h10a0ffff;
      60422: inst = 32'hca0fff2;
      60423: inst = 32'h24822800;
      60424: inst = 32'h10a00000;
      60425: inst = 32'hca00004;
      60426: inst = 32'h38632800;
      60427: inst = 32'h38842800;
      60428: inst = 32'h10a00000;
      60429: inst = 32'hca0ec11;
      60430: inst = 32'h13e00001;
      60431: inst = 32'hfe0d96a;
      60432: inst = 32'h5be00000;
      60433: inst = 32'h8c50000;
      60434: inst = 32'h24612800;
      60435: inst = 32'h10a0ffff;
      60436: inst = 32'hca0fff2;
      60437: inst = 32'h24822800;
      60438: inst = 32'h10a00000;
      60439: inst = 32'hca00004;
      60440: inst = 32'h38632800;
      60441: inst = 32'h38842800;
      60442: inst = 32'h10a00000;
      60443: inst = 32'hca0ec1f;
      60444: inst = 32'h13e00001;
      60445: inst = 32'hfe0d96a;
      60446: inst = 32'h5be00000;
      60447: inst = 32'h8c50000;
      60448: inst = 32'h24612800;
      60449: inst = 32'h10a0ffff;
      60450: inst = 32'hca0fff2;
      60451: inst = 32'h24822800;
      60452: inst = 32'h10a00000;
      60453: inst = 32'hca00004;
      60454: inst = 32'h38632800;
      60455: inst = 32'h38842800;
      60456: inst = 32'h10a00000;
      60457: inst = 32'hca0ec2d;
      60458: inst = 32'h13e00001;
      60459: inst = 32'hfe0d96a;
      60460: inst = 32'h5be00000;
      60461: inst = 32'h8c50000;
      60462: inst = 32'h24612800;
      60463: inst = 32'h10a0ffff;
      60464: inst = 32'hca0fff2;
      60465: inst = 32'h24822800;
      60466: inst = 32'h10a00000;
      60467: inst = 32'hca00004;
      60468: inst = 32'h38632800;
      60469: inst = 32'h38842800;
      60470: inst = 32'h10a00000;
      60471: inst = 32'hca0ec3b;
      60472: inst = 32'h13e00001;
      60473: inst = 32'hfe0d96a;
      60474: inst = 32'h5be00000;
      60475: inst = 32'h8c50000;
      60476: inst = 32'h24612800;
      60477: inst = 32'h10a0ffff;
      60478: inst = 32'hca0fff2;
      60479: inst = 32'h24822800;
      60480: inst = 32'h10a00000;
      60481: inst = 32'hca00004;
      60482: inst = 32'h38632800;
      60483: inst = 32'h38842800;
      60484: inst = 32'h10a00000;
      60485: inst = 32'hca0ec49;
      60486: inst = 32'h13e00001;
      60487: inst = 32'hfe0d96a;
      60488: inst = 32'h5be00000;
      60489: inst = 32'h8c50000;
      60490: inst = 32'h24612800;
      60491: inst = 32'h10a0ffff;
      60492: inst = 32'hca0fff2;
      60493: inst = 32'h24822800;
      60494: inst = 32'h10a00000;
      60495: inst = 32'hca00004;
      60496: inst = 32'h38632800;
      60497: inst = 32'h38842800;
      60498: inst = 32'h10a00000;
      60499: inst = 32'hca0ec57;
      60500: inst = 32'h13e00001;
      60501: inst = 32'hfe0d96a;
      60502: inst = 32'h5be00000;
      60503: inst = 32'h8c50000;
      60504: inst = 32'h24612800;
      60505: inst = 32'h10a0ffff;
      60506: inst = 32'hca0fff2;
      60507: inst = 32'h24822800;
      60508: inst = 32'h10a00000;
      60509: inst = 32'hca00004;
      60510: inst = 32'h38632800;
      60511: inst = 32'h38842800;
      60512: inst = 32'h10a00000;
      60513: inst = 32'hca0ec65;
      60514: inst = 32'h13e00001;
      60515: inst = 32'hfe0d96a;
      60516: inst = 32'h5be00000;
      60517: inst = 32'h8c50000;
      60518: inst = 32'h24612800;
      60519: inst = 32'h10a0ffff;
      60520: inst = 32'hca0fff2;
      60521: inst = 32'h24822800;
      60522: inst = 32'h10a00000;
      60523: inst = 32'hca00004;
      60524: inst = 32'h38632800;
      60525: inst = 32'h38842800;
      60526: inst = 32'h10a00000;
      60527: inst = 32'hca0ec73;
      60528: inst = 32'h13e00001;
      60529: inst = 32'hfe0d96a;
      60530: inst = 32'h5be00000;
      60531: inst = 32'h8c50000;
      60532: inst = 32'h24612800;
      60533: inst = 32'h10a0ffff;
      60534: inst = 32'hca0fff2;
      60535: inst = 32'h24822800;
      60536: inst = 32'h10a00000;
      60537: inst = 32'hca00004;
      60538: inst = 32'h38632800;
      60539: inst = 32'h38842800;
      60540: inst = 32'h10a00000;
      60541: inst = 32'hca0ec81;
      60542: inst = 32'h13e00001;
      60543: inst = 32'hfe0d96a;
      60544: inst = 32'h5be00000;
      60545: inst = 32'h8c50000;
      60546: inst = 32'h24612800;
      60547: inst = 32'h10a0ffff;
      60548: inst = 32'hca0fff2;
      60549: inst = 32'h24822800;
      60550: inst = 32'h10a00000;
      60551: inst = 32'hca00004;
      60552: inst = 32'h38632800;
      60553: inst = 32'h38842800;
      60554: inst = 32'h10a00000;
      60555: inst = 32'hca0ec8f;
      60556: inst = 32'h13e00001;
      60557: inst = 32'hfe0d96a;
      60558: inst = 32'h5be00000;
      60559: inst = 32'h8c50000;
      60560: inst = 32'h24612800;
      60561: inst = 32'h10a0ffff;
      60562: inst = 32'hca0fff2;
      60563: inst = 32'h24822800;
      60564: inst = 32'h10a00000;
      60565: inst = 32'hca00004;
      60566: inst = 32'h38632800;
      60567: inst = 32'h38842800;
      60568: inst = 32'h10a00000;
      60569: inst = 32'hca0ec9d;
      60570: inst = 32'h13e00001;
      60571: inst = 32'hfe0d96a;
      60572: inst = 32'h5be00000;
      60573: inst = 32'h8c50000;
      60574: inst = 32'h24612800;
      60575: inst = 32'h10a0ffff;
      60576: inst = 32'hca0fff2;
      60577: inst = 32'h24822800;
      60578: inst = 32'h10a00000;
      60579: inst = 32'hca00004;
      60580: inst = 32'h38632800;
      60581: inst = 32'h38842800;
      60582: inst = 32'h10a00000;
      60583: inst = 32'hca0ecab;
      60584: inst = 32'h13e00001;
      60585: inst = 32'hfe0d96a;
      60586: inst = 32'h5be00000;
      60587: inst = 32'h8c50000;
      60588: inst = 32'h24612800;
      60589: inst = 32'h10a0ffff;
      60590: inst = 32'hca0fff2;
      60591: inst = 32'h24822800;
      60592: inst = 32'h10a00000;
      60593: inst = 32'hca00004;
      60594: inst = 32'h38632800;
      60595: inst = 32'h38842800;
      60596: inst = 32'h10a00000;
      60597: inst = 32'hca0ecb9;
      60598: inst = 32'h13e00001;
      60599: inst = 32'hfe0d96a;
      60600: inst = 32'h5be00000;
      60601: inst = 32'h8c50000;
      60602: inst = 32'h24612800;
      60603: inst = 32'h10a0ffff;
      60604: inst = 32'hca0fff2;
      60605: inst = 32'h24822800;
      60606: inst = 32'h10a00000;
      60607: inst = 32'hca00004;
      60608: inst = 32'h38632800;
      60609: inst = 32'h38842800;
      60610: inst = 32'h10a00000;
      60611: inst = 32'hca0ecc7;
      60612: inst = 32'h13e00001;
      60613: inst = 32'hfe0d96a;
      60614: inst = 32'h5be00000;
      60615: inst = 32'h8c50000;
      60616: inst = 32'h24612800;
      60617: inst = 32'h10a0ffff;
      60618: inst = 32'hca0fff2;
      60619: inst = 32'h24822800;
      60620: inst = 32'h10a00000;
      60621: inst = 32'hca00004;
      60622: inst = 32'h38632800;
      60623: inst = 32'h38842800;
      60624: inst = 32'h10a00000;
      60625: inst = 32'hca0ecd5;
      60626: inst = 32'h13e00001;
      60627: inst = 32'hfe0d96a;
      60628: inst = 32'h5be00000;
      60629: inst = 32'h8c50000;
      60630: inst = 32'h24612800;
      60631: inst = 32'h10a0ffff;
      60632: inst = 32'hca0fff2;
      60633: inst = 32'h24822800;
      60634: inst = 32'h10a00000;
      60635: inst = 32'hca00004;
      60636: inst = 32'h38632800;
      60637: inst = 32'h38842800;
      60638: inst = 32'h10a00000;
      60639: inst = 32'hca0ece3;
      60640: inst = 32'h13e00001;
      60641: inst = 32'hfe0d96a;
      60642: inst = 32'h5be00000;
      60643: inst = 32'h8c50000;
      60644: inst = 32'h24612800;
      60645: inst = 32'h10a0ffff;
      60646: inst = 32'hca0fff2;
      60647: inst = 32'h24822800;
      60648: inst = 32'h10a00000;
      60649: inst = 32'hca00004;
      60650: inst = 32'h38632800;
      60651: inst = 32'h38842800;
      60652: inst = 32'h10a00000;
      60653: inst = 32'hca0ecf1;
      60654: inst = 32'h13e00001;
      60655: inst = 32'hfe0d96a;
      60656: inst = 32'h5be00000;
      60657: inst = 32'h8c50000;
      60658: inst = 32'h24612800;
      60659: inst = 32'h10a0ffff;
      60660: inst = 32'hca0fff2;
      60661: inst = 32'h24822800;
      60662: inst = 32'h10a00000;
      60663: inst = 32'hca00004;
      60664: inst = 32'h38632800;
      60665: inst = 32'h38842800;
      60666: inst = 32'h10a00000;
      60667: inst = 32'hca0ecff;
      60668: inst = 32'h13e00001;
      60669: inst = 32'hfe0d96a;
      60670: inst = 32'h5be00000;
      60671: inst = 32'h8c50000;
      60672: inst = 32'h24612800;
      60673: inst = 32'h10a0ffff;
      60674: inst = 32'hca0fff2;
      60675: inst = 32'h24822800;
      60676: inst = 32'h10a00000;
      60677: inst = 32'hca00004;
      60678: inst = 32'h38632800;
      60679: inst = 32'h38842800;
      60680: inst = 32'h10a00000;
      60681: inst = 32'hca0ed0d;
      60682: inst = 32'h13e00001;
      60683: inst = 32'hfe0d96a;
      60684: inst = 32'h5be00000;
      60685: inst = 32'h8c50000;
      60686: inst = 32'h24612800;
      60687: inst = 32'h10a0ffff;
      60688: inst = 32'hca0fff2;
      60689: inst = 32'h24822800;
      60690: inst = 32'h10a00000;
      60691: inst = 32'hca00004;
      60692: inst = 32'h38632800;
      60693: inst = 32'h38842800;
      60694: inst = 32'h10a00000;
      60695: inst = 32'hca0ed1b;
      60696: inst = 32'h13e00001;
      60697: inst = 32'hfe0d96a;
      60698: inst = 32'h5be00000;
      60699: inst = 32'h8c50000;
      60700: inst = 32'h24612800;
      60701: inst = 32'h10a0ffff;
      60702: inst = 32'hca0fff2;
      60703: inst = 32'h24822800;
      60704: inst = 32'h10a00000;
      60705: inst = 32'hca00004;
      60706: inst = 32'h38632800;
      60707: inst = 32'h38842800;
      60708: inst = 32'h10a00000;
      60709: inst = 32'hca0ed29;
      60710: inst = 32'h13e00001;
      60711: inst = 32'hfe0d96a;
      60712: inst = 32'h5be00000;
      60713: inst = 32'h8c50000;
      60714: inst = 32'h24612800;
      60715: inst = 32'h10a0ffff;
      60716: inst = 32'hca0fff3;
      60717: inst = 32'h24822800;
      60718: inst = 32'h10a00000;
      60719: inst = 32'hca00004;
      60720: inst = 32'h38632800;
      60721: inst = 32'h38842800;
      60722: inst = 32'h10a00000;
      60723: inst = 32'hca0ed37;
      60724: inst = 32'h13e00001;
      60725: inst = 32'hfe0d96a;
      60726: inst = 32'h5be00000;
      60727: inst = 32'h8c50000;
      60728: inst = 32'h24612800;
      60729: inst = 32'h10a0ffff;
      60730: inst = 32'hca0fff3;
      60731: inst = 32'h24822800;
      60732: inst = 32'h10a00000;
      60733: inst = 32'hca00004;
      60734: inst = 32'h38632800;
      60735: inst = 32'h38842800;
      60736: inst = 32'h10a00000;
      60737: inst = 32'hca0ed45;
      60738: inst = 32'h13e00001;
      60739: inst = 32'hfe0d96a;
      60740: inst = 32'h5be00000;
      60741: inst = 32'h8c50000;
      60742: inst = 32'h24612800;
      60743: inst = 32'h10a0ffff;
      60744: inst = 32'hca0fff3;
      60745: inst = 32'h24822800;
      60746: inst = 32'h10a00000;
      60747: inst = 32'hca00004;
      60748: inst = 32'h38632800;
      60749: inst = 32'h38842800;
      60750: inst = 32'h10a00000;
      60751: inst = 32'hca0ed53;
      60752: inst = 32'h13e00001;
      60753: inst = 32'hfe0d96a;
      60754: inst = 32'h5be00000;
      60755: inst = 32'h8c50000;
      60756: inst = 32'h24612800;
      60757: inst = 32'h10a0ffff;
      60758: inst = 32'hca0fff3;
      60759: inst = 32'h24822800;
      60760: inst = 32'h10a00000;
      60761: inst = 32'hca00004;
      60762: inst = 32'h38632800;
      60763: inst = 32'h38842800;
      60764: inst = 32'h10a00000;
      60765: inst = 32'hca0ed61;
      60766: inst = 32'h13e00001;
      60767: inst = 32'hfe0d96a;
      60768: inst = 32'h5be00000;
      60769: inst = 32'h8c50000;
      60770: inst = 32'h24612800;
      60771: inst = 32'h10a0ffff;
      60772: inst = 32'hca0fff3;
      60773: inst = 32'h24822800;
      60774: inst = 32'h10a00000;
      60775: inst = 32'hca00004;
      60776: inst = 32'h38632800;
      60777: inst = 32'h38842800;
      60778: inst = 32'h10a00000;
      60779: inst = 32'hca0ed6f;
      60780: inst = 32'h13e00001;
      60781: inst = 32'hfe0d96a;
      60782: inst = 32'h5be00000;
      60783: inst = 32'h8c50000;
      60784: inst = 32'h24612800;
      60785: inst = 32'h10a0ffff;
      60786: inst = 32'hca0fff3;
      60787: inst = 32'h24822800;
      60788: inst = 32'h10a00000;
      60789: inst = 32'hca00004;
      60790: inst = 32'h38632800;
      60791: inst = 32'h38842800;
      60792: inst = 32'h10a00000;
      60793: inst = 32'hca0ed7d;
      60794: inst = 32'h13e00001;
      60795: inst = 32'hfe0d96a;
      60796: inst = 32'h5be00000;
      60797: inst = 32'h8c50000;
      60798: inst = 32'h24612800;
      60799: inst = 32'h10a0ffff;
      60800: inst = 32'hca0fff3;
      60801: inst = 32'h24822800;
      60802: inst = 32'h10a00000;
      60803: inst = 32'hca00004;
      60804: inst = 32'h38632800;
      60805: inst = 32'h38842800;
      60806: inst = 32'h10a00000;
      60807: inst = 32'hca0ed8b;
      60808: inst = 32'h13e00001;
      60809: inst = 32'hfe0d96a;
      60810: inst = 32'h5be00000;
      60811: inst = 32'h8c50000;
      60812: inst = 32'h24612800;
      60813: inst = 32'h10a0ffff;
      60814: inst = 32'hca0fff3;
      60815: inst = 32'h24822800;
      60816: inst = 32'h10a00000;
      60817: inst = 32'hca00004;
      60818: inst = 32'h38632800;
      60819: inst = 32'h38842800;
      60820: inst = 32'h10a00000;
      60821: inst = 32'hca0ed99;
      60822: inst = 32'h13e00001;
      60823: inst = 32'hfe0d96a;
      60824: inst = 32'h5be00000;
      60825: inst = 32'h8c50000;
      60826: inst = 32'h24612800;
      60827: inst = 32'h10a0ffff;
      60828: inst = 32'hca0fff3;
      60829: inst = 32'h24822800;
      60830: inst = 32'h10a00000;
      60831: inst = 32'hca00004;
      60832: inst = 32'h38632800;
      60833: inst = 32'h38842800;
      60834: inst = 32'h10a00000;
      60835: inst = 32'hca0eda7;
      60836: inst = 32'h13e00001;
      60837: inst = 32'hfe0d96a;
      60838: inst = 32'h5be00000;
      60839: inst = 32'h8c50000;
      60840: inst = 32'h24612800;
      60841: inst = 32'h10a0ffff;
      60842: inst = 32'hca0fff3;
      60843: inst = 32'h24822800;
      60844: inst = 32'h10a00000;
      60845: inst = 32'hca00004;
      60846: inst = 32'h38632800;
      60847: inst = 32'h38842800;
      60848: inst = 32'h10a00000;
      60849: inst = 32'hca0edb5;
      60850: inst = 32'h13e00001;
      60851: inst = 32'hfe0d96a;
      60852: inst = 32'h5be00000;
      60853: inst = 32'h8c50000;
      60854: inst = 32'h24612800;
      60855: inst = 32'h10a0ffff;
      60856: inst = 32'hca0fff3;
      60857: inst = 32'h24822800;
      60858: inst = 32'h10a00000;
      60859: inst = 32'hca00004;
      60860: inst = 32'h38632800;
      60861: inst = 32'h38842800;
      60862: inst = 32'h10a00000;
      60863: inst = 32'hca0edc3;
      60864: inst = 32'h13e00001;
      60865: inst = 32'hfe0d96a;
      60866: inst = 32'h5be00000;
      60867: inst = 32'h8c50000;
      60868: inst = 32'h24612800;
      60869: inst = 32'h10a0ffff;
      60870: inst = 32'hca0fff3;
      60871: inst = 32'h24822800;
      60872: inst = 32'h10a00000;
      60873: inst = 32'hca00004;
      60874: inst = 32'h38632800;
      60875: inst = 32'h38842800;
      60876: inst = 32'h10a00000;
      60877: inst = 32'hca0edd1;
      60878: inst = 32'h13e00001;
      60879: inst = 32'hfe0d96a;
      60880: inst = 32'h5be00000;
      60881: inst = 32'h8c50000;
      60882: inst = 32'h24612800;
      60883: inst = 32'h10a0ffff;
      60884: inst = 32'hca0fff3;
      60885: inst = 32'h24822800;
      60886: inst = 32'h10a00000;
      60887: inst = 32'hca00004;
      60888: inst = 32'h38632800;
      60889: inst = 32'h38842800;
      60890: inst = 32'h10a00000;
      60891: inst = 32'hca0eddf;
      60892: inst = 32'h13e00001;
      60893: inst = 32'hfe0d96a;
      60894: inst = 32'h5be00000;
      60895: inst = 32'h8c50000;
      60896: inst = 32'h24612800;
      60897: inst = 32'h10a0ffff;
      60898: inst = 32'hca0fff3;
      60899: inst = 32'h24822800;
      60900: inst = 32'h10a00000;
      60901: inst = 32'hca00004;
      60902: inst = 32'h38632800;
      60903: inst = 32'h38842800;
      60904: inst = 32'h10a00000;
      60905: inst = 32'hca0eded;
      60906: inst = 32'h13e00001;
      60907: inst = 32'hfe0d96a;
      60908: inst = 32'h5be00000;
      60909: inst = 32'h8c50000;
      60910: inst = 32'h24612800;
      60911: inst = 32'h10a0ffff;
      60912: inst = 32'hca0fff3;
      60913: inst = 32'h24822800;
      60914: inst = 32'h10a00000;
      60915: inst = 32'hca00004;
      60916: inst = 32'h38632800;
      60917: inst = 32'h38842800;
      60918: inst = 32'h10a00000;
      60919: inst = 32'hca0edfb;
      60920: inst = 32'h13e00001;
      60921: inst = 32'hfe0d96a;
      60922: inst = 32'h5be00000;
      60923: inst = 32'h8c50000;
      60924: inst = 32'h24612800;
      60925: inst = 32'h10a0ffff;
      60926: inst = 32'hca0fff3;
      60927: inst = 32'h24822800;
      60928: inst = 32'h10a00000;
      60929: inst = 32'hca00004;
      60930: inst = 32'h38632800;
      60931: inst = 32'h38842800;
      60932: inst = 32'h10a00000;
      60933: inst = 32'hca0ee09;
      60934: inst = 32'h13e00001;
      60935: inst = 32'hfe0d96a;
      60936: inst = 32'h5be00000;
      60937: inst = 32'h8c50000;
      60938: inst = 32'h24612800;
      60939: inst = 32'h10a0ffff;
      60940: inst = 32'hca0fff3;
      60941: inst = 32'h24822800;
      60942: inst = 32'h10a00000;
      60943: inst = 32'hca00004;
      60944: inst = 32'h38632800;
      60945: inst = 32'h38842800;
      60946: inst = 32'h10a00000;
      60947: inst = 32'hca0ee17;
      60948: inst = 32'h13e00001;
      60949: inst = 32'hfe0d96a;
      60950: inst = 32'h5be00000;
      60951: inst = 32'h8c50000;
      60952: inst = 32'h24612800;
      60953: inst = 32'h10a0ffff;
      60954: inst = 32'hca0fff3;
      60955: inst = 32'h24822800;
      60956: inst = 32'h10a00000;
      60957: inst = 32'hca00004;
      60958: inst = 32'h38632800;
      60959: inst = 32'h38842800;
      60960: inst = 32'h10a00000;
      60961: inst = 32'hca0ee25;
      60962: inst = 32'h13e00001;
      60963: inst = 32'hfe0d96a;
      60964: inst = 32'h5be00000;
      60965: inst = 32'h8c50000;
      60966: inst = 32'h24612800;
      60967: inst = 32'h10a0ffff;
      60968: inst = 32'hca0fff3;
      60969: inst = 32'h24822800;
      60970: inst = 32'h10a00000;
      60971: inst = 32'hca00004;
      60972: inst = 32'h38632800;
      60973: inst = 32'h38842800;
      60974: inst = 32'h10a00000;
      60975: inst = 32'hca0ee33;
      60976: inst = 32'h13e00001;
      60977: inst = 32'hfe0d96a;
      60978: inst = 32'h5be00000;
      60979: inst = 32'h8c50000;
      60980: inst = 32'h24612800;
      60981: inst = 32'h10a0ffff;
      60982: inst = 32'hca0fff3;
      60983: inst = 32'h24822800;
      60984: inst = 32'h10a00000;
      60985: inst = 32'hca00004;
      60986: inst = 32'h38632800;
      60987: inst = 32'h38842800;
      60988: inst = 32'h10a00000;
      60989: inst = 32'hca0ee41;
      60990: inst = 32'h13e00001;
      60991: inst = 32'hfe0d96a;
      60992: inst = 32'h5be00000;
      60993: inst = 32'h8c50000;
      60994: inst = 32'h24612800;
      60995: inst = 32'h10a0ffff;
      60996: inst = 32'hca0fff3;
      60997: inst = 32'h24822800;
      60998: inst = 32'h10a00000;
      60999: inst = 32'hca00004;
      61000: inst = 32'h38632800;
      61001: inst = 32'h38842800;
      61002: inst = 32'h10a00000;
      61003: inst = 32'hca0ee4f;
      61004: inst = 32'h13e00001;
      61005: inst = 32'hfe0d96a;
      61006: inst = 32'h5be00000;
      61007: inst = 32'h8c50000;
      61008: inst = 32'h24612800;
      61009: inst = 32'h10a0ffff;
      61010: inst = 32'hca0fff3;
      61011: inst = 32'h24822800;
      61012: inst = 32'h10a00000;
      61013: inst = 32'hca00004;
      61014: inst = 32'h38632800;
      61015: inst = 32'h38842800;
      61016: inst = 32'h10a00000;
      61017: inst = 32'hca0ee5d;
      61018: inst = 32'h13e00001;
      61019: inst = 32'hfe0d96a;
      61020: inst = 32'h5be00000;
      61021: inst = 32'h8c50000;
      61022: inst = 32'h24612800;
      61023: inst = 32'h10a0ffff;
      61024: inst = 32'hca0fff3;
      61025: inst = 32'h24822800;
      61026: inst = 32'h10a00000;
      61027: inst = 32'hca00004;
      61028: inst = 32'h38632800;
      61029: inst = 32'h38842800;
      61030: inst = 32'h10a00000;
      61031: inst = 32'hca0ee6b;
      61032: inst = 32'h13e00001;
      61033: inst = 32'hfe0d96a;
      61034: inst = 32'h5be00000;
      61035: inst = 32'h8c50000;
      61036: inst = 32'h24612800;
      61037: inst = 32'h10a0ffff;
      61038: inst = 32'hca0fff3;
      61039: inst = 32'h24822800;
      61040: inst = 32'h10a00000;
      61041: inst = 32'hca00004;
      61042: inst = 32'h38632800;
      61043: inst = 32'h38842800;
      61044: inst = 32'h10a00000;
      61045: inst = 32'hca0ee79;
      61046: inst = 32'h13e00001;
      61047: inst = 32'hfe0d96a;
      61048: inst = 32'h5be00000;
      61049: inst = 32'h8c50000;
      61050: inst = 32'h24612800;
      61051: inst = 32'h10a0ffff;
      61052: inst = 32'hca0fff3;
      61053: inst = 32'h24822800;
      61054: inst = 32'h10a00000;
      61055: inst = 32'hca00004;
      61056: inst = 32'h38632800;
      61057: inst = 32'h38842800;
      61058: inst = 32'h10a00000;
      61059: inst = 32'hca0ee87;
      61060: inst = 32'h13e00001;
      61061: inst = 32'hfe0d96a;
      61062: inst = 32'h5be00000;
      61063: inst = 32'h8c50000;
      61064: inst = 32'h24612800;
      61065: inst = 32'h10a0ffff;
      61066: inst = 32'hca0fff3;
      61067: inst = 32'h24822800;
      61068: inst = 32'h10a00000;
      61069: inst = 32'hca00004;
      61070: inst = 32'h38632800;
      61071: inst = 32'h38842800;
      61072: inst = 32'h10a00000;
      61073: inst = 32'hca0ee95;
      61074: inst = 32'h13e00001;
      61075: inst = 32'hfe0d96a;
      61076: inst = 32'h5be00000;
      61077: inst = 32'h8c50000;
      61078: inst = 32'h24612800;
      61079: inst = 32'h10a0ffff;
      61080: inst = 32'hca0fff3;
      61081: inst = 32'h24822800;
      61082: inst = 32'h10a00000;
      61083: inst = 32'hca00004;
      61084: inst = 32'h38632800;
      61085: inst = 32'h38842800;
      61086: inst = 32'h10a00000;
      61087: inst = 32'hca0eea3;
      61088: inst = 32'h13e00001;
      61089: inst = 32'hfe0d96a;
      61090: inst = 32'h5be00000;
      61091: inst = 32'h8c50000;
      61092: inst = 32'h24612800;
      61093: inst = 32'h10a0ffff;
      61094: inst = 32'hca0fff3;
      61095: inst = 32'h24822800;
      61096: inst = 32'h10a00000;
      61097: inst = 32'hca00004;
      61098: inst = 32'h38632800;
      61099: inst = 32'h38842800;
      61100: inst = 32'h10a00000;
      61101: inst = 32'hca0eeb1;
      61102: inst = 32'h13e00001;
      61103: inst = 32'hfe0d96a;
      61104: inst = 32'h5be00000;
      61105: inst = 32'h8c50000;
      61106: inst = 32'h24612800;
      61107: inst = 32'h10a0ffff;
      61108: inst = 32'hca0fff3;
      61109: inst = 32'h24822800;
      61110: inst = 32'h10a00000;
      61111: inst = 32'hca00004;
      61112: inst = 32'h38632800;
      61113: inst = 32'h38842800;
      61114: inst = 32'h10a00000;
      61115: inst = 32'hca0eebf;
      61116: inst = 32'h13e00001;
      61117: inst = 32'hfe0d96a;
      61118: inst = 32'h5be00000;
      61119: inst = 32'h8c50000;
      61120: inst = 32'h24612800;
      61121: inst = 32'h10a0ffff;
      61122: inst = 32'hca0fff3;
      61123: inst = 32'h24822800;
      61124: inst = 32'h10a00000;
      61125: inst = 32'hca00004;
      61126: inst = 32'h38632800;
      61127: inst = 32'h38842800;
      61128: inst = 32'h10a00000;
      61129: inst = 32'hca0eecd;
      61130: inst = 32'h13e00001;
      61131: inst = 32'hfe0d96a;
      61132: inst = 32'h5be00000;
      61133: inst = 32'h8c50000;
      61134: inst = 32'h24612800;
      61135: inst = 32'h10a0ffff;
      61136: inst = 32'hca0fff3;
      61137: inst = 32'h24822800;
      61138: inst = 32'h10a00000;
      61139: inst = 32'hca00004;
      61140: inst = 32'h38632800;
      61141: inst = 32'h38842800;
      61142: inst = 32'h10a00000;
      61143: inst = 32'hca0eedb;
      61144: inst = 32'h13e00001;
      61145: inst = 32'hfe0d96a;
      61146: inst = 32'h5be00000;
      61147: inst = 32'h8c50000;
      61148: inst = 32'h24612800;
      61149: inst = 32'h10a0ffff;
      61150: inst = 32'hca0fff3;
      61151: inst = 32'h24822800;
      61152: inst = 32'h10a00000;
      61153: inst = 32'hca00004;
      61154: inst = 32'h38632800;
      61155: inst = 32'h38842800;
      61156: inst = 32'h10a00000;
      61157: inst = 32'hca0eee9;
      61158: inst = 32'h13e00001;
      61159: inst = 32'hfe0d96a;
      61160: inst = 32'h5be00000;
      61161: inst = 32'h8c50000;
      61162: inst = 32'h24612800;
      61163: inst = 32'h10a0ffff;
      61164: inst = 32'hca0fff3;
      61165: inst = 32'h24822800;
      61166: inst = 32'h10a00000;
      61167: inst = 32'hca00004;
      61168: inst = 32'h38632800;
      61169: inst = 32'h38842800;
      61170: inst = 32'h10a00000;
      61171: inst = 32'hca0eef7;
      61172: inst = 32'h13e00001;
      61173: inst = 32'hfe0d96a;
      61174: inst = 32'h5be00000;
      61175: inst = 32'h8c50000;
      61176: inst = 32'h24612800;
      61177: inst = 32'h10a0ffff;
      61178: inst = 32'hca0fff3;
      61179: inst = 32'h24822800;
      61180: inst = 32'h10a00000;
      61181: inst = 32'hca00004;
      61182: inst = 32'h38632800;
      61183: inst = 32'h38842800;
      61184: inst = 32'h10a00000;
      61185: inst = 32'hca0ef05;
      61186: inst = 32'h13e00001;
      61187: inst = 32'hfe0d96a;
      61188: inst = 32'h5be00000;
      61189: inst = 32'h8c50000;
      61190: inst = 32'h24612800;
      61191: inst = 32'h10a0ffff;
      61192: inst = 32'hca0fff3;
      61193: inst = 32'h24822800;
      61194: inst = 32'h10a00000;
      61195: inst = 32'hca00004;
      61196: inst = 32'h38632800;
      61197: inst = 32'h38842800;
      61198: inst = 32'h10a00000;
      61199: inst = 32'hca0ef13;
      61200: inst = 32'h13e00001;
      61201: inst = 32'hfe0d96a;
      61202: inst = 32'h5be00000;
      61203: inst = 32'h8c50000;
      61204: inst = 32'h24612800;
      61205: inst = 32'h10a0ffff;
      61206: inst = 32'hca0fff3;
      61207: inst = 32'h24822800;
      61208: inst = 32'h10a00000;
      61209: inst = 32'hca00004;
      61210: inst = 32'h38632800;
      61211: inst = 32'h38842800;
      61212: inst = 32'h10a00000;
      61213: inst = 32'hca0ef21;
      61214: inst = 32'h13e00001;
      61215: inst = 32'hfe0d96a;
      61216: inst = 32'h5be00000;
      61217: inst = 32'h8c50000;
      61218: inst = 32'h24612800;
      61219: inst = 32'h10a0ffff;
      61220: inst = 32'hca0fff3;
      61221: inst = 32'h24822800;
      61222: inst = 32'h10a00000;
      61223: inst = 32'hca00004;
      61224: inst = 32'h38632800;
      61225: inst = 32'h38842800;
      61226: inst = 32'h10a00000;
      61227: inst = 32'hca0ef2f;
      61228: inst = 32'h13e00001;
      61229: inst = 32'hfe0d96a;
      61230: inst = 32'h5be00000;
      61231: inst = 32'h8c50000;
      61232: inst = 32'h24612800;
      61233: inst = 32'h10a0ffff;
      61234: inst = 32'hca0fff3;
      61235: inst = 32'h24822800;
      61236: inst = 32'h10a00000;
      61237: inst = 32'hca00004;
      61238: inst = 32'h38632800;
      61239: inst = 32'h38842800;
      61240: inst = 32'h10a00000;
      61241: inst = 32'hca0ef3d;
      61242: inst = 32'h13e00001;
      61243: inst = 32'hfe0d96a;
      61244: inst = 32'h5be00000;
      61245: inst = 32'h8c50000;
      61246: inst = 32'h24612800;
      61247: inst = 32'h10a0ffff;
      61248: inst = 32'hca0fff3;
      61249: inst = 32'h24822800;
      61250: inst = 32'h10a00000;
      61251: inst = 32'hca00004;
      61252: inst = 32'h38632800;
      61253: inst = 32'h38842800;
      61254: inst = 32'h10a00000;
      61255: inst = 32'hca0ef4b;
      61256: inst = 32'h13e00001;
      61257: inst = 32'hfe0d96a;
      61258: inst = 32'h5be00000;
      61259: inst = 32'h8c50000;
      61260: inst = 32'h24612800;
      61261: inst = 32'h10a0ffff;
      61262: inst = 32'hca0fff3;
      61263: inst = 32'h24822800;
      61264: inst = 32'h10a00000;
      61265: inst = 32'hca00004;
      61266: inst = 32'h38632800;
      61267: inst = 32'h38842800;
      61268: inst = 32'h10a00000;
      61269: inst = 32'hca0ef59;
      61270: inst = 32'h13e00001;
      61271: inst = 32'hfe0d96a;
      61272: inst = 32'h5be00000;
      61273: inst = 32'h8c50000;
      61274: inst = 32'h24612800;
      61275: inst = 32'h10a0ffff;
      61276: inst = 32'hca0fff3;
      61277: inst = 32'h24822800;
      61278: inst = 32'h10a00000;
      61279: inst = 32'hca00004;
      61280: inst = 32'h38632800;
      61281: inst = 32'h38842800;
      61282: inst = 32'h10a00000;
      61283: inst = 32'hca0ef67;
      61284: inst = 32'h13e00001;
      61285: inst = 32'hfe0d96a;
      61286: inst = 32'h5be00000;
      61287: inst = 32'h8c50000;
      61288: inst = 32'h24612800;
      61289: inst = 32'h10a0ffff;
      61290: inst = 32'hca0fff3;
      61291: inst = 32'h24822800;
      61292: inst = 32'h10a00000;
      61293: inst = 32'hca00004;
      61294: inst = 32'h38632800;
      61295: inst = 32'h38842800;
      61296: inst = 32'h10a00000;
      61297: inst = 32'hca0ef75;
      61298: inst = 32'h13e00001;
      61299: inst = 32'hfe0d96a;
      61300: inst = 32'h5be00000;
      61301: inst = 32'h8c50000;
      61302: inst = 32'h24612800;
      61303: inst = 32'h10a0ffff;
      61304: inst = 32'hca0fff3;
      61305: inst = 32'h24822800;
      61306: inst = 32'h10a00000;
      61307: inst = 32'hca00004;
      61308: inst = 32'h38632800;
      61309: inst = 32'h38842800;
      61310: inst = 32'h10a00000;
      61311: inst = 32'hca0ef83;
      61312: inst = 32'h13e00001;
      61313: inst = 32'hfe0d96a;
      61314: inst = 32'h5be00000;
      61315: inst = 32'h8c50000;
      61316: inst = 32'h24612800;
      61317: inst = 32'h10a0ffff;
      61318: inst = 32'hca0fff3;
      61319: inst = 32'h24822800;
      61320: inst = 32'h10a00000;
      61321: inst = 32'hca00004;
      61322: inst = 32'h38632800;
      61323: inst = 32'h38842800;
      61324: inst = 32'h10a00000;
      61325: inst = 32'hca0ef91;
      61326: inst = 32'h13e00001;
      61327: inst = 32'hfe0d96a;
      61328: inst = 32'h5be00000;
      61329: inst = 32'h8c50000;
      61330: inst = 32'h24612800;
      61331: inst = 32'h10a0ffff;
      61332: inst = 32'hca0fff3;
      61333: inst = 32'h24822800;
      61334: inst = 32'h10a00000;
      61335: inst = 32'hca00004;
      61336: inst = 32'h38632800;
      61337: inst = 32'h38842800;
      61338: inst = 32'h10a00000;
      61339: inst = 32'hca0ef9f;
      61340: inst = 32'h13e00001;
      61341: inst = 32'hfe0d96a;
      61342: inst = 32'h5be00000;
      61343: inst = 32'h8c50000;
      61344: inst = 32'h24612800;
      61345: inst = 32'h10a0ffff;
      61346: inst = 32'hca0fff3;
      61347: inst = 32'h24822800;
      61348: inst = 32'h10a00000;
      61349: inst = 32'hca00004;
      61350: inst = 32'h38632800;
      61351: inst = 32'h38842800;
      61352: inst = 32'h10a00000;
      61353: inst = 32'hca0efad;
      61354: inst = 32'h13e00001;
      61355: inst = 32'hfe0d96a;
      61356: inst = 32'h5be00000;
      61357: inst = 32'h8c50000;
      61358: inst = 32'h24612800;
      61359: inst = 32'h10a0ffff;
      61360: inst = 32'hca0fff3;
      61361: inst = 32'h24822800;
      61362: inst = 32'h10a00000;
      61363: inst = 32'hca00004;
      61364: inst = 32'h38632800;
      61365: inst = 32'h38842800;
      61366: inst = 32'h10a00000;
      61367: inst = 32'hca0efbb;
      61368: inst = 32'h13e00001;
      61369: inst = 32'hfe0d96a;
      61370: inst = 32'h5be00000;
      61371: inst = 32'h8c50000;
      61372: inst = 32'h24612800;
      61373: inst = 32'h10a0ffff;
      61374: inst = 32'hca0fff3;
      61375: inst = 32'h24822800;
      61376: inst = 32'h10a00000;
      61377: inst = 32'hca00004;
      61378: inst = 32'h38632800;
      61379: inst = 32'h38842800;
      61380: inst = 32'h10a00000;
      61381: inst = 32'hca0efc9;
      61382: inst = 32'h13e00001;
      61383: inst = 32'hfe0d96a;
      61384: inst = 32'h5be00000;
      61385: inst = 32'h8c50000;
      61386: inst = 32'h24612800;
      61387: inst = 32'h10a0ffff;
      61388: inst = 32'hca0fff3;
      61389: inst = 32'h24822800;
      61390: inst = 32'h10a00000;
      61391: inst = 32'hca00004;
      61392: inst = 32'h38632800;
      61393: inst = 32'h38842800;
      61394: inst = 32'h10a00000;
      61395: inst = 32'hca0efd7;
      61396: inst = 32'h13e00001;
      61397: inst = 32'hfe0d96a;
      61398: inst = 32'h5be00000;
      61399: inst = 32'h8c50000;
      61400: inst = 32'h24612800;
      61401: inst = 32'h10a0ffff;
      61402: inst = 32'hca0fff3;
      61403: inst = 32'h24822800;
      61404: inst = 32'h10a00000;
      61405: inst = 32'hca00004;
      61406: inst = 32'h38632800;
      61407: inst = 32'h38842800;
      61408: inst = 32'h10a00000;
      61409: inst = 32'hca0efe5;
      61410: inst = 32'h13e00001;
      61411: inst = 32'hfe0d96a;
      61412: inst = 32'h5be00000;
      61413: inst = 32'h8c50000;
      61414: inst = 32'h24612800;
      61415: inst = 32'h10a0ffff;
      61416: inst = 32'hca0fff3;
      61417: inst = 32'h24822800;
      61418: inst = 32'h10a00000;
      61419: inst = 32'hca00004;
      61420: inst = 32'h38632800;
      61421: inst = 32'h38842800;
      61422: inst = 32'h10a00000;
      61423: inst = 32'hca0eff3;
      61424: inst = 32'h13e00001;
      61425: inst = 32'hfe0d96a;
      61426: inst = 32'h5be00000;
      61427: inst = 32'h8c50000;
      61428: inst = 32'h24612800;
      61429: inst = 32'h10a0ffff;
      61430: inst = 32'hca0fff3;
      61431: inst = 32'h24822800;
      61432: inst = 32'h10a00000;
      61433: inst = 32'hca00004;
      61434: inst = 32'h38632800;
      61435: inst = 32'h38842800;
      61436: inst = 32'h10a00000;
      61437: inst = 32'hca0f001;
      61438: inst = 32'h13e00001;
      61439: inst = 32'hfe0d96a;
      61440: inst = 32'h5be00000;
      61441: inst = 32'h8c50000;
      61442: inst = 32'h24612800;
      61443: inst = 32'h10a0ffff;
      61444: inst = 32'hca0fff3;
      61445: inst = 32'h24822800;
      61446: inst = 32'h10a00000;
      61447: inst = 32'hca00004;
      61448: inst = 32'h38632800;
      61449: inst = 32'h38842800;
      61450: inst = 32'h10a00000;
      61451: inst = 32'hca0f00f;
      61452: inst = 32'h13e00001;
      61453: inst = 32'hfe0d96a;
      61454: inst = 32'h5be00000;
      61455: inst = 32'h8c50000;
      61456: inst = 32'h24612800;
      61457: inst = 32'h10a0ffff;
      61458: inst = 32'hca0fff3;
      61459: inst = 32'h24822800;
      61460: inst = 32'h10a00000;
      61461: inst = 32'hca00004;
      61462: inst = 32'h38632800;
      61463: inst = 32'h38842800;
      61464: inst = 32'h10a00000;
      61465: inst = 32'hca0f01d;
      61466: inst = 32'h13e00001;
      61467: inst = 32'hfe0d96a;
      61468: inst = 32'h5be00000;
      61469: inst = 32'h8c50000;
      61470: inst = 32'h24612800;
      61471: inst = 32'h10a0ffff;
      61472: inst = 32'hca0fff3;
      61473: inst = 32'h24822800;
      61474: inst = 32'h10a00000;
      61475: inst = 32'hca00004;
      61476: inst = 32'h38632800;
      61477: inst = 32'h38842800;
      61478: inst = 32'h10a00000;
      61479: inst = 32'hca0f02b;
      61480: inst = 32'h13e00001;
      61481: inst = 32'hfe0d96a;
      61482: inst = 32'h5be00000;
      61483: inst = 32'h8c50000;
      61484: inst = 32'h24612800;
      61485: inst = 32'h10a0ffff;
      61486: inst = 32'hca0fff3;
      61487: inst = 32'h24822800;
      61488: inst = 32'h10a00000;
      61489: inst = 32'hca00004;
      61490: inst = 32'h38632800;
      61491: inst = 32'h38842800;
      61492: inst = 32'h10a00000;
      61493: inst = 32'hca0f039;
      61494: inst = 32'h13e00001;
      61495: inst = 32'hfe0d96a;
      61496: inst = 32'h5be00000;
      61497: inst = 32'h8c50000;
      61498: inst = 32'h24612800;
      61499: inst = 32'h10a0ffff;
      61500: inst = 32'hca0fff3;
      61501: inst = 32'h24822800;
      61502: inst = 32'h10a00000;
      61503: inst = 32'hca00004;
      61504: inst = 32'h38632800;
      61505: inst = 32'h38842800;
      61506: inst = 32'h10a00000;
      61507: inst = 32'hca0f047;
      61508: inst = 32'h13e00001;
      61509: inst = 32'hfe0d96a;
      61510: inst = 32'h5be00000;
      61511: inst = 32'h8c50000;
      61512: inst = 32'h24612800;
      61513: inst = 32'h10a0ffff;
      61514: inst = 32'hca0fff3;
      61515: inst = 32'h24822800;
      61516: inst = 32'h10a00000;
      61517: inst = 32'hca00004;
      61518: inst = 32'h38632800;
      61519: inst = 32'h38842800;
      61520: inst = 32'h10a00000;
      61521: inst = 32'hca0f055;
      61522: inst = 32'h13e00001;
      61523: inst = 32'hfe0d96a;
      61524: inst = 32'h5be00000;
      61525: inst = 32'h8c50000;
      61526: inst = 32'h24612800;
      61527: inst = 32'h10a0ffff;
      61528: inst = 32'hca0fff3;
      61529: inst = 32'h24822800;
      61530: inst = 32'h10a00000;
      61531: inst = 32'hca00004;
      61532: inst = 32'h38632800;
      61533: inst = 32'h38842800;
      61534: inst = 32'h10a00000;
      61535: inst = 32'hca0f063;
      61536: inst = 32'h13e00001;
      61537: inst = 32'hfe0d96a;
      61538: inst = 32'h5be00000;
      61539: inst = 32'h8c50000;
      61540: inst = 32'h24612800;
      61541: inst = 32'h10a0ffff;
      61542: inst = 32'hca0fff3;
      61543: inst = 32'h24822800;
      61544: inst = 32'h10a00000;
      61545: inst = 32'hca00004;
      61546: inst = 32'h38632800;
      61547: inst = 32'h38842800;
      61548: inst = 32'h10a00000;
      61549: inst = 32'hca0f071;
      61550: inst = 32'h13e00001;
      61551: inst = 32'hfe0d96a;
      61552: inst = 32'h5be00000;
      61553: inst = 32'h8c50000;
      61554: inst = 32'h24612800;
      61555: inst = 32'h10a0ffff;
      61556: inst = 32'hca0fff3;
      61557: inst = 32'h24822800;
      61558: inst = 32'h10a00000;
      61559: inst = 32'hca00004;
      61560: inst = 32'h38632800;
      61561: inst = 32'h38842800;
      61562: inst = 32'h10a00000;
      61563: inst = 32'hca0f07f;
      61564: inst = 32'h13e00001;
      61565: inst = 32'hfe0d96a;
      61566: inst = 32'h5be00000;
      61567: inst = 32'h8c50000;
      61568: inst = 32'h24612800;
      61569: inst = 32'h10a0ffff;
      61570: inst = 32'hca0fff3;
      61571: inst = 32'h24822800;
      61572: inst = 32'h10a00000;
      61573: inst = 32'hca00004;
      61574: inst = 32'h38632800;
      61575: inst = 32'h38842800;
      61576: inst = 32'h10a00000;
      61577: inst = 32'hca0f08d;
      61578: inst = 32'h13e00001;
      61579: inst = 32'hfe0d96a;
      61580: inst = 32'h5be00000;
      61581: inst = 32'h8c50000;
      61582: inst = 32'h24612800;
      61583: inst = 32'h10a0ffff;
      61584: inst = 32'hca0fff3;
      61585: inst = 32'h24822800;
      61586: inst = 32'h10a00000;
      61587: inst = 32'hca00004;
      61588: inst = 32'h38632800;
      61589: inst = 32'h38842800;
      61590: inst = 32'h10a00000;
      61591: inst = 32'hca0f09b;
      61592: inst = 32'h13e00001;
      61593: inst = 32'hfe0d96a;
      61594: inst = 32'h5be00000;
      61595: inst = 32'h8c50000;
      61596: inst = 32'h24612800;
      61597: inst = 32'h10a0ffff;
      61598: inst = 32'hca0fff3;
      61599: inst = 32'h24822800;
      61600: inst = 32'h10a00000;
      61601: inst = 32'hca00004;
      61602: inst = 32'h38632800;
      61603: inst = 32'h38842800;
      61604: inst = 32'h10a00000;
      61605: inst = 32'hca0f0a9;
      61606: inst = 32'h13e00001;
      61607: inst = 32'hfe0d96a;
      61608: inst = 32'h5be00000;
      61609: inst = 32'h8c50000;
      61610: inst = 32'h24612800;
      61611: inst = 32'h10a0ffff;
      61612: inst = 32'hca0fff3;
      61613: inst = 32'h24822800;
      61614: inst = 32'h10a00000;
      61615: inst = 32'hca00004;
      61616: inst = 32'h38632800;
      61617: inst = 32'h38842800;
      61618: inst = 32'h10a00000;
      61619: inst = 32'hca0f0b7;
      61620: inst = 32'h13e00001;
      61621: inst = 32'hfe0d96a;
      61622: inst = 32'h5be00000;
      61623: inst = 32'h8c50000;
      61624: inst = 32'h24612800;
      61625: inst = 32'h10a0ffff;
      61626: inst = 32'hca0fff3;
      61627: inst = 32'h24822800;
      61628: inst = 32'h10a00000;
      61629: inst = 32'hca00004;
      61630: inst = 32'h38632800;
      61631: inst = 32'h38842800;
      61632: inst = 32'h10a00000;
      61633: inst = 32'hca0f0c5;
      61634: inst = 32'h13e00001;
      61635: inst = 32'hfe0d96a;
      61636: inst = 32'h5be00000;
      61637: inst = 32'h8c50000;
      61638: inst = 32'h24612800;
      61639: inst = 32'h10a0ffff;
      61640: inst = 32'hca0fff3;
      61641: inst = 32'h24822800;
      61642: inst = 32'h10a00000;
      61643: inst = 32'hca00004;
      61644: inst = 32'h38632800;
      61645: inst = 32'h38842800;
      61646: inst = 32'h10a00000;
      61647: inst = 32'hca0f0d3;
      61648: inst = 32'h13e00001;
      61649: inst = 32'hfe0d96a;
      61650: inst = 32'h5be00000;
      61651: inst = 32'h8c50000;
      61652: inst = 32'h24612800;
      61653: inst = 32'h10a0ffff;
      61654: inst = 32'hca0fff3;
      61655: inst = 32'h24822800;
      61656: inst = 32'h10a00000;
      61657: inst = 32'hca00004;
      61658: inst = 32'h38632800;
      61659: inst = 32'h38842800;
      61660: inst = 32'h10a00000;
      61661: inst = 32'hca0f0e1;
      61662: inst = 32'h13e00001;
      61663: inst = 32'hfe0d96a;
      61664: inst = 32'h5be00000;
      61665: inst = 32'h8c50000;
      61666: inst = 32'h24612800;
      61667: inst = 32'h10a0ffff;
      61668: inst = 32'hca0fff3;
      61669: inst = 32'h24822800;
      61670: inst = 32'h10a00000;
      61671: inst = 32'hca00004;
      61672: inst = 32'h38632800;
      61673: inst = 32'h38842800;
      61674: inst = 32'h10a00000;
      61675: inst = 32'hca0f0ef;
      61676: inst = 32'h13e00001;
      61677: inst = 32'hfe0d96a;
      61678: inst = 32'h5be00000;
      61679: inst = 32'h8c50000;
      61680: inst = 32'h24612800;
      61681: inst = 32'h10a0ffff;
      61682: inst = 32'hca0fff3;
      61683: inst = 32'h24822800;
      61684: inst = 32'h10a00000;
      61685: inst = 32'hca00004;
      61686: inst = 32'h38632800;
      61687: inst = 32'h38842800;
      61688: inst = 32'h10a00000;
      61689: inst = 32'hca0f0fd;
      61690: inst = 32'h13e00001;
      61691: inst = 32'hfe0d96a;
      61692: inst = 32'h5be00000;
      61693: inst = 32'h8c50000;
      61694: inst = 32'h24612800;
      61695: inst = 32'h10a0ffff;
      61696: inst = 32'hca0fff3;
      61697: inst = 32'h24822800;
      61698: inst = 32'h10a00000;
      61699: inst = 32'hca00004;
      61700: inst = 32'h38632800;
      61701: inst = 32'h38842800;
      61702: inst = 32'h10a00000;
      61703: inst = 32'hca0f10b;
      61704: inst = 32'h13e00001;
      61705: inst = 32'hfe0d96a;
      61706: inst = 32'h5be00000;
      61707: inst = 32'h8c50000;
      61708: inst = 32'h24612800;
      61709: inst = 32'h10a0ffff;
      61710: inst = 32'hca0fff3;
      61711: inst = 32'h24822800;
      61712: inst = 32'h10a00000;
      61713: inst = 32'hca00004;
      61714: inst = 32'h38632800;
      61715: inst = 32'h38842800;
      61716: inst = 32'h10a00000;
      61717: inst = 32'hca0f119;
      61718: inst = 32'h13e00001;
      61719: inst = 32'hfe0d96a;
      61720: inst = 32'h5be00000;
      61721: inst = 32'h8c50000;
      61722: inst = 32'h24612800;
      61723: inst = 32'h10a0ffff;
      61724: inst = 32'hca0fff3;
      61725: inst = 32'h24822800;
      61726: inst = 32'h10a00000;
      61727: inst = 32'hca00004;
      61728: inst = 32'h38632800;
      61729: inst = 32'h38842800;
      61730: inst = 32'h10a00000;
      61731: inst = 32'hca0f127;
      61732: inst = 32'h13e00001;
      61733: inst = 32'hfe0d96a;
      61734: inst = 32'h5be00000;
      61735: inst = 32'h8c50000;
      61736: inst = 32'h24612800;
      61737: inst = 32'h10a0ffff;
      61738: inst = 32'hca0fff3;
      61739: inst = 32'h24822800;
      61740: inst = 32'h10a00000;
      61741: inst = 32'hca00004;
      61742: inst = 32'h38632800;
      61743: inst = 32'h38842800;
      61744: inst = 32'h10a00000;
      61745: inst = 32'hca0f135;
      61746: inst = 32'h13e00001;
      61747: inst = 32'hfe0d96a;
      61748: inst = 32'h5be00000;
      61749: inst = 32'h8c50000;
      61750: inst = 32'h24612800;
      61751: inst = 32'h10a0ffff;
      61752: inst = 32'hca0fff3;
      61753: inst = 32'h24822800;
      61754: inst = 32'h10a00000;
      61755: inst = 32'hca00004;
      61756: inst = 32'h38632800;
      61757: inst = 32'h38842800;
      61758: inst = 32'h10a00000;
      61759: inst = 32'hca0f143;
      61760: inst = 32'h13e00001;
      61761: inst = 32'hfe0d96a;
      61762: inst = 32'h5be00000;
      61763: inst = 32'h8c50000;
      61764: inst = 32'h24612800;
      61765: inst = 32'h10a0ffff;
      61766: inst = 32'hca0fff3;
      61767: inst = 32'h24822800;
      61768: inst = 32'h10a00000;
      61769: inst = 32'hca00004;
      61770: inst = 32'h38632800;
      61771: inst = 32'h38842800;
      61772: inst = 32'h10a00000;
      61773: inst = 32'hca0f151;
      61774: inst = 32'h13e00001;
      61775: inst = 32'hfe0d96a;
      61776: inst = 32'h5be00000;
      61777: inst = 32'h8c50000;
      61778: inst = 32'h24612800;
      61779: inst = 32'h10a0ffff;
      61780: inst = 32'hca0fff3;
      61781: inst = 32'h24822800;
      61782: inst = 32'h10a00000;
      61783: inst = 32'hca00004;
      61784: inst = 32'h38632800;
      61785: inst = 32'h38842800;
      61786: inst = 32'h10a00000;
      61787: inst = 32'hca0f15f;
      61788: inst = 32'h13e00001;
      61789: inst = 32'hfe0d96a;
      61790: inst = 32'h5be00000;
      61791: inst = 32'h8c50000;
      61792: inst = 32'h24612800;
      61793: inst = 32'h10a0ffff;
      61794: inst = 32'hca0fff3;
      61795: inst = 32'h24822800;
      61796: inst = 32'h10a00000;
      61797: inst = 32'hca00004;
      61798: inst = 32'h38632800;
      61799: inst = 32'h38842800;
      61800: inst = 32'h10a00000;
      61801: inst = 32'hca0f16d;
      61802: inst = 32'h13e00001;
      61803: inst = 32'hfe0d96a;
      61804: inst = 32'h5be00000;
      61805: inst = 32'h8c50000;
      61806: inst = 32'h24612800;
      61807: inst = 32'h10a0ffff;
      61808: inst = 32'hca0fff3;
      61809: inst = 32'h24822800;
      61810: inst = 32'h10a00000;
      61811: inst = 32'hca00004;
      61812: inst = 32'h38632800;
      61813: inst = 32'h38842800;
      61814: inst = 32'h10a00000;
      61815: inst = 32'hca0f17b;
      61816: inst = 32'h13e00001;
      61817: inst = 32'hfe0d96a;
      61818: inst = 32'h5be00000;
      61819: inst = 32'h8c50000;
      61820: inst = 32'h24612800;
      61821: inst = 32'h10a0ffff;
      61822: inst = 32'hca0fff3;
      61823: inst = 32'h24822800;
      61824: inst = 32'h10a00000;
      61825: inst = 32'hca00004;
      61826: inst = 32'h38632800;
      61827: inst = 32'h38842800;
      61828: inst = 32'h10a00000;
      61829: inst = 32'hca0f189;
      61830: inst = 32'h13e00001;
      61831: inst = 32'hfe0d96a;
      61832: inst = 32'h5be00000;
      61833: inst = 32'h8c50000;
      61834: inst = 32'h24612800;
      61835: inst = 32'h10a0ffff;
      61836: inst = 32'hca0fff3;
      61837: inst = 32'h24822800;
      61838: inst = 32'h10a00000;
      61839: inst = 32'hca00004;
      61840: inst = 32'h38632800;
      61841: inst = 32'h38842800;
      61842: inst = 32'h10a00000;
      61843: inst = 32'hca0f197;
      61844: inst = 32'h13e00001;
      61845: inst = 32'hfe0d96a;
      61846: inst = 32'h5be00000;
      61847: inst = 32'h8c50000;
      61848: inst = 32'h24612800;
      61849: inst = 32'h10a0ffff;
      61850: inst = 32'hca0fff3;
      61851: inst = 32'h24822800;
      61852: inst = 32'h10a00000;
      61853: inst = 32'hca00004;
      61854: inst = 32'h38632800;
      61855: inst = 32'h38842800;
      61856: inst = 32'h10a00000;
      61857: inst = 32'hca0f1a5;
      61858: inst = 32'h13e00001;
      61859: inst = 32'hfe0d96a;
      61860: inst = 32'h5be00000;
      61861: inst = 32'h8c50000;
      61862: inst = 32'h24612800;
      61863: inst = 32'h10a0ffff;
      61864: inst = 32'hca0fff3;
      61865: inst = 32'h24822800;
      61866: inst = 32'h10a00000;
      61867: inst = 32'hca00004;
      61868: inst = 32'h38632800;
      61869: inst = 32'h38842800;
      61870: inst = 32'h10a00000;
      61871: inst = 32'hca0f1b3;
      61872: inst = 32'h13e00001;
      61873: inst = 32'hfe0d96a;
      61874: inst = 32'h5be00000;
      61875: inst = 32'h8c50000;
      61876: inst = 32'h24612800;
      61877: inst = 32'h10a0ffff;
      61878: inst = 32'hca0fff3;
      61879: inst = 32'h24822800;
      61880: inst = 32'h10a00000;
      61881: inst = 32'hca00004;
      61882: inst = 32'h38632800;
      61883: inst = 32'h38842800;
      61884: inst = 32'h10a00000;
      61885: inst = 32'hca0f1c1;
      61886: inst = 32'h13e00001;
      61887: inst = 32'hfe0d96a;
      61888: inst = 32'h5be00000;
      61889: inst = 32'h8c50000;
      61890: inst = 32'h24612800;
      61891: inst = 32'h10a0ffff;
      61892: inst = 32'hca0fff3;
      61893: inst = 32'h24822800;
      61894: inst = 32'h10a00000;
      61895: inst = 32'hca00004;
      61896: inst = 32'h38632800;
      61897: inst = 32'h38842800;
      61898: inst = 32'h10a00000;
      61899: inst = 32'hca0f1cf;
      61900: inst = 32'h13e00001;
      61901: inst = 32'hfe0d96a;
      61902: inst = 32'h5be00000;
      61903: inst = 32'h8c50000;
      61904: inst = 32'h24612800;
      61905: inst = 32'h10a0ffff;
      61906: inst = 32'hca0fff3;
      61907: inst = 32'h24822800;
      61908: inst = 32'h10a00000;
      61909: inst = 32'hca00004;
      61910: inst = 32'h38632800;
      61911: inst = 32'h38842800;
      61912: inst = 32'h10a00000;
      61913: inst = 32'hca0f1dd;
      61914: inst = 32'h13e00001;
      61915: inst = 32'hfe0d96a;
      61916: inst = 32'h5be00000;
      61917: inst = 32'h8c50000;
      61918: inst = 32'h24612800;
      61919: inst = 32'h10a0ffff;
      61920: inst = 32'hca0fff3;
      61921: inst = 32'h24822800;
      61922: inst = 32'h10a00000;
      61923: inst = 32'hca00004;
      61924: inst = 32'h38632800;
      61925: inst = 32'h38842800;
      61926: inst = 32'h10a00000;
      61927: inst = 32'hca0f1eb;
      61928: inst = 32'h13e00001;
      61929: inst = 32'hfe0d96a;
      61930: inst = 32'h5be00000;
      61931: inst = 32'h8c50000;
      61932: inst = 32'h24612800;
      61933: inst = 32'h10a0ffff;
      61934: inst = 32'hca0fff3;
      61935: inst = 32'h24822800;
      61936: inst = 32'h10a00000;
      61937: inst = 32'hca00004;
      61938: inst = 32'h38632800;
      61939: inst = 32'h38842800;
      61940: inst = 32'h10a00000;
      61941: inst = 32'hca0f1f9;
      61942: inst = 32'h13e00001;
      61943: inst = 32'hfe0d96a;
      61944: inst = 32'h5be00000;
      61945: inst = 32'h8c50000;
      61946: inst = 32'h24612800;
      61947: inst = 32'h10a0ffff;
      61948: inst = 32'hca0fff3;
      61949: inst = 32'h24822800;
      61950: inst = 32'h10a00000;
      61951: inst = 32'hca00004;
      61952: inst = 32'h38632800;
      61953: inst = 32'h38842800;
      61954: inst = 32'h10a00000;
      61955: inst = 32'hca0f207;
      61956: inst = 32'h13e00001;
      61957: inst = 32'hfe0d96a;
      61958: inst = 32'h5be00000;
      61959: inst = 32'h8c50000;
      61960: inst = 32'h24612800;
      61961: inst = 32'h10a0ffff;
      61962: inst = 32'hca0fff3;
      61963: inst = 32'h24822800;
      61964: inst = 32'h10a00000;
      61965: inst = 32'hca00004;
      61966: inst = 32'h38632800;
      61967: inst = 32'h38842800;
      61968: inst = 32'h10a00000;
      61969: inst = 32'hca0f215;
      61970: inst = 32'h13e00001;
      61971: inst = 32'hfe0d96a;
      61972: inst = 32'h5be00000;
      61973: inst = 32'h8c50000;
      61974: inst = 32'h24612800;
      61975: inst = 32'h10a0ffff;
      61976: inst = 32'hca0fff3;
      61977: inst = 32'h24822800;
      61978: inst = 32'h10a00000;
      61979: inst = 32'hca00004;
      61980: inst = 32'h38632800;
      61981: inst = 32'h38842800;
      61982: inst = 32'h10a00000;
      61983: inst = 32'hca0f223;
      61984: inst = 32'h13e00001;
      61985: inst = 32'hfe0d96a;
      61986: inst = 32'h5be00000;
      61987: inst = 32'h8c50000;
      61988: inst = 32'h24612800;
      61989: inst = 32'h10a0ffff;
      61990: inst = 32'hca0fff3;
      61991: inst = 32'h24822800;
      61992: inst = 32'h10a00000;
      61993: inst = 32'hca00004;
      61994: inst = 32'h38632800;
      61995: inst = 32'h38842800;
      61996: inst = 32'h10a00000;
      61997: inst = 32'hca0f231;
      61998: inst = 32'h13e00001;
      61999: inst = 32'hfe0d96a;
      62000: inst = 32'h5be00000;
      62001: inst = 32'h8c50000;
      62002: inst = 32'h24612800;
      62003: inst = 32'h10a0ffff;
      62004: inst = 32'hca0fff3;
      62005: inst = 32'h24822800;
      62006: inst = 32'h10a00000;
      62007: inst = 32'hca00004;
      62008: inst = 32'h38632800;
      62009: inst = 32'h38842800;
      62010: inst = 32'h10a00000;
      62011: inst = 32'hca0f23f;
      62012: inst = 32'h13e00001;
      62013: inst = 32'hfe0d96a;
      62014: inst = 32'h5be00000;
      62015: inst = 32'h8c50000;
      62016: inst = 32'h24612800;
      62017: inst = 32'h10a0ffff;
      62018: inst = 32'hca0fff3;
      62019: inst = 32'h24822800;
      62020: inst = 32'h10a00000;
      62021: inst = 32'hca00004;
      62022: inst = 32'h38632800;
      62023: inst = 32'h38842800;
      62024: inst = 32'h10a00000;
      62025: inst = 32'hca0f24d;
      62026: inst = 32'h13e00001;
      62027: inst = 32'hfe0d96a;
      62028: inst = 32'h5be00000;
      62029: inst = 32'h8c50000;
      62030: inst = 32'h24612800;
      62031: inst = 32'h10a0ffff;
      62032: inst = 32'hca0fff3;
      62033: inst = 32'h24822800;
      62034: inst = 32'h10a00000;
      62035: inst = 32'hca00004;
      62036: inst = 32'h38632800;
      62037: inst = 32'h38842800;
      62038: inst = 32'h10a00000;
      62039: inst = 32'hca0f25b;
      62040: inst = 32'h13e00001;
      62041: inst = 32'hfe0d96a;
      62042: inst = 32'h5be00000;
      62043: inst = 32'h8c50000;
      62044: inst = 32'h24612800;
      62045: inst = 32'h10a0ffff;
      62046: inst = 32'hca0fff3;
      62047: inst = 32'h24822800;
      62048: inst = 32'h10a00000;
      62049: inst = 32'hca00004;
      62050: inst = 32'h38632800;
      62051: inst = 32'h38842800;
      62052: inst = 32'h10a00000;
      62053: inst = 32'hca0f269;
      62054: inst = 32'h13e00001;
      62055: inst = 32'hfe0d96a;
      62056: inst = 32'h5be00000;
      62057: inst = 32'h8c50000;
      62058: inst = 32'h24612800;
      62059: inst = 32'h10a0ffff;
      62060: inst = 32'hca0fff4;
      62061: inst = 32'h24822800;
      62062: inst = 32'h10a00000;
      62063: inst = 32'hca00004;
      62064: inst = 32'h38632800;
      62065: inst = 32'h38842800;
      62066: inst = 32'h10a00000;
      62067: inst = 32'hca0f277;
      62068: inst = 32'h13e00001;
      62069: inst = 32'hfe0d96a;
      62070: inst = 32'h5be00000;
      62071: inst = 32'h8c50000;
      62072: inst = 32'h24612800;
      62073: inst = 32'h10a0ffff;
      62074: inst = 32'hca0fff4;
      62075: inst = 32'h24822800;
      62076: inst = 32'h10a00000;
      62077: inst = 32'hca00004;
      62078: inst = 32'h38632800;
      62079: inst = 32'h38842800;
      62080: inst = 32'h10a00000;
      62081: inst = 32'hca0f285;
      62082: inst = 32'h13e00001;
      62083: inst = 32'hfe0d96a;
      62084: inst = 32'h5be00000;
      62085: inst = 32'h8c50000;
      62086: inst = 32'h24612800;
      62087: inst = 32'h10a0ffff;
      62088: inst = 32'hca0fff4;
      62089: inst = 32'h24822800;
      62090: inst = 32'h10a00000;
      62091: inst = 32'hca00004;
      62092: inst = 32'h38632800;
      62093: inst = 32'h38842800;
      62094: inst = 32'h10a00000;
      62095: inst = 32'hca0f293;
      62096: inst = 32'h13e00001;
      62097: inst = 32'hfe0d96a;
      62098: inst = 32'h5be00000;
      62099: inst = 32'h8c50000;
      62100: inst = 32'h24612800;
      62101: inst = 32'h10a0ffff;
      62102: inst = 32'hca0fff4;
      62103: inst = 32'h24822800;
      62104: inst = 32'h10a00000;
      62105: inst = 32'hca00004;
      62106: inst = 32'h38632800;
      62107: inst = 32'h38842800;
      62108: inst = 32'h10a00000;
      62109: inst = 32'hca0f2a1;
      62110: inst = 32'h13e00001;
      62111: inst = 32'hfe0d96a;
      62112: inst = 32'h5be00000;
      62113: inst = 32'h8c50000;
      62114: inst = 32'h24612800;
      62115: inst = 32'h10a0ffff;
      62116: inst = 32'hca0fff4;
      62117: inst = 32'h24822800;
      62118: inst = 32'h10a00000;
      62119: inst = 32'hca00004;
      62120: inst = 32'h38632800;
      62121: inst = 32'h38842800;
      62122: inst = 32'h10a00000;
      62123: inst = 32'hca0f2af;
      62124: inst = 32'h13e00001;
      62125: inst = 32'hfe0d96a;
      62126: inst = 32'h5be00000;
      62127: inst = 32'h8c50000;
      62128: inst = 32'h24612800;
      62129: inst = 32'h10a0ffff;
      62130: inst = 32'hca0fff4;
      62131: inst = 32'h24822800;
      62132: inst = 32'h10a00000;
      62133: inst = 32'hca00004;
      62134: inst = 32'h38632800;
      62135: inst = 32'h38842800;
      62136: inst = 32'h10a00000;
      62137: inst = 32'hca0f2bd;
      62138: inst = 32'h13e00001;
      62139: inst = 32'hfe0d96a;
      62140: inst = 32'h5be00000;
      62141: inst = 32'h8c50000;
      62142: inst = 32'h24612800;
      62143: inst = 32'h10a0ffff;
      62144: inst = 32'hca0fff4;
      62145: inst = 32'h24822800;
      62146: inst = 32'h10a00000;
      62147: inst = 32'hca00004;
      62148: inst = 32'h38632800;
      62149: inst = 32'h38842800;
      62150: inst = 32'h10a00000;
      62151: inst = 32'hca0f2cb;
      62152: inst = 32'h13e00001;
      62153: inst = 32'hfe0d96a;
      62154: inst = 32'h5be00000;
      62155: inst = 32'h8c50000;
      62156: inst = 32'h24612800;
      62157: inst = 32'h10a0ffff;
      62158: inst = 32'hca0fff4;
      62159: inst = 32'h24822800;
      62160: inst = 32'h10a00000;
      62161: inst = 32'hca00004;
      62162: inst = 32'h38632800;
      62163: inst = 32'h38842800;
      62164: inst = 32'h10a00000;
      62165: inst = 32'hca0f2d9;
      62166: inst = 32'h13e00001;
      62167: inst = 32'hfe0d96a;
      62168: inst = 32'h5be00000;
      62169: inst = 32'h8c50000;
      62170: inst = 32'h24612800;
      62171: inst = 32'h10a0ffff;
      62172: inst = 32'hca0fff4;
      62173: inst = 32'h24822800;
      62174: inst = 32'h10a00000;
      62175: inst = 32'hca00004;
      62176: inst = 32'h38632800;
      62177: inst = 32'h38842800;
      62178: inst = 32'h10a00000;
      62179: inst = 32'hca0f2e7;
      62180: inst = 32'h13e00001;
      62181: inst = 32'hfe0d96a;
      62182: inst = 32'h5be00000;
      62183: inst = 32'h8c50000;
      62184: inst = 32'h24612800;
      62185: inst = 32'h10a0ffff;
      62186: inst = 32'hca0fff4;
      62187: inst = 32'h24822800;
      62188: inst = 32'h10a00000;
      62189: inst = 32'hca00004;
      62190: inst = 32'h38632800;
      62191: inst = 32'h38842800;
      62192: inst = 32'h10a00000;
      62193: inst = 32'hca0f2f5;
      62194: inst = 32'h13e00001;
      62195: inst = 32'hfe0d96a;
      62196: inst = 32'h5be00000;
      62197: inst = 32'h8c50000;
      62198: inst = 32'h24612800;
      62199: inst = 32'h10a0ffff;
      62200: inst = 32'hca0fff4;
      62201: inst = 32'h24822800;
      62202: inst = 32'h10a00000;
      62203: inst = 32'hca00004;
      62204: inst = 32'h38632800;
      62205: inst = 32'h38842800;
      62206: inst = 32'h10a00000;
      62207: inst = 32'hca0f303;
      62208: inst = 32'h13e00001;
      62209: inst = 32'hfe0d96a;
      62210: inst = 32'h5be00000;
      62211: inst = 32'h8c50000;
      62212: inst = 32'h24612800;
      62213: inst = 32'h10a0ffff;
      62214: inst = 32'hca0fff4;
      62215: inst = 32'h24822800;
      62216: inst = 32'h10a00000;
      62217: inst = 32'hca00004;
      62218: inst = 32'h38632800;
      62219: inst = 32'h38842800;
      62220: inst = 32'h10a00000;
      62221: inst = 32'hca0f311;
      62222: inst = 32'h13e00001;
      62223: inst = 32'hfe0d96a;
      62224: inst = 32'h5be00000;
      62225: inst = 32'h8c50000;
      62226: inst = 32'h24612800;
      62227: inst = 32'h10a0ffff;
      62228: inst = 32'hca0fff4;
      62229: inst = 32'h24822800;
      62230: inst = 32'h10a00000;
      62231: inst = 32'hca00004;
      62232: inst = 32'h38632800;
      62233: inst = 32'h38842800;
      62234: inst = 32'h10a00000;
      62235: inst = 32'hca0f31f;
      62236: inst = 32'h13e00001;
      62237: inst = 32'hfe0d96a;
      62238: inst = 32'h5be00000;
      62239: inst = 32'h8c50000;
      62240: inst = 32'h24612800;
      62241: inst = 32'h10a0ffff;
      62242: inst = 32'hca0fff4;
      62243: inst = 32'h24822800;
      62244: inst = 32'h10a00000;
      62245: inst = 32'hca00004;
      62246: inst = 32'h38632800;
      62247: inst = 32'h38842800;
      62248: inst = 32'h10a00000;
      62249: inst = 32'hca0f32d;
      62250: inst = 32'h13e00001;
      62251: inst = 32'hfe0d96a;
      62252: inst = 32'h5be00000;
      62253: inst = 32'h8c50000;
      62254: inst = 32'h24612800;
      62255: inst = 32'h10a0ffff;
      62256: inst = 32'hca0fff4;
      62257: inst = 32'h24822800;
      62258: inst = 32'h10a00000;
      62259: inst = 32'hca00004;
      62260: inst = 32'h38632800;
      62261: inst = 32'h38842800;
      62262: inst = 32'h10a00000;
      62263: inst = 32'hca0f33b;
      62264: inst = 32'h13e00001;
      62265: inst = 32'hfe0d96a;
      62266: inst = 32'h5be00000;
      62267: inst = 32'h8c50000;
      62268: inst = 32'h24612800;
      62269: inst = 32'h10a0ffff;
      62270: inst = 32'hca0fff4;
      62271: inst = 32'h24822800;
      62272: inst = 32'h10a00000;
      62273: inst = 32'hca00004;
      62274: inst = 32'h38632800;
      62275: inst = 32'h38842800;
      62276: inst = 32'h10a00000;
      62277: inst = 32'hca0f349;
      62278: inst = 32'h13e00001;
      62279: inst = 32'hfe0d96a;
      62280: inst = 32'h5be00000;
      62281: inst = 32'h8c50000;
      62282: inst = 32'h24612800;
      62283: inst = 32'h10a0ffff;
      62284: inst = 32'hca0fff4;
      62285: inst = 32'h24822800;
      62286: inst = 32'h10a00000;
      62287: inst = 32'hca00004;
      62288: inst = 32'h38632800;
      62289: inst = 32'h38842800;
      62290: inst = 32'h10a00000;
      62291: inst = 32'hca0f357;
      62292: inst = 32'h13e00001;
      62293: inst = 32'hfe0d96a;
      62294: inst = 32'h5be00000;
      62295: inst = 32'h8c50000;
      62296: inst = 32'h24612800;
      62297: inst = 32'h10a0ffff;
      62298: inst = 32'hca0fff4;
      62299: inst = 32'h24822800;
      62300: inst = 32'h10a00000;
      62301: inst = 32'hca00004;
      62302: inst = 32'h38632800;
      62303: inst = 32'h38842800;
      62304: inst = 32'h10a00000;
      62305: inst = 32'hca0f365;
      62306: inst = 32'h13e00001;
      62307: inst = 32'hfe0d96a;
      62308: inst = 32'h5be00000;
      62309: inst = 32'h8c50000;
      62310: inst = 32'h24612800;
      62311: inst = 32'h10a0ffff;
      62312: inst = 32'hca0fff4;
      62313: inst = 32'h24822800;
      62314: inst = 32'h10a00000;
      62315: inst = 32'hca00004;
      62316: inst = 32'h38632800;
      62317: inst = 32'h38842800;
      62318: inst = 32'h10a00000;
      62319: inst = 32'hca0f373;
      62320: inst = 32'h13e00001;
      62321: inst = 32'hfe0d96a;
      62322: inst = 32'h5be00000;
      62323: inst = 32'h8c50000;
      62324: inst = 32'h24612800;
      62325: inst = 32'h10a0ffff;
      62326: inst = 32'hca0fff4;
      62327: inst = 32'h24822800;
      62328: inst = 32'h10a00000;
      62329: inst = 32'hca00004;
      62330: inst = 32'h38632800;
      62331: inst = 32'h38842800;
      62332: inst = 32'h10a00000;
      62333: inst = 32'hca0f381;
      62334: inst = 32'h13e00001;
      62335: inst = 32'hfe0d96a;
      62336: inst = 32'h5be00000;
      62337: inst = 32'h8c50000;
      62338: inst = 32'h24612800;
      62339: inst = 32'h10a0ffff;
      62340: inst = 32'hca0fff4;
      62341: inst = 32'h24822800;
      62342: inst = 32'h10a00000;
      62343: inst = 32'hca00004;
      62344: inst = 32'h38632800;
      62345: inst = 32'h38842800;
      62346: inst = 32'h10a00000;
      62347: inst = 32'hca0f38f;
      62348: inst = 32'h13e00001;
      62349: inst = 32'hfe0d96a;
      62350: inst = 32'h5be00000;
      62351: inst = 32'h8c50000;
      62352: inst = 32'h24612800;
      62353: inst = 32'h10a0ffff;
      62354: inst = 32'hca0fff4;
      62355: inst = 32'h24822800;
      62356: inst = 32'h10a00000;
      62357: inst = 32'hca00004;
      62358: inst = 32'h38632800;
      62359: inst = 32'h38842800;
      62360: inst = 32'h10a00000;
      62361: inst = 32'hca0f39d;
      62362: inst = 32'h13e00001;
      62363: inst = 32'hfe0d96a;
      62364: inst = 32'h5be00000;
      62365: inst = 32'h8c50000;
      62366: inst = 32'h24612800;
      62367: inst = 32'h10a0ffff;
      62368: inst = 32'hca0fff4;
      62369: inst = 32'h24822800;
      62370: inst = 32'h10a00000;
      62371: inst = 32'hca00004;
      62372: inst = 32'h38632800;
      62373: inst = 32'h38842800;
      62374: inst = 32'h10a00000;
      62375: inst = 32'hca0f3ab;
      62376: inst = 32'h13e00001;
      62377: inst = 32'hfe0d96a;
      62378: inst = 32'h5be00000;
      62379: inst = 32'h8c50000;
      62380: inst = 32'h24612800;
      62381: inst = 32'h10a0ffff;
      62382: inst = 32'hca0fff4;
      62383: inst = 32'h24822800;
      62384: inst = 32'h10a00000;
      62385: inst = 32'hca00004;
      62386: inst = 32'h38632800;
      62387: inst = 32'h38842800;
      62388: inst = 32'h10a00000;
      62389: inst = 32'hca0f3b9;
      62390: inst = 32'h13e00001;
      62391: inst = 32'hfe0d96a;
      62392: inst = 32'h5be00000;
      62393: inst = 32'h8c50000;
      62394: inst = 32'h24612800;
      62395: inst = 32'h10a0ffff;
      62396: inst = 32'hca0fff4;
      62397: inst = 32'h24822800;
      62398: inst = 32'h10a00000;
      62399: inst = 32'hca00004;
      62400: inst = 32'h38632800;
      62401: inst = 32'h38842800;
      62402: inst = 32'h10a00000;
      62403: inst = 32'hca0f3c7;
      62404: inst = 32'h13e00001;
      62405: inst = 32'hfe0d96a;
      62406: inst = 32'h5be00000;
      62407: inst = 32'h8c50000;
      62408: inst = 32'h24612800;
      62409: inst = 32'h10a0ffff;
      62410: inst = 32'hca0fff4;
      62411: inst = 32'h24822800;
      62412: inst = 32'h10a00000;
      62413: inst = 32'hca00004;
      62414: inst = 32'h38632800;
      62415: inst = 32'h38842800;
      62416: inst = 32'h10a00000;
      62417: inst = 32'hca0f3d5;
      62418: inst = 32'h13e00001;
      62419: inst = 32'hfe0d96a;
      62420: inst = 32'h5be00000;
      62421: inst = 32'h8c50000;
      62422: inst = 32'h24612800;
      62423: inst = 32'h10a0ffff;
      62424: inst = 32'hca0fff4;
      62425: inst = 32'h24822800;
      62426: inst = 32'h10a00000;
      62427: inst = 32'hca00004;
      62428: inst = 32'h38632800;
      62429: inst = 32'h38842800;
      62430: inst = 32'h10a00000;
      62431: inst = 32'hca0f3e3;
      62432: inst = 32'h13e00001;
      62433: inst = 32'hfe0d96a;
      62434: inst = 32'h5be00000;
      62435: inst = 32'h8c50000;
      62436: inst = 32'h24612800;
      62437: inst = 32'h10a0ffff;
      62438: inst = 32'hca0fff4;
      62439: inst = 32'h24822800;
      62440: inst = 32'h10a00000;
      62441: inst = 32'hca00004;
      62442: inst = 32'h38632800;
      62443: inst = 32'h38842800;
      62444: inst = 32'h10a00000;
      62445: inst = 32'hca0f3f1;
      62446: inst = 32'h13e00001;
      62447: inst = 32'hfe0d96a;
      62448: inst = 32'h5be00000;
      62449: inst = 32'h8c50000;
      62450: inst = 32'h24612800;
      62451: inst = 32'h10a0ffff;
      62452: inst = 32'hca0fff4;
      62453: inst = 32'h24822800;
      62454: inst = 32'h10a00000;
      62455: inst = 32'hca00004;
      62456: inst = 32'h38632800;
      62457: inst = 32'h38842800;
      62458: inst = 32'h10a00000;
      62459: inst = 32'hca0f3ff;
      62460: inst = 32'h13e00001;
      62461: inst = 32'hfe0d96a;
      62462: inst = 32'h5be00000;
      62463: inst = 32'h8c50000;
      62464: inst = 32'h24612800;
      62465: inst = 32'h10a0ffff;
      62466: inst = 32'hca0fff4;
      62467: inst = 32'h24822800;
      62468: inst = 32'h10a00000;
      62469: inst = 32'hca00004;
      62470: inst = 32'h38632800;
      62471: inst = 32'h38842800;
      62472: inst = 32'h10a00000;
      62473: inst = 32'hca0f40d;
      62474: inst = 32'h13e00001;
      62475: inst = 32'hfe0d96a;
      62476: inst = 32'h5be00000;
      62477: inst = 32'h8c50000;
      62478: inst = 32'h24612800;
      62479: inst = 32'h10a0ffff;
      62480: inst = 32'hca0fff4;
      62481: inst = 32'h24822800;
      62482: inst = 32'h10a00000;
      62483: inst = 32'hca00004;
      62484: inst = 32'h38632800;
      62485: inst = 32'h38842800;
      62486: inst = 32'h10a00000;
      62487: inst = 32'hca0f41b;
      62488: inst = 32'h13e00001;
      62489: inst = 32'hfe0d96a;
      62490: inst = 32'h5be00000;
      62491: inst = 32'h8c50000;
      62492: inst = 32'h24612800;
      62493: inst = 32'h10a0ffff;
      62494: inst = 32'hca0fff4;
      62495: inst = 32'h24822800;
      62496: inst = 32'h10a00000;
      62497: inst = 32'hca00004;
      62498: inst = 32'h38632800;
      62499: inst = 32'h38842800;
      62500: inst = 32'h10a00000;
      62501: inst = 32'hca0f429;
      62502: inst = 32'h13e00001;
      62503: inst = 32'hfe0d96a;
      62504: inst = 32'h5be00000;
      62505: inst = 32'h8c50000;
      62506: inst = 32'h24612800;
      62507: inst = 32'h10a0ffff;
      62508: inst = 32'hca0fff4;
      62509: inst = 32'h24822800;
      62510: inst = 32'h10a00000;
      62511: inst = 32'hca00004;
      62512: inst = 32'h38632800;
      62513: inst = 32'h38842800;
      62514: inst = 32'h10a00000;
      62515: inst = 32'hca0f437;
      62516: inst = 32'h13e00001;
      62517: inst = 32'hfe0d96a;
      62518: inst = 32'h5be00000;
      62519: inst = 32'h8c50000;
      62520: inst = 32'h24612800;
      62521: inst = 32'h10a0ffff;
      62522: inst = 32'hca0fff4;
      62523: inst = 32'h24822800;
      62524: inst = 32'h10a00000;
      62525: inst = 32'hca00004;
      62526: inst = 32'h38632800;
      62527: inst = 32'h38842800;
      62528: inst = 32'h10a00000;
      62529: inst = 32'hca0f445;
      62530: inst = 32'h13e00001;
      62531: inst = 32'hfe0d96a;
      62532: inst = 32'h5be00000;
      62533: inst = 32'h8c50000;
      62534: inst = 32'h24612800;
      62535: inst = 32'h10a0ffff;
      62536: inst = 32'hca0fff4;
      62537: inst = 32'h24822800;
      62538: inst = 32'h10a00000;
      62539: inst = 32'hca00004;
      62540: inst = 32'h38632800;
      62541: inst = 32'h38842800;
      62542: inst = 32'h10a00000;
      62543: inst = 32'hca0f453;
      62544: inst = 32'h13e00001;
      62545: inst = 32'hfe0d96a;
      62546: inst = 32'h5be00000;
      62547: inst = 32'h8c50000;
      62548: inst = 32'h24612800;
      62549: inst = 32'h10a0ffff;
      62550: inst = 32'hca0fff4;
      62551: inst = 32'h24822800;
      62552: inst = 32'h10a00000;
      62553: inst = 32'hca00004;
      62554: inst = 32'h38632800;
      62555: inst = 32'h38842800;
      62556: inst = 32'h10a00000;
      62557: inst = 32'hca0f461;
      62558: inst = 32'h13e00001;
      62559: inst = 32'hfe0d96a;
      62560: inst = 32'h5be00000;
      62561: inst = 32'h8c50000;
      62562: inst = 32'h24612800;
      62563: inst = 32'h10a0ffff;
      62564: inst = 32'hca0fff4;
      62565: inst = 32'h24822800;
      62566: inst = 32'h10a00000;
      62567: inst = 32'hca00004;
      62568: inst = 32'h38632800;
      62569: inst = 32'h38842800;
      62570: inst = 32'h10a00000;
      62571: inst = 32'hca0f46f;
      62572: inst = 32'h13e00001;
      62573: inst = 32'hfe0d96a;
      62574: inst = 32'h5be00000;
      62575: inst = 32'h8c50000;
      62576: inst = 32'h24612800;
      62577: inst = 32'h10a0ffff;
      62578: inst = 32'hca0fff4;
      62579: inst = 32'h24822800;
      62580: inst = 32'h10a00000;
      62581: inst = 32'hca00004;
      62582: inst = 32'h38632800;
      62583: inst = 32'h38842800;
      62584: inst = 32'h10a00000;
      62585: inst = 32'hca0f47d;
      62586: inst = 32'h13e00001;
      62587: inst = 32'hfe0d96a;
      62588: inst = 32'h5be00000;
      62589: inst = 32'h8c50000;
      62590: inst = 32'h24612800;
      62591: inst = 32'h10a0ffff;
      62592: inst = 32'hca0fff4;
      62593: inst = 32'h24822800;
      62594: inst = 32'h10a00000;
      62595: inst = 32'hca00004;
      62596: inst = 32'h38632800;
      62597: inst = 32'h38842800;
      62598: inst = 32'h10a00000;
      62599: inst = 32'hca0f48b;
      62600: inst = 32'h13e00001;
      62601: inst = 32'hfe0d96a;
      62602: inst = 32'h5be00000;
      62603: inst = 32'h8c50000;
      62604: inst = 32'h24612800;
      62605: inst = 32'h10a0ffff;
      62606: inst = 32'hca0fff4;
      62607: inst = 32'h24822800;
      62608: inst = 32'h10a00000;
      62609: inst = 32'hca00004;
      62610: inst = 32'h38632800;
      62611: inst = 32'h38842800;
      62612: inst = 32'h10a00000;
      62613: inst = 32'hca0f499;
      62614: inst = 32'h13e00001;
      62615: inst = 32'hfe0d96a;
      62616: inst = 32'h5be00000;
      62617: inst = 32'h8c50000;
      62618: inst = 32'h24612800;
      62619: inst = 32'h10a0ffff;
      62620: inst = 32'hca0fff4;
      62621: inst = 32'h24822800;
      62622: inst = 32'h10a00000;
      62623: inst = 32'hca00004;
      62624: inst = 32'h38632800;
      62625: inst = 32'h38842800;
      62626: inst = 32'h10a00000;
      62627: inst = 32'hca0f4a7;
      62628: inst = 32'h13e00001;
      62629: inst = 32'hfe0d96a;
      62630: inst = 32'h5be00000;
      62631: inst = 32'h8c50000;
      62632: inst = 32'h24612800;
      62633: inst = 32'h10a0ffff;
      62634: inst = 32'hca0fff4;
      62635: inst = 32'h24822800;
      62636: inst = 32'h10a00000;
      62637: inst = 32'hca00004;
      62638: inst = 32'h38632800;
      62639: inst = 32'h38842800;
      62640: inst = 32'h10a00000;
      62641: inst = 32'hca0f4b5;
      62642: inst = 32'h13e00001;
      62643: inst = 32'hfe0d96a;
      62644: inst = 32'h5be00000;
      62645: inst = 32'h8c50000;
      62646: inst = 32'h24612800;
      62647: inst = 32'h10a0ffff;
      62648: inst = 32'hca0fff4;
      62649: inst = 32'h24822800;
      62650: inst = 32'h10a00000;
      62651: inst = 32'hca00004;
      62652: inst = 32'h38632800;
      62653: inst = 32'h38842800;
      62654: inst = 32'h10a00000;
      62655: inst = 32'hca0f4c3;
      62656: inst = 32'h13e00001;
      62657: inst = 32'hfe0d96a;
      62658: inst = 32'h5be00000;
      62659: inst = 32'h8c50000;
      62660: inst = 32'h24612800;
      62661: inst = 32'h10a0ffff;
      62662: inst = 32'hca0fff4;
      62663: inst = 32'h24822800;
      62664: inst = 32'h10a00000;
      62665: inst = 32'hca00004;
      62666: inst = 32'h38632800;
      62667: inst = 32'h38842800;
      62668: inst = 32'h10a00000;
      62669: inst = 32'hca0f4d1;
      62670: inst = 32'h13e00001;
      62671: inst = 32'hfe0d96a;
      62672: inst = 32'h5be00000;
      62673: inst = 32'h8c50000;
      62674: inst = 32'h24612800;
      62675: inst = 32'h10a0ffff;
      62676: inst = 32'hca0fff4;
      62677: inst = 32'h24822800;
      62678: inst = 32'h10a00000;
      62679: inst = 32'hca00004;
      62680: inst = 32'h38632800;
      62681: inst = 32'h38842800;
      62682: inst = 32'h10a00000;
      62683: inst = 32'hca0f4df;
      62684: inst = 32'h13e00001;
      62685: inst = 32'hfe0d96a;
      62686: inst = 32'h5be00000;
      62687: inst = 32'h8c50000;
      62688: inst = 32'h24612800;
      62689: inst = 32'h10a0ffff;
      62690: inst = 32'hca0fff4;
      62691: inst = 32'h24822800;
      62692: inst = 32'h10a00000;
      62693: inst = 32'hca00004;
      62694: inst = 32'h38632800;
      62695: inst = 32'h38842800;
      62696: inst = 32'h10a00000;
      62697: inst = 32'hca0f4ed;
      62698: inst = 32'h13e00001;
      62699: inst = 32'hfe0d96a;
      62700: inst = 32'h5be00000;
      62701: inst = 32'h8c50000;
      62702: inst = 32'h24612800;
      62703: inst = 32'h10a0ffff;
      62704: inst = 32'hca0fff4;
      62705: inst = 32'h24822800;
      62706: inst = 32'h10a00000;
      62707: inst = 32'hca00004;
      62708: inst = 32'h38632800;
      62709: inst = 32'h38842800;
      62710: inst = 32'h10a00000;
      62711: inst = 32'hca0f4fb;
      62712: inst = 32'h13e00001;
      62713: inst = 32'hfe0d96a;
      62714: inst = 32'h5be00000;
      62715: inst = 32'h8c50000;
      62716: inst = 32'h24612800;
      62717: inst = 32'h10a0ffff;
      62718: inst = 32'hca0fff4;
      62719: inst = 32'h24822800;
      62720: inst = 32'h10a00000;
      62721: inst = 32'hca00004;
      62722: inst = 32'h38632800;
      62723: inst = 32'h38842800;
      62724: inst = 32'h10a00000;
      62725: inst = 32'hca0f509;
      62726: inst = 32'h13e00001;
      62727: inst = 32'hfe0d96a;
      62728: inst = 32'h5be00000;
      62729: inst = 32'h8c50000;
      62730: inst = 32'h24612800;
      62731: inst = 32'h10a0ffff;
      62732: inst = 32'hca0fff4;
      62733: inst = 32'h24822800;
      62734: inst = 32'h10a00000;
      62735: inst = 32'hca00004;
      62736: inst = 32'h38632800;
      62737: inst = 32'h38842800;
      62738: inst = 32'h10a00000;
      62739: inst = 32'hca0f517;
      62740: inst = 32'h13e00001;
      62741: inst = 32'hfe0d96a;
      62742: inst = 32'h5be00000;
      62743: inst = 32'h8c50000;
      62744: inst = 32'h24612800;
      62745: inst = 32'h10a0ffff;
      62746: inst = 32'hca0fff4;
      62747: inst = 32'h24822800;
      62748: inst = 32'h10a00000;
      62749: inst = 32'hca00004;
      62750: inst = 32'h38632800;
      62751: inst = 32'h38842800;
      62752: inst = 32'h10a00000;
      62753: inst = 32'hca0f525;
      62754: inst = 32'h13e00001;
      62755: inst = 32'hfe0d96a;
      62756: inst = 32'h5be00000;
      62757: inst = 32'h8c50000;
      62758: inst = 32'h24612800;
      62759: inst = 32'h10a0ffff;
      62760: inst = 32'hca0fff4;
      62761: inst = 32'h24822800;
      62762: inst = 32'h10a00000;
      62763: inst = 32'hca00004;
      62764: inst = 32'h38632800;
      62765: inst = 32'h38842800;
      62766: inst = 32'h10a00000;
      62767: inst = 32'hca0f533;
      62768: inst = 32'h13e00001;
      62769: inst = 32'hfe0d96a;
      62770: inst = 32'h5be00000;
      62771: inst = 32'h8c50000;
      62772: inst = 32'h24612800;
      62773: inst = 32'h10a0ffff;
      62774: inst = 32'hca0fff4;
      62775: inst = 32'h24822800;
      62776: inst = 32'h10a00000;
      62777: inst = 32'hca00004;
      62778: inst = 32'h38632800;
      62779: inst = 32'h38842800;
      62780: inst = 32'h10a00000;
      62781: inst = 32'hca0f541;
      62782: inst = 32'h13e00001;
      62783: inst = 32'hfe0d96a;
      62784: inst = 32'h5be00000;
      62785: inst = 32'h8c50000;
      62786: inst = 32'h24612800;
      62787: inst = 32'h10a0ffff;
      62788: inst = 32'hca0fff4;
      62789: inst = 32'h24822800;
      62790: inst = 32'h10a00000;
      62791: inst = 32'hca00004;
      62792: inst = 32'h38632800;
      62793: inst = 32'h38842800;
      62794: inst = 32'h10a00000;
      62795: inst = 32'hca0f54f;
      62796: inst = 32'h13e00001;
      62797: inst = 32'hfe0d96a;
      62798: inst = 32'h5be00000;
      62799: inst = 32'h8c50000;
      62800: inst = 32'h24612800;
      62801: inst = 32'h10a0ffff;
      62802: inst = 32'hca0fff4;
      62803: inst = 32'h24822800;
      62804: inst = 32'h10a00000;
      62805: inst = 32'hca00004;
      62806: inst = 32'h38632800;
      62807: inst = 32'h38842800;
      62808: inst = 32'h10a00000;
      62809: inst = 32'hca0f55d;
      62810: inst = 32'h13e00001;
      62811: inst = 32'hfe0d96a;
      62812: inst = 32'h5be00000;
      62813: inst = 32'h8c50000;
      62814: inst = 32'h24612800;
      62815: inst = 32'h10a0ffff;
      62816: inst = 32'hca0fff4;
      62817: inst = 32'h24822800;
      62818: inst = 32'h10a00000;
      62819: inst = 32'hca00004;
      62820: inst = 32'h38632800;
      62821: inst = 32'h38842800;
      62822: inst = 32'h10a00000;
      62823: inst = 32'hca0f56b;
      62824: inst = 32'h13e00001;
      62825: inst = 32'hfe0d96a;
      62826: inst = 32'h5be00000;
      62827: inst = 32'h8c50000;
      62828: inst = 32'h24612800;
      62829: inst = 32'h10a0ffff;
      62830: inst = 32'hca0fff4;
      62831: inst = 32'h24822800;
      62832: inst = 32'h10a00000;
      62833: inst = 32'hca00004;
      62834: inst = 32'h38632800;
      62835: inst = 32'h38842800;
      62836: inst = 32'h10a00000;
      62837: inst = 32'hca0f579;
      62838: inst = 32'h13e00001;
      62839: inst = 32'hfe0d96a;
      62840: inst = 32'h5be00000;
      62841: inst = 32'h8c50000;
      62842: inst = 32'h24612800;
      62843: inst = 32'h10a0ffff;
      62844: inst = 32'hca0fff4;
      62845: inst = 32'h24822800;
      62846: inst = 32'h10a00000;
      62847: inst = 32'hca00004;
      62848: inst = 32'h38632800;
      62849: inst = 32'h38842800;
      62850: inst = 32'h10a00000;
      62851: inst = 32'hca0f587;
      62852: inst = 32'h13e00001;
      62853: inst = 32'hfe0d96a;
      62854: inst = 32'h5be00000;
      62855: inst = 32'h8c50000;
      62856: inst = 32'h24612800;
      62857: inst = 32'h10a0ffff;
      62858: inst = 32'hca0fff4;
      62859: inst = 32'h24822800;
      62860: inst = 32'h10a00000;
      62861: inst = 32'hca00004;
      62862: inst = 32'h38632800;
      62863: inst = 32'h38842800;
      62864: inst = 32'h10a00000;
      62865: inst = 32'hca0f595;
      62866: inst = 32'h13e00001;
      62867: inst = 32'hfe0d96a;
      62868: inst = 32'h5be00000;
      62869: inst = 32'h8c50000;
      62870: inst = 32'h24612800;
      62871: inst = 32'h10a0ffff;
      62872: inst = 32'hca0fff4;
      62873: inst = 32'h24822800;
      62874: inst = 32'h10a00000;
      62875: inst = 32'hca00004;
      62876: inst = 32'h38632800;
      62877: inst = 32'h38842800;
      62878: inst = 32'h10a00000;
      62879: inst = 32'hca0f5a3;
      62880: inst = 32'h13e00001;
      62881: inst = 32'hfe0d96a;
      62882: inst = 32'h5be00000;
      62883: inst = 32'h8c50000;
      62884: inst = 32'h24612800;
      62885: inst = 32'h10a0ffff;
      62886: inst = 32'hca0fff4;
      62887: inst = 32'h24822800;
      62888: inst = 32'h10a00000;
      62889: inst = 32'hca00004;
      62890: inst = 32'h38632800;
      62891: inst = 32'h38842800;
      62892: inst = 32'h10a00000;
      62893: inst = 32'hca0f5b1;
      62894: inst = 32'h13e00001;
      62895: inst = 32'hfe0d96a;
      62896: inst = 32'h5be00000;
      62897: inst = 32'h8c50000;
      62898: inst = 32'h24612800;
      62899: inst = 32'h10a0ffff;
      62900: inst = 32'hca0fff4;
      62901: inst = 32'h24822800;
      62902: inst = 32'h10a00000;
      62903: inst = 32'hca00004;
      62904: inst = 32'h38632800;
      62905: inst = 32'h38842800;
      62906: inst = 32'h10a00000;
      62907: inst = 32'hca0f5bf;
      62908: inst = 32'h13e00001;
      62909: inst = 32'hfe0d96a;
      62910: inst = 32'h5be00000;
      62911: inst = 32'h8c50000;
      62912: inst = 32'h24612800;
      62913: inst = 32'h10a0ffff;
      62914: inst = 32'hca0fff4;
      62915: inst = 32'h24822800;
      62916: inst = 32'h10a00000;
      62917: inst = 32'hca00004;
      62918: inst = 32'h38632800;
      62919: inst = 32'h38842800;
      62920: inst = 32'h10a00000;
      62921: inst = 32'hca0f5cd;
      62922: inst = 32'h13e00001;
      62923: inst = 32'hfe0d96a;
      62924: inst = 32'h5be00000;
      62925: inst = 32'h8c50000;
      62926: inst = 32'h24612800;
      62927: inst = 32'h10a0ffff;
      62928: inst = 32'hca0fff4;
      62929: inst = 32'h24822800;
      62930: inst = 32'h10a00000;
      62931: inst = 32'hca00004;
      62932: inst = 32'h38632800;
      62933: inst = 32'h38842800;
      62934: inst = 32'h10a00000;
      62935: inst = 32'hca0f5db;
      62936: inst = 32'h13e00001;
      62937: inst = 32'hfe0d96a;
      62938: inst = 32'h5be00000;
      62939: inst = 32'h8c50000;
      62940: inst = 32'h24612800;
      62941: inst = 32'h10a0ffff;
      62942: inst = 32'hca0fff4;
      62943: inst = 32'h24822800;
      62944: inst = 32'h10a00000;
      62945: inst = 32'hca00004;
      62946: inst = 32'h38632800;
      62947: inst = 32'h38842800;
      62948: inst = 32'h10a00000;
      62949: inst = 32'hca0f5e9;
      62950: inst = 32'h13e00001;
      62951: inst = 32'hfe0d96a;
      62952: inst = 32'h5be00000;
      62953: inst = 32'h8c50000;
      62954: inst = 32'h24612800;
      62955: inst = 32'h10a0ffff;
      62956: inst = 32'hca0fff4;
      62957: inst = 32'h24822800;
      62958: inst = 32'h10a00000;
      62959: inst = 32'hca00004;
      62960: inst = 32'h38632800;
      62961: inst = 32'h38842800;
      62962: inst = 32'h10a00000;
      62963: inst = 32'hca0f5f7;
      62964: inst = 32'h13e00001;
      62965: inst = 32'hfe0d96a;
      62966: inst = 32'h5be00000;
      62967: inst = 32'h8c50000;
      62968: inst = 32'h24612800;
      62969: inst = 32'h10a0ffff;
      62970: inst = 32'hca0fff4;
      62971: inst = 32'h24822800;
      62972: inst = 32'h10a00000;
      62973: inst = 32'hca00004;
      62974: inst = 32'h38632800;
      62975: inst = 32'h38842800;
      62976: inst = 32'h10a00000;
      62977: inst = 32'hca0f605;
      62978: inst = 32'h13e00001;
      62979: inst = 32'hfe0d96a;
      62980: inst = 32'h5be00000;
      62981: inst = 32'h8c50000;
      62982: inst = 32'h24612800;
      62983: inst = 32'h10a0ffff;
      62984: inst = 32'hca0fff4;
      62985: inst = 32'h24822800;
      62986: inst = 32'h10a00000;
      62987: inst = 32'hca00004;
      62988: inst = 32'h38632800;
      62989: inst = 32'h38842800;
      62990: inst = 32'h10a00000;
      62991: inst = 32'hca0f613;
      62992: inst = 32'h13e00001;
      62993: inst = 32'hfe0d96a;
      62994: inst = 32'h5be00000;
      62995: inst = 32'h8c50000;
      62996: inst = 32'h24612800;
      62997: inst = 32'h10a0ffff;
      62998: inst = 32'hca0fff4;
      62999: inst = 32'h24822800;
      63000: inst = 32'h10a00000;
      63001: inst = 32'hca00004;
      63002: inst = 32'h38632800;
      63003: inst = 32'h38842800;
      63004: inst = 32'h10a00000;
      63005: inst = 32'hca0f621;
      63006: inst = 32'h13e00001;
      63007: inst = 32'hfe0d96a;
      63008: inst = 32'h5be00000;
      63009: inst = 32'h8c50000;
      63010: inst = 32'h24612800;
      63011: inst = 32'h10a0ffff;
      63012: inst = 32'hca0fff4;
      63013: inst = 32'h24822800;
      63014: inst = 32'h10a00000;
      63015: inst = 32'hca00004;
      63016: inst = 32'h38632800;
      63017: inst = 32'h38842800;
      63018: inst = 32'h10a00000;
      63019: inst = 32'hca0f62f;
      63020: inst = 32'h13e00001;
      63021: inst = 32'hfe0d96a;
      63022: inst = 32'h5be00000;
      63023: inst = 32'h8c50000;
      63024: inst = 32'h24612800;
      63025: inst = 32'h10a0ffff;
      63026: inst = 32'hca0fff4;
      63027: inst = 32'h24822800;
      63028: inst = 32'h10a00000;
      63029: inst = 32'hca00004;
      63030: inst = 32'h38632800;
      63031: inst = 32'h38842800;
      63032: inst = 32'h10a00000;
      63033: inst = 32'hca0f63d;
      63034: inst = 32'h13e00001;
      63035: inst = 32'hfe0d96a;
      63036: inst = 32'h5be00000;
      63037: inst = 32'h8c50000;
      63038: inst = 32'h24612800;
      63039: inst = 32'h10a0ffff;
      63040: inst = 32'hca0fff4;
      63041: inst = 32'h24822800;
      63042: inst = 32'h10a00000;
      63043: inst = 32'hca00004;
      63044: inst = 32'h38632800;
      63045: inst = 32'h38842800;
      63046: inst = 32'h10a00000;
      63047: inst = 32'hca0f64b;
      63048: inst = 32'h13e00001;
      63049: inst = 32'hfe0d96a;
      63050: inst = 32'h5be00000;
      63051: inst = 32'h8c50000;
      63052: inst = 32'h24612800;
      63053: inst = 32'h10a0ffff;
      63054: inst = 32'hca0fff4;
      63055: inst = 32'h24822800;
      63056: inst = 32'h10a00000;
      63057: inst = 32'hca00004;
      63058: inst = 32'h38632800;
      63059: inst = 32'h38842800;
      63060: inst = 32'h10a00000;
      63061: inst = 32'hca0f659;
      63062: inst = 32'h13e00001;
      63063: inst = 32'hfe0d96a;
      63064: inst = 32'h5be00000;
      63065: inst = 32'h8c50000;
      63066: inst = 32'h24612800;
      63067: inst = 32'h10a0ffff;
      63068: inst = 32'hca0fff4;
      63069: inst = 32'h24822800;
      63070: inst = 32'h10a00000;
      63071: inst = 32'hca00004;
      63072: inst = 32'h38632800;
      63073: inst = 32'h38842800;
      63074: inst = 32'h10a00000;
      63075: inst = 32'hca0f667;
      63076: inst = 32'h13e00001;
      63077: inst = 32'hfe0d96a;
      63078: inst = 32'h5be00000;
      63079: inst = 32'h8c50000;
      63080: inst = 32'h24612800;
      63081: inst = 32'h10a0ffff;
      63082: inst = 32'hca0fff4;
      63083: inst = 32'h24822800;
      63084: inst = 32'h10a00000;
      63085: inst = 32'hca00004;
      63086: inst = 32'h38632800;
      63087: inst = 32'h38842800;
      63088: inst = 32'h10a00000;
      63089: inst = 32'hca0f675;
      63090: inst = 32'h13e00001;
      63091: inst = 32'hfe0d96a;
      63092: inst = 32'h5be00000;
      63093: inst = 32'h8c50000;
      63094: inst = 32'h24612800;
      63095: inst = 32'h10a0ffff;
      63096: inst = 32'hca0fff4;
      63097: inst = 32'h24822800;
      63098: inst = 32'h10a00000;
      63099: inst = 32'hca00004;
      63100: inst = 32'h38632800;
      63101: inst = 32'h38842800;
      63102: inst = 32'h10a00000;
      63103: inst = 32'hca0f683;
      63104: inst = 32'h13e00001;
      63105: inst = 32'hfe0d96a;
      63106: inst = 32'h5be00000;
      63107: inst = 32'h8c50000;
      63108: inst = 32'h24612800;
      63109: inst = 32'h10a0ffff;
      63110: inst = 32'hca0fff4;
      63111: inst = 32'h24822800;
      63112: inst = 32'h10a00000;
      63113: inst = 32'hca00004;
      63114: inst = 32'h38632800;
      63115: inst = 32'h38842800;
      63116: inst = 32'h10a00000;
      63117: inst = 32'hca0f691;
      63118: inst = 32'h13e00001;
      63119: inst = 32'hfe0d96a;
      63120: inst = 32'h5be00000;
      63121: inst = 32'h8c50000;
      63122: inst = 32'h24612800;
      63123: inst = 32'h10a0ffff;
      63124: inst = 32'hca0fff4;
      63125: inst = 32'h24822800;
      63126: inst = 32'h10a00000;
      63127: inst = 32'hca00004;
      63128: inst = 32'h38632800;
      63129: inst = 32'h38842800;
      63130: inst = 32'h10a00000;
      63131: inst = 32'hca0f69f;
      63132: inst = 32'h13e00001;
      63133: inst = 32'hfe0d96a;
      63134: inst = 32'h5be00000;
      63135: inst = 32'h8c50000;
      63136: inst = 32'h24612800;
      63137: inst = 32'h10a0ffff;
      63138: inst = 32'hca0fff4;
      63139: inst = 32'h24822800;
      63140: inst = 32'h10a00000;
      63141: inst = 32'hca00004;
      63142: inst = 32'h38632800;
      63143: inst = 32'h38842800;
      63144: inst = 32'h10a00000;
      63145: inst = 32'hca0f6ad;
      63146: inst = 32'h13e00001;
      63147: inst = 32'hfe0d96a;
      63148: inst = 32'h5be00000;
      63149: inst = 32'h8c50000;
      63150: inst = 32'h24612800;
      63151: inst = 32'h10a0ffff;
      63152: inst = 32'hca0fff4;
      63153: inst = 32'h24822800;
      63154: inst = 32'h10a00000;
      63155: inst = 32'hca00004;
      63156: inst = 32'h38632800;
      63157: inst = 32'h38842800;
      63158: inst = 32'h10a00000;
      63159: inst = 32'hca0f6bb;
      63160: inst = 32'h13e00001;
      63161: inst = 32'hfe0d96a;
      63162: inst = 32'h5be00000;
      63163: inst = 32'h8c50000;
      63164: inst = 32'h24612800;
      63165: inst = 32'h10a0ffff;
      63166: inst = 32'hca0fff4;
      63167: inst = 32'h24822800;
      63168: inst = 32'h10a00000;
      63169: inst = 32'hca00004;
      63170: inst = 32'h38632800;
      63171: inst = 32'h38842800;
      63172: inst = 32'h10a00000;
      63173: inst = 32'hca0f6c9;
      63174: inst = 32'h13e00001;
      63175: inst = 32'hfe0d96a;
      63176: inst = 32'h5be00000;
      63177: inst = 32'h8c50000;
      63178: inst = 32'h24612800;
      63179: inst = 32'h10a0ffff;
      63180: inst = 32'hca0fff4;
      63181: inst = 32'h24822800;
      63182: inst = 32'h10a00000;
      63183: inst = 32'hca00004;
      63184: inst = 32'h38632800;
      63185: inst = 32'h38842800;
      63186: inst = 32'h10a00000;
      63187: inst = 32'hca0f6d7;
      63188: inst = 32'h13e00001;
      63189: inst = 32'hfe0d96a;
      63190: inst = 32'h5be00000;
      63191: inst = 32'h8c50000;
      63192: inst = 32'h24612800;
      63193: inst = 32'h10a0ffff;
      63194: inst = 32'hca0fff4;
      63195: inst = 32'h24822800;
      63196: inst = 32'h10a00000;
      63197: inst = 32'hca00004;
      63198: inst = 32'h38632800;
      63199: inst = 32'h38842800;
      63200: inst = 32'h10a00000;
      63201: inst = 32'hca0f6e5;
      63202: inst = 32'h13e00001;
      63203: inst = 32'hfe0d96a;
      63204: inst = 32'h5be00000;
      63205: inst = 32'h8c50000;
      63206: inst = 32'h24612800;
      63207: inst = 32'h10a0ffff;
      63208: inst = 32'hca0fff4;
      63209: inst = 32'h24822800;
      63210: inst = 32'h10a00000;
      63211: inst = 32'hca00004;
      63212: inst = 32'h38632800;
      63213: inst = 32'h38842800;
      63214: inst = 32'h10a00000;
      63215: inst = 32'hca0f6f3;
      63216: inst = 32'h13e00001;
      63217: inst = 32'hfe0d96a;
      63218: inst = 32'h5be00000;
      63219: inst = 32'h8c50000;
      63220: inst = 32'h24612800;
      63221: inst = 32'h10a0ffff;
      63222: inst = 32'hca0fff4;
      63223: inst = 32'h24822800;
      63224: inst = 32'h10a00000;
      63225: inst = 32'hca00004;
      63226: inst = 32'h38632800;
      63227: inst = 32'h38842800;
      63228: inst = 32'h10a00000;
      63229: inst = 32'hca0f701;
      63230: inst = 32'h13e00001;
      63231: inst = 32'hfe0d96a;
      63232: inst = 32'h5be00000;
      63233: inst = 32'h8c50000;
      63234: inst = 32'h24612800;
      63235: inst = 32'h10a0ffff;
      63236: inst = 32'hca0fff4;
      63237: inst = 32'h24822800;
      63238: inst = 32'h10a00000;
      63239: inst = 32'hca00004;
      63240: inst = 32'h38632800;
      63241: inst = 32'h38842800;
      63242: inst = 32'h10a00000;
      63243: inst = 32'hca0f70f;
      63244: inst = 32'h13e00001;
      63245: inst = 32'hfe0d96a;
      63246: inst = 32'h5be00000;
      63247: inst = 32'h8c50000;
      63248: inst = 32'h24612800;
      63249: inst = 32'h10a0ffff;
      63250: inst = 32'hca0fff4;
      63251: inst = 32'h24822800;
      63252: inst = 32'h10a00000;
      63253: inst = 32'hca00004;
      63254: inst = 32'h38632800;
      63255: inst = 32'h38842800;
      63256: inst = 32'h10a00000;
      63257: inst = 32'hca0f71d;
      63258: inst = 32'h13e00001;
      63259: inst = 32'hfe0d96a;
      63260: inst = 32'h5be00000;
      63261: inst = 32'h8c50000;
      63262: inst = 32'h24612800;
      63263: inst = 32'h10a0ffff;
      63264: inst = 32'hca0fff4;
      63265: inst = 32'h24822800;
      63266: inst = 32'h10a00000;
      63267: inst = 32'hca00004;
      63268: inst = 32'h38632800;
      63269: inst = 32'h38842800;
      63270: inst = 32'h10a00000;
      63271: inst = 32'hca0f72b;
      63272: inst = 32'h13e00001;
      63273: inst = 32'hfe0d96a;
      63274: inst = 32'h5be00000;
      63275: inst = 32'h8c50000;
      63276: inst = 32'h24612800;
      63277: inst = 32'h10a0ffff;
      63278: inst = 32'hca0fff4;
      63279: inst = 32'h24822800;
      63280: inst = 32'h10a00000;
      63281: inst = 32'hca00004;
      63282: inst = 32'h38632800;
      63283: inst = 32'h38842800;
      63284: inst = 32'h10a00000;
      63285: inst = 32'hca0f739;
      63286: inst = 32'h13e00001;
      63287: inst = 32'hfe0d96a;
      63288: inst = 32'h5be00000;
      63289: inst = 32'h8c50000;
      63290: inst = 32'h24612800;
      63291: inst = 32'h10a0ffff;
      63292: inst = 32'hca0fff4;
      63293: inst = 32'h24822800;
      63294: inst = 32'h10a00000;
      63295: inst = 32'hca00004;
      63296: inst = 32'h38632800;
      63297: inst = 32'h38842800;
      63298: inst = 32'h10a00000;
      63299: inst = 32'hca0f747;
      63300: inst = 32'h13e00001;
      63301: inst = 32'hfe0d96a;
      63302: inst = 32'h5be00000;
      63303: inst = 32'h8c50000;
      63304: inst = 32'h24612800;
      63305: inst = 32'h10a0ffff;
      63306: inst = 32'hca0fff4;
      63307: inst = 32'h24822800;
      63308: inst = 32'h10a00000;
      63309: inst = 32'hca00004;
      63310: inst = 32'h38632800;
      63311: inst = 32'h38842800;
      63312: inst = 32'h10a00000;
      63313: inst = 32'hca0f755;
      63314: inst = 32'h13e00001;
      63315: inst = 32'hfe0d96a;
      63316: inst = 32'h5be00000;
      63317: inst = 32'h8c50000;
      63318: inst = 32'h24612800;
      63319: inst = 32'h10a0ffff;
      63320: inst = 32'hca0fff4;
      63321: inst = 32'h24822800;
      63322: inst = 32'h10a00000;
      63323: inst = 32'hca00004;
      63324: inst = 32'h38632800;
      63325: inst = 32'h38842800;
      63326: inst = 32'h10a00000;
      63327: inst = 32'hca0f763;
      63328: inst = 32'h13e00001;
      63329: inst = 32'hfe0d96a;
      63330: inst = 32'h5be00000;
      63331: inst = 32'h8c50000;
      63332: inst = 32'h24612800;
      63333: inst = 32'h10a0ffff;
      63334: inst = 32'hca0fff4;
      63335: inst = 32'h24822800;
      63336: inst = 32'h10a00000;
      63337: inst = 32'hca00004;
      63338: inst = 32'h38632800;
      63339: inst = 32'h38842800;
      63340: inst = 32'h10a00000;
      63341: inst = 32'hca0f771;
      63342: inst = 32'h13e00001;
      63343: inst = 32'hfe0d96a;
      63344: inst = 32'h5be00000;
      63345: inst = 32'h8c50000;
      63346: inst = 32'h24612800;
      63347: inst = 32'h10a0ffff;
      63348: inst = 32'hca0fff4;
      63349: inst = 32'h24822800;
      63350: inst = 32'h10a00000;
      63351: inst = 32'hca00004;
      63352: inst = 32'h38632800;
      63353: inst = 32'h38842800;
      63354: inst = 32'h10a00000;
      63355: inst = 32'hca0f77f;
      63356: inst = 32'h13e00001;
      63357: inst = 32'hfe0d96a;
      63358: inst = 32'h5be00000;
      63359: inst = 32'h8c50000;
      63360: inst = 32'h24612800;
      63361: inst = 32'h10a0ffff;
      63362: inst = 32'hca0fff4;
      63363: inst = 32'h24822800;
      63364: inst = 32'h10a00000;
      63365: inst = 32'hca00004;
      63366: inst = 32'h38632800;
      63367: inst = 32'h38842800;
      63368: inst = 32'h10a00000;
      63369: inst = 32'hca0f78d;
      63370: inst = 32'h13e00001;
      63371: inst = 32'hfe0d96a;
      63372: inst = 32'h5be00000;
      63373: inst = 32'h8c50000;
      63374: inst = 32'h24612800;
      63375: inst = 32'h10a0ffff;
      63376: inst = 32'hca0fff4;
      63377: inst = 32'h24822800;
      63378: inst = 32'h10a00000;
      63379: inst = 32'hca00004;
      63380: inst = 32'h38632800;
      63381: inst = 32'h38842800;
      63382: inst = 32'h10a00000;
      63383: inst = 32'hca0f79b;
      63384: inst = 32'h13e00001;
      63385: inst = 32'hfe0d96a;
      63386: inst = 32'h5be00000;
      63387: inst = 32'h8c50000;
      63388: inst = 32'h24612800;
      63389: inst = 32'h10a0ffff;
      63390: inst = 32'hca0fff4;
      63391: inst = 32'h24822800;
      63392: inst = 32'h10a00000;
      63393: inst = 32'hca00004;
      63394: inst = 32'h38632800;
      63395: inst = 32'h38842800;
      63396: inst = 32'h10a00000;
      63397: inst = 32'hca0f7a9;
      63398: inst = 32'h13e00001;
      63399: inst = 32'hfe0d96a;
      63400: inst = 32'h5be00000;
      63401: inst = 32'h8c50000;
      63402: inst = 32'h24612800;
      63403: inst = 32'h10a0ffff;
      63404: inst = 32'hca0fff5;
      63405: inst = 32'h24822800;
      63406: inst = 32'h10a00000;
      63407: inst = 32'hca00004;
      63408: inst = 32'h38632800;
      63409: inst = 32'h38842800;
      63410: inst = 32'h10a00000;
      63411: inst = 32'hca0f7b7;
      63412: inst = 32'h13e00001;
      63413: inst = 32'hfe0d96a;
      63414: inst = 32'h5be00000;
      63415: inst = 32'h8c50000;
      63416: inst = 32'h24612800;
      63417: inst = 32'h10a0ffff;
      63418: inst = 32'hca0fff5;
      63419: inst = 32'h24822800;
      63420: inst = 32'h10a00000;
      63421: inst = 32'hca00004;
      63422: inst = 32'h38632800;
      63423: inst = 32'h38842800;
      63424: inst = 32'h10a00000;
      63425: inst = 32'hca0f7c5;
      63426: inst = 32'h13e00001;
      63427: inst = 32'hfe0d96a;
      63428: inst = 32'h5be00000;
      63429: inst = 32'h8c50000;
      63430: inst = 32'h24612800;
      63431: inst = 32'h10a0ffff;
      63432: inst = 32'hca0fff5;
      63433: inst = 32'h24822800;
      63434: inst = 32'h10a00000;
      63435: inst = 32'hca00004;
      63436: inst = 32'h38632800;
      63437: inst = 32'h38842800;
      63438: inst = 32'h10a00000;
      63439: inst = 32'hca0f7d3;
      63440: inst = 32'h13e00001;
      63441: inst = 32'hfe0d96a;
      63442: inst = 32'h5be00000;
      63443: inst = 32'h8c50000;
      63444: inst = 32'h24612800;
      63445: inst = 32'h10a0ffff;
      63446: inst = 32'hca0fff5;
      63447: inst = 32'h24822800;
      63448: inst = 32'h10a00000;
      63449: inst = 32'hca00004;
      63450: inst = 32'h38632800;
      63451: inst = 32'h38842800;
      63452: inst = 32'h10a00000;
      63453: inst = 32'hca0f7e1;
      63454: inst = 32'h13e00001;
      63455: inst = 32'hfe0d96a;
      63456: inst = 32'h5be00000;
      63457: inst = 32'h8c50000;
      63458: inst = 32'h24612800;
      63459: inst = 32'h10a0ffff;
      63460: inst = 32'hca0fff5;
      63461: inst = 32'h24822800;
      63462: inst = 32'h10a00000;
      63463: inst = 32'hca00004;
      63464: inst = 32'h38632800;
      63465: inst = 32'h38842800;
      63466: inst = 32'h10a00000;
      63467: inst = 32'hca0f7ef;
      63468: inst = 32'h13e00001;
      63469: inst = 32'hfe0d96a;
      63470: inst = 32'h5be00000;
      63471: inst = 32'h8c50000;
      63472: inst = 32'h24612800;
      63473: inst = 32'h10a0ffff;
      63474: inst = 32'hca0fff5;
      63475: inst = 32'h24822800;
      63476: inst = 32'h10a00000;
      63477: inst = 32'hca00004;
      63478: inst = 32'h38632800;
      63479: inst = 32'h38842800;
      63480: inst = 32'h10a00000;
      63481: inst = 32'hca0f7fd;
      63482: inst = 32'h13e00001;
      63483: inst = 32'hfe0d96a;
      63484: inst = 32'h5be00000;
      63485: inst = 32'h8c50000;
      63486: inst = 32'h24612800;
      63487: inst = 32'h10a0ffff;
      63488: inst = 32'hca0fff5;
      63489: inst = 32'h24822800;
      63490: inst = 32'h10a00000;
      63491: inst = 32'hca00004;
      63492: inst = 32'h38632800;
      63493: inst = 32'h38842800;
      63494: inst = 32'h10a00000;
      63495: inst = 32'hca0f80b;
      63496: inst = 32'h13e00001;
      63497: inst = 32'hfe0d96a;
      63498: inst = 32'h5be00000;
      63499: inst = 32'h8c50000;
      63500: inst = 32'h24612800;
      63501: inst = 32'h10a0ffff;
      63502: inst = 32'hca0fff5;
      63503: inst = 32'h24822800;
      63504: inst = 32'h10a00000;
      63505: inst = 32'hca00004;
      63506: inst = 32'h38632800;
      63507: inst = 32'h38842800;
      63508: inst = 32'h10a00000;
      63509: inst = 32'hca0f819;
      63510: inst = 32'h13e00001;
      63511: inst = 32'hfe0d96a;
      63512: inst = 32'h5be00000;
      63513: inst = 32'h8c50000;
      63514: inst = 32'h24612800;
      63515: inst = 32'h10a0ffff;
      63516: inst = 32'hca0fff5;
      63517: inst = 32'h24822800;
      63518: inst = 32'h10a00000;
      63519: inst = 32'hca00004;
      63520: inst = 32'h38632800;
      63521: inst = 32'h38842800;
      63522: inst = 32'h10a00000;
      63523: inst = 32'hca0f827;
      63524: inst = 32'h13e00001;
      63525: inst = 32'hfe0d96a;
      63526: inst = 32'h5be00000;
      63527: inst = 32'h8c50000;
      63528: inst = 32'h24612800;
      63529: inst = 32'h10a0ffff;
      63530: inst = 32'hca0fff5;
      63531: inst = 32'h24822800;
      63532: inst = 32'h10a00000;
      63533: inst = 32'hca00004;
      63534: inst = 32'h38632800;
      63535: inst = 32'h38842800;
      63536: inst = 32'h10a00000;
      63537: inst = 32'hca0f835;
      63538: inst = 32'h13e00001;
      63539: inst = 32'hfe0d96a;
      63540: inst = 32'h5be00000;
      63541: inst = 32'h8c50000;
      63542: inst = 32'h24612800;
      63543: inst = 32'h10a0ffff;
      63544: inst = 32'hca0fff5;
      63545: inst = 32'h24822800;
      63546: inst = 32'h10a00000;
      63547: inst = 32'hca00004;
      63548: inst = 32'h38632800;
      63549: inst = 32'h38842800;
      63550: inst = 32'h10a00000;
      63551: inst = 32'hca0f843;
      63552: inst = 32'h13e00001;
      63553: inst = 32'hfe0d96a;
      63554: inst = 32'h5be00000;
      63555: inst = 32'h8c50000;
      63556: inst = 32'h24612800;
      63557: inst = 32'h10a0ffff;
      63558: inst = 32'hca0fff5;
      63559: inst = 32'h24822800;
      63560: inst = 32'h10a00000;
      63561: inst = 32'hca00004;
      63562: inst = 32'h38632800;
      63563: inst = 32'h38842800;
      63564: inst = 32'h10a00000;
      63565: inst = 32'hca0f851;
      63566: inst = 32'h13e00001;
      63567: inst = 32'hfe0d96a;
      63568: inst = 32'h5be00000;
      63569: inst = 32'h8c50000;
      63570: inst = 32'h24612800;
      63571: inst = 32'h10a0ffff;
      63572: inst = 32'hca0fff5;
      63573: inst = 32'h24822800;
      63574: inst = 32'h10a00000;
      63575: inst = 32'hca00004;
      63576: inst = 32'h38632800;
      63577: inst = 32'h38842800;
      63578: inst = 32'h10a00000;
      63579: inst = 32'hca0f85f;
      63580: inst = 32'h13e00001;
      63581: inst = 32'hfe0d96a;
      63582: inst = 32'h5be00000;
      63583: inst = 32'h8c50000;
      63584: inst = 32'h24612800;
      63585: inst = 32'h10a0ffff;
      63586: inst = 32'hca0fff5;
      63587: inst = 32'h24822800;
      63588: inst = 32'h10a00000;
      63589: inst = 32'hca00004;
      63590: inst = 32'h38632800;
      63591: inst = 32'h38842800;
      63592: inst = 32'h10a00000;
      63593: inst = 32'hca0f86d;
      63594: inst = 32'h13e00001;
      63595: inst = 32'hfe0d96a;
      63596: inst = 32'h5be00000;
      63597: inst = 32'h8c50000;
      63598: inst = 32'h24612800;
      63599: inst = 32'h10a0ffff;
      63600: inst = 32'hca0fff5;
      63601: inst = 32'h24822800;
      63602: inst = 32'h10a00000;
      63603: inst = 32'hca00004;
      63604: inst = 32'h38632800;
      63605: inst = 32'h38842800;
      63606: inst = 32'h10a00000;
      63607: inst = 32'hca0f87b;
      63608: inst = 32'h13e00001;
      63609: inst = 32'hfe0d96a;
      63610: inst = 32'h5be00000;
      63611: inst = 32'h8c50000;
      63612: inst = 32'h24612800;
      63613: inst = 32'h10a0ffff;
      63614: inst = 32'hca0fff5;
      63615: inst = 32'h24822800;
      63616: inst = 32'h10a00000;
      63617: inst = 32'hca00004;
      63618: inst = 32'h38632800;
      63619: inst = 32'h38842800;
      63620: inst = 32'h10a00000;
      63621: inst = 32'hca0f889;
      63622: inst = 32'h13e00001;
      63623: inst = 32'hfe0d96a;
      63624: inst = 32'h5be00000;
      63625: inst = 32'h8c50000;
      63626: inst = 32'h24612800;
      63627: inst = 32'h10a0ffff;
      63628: inst = 32'hca0fff5;
      63629: inst = 32'h24822800;
      63630: inst = 32'h10a00000;
      63631: inst = 32'hca00004;
      63632: inst = 32'h38632800;
      63633: inst = 32'h38842800;
      63634: inst = 32'h10a00000;
      63635: inst = 32'hca0f897;
      63636: inst = 32'h13e00001;
      63637: inst = 32'hfe0d96a;
      63638: inst = 32'h5be00000;
      63639: inst = 32'h8c50000;
      63640: inst = 32'h24612800;
      63641: inst = 32'h10a0ffff;
      63642: inst = 32'hca0fff5;
      63643: inst = 32'h24822800;
      63644: inst = 32'h10a00000;
      63645: inst = 32'hca00004;
      63646: inst = 32'h38632800;
      63647: inst = 32'h38842800;
      63648: inst = 32'h10a00000;
      63649: inst = 32'hca0f8a5;
      63650: inst = 32'h13e00001;
      63651: inst = 32'hfe0d96a;
      63652: inst = 32'h5be00000;
      63653: inst = 32'h8c50000;
      63654: inst = 32'h24612800;
      63655: inst = 32'h10a0ffff;
      63656: inst = 32'hca0fff5;
      63657: inst = 32'h24822800;
      63658: inst = 32'h10a00000;
      63659: inst = 32'hca00004;
      63660: inst = 32'h38632800;
      63661: inst = 32'h38842800;
      63662: inst = 32'h10a00000;
      63663: inst = 32'hca0f8b3;
      63664: inst = 32'h13e00001;
      63665: inst = 32'hfe0d96a;
      63666: inst = 32'h5be00000;
      63667: inst = 32'h8c50000;
      63668: inst = 32'h24612800;
      63669: inst = 32'h10a0ffff;
      63670: inst = 32'hca0fff5;
      63671: inst = 32'h24822800;
      63672: inst = 32'h10a00000;
      63673: inst = 32'hca00004;
      63674: inst = 32'h38632800;
      63675: inst = 32'h38842800;
      63676: inst = 32'h10a00000;
      63677: inst = 32'hca0f8c1;
      63678: inst = 32'h13e00001;
      63679: inst = 32'hfe0d96a;
      63680: inst = 32'h5be00000;
      63681: inst = 32'h8c50000;
      63682: inst = 32'h24612800;
      63683: inst = 32'h10a0ffff;
      63684: inst = 32'hca0fff5;
      63685: inst = 32'h24822800;
      63686: inst = 32'h10a00000;
      63687: inst = 32'hca00004;
      63688: inst = 32'h38632800;
      63689: inst = 32'h38842800;
      63690: inst = 32'h10a00000;
      63691: inst = 32'hca0f8cf;
      63692: inst = 32'h13e00001;
      63693: inst = 32'hfe0d96a;
      63694: inst = 32'h5be00000;
      63695: inst = 32'h8c50000;
      63696: inst = 32'h24612800;
      63697: inst = 32'h10a0ffff;
      63698: inst = 32'hca0fff5;
      63699: inst = 32'h24822800;
      63700: inst = 32'h10a00000;
      63701: inst = 32'hca00004;
      63702: inst = 32'h38632800;
      63703: inst = 32'h38842800;
      63704: inst = 32'h10a00000;
      63705: inst = 32'hca0f8dd;
      63706: inst = 32'h13e00001;
      63707: inst = 32'hfe0d96a;
      63708: inst = 32'h5be00000;
      63709: inst = 32'h8c50000;
      63710: inst = 32'h24612800;
      63711: inst = 32'h10a0ffff;
      63712: inst = 32'hca0fff5;
      63713: inst = 32'h24822800;
      63714: inst = 32'h10a00000;
      63715: inst = 32'hca00004;
      63716: inst = 32'h38632800;
      63717: inst = 32'h38842800;
      63718: inst = 32'h10a00000;
      63719: inst = 32'hca0f8eb;
      63720: inst = 32'h13e00001;
      63721: inst = 32'hfe0d96a;
      63722: inst = 32'h5be00000;
      63723: inst = 32'h8c50000;
      63724: inst = 32'h24612800;
      63725: inst = 32'h10a0ffff;
      63726: inst = 32'hca0fff5;
      63727: inst = 32'h24822800;
      63728: inst = 32'h10a00000;
      63729: inst = 32'hca00004;
      63730: inst = 32'h38632800;
      63731: inst = 32'h38842800;
      63732: inst = 32'h10a00000;
      63733: inst = 32'hca0f8f9;
      63734: inst = 32'h13e00001;
      63735: inst = 32'hfe0d96a;
      63736: inst = 32'h5be00000;
      63737: inst = 32'h8c50000;
      63738: inst = 32'h24612800;
      63739: inst = 32'h10a0ffff;
      63740: inst = 32'hca0fff5;
      63741: inst = 32'h24822800;
      63742: inst = 32'h10a00000;
      63743: inst = 32'hca00004;
      63744: inst = 32'h38632800;
      63745: inst = 32'h38842800;
      63746: inst = 32'h10a00000;
      63747: inst = 32'hca0f907;
      63748: inst = 32'h13e00001;
      63749: inst = 32'hfe0d96a;
      63750: inst = 32'h5be00000;
      63751: inst = 32'h8c50000;
      63752: inst = 32'h24612800;
      63753: inst = 32'h10a0ffff;
      63754: inst = 32'hca0fff5;
      63755: inst = 32'h24822800;
      63756: inst = 32'h10a00000;
      63757: inst = 32'hca00004;
      63758: inst = 32'h38632800;
      63759: inst = 32'h38842800;
      63760: inst = 32'h10a00000;
      63761: inst = 32'hca0f915;
      63762: inst = 32'h13e00001;
      63763: inst = 32'hfe0d96a;
      63764: inst = 32'h5be00000;
      63765: inst = 32'h8c50000;
      63766: inst = 32'h24612800;
      63767: inst = 32'h10a0ffff;
      63768: inst = 32'hca0fff5;
      63769: inst = 32'h24822800;
      63770: inst = 32'h10a00000;
      63771: inst = 32'hca00004;
      63772: inst = 32'h38632800;
      63773: inst = 32'h38842800;
      63774: inst = 32'h10a00000;
      63775: inst = 32'hca0f923;
      63776: inst = 32'h13e00001;
      63777: inst = 32'hfe0d96a;
      63778: inst = 32'h5be00000;
      63779: inst = 32'h8c50000;
      63780: inst = 32'h24612800;
      63781: inst = 32'h10a0ffff;
      63782: inst = 32'hca0fff5;
      63783: inst = 32'h24822800;
      63784: inst = 32'h10a00000;
      63785: inst = 32'hca00004;
      63786: inst = 32'h38632800;
      63787: inst = 32'h38842800;
      63788: inst = 32'h10a00000;
      63789: inst = 32'hca0f931;
      63790: inst = 32'h13e00001;
      63791: inst = 32'hfe0d96a;
      63792: inst = 32'h5be00000;
      63793: inst = 32'h8c50000;
      63794: inst = 32'h24612800;
      63795: inst = 32'h10a0ffff;
      63796: inst = 32'hca0fff5;
      63797: inst = 32'h24822800;
      63798: inst = 32'h10a00000;
      63799: inst = 32'hca00004;
      63800: inst = 32'h38632800;
      63801: inst = 32'h38842800;
      63802: inst = 32'h10a00000;
      63803: inst = 32'hca0f93f;
      63804: inst = 32'h13e00001;
      63805: inst = 32'hfe0d96a;
      63806: inst = 32'h5be00000;
      63807: inst = 32'h8c50000;
      63808: inst = 32'h24612800;
      63809: inst = 32'h10a0ffff;
      63810: inst = 32'hca0fff5;
      63811: inst = 32'h24822800;
      63812: inst = 32'h10a00000;
      63813: inst = 32'hca00004;
      63814: inst = 32'h38632800;
      63815: inst = 32'h38842800;
      63816: inst = 32'h10a00000;
      63817: inst = 32'hca0f94d;
      63818: inst = 32'h13e00001;
      63819: inst = 32'hfe0d96a;
      63820: inst = 32'h5be00000;
      63821: inst = 32'h8c50000;
      63822: inst = 32'h24612800;
      63823: inst = 32'h10a0ffff;
      63824: inst = 32'hca0fff5;
      63825: inst = 32'h24822800;
      63826: inst = 32'h10a00000;
      63827: inst = 32'hca00004;
      63828: inst = 32'h38632800;
      63829: inst = 32'h38842800;
      63830: inst = 32'h10a00000;
      63831: inst = 32'hca0f95b;
      63832: inst = 32'h13e00001;
      63833: inst = 32'hfe0d96a;
      63834: inst = 32'h5be00000;
      63835: inst = 32'h8c50000;
      63836: inst = 32'h24612800;
      63837: inst = 32'h10a0ffff;
      63838: inst = 32'hca0fff5;
      63839: inst = 32'h24822800;
      63840: inst = 32'h10a00000;
      63841: inst = 32'hca00004;
      63842: inst = 32'h38632800;
      63843: inst = 32'h38842800;
      63844: inst = 32'h10a00000;
      63845: inst = 32'hca0f969;
      63846: inst = 32'h13e00001;
      63847: inst = 32'hfe0d96a;
      63848: inst = 32'h5be00000;
      63849: inst = 32'h8c50000;
      63850: inst = 32'h24612800;
      63851: inst = 32'h10a0ffff;
      63852: inst = 32'hca0fff5;
      63853: inst = 32'h24822800;
      63854: inst = 32'h10a00000;
      63855: inst = 32'hca00004;
      63856: inst = 32'h38632800;
      63857: inst = 32'h38842800;
      63858: inst = 32'h10a00000;
      63859: inst = 32'hca0f977;
      63860: inst = 32'h13e00001;
      63861: inst = 32'hfe0d96a;
      63862: inst = 32'h5be00000;
      63863: inst = 32'h8c50000;
      63864: inst = 32'h24612800;
      63865: inst = 32'h10a0ffff;
      63866: inst = 32'hca0fff5;
      63867: inst = 32'h24822800;
      63868: inst = 32'h10a00000;
      63869: inst = 32'hca00004;
      63870: inst = 32'h38632800;
      63871: inst = 32'h38842800;
      63872: inst = 32'h10a00000;
      63873: inst = 32'hca0f985;
      63874: inst = 32'h13e00001;
      63875: inst = 32'hfe0d96a;
      63876: inst = 32'h5be00000;
      63877: inst = 32'h8c50000;
      63878: inst = 32'h24612800;
      63879: inst = 32'h10a0ffff;
      63880: inst = 32'hca0fff5;
      63881: inst = 32'h24822800;
      63882: inst = 32'h10a00000;
      63883: inst = 32'hca00004;
      63884: inst = 32'h38632800;
      63885: inst = 32'h38842800;
      63886: inst = 32'h10a00000;
      63887: inst = 32'hca0f993;
      63888: inst = 32'h13e00001;
      63889: inst = 32'hfe0d96a;
      63890: inst = 32'h5be00000;
      63891: inst = 32'h8c50000;
      63892: inst = 32'h24612800;
      63893: inst = 32'h10a0ffff;
      63894: inst = 32'hca0fff5;
      63895: inst = 32'h24822800;
      63896: inst = 32'h10a00000;
      63897: inst = 32'hca00004;
      63898: inst = 32'h38632800;
      63899: inst = 32'h38842800;
      63900: inst = 32'h10a00000;
      63901: inst = 32'hca0f9a1;
      63902: inst = 32'h13e00001;
      63903: inst = 32'hfe0d96a;
      63904: inst = 32'h5be00000;
      63905: inst = 32'h8c50000;
      63906: inst = 32'h24612800;
      63907: inst = 32'h10a0ffff;
      63908: inst = 32'hca0fff5;
      63909: inst = 32'h24822800;
      63910: inst = 32'h10a00000;
      63911: inst = 32'hca00004;
      63912: inst = 32'h38632800;
      63913: inst = 32'h38842800;
      63914: inst = 32'h10a00000;
      63915: inst = 32'hca0f9af;
      63916: inst = 32'h13e00001;
      63917: inst = 32'hfe0d96a;
      63918: inst = 32'h5be00000;
      63919: inst = 32'h8c50000;
      63920: inst = 32'h24612800;
      63921: inst = 32'h10a0ffff;
      63922: inst = 32'hca0fff5;
      63923: inst = 32'h24822800;
      63924: inst = 32'h10a00000;
      63925: inst = 32'hca00004;
      63926: inst = 32'h38632800;
      63927: inst = 32'h38842800;
      63928: inst = 32'h10a00000;
      63929: inst = 32'hca0f9bd;
      63930: inst = 32'h13e00001;
      63931: inst = 32'hfe0d96a;
      63932: inst = 32'h5be00000;
      63933: inst = 32'h8c50000;
      63934: inst = 32'h24612800;
      63935: inst = 32'h10a0ffff;
      63936: inst = 32'hca0fff5;
      63937: inst = 32'h24822800;
      63938: inst = 32'h10a00000;
      63939: inst = 32'hca00004;
      63940: inst = 32'h38632800;
      63941: inst = 32'h38842800;
      63942: inst = 32'h10a00000;
      63943: inst = 32'hca0f9cb;
      63944: inst = 32'h13e00001;
      63945: inst = 32'hfe0d96a;
      63946: inst = 32'h5be00000;
      63947: inst = 32'h8c50000;
      63948: inst = 32'h24612800;
      63949: inst = 32'h10a0ffff;
      63950: inst = 32'hca0fff5;
      63951: inst = 32'h24822800;
      63952: inst = 32'h10a00000;
      63953: inst = 32'hca00004;
      63954: inst = 32'h38632800;
      63955: inst = 32'h38842800;
      63956: inst = 32'h10a00000;
      63957: inst = 32'hca0f9d9;
      63958: inst = 32'h13e00001;
      63959: inst = 32'hfe0d96a;
      63960: inst = 32'h5be00000;
      63961: inst = 32'h8c50000;
      63962: inst = 32'h24612800;
      63963: inst = 32'h10a0ffff;
      63964: inst = 32'hca0fff5;
      63965: inst = 32'h24822800;
      63966: inst = 32'h10a00000;
      63967: inst = 32'hca00004;
      63968: inst = 32'h38632800;
      63969: inst = 32'h38842800;
      63970: inst = 32'h10a00000;
      63971: inst = 32'hca0f9e7;
      63972: inst = 32'h13e00001;
      63973: inst = 32'hfe0d96a;
      63974: inst = 32'h5be00000;
      63975: inst = 32'h8c50000;
      63976: inst = 32'h24612800;
      63977: inst = 32'h10a0ffff;
      63978: inst = 32'hca0fff5;
      63979: inst = 32'h24822800;
      63980: inst = 32'h10a00000;
      63981: inst = 32'hca00004;
      63982: inst = 32'h38632800;
      63983: inst = 32'h38842800;
      63984: inst = 32'h10a00000;
      63985: inst = 32'hca0f9f5;
      63986: inst = 32'h13e00001;
      63987: inst = 32'hfe0d96a;
      63988: inst = 32'h5be00000;
      63989: inst = 32'h8c50000;
      63990: inst = 32'h24612800;
      63991: inst = 32'h10a0ffff;
      63992: inst = 32'hca0fff5;
      63993: inst = 32'h24822800;
      63994: inst = 32'h10a00000;
      63995: inst = 32'hca00004;
      63996: inst = 32'h38632800;
      63997: inst = 32'h38842800;
      63998: inst = 32'h10a00000;
      63999: inst = 32'hca0fa03;
      64000: inst = 32'h13e00001;
      64001: inst = 32'hfe0d96a;
      64002: inst = 32'h5be00000;
      64003: inst = 32'h8c50000;
      64004: inst = 32'h24612800;
      64005: inst = 32'h10a0ffff;
      64006: inst = 32'hca0fff5;
      64007: inst = 32'h24822800;
      64008: inst = 32'h10a00000;
      64009: inst = 32'hca00004;
      64010: inst = 32'h38632800;
      64011: inst = 32'h38842800;
      64012: inst = 32'h10a00000;
      64013: inst = 32'hca0fa11;
      64014: inst = 32'h13e00001;
      64015: inst = 32'hfe0d96a;
      64016: inst = 32'h5be00000;
      64017: inst = 32'h8c50000;
      64018: inst = 32'h24612800;
      64019: inst = 32'h10a0ffff;
      64020: inst = 32'hca0fff5;
      64021: inst = 32'h24822800;
      64022: inst = 32'h10a00000;
      64023: inst = 32'hca00004;
      64024: inst = 32'h38632800;
      64025: inst = 32'h38842800;
      64026: inst = 32'h10a00000;
      64027: inst = 32'hca0fa1f;
      64028: inst = 32'h13e00001;
      64029: inst = 32'hfe0d96a;
      64030: inst = 32'h5be00000;
      64031: inst = 32'h8c50000;
      64032: inst = 32'h24612800;
      64033: inst = 32'h10a0ffff;
      64034: inst = 32'hca0fff5;
      64035: inst = 32'h24822800;
      64036: inst = 32'h10a00000;
      64037: inst = 32'hca00004;
      64038: inst = 32'h38632800;
      64039: inst = 32'h38842800;
      64040: inst = 32'h10a00000;
      64041: inst = 32'hca0fa2d;
      64042: inst = 32'h13e00001;
      64043: inst = 32'hfe0d96a;
      64044: inst = 32'h5be00000;
      64045: inst = 32'h8c50000;
      64046: inst = 32'h24612800;
      64047: inst = 32'h10a0ffff;
      64048: inst = 32'hca0fff5;
      64049: inst = 32'h24822800;
      64050: inst = 32'h10a00000;
      64051: inst = 32'hca00004;
      64052: inst = 32'h38632800;
      64053: inst = 32'h38842800;
      64054: inst = 32'h10a00000;
      64055: inst = 32'hca0fa3b;
      64056: inst = 32'h13e00001;
      64057: inst = 32'hfe0d96a;
      64058: inst = 32'h5be00000;
      64059: inst = 32'h8c50000;
      64060: inst = 32'h24612800;
      64061: inst = 32'h10a0ffff;
      64062: inst = 32'hca0fff5;
      64063: inst = 32'h24822800;
      64064: inst = 32'h10a00000;
      64065: inst = 32'hca00004;
      64066: inst = 32'h38632800;
      64067: inst = 32'h38842800;
      64068: inst = 32'h10a00000;
      64069: inst = 32'hca0fa49;
      64070: inst = 32'h13e00001;
      64071: inst = 32'hfe0d96a;
      64072: inst = 32'h5be00000;
      64073: inst = 32'h8c50000;
      64074: inst = 32'h24612800;
      64075: inst = 32'h10a0ffff;
      64076: inst = 32'hca0fff5;
      64077: inst = 32'h24822800;
      64078: inst = 32'h10a00000;
      64079: inst = 32'hca00004;
      64080: inst = 32'h38632800;
      64081: inst = 32'h38842800;
      64082: inst = 32'h10a00000;
      64083: inst = 32'hca0fa57;
      64084: inst = 32'h13e00001;
      64085: inst = 32'hfe0d96a;
      64086: inst = 32'h5be00000;
      64087: inst = 32'h8c50000;
      64088: inst = 32'h24612800;
      64089: inst = 32'h10a0ffff;
      64090: inst = 32'hca0fff5;
      64091: inst = 32'h24822800;
      64092: inst = 32'h10a00000;
      64093: inst = 32'hca00004;
      64094: inst = 32'h38632800;
      64095: inst = 32'h38842800;
      64096: inst = 32'h10a00000;
      64097: inst = 32'hca0fa65;
      64098: inst = 32'h13e00001;
      64099: inst = 32'hfe0d96a;
      64100: inst = 32'h5be00000;
      64101: inst = 32'h8c50000;
      64102: inst = 32'h24612800;
      64103: inst = 32'h10a0ffff;
      64104: inst = 32'hca0fff5;
      64105: inst = 32'h24822800;
      64106: inst = 32'h10a00000;
      64107: inst = 32'hca00004;
      64108: inst = 32'h38632800;
      64109: inst = 32'h38842800;
      64110: inst = 32'h10a00000;
      64111: inst = 32'hca0fa73;
      64112: inst = 32'h13e00001;
      64113: inst = 32'hfe0d96a;
      64114: inst = 32'h5be00000;
      64115: inst = 32'h8c50000;
      64116: inst = 32'h24612800;
      64117: inst = 32'h10a0ffff;
      64118: inst = 32'hca0fff5;
      64119: inst = 32'h24822800;
      64120: inst = 32'h10a00000;
      64121: inst = 32'hca00004;
      64122: inst = 32'h38632800;
      64123: inst = 32'h38842800;
      64124: inst = 32'h10a00000;
      64125: inst = 32'hca0fa81;
      64126: inst = 32'h13e00001;
      64127: inst = 32'hfe0d96a;
      64128: inst = 32'h5be00000;
      64129: inst = 32'h8c50000;
      64130: inst = 32'h24612800;
      64131: inst = 32'h10a0ffff;
      64132: inst = 32'hca0fff5;
      64133: inst = 32'h24822800;
      64134: inst = 32'h10a00000;
      64135: inst = 32'hca00004;
      64136: inst = 32'h38632800;
      64137: inst = 32'h38842800;
      64138: inst = 32'h10a00000;
      64139: inst = 32'hca0fa8f;
      64140: inst = 32'h13e00001;
      64141: inst = 32'hfe0d96a;
      64142: inst = 32'h5be00000;
      64143: inst = 32'h8c50000;
      64144: inst = 32'h24612800;
      64145: inst = 32'h10a0ffff;
      64146: inst = 32'hca0fff5;
      64147: inst = 32'h24822800;
      64148: inst = 32'h10a00000;
      64149: inst = 32'hca00004;
      64150: inst = 32'h38632800;
      64151: inst = 32'h38842800;
      64152: inst = 32'h10a00000;
      64153: inst = 32'hca0fa9d;
      64154: inst = 32'h13e00001;
      64155: inst = 32'hfe0d96a;
      64156: inst = 32'h5be00000;
      64157: inst = 32'h8c50000;
      64158: inst = 32'h24612800;
      64159: inst = 32'h10a0ffff;
      64160: inst = 32'hca0fff5;
      64161: inst = 32'h24822800;
      64162: inst = 32'h10a00000;
      64163: inst = 32'hca00004;
      64164: inst = 32'h38632800;
      64165: inst = 32'h38842800;
      64166: inst = 32'h10a00000;
      64167: inst = 32'hca0faab;
      64168: inst = 32'h13e00001;
      64169: inst = 32'hfe0d96a;
      64170: inst = 32'h5be00000;
      64171: inst = 32'h8c50000;
      64172: inst = 32'h24612800;
      64173: inst = 32'h10a0ffff;
      64174: inst = 32'hca0fff5;
      64175: inst = 32'h24822800;
      64176: inst = 32'h10a00000;
      64177: inst = 32'hca00004;
      64178: inst = 32'h38632800;
      64179: inst = 32'h38842800;
      64180: inst = 32'h10a00000;
      64181: inst = 32'hca0fab9;
      64182: inst = 32'h13e00001;
      64183: inst = 32'hfe0d96a;
      64184: inst = 32'h5be00000;
      64185: inst = 32'h8c50000;
      64186: inst = 32'h24612800;
      64187: inst = 32'h10a0ffff;
      64188: inst = 32'hca0fff5;
      64189: inst = 32'h24822800;
      64190: inst = 32'h10a00000;
      64191: inst = 32'hca00004;
      64192: inst = 32'h38632800;
      64193: inst = 32'h38842800;
      64194: inst = 32'h10a00000;
      64195: inst = 32'hca0fac7;
      64196: inst = 32'h13e00001;
      64197: inst = 32'hfe0d96a;
      64198: inst = 32'h5be00000;
      64199: inst = 32'h8c50000;
      64200: inst = 32'h24612800;
      64201: inst = 32'h10a0ffff;
      64202: inst = 32'hca0fff5;
      64203: inst = 32'h24822800;
      64204: inst = 32'h10a00000;
      64205: inst = 32'hca00004;
      64206: inst = 32'h38632800;
      64207: inst = 32'h38842800;
      64208: inst = 32'h10a00000;
      64209: inst = 32'hca0fad5;
      64210: inst = 32'h13e00001;
      64211: inst = 32'hfe0d96a;
      64212: inst = 32'h5be00000;
      64213: inst = 32'h8c50000;
      64214: inst = 32'h24612800;
      64215: inst = 32'h10a0ffff;
      64216: inst = 32'hca0fff5;
      64217: inst = 32'h24822800;
      64218: inst = 32'h10a00000;
      64219: inst = 32'hca00004;
      64220: inst = 32'h38632800;
      64221: inst = 32'h38842800;
      64222: inst = 32'h10a00000;
      64223: inst = 32'hca0fae3;
      64224: inst = 32'h13e00001;
      64225: inst = 32'hfe0d96a;
      64226: inst = 32'h5be00000;
      64227: inst = 32'h8c50000;
      64228: inst = 32'h24612800;
      64229: inst = 32'h10a0ffff;
      64230: inst = 32'hca0fff5;
      64231: inst = 32'h24822800;
      64232: inst = 32'h10a00000;
      64233: inst = 32'hca00004;
      64234: inst = 32'h38632800;
      64235: inst = 32'h38842800;
      64236: inst = 32'h10a00000;
      64237: inst = 32'hca0faf1;
      64238: inst = 32'h13e00001;
      64239: inst = 32'hfe0d96a;
      64240: inst = 32'h5be00000;
      64241: inst = 32'h8c50000;
      64242: inst = 32'h24612800;
      64243: inst = 32'h10a0ffff;
      64244: inst = 32'hca0fff5;
      64245: inst = 32'h24822800;
      64246: inst = 32'h10a00000;
      64247: inst = 32'hca00004;
      64248: inst = 32'h38632800;
      64249: inst = 32'h38842800;
      64250: inst = 32'h10a00000;
      64251: inst = 32'hca0faff;
      64252: inst = 32'h13e00001;
      64253: inst = 32'hfe0d96a;
      64254: inst = 32'h5be00000;
      64255: inst = 32'h8c50000;
      64256: inst = 32'h24612800;
      64257: inst = 32'h10a0ffff;
      64258: inst = 32'hca0fff5;
      64259: inst = 32'h24822800;
      64260: inst = 32'h10a00000;
      64261: inst = 32'hca00004;
      64262: inst = 32'h38632800;
      64263: inst = 32'h38842800;
      64264: inst = 32'h10a00000;
      64265: inst = 32'hca0fb0d;
      64266: inst = 32'h13e00001;
      64267: inst = 32'hfe0d96a;
      64268: inst = 32'h5be00000;
      64269: inst = 32'h8c50000;
      64270: inst = 32'h24612800;
      64271: inst = 32'h10a0ffff;
      64272: inst = 32'hca0fff5;
      64273: inst = 32'h24822800;
      64274: inst = 32'h10a00000;
      64275: inst = 32'hca00004;
      64276: inst = 32'h38632800;
      64277: inst = 32'h38842800;
      64278: inst = 32'h10a00000;
      64279: inst = 32'hca0fb1b;
      64280: inst = 32'h13e00001;
      64281: inst = 32'hfe0d96a;
      64282: inst = 32'h5be00000;
      64283: inst = 32'h8c50000;
      64284: inst = 32'h24612800;
      64285: inst = 32'h10a0ffff;
      64286: inst = 32'hca0fff5;
      64287: inst = 32'h24822800;
      64288: inst = 32'h10a00000;
      64289: inst = 32'hca00004;
      64290: inst = 32'h38632800;
      64291: inst = 32'h38842800;
      64292: inst = 32'h10a00000;
      64293: inst = 32'hca0fb29;
      64294: inst = 32'h13e00001;
      64295: inst = 32'hfe0d96a;
      64296: inst = 32'h5be00000;
      64297: inst = 32'h8c50000;
      64298: inst = 32'h24612800;
      64299: inst = 32'h10a0ffff;
      64300: inst = 32'hca0fff5;
      64301: inst = 32'h24822800;
      64302: inst = 32'h10a00000;
      64303: inst = 32'hca00004;
      64304: inst = 32'h38632800;
      64305: inst = 32'h38842800;
      64306: inst = 32'h10a00000;
      64307: inst = 32'hca0fb37;
      64308: inst = 32'h13e00001;
      64309: inst = 32'hfe0d96a;
      64310: inst = 32'h5be00000;
      64311: inst = 32'h8c50000;
      64312: inst = 32'h24612800;
      64313: inst = 32'h10a0ffff;
      64314: inst = 32'hca0fff5;
      64315: inst = 32'h24822800;
      64316: inst = 32'h10a00000;
      64317: inst = 32'hca00004;
      64318: inst = 32'h38632800;
      64319: inst = 32'h38842800;
      64320: inst = 32'h10a00000;
      64321: inst = 32'hca0fb45;
      64322: inst = 32'h13e00001;
      64323: inst = 32'hfe0d96a;
      64324: inst = 32'h5be00000;
      64325: inst = 32'h8c50000;
      64326: inst = 32'h24612800;
      64327: inst = 32'h10a0ffff;
      64328: inst = 32'hca0fff5;
      64329: inst = 32'h24822800;
      64330: inst = 32'h10a00000;
      64331: inst = 32'hca00004;
      64332: inst = 32'h38632800;
      64333: inst = 32'h38842800;
      64334: inst = 32'h10a00000;
      64335: inst = 32'hca0fb53;
      64336: inst = 32'h13e00001;
      64337: inst = 32'hfe0d96a;
      64338: inst = 32'h5be00000;
      64339: inst = 32'h8c50000;
      64340: inst = 32'h24612800;
      64341: inst = 32'h10a0ffff;
      64342: inst = 32'hca0fff5;
      64343: inst = 32'h24822800;
      64344: inst = 32'h10a00000;
      64345: inst = 32'hca00004;
      64346: inst = 32'h38632800;
      64347: inst = 32'h38842800;
      64348: inst = 32'h10a00000;
      64349: inst = 32'hca0fb61;
      64350: inst = 32'h13e00001;
      64351: inst = 32'hfe0d96a;
      64352: inst = 32'h5be00000;
      64353: inst = 32'h8c50000;
      64354: inst = 32'h24612800;
      64355: inst = 32'h10a0ffff;
      64356: inst = 32'hca0fff5;
      64357: inst = 32'h24822800;
      64358: inst = 32'h10a00000;
      64359: inst = 32'hca00004;
      64360: inst = 32'h38632800;
      64361: inst = 32'h38842800;
      64362: inst = 32'h10a00000;
      64363: inst = 32'hca0fb6f;
      64364: inst = 32'h13e00001;
      64365: inst = 32'hfe0d96a;
      64366: inst = 32'h5be00000;
      64367: inst = 32'h8c50000;
      64368: inst = 32'h24612800;
      64369: inst = 32'h10a0ffff;
      64370: inst = 32'hca0fff5;
      64371: inst = 32'h24822800;
      64372: inst = 32'h10a00000;
      64373: inst = 32'hca00004;
      64374: inst = 32'h38632800;
      64375: inst = 32'h38842800;
      64376: inst = 32'h10a00000;
      64377: inst = 32'hca0fb7d;
      64378: inst = 32'h13e00001;
      64379: inst = 32'hfe0d96a;
      64380: inst = 32'h5be00000;
      64381: inst = 32'h8c50000;
      64382: inst = 32'h24612800;
      64383: inst = 32'h10a0ffff;
      64384: inst = 32'hca0fff5;
      64385: inst = 32'h24822800;
      64386: inst = 32'h10a00000;
      64387: inst = 32'hca00004;
      64388: inst = 32'h38632800;
      64389: inst = 32'h38842800;
      64390: inst = 32'h10a00000;
      64391: inst = 32'hca0fb8b;
      64392: inst = 32'h13e00001;
      64393: inst = 32'hfe0d96a;
      64394: inst = 32'h5be00000;
      64395: inst = 32'h8c50000;
      64396: inst = 32'h24612800;
      64397: inst = 32'h10a0ffff;
      64398: inst = 32'hca0fff5;
      64399: inst = 32'h24822800;
      64400: inst = 32'h10a00000;
      64401: inst = 32'hca00004;
      64402: inst = 32'h38632800;
      64403: inst = 32'h38842800;
      64404: inst = 32'h10a00000;
      64405: inst = 32'hca0fb99;
      64406: inst = 32'h13e00001;
      64407: inst = 32'hfe0d96a;
      64408: inst = 32'h5be00000;
      64409: inst = 32'h8c50000;
      64410: inst = 32'h24612800;
      64411: inst = 32'h10a0ffff;
      64412: inst = 32'hca0fff5;
      64413: inst = 32'h24822800;
      64414: inst = 32'h10a00000;
      64415: inst = 32'hca00004;
      64416: inst = 32'h38632800;
      64417: inst = 32'h38842800;
      64418: inst = 32'h10a00000;
      64419: inst = 32'hca0fba7;
      64420: inst = 32'h13e00001;
      64421: inst = 32'hfe0d96a;
      64422: inst = 32'h5be00000;
      64423: inst = 32'h8c50000;
      64424: inst = 32'h24612800;
      64425: inst = 32'h10a0ffff;
      64426: inst = 32'hca0fff5;
      64427: inst = 32'h24822800;
      64428: inst = 32'h10a00000;
      64429: inst = 32'hca00004;
      64430: inst = 32'h38632800;
      64431: inst = 32'h38842800;
      64432: inst = 32'h10a00000;
      64433: inst = 32'hca0fbb5;
      64434: inst = 32'h13e00001;
      64435: inst = 32'hfe0d96a;
      64436: inst = 32'h5be00000;
      64437: inst = 32'h8c50000;
      64438: inst = 32'h24612800;
      64439: inst = 32'h10a0ffff;
      64440: inst = 32'hca0fff5;
      64441: inst = 32'h24822800;
      64442: inst = 32'h10a00000;
      64443: inst = 32'hca00004;
      64444: inst = 32'h38632800;
      64445: inst = 32'h38842800;
      64446: inst = 32'h10a00000;
      64447: inst = 32'hca0fbc3;
      64448: inst = 32'h13e00001;
      64449: inst = 32'hfe0d96a;
      64450: inst = 32'h5be00000;
      64451: inst = 32'h8c50000;
      64452: inst = 32'h24612800;
      64453: inst = 32'h10a0ffff;
      64454: inst = 32'hca0fff5;
      64455: inst = 32'h24822800;
      64456: inst = 32'h10a00000;
      64457: inst = 32'hca00004;
      64458: inst = 32'h38632800;
      64459: inst = 32'h38842800;
      64460: inst = 32'h10a00000;
      64461: inst = 32'hca0fbd1;
      64462: inst = 32'h13e00001;
      64463: inst = 32'hfe0d96a;
      64464: inst = 32'h5be00000;
      64465: inst = 32'h8c50000;
      64466: inst = 32'h24612800;
      64467: inst = 32'h10a0ffff;
      64468: inst = 32'hca0fff5;
      64469: inst = 32'h24822800;
      64470: inst = 32'h10a00000;
      64471: inst = 32'hca00004;
      64472: inst = 32'h38632800;
      64473: inst = 32'h38842800;
      64474: inst = 32'h10a00000;
      64475: inst = 32'hca0fbdf;
      64476: inst = 32'h13e00001;
      64477: inst = 32'hfe0d96a;
      64478: inst = 32'h5be00000;
      64479: inst = 32'h8c50000;
      64480: inst = 32'h24612800;
      64481: inst = 32'h10a0ffff;
      64482: inst = 32'hca0fff5;
      64483: inst = 32'h24822800;
      64484: inst = 32'h10a00000;
      64485: inst = 32'hca00004;
      64486: inst = 32'h38632800;
      64487: inst = 32'h38842800;
      64488: inst = 32'h10a00000;
      64489: inst = 32'hca0fbed;
      64490: inst = 32'h13e00001;
      64491: inst = 32'hfe0d96a;
      64492: inst = 32'h5be00000;
      64493: inst = 32'h8c50000;
      64494: inst = 32'h24612800;
      64495: inst = 32'h10a0ffff;
      64496: inst = 32'hca0fff5;
      64497: inst = 32'h24822800;
      64498: inst = 32'h10a00000;
      64499: inst = 32'hca00004;
      64500: inst = 32'h38632800;
      64501: inst = 32'h38842800;
      64502: inst = 32'h10a00000;
      64503: inst = 32'hca0fbfb;
      64504: inst = 32'h13e00001;
      64505: inst = 32'hfe0d96a;
      64506: inst = 32'h5be00000;
      64507: inst = 32'h8c50000;
      64508: inst = 32'h24612800;
      64509: inst = 32'h10a0ffff;
      64510: inst = 32'hca0fff5;
      64511: inst = 32'h24822800;
      64512: inst = 32'h10a00000;
      64513: inst = 32'hca00004;
      64514: inst = 32'h38632800;
      64515: inst = 32'h38842800;
      64516: inst = 32'h10a00000;
      64517: inst = 32'hca0fc09;
      64518: inst = 32'h13e00001;
      64519: inst = 32'hfe0d96a;
      64520: inst = 32'h5be00000;
      64521: inst = 32'h8c50000;
      64522: inst = 32'h24612800;
      64523: inst = 32'h10a0ffff;
      64524: inst = 32'hca0fff5;
      64525: inst = 32'h24822800;
      64526: inst = 32'h10a00000;
      64527: inst = 32'hca00004;
      64528: inst = 32'h38632800;
      64529: inst = 32'h38842800;
      64530: inst = 32'h10a00000;
      64531: inst = 32'hca0fc17;
      64532: inst = 32'h13e00001;
      64533: inst = 32'hfe0d96a;
      64534: inst = 32'h5be00000;
      64535: inst = 32'h8c50000;
      64536: inst = 32'h24612800;
      64537: inst = 32'h10a0ffff;
      64538: inst = 32'hca0fff5;
      64539: inst = 32'h24822800;
      64540: inst = 32'h10a00000;
      64541: inst = 32'hca00004;
      64542: inst = 32'h38632800;
      64543: inst = 32'h38842800;
      64544: inst = 32'h10a00000;
      64545: inst = 32'hca0fc25;
      64546: inst = 32'h13e00001;
      64547: inst = 32'hfe0d96a;
      64548: inst = 32'h5be00000;
      64549: inst = 32'h8c50000;
      64550: inst = 32'h24612800;
      64551: inst = 32'h10a0ffff;
      64552: inst = 32'hca0fff5;
      64553: inst = 32'h24822800;
      64554: inst = 32'h10a00000;
      64555: inst = 32'hca00004;
      64556: inst = 32'h38632800;
      64557: inst = 32'h38842800;
      64558: inst = 32'h10a00000;
      64559: inst = 32'hca0fc33;
      64560: inst = 32'h13e00001;
      64561: inst = 32'hfe0d96a;
      64562: inst = 32'h5be00000;
      64563: inst = 32'h8c50000;
      64564: inst = 32'h24612800;
      64565: inst = 32'h10a0ffff;
      64566: inst = 32'hca0fff5;
      64567: inst = 32'h24822800;
      64568: inst = 32'h10a00000;
      64569: inst = 32'hca00004;
      64570: inst = 32'h38632800;
      64571: inst = 32'h38842800;
      64572: inst = 32'h10a00000;
      64573: inst = 32'hca0fc41;
      64574: inst = 32'h13e00001;
      64575: inst = 32'hfe0d96a;
      64576: inst = 32'h5be00000;
      64577: inst = 32'h8c50000;
      64578: inst = 32'h24612800;
      64579: inst = 32'h10a0ffff;
      64580: inst = 32'hca0fff5;
      64581: inst = 32'h24822800;
      64582: inst = 32'h10a00000;
      64583: inst = 32'hca00004;
      64584: inst = 32'h38632800;
      64585: inst = 32'h38842800;
      64586: inst = 32'h10a00000;
      64587: inst = 32'hca0fc4f;
      64588: inst = 32'h13e00001;
      64589: inst = 32'hfe0d96a;
      64590: inst = 32'h5be00000;
      64591: inst = 32'h8c50000;
      64592: inst = 32'h24612800;
      64593: inst = 32'h10a0ffff;
      64594: inst = 32'hca0fff5;
      64595: inst = 32'h24822800;
      64596: inst = 32'h10a00000;
      64597: inst = 32'hca00004;
      64598: inst = 32'h38632800;
      64599: inst = 32'h38842800;
      64600: inst = 32'h10a00000;
      64601: inst = 32'hca0fc5d;
      64602: inst = 32'h13e00001;
      64603: inst = 32'hfe0d96a;
      64604: inst = 32'h5be00000;
      64605: inst = 32'h8c50000;
      64606: inst = 32'h24612800;
      64607: inst = 32'h10a0ffff;
      64608: inst = 32'hca0fff5;
      64609: inst = 32'h24822800;
      64610: inst = 32'h10a00000;
      64611: inst = 32'hca00004;
      64612: inst = 32'h38632800;
      64613: inst = 32'h38842800;
      64614: inst = 32'h10a00000;
      64615: inst = 32'hca0fc6b;
      64616: inst = 32'h13e00001;
      64617: inst = 32'hfe0d96a;
      64618: inst = 32'h5be00000;
      64619: inst = 32'h8c50000;
      64620: inst = 32'h24612800;
      64621: inst = 32'h10a0ffff;
      64622: inst = 32'hca0fff5;
      64623: inst = 32'h24822800;
      64624: inst = 32'h10a00000;
      64625: inst = 32'hca00004;
      64626: inst = 32'h38632800;
      64627: inst = 32'h38842800;
      64628: inst = 32'h10a00000;
      64629: inst = 32'hca0fc79;
      64630: inst = 32'h13e00001;
      64631: inst = 32'hfe0d96a;
      64632: inst = 32'h5be00000;
      64633: inst = 32'h8c50000;
      64634: inst = 32'h24612800;
      64635: inst = 32'h10a0ffff;
      64636: inst = 32'hca0fff5;
      64637: inst = 32'h24822800;
      64638: inst = 32'h10a00000;
      64639: inst = 32'hca00004;
      64640: inst = 32'h38632800;
      64641: inst = 32'h38842800;
      64642: inst = 32'h10a00000;
      64643: inst = 32'hca0fc87;
      64644: inst = 32'h13e00001;
      64645: inst = 32'hfe0d96a;
      64646: inst = 32'h5be00000;
      64647: inst = 32'h8c50000;
      64648: inst = 32'h24612800;
      64649: inst = 32'h10a0ffff;
      64650: inst = 32'hca0fff5;
      64651: inst = 32'h24822800;
      64652: inst = 32'h10a00000;
      64653: inst = 32'hca00004;
      64654: inst = 32'h38632800;
      64655: inst = 32'h38842800;
      64656: inst = 32'h10a00000;
      64657: inst = 32'hca0fc95;
      64658: inst = 32'h13e00001;
      64659: inst = 32'hfe0d96a;
      64660: inst = 32'h5be00000;
      64661: inst = 32'h8c50000;
      64662: inst = 32'h24612800;
      64663: inst = 32'h10a0ffff;
      64664: inst = 32'hca0fff5;
      64665: inst = 32'h24822800;
      64666: inst = 32'h10a00000;
      64667: inst = 32'hca00004;
      64668: inst = 32'h38632800;
      64669: inst = 32'h38842800;
      64670: inst = 32'h10a00000;
      64671: inst = 32'hca0fca3;
      64672: inst = 32'h13e00001;
      64673: inst = 32'hfe0d96a;
      64674: inst = 32'h5be00000;
      64675: inst = 32'h8c50000;
      64676: inst = 32'h24612800;
      64677: inst = 32'h10a0ffff;
      64678: inst = 32'hca0fff5;
      64679: inst = 32'h24822800;
      64680: inst = 32'h10a00000;
      64681: inst = 32'hca00004;
      64682: inst = 32'h38632800;
      64683: inst = 32'h38842800;
      64684: inst = 32'h10a00000;
      64685: inst = 32'hca0fcb1;
      64686: inst = 32'h13e00001;
      64687: inst = 32'hfe0d96a;
      64688: inst = 32'h5be00000;
      64689: inst = 32'h8c50000;
      64690: inst = 32'h24612800;
      64691: inst = 32'h10a0ffff;
      64692: inst = 32'hca0fff5;
      64693: inst = 32'h24822800;
      64694: inst = 32'h10a00000;
      64695: inst = 32'hca00004;
      64696: inst = 32'h38632800;
      64697: inst = 32'h38842800;
      64698: inst = 32'h10a00000;
      64699: inst = 32'hca0fcbf;
      64700: inst = 32'h13e00001;
      64701: inst = 32'hfe0d96a;
      64702: inst = 32'h5be00000;
      64703: inst = 32'h8c50000;
      64704: inst = 32'h24612800;
      64705: inst = 32'h10a0ffff;
      64706: inst = 32'hca0fff5;
      64707: inst = 32'h24822800;
      64708: inst = 32'h10a00000;
      64709: inst = 32'hca00004;
      64710: inst = 32'h38632800;
      64711: inst = 32'h38842800;
      64712: inst = 32'h10a00000;
      64713: inst = 32'hca0fccd;
      64714: inst = 32'h13e00001;
      64715: inst = 32'hfe0d96a;
      64716: inst = 32'h5be00000;
      64717: inst = 32'h8c50000;
      64718: inst = 32'h24612800;
      64719: inst = 32'h10a0ffff;
      64720: inst = 32'hca0fff5;
      64721: inst = 32'h24822800;
      64722: inst = 32'h10a00000;
      64723: inst = 32'hca00004;
      64724: inst = 32'h38632800;
      64725: inst = 32'h38842800;
      64726: inst = 32'h10a00000;
      64727: inst = 32'hca0fcdb;
      64728: inst = 32'h13e00001;
      64729: inst = 32'hfe0d96a;
      64730: inst = 32'h5be00000;
      64731: inst = 32'h8c50000;
      64732: inst = 32'h24612800;
      64733: inst = 32'h10a0ffff;
      64734: inst = 32'hca0fff5;
      64735: inst = 32'h24822800;
      64736: inst = 32'h10a00000;
      64737: inst = 32'hca00004;
      64738: inst = 32'h38632800;
      64739: inst = 32'h38842800;
      64740: inst = 32'h10a00000;
      64741: inst = 32'hca0fce9;
      64742: inst = 32'h13e00001;
      64743: inst = 32'hfe0d96a;
      64744: inst = 32'h5be00000;
      64745: inst = 32'h8c50000;
      64746: inst = 32'h24612800;
      64747: inst = 32'h10a0ffff;
      64748: inst = 32'hca0fff6;
      64749: inst = 32'h24822800;
      64750: inst = 32'h10a00000;
      64751: inst = 32'hca00004;
      64752: inst = 32'h38632800;
      64753: inst = 32'h38842800;
      64754: inst = 32'h10a00000;
      64755: inst = 32'hca0fcf7;
      64756: inst = 32'h13e00001;
      64757: inst = 32'hfe0d96a;
      64758: inst = 32'h5be00000;
      64759: inst = 32'h8c50000;
      64760: inst = 32'h24612800;
      64761: inst = 32'h10a0ffff;
      64762: inst = 32'hca0fff6;
      64763: inst = 32'h24822800;
      64764: inst = 32'h10a00000;
      64765: inst = 32'hca00004;
      64766: inst = 32'h38632800;
      64767: inst = 32'h38842800;
      64768: inst = 32'h10a00000;
      64769: inst = 32'hca0fd05;
      64770: inst = 32'h13e00001;
      64771: inst = 32'hfe0d96a;
      64772: inst = 32'h5be00000;
      64773: inst = 32'h8c50000;
      64774: inst = 32'h24612800;
      64775: inst = 32'h10a0ffff;
      64776: inst = 32'hca0fff6;
      64777: inst = 32'h24822800;
      64778: inst = 32'h10a00000;
      64779: inst = 32'hca00004;
      64780: inst = 32'h38632800;
      64781: inst = 32'h38842800;
      64782: inst = 32'h10a00000;
      64783: inst = 32'hca0fd13;
      64784: inst = 32'h13e00001;
      64785: inst = 32'hfe0d96a;
      64786: inst = 32'h5be00000;
      64787: inst = 32'h8c50000;
      64788: inst = 32'h24612800;
      64789: inst = 32'h10a0ffff;
      64790: inst = 32'hca0fff6;
      64791: inst = 32'h24822800;
      64792: inst = 32'h10a00000;
      64793: inst = 32'hca00004;
      64794: inst = 32'h38632800;
      64795: inst = 32'h38842800;
      64796: inst = 32'h10a00000;
      64797: inst = 32'hca0fd21;
      64798: inst = 32'h13e00001;
      64799: inst = 32'hfe0d96a;
      64800: inst = 32'h5be00000;
      64801: inst = 32'h8c50000;
      64802: inst = 32'h24612800;
      64803: inst = 32'h10a0ffff;
      64804: inst = 32'hca0fff6;
      64805: inst = 32'h24822800;
      64806: inst = 32'h10a00000;
      64807: inst = 32'hca00004;
      64808: inst = 32'h38632800;
      64809: inst = 32'h38842800;
      64810: inst = 32'h10a00000;
      64811: inst = 32'hca0fd2f;
      64812: inst = 32'h13e00001;
      64813: inst = 32'hfe0d96a;
      64814: inst = 32'h5be00000;
      64815: inst = 32'h8c50000;
      64816: inst = 32'h24612800;
      64817: inst = 32'h10a0ffff;
      64818: inst = 32'hca0fff6;
      64819: inst = 32'h24822800;
      64820: inst = 32'h10a00000;
      64821: inst = 32'hca00004;
      64822: inst = 32'h38632800;
      64823: inst = 32'h38842800;
      64824: inst = 32'h10a00000;
      64825: inst = 32'hca0fd3d;
      64826: inst = 32'h13e00001;
      64827: inst = 32'hfe0d96a;
      64828: inst = 32'h5be00000;
      64829: inst = 32'h8c50000;
      64830: inst = 32'h24612800;
      64831: inst = 32'h10a0ffff;
      64832: inst = 32'hca0fff6;
      64833: inst = 32'h24822800;
      64834: inst = 32'h10a00000;
      64835: inst = 32'hca00004;
      64836: inst = 32'h38632800;
      64837: inst = 32'h38842800;
      64838: inst = 32'h10a00000;
      64839: inst = 32'hca0fd4b;
      64840: inst = 32'h13e00001;
      64841: inst = 32'hfe0d96a;
      64842: inst = 32'h5be00000;
      64843: inst = 32'h8c50000;
      64844: inst = 32'h24612800;
      64845: inst = 32'h10a0ffff;
      64846: inst = 32'hca0fff6;
      64847: inst = 32'h24822800;
      64848: inst = 32'h10a00000;
      64849: inst = 32'hca00004;
      64850: inst = 32'h38632800;
      64851: inst = 32'h38842800;
      64852: inst = 32'h10a00000;
      64853: inst = 32'hca0fd59;
      64854: inst = 32'h13e00001;
      64855: inst = 32'hfe0d96a;
      64856: inst = 32'h5be00000;
      64857: inst = 32'h8c50000;
      64858: inst = 32'h24612800;
      64859: inst = 32'h10a0ffff;
      64860: inst = 32'hca0fff6;
      64861: inst = 32'h24822800;
      64862: inst = 32'h10a00000;
      64863: inst = 32'hca00004;
      64864: inst = 32'h38632800;
      64865: inst = 32'h38842800;
      64866: inst = 32'h10a00000;
      64867: inst = 32'hca0fd67;
      64868: inst = 32'h13e00001;
      64869: inst = 32'hfe0d96a;
      64870: inst = 32'h5be00000;
      64871: inst = 32'h8c50000;
      64872: inst = 32'h24612800;
      64873: inst = 32'h10a0ffff;
      64874: inst = 32'hca0fff6;
      64875: inst = 32'h24822800;
      64876: inst = 32'h10a00000;
      64877: inst = 32'hca00004;
      64878: inst = 32'h38632800;
      64879: inst = 32'h38842800;
      64880: inst = 32'h10a00000;
      64881: inst = 32'hca0fd75;
      64882: inst = 32'h13e00001;
      64883: inst = 32'hfe0d96a;
      64884: inst = 32'h5be00000;
      64885: inst = 32'h8c50000;
      64886: inst = 32'h24612800;
      64887: inst = 32'h10a0ffff;
      64888: inst = 32'hca0fff6;
      64889: inst = 32'h24822800;
      64890: inst = 32'h10a00000;
      64891: inst = 32'hca00004;
      64892: inst = 32'h38632800;
      64893: inst = 32'h38842800;
      64894: inst = 32'h10a00000;
      64895: inst = 32'hca0fd83;
      64896: inst = 32'h13e00001;
      64897: inst = 32'hfe0d96a;
      64898: inst = 32'h5be00000;
      64899: inst = 32'h8c50000;
      64900: inst = 32'h24612800;
      64901: inst = 32'h10a0ffff;
      64902: inst = 32'hca0fff6;
      64903: inst = 32'h24822800;
      64904: inst = 32'h10a00000;
      64905: inst = 32'hca00004;
      64906: inst = 32'h38632800;
      64907: inst = 32'h38842800;
      64908: inst = 32'h10a00000;
      64909: inst = 32'hca0fd91;
      64910: inst = 32'h13e00001;
      64911: inst = 32'hfe0d96a;
      64912: inst = 32'h5be00000;
      64913: inst = 32'h8c50000;
      64914: inst = 32'h24612800;
      64915: inst = 32'h10a0ffff;
      64916: inst = 32'hca0fff6;
      64917: inst = 32'h24822800;
      64918: inst = 32'h10a00000;
      64919: inst = 32'hca00004;
      64920: inst = 32'h38632800;
      64921: inst = 32'h38842800;
      64922: inst = 32'h10a00000;
      64923: inst = 32'hca0fd9f;
      64924: inst = 32'h13e00001;
      64925: inst = 32'hfe0d96a;
      64926: inst = 32'h5be00000;
      64927: inst = 32'h8c50000;
      64928: inst = 32'h24612800;
      64929: inst = 32'h10a0ffff;
      64930: inst = 32'hca0fff6;
      64931: inst = 32'h24822800;
      64932: inst = 32'h10a00000;
      64933: inst = 32'hca00004;
      64934: inst = 32'h38632800;
      64935: inst = 32'h38842800;
      64936: inst = 32'h10a00000;
      64937: inst = 32'hca0fdad;
      64938: inst = 32'h13e00001;
      64939: inst = 32'hfe0d96a;
      64940: inst = 32'h5be00000;
      64941: inst = 32'h8c50000;
      64942: inst = 32'h24612800;
      64943: inst = 32'h10a0ffff;
      64944: inst = 32'hca0fff6;
      64945: inst = 32'h24822800;
      64946: inst = 32'h10a00000;
      64947: inst = 32'hca00004;
      64948: inst = 32'h38632800;
      64949: inst = 32'h38842800;
      64950: inst = 32'h10a00000;
      64951: inst = 32'hca0fdbb;
      64952: inst = 32'h13e00001;
      64953: inst = 32'hfe0d96a;
      64954: inst = 32'h5be00000;
      64955: inst = 32'h8c50000;
      64956: inst = 32'h24612800;
      64957: inst = 32'h10a0ffff;
      64958: inst = 32'hca0fff6;
      64959: inst = 32'h24822800;
      64960: inst = 32'h10a00000;
      64961: inst = 32'hca00004;
      64962: inst = 32'h38632800;
      64963: inst = 32'h38842800;
      64964: inst = 32'h10a00000;
      64965: inst = 32'hca0fdc9;
      64966: inst = 32'h13e00001;
      64967: inst = 32'hfe0d96a;
      64968: inst = 32'h5be00000;
      64969: inst = 32'h8c50000;
      64970: inst = 32'h24612800;
      64971: inst = 32'h10a0ffff;
      64972: inst = 32'hca0fff6;
      64973: inst = 32'h24822800;
      64974: inst = 32'h10a00000;
      64975: inst = 32'hca00004;
      64976: inst = 32'h38632800;
      64977: inst = 32'h38842800;
      64978: inst = 32'h10a00000;
      64979: inst = 32'hca0fdd7;
      64980: inst = 32'h13e00001;
      64981: inst = 32'hfe0d96a;
      64982: inst = 32'h5be00000;
      64983: inst = 32'h8c50000;
      64984: inst = 32'h24612800;
      64985: inst = 32'h10a0ffff;
      64986: inst = 32'hca0fff6;
      64987: inst = 32'h24822800;
      64988: inst = 32'h10a00000;
      64989: inst = 32'hca00004;
      64990: inst = 32'h38632800;
      64991: inst = 32'h38842800;
      64992: inst = 32'h10a00000;
      64993: inst = 32'hca0fde5;
      64994: inst = 32'h13e00001;
      64995: inst = 32'hfe0d96a;
      64996: inst = 32'h5be00000;
      64997: inst = 32'h8c50000;
      64998: inst = 32'h24612800;
      64999: inst = 32'h10a0ffff;
      65000: inst = 32'hca0fff6;
      65001: inst = 32'h24822800;
      65002: inst = 32'h10a00000;
      65003: inst = 32'hca00004;
      65004: inst = 32'h38632800;
      65005: inst = 32'h38842800;
      65006: inst = 32'h10a00000;
      65007: inst = 32'hca0fdf3;
      65008: inst = 32'h13e00001;
      65009: inst = 32'hfe0d96a;
      65010: inst = 32'h5be00000;
      65011: inst = 32'h8c50000;
      65012: inst = 32'h24612800;
      65013: inst = 32'h10a0ffff;
      65014: inst = 32'hca0fff6;
      65015: inst = 32'h24822800;
      65016: inst = 32'h10a00000;
      65017: inst = 32'hca00004;
      65018: inst = 32'h38632800;
      65019: inst = 32'h38842800;
      65020: inst = 32'h10a00000;
      65021: inst = 32'hca0fe01;
      65022: inst = 32'h13e00001;
      65023: inst = 32'hfe0d96a;
      65024: inst = 32'h5be00000;
      65025: inst = 32'h8c50000;
      65026: inst = 32'h24612800;
      65027: inst = 32'h10a0ffff;
      65028: inst = 32'hca0fff6;
      65029: inst = 32'h24822800;
      65030: inst = 32'h10a00000;
      65031: inst = 32'hca00004;
      65032: inst = 32'h38632800;
      65033: inst = 32'h38842800;
      65034: inst = 32'h10a00000;
      65035: inst = 32'hca0fe0f;
      65036: inst = 32'h13e00001;
      65037: inst = 32'hfe0d96a;
      65038: inst = 32'h5be00000;
      65039: inst = 32'h8c50000;
      65040: inst = 32'h24612800;
      65041: inst = 32'h10a0ffff;
      65042: inst = 32'hca0fff6;
      65043: inst = 32'h24822800;
      65044: inst = 32'h10a00000;
      65045: inst = 32'hca00004;
      65046: inst = 32'h38632800;
      65047: inst = 32'h38842800;
      65048: inst = 32'h10a00000;
      65049: inst = 32'hca0fe1d;
      65050: inst = 32'h13e00001;
      65051: inst = 32'hfe0d96a;
      65052: inst = 32'h5be00000;
      65053: inst = 32'h8c50000;
      65054: inst = 32'h24612800;
      65055: inst = 32'h10a0ffff;
      65056: inst = 32'hca0fff6;
      65057: inst = 32'h24822800;
      65058: inst = 32'h10a00000;
      65059: inst = 32'hca00004;
      65060: inst = 32'h38632800;
      65061: inst = 32'h38842800;
      65062: inst = 32'h10a00000;
      65063: inst = 32'hca0fe2b;
      65064: inst = 32'h13e00001;
      65065: inst = 32'hfe0d96a;
      65066: inst = 32'h5be00000;
      65067: inst = 32'h8c50000;
      65068: inst = 32'h24612800;
      65069: inst = 32'h10a0ffff;
      65070: inst = 32'hca0fff6;
      65071: inst = 32'h24822800;
      65072: inst = 32'h10a00000;
      65073: inst = 32'hca00004;
      65074: inst = 32'h38632800;
      65075: inst = 32'h38842800;
      65076: inst = 32'h10a00000;
      65077: inst = 32'hca0fe39;
      65078: inst = 32'h13e00001;
      65079: inst = 32'hfe0d96a;
      65080: inst = 32'h5be00000;
      65081: inst = 32'h8c50000;
      65082: inst = 32'h24612800;
      65083: inst = 32'h10a0ffff;
      65084: inst = 32'hca0fff6;
      65085: inst = 32'h24822800;
      65086: inst = 32'h10a00000;
      65087: inst = 32'hca00004;
      65088: inst = 32'h38632800;
      65089: inst = 32'h38842800;
      65090: inst = 32'h10a00000;
      65091: inst = 32'hca0fe47;
      65092: inst = 32'h13e00001;
      65093: inst = 32'hfe0d96a;
      65094: inst = 32'h5be00000;
      65095: inst = 32'h8c50000;
      65096: inst = 32'h24612800;
      65097: inst = 32'h10a0ffff;
      65098: inst = 32'hca0fff6;
      65099: inst = 32'h24822800;
      65100: inst = 32'h10a00000;
      65101: inst = 32'hca00004;
      65102: inst = 32'h38632800;
      65103: inst = 32'h38842800;
      65104: inst = 32'h10a00000;
      65105: inst = 32'hca0fe55;
      65106: inst = 32'h13e00001;
      65107: inst = 32'hfe0d96a;
      65108: inst = 32'h5be00000;
      65109: inst = 32'h8c50000;
      65110: inst = 32'h24612800;
      65111: inst = 32'h10a0ffff;
      65112: inst = 32'hca0fff6;
      65113: inst = 32'h24822800;
      65114: inst = 32'h10a00000;
      65115: inst = 32'hca00004;
      65116: inst = 32'h38632800;
      65117: inst = 32'h38842800;
      65118: inst = 32'h10a00000;
      65119: inst = 32'hca0fe63;
      65120: inst = 32'h13e00001;
      65121: inst = 32'hfe0d96a;
      65122: inst = 32'h5be00000;
      65123: inst = 32'h8c50000;
      65124: inst = 32'h24612800;
      65125: inst = 32'h10a0ffff;
      65126: inst = 32'hca0fff6;
      65127: inst = 32'h24822800;
      65128: inst = 32'h10a00000;
      65129: inst = 32'hca00004;
      65130: inst = 32'h38632800;
      65131: inst = 32'h38842800;
      65132: inst = 32'h10a00000;
      65133: inst = 32'hca0fe71;
      65134: inst = 32'h13e00001;
      65135: inst = 32'hfe0d96a;
      65136: inst = 32'h5be00000;
      65137: inst = 32'h8c50000;
      65138: inst = 32'h24612800;
      65139: inst = 32'h10a0ffff;
      65140: inst = 32'hca0fff6;
      65141: inst = 32'h24822800;
      65142: inst = 32'h10a00000;
      65143: inst = 32'hca00004;
      65144: inst = 32'h38632800;
      65145: inst = 32'h38842800;
      65146: inst = 32'h10a00000;
      65147: inst = 32'hca0fe7f;
      65148: inst = 32'h13e00001;
      65149: inst = 32'hfe0d96a;
      65150: inst = 32'h5be00000;
      65151: inst = 32'h8c50000;
      65152: inst = 32'h24612800;
      65153: inst = 32'h10a0ffff;
      65154: inst = 32'hca0fff6;
      65155: inst = 32'h24822800;
      65156: inst = 32'h10a00000;
      65157: inst = 32'hca00004;
      65158: inst = 32'h38632800;
      65159: inst = 32'h38842800;
      65160: inst = 32'h10a00000;
      65161: inst = 32'hca0fe8d;
      65162: inst = 32'h13e00001;
      65163: inst = 32'hfe0d96a;
      65164: inst = 32'h5be00000;
      65165: inst = 32'h8c50000;
      65166: inst = 32'h24612800;
      65167: inst = 32'h10a0ffff;
      65168: inst = 32'hca0fff6;
      65169: inst = 32'h24822800;
      65170: inst = 32'h10a00000;
      65171: inst = 32'hca00004;
      65172: inst = 32'h38632800;
      65173: inst = 32'h38842800;
      65174: inst = 32'h10a00000;
      65175: inst = 32'hca0fe9b;
      65176: inst = 32'h13e00001;
      65177: inst = 32'hfe0d96a;
      65178: inst = 32'h5be00000;
      65179: inst = 32'h8c50000;
      65180: inst = 32'h24612800;
      65181: inst = 32'h10a0ffff;
      65182: inst = 32'hca0fff6;
      65183: inst = 32'h24822800;
      65184: inst = 32'h10a00000;
      65185: inst = 32'hca00004;
      65186: inst = 32'h38632800;
      65187: inst = 32'h38842800;
      65188: inst = 32'h10a00000;
      65189: inst = 32'hca0fea9;
      65190: inst = 32'h13e00001;
      65191: inst = 32'hfe0d96a;
      65192: inst = 32'h5be00000;
      65193: inst = 32'h8c50000;
      65194: inst = 32'h24612800;
      65195: inst = 32'h10a0ffff;
      65196: inst = 32'hca0fff6;
      65197: inst = 32'h24822800;
      65198: inst = 32'h10a00000;
      65199: inst = 32'hca00004;
      65200: inst = 32'h38632800;
      65201: inst = 32'h38842800;
      65202: inst = 32'h10a00000;
      65203: inst = 32'hca0feb7;
      65204: inst = 32'h13e00001;
      65205: inst = 32'hfe0d96a;
      65206: inst = 32'h5be00000;
      65207: inst = 32'h8c50000;
      65208: inst = 32'h24612800;
      65209: inst = 32'h10a0ffff;
      65210: inst = 32'hca0fff6;
      65211: inst = 32'h24822800;
      65212: inst = 32'h10a00000;
      65213: inst = 32'hca00004;
      65214: inst = 32'h38632800;
      65215: inst = 32'h38842800;
      65216: inst = 32'h10a00000;
      65217: inst = 32'hca0fec5;
      65218: inst = 32'h13e00001;
      65219: inst = 32'hfe0d96a;
      65220: inst = 32'h5be00000;
      65221: inst = 32'h8c50000;
      65222: inst = 32'h24612800;
      65223: inst = 32'h10a0ffff;
      65224: inst = 32'hca0fff6;
      65225: inst = 32'h24822800;
      65226: inst = 32'h10a00000;
      65227: inst = 32'hca00004;
      65228: inst = 32'h38632800;
      65229: inst = 32'h38842800;
      65230: inst = 32'h10a00000;
      65231: inst = 32'hca0fed3;
      65232: inst = 32'h13e00001;
      65233: inst = 32'hfe0d96a;
      65234: inst = 32'h5be00000;
      65235: inst = 32'h8c50000;
      65236: inst = 32'h24612800;
      65237: inst = 32'h10a0ffff;
      65238: inst = 32'hca0fff6;
      65239: inst = 32'h24822800;
      65240: inst = 32'h10a00000;
      65241: inst = 32'hca00004;
      65242: inst = 32'h38632800;
      65243: inst = 32'h38842800;
      65244: inst = 32'h10a00000;
      65245: inst = 32'hca0fee1;
      65246: inst = 32'h13e00001;
      65247: inst = 32'hfe0d96a;
      65248: inst = 32'h5be00000;
      65249: inst = 32'h8c50000;
      65250: inst = 32'h24612800;
      65251: inst = 32'h10a0ffff;
      65252: inst = 32'hca0fff6;
      65253: inst = 32'h24822800;
      65254: inst = 32'h10a00000;
      65255: inst = 32'hca00004;
      65256: inst = 32'h38632800;
      65257: inst = 32'h38842800;
      65258: inst = 32'h10a00000;
      65259: inst = 32'hca0feef;
      65260: inst = 32'h13e00001;
      65261: inst = 32'hfe0d96a;
      65262: inst = 32'h5be00000;
      65263: inst = 32'h8c50000;
      65264: inst = 32'h24612800;
      65265: inst = 32'h10a0ffff;
      65266: inst = 32'hca0fff6;
      65267: inst = 32'h24822800;
      65268: inst = 32'h10a00000;
      65269: inst = 32'hca00004;
      65270: inst = 32'h38632800;
      65271: inst = 32'h38842800;
      65272: inst = 32'h10a00000;
      65273: inst = 32'hca0fefd;
      65274: inst = 32'h13e00001;
      65275: inst = 32'hfe0d96a;
      65276: inst = 32'h5be00000;
      65277: inst = 32'h8c50000;
      65278: inst = 32'h24612800;
      65279: inst = 32'h10a0ffff;
      65280: inst = 32'hca0fff6;
      65281: inst = 32'h24822800;
      65282: inst = 32'h10a00000;
      65283: inst = 32'hca00004;
      65284: inst = 32'h38632800;
      65285: inst = 32'h38842800;
      65286: inst = 32'h10a00000;
      65287: inst = 32'hca0ff0b;
      65288: inst = 32'h13e00001;
      65289: inst = 32'hfe0d96a;
      65290: inst = 32'h5be00000;
      65291: inst = 32'h8c50000;
      65292: inst = 32'h24612800;
      65293: inst = 32'h10a0ffff;
      65294: inst = 32'hca0fff6;
      65295: inst = 32'h24822800;
      65296: inst = 32'h10a00000;
      65297: inst = 32'hca00004;
      65298: inst = 32'h38632800;
      65299: inst = 32'h38842800;
      65300: inst = 32'h10a00000;
      65301: inst = 32'hca0ff19;
      65302: inst = 32'h13e00001;
      65303: inst = 32'hfe0d96a;
      65304: inst = 32'h5be00000;
      65305: inst = 32'h8c50000;
      65306: inst = 32'h24612800;
      65307: inst = 32'h10a0ffff;
      65308: inst = 32'hca0fff6;
      65309: inst = 32'h24822800;
      65310: inst = 32'h10a00000;
      65311: inst = 32'hca00004;
      65312: inst = 32'h38632800;
      65313: inst = 32'h38842800;
      65314: inst = 32'h10a00000;
      65315: inst = 32'hca0ff27;
      65316: inst = 32'h13e00001;
      65317: inst = 32'hfe0d96a;
      65318: inst = 32'h5be00000;
      65319: inst = 32'h8c50000;
      65320: inst = 32'h24612800;
      65321: inst = 32'h10a0ffff;
      65322: inst = 32'hca0fff6;
      65323: inst = 32'h24822800;
      65324: inst = 32'h10a00000;
      65325: inst = 32'hca00004;
      65326: inst = 32'h38632800;
      65327: inst = 32'h38842800;
      65328: inst = 32'h10a00000;
      65329: inst = 32'hca0ff35;
      65330: inst = 32'h13e00001;
      65331: inst = 32'hfe0d96a;
      65332: inst = 32'h5be00000;
      65333: inst = 32'h8c50000;
      65334: inst = 32'h24612800;
      65335: inst = 32'h10a0ffff;
      65336: inst = 32'hca0fff6;
      65337: inst = 32'h24822800;
      65338: inst = 32'h10a00000;
      65339: inst = 32'hca00004;
      65340: inst = 32'h38632800;
      65341: inst = 32'h38842800;
      65342: inst = 32'h10a00000;
      65343: inst = 32'hca0ff43;
      65344: inst = 32'h13e00001;
      65345: inst = 32'hfe0d96a;
      65346: inst = 32'h5be00000;
      65347: inst = 32'h8c50000;
      65348: inst = 32'h24612800;
      65349: inst = 32'h10a0ffff;
      65350: inst = 32'hca0fff6;
      65351: inst = 32'h24822800;
      65352: inst = 32'h10a00000;
      65353: inst = 32'hca00004;
      65354: inst = 32'h38632800;
      65355: inst = 32'h38842800;
      65356: inst = 32'h10a00000;
      65357: inst = 32'hca0ff51;
      65358: inst = 32'h13e00001;
      65359: inst = 32'hfe0d96a;
      65360: inst = 32'h5be00000;
      65361: inst = 32'h8c50000;
      65362: inst = 32'h24612800;
      65363: inst = 32'h10a0ffff;
      65364: inst = 32'hca0fff6;
      65365: inst = 32'h24822800;
      65366: inst = 32'h10a00000;
      65367: inst = 32'hca00004;
      65368: inst = 32'h38632800;
      65369: inst = 32'h38842800;
      65370: inst = 32'h10a00000;
      65371: inst = 32'hca0ff5f;
      65372: inst = 32'h13e00001;
      65373: inst = 32'hfe0d96a;
      65374: inst = 32'h5be00000;
      65375: inst = 32'h8c50000;
      65376: inst = 32'h24612800;
      65377: inst = 32'h10a0ffff;
      65378: inst = 32'hca0fff6;
      65379: inst = 32'h24822800;
      65380: inst = 32'h10a00000;
      65381: inst = 32'hca00004;
      65382: inst = 32'h38632800;
      65383: inst = 32'h38842800;
      65384: inst = 32'h10a00000;
      65385: inst = 32'hca0ff6d;
      65386: inst = 32'h13e00001;
      65387: inst = 32'hfe0d96a;
      65388: inst = 32'h5be00000;
      65389: inst = 32'h8c50000;
      65390: inst = 32'h24612800;
      65391: inst = 32'h10a0ffff;
      65392: inst = 32'hca0fff6;
      65393: inst = 32'h24822800;
      65394: inst = 32'h10a00000;
      65395: inst = 32'hca00004;
      65396: inst = 32'h38632800;
      65397: inst = 32'h38842800;
      65398: inst = 32'h10a00000;
      65399: inst = 32'hca0ff7b;
      65400: inst = 32'h13e00001;
      65401: inst = 32'hfe0d96a;
      65402: inst = 32'h5be00000;
      65403: inst = 32'h8c50000;
      65404: inst = 32'h24612800;
      65405: inst = 32'h10a0ffff;
      65406: inst = 32'hca0fff6;
      65407: inst = 32'h24822800;
      65408: inst = 32'h10a00000;
      65409: inst = 32'hca00004;
      65410: inst = 32'h38632800;
      65411: inst = 32'h38842800;
      65412: inst = 32'h10a00000;
      65413: inst = 32'hca0ff89;
      65414: inst = 32'h13e00001;
      65415: inst = 32'hfe0d96a;
      65416: inst = 32'h5be00000;
      65417: inst = 32'h8c50000;
      65418: inst = 32'h24612800;
      65419: inst = 32'h10a0ffff;
      65420: inst = 32'hca0fff6;
      65421: inst = 32'h24822800;
      65422: inst = 32'h10a00000;
      65423: inst = 32'hca00004;
      65424: inst = 32'h38632800;
      65425: inst = 32'h38842800;
      65426: inst = 32'h10a00000;
      65427: inst = 32'hca0ff97;
      65428: inst = 32'h13e00001;
      65429: inst = 32'hfe0d96a;
      65430: inst = 32'h5be00000;
      65431: inst = 32'h8c50000;
      65432: inst = 32'h24612800;
      65433: inst = 32'h10a0ffff;
      65434: inst = 32'hca0fff6;
      65435: inst = 32'h24822800;
      65436: inst = 32'h10a00000;
      65437: inst = 32'hca00004;
      65438: inst = 32'h38632800;
      65439: inst = 32'h38842800;
      65440: inst = 32'h10a00000;
      65441: inst = 32'hca0ffa5;
      65442: inst = 32'h13e00001;
      65443: inst = 32'hfe0d96a;
      65444: inst = 32'h5be00000;
      65445: inst = 32'h8c50000;
      65446: inst = 32'h24612800;
      65447: inst = 32'h10a0ffff;
      65448: inst = 32'hca0fff6;
      65449: inst = 32'h24822800;
      65450: inst = 32'h10a00000;
      65451: inst = 32'hca00004;
      65452: inst = 32'h38632800;
      65453: inst = 32'h38842800;
      65454: inst = 32'h10a00000;
      65455: inst = 32'hca0ffb3;
      65456: inst = 32'h13e00001;
      65457: inst = 32'hfe0d96a;
      65458: inst = 32'h5be00000;
      65459: inst = 32'h8c50000;
      65460: inst = 32'h24612800;
      65461: inst = 32'h10a0ffff;
      65462: inst = 32'hca0fff6;
      65463: inst = 32'h24822800;
      65464: inst = 32'h10a00000;
      65465: inst = 32'hca00004;
      65466: inst = 32'h38632800;
      65467: inst = 32'h38842800;
      65468: inst = 32'h10a00000;
      65469: inst = 32'hca0ffc1;
      65470: inst = 32'h13e00001;
      65471: inst = 32'hfe0d96a;
      65472: inst = 32'h5be00000;
      65473: inst = 32'h8c50000;
      65474: inst = 32'h24612800;
      65475: inst = 32'h10a0ffff;
      65476: inst = 32'hca0fff6;
      65477: inst = 32'h24822800;
      65478: inst = 32'h10a00000;
      65479: inst = 32'hca00004;
      65480: inst = 32'h38632800;
      65481: inst = 32'h38842800;
      65482: inst = 32'h10a00000;
      65483: inst = 32'hca0ffcf;
      65484: inst = 32'h13e00001;
      65485: inst = 32'hfe0d96a;
      65486: inst = 32'h5be00000;
      65487: inst = 32'h8c50000;
      65488: inst = 32'h24612800;
      65489: inst = 32'h10a0ffff;
      65490: inst = 32'hca0fff6;
      65491: inst = 32'h24822800;
      65492: inst = 32'h10a00000;
      65493: inst = 32'hca00004;
      65494: inst = 32'h38632800;
      65495: inst = 32'h38842800;
      65496: inst = 32'h10a00000;
      65497: inst = 32'hca0ffdd;
      65498: inst = 32'h13e00001;
      65499: inst = 32'hfe0d96a;
      65500: inst = 32'h5be00000;
      65501: inst = 32'h8c50000;
      65502: inst = 32'h24612800;
      65503: inst = 32'h10a0ffff;
      65504: inst = 32'hca0fff6;
      65505: inst = 32'h24822800;
      65506: inst = 32'h10a00000;
      65507: inst = 32'hca00004;
      65508: inst = 32'h38632800;
      65509: inst = 32'h38842800;
      65510: inst = 32'h10a00000;
      65511: inst = 32'hca0ffeb;
      65512: inst = 32'h13e00001;
      65513: inst = 32'hfe0d96a;
      65514: inst = 32'h5be00000;
      65515: inst = 32'h8c50000;
      65516: inst = 32'h24612800;
      65517: inst = 32'h10a0ffff;
      65518: inst = 32'hca0fff6;
      65519: inst = 32'h24822800;
      65520: inst = 32'h10a00000;
      65521: inst = 32'hca00004;
      65522: inst = 32'h38632800;
      65523: inst = 32'h38842800;
      65524: inst = 32'h10a00000;
      65525: inst = 32'hca0fff9;
      65526: inst = 32'h13e00001;
      65527: inst = 32'hfe0d96a;
      65528: inst = 32'h5be00000;
      65529: inst = 32'h8c50000;
      65530: inst = 32'h24612800;
      65531: inst = 32'h10a0ffff;
      65532: inst = 32'hca0fff6;
      65533: inst = 32'h24822800;
      65534: inst = 32'h10a00000;
      65535: inst = 32'hca00004;
      65536: inst = 32'h38632800;
      65537: inst = 32'h38842800;
      65538: inst = 32'h10a00001;
      65539: inst = 32'hca00007;
      65540: inst = 32'h13e00001;
      65541: inst = 32'hfe0d96a;
      65542: inst = 32'h5be00000;
      65543: inst = 32'h8c50000;
      65544: inst = 32'h24612800;
      65545: inst = 32'h10a0ffff;
      65546: inst = 32'hca0fff6;
      65547: inst = 32'h24822800;
      65548: inst = 32'h10a00000;
      65549: inst = 32'hca00004;
      65550: inst = 32'h38632800;
      65551: inst = 32'h38842800;
      65552: inst = 32'h10a00001;
      65553: inst = 32'hca00015;
      65554: inst = 32'h13e00001;
      65555: inst = 32'hfe0d96a;
      65556: inst = 32'h5be00000;
      65557: inst = 32'h8c50000;
      65558: inst = 32'h24612800;
      65559: inst = 32'h10a0ffff;
      65560: inst = 32'hca0fff6;
      65561: inst = 32'h24822800;
      65562: inst = 32'h10a00000;
      65563: inst = 32'hca00004;
      65564: inst = 32'h38632800;
      65565: inst = 32'h38842800;
      65566: inst = 32'h10a00001;
      65567: inst = 32'hca00023;
      65568: inst = 32'h13e00001;
      65569: inst = 32'hfe0d96a;
      65570: inst = 32'h5be00000;
      65571: inst = 32'h8c50000;
      65572: inst = 32'h24612800;
      65573: inst = 32'h10a0ffff;
      65574: inst = 32'hca0fff6;
      65575: inst = 32'h24822800;
      65576: inst = 32'h10a00000;
      65577: inst = 32'hca00004;
      65578: inst = 32'h38632800;
      65579: inst = 32'h38842800;
      65580: inst = 32'h10a00001;
      65581: inst = 32'hca00031;
      65582: inst = 32'h13e00001;
      65583: inst = 32'hfe0d96a;
      65584: inst = 32'h5be00000;
      65585: inst = 32'h8c50000;
      65586: inst = 32'h24612800;
      65587: inst = 32'h10a0ffff;
      65588: inst = 32'hca0fff6;
      65589: inst = 32'h24822800;
      65590: inst = 32'h10a00000;
      65591: inst = 32'hca00004;
      65592: inst = 32'h38632800;
      65593: inst = 32'h38842800;
      65594: inst = 32'h10a00001;
      65595: inst = 32'hca0003f;
      65596: inst = 32'h13e00001;
      65597: inst = 32'hfe0d96a;
      65598: inst = 32'h5be00000;
      65599: inst = 32'h8c50000;
      65600: inst = 32'h24612800;
      65601: inst = 32'h10a0ffff;
      65602: inst = 32'hca0fff6;
      65603: inst = 32'h24822800;
      65604: inst = 32'h10a00000;
      65605: inst = 32'hca00004;
      65606: inst = 32'h38632800;
      65607: inst = 32'h38842800;
      65608: inst = 32'h10a00001;
      65609: inst = 32'hca0004d;
      65610: inst = 32'h13e00001;
      65611: inst = 32'hfe0d96a;
      65612: inst = 32'h5be00000;
      65613: inst = 32'h8c50000;
      65614: inst = 32'h24612800;
      65615: inst = 32'h10a0ffff;
      65616: inst = 32'hca0fff6;
      65617: inst = 32'h24822800;
      65618: inst = 32'h10a00000;
      65619: inst = 32'hca00004;
      65620: inst = 32'h38632800;
      65621: inst = 32'h38842800;
      65622: inst = 32'h10a00001;
      65623: inst = 32'hca0005b;
      65624: inst = 32'h13e00001;
      65625: inst = 32'hfe0d96a;
      65626: inst = 32'h5be00000;
      65627: inst = 32'h8c50000;
      65628: inst = 32'h24612800;
      65629: inst = 32'h10a0ffff;
      65630: inst = 32'hca0fff6;
      65631: inst = 32'h24822800;
      65632: inst = 32'h10a00000;
      65633: inst = 32'hca00004;
      65634: inst = 32'h38632800;
      65635: inst = 32'h38842800;
      65636: inst = 32'h10a00001;
      65637: inst = 32'hca00069;
      65638: inst = 32'h13e00001;
      65639: inst = 32'hfe0d96a;
      65640: inst = 32'h5be00000;
      65641: inst = 32'h8c50000;
      65642: inst = 32'h24612800;
      65643: inst = 32'h10a0ffff;
      65644: inst = 32'hca0fff6;
      65645: inst = 32'h24822800;
      65646: inst = 32'h10a00000;
      65647: inst = 32'hca00004;
      65648: inst = 32'h38632800;
      65649: inst = 32'h38842800;
      65650: inst = 32'h10a00001;
      65651: inst = 32'hca00077;
      65652: inst = 32'h13e00001;
      65653: inst = 32'hfe0d96a;
      65654: inst = 32'h5be00000;
      65655: inst = 32'h8c50000;
      65656: inst = 32'h24612800;
      65657: inst = 32'h10a0ffff;
      65658: inst = 32'hca0fff6;
      65659: inst = 32'h24822800;
      65660: inst = 32'h10a00000;
      65661: inst = 32'hca00004;
      65662: inst = 32'h38632800;
      65663: inst = 32'h38842800;
      65664: inst = 32'h10a00001;
      65665: inst = 32'hca00085;
      65666: inst = 32'h13e00001;
      65667: inst = 32'hfe0d96a;
      65668: inst = 32'h5be00000;
      65669: inst = 32'h8c50000;
      65670: inst = 32'h24612800;
      65671: inst = 32'h10a0ffff;
      65672: inst = 32'hca0fff6;
      65673: inst = 32'h24822800;
      65674: inst = 32'h10a00000;
      65675: inst = 32'hca00004;
      65676: inst = 32'h38632800;
      65677: inst = 32'h38842800;
      65678: inst = 32'h10a00001;
      65679: inst = 32'hca00093;
      65680: inst = 32'h13e00001;
      65681: inst = 32'hfe0d96a;
      65682: inst = 32'h5be00000;
      65683: inst = 32'h8c50000;
      65684: inst = 32'h24612800;
      65685: inst = 32'h10a0ffff;
      65686: inst = 32'hca0fff6;
      65687: inst = 32'h24822800;
      65688: inst = 32'h10a00000;
      65689: inst = 32'hca00004;
      65690: inst = 32'h38632800;
      65691: inst = 32'h38842800;
      65692: inst = 32'h10a00001;
      65693: inst = 32'hca000a1;
      65694: inst = 32'h13e00001;
      65695: inst = 32'hfe0d96a;
      65696: inst = 32'h5be00000;
      65697: inst = 32'h8c50000;
      65698: inst = 32'h24612800;
      65699: inst = 32'h10a0ffff;
      65700: inst = 32'hca0fff6;
      65701: inst = 32'h24822800;
      65702: inst = 32'h10a00000;
      65703: inst = 32'hca00004;
      65704: inst = 32'h38632800;
      65705: inst = 32'h38842800;
      65706: inst = 32'h10a00001;
      65707: inst = 32'hca000af;
      65708: inst = 32'h13e00001;
      65709: inst = 32'hfe0d96a;
      65710: inst = 32'h5be00000;
      65711: inst = 32'h8c50000;
      65712: inst = 32'h24612800;
      65713: inst = 32'h10a0ffff;
      65714: inst = 32'hca0fff6;
      65715: inst = 32'h24822800;
      65716: inst = 32'h10a00000;
      65717: inst = 32'hca00004;
      65718: inst = 32'h38632800;
      65719: inst = 32'h38842800;
      65720: inst = 32'h10a00001;
      65721: inst = 32'hca000bd;
      65722: inst = 32'h13e00001;
      65723: inst = 32'hfe0d96a;
      65724: inst = 32'h5be00000;
      65725: inst = 32'h8c50000;
      65726: inst = 32'h24612800;
      65727: inst = 32'h10a0ffff;
      65728: inst = 32'hca0fff6;
      65729: inst = 32'h24822800;
      65730: inst = 32'h10a00000;
      65731: inst = 32'hca00004;
      65732: inst = 32'h38632800;
      65733: inst = 32'h38842800;
      65734: inst = 32'h10a00001;
      65735: inst = 32'hca000cb;
      65736: inst = 32'h13e00001;
      65737: inst = 32'hfe0d96a;
      65738: inst = 32'h5be00000;
      65739: inst = 32'h8c50000;
      65740: inst = 32'h24612800;
      65741: inst = 32'h10a0ffff;
      65742: inst = 32'hca0fff6;
      65743: inst = 32'h24822800;
      65744: inst = 32'h10a00000;
      65745: inst = 32'hca00004;
      65746: inst = 32'h38632800;
      65747: inst = 32'h38842800;
      65748: inst = 32'h10a00001;
      65749: inst = 32'hca000d9;
      65750: inst = 32'h13e00001;
      65751: inst = 32'hfe0d96a;
      65752: inst = 32'h5be00000;
      65753: inst = 32'h8c50000;
      65754: inst = 32'h24612800;
      65755: inst = 32'h10a0ffff;
      65756: inst = 32'hca0fff6;
      65757: inst = 32'h24822800;
      65758: inst = 32'h10a00000;
      65759: inst = 32'hca00004;
      65760: inst = 32'h38632800;
      65761: inst = 32'h38842800;
      65762: inst = 32'h10a00001;
      65763: inst = 32'hca000e7;
      65764: inst = 32'h13e00001;
      65765: inst = 32'hfe0d96a;
      65766: inst = 32'h5be00000;
      65767: inst = 32'h8c50000;
      65768: inst = 32'h24612800;
      65769: inst = 32'h10a0ffff;
      65770: inst = 32'hca0fff6;
      65771: inst = 32'h24822800;
      65772: inst = 32'h10a00000;
      65773: inst = 32'hca00004;
      65774: inst = 32'h38632800;
      65775: inst = 32'h38842800;
      65776: inst = 32'h10a00001;
      65777: inst = 32'hca000f5;
      65778: inst = 32'h13e00001;
      65779: inst = 32'hfe0d96a;
      65780: inst = 32'h5be00000;
      65781: inst = 32'h8c50000;
      65782: inst = 32'h24612800;
      65783: inst = 32'h10a0ffff;
      65784: inst = 32'hca0fff6;
      65785: inst = 32'h24822800;
      65786: inst = 32'h10a00000;
      65787: inst = 32'hca00004;
      65788: inst = 32'h38632800;
      65789: inst = 32'h38842800;
      65790: inst = 32'h10a00001;
      65791: inst = 32'hca00103;
      65792: inst = 32'h13e00001;
      65793: inst = 32'hfe0d96a;
      65794: inst = 32'h5be00000;
      65795: inst = 32'h8c50000;
      65796: inst = 32'h24612800;
      65797: inst = 32'h10a0ffff;
      65798: inst = 32'hca0fff6;
      65799: inst = 32'h24822800;
      65800: inst = 32'h10a00000;
      65801: inst = 32'hca00004;
      65802: inst = 32'h38632800;
      65803: inst = 32'h38842800;
      65804: inst = 32'h10a00001;
      65805: inst = 32'hca00111;
      65806: inst = 32'h13e00001;
      65807: inst = 32'hfe0d96a;
      65808: inst = 32'h5be00000;
      65809: inst = 32'h8c50000;
      65810: inst = 32'h24612800;
      65811: inst = 32'h10a0ffff;
      65812: inst = 32'hca0fff6;
      65813: inst = 32'h24822800;
      65814: inst = 32'h10a00000;
      65815: inst = 32'hca00004;
      65816: inst = 32'h38632800;
      65817: inst = 32'h38842800;
      65818: inst = 32'h10a00001;
      65819: inst = 32'hca0011f;
      65820: inst = 32'h13e00001;
      65821: inst = 32'hfe0d96a;
      65822: inst = 32'h5be00000;
      65823: inst = 32'h8c50000;
      65824: inst = 32'h24612800;
      65825: inst = 32'h10a0ffff;
      65826: inst = 32'hca0fff6;
      65827: inst = 32'h24822800;
      65828: inst = 32'h10a00000;
      65829: inst = 32'hca00004;
      65830: inst = 32'h38632800;
      65831: inst = 32'h38842800;
      65832: inst = 32'h10a00001;
      65833: inst = 32'hca0012d;
      65834: inst = 32'h13e00001;
      65835: inst = 32'hfe0d96a;
      65836: inst = 32'h5be00000;
      65837: inst = 32'h8c50000;
      65838: inst = 32'h24612800;
      65839: inst = 32'h10a0ffff;
      65840: inst = 32'hca0fff6;
      65841: inst = 32'h24822800;
      65842: inst = 32'h10a00000;
      65843: inst = 32'hca00004;
      65844: inst = 32'h38632800;
      65845: inst = 32'h38842800;
      65846: inst = 32'h10a00001;
      65847: inst = 32'hca0013b;
      65848: inst = 32'h13e00001;
      65849: inst = 32'hfe0d96a;
      65850: inst = 32'h5be00000;
      65851: inst = 32'h8c50000;
      65852: inst = 32'h24612800;
      65853: inst = 32'h10a0ffff;
      65854: inst = 32'hca0fff6;
      65855: inst = 32'h24822800;
      65856: inst = 32'h10a00000;
      65857: inst = 32'hca00004;
      65858: inst = 32'h38632800;
      65859: inst = 32'h38842800;
      65860: inst = 32'h10a00001;
      65861: inst = 32'hca00149;
      65862: inst = 32'h13e00001;
      65863: inst = 32'hfe0d96a;
      65864: inst = 32'h5be00000;
      65865: inst = 32'h8c50000;
      65866: inst = 32'h24612800;
      65867: inst = 32'h10a0ffff;
      65868: inst = 32'hca0fff6;
      65869: inst = 32'h24822800;
      65870: inst = 32'h10a00000;
      65871: inst = 32'hca00004;
      65872: inst = 32'h38632800;
      65873: inst = 32'h38842800;
      65874: inst = 32'h10a00001;
      65875: inst = 32'hca00157;
      65876: inst = 32'h13e00001;
      65877: inst = 32'hfe0d96a;
      65878: inst = 32'h5be00000;
      65879: inst = 32'h8c50000;
      65880: inst = 32'h24612800;
      65881: inst = 32'h10a0ffff;
      65882: inst = 32'hca0fff6;
      65883: inst = 32'h24822800;
      65884: inst = 32'h10a00000;
      65885: inst = 32'hca00004;
      65886: inst = 32'h38632800;
      65887: inst = 32'h38842800;
      65888: inst = 32'h10a00001;
      65889: inst = 32'hca00165;
      65890: inst = 32'h13e00001;
      65891: inst = 32'hfe0d96a;
      65892: inst = 32'h5be00000;
      65893: inst = 32'h8c50000;
      65894: inst = 32'h24612800;
      65895: inst = 32'h10a0ffff;
      65896: inst = 32'hca0fff6;
      65897: inst = 32'h24822800;
      65898: inst = 32'h10a00000;
      65899: inst = 32'hca00004;
      65900: inst = 32'h38632800;
      65901: inst = 32'h38842800;
      65902: inst = 32'h10a00001;
      65903: inst = 32'hca00173;
      65904: inst = 32'h13e00001;
      65905: inst = 32'hfe0d96a;
      65906: inst = 32'h5be00000;
      65907: inst = 32'h8c50000;
      65908: inst = 32'h24612800;
      65909: inst = 32'h10a0ffff;
      65910: inst = 32'hca0fff6;
      65911: inst = 32'h24822800;
      65912: inst = 32'h10a00000;
      65913: inst = 32'hca00004;
      65914: inst = 32'h38632800;
      65915: inst = 32'h38842800;
      65916: inst = 32'h10a00001;
      65917: inst = 32'hca00181;
      65918: inst = 32'h13e00001;
      65919: inst = 32'hfe0d96a;
      65920: inst = 32'h5be00000;
      65921: inst = 32'h8c50000;
      65922: inst = 32'h24612800;
      65923: inst = 32'h10a0ffff;
      65924: inst = 32'hca0fff6;
      65925: inst = 32'h24822800;
      65926: inst = 32'h10a00000;
      65927: inst = 32'hca00004;
      65928: inst = 32'h38632800;
      65929: inst = 32'h38842800;
      65930: inst = 32'h10a00001;
      65931: inst = 32'hca0018f;
      65932: inst = 32'h13e00001;
      65933: inst = 32'hfe0d96a;
      65934: inst = 32'h5be00000;
      65935: inst = 32'h8c50000;
      65936: inst = 32'h24612800;
      65937: inst = 32'h10a0ffff;
      65938: inst = 32'hca0fff6;
      65939: inst = 32'h24822800;
      65940: inst = 32'h10a00000;
      65941: inst = 32'hca00004;
      65942: inst = 32'h38632800;
      65943: inst = 32'h38842800;
      65944: inst = 32'h10a00001;
      65945: inst = 32'hca0019d;
      65946: inst = 32'h13e00001;
      65947: inst = 32'hfe0d96a;
      65948: inst = 32'h5be00000;
      65949: inst = 32'h8c50000;
      65950: inst = 32'h24612800;
      65951: inst = 32'h10a0ffff;
      65952: inst = 32'hca0fff6;
      65953: inst = 32'h24822800;
      65954: inst = 32'h10a00000;
      65955: inst = 32'hca00004;
      65956: inst = 32'h38632800;
      65957: inst = 32'h38842800;
      65958: inst = 32'h10a00001;
      65959: inst = 32'hca001ab;
      65960: inst = 32'h13e00001;
      65961: inst = 32'hfe0d96a;
      65962: inst = 32'h5be00000;
      65963: inst = 32'h8c50000;
      65964: inst = 32'h24612800;
      65965: inst = 32'h10a0ffff;
      65966: inst = 32'hca0fff6;
      65967: inst = 32'h24822800;
      65968: inst = 32'h10a00000;
      65969: inst = 32'hca00004;
      65970: inst = 32'h38632800;
      65971: inst = 32'h38842800;
      65972: inst = 32'h10a00001;
      65973: inst = 32'hca001b9;
      65974: inst = 32'h13e00001;
      65975: inst = 32'hfe0d96a;
      65976: inst = 32'h5be00000;
      65977: inst = 32'h8c50000;
      65978: inst = 32'h24612800;
      65979: inst = 32'h10a0ffff;
      65980: inst = 32'hca0fff6;
      65981: inst = 32'h24822800;
      65982: inst = 32'h10a00000;
      65983: inst = 32'hca00004;
      65984: inst = 32'h38632800;
      65985: inst = 32'h38842800;
      65986: inst = 32'h10a00001;
      65987: inst = 32'hca001c7;
      65988: inst = 32'h13e00001;
      65989: inst = 32'hfe0d96a;
      65990: inst = 32'h5be00000;
      65991: inst = 32'h8c50000;
      65992: inst = 32'h24612800;
      65993: inst = 32'h10a0ffff;
      65994: inst = 32'hca0fff6;
      65995: inst = 32'h24822800;
      65996: inst = 32'h10a00000;
      65997: inst = 32'hca00004;
      65998: inst = 32'h38632800;
      65999: inst = 32'h38842800;
      66000: inst = 32'h10a00001;
      66001: inst = 32'hca001d5;
      66002: inst = 32'h13e00001;
      66003: inst = 32'hfe0d96a;
      66004: inst = 32'h5be00000;
      66005: inst = 32'h8c50000;
      66006: inst = 32'h24612800;
      66007: inst = 32'h10a0ffff;
      66008: inst = 32'hca0fff6;
      66009: inst = 32'h24822800;
      66010: inst = 32'h10a00000;
      66011: inst = 32'hca00004;
      66012: inst = 32'h38632800;
      66013: inst = 32'h38842800;
      66014: inst = 32'h10a00001;
      66015: inst = 32'hca001e3;
      66016: inst = 32'h13e00001;
      66017: inst = 32'hfe0d96a;
      66018: inst = 32'h5be00000;
      66019: inst = 32'h8c50000;
      66020: inst = 32'h24612800;
      66021: inst = 32'h10a0ffff;
      66022: inst = 32'hca0fff6;
      66023: inst = 32'h24822800;
      66024: inst = 32'h10a00000;
      66025: inst = 32'hca00004;
      66026: inst = 32'h38632800;
      66027: inst = 32'h38842800;
      66028: inst = 32'h10a00001;
      66029: inst = 32'hca001f1;
      66030: inst = 32'h13e00001;
      66031: inst = 32'hfe0d96a;
      66032: inst = 32'h5be00000;
      66033: inst = 32'h8c50000;
      66034: inst = 32'h24612800;
      66035: inst = 32'h10a0ffff;
      66036: inst = 32'hca0fff6;
      66037: inst = 32'h24822800;
      66038: inst = 32'h10a00000;
      66039: inst = 32'hca00004;
      66040: inst = 32'h38632800;
      66041: inst = 32'h38842800;
      66042: inst = 32'h10a00001;
      66043: inst = 32'hca001ff;
      66044: inst = 32'h13e00001;
      66045: inst = 32'hfe0d96a;
      66046: inst = 32'h5be00000;
      66047: inst = 32'h8c50000;
      66048: inst = 32'h24612800;
      66049: inst = 32'h10a0ffff;
      66050: inst = 32'hca0fff6;
      66051: inst = 32'h24822800;
      66052: inst = 32'h10a00000;
      66053: inst = 32'hca00004;
      66054: inst = 32'h38632800;
      66055: inst = 32'h38842800;
      66056: inst = 32'h10a00001;
      66057: inst = 32'hca0020d;
      66058: inst = 32'h13e00001;
      66059: inst = 32'hfe0d96a;
      66060: inst = 32'h5be00000;
      66061: inst = 32'h8c50000;
      66062: inst = 32'h24612800;
      66063: inst = 32'h10a0ffff;
      66064: inst = 32'hca0fff6;
      66065: inst = 32'h24822800;
      66066: inst = 32'h10a00000;
      66067: inst = 32'hca00004;
      66068: inst = 32'h38632800;
      66069: inst = 32'h38842800;
      66070: inst = 32'h10a00001;
      66071: inst = 32'hca0021b;
      66072: inst = 32'h13e00001;
      66073: inst = 32'hfe0d96a;
      66074: inst = 32'h5be00000;
      66075: inst = 32'h8c50000;
      66076: inst = 32'h24612800;
      66077: inst = 32'h10a0ffff;
      66078: inst = 32'hca0fff6;
      66079: inst = 32'h24822800;
      66080: inst = 32'h10a00000;
      66081: inst = 32'hca00004;
      66082: inst = 32'h38632800;
      66083: inst = 32'h38842800;
      66084: inst = 32'h10a00001;
      66085: inst = 32'hca00229;
      66086: inst = 32'h13e00001;
      66087: inst = 32'hfe0d96a;
      66088: inst = 32'h5be00000;
      66089: inst = 32'h8c50000;
      66090: inst = 32'h24612800;
      66091: inst = 32'h10a0ffff;
      66092: inst = 32'hca0fff7;
      66093: inst = 32'h24822800;
      66094: inst = 32'h10a00000;
      66095: inst = 32'hca00004;
      66096: inst = 32'h38632800;
      66097: inst = 32'h38842800;
      66098: inst = 32'h10a00001;
      66099: inst = 32'hca00237;
      66100: inst = 32'h13e00001;
      66101: inst = 32'hfe0d96a;
      66102: inst = 32'h5be00000;
      66103: inst = 32'h8c50000;
      66104: inst = 32'h24612800;
      66105: inst = 32'h10a0ffff;
      66106: inst = 32'hca0fff7;
      66107: inst = 32'h24822800;
      66108: inst = 32'h10a00000;
      66109: inst = 32'hca00004;
      66110: inst = 32'h38632800;
      66111: inst = 32'h38842800;
      66112: inst = 32'h10a00001;
      66113: inst = 32'hca00245;
      66114: inst = 32'h13e00001;
      66115: inst = 32'hfe0d96a;
      66116: inst = 32'h5be00000;
      66117: inst = 32'h8c50000;
      66118: inst = 32'h24612800;
      66119: inst = 32'h10a0ffff;
      66120: inst = 32'hca0fff7;
      66121: inst = 32'h24822800;
      66122: inst = 32'h10a00000;
      66123: inst = 32'hca00004;
      66124: inst = 32'h38632800;
      66125: inst = 32'h38842800;
      66126: inst = 32'h10a00001;
      66127: inst = 32'hca00253;
      66128: inst = 32'h13e00001;
      66129: inst = 32'hfe0d96a;
      66130: inst = 32'h5be00000;
      66131: inst = 32'h8c50000;
      66132: inst = 32'h24612800;
      66133: inst = 32'h10a0ffff;
      66134: inst = 32'hca0fff7;
      66135: inst = 32'h24822800;
      66136: inst = 32'h10a00000;
      66137: inst = 32'hca00004;
      66138: inst = 32'h38632800;
      66139: inst = 32'h38842800;
      66140: inst = 32'h10a00001;
      66141: inst = 32'hca00261;
      66142: inst = 32'h13e00001;
      66143: inst = 32'hfe0d96a;
      66144: inst = 32'h5be00000;
      66145: inst = 32'h8c50000;
      66146: inst = 32'h24612800;
      66147: inst = 32'h10a0ffff;
      66148: inst = 32'hca0fff7;
      66149: inst = 32'h24822800;
      66150: inst = 32'h10a00000;
      66151: inst = 32'hca00004;
      66152: inst = 32'h38632800;
      66153: inst = 32'h38842800;
      66154: inst = 32'h10a00001;
      66155: inst = 32'hca0026f;
      66156: inst = 32'h13e00001;
      66157: inst = 32'hfe0d96a;
      66158: inst = 32'h5be00000;
      66159: inst = 32'h8c50000;
      66160: inst = 32'h24612800;
      66161: inst = 32'h10a0ffff;
      66162: inst = 32'hca0fff7;
      66163: inst = 32'h24822800;
      66164: inst = 32'h10a00000;
      66165: inst = 32'hca00004;
      66166: inst = 32'h38632800;
      66167: inst = 32'h38842800;
      66168: inst = 32'h10a00001;
      66169: inst = 32'hca0027d;
      66170: inst = 32'h13e00001;
      66171: inst = 32'hfe0d96a;
      66172: inst = 32'h5be00000;
      66173: inst = 32'h8c50000;
      66174: inst = 32'h24612800;
      66175: inst = 32'h10a0ffff;
      66176: inst = 32'hca0fff7;
      66177: inst = 32'h24822800;
      66178: inst = 32'h10a00000;
      66179: inst = 32'hca00004;
      66180: inst = 32'h38632800;
      66181: inst = 32'h38842800;
      66182: inst = 32'h10a00001;
      66183: inst = 32'hca0028b;
      66184: inst = 32'h13e00001;
      66185: inst = 32'hfe0d96a;
      66186: inst = 32'h5be00000;
      66187: inst = 32'h8c50000;
      66188: inst = 32'h24612800;
      66189: inst = 32'h10a0ffff;
      66190: inst = 32'hca0fff7;
      66191: inst = 32'h24822800;
      66192: inst = 32'h10a00000;
      66193: inst = 32'hca00004;
      66194: inst = 32'h38632800;
      66195: inst = 32'h38842800;
      66196: inst = 32'h10a00001;
      66197: inst = 32'hca00299;
      66198: inst = 32'h13e00001;
      66199: inst = 32'hfe0d96a;
      66200: inst = 32'h5be00000;
      66201: inst = 32'h8c50000;
      66202: inst = 32'h24612800;
      66203: inst = 32'h10a0ffff;
      66204: inst = 32'hca0fff7;
      66205: inst = 32'h24822800;
      66206: inst = 32'h10a00000;
      66207: inst = 32'hca00004;
      66208: inst = 32'h38632800;
      66209: inst = 32'h38842800;
      66210: inst = 32'h10a00001;
      66211: inst = 32'hca002a7;
      66212: inst = 32'h13e00001;
      66213: inst = 32'hfe0d96a;
      66214: inst = 32'h5be00000;
      66215: inst = 32'h8c50000;
      66216: inst = 32'h24612800;
      66217: inst = 32'h10a0ffff;
      66218: inst = 32'hca0fff7;
      66219: inst = 32'h24822800;
      66220: inst = 32'h10a00000;
      66221: inst = 32'hca00004;
      66222: inst = 32'h38632800;
      66223: inst = 32'h38842800;
      66224: inst = 32'h10a00001;
      66225: inst = 32'hca002b5;
      66226: inst = 32'h13e00001;
      66227: inst = 32'hfe0d96a;
      66228: inst = 32'h5be00000;
      66229: inst = 32'h8c50000;
      66230: inst = 32'h24612800;
      66231: inst = 32'h10a0ffff;
      66232: inst = 32'hca0fff7;
      66233: inst = 32'h24822800;
      66234: inst = 32'h10a00000;
      66235: inst = 32'hca00004;
      66236: inst = 32'h38632800;
      66237: inst = 32'h38842800;
      66238: inst = 32'h10a00001;
      66239: inst = 32'hca002c3;
      66240: inst = 32'h13e00001;
      66241: inst = 32'hfe0d96a;
      66242: inst = 32'h5be00000;
      66243: inst = 32'h8c50000;
      66244: inst = 32'h24612800;
      66245: inst = 32'h10a0ffff;
      66246: inst = 32'hca0fff7;
      66247: inst = 32'h24822800;
      66248: inst = 32'h10a00000;
      66249: inst = 32'hca00004;
      66250: inst = 32'h38632800;
      66251: inst = 32'h38842800;
      66252: inst = 32'h10a00001;
      66253: inst = 32'hca002d1;
      66254: inst = 32'h13e00001;
      66255: inst = 32'hfe0d96a;
      66256: inst = 32'h5be00000;
      66257: inst = 32'h8c50000;
      66258: inst = 32'h24612800;
      66259: inst = 32'h10a0ffff;
      66260: inst = 32'hca0fff7;
      66261: inst = 32'h24822800;
      66262: inst = 32'h10a00000;
      66263: inst = 32'hca00004;
      66264: inst = 32'h38632800;
      66265: inst = 32'h38842800;
      66266: inst = 32'h10a00001;
      66267: inst = 32'hca002df;
      66268: inst = 32'h13e00001;
      66269: inst = 32'hfe0d96a;
      66270: inst = 32'h5be00000;
      66271: inst = 32'h8c50000;
      66272: inst = 32'h24612800;
      66273: inst = 32'h10a0ffff;
      66274: inst = 32'hca0fff7;
      66275: inst = 32'h24822800;
      66276: inst = 32'h10a00000;
      66277: inst = 32'hca00004;
      66278: inst = 32'h38632800;
      66279: inst = 32'h38842800;
      66280: inst = 32'h10a00001;
      66281: inst = 32'hca002ed;
      66282: inst = 32'h13e00001;
      66283: inst = 32'hfe0d96a;
      66284: inst = 32'h5be00000;
      66285: inst = 32'h8c50000;
      66286: inst = 32'h24612800;
      66287: inst = 32'h10a0ffff;
      66288: inst = 32'hca0fff7;
      66289: inst = 32'h24822800;
      66290: inst = 32'h10a00000;
      66291: inst = 32'hca00004;
      66292: inst = 32'h38632800;
      66293: inst = 32'h38842800;
      66294: inst = 32'h10a00001;
      66295: inst = 32'hca002fb;
      66296: inst = 32'h13e00001;
      66297: inst = 32'hfe0d96a;
      66298: inst = 32'h5be00000;
      66299: inst = 32'h8c50000;
      66300: inst = 32'h24612800;
      66301: inst = 32'h10a0ffff;
      66302: inst = 32'hca0fff7;
      66303: inst = 32'h24822800;
      66304: inst = 32'h10a00000;
      66305: inst = 32'hca00004;
      66306: inst = 32'h38632800;
      66307: inst = 32'h38842800;
      66308: inst = 32'h10a00001;
      66309: inst = 32'hca00309;
      66310: inst = 32'h13e00001;
      66311: inst = 32'hfe0d96a;
      66312: inst = 32'h5be00000;
      66313: inst = 32'h8c50000;
      66314: inst = 32'h24612800;
      66315: inst = 32'h10a0ffff;
      66316: inst = 32'hca0fff7;
      66317: inst = 32'h24822800;
      66318: inst = 32'h10a00000;
      66319: inst = 32'hca00004;
      66320: inst = 32'h38632800;
      66321: inst = 32'h38842800;
      66322: inst = 32'h10a00001;
      66323: inst = 32'hca00317;
      66324: inst = 32'h13e00001;
      66325: inst = 32'hfe0d96a;
      66326: inst = 32'h5be00000;
      66327: inst = 32'h8c50000;
      66328: inst = 32'h24612800;
      66329: inst = 32'h10a0ffff;
      66330: inst = 32'hca0fff7;
      66331: inst = 32'h24822800;
      66332: inst = 32'h10a00000;
      66333: inst = 32'hca00004;
      66334: inst = 32'h38632800;
      66335: inst = 32'h38842800;
      66336: inst = 32'h10a00001;
      66337: inst = 32'hca00325;
      66338: inst = 32'h13e00001;
      66339: inst = 32'hfe0d96a;
      66340: inst = 32'h5be00000;
      66341: inst = 32'h8c50000;
      66342: inst = 32'h24612800;
      66343: inst = 32'h10a0ffff;
      66344: inst = 32'hca0fff7;
      66345: inst = 32'h24822800;
      66346: inst = 32'h10a00000;
      66347: inst = 32'hca00004;
      66348: inst = 32'h38632800;
      66349: inst = 32'h38842800;
      66350: inst = 32'h10a00001;
      66351: inst = 32'hca00333;
      66352: inst = 32'h13e00001;
      66353: inst = 32'hfe0d96a;
      66354: inst = 32'h5be00000;
      66355: inst = 32'h8c50000;
      66356: inst = 32'h24612800;
      66357: inst = 32'h10a0ffff;
      66358: inst = 32'hca0fff7;
      66359: inst = 32'h24822800;
      66360: inst = 32'h10a00000;
      66361: inst = 32'hca00004;
      66362: inst = 32'h38632800;
      66363: inst = 32'h38842800;
      66364: inst = 32'h10a00001;
      66365: inst = 32'hca00341;
      66366: inst = 32'h13e00001;
      66367: inst = 32'hfe0d96a;
      66368: inst = 32'h5be00000;
      66369: inst = 32'h8c50000;
      66370: inst = 32'h24612800;
      66371: inst = 32'h10a0ffff;
      66372: inst = 32'hca0fff7;
      66373: inst = 32'h24822800;
      66374: inst = 32'h10a00000;
      66375: inst = 32'hca00004;
      66376: inst = 32'h38632800;
      66377: inst = 32'h38842800;
      66378: inst = 32'h10a00001;
      66379: inst = 32'hca0034f;
      66380: inst = 32'h13e00001;
      66381: inst = 32'hfe0d96a;
      66382: inst = 32'h5be00000;
      66383: inst = 32'h8c50000;
      66384: inst = 32'h24612800;
      66385: inst = 32'h10a0ffff;
      66386: inst = 32'hca0fff7;
      66387: inst = 32'h24822800;
      66388: inst = 32'h10a00000;
      66389: inst = 32'hca00004;
      66390: inst = 32'h38632800;
      66391: inst = 32'h38842800;
      66392: inst = 32'h10a00001;
      66393: inst = 32'hca0035d;
      66394: inst = 32'h13e00001;
      66395: inst = 32'hfe0d96a;
      66396: inst = 32'h5be00000;
      66397: inst = 32'h8c50000;
      66398: inst = 32'h24612800;
      66399: inst = 32'h10a0ffff;
      66400: inst = 32'hca0fff7;
      66401: inst = 32'h24822800;
      66402: inst = 32'h10a00000;
      66403: inst = 32'hca00004;
      66404: inst = 32'h38632800;
      66405: inst = 32'h38842800;
      66406: inst = 32'h10a00001;
      66407: inst = 32'hca0036b;
      66408: inst = 32'h13e00001;
      66409: inst = 32'hfe0d96a;
      66410: inst = 32'h5be00000;
      66411: inst = 32'h8c50000;
      66412: inst = 32'h24612800;
      66413: inst = 32'h10a0ffff;
      66414: inst = 32'hca0fff7;
      66415: inst = 32'h24822800;
      66416: inst = 32'h10a00000;
      66417: inst = 32'hca00004;
      66418: inst = 32'h38632800;
      66419: inst = 32'h38842800;
      66420: inst = 32'h10a00001;
      66421: inst = 32'hca00379;
      66422: inst = 32'h13e00001;
      66423: inst = 32'hfe0d96a;
      66424: inst = 32'h5be00000;
      66425: inst = 32'h8c50000;
      66426: inst = 32'h24612800;
      66427: inst = 32'h10a0ffff;
      66428: inst = 32'hca0fff7;
      66429: inst = 32'h24822800;
      66430: inst = 32'h10a00000;
      66431: inst = 32'hca00004;
      66432: inst = 32'h38632800;
      66433: inst = 32'h38842800;
      66434: inst = 32'h10a00001;
      66435: inst = 32'hca00387;
      66436: inst = 32'h13e00001;
      66437: inst = 32'hfe0d96a;
      66438: inst = 32'h5be00000;
      66439: inst = 32'h8c50000;
      66440: inst = 32'h24612800;
      66441: inst = 32'h10a0ffff;
      66442: inst = 32'hca0fff7;
      66443: inst = 32'h24822800;
      66444: inst = 32'h10a00000;
      66445: inst = 32'hca00004;
      66446: inst = 32'h38632800;
      66447: inst = 32'h38842800;
      66448: inst = 32'h10a00001;
      66449: inst = 32'hca00395;
      66450: inst = 32'h13e00001;
      66451: inst = 32'hfe0d96a;
      66452: inst = 32'h5be00000;
      66453: inst = 32'h8c50000;
      66454: inst = 32'h24612800;
      66455: inst = 32'h10a0ffff;
      66456: inst = 32'hca0fff7;
      66457: inst = 32'h24822800;
      66458: inst = 32'h10a00000;
      66459: inst = 32'hca00004;
      66460: inst = 32'h38632800;
      66461: inst = 32'h38842800;
      66462: inst = 32'h10a00001;
      66463: inst = 32'hca003a3;
      66464: inst = 32'h13e00001;
      66465: inst = 32'hfe0d96a;
      66466: inst = 32'h5be00000;
      66467: inst = 32'h8c50000;
      66468: inst = 32'h24612800;
      66469: inst = 32'h10a0ffff;
      66470: inst = 32'hca0fff7;
      66471: inst = 32'h24822800;
      66472: inst = 32'h10a00000;
      66473: inst = 32'hca00004;
      66474: inst = 32'h38632800;
      66475: inst = 32'h38842800;
      66476: inst = 32'h10a00001;
      66477: inst = 32'hca003b1;
      66478: inst = 32'h13e00001;
      66479: inst = 32'hfe0d96a;
      66480: inst = 32'h5be00000;
      66481: inst = 32'h8c50000;
      66482: inst = 32'h24612800;
      66483: inst = 32'h10a0ffff;
      66484: inst = 32'hca0fff7;
      66485: inst = 32'h24822800;
      66486: inst = 32'h10a00000;
      66487: inst = 32'hca00004;
      66488: inst = 32'h38632800;
      66489: inst = 32'h38842800;
      66490: inst = 32'h10a00001;
      66491: inst = 32'hca003bf;
      66492: inst = 32'h13e00001;
      66493: inst = 32'hfe0d96a;
      66494: inst = 32'h5be00000;
      66495: inst = 32'h8c50000;
      66496: inst = 32'h24612800;
      66497: inst = 32'h10a0ffff;
      66498: inst = 32'hca0fff7;
      66499: inst = 32'h24822800;
      66500: inst = 32'h10a00000;
      66501: inst = 32'hca00004;
      66502: inst = 32'h38632800;
      66503: inst = 32'h38842800;
      66504: inst = 32'h10a00001;
      66505: inst = 32'hca003cd;
      66506: inst = 32'h13e00001;
      66507: inst = 32'hfe0d96a;
      66508: inst = 32'h5be00000;
      66509: inst = 32'h8c50000;
      66510: inst = 32'h24612800;
      66511: inst = 32'h10a0ffff;
      66512: inst = 32'hca0fff7;
      66513: inst = 32'h24822800;
      66514: inst = 32'h10a00000;
      66515: inst = 32'hca00004;
      66516: inst = 32'h38632800;
      66517: inst = 32'h38842800;
      66518: inst = 32'h10a00001;
      66519: inst = 32'hca003db;
      66520: inst = 32'h13e00001;
      66521: inst = 32'hfe0d96a;
      66522: inst = 32'h5be00000;
      66523: inst = 32'h8c50000;
      66524: inst = 32'h24612800;
      66525: inst = 32'h10a0ffff;
      66526: inst = 32'hca0fff7;
      66527: inst = 32'h24822800;
      66528: inst = 32'h10a00000;
      66529: inst = 32'hca00004;
      66530: inst = 32'h38632800;
      66531: inst = 32'h38842800;
      66532: inst = 32'h10a00001;
      66533: inst = 32'hca003e9;
      66534: inst = 32'h13e00001;
      66535: inst = 32'hfe0d96a;
      66536: inst = 32'h5be00000;
      66537: inst = 32'h8c50000;
      66538: inst = 32'h24612800;
      66539: inst = 32'h10a0ffff;
      66540: inst = 32'hca0fff7;
      66541: inst = 32'h24822800;
      66542: inst = 32'h10a00000;
      66543: inst = 32'hca00004;
      66544: inst = 32'h38632800;
      66545: inst = 32'h38842800;
      66546: inst = 32'h10a00001;
      66547: inst = 32'hca003f7;
      66548: inst = 32'h13e00001;
      66549: inst = 32'hfe0d96a;
      66550: inst = 32'h5be00000;
      66551: inst = 32'h8c50000;
      66552: inst = 32'h24612800;
      66553: inst = 32'h10a0ffff;
      66554: inst = 32'hca0fff7;
      66555: inst = 32'h24822800;
      66556: inst = 32'h10a00000;
      66557: inst = 32'hca00004;
      66558: inst = 32'h38632800;
      66559: inst = 32'h38842800;
      66560: inst = 32'h10a00001;
      66561: inst = 32'hca00405;
      66562: inst = 32'h13e00001;
      66563: inst = 32'hfe0d96a;
      66564: inst = 32'h5be00000;
      66565: inst = 32'h8c50000;
      66566: inst = 32'h24612800;
      66567: inst = 32'h10a0ffff;
      66568: inst = 32'hca0fff7;
      66569: inst = 32'h24822800;
      66570: inst = 32'h10a00000;
      66571: inst = 32'hca00004;
      66572: inst = 32'h38632800;
      66573: inst = 32'h38842800;
      66574: inst = 32'h10a00001;
      66575: inst = 32'hca00413;
      66576: inst = 32'h13e00001;
      66577: inst = 32'hfe0d96a;
      66578: inst = 32'h5be00000;
      66579: inst = 32'h8c50000;
      66580: inst = 32'h24612800;
      66581: inst = 32'h10a0ffff;
      66582: inst = 32'hca0fff7;
      66583: inst = 32'h24822800;
      66584: inst = 32'h10a00000;
      66585: inst = 32'hca00004;
      66586: inst = 32'h38632800;
      66587: inst = 32'h38842800;
      66588: inst = 32'h10a00001;
      66589: inst = 32'hca00421;
      66590: inst = 32'h13e00001;
      66591: inst = 32'hfe0d96a;
      66592: inst = 32'h5be00000;
      66593: inst = 32'h8c50000;
      66594: inst = 32'h24612800;
      66595: inst = 32'h10a0ffff;
      66596: inst = 32'hca0fff7;
      66597: inst = 32'h24822800;
      66598: inst = 32'h10a00000;
      66599: inst = 32'hca00004;
      66600: inst = 32'h38632800;
      66601: inst = 32'h38842800;
      66602: inst = 32'h10a00001;
      66603: inst = 32'hca0042f;
      66604: inst = 32'h13e00001;
      66605: inst = 32'hfe0d96a;
      66606: inst = 32'h5be00000;
      66607: inst = 32'h8c50000;
      66608: inst = 32'h24612800;
      66609: inst = 32'h10a0ffff;
      66610: inst = 32'hca0fff7;
      66611: inst = 32'h24822800;
      66612: inst = 32'h10a00000;
      66613: inst = 32'hca00004;
      66614: inst = 32'h38632800;
      66615: inst = 32'h38842800;
      66616: inst = 32'h10a00001;
      66617: inst = 32'hca0043d;
      66618: inst = 32'h13e00001;
      66619: inst = 32'hfe0d96a;
      66620: inst = 32'h5be00000;
      66621: inst = 32'h8c50000;
      66622: inst = 32'h24612800;
      66623: inst = 32'h10a0ffff;
      66624: inst = 32'hca0fff7;
      66625: inst = 32'h24822800;
      66626: inst = 32'h10a00000;
      66627: inst = 32'hca00004;
      66628: inst = 32'h38632800;
      66629: inst = 32'h38842800;
      66630: inst = 32'h10a00001;
      66631: inst = 32'hca0044b;
      66632: inst = 32'h13e00001;
      66633: inst = 32'hfe0d96a;
      66634: inst = 32'h5be00000;
      66635: inst = 32'h8c50000;
      66636: inst = 32'h24612800;
      66637: inst = 32'h10a0ffff;
      66638: inst = 32'hca0fff7;
      66639: inst = 32'h24822800;
      66640: inst = 32'h10a00000;
      66641: inst = 32'hca00004;
      66642: inst = 32'h38632800;
      66643: inst = 32'h38842800;
      66644: inst = 32'h10a00001;
      66645: inst = 32'hca00459;
      66646: inst = 32'h13e00001;
      66647: inst = 32'hfe0d96a;
      66648: inst = 32'h5be00000;
      66649: inst = 32'h8c50000;
      66650: inst = 32'h24612800;
      66651: inst = 32'h10a0ffff;
      66652: inst = 32'hca0fff7;
      66653: inst = 32'h24822800;
      66654: inst = 32'h10a00000;
      66655: inst = 32'hca00004;
      66656: inst = 32'h38632800;
      66657: inst = 32'h38842800;
      66658: inst = 32'h10a00001;
      66659: inst = 32'hca00467;
      66660: inst = 32'h13e00001;
      66661: inst = 32'hfe0d96a;
      66662: inst = 32'h5be00000;
      66663: inst = 32'h8c50000;
      66664: inst = 32'h24612800;
      66665: inst = 32'h10a0ffff;
      66666: inst = 32'hca0fff7;
      66667: inst = 32'h24822800;
      66668: inst = 32'h10a00000;
      66669: inst = 32'hca00004;
      66670: inst = 32'h38632800;
      66671: inst = 32'h38842800;
      66672: inst = 32'h10a00001;
      66673: inst = 32'hca00475;
      66674: inst = 32'h13e00001;
      66675: inst = 32'hfe0d96a;
      66676: inst = 32'h5be00000;
      66677: inst = 32'h8c50000;
      66678: inst = 32'h24612800;
      66679: inst = 32'h10a0ffff;
      66680: inst = 32'hca0fff7;
      66681: inst = 32'h24822800;
      66682: inst = 32'h10a00000;
      66683: inst = 32'hca00004;
      66684: inst = 32'h38632800;
      66685: inst = 32'h38842800;
      66686: inst = 32'h10a00001;
      66687: inst = 32'hca00483;
      66688: inst = 32'h13e00001;
      66689: inst = 32'hfe0d96a;
      66690: inst = 32'h5be00000;
      66691: inst = 32'h8c50000;
      66692: inst = 32'h24612800;
      66693: inst = 32'h10a0ffff;
      66694: inst = 32'hca0fff7;
      66695: inst = 32'h24822800;
      66696: inst = 32'h10a00000;
      66697: inst = 32'hca00004;
      66698: inst = 32'h38632800;
      66699: inst = 32'h38842800;
      66700: inst = 32'h10a00001;
      66701: inst = 32'hca00491;
      66702: inst = 32'h13e00001;
      66703: inst = 32'hfe0d96a;
      66704: inst = 32'h5be00000;
      66705: inst = 32'h8c50000;
      66706: inst = 32'h24612800;
      66707: inst = 32'h10a0ffff;
      66708: inst = 32'hca0fff7;
      66709: inst = 32'h24822800;
      66710: inst = 32'h10a00000;
      66711: inst = 32'hca00004;
      66712: inst = 32'h38632800;
      66713: inst = 32'h38842800;
      66714: inst = 32'h10a00001;
      66715: inst = 32'hca0049f;
      66716: inst = 32'h13e00001;
      66717: inst = 32'hfe0d96a;
      66718: inst = 32'h5be00000;
      66719: inst = 32'h8c50000;
      66720: inst = 32'h24612800;
      66721: inst = 32'h10a0ffff;
      66722: inst = 32'hca0fff7;
      66723: inst = 32'h24822800;
      66724: inst = 32'h10a00000;
      66725: inst = 32'hca00004;
      66726: inst = 32'h38632800;
      66727: inst = 32'h38842800;
      66728: inst = 32'h10a00001;
      66729: inst = 32'hca004ad;
      66730: inst = 32'h13e00001;
      66731: inst = 32'hfe0d96a;
      66732: inst = 32'h5be00000;
      66733: inst = 32'h8c50000;
      66734: inst = 32'h24612800;
      66735: inst = 32'h10a0ffff;
      66736: inst = 32'hca0fff7;
      66737: inst = 32'h24822800;
      66738: inst = 32'h10a00000;
      66739: inst = 32'hca00004;
      66740: inst = 32'h38632800;
      66741: inst = 32'h38842800;
      66742: inst = 32'h10a00001;
      66743: inst = 32'hca004bb;
      66744: inst = 32'h13e00001;
      66745: inst = 32'hfe0d96a;
      66746: inst = 32'h5be00000;
      66747: inst = 32'h8c50000;
      66748: inst = 32'h24612800;
      66749: inst = 32'h10a0ffff;
      66750: inst = 32'hca0fff7;
      66751: inst = 32'h24822800;
      66752: inst = 32'h10a00000;
      66753: inst = 32'hca00004;
      66754: inst = 32'h38632800;
      66755: inst = 32'h38842800;
      66756: inst = 32'h10a00001;
      66757: inst = 32'hca004c9;
      66758: inst = 32'h13e00001;
      66759: inst = 32'hfe0d96a;
      66760: inst = 32'h5be00000;
      66761: inst = 32'h8c50000;
      66762: inst = 32'h24612800;
      66763: inst = 32'h10a0ffff;
      66764: inst = 32'hca0fff7;
      66765: inst = 32'h24822800;
      66766: inst = 32'h10a00000;
      66767: inst = 32'hca00004;
      66768: inst = 32'h38632800;
      66769: inst = 32'h38842800;
      66770: inst = 32'h10a00001;
      66771: inst = 32'hca004d7;
      66772: inst = 32'h13e00001;
      66773: inst = 32'hfe0d96a;
      66774: inst = 32'h5be00000;
      66775: inst = 32'h8c50000;
      66776: inst = 32'h24612800;
      66777: inst = 32'h10a0ffff;
      66778: inst = 32'hca0fff7;
      66779: inst = 32'h24822800;
      66780: inst = 32'h10a00000;
      66781: inst = 32'hca00004;
      66782: inst = 32'h38632800;
      66783: inst = 32'h38842800;
      66784: inst = 32'h10a00001;
      66785: inst = 32'hca004e5;
      66786: inst = 32'h13e00001;
      66787: inst = 32'hfe0d96a;
      66788: inst = 32'h5be00000;
      66789: inst = 32'h8c50000;
      66790: inst = 32'h24612800;
      66791: inst = 32'h10a0ffff;
      66792: inst = 32'hca0fff7;
      66793: inst = 32'h24822800;
      66794: inst = 32'h10a00000;
      66795: inst = 32'hca00004;
      66796: inst = 32'h38632800;
      66797: inst = 32'h38842800;
      66798: inst = 32'h10a00001;
      66799: inst = 32'hca004f3;
      66800: inst = 32'h13e00001;
      66801: inst = 32'hfe0d96a;
      66802: inst = 32'h5be00000;
      66803: inst = 32'h8c50000;
      66804: inst = 32'h24612800;
      66805: inst = 32'h10a0ffff;
      66806: inst = 32'hca0fff7;
      66807: inst = 32'h24822800;
      66808: inst = 32'h10a00000;
      66809: inst = 32'hca00004;
      66810: inst = 32'h38632800;
      66811: inst = 32'h38842800;
      66812: inst = 32'h10a00001;
      66813: inst = 32'hca00501;
      66814: inst = 32'h13e00001;
      66815: inst = 32'hfe0d96a;
      66816: inst = 32'h5be00000;
      66817: inst = 32'h8c50000;
      66818: inst = 32'h24612800;
      66819: inst = 32'h10a0ffff;
      66820: inst = 32'hca0fff7;
      66821: inst = 32'h24822800;
      66822: inst = 32'h10a00000;
      66823: inst = 32'hca00004;
      66824: inst = 32'h38632800;
      66825: inst = 32'h38842800;
      66826: inst = 32'h10a00001;
      66827: inst = 32'hca0050f;
      66828: inst = 32'h13e00001;
      66829: inst = 32'hfe0d96a;
      66830: inst = 32'h5be00000;
      66831: inst = 32'h8c50000;
      66832: inst = 32'h24612800;
      66833: inst = 32'h10a0ffff;
      66834: inst = 32'hca0fff7;
      66835: inst = 32'h24822800;
      66836: inst = 32'h10a00000;
      66837: inst = 32'hca00004;
      66838: inst = 32'h38632800;
      66839: inst = 32'h38842800;
      66840: inst = 32'h10a00001;
      66841: inst = 32'hca0051d;
      66842: inst = 32'h13e00001;
      66843: inst = 32'hfe0d96a;
      66844: inst = 32'h5be00000;
      66845: inst = 32'h8c50000;
      66846: inst = 32'h24612800;
      66847: inst = 32'h10a0ffff;
      66848: inst = 32'hca0fff7;
      66849: inst = 32'h24822800;
      66850: inst = 32'h10a00000;
      66851: inst = 32'hca00004;
      66852: inst = 32'h38632800;
      66853: inst = 32'h38842800;
      66854: inst = 32'h10a00001;
      66855: inst = 32'hca0052b;
      66856: inst = 32'h13e00001;
      66857: inst = 32'hfe0d96a;
      66858: inst = 32'h5be00000;
      66859: inst = 32'h8c50000;
      66860: inst = 32'h24612800;
      66861: inst = 32'h10a0ffff;
      66862: inst = 32'hca0fff7;
      66863: inst = 32'h24822800;
      66864: inst = 32'h10a00000;
      66865: inst = 32'hca00004;
      66866: inst = 32'h38632800;
      66867: inst = 32'h38842800;
      66868: inst = 32'h10a00001;
      66869: inst = 32'hca00539;
      66870: inst = 32'h13e00001;
      66871: inst = 32'hfe0d96a;
      66872: inst = 32'h5be00000;
      66873: inst = 32'h8c50000;
      66874: inst = 32'h24612800;
      66875: inst = 32'h10a0ffff;
      66876: inst = 32'hca0fff7;
      66877: inst = 32'h24822800;
      66878: inst = 32'h10a00000;
      66879: inst = 32'hca00004;
      66880: inst = 32'h38632800;
      66881: inst = 32'h38842800;
      66882: inst = 32'h10a00001;
      66883: inst = 32'hca00547;
      66884: inst = 32'h13e00001;
      66885: inst = 32'hfe0d96a;
      66886: inst = 32'h5be00000;
      66887: inst = 32'h8c50000;
      66888: inst = 32'h24612800;
      66889: inst = 32'h10a0ffff;
      66890: inst = 32'hca0fff7;
      66891: inst = 32'h24822800;
      66892: inst = 32'h10a00000;
      66893: inst = 32'hca00004;
      66894: inst = 32'h38632800;
      66895: inst = 32'h38842800;
      66896: inst = 32'h10a00001;
      66897: inst = 32'hca00555;
      66898: inst = 32'h13e00001;
      66899: inst = 32'hfe0d96a;
      66900: inst = 32'h5be00000;
      66901: inst = 32'h8c50000;
      66902: inst = 32'h24612800;
      66903: inst = 32'h10a0ffff;
      66904: inst = 32'hca0fff7;
      66905: inst = 32'h24822800;
      66906: inst = 32'h10a00000;
      66907: inst = 32'hca00004;
      66908: inst = 32'h38632800;
      66909: inst = 32'h38842800;
      66910: inst = 32'h10a00001;
      66911: inst = 32'hca00563;
      66912: inst = 32'h13e00001;
      66913: inst = 32'hfe0d96a;
      66914: inst = 32'h5be00000;
      66915: inst = 32'h8c50000;
      66916: inst = 32'h24612800;
      66917: inst = 32'h10a0ffff;
      66918: inst = 32'hca0fff7;
      66919: inst = 32'h24822800;
      66920: inst = 32'h10a00000;
      66921: inst = 32'hca00004;
      66922: inst = 32'h38632800;
      66923: inst = 32'h38842800;
      66924: inst = 32'h10a00001;
      66925: inst = 32'hca00571;
      66926: inst = 32'h13e00001;
      66927: inst = 32'hfe0d96a;
      66928: inst = 32'h5be00000;
      66929: inst = 32'h8c50000;
      66930: inst = 32'h24612800;
      66931: inst = 32'h10a0ffff;
      66932: inst = 32'hca0fff7;
      66933: inst = 32'h24822800;
      66934: inst = 32'h10a00000;
      66935: inst = 32'hca00004;
      66936: inst = 32'h38632800;
      66937: inst = 32'h38842800;
      66938: inst = 32'h10a00001;
      66939: inst = 32'hca0057f;
      66940: inst = 32'h13e00001;
      66941: inst = 32'hfe0d96a;
      66942: inst = 32'h5be00000;
      66943: inst = 32'h8c50000;
      66944: inst = 32'h24612800;
      66945: inst = 32'h10a0ffff;
      66946: inst = 32'hca0fff7;
      66947: inst = 32'h24822800;
      66948: inst = 32'h10a00000;
      66949: inst = 32'hca00004;
      66950: inst = 32'h38632800;
      66951: inst = 32'h38842800;
      66952: inst = 32'h10a00001;
      66953: inst = 32'hca0058d;
      66954: inst = 32'h13e00001;
      66955: inst = 32'hfe0d96a;
      66956: inst = 32'h5be00000;
      66957: inst = 32'h8c50000;
      66958: inst = 32'h24612800;
      66959: inst = 32'h10a0ffff;
      66960: inst = 32'hca0fff7;
      66961: inst = 32'h24822800;
      66962: inst = 32'h10a00000;
      66963: inst = 32'hca00004;
      66964: inst = 32'h38632800;
      66965: inst = 32'h38842800;
      66966: inst = 32'h10a00001;
      66967: inst = 32'hca0059b;
      66968: inst = 32'h13e00001;
      66969: inst = 32'hfe0d96a;
      66970: inst = 32'h5be00000;
      66971: inst = 32'h8c50000;
      66972: inst = 32'h24612800;
      66973: inst = 32'h10a0ffff;
      66974: inst = 32'hca0fff7;
      66975: inst = 32'h24822800;
      66976: inst = 32'h10a00000;
      66977: inst = 32'hca00004;
      66978: inst = 32'h38632800;
      66979: inst = 32'h38842800;
      66980: inst = 32'h10a00001;
      66981: inst = 32'hca005a9;
      66982: inst = 32'h13e00001;
      66983: inst = 32'hfe0d96a;
      66984: inst = 32'h5be00000;
      66985: inst = 32'h8c50000;
      66986: inst = 32'h24612800;
      66987: inst = 32'h10a0ffff;
      66988: inst = 32'hca0fff7;
      66989: inst = 32'h24822800;
      66990: inst = 32'h10a00000;
      66991: inst = 32'hca00004;
      66992: inst = 32'h38632800;
      66993: inst = 32'h38842800;
      66994: inst = 32'h10a00001;
      66995: inst = 32'hca005b7;
      66996: inst = 32'h13e00001;
      66997: inst = 32'hfe0d96a;
      66998: inst = 32'h5be00000;
      66999: inst = 32'h8c50000;
      67000: inst = 32'h24612800;
      67001: inst = 32'h10a0ffff;
      67002: inst = 32'hca0fff7;
      67003: inst = 32'h24822800;
      67004: inst = 32'h10a00000;
      67005: inst = 32'hca00004;
      67006: inst = 32'h38632800;
      67007: inst = 32'h38842800;
      67008: inst = 32'h10a00001;
      67009: inst = 32'hca005c5;
      67010: inst = 32'h13e00001;
      67011: inst = 32'hfe0d96a;
      67012: inst = 32'h5be00000;
      67013: inst = 32'h8c50000;
      67014: inst = 32'h24612800;
      67015: inst = 32'h10a0ffff;
      67016: inst = 32'hca0fff7;
      67017: inst = 32'h24822800;
      67018: inst = 32'h10a00000;
      67019: inst = 32'hca00004;
      67020: inst = 32'h38632800;
      67021: inst = 32'h38842800;
      67022: inst = 32'h10a00001;
      67023: inst = 32'hca005d3;
      67024: inst = 32'h13e00001;
      67025: inst = 32'hfe0d96a;
      67026: inst = 32'h5be00000;
      67027: inst = 32'h8c50000;
      67028: inst = 32'h24612800;
      67029: inst = 32'h10a0ffff;
      67030: inst = 32'hca0fff7;
      67031: inst = 32'h24822800;
      67032: inst = 32'h10a00000;
      67033: inst = 32'hca00004;
      67034: inst = 32'h38632800;
      67035: inst = 32'h38842800;
      67036: inst = 32'h10a00001;
      67037: inst = 32'hca005e1;
      67038: inst = 32'h13e00001;
      67039: inst = 32'hfe0d96a;
      67040: inst = 32'h5be00000;
      67041: inst = 32'h8c50000;
      67042: inst = 32'h24612800;
      67043: inst = 32'h10a0ffff;
      67044: inst = 32'hca0fff7;
      67045: inst = 32'h24822800;
      67046: inst = 32'h10a00000;
      67047: inst = 32'hca00004;
      67048: inst = 32'h38632800;
      67049: inst = 32'h38842800;
      67050: inst = 32'h10a00001;
      67051: inst = 32'hca005ef;
      67052: inst = 32'h13e00001;
      67053: inst = 32'hfe0d96a;
      67054: inst = 32'h5be00000;
      67055: inst = 32'h8c50000;
      67056: inst = 32'h24612800;
      67057: inst = 32'h10a0ffff;
      67058: inst = 32'hca0fff7;
      67059: inst = 32'h24822800;
      67060: inst = 32'h10a00000;
      67061: inst = 32'hca00004;
      67062: inst = 32'h38632800;
      67063: inst = 32'h38842800;
      67064: inst = 32'h10a00001;
      67065: inst = 32'hca005fd;
      67066: inst = 32'h13e00001;
      67067: inst = 32'hfe0d96a;
      67068: inst = 32'h5be00000;
      67069: inst = 32'h8c50000;
      67070: inst = 32'h24612800;
      67071: inst = 32'h10a0ffff;
      67072: inst = 32'hca0fff7;
      67073: inst = 32'h24822800;
      67074: inst = 32'h10a00000;
      67075: inst = 32'hca00004;
      67076: inst = 32'h38632800;
      67077: inst = 32'h38842800;
      67078: inst = 32'h10a00001;
      67079: inst = 32'hca0060b;
      67080: inst = 32'h13e00001;
      67081: inst = 32'hfe0d96a;
      67082: inst = 32'h5be00000;
      67083: inst = 32'h8c50000;
      67084: inst = 32'h24612800;
      67085: inst = 32'h10a0ffff;
      67086: inst = 32'hca0fff7;
      67087: inst = 32'h24822800;
      67088: inst = 32'h10a00000;
      67089: inst = 32'hca00004;
      67090: inst = 32'h38632800;
      67091: inst = 32'h38842800;
      67092: inst = 32'h10a00001;
      67093: inst = 32'hca00619;
      67094: inst = 32'h13e00001;
      67095: inst = 32'hfe0d96a;
      67096: inst = 32'h5be00000;
      67097: inst = 32'h8c50000;
      67098: inst = 32'h24612800;
      67099: inst = 32'h10a0ffff;
      67100: inst = 32'hca0fff7;
      67101: inst = 32'h24822800;
      67102: inst = 32'h10a00000;
      67103: inst = 32'hca00004;
      67104: inst = 32'h38632800;
      67105: inst = 32'h38842800;
      67106: inst = 32'h10a00001;
      67107: inst = 32'hca00627;
      67108: inst = 32'h13e00001;
      67109: inst = 32'hfe0d96a;
      67110: inst = 32'h5be00000;
      67111: inst = 32'h8c50000;
      67112: inst = 32'h24612800;
      67113: inst = 32'h10a0ffff;
      67114: inst = 32'hca0fff7;
      67115: inst = 32'h24822800;
      67116: inst = 32'h10a00000;
      67117: inst = 32'hca00004;
      67118: inst = 32'h38632800;
      67119: inst = 32'h38842800;
      67120: inst = 32'h10a00001;
      67121: inst = 32'hca00635;
      67122: inst = 32'h13e00001;
      67123: inst = 32'hfe0d96a;
      67124: inst = 32'h5be00000;
      67125: inst = 32'h8c50000;
      67126: inst = 32'h24612800;
      67127: inst = 32'h10a0ffff;
      67128: inst = 32'hca0fff7;
      67129: inst = 32'h24822800;
      67130: inst = 32'h10a00000;
      67131: inst = 32'hca00004;
      67132: inst = 32'h38632800;
      67133: inst = 32'h38842800;
      67134: inst = 32'h10a00001;
      67135: inst = 32'hca00643;
      67136: inst = 32'h13e00001;
      67137: inst = 32'hfe0d96a;
      67138: inst = 32'h5be00000;
      67139: inst = 32'h8c50000;
      67140: inst = 32'h24612800;
      67141: inst = 32'h10a0ffff;
      67142: inst = 32'hca0fff7;
      67143: inst = 32'h24822800;
      67144: inst = 32'h10a00000;
      67145: inst = 32'hca00004;
      67146: inst = 32'h38632800;
      67147: inst = 32'h38842800;
      67148: inst = 32'h10a00001;
      67149: inst = 32'hca00651;
      67150: inst = 32'h13e00001;
      67151: inst = 32'hfe0d96a;
      67152: inst = 32'h5be00000;
      67153: inst = 32'h8c50000;
      67154: inst = 32'h24612800;
      67155: inst = 32'h10a0ffff;
      67156: inst = 32'hca0fff7;
      67157: inst = 32'h24822800;
      67158: inst = 32'h10a00000;
      67159: inst = 32'hca00004;
      67160: inst = 32'h38632800;
      67161: inst = 32'h38842800;
      67162: inst = 32'h10a00001;
      67163: inst = 32'hca0065f;
      67164: inst = 32'h13e00001;
      67165: inst = 32'hfe0d96a;
      67166: inst = 32'h5be00000;
      67167: inst = 32'h8c50000;
      67168: inst = 32'h24612800;
      67169: inst = 32'h10a0ffff;
      67170: inst = 32'hca0fff7;
      67171: inst = 32'h24822800;
      67172: inst = 32'h10a00000;
      67173: inst = 32'hca00004;
      67174: inst = 32'h38632800;
      67175: inst = 32'h38842800;
      67176: inst = 32'h10a00001;
      67177: inst = 32'hca0066d;
      67178: inst = 32'h13e00001;
      67179: inst = 32'hfe0d96a;
      67180: inst = 32'h5be00000;
      67181: inst = 32'h8c50000;
      67182: inst = 32'h24612800;
      67183: inst = 32'h10a0ffff;
      67184: inst = 32'hca0fff7;
      67185: inst = 32'h24822800;
      67186: inst = 32'h10a00000;
      67187: inst = 32'hca00004;
      67188: inst = 32'h38632800;
      67189: inst = 32'h38842800;
      67190: inst = 32'h10a00001;
      67191: inst = 32'hca0067b;
      67192: inst = 32'h13e00001;
      67193: inst = 32'hfe0d96a;
      67194: inst = 32'h5be00000;
      67195: inst = 32'h8c50000;
      67196: inst = 32'h24612800;
      67197: inst = 32'h10a0ffff;
      67198: inst = 32'hca0fff7;
      67199: inst = 32'h24822800;
      67200: inst = 32'h10a00000;
      67201: inst = 32'hca00004;
      67202: inst = 32'h38632800;
      67203: inst = 32'h38842800;
      67204: inst = 32'h10a00001;
      67205: inst = 32'hca00689;
      67206: inst = 32'h13e00001;
      67207: inst = 32'hfe0d96a;
      67208: inst = 32'h5be00000;
      67209: inst = 32'h8c50000;
      67210: inst = 32'h24612800;
      67211: inst = 32'h10a0ffff;
      67212: inst = 32'hca0fff7;
      67213: inst = 32'h24822800;
      67214: inst = 32'h10a00000;
      67215: inst = 32'hca00004;
      67216: inst = 32'h38632800;
      67217: inst = 32'h38842800;
      67218: inst = 32'h10a00001;
      67219: inst = 32'hca00697;
      67220: inst = 32'h13e00001;
      67221: inst = 32'hfe0d96a;
      67222: inst = 32'h5be00000;
      67223: inst = 32'h8c50000;
      67224: inst = 32'h24612800;
      67225: inst = 32'h10a0ffff;
      67226: inst = 32'hca0fff7;
      67227: inst = 32'h24822800;
      67228: inst = 32'h10a00000;
      67229: inst = 32'hca00004;
      67230: inst = 32'h38632800;
      67231: inst = 32'h38842800;
      67232: inst = 32'h10a00001;
      67233: inst = 32'hca006a5;
      67234: inst = 32'h13e00001;
      67235: inst = 32'hfe0d96a;
      67236: inst = 32'h5be00000;
      67237: inst = 32'h8c50000;
      67238: inst = 32'h24612800;
      67239: inst = 32'h10a0ffff;
      67240: inst = 32'hca0fff7;
      67241: inst = 32'h24822800;
      67242: inst = 32'h10a00000;
      67243: inst = 32'hca00004;
      67244: inst = 32'h38632800;
      67245: inst = 32'h38842800;
      67246: inst = 32'h10a00001;
      67247: inst = 32'hca006b3;
      67248: inst = 32'h13e00001;
      67249: inst = 32'hfe0d96a;
      67250: inst = 32'h5be00000;
      67251: inst = 32'h8c50000;
      67252: inst = 32'h24612800;
      67253: inst = 32'h10a0ffff;
      67254: inst = 32'hca0fff7;
      67255: inst = 32'h24822800;
      67256: inst = 32'h10a00000;
      67257: inst = 32'hca00004;
      67258: inst = 32'h38632800;
      67259: inst = 32'h38842800;
      67260: inst = 32'h10a00001;
      67261: inst = 32'hca006c1;
      67262: inst = 32'h13e00001;
      67263: inst = 32'hfe0d96a;
      67264: inst = 32'h5be00000;
      67265: inst = 32'h8c50000;
      67266: inst = 32'h24612800;
      67267: inst = 32'h10a0ffff;
      67268: inst = 32'hca0fff7;
      67269: inst = 32'h24822800;
      67270: inst = 32'h10a00000;
      67271: inst = 32'hca00004;
      67272: inst = 32'h38632800;
      67273: inst = 32'h38842800;
      67274: inst = 32'h10a00001;
      67275: inst = 32'hca006cf;
      67276: inst = 32'h13e00001;
      67277: inst = 32'hfe0d96a;
      67278: inst = 32'h5be00000;
      67279: inst = 32'h8c50000;
      67280: inst = 32'h24612800;
      67281: inst = 32'h10a0ffff;
      67282: inst = 32'hca0fff7;
      67283: inst = 32'h24822800;
      67284: inst = 32'h10a00000;
      67285: inst = 32'hca00004;
      67286: inst = 32'h38632800;
      67287: inst = 32'h38842800;
      67288: inst = 32'h10a00001;
      67289: inst = 32'hca006dd;
      67290: inst = 32'h13e00001;
      67291: inst = 32'hfe0d96a;
      67292: inst = 32'h5be00000;
      67293: inst = 32'h8c50000;
      67294: inst = 32'h24612800;
      67295: inst = 32'h10a0ffff;
      67296: inst = 32'hca0fff7;
      67297: inst = 32'h24822800;
      67298: inst = 32'h10a00000;
      67299: inst = 32'hca00004;
      67300: inst = 32'h38632800;
      67301: inst = 32'h38842800;
      67302: inst = 32'h10a00001;
      67303: inst = 32'hca006eb;
      67304: inst = 32'h13e00001;
      67305: inst = 32'hfe0d96a;
      67306: inst = 32'h5be00000;
      67307: inst = 32'h8c50000;
      67308: inst = 32'h24612800;
      67309: inst = 32'h10a0ffff;
      67310: inst = 32'hca0fff7;
      67311: inst = 32'h24822800;
      67312: inst = 32'h10a00000;
      67313: inst = 32'hca00004;
      67314: inst = 32'h38632800;
      67315: inst = 32'h38842800;
      67316: inst = 32'h10a00001;
      67317: inst = 32'hca006f9;
      67318: inst = 32'h13e00001;
      67319: inst = 32'hfe0d96a;
      67320: inst = 32'h5be00000;
      67321: inst = 32'h8c50000;
      67322: inst = 32'h24612800;
      67323: inst = 32'h10a0ffff;
      67324: inst = 32'hca0fff7;
      67325: inst = 32'h24822800;
      67326: inst = 32'h10a00000;
      67327: inst = 32'hca00004;
      67328: inst = 32'h38632800;
      67329: inst = 32'h38842800;
      67330: inst = 32'h10a00001;
      67331: inst = 32'hca00707;
      67332: inst = 32'h13e00001;
      67333: inst = 32'hfe0d96a;
      67334: inst = 32'h5be00000;
      67335: inst = 32'h8c50000;
      67336: inst = 32'h24612800;
      67337: inst = 32'h10a0ffff;
      67338: inst = 32'hca0fff7;
      67339: inst = 32'h24822800;
      67340: inst = 32'h10a00000;
      67341: inst = 32'hca00004;
      67342: inst = 32'h38632800;
      67343: inst = 32'h38842800;
      67344: inst = 32'h10a00001;
      67345: inst = 32'hca00715;
      67346: inst = 32'h13e00001;
      67347: inst = 32'hfe0d96a;
      67348: inst = 32'h5be00000;
      67349: inst = 32'h8c50000;
      67350: inst = 32'h24612800;
      67351: inst = 32'h10a0ffff;
      67352: inst = 32'hca0fff7;
      67353: inst = 32'h24822800;
      67354: inst = 32'h10a00000;
      67355: inst = 32'hca00004;
      67356: inst = 32'h38632800;
      67357: inst = 32'h38842800;
      67358: inst = 32'h10a00001;
      67359: inst = 32'hca00723;
      67360: inst = 32'h13e00001;
      67361: inst = 32'hfe0d96a;
      67362: inst = 32'h5be00000;
      67363: inst = 32'h8c50000;
      67364: inst = 32'h24612800;
      67365: inst = 32'h10a0ffff;
      67366: inst = 32'hca0fff7;
      67367: inst = 32'h24822800;
      67368: inst = 32'h10a00000;
      67369: inst = 32'hca00004;
      67370: inst = 32'h38632800;
      67371: inst = 32'h38842800;
      67372: inst = 32'h10a00001;
      67373: inst = 32'hca00731;
      67374: inst = 32'h13e00001;
      67375: inst = 32'hfe0d96a;
      67376: inst = 32'h5be00000;
      67377: inst = 32'h8c50000;
      67378: inst = 32'h24612800;
      67379: inst = 32'h10a0ffff;
      67380: inst = 32'hca0fff7;
      67381: inst = 32'h24822800;
      67382: inst = 32'h10a00000;
      67383: inst = 32'hca00004;
      67384: inst = 32'h38632800;
      67385: inst = 32'h38842800;
      67386: inst = 32'h10a00001;
      67387: inst = 32'hca0073f;
      67388: inst = 32'h13e00001;
      67389: inst = 32'hfe0d96a;
      67390: inst = 32'h5be00000;
      67391: inst = 32'h8c50000;
      67392: inst = 32'h24612800;
      67393: inst = 32'h10a0ffff;
      67394: inst = 32'hca0fff7;
      67395: inst = 32'h24822800;
      67396: inst = 32'h10a00000;
      67397: inst = 32'hca00004;
      67398: inst = 32'h38632800;
      67399: inst = 32'h38842800;
      67400: inst = 32'h10a00001;
      67401: inst = 32'hca0074d;
      67402: inst = 32'h13e00001;
      67403: inst = 32'hfe0d96a;
      67404: inst = 32'h5be00000;
      67405: inst = 32'h8c50000;
      67406: inst = 32'h24612800;
      67407: inst = 32'h10a0ffff;
      67408: inst = 32'hca0fff7;
      67409: inst = 32'h24822800;
      67410: inst = 32'h10a00000;
      67411: inst = 32'hca00004;
      67412: inst = 32'h38632800;
      67413: inst = 32'h38842800;
      67414: inst = 32'h10a00001;
      67415: inst = 32'hca0075b;
      67416: inst = 32'h13e00001;
      67417: inst = 32'hfe0d96a;
      67418: inst = 32'h5be00000;
      67419: inst = 32'h8c50000;
      67420: inst = 32'h24612800;
      67421: inst = 32'h10a0ffff;
      67422: inst = 32'hca0fff7;
      67423: inst = 32'h24822800;
      67424: inst = 32'h10a00000;
      67425: inst = 32'hca00004;
      67426: inst = 32'h38632800;
      67427: inst = 32'h38842800;
      67428: inst = 32'h10a00001;
      67429: inst = 32'hca00769;
      67430: inst = 32'h13e00001;
      67431: inst = 32'hfe0d96a;
      67432: inst = 32'h5be00000;
      67433: inst = 32'h8c50000;
      67434: inst = 32'h24612800;
      67435: inst = 32'h10a0ffff;
      67436: inst = 32'hca0fff8;
      67437: inst = 32'h24822800;
      67438: inst = 32'h10a00000;
      67439: inst = 32'hca00004;
      67440: inst = 32'h38632800;
      67441: inst = 32'h38842800;
      67442: inst = 32'h10a00001;
      67443: inst = 32'hca00777;
      67444: inst = 32'h13e00001;
      67445: inst = 32'hfe0d96a;
      67446: inst = 32'h5be00000;
      67447: inst = 32'h8c50000;
      67448: inst = 32'h24612800;
      67449: inst = 32'h10a0ffff;
      67450: inst = 32'hca0fff8;
      67451: inst = 32'h24822800;
      67452: inst = 32'h10a00000;
      67453: inst = 32'hca00004;
      67454: inst = 32'h38632800;
      67455: inst = 32'h38842800;
      67456: inst = 32'h10a00001;
      67457: inst = 32'hca00785;
      67458: inst = 32'h13e00001;
      67459: inst = 32'hfe0d96a;
      67460: inst = 32'h5be00000;
      67461: inst = 32'h8c50000;
      67462: inst = 32'h24612800;
      67463: inst = 32'h10a0ffff;
      67464: inst = 32'hca0fff8;
      67465: inst = 32'h24822800;
      67466: inst = 32'h10a00000;
      67467: inst = 32'hca00004;
      67468: inst = 32'h38632800;
      67469: inst = 32'h38842800;
      67470: inst = 32'h10a00001;
      67471: inst = 32'hca00793;
      67472: inst = 32'h13e00001;
      67473: inst = 32'hfe0d96a;
      67474: inst = 32'h5be00000;
      67475: inst = 32'h8c50000;
      67476: inst = 32'h24612800;
      67477: inst = 32'h10a0ffff;
      67478: inst = 32'hca0fff8;
      67479: inst = 32'h24822800;
      67480: inst = 32'h10a00000;
      67481: inst = 32'hca00004;
      67482: inst = 32'h38632800;
      67483: inst = 32'h38842800;
      67484: inst = 32'h10a00001;
      67485: inst = 32'hca007a1;
      67486: inst = 32'h13e00001;
      67487: inst = 32'hfe0d96a;
      67488: inst = 32'h5be00000;
      67489: inst = 32'h8c50000;
      67490: inst = 32'h24612800;
      67491: inst = 32'h10a0ffff;
      67492: inst = 32'hca0fff8;
      67493: inst = 32'h24822800;
      67494: inst = 32'h10a00000;
      67495: inst = 32'hca00004;
      67496: inst = 32'h38632800;
      67497: inst = 32'h38842800;
      67498: inst = 32'h10a00001;
      67499: inst = 32'hca007af;
      67500: inst = 32'h13e00001;
      67501: inst = 32'hfe0d96a;
      67502: inst = 32'h5be00000;
      67503: inst = 32'h8c50000;
      67504: inst = 32'h24612800;
      67505: inst = 32'h10a0ffff;
      67506: inst = 32'hca0fff8;
      67507: inst = 32'h24822800;
      67508: inst = 32'h10a00000;
      67509: inst = 32'hca00004;
      67510: inst = 32'h38632800;
      67511: inst = 32'h38842800;
      67512: inst = 32'h10a00001;
      67513: inst = 32'hca007bd;
      67514: inst = 32'h13e00001;
      67515: inst = 32'hfe0d96a;
      67516: inst = 32'h5be00000;
      67517: inst = 32'h8c50000;
      67518: inst = 32'h24612800;
      67519: inst = 32'h10a0ffff;
      67520: inst = 32'hca0fff8;
      67521: inst = 32'h24822800;
      67522: inst = 32'h10a00000;
      67523: inst = 32'hca00004;
      67524: inst = 32'h38632800;
      67525: inst = 32'h38842800;
      67526: inst = 32'h10a00001;
      67527: inst = 32'hca007cb;
      67528: inst = 32'h13e00001;
      67529: inst = 32'hfe0d96a;
      67530: inst = 32'h5be00000;
      67531: inst = 32'h8c50000;
      67532: inst = 32'h24612800;
      67533: inst = 32'h10a0ffff;
      67534: inst = 32'hca0fff8;
      67535: inst = 32'h24822800;
      67536: inst = 32'h10a00000;
      67537: inst = 32'hca00004;
      67538: inst = 32'h38632800;
      67539: inst = 32'h38842800;
      67540: inst = 32'h10a00001;
      67541: inst = 32'hca007d9;
      67542: inst = 32'h13e00001;
      67543: inst = 32'hfe0d96a;
      67544: inst = 32'h5be00000;
      67545: inst = 32'h8c50000;
      67546: inst = 32'h24612800;
      67547: inst = 32'h10a0ffff;
      67548: inst = 32'hca0fff8;
      67549: inst = 32'h24822800;
      67550: inst = 32'h10a00000;
      67551: inst = 32'hca00004;
      67552: inst = 32'h38632800;
      67553: inst = 32'h38842800;
      67554: inst = 32'h10a00001;
      67555: inst = 32'hca007e7;
      67556: inst = 32'h13e00001;
      67557: inst = 32'hfe0d96a;
      67558: inst = 32'h5be00000;
      67559: inst = 32'h8c50000;
      67560: inst = 32'h24612800;
      67561: inst = 32'h10a0ffff;
      67562: inst = 32'hca0fff8;
      67563: inst = 32'h24822800;
      67564: inst = 32'h10a00000;
      67565: inst = 32'hca00004;
      67566: inst = 32'h38632800;
      67567: inst = 32'h38842800;
      67568: inst = 32'h10a00001;
      67569: inst = 32'hca007f5;
      67570: inst = 32'h13e00001;
      67571: inst = 32'hfe0d96a;
      67572: inst = 32'h5be00000;
      67573: inst = 32'h8c50000;
      67574: inst = 32'h24612800;
      67575: inst = 32'h10a0ffff;
      67576: inst = 32'hca0fff8;
      67577: inst = 32'h24822800;
      67578: inst = 32'h10a00000;
      67579: inst = 32'hca00004;
      67580: inst = 32'h38632800;
      67581: inst = 32'h38842800;
      67582: inst = 32'h10a00001;
      67583: inst = 32'hca00803;
      67584: inst = 32'h13e00001;
      67585: inst = 32'hfe0d96a;
      67586: inst = 32'h5be00000;
      67587: inst = 32'h8c50000;
      67588: inst = 32'h24612800;
      67589: inst = 32'h10a0ffff;
      67590: inst = 32'hca0fff8;
      67591: inst = 32'h24822800;
      67592: inst = 32'h10a00000;
      67593: inst = 32'hca00004;
      67594: inst = 32'h38632800;
      67595: inst = 32'h38842800;
      67596: inst = 32'h10a00001;
      67597: inst = 32'hca00811;
      67598: inst = 32'h13e00001;
      67599: inst = 32'hfe0d96a;
      67600: inst = 32'h5be00000;
      67601: inst = 32'h8c50000;
      67602: inst = 32'h24612800;
      67603: inst = 32'h10a0ffff;
      67604: inst = 32'hca0fff8;
      67605: inst = 32'h24822800;
      67606: inst = 32'h10a00000;
      67607: inst = 32'hca00004;
      67608: inst = 32'h38632800;
      67609: inst = 32'h38842800;
      67610: inst = 32'h10a00001;
      67611: inst = 32'hca0081f;
      67612: inst = 32'h13e00001;
      67613: inst = 32'hfe0d96a;
      67614: inst = 32'h5be00000;
      67615: inst = 32'h8c50000;
      67616: inst = 32'h24612800;
      67617: inst = 32'h10a0ffff;
      67618: inst = 32'hca0fff8;
      67619: inst = 32'h24822800;
      67620: inst = 32'h10a00000;
      67621: inst = 32'hca00004;
      67622: inst = 32'h38632800;
      67623: inst = 32'h38842800;
      67624: inst = 32'h10a00001;
      67625: inst = 32'hca0082d;
      67626: inst = 32'h13e00001;
      67627: inst = 32'hfe0d96a;
      67628: inst = 32'h5be00000;
      67629: inst = 32'h8c50000;
      67630: inst = 32'h24612800;
      67631: inst = 32'h10a0ffff;
      67632: inst = 32'hca0fff8;
      67633: inst = 32'h24822800;
      67634: inst = 32'h10a00000;
      67635: inst = 32'hca00004;
      67636: inst = 32'h38632800;
      67637: inst = 32'h38842800;
      67638: inst = 32'h10a00001;
      67639: inst = 32'hca0083b;
      67640: inst = 32'h13e00001;
      67641: inst = 32'hfe0d96a;
      67642: inst = 32'h5be00000;
      67643: inst = 32'h8c50000;
      67644: inst = 32'h24612800;
      67645: inst = 32'h10a0ffff;
      67646: inst = 32'hca0fff8;
      67647: inst = 32'h24822800;
      67648: inst = 32'h10a00000;
      67649: inst = 32'hca00004;
      67650: inst = 32'h38632800;
      67651: inst = 32'h38842800;
      67652: inst = 32'h10a00001;
      67653: inst = 32'hca00849;
      67654: inst = 32'h13e00001;
      67655: inst = 32'hfe0d96a;
      67656: inst = 32'h5be00000;
      67657: inst = 32'h8c50000;
      67658: inst = 32'h24612800;
      67659: inst = 32'h10a0ffff;
      67660: inst = 32'hca0fff8;
      67661: inst = 32'h24822800;
      67662: inst = 32'h10a00000;
      67663: inst = 32'hca00004;
      67664: inst = 32'h38632800;
      67665: inst = 32'h38842800;
      67666: inst = 32'h10a00001;
      67667: inst = 32'hca00857;
      67668: inst = 32'h13e00001;
      67669: inst = 32'hfe0d96a;
      67670: inst = 32'h5be00000;
      67671: inst = 32'h8c50000;
      67672: inst = 32'h24612800;
      67673: inst = 32'h10a0ffff;
      67674: inst = 32'hca0fff8;
      67675: inst = 32'h24822800;
      67676: inst = 32'h10a00000;
      67677: inst = 32'hca00004;
      67678: inst = 32'h38632800;
      67679: inst = 32'h38842800;
      67680: inst = 32'h10a00001;
      67681: inst = 32'hca00865;
      67682: inst = 32'h13e00001;
      67683: inst = 32'hfe0d96a;
      67684: inst = 32'h5be00000;
      67685: inst = 32'h8c50000;
      67686: inst = 32'h24612800;
      67687: inst = 32'h10a0ffff;
      67688: inst = 32'hca0fff8;
      67689: inst = 32'h24822800;
      67690: inst = 32'h10a00000;
      67691: inst = 32'hca00004;
      67692: inst = 32'h38632800;
      67693: inst = 32'h38842800;
      67694: inst = 32'h10a00001;
      67695: inst = 32'hca00873;
      67696: inst = 32'h13e00001;
      67697: inst = 32'hfe0d96a;
      67698: inst = 32'h5be00000;
      67699: inst = 32'h8c50000;
      67700: inst = 32'h24612800;
      67701: inst = 32'h10a0ffff;
      67702: inst = 32'hca0fff8;
      67703: inst = 32'h24822800;
      67704: inst = 32'h10a00000;
      67705: inst = 32'hca00004;
      67706: inst = 32'h38632800;
      67707: inst = 32'h38842800;
      67708: inst = 32'h10a00001;
      67709: inst = 32'hca00881;
      67710: inst = 32'h13e00001;
      67711: inst = 32'hfe0d96a;
      67712: inst = 32'h5be00000;
      67713: inst = 32'h8c50000;
      67714: inst = 32'h24612800;
      67715: inst = 32'h10a0ffff;
      67716: inst = 32'hca0fff8;
      67717: inst = 32'h24822800;
      67718: inst = 32'h10a00000;
      67719: inst = 32'hca00004;
      67720: inst = 32'h38632800;
      67721: inst = 32'h38842800;
      67722: inst = 32'h10a00001;
      67723: inst = 32'hca0088f;
      67724: inst = 32'h13e00001;
      67725: inst = 32'hfe0d96a;
      67726: inst = 32'h5be00000;
      67727: inst = 32'h8c50000;
      67728: inst = 32'h24612800;
      67729: inst = 32'h10a0ffff;
      67730: inst = 32'hca0fff8;
      67731: inst = 32'h24822800;
      67732: inst = 32'h10a00000;
      67733: inst = 32'hca00004;
      67734: inst = 32'h38632800;
      67735: inst = 32'h38842800;
      67736: inst = 32'h10a00001;
      67737: inst = 32'hca0089d;
      67738: inst = 32'h13e00001;
      67739: inst = 32'hfe0d96a;
      67740: inst = 32'h5be00000;
      67741: inst = 32'h8c50000;
      67742: inst = 32'h24612800;
      67743: inst = 32'h10a0ffff;
      67744: inst = 32'hca0fff8;
      67745: inst = 32'h24822800;
      67746: inst = 32'h10a00000;
      67747: inst = 32'hca00004;
      67748: inst = 32'h38632800;
      67749: inst = 32'h38842800;
      67750: inst = 32'h10a00001;
      67751: inst = 32'hca008ab;
      67752: inst = 32'h13e00001;
      67753: inst = 32'hfe0d96a;
      67754: inst = 32'h5be00000;
      67755: inst = 32'h8c50000;
      67756: inst = 32'h24612800;
      67757: inst = 32'h10a0ffff;
      67758: inst = 32'hca0fff8;
      67759: inst = 32'h24822800;
      67760: inst = 32'h10a00000;
      67761: inst = 32'hca00004;
      67762: inst = 32'h38632800;
      67763: inst = 32'h38842800;
      67764: inst = 32'h10a00001;
      67765: inst = 32'hca008b9;
      67766: inst = 32'h13e00001;
      67767: inst = 32'hfe0d96a;
      67768: inst = 32'h5be00000;
      67769: inst = 32'h8c50000;
      67770: inst = 32'h24612800;
      67771: inst = 32'h10a0ffff;
      67772: inst = 32'hca0fff8;
      67773: inst = 32'h24822800;
      67774: inst = 32'h10a00000;
      67775: inst = 32'hca00004;
      67776: inst = 32'h38632800;
      67777: inst = 32'h38842800;
      67778: inst = 32'h10a00001;
      67779: inst = 32'hca008c7;
      67780: inst = 32'h13e00001;
      67781: inst = 32'hfe0d96a;
      67782: inst = 32'h5be00000;
      67783: inst = 32'h8c50000;
      67784: inst = 32'h24612800;
      67785: inst = 32'h10a0ffff;
      67786: inst = 32'hca0fff8;
      67787: inst = 32'h24822800;
      67788: inst = 32'h10a00000;
      67789: inst = 32'hca00004;
      67790: inst = 32'h38632800;
      67791: inst = 32'h38842800;
      67792: inst = 32'h10a00001;
      67793: inst = 32'hca008d5;
      67794: inst = 32'h13e00001;
      67795: inst = 32'hfe0d96a;
      67796: inst = 32'h5be00000;
      67797: inst = 32'h8c50000;
      67798: inst = 32'h24612800;
      67799: inst = 32'h10a0ffff;
      67800: inst = 32'hca0fff8;
      67801: inst = 32'h24822800;
      67802: inst = 32'h10a00000;
      67803: inst = 32'hca00004;
      67804: inst = 32'h38632800;
      67805: inst = 32'h38842800;
      67806: inst = 32'h10a00001;
      67807: inst = 32'hca008e3;
      67808: inst = 32'h13e00001;
      67809: inst = 32'hfe0d96a;
      67810: inst = 32'h5be00000;
      67811: inst = 32'h8c50000;
      67812: inst = 32'h24612800;
      67813: inst = 32'h10a0ffff;
      67814: inst = 32'hca0fff8;
      67815: inst = 32'h24822800;
      67816: inst = 32'h10a00000;
      67817: inst = 32'hca00004;
      67818: inst = 32'h38632800;
      67819: inst = 32'h38842800;
      67820: inst = 32'h10a00001;
      67821: inst = 32'hca008f1;
      67822: inst = 32'h13e00001;
      67823: inst = 32'hfe0d96a;
      67824: inst = 32'h5be00000;
      67825: inst = 32'h8c50000;
      67826: inst = 32'h24612800;
      67827: inst = 32'h10a0ffff;
      67828: inst = 32'hca0fff8;
      67829: inst = 32'h24822800;
      67830: inst = 32'h10a00000;
      67831: inst = 32'hca00004;
      67832: inst = 32'h38632800;
      67833: inst = 32'h38842800;
      67834: inst = 32'h10a00001;
      67835: inst = 32'hca008ff;
      67836: inst = 32'h13e00001;
      67837: inst = 32'hfe0d96a;
      67838: inst = 32'h5be00000;
      67839: inst = 32'h8c50000;
      67840: inst = 32'h24612800;
      67841: inst = 32'h10a0ffff;
      67842: inst = 32'hca0fff8;
      67843: inst = 32'h24822800;
      67844: inst = 32'h10a00000;
      67845: inst = 32'hca00004;
      67846: inst = 32'h38632800;
      67847: inst = 32'h38842800;
      67848: inst = 32'h10a00001;
      67849: inst = 32'hca0090d;
      67850: inst = 32'h13e00001;
      67851: inst = 32'hfe0d96a;
      67852: inst = 32'h5be00000;
      67853: inst = 32'h8c50000;
      67854: inst = 32'h24612800;
      67855: inst = 32'h10a0ffff;
      67856: inst = 32'hca0fff8;
      67857: inst = 32'h24822800;
      67858: inst = 32'h10a00000;
      67859: inst = 32'hca00004;
      67860: inst = 32'h38632800;
      67861: inst = 32'h38842800;
      67862: inst = 32'h10a00001;
      67863: inst = 32'hca0091b;
      67864: inst = 32'h13e00001;
      67865: inst = 32'hfe0d96a;
      67866: inst = 32'h5be00000;
      67867: inst = 32'h8c50000;
      67868: inst = 32'h24612800;
      67869: inst = 32'h10a0ffff;
      67870: inst = 32'hca0fff8;
      67871: inst = 32'h24822800;
      67872: inst = 32'h10a00000;
      67873: inst = 32'hca00004;
      67874: inst = 32'h38632800;
      67875: inst = 32'h38842800;
      67876: inst = 32'h10a00001;
      67877: inst = 32'hca00929;
      67878: inst = 32'h13e00001;
      67879: inst = 32'hfe0d96a;
      67880: inst = 32'h5be00000;
      67881: inst = 32'h8c50000;
      67882: inst = 32'h24612800;
      67883: inst = 32'h10a0ffff;
      67884: inst = 32'hca0fff8;
      67885: inst = 32'h24822800;
      67886: inst = 32'h10a00000;
      67887: inst = 32'hca00004;
      67888: inst = 32'h38632800;
      67889: inst = 32'h38842800;
      67890: inst = 32'h10a00001;
      67891: inst = 32'hca00937;
      67892: inst = 32'h13e00001;
      67893: inst = 32'hfe0d96a;
      67894: inst = 32'h5be00000;
      67895: inst = 32'h8c50000;
      67896: inst = 32'h24612800;
      67897: inst = 32'h10a0ffff;
      67898: inst = 32'hca0fff8;
      67899: inst = 32'h24822800;
      67900: inst = 32'h10a00000;
      67901: inst = 32'hca00004;
      67902: inst = 32'h38632800;
      67903: inst = 32'h38842800;
      67904: inst = 32'h10a00001;
      67905: inst = 32'hca00945;
      67906: inst = 32'h13e00001;
      67907: inst = 32'hfe0d96a;
      67908: inst = 32'h5be00000;
      67909: inst = 32'h8c50000;
      67910: inst = 32'h24612800;
      67911: inst = 32'h10a0ffff;
      67912: inst = 32'hca0fff8;
      67913: inst = 32'h24822800;
      67914: inst = 32'h10a00000;
      67915: inst = 32'hca00004;
      67916: inst = 32'h38632800;
      67917: inst = 32'h38842800;
      67918: inst = 32'h10a00001;
      67919: inst = 32'hca00953;
      67920: inst = 32'h13e00001;
      67921: inst = 32'hfe0d96a;
      67922: inst = 32'h5be00000;
      67923: inst = 32'h8c50000;
      67924: inst = 32'h24612800;
      67925: inst = 32'h10a0ffff;
      67926: inst = 32'hca0fff8;
      67927: inst = 32'h24822800;
      67928: inst = 32'h10a00000;
      67929: inst = 32'hca00004;
      67930: inst = 32'h38632800;
      67931: inst = 32'h38842800;
      67932: inst = 32'h10a00001;
      67933: inst = 32'hca00961;
      67934: inst = 32'h13e00001;
      67935: inst = 32'hfe0d96a;
      67936: inst = 32'h5be00000;
      67937: inst = 32'h8c50000;
      67938: inst = 32'h24612800;
      67939: inst = 32'h10a0ffff;
      67940: inst = 32'hca0fff8;
      67941: inst = 32'h24822800;
      67942: inst = 32'h10a00000;
      67943: inst = 32'hca00004;
      67944: inst = 32'h38632800;
      67945: inst = 32'h38842800;
      67946: inst = 32'h10a00001;
      67947: inst = 32'hca0096f;
      67948: inst = 32'h13e00001;
      67949: inst = 32'hfe0d96a;
      67950: inst = 32'h5be00000;
      67951: inst = 32'h8c50000;
      67952: inst = 32'h24612800;
      67953: inst = 32'h10a0ffff;
      67954: inst = 32'hca0fff8;
      67955: inst = 32'h24822800;
      67956: inst = 32'h10a00000;
      67957: inst = 32'hca00004;
      67958: inst = 32'h38632800;
      67959: inst = 32'h38842800;
      67960: inst = 32'h10a00001;
      67961: inst = 32'hca0097d;
      67962: inst = 32'h13e00001;
      67963: inst = 32'hfe0d96a;
      67964: inst = 32'h5be00000;
      67965: inst = 32'h8c50000;
      67966: inst = 32'h24612800;
      67967: inst = 32'h10a0ffff;
      67968: inst = 32'hca0fff8;
      67969: inst = 32'h24822800;
      67970: inst = 32'h10a00000;
      67971: inst = 32'hca00004;
      67972: inst = 32'h38632800;
      67973: inst = 32'h38842800;
      67974: inst = 32'h10a00001;
      67975: inst = 32'hca0098b;
      67976: inst = 32'h13e00001;
      67977: inst = 32'hfe0d96a;
      67978: inst = 32'h5be00000;
      67979: inst = 32'h8c50000;
      67980: inst = 32'h24612800;
      67981: inst = 32'h10a0ffff;
      67982: inst = 32'hca0fff8;
      67983: inst = 32'h24822800;
      67984: inst = 32'h10a00000;
      67985: inst = 32'hca00004;
      67986: inst = 32'h38632800;
      67987: inst = 32'h38842800;
      67988: inst = 32'h10a00001;
      67989: inst = 32'hca00999;
      67990: inst = 32'h13e00001;
      67991: inst = 32'hfe0d96a;
      67992: inst = 32'h5be00000;
      67993: inst = 32'h8c50000;
      67994: inst = 32'h24612800;
      67995: inst = 32'h10a0ffff;
      67996: inst = 32'hca0fff8;
      67997: inst = 32'h24822800;
      67998: inst = 32'h10a00000;
      67999: inst = 32'hca00004;
      68000: inst = 32'h38632800;
      68001: inst = 32'h38842800;
      68002: inst = 32'h10a00001;
      68003: inst = 32'hca009a7;
      68004: inst = 32'h13e00001;
      68005: inst = 32'hfe0d96a;
      68006: inst = 32'h5be00000;
      68007: inst = 32'h8c50000;
      68008: inst = 32'h24612800;
      68009: inst = 32'h10a0ffff;
      68010: inst = 32'hca0fff8;
      68011: inst = 32'h24822800;
      68012: inst = 32'h10a00000;
      68013: inst = 32'hca00004;
      68014: inst = 32'h38632800;
      68015: inst = 32'h38842800;
      68016: inst = 32'h10a00001;
      68017: inst = 32'hca009b5;
      68018: inst = 32'h13e00001;
      68019: inst = 32'hfe0d96a;
      68020: inst = 32'h5be00000;
      68021: inst = 32'h8c50000;
      68022: inst = 32'h24612800;
      68023: inst = 32'h10a0ffff;
      68024: inst = 32'hca0fff8;
      68025: inst = 32'h24822800;
      68026: inst = 32'h10a00000;
      68027: inst = 32'hca00004;
      68028: inst = 32'h38632800;
      68029: inst = 32'h38842800;
      68030: inst = 32'h10a00001;
      68031: inst = 32'hca009c3;
      68032: inst = 32'h13e00001;
      68033: inst = 32'hfe0d96a;
      68034: inst = 32'h5be00000;
      68035: inst = 32'h8c50000;
      68036: inst = 32'h24612800;
      68037: inst = 32'h10a0ffff;
      68038: inst = 32'hca0fff8;
      68039: inst = 32'h24822800;
      68040: inst = 32'h10a00000;
      68041: inst = 32'hca00004;
      68042: inst = 32'h38632800;
      68043: inst = 32'h38842800;
      68044: inst = 32'h10a00001;
      68045: inst = 32'hca009d1;
      68046: inst = 32'h13e00001;
      68047: inst = 32'hfe0d96a;
      68048: inst = 32'h5be00000;
      68049: inst = 32'h8c50000;
      68050: inst = 32'h24612800;
      68051: inst = 32'h10a0ffff;
      68052: inst = 32'hca0fff8;
      68053: inst = 32'h24822800;
      68054: inst = 32'h10a00000;
      68055: inst = 32'hca00004;
      68056: inst = 32'h38632800;
      68057: inst = 32'h38842800;
      68058: inst = 32'h10a00001;
      68059: inst = 32'hca009df;
      68060: inst = 32'h13e00001;
      68061: inst = 32'hfe0d96a;
      68062: inst = 32'h5be00000;
      68063: inst = 32'h8c50000;
      68064: inst = 32'h24612800;
      68065: inst = 32'h10a0ffff;
      68066: inst = 32'hca0fff8;
      68067: inst = 32'h24822800;
      68068: inst = 32'h10a00000;
      68069: inst = 32'hca00004;
      68070: inst = 32'h38632800;
      68071: inst = 32'h38842800;
      68072: inst = 32'h10a00001;
      68073: inst = 32'hca009ed;
      68074: inst = 32'h13e00001;
      68075: inst = 32'hfe0d96a;
      68076: inst = 32'h5be00000;
      68077: inst = 32'h8c50000;
      68078: inst = 32'h24612800;
      68079: inst = 32'h10a0ffff;
      68080: inst = 32'hca0fff8;
      68081: inst = 32'h24822800;
      68082: inst = 32'h10a00000;
      68083: inst = 32'hca00004;
      68084: inst = 32'h38632800;
      68085: inst = 32'h38842800;
      68086: inst = 32'h10a00001;
      68087: inst = 32'hca009fb;
      68088: inst = 32'h13e00001;
      68089: inst = 32'hfe0d96a;
      68090: inst = 32'h5be00000;
      68091: inst = 32'h8c50000;
      68092: inst = 32'h24612800;
      68093: inst = 32'h10a0ffff;
      68094: inst = 32'hca0fff8;
      68095: inst = 32'h24822800;
      68096: inst = 32'h10a00000;
      68097: inst = 32'hca00004;
      68098: inst = 32'h38632800;
      68099: inst = 32'h38842800;
      68100: inst = 32'h10a00001;
      68101: inst = 32'hca00a09;
      68102: inst = 32'h13e00001;
      68103: inst = 32'hfe0d96a;
      68104: inst = 32'h5be00000;
      68105: inst = 32'h8c50000;
      68106: inst = 32'h24612800;
      68107: inst = 32'h10a0ffff;
      68108: inst = 32'hca0fff8;
      68109: inst = 32'h24822800;
      68110: inst = 32'h10a00000;
      68111: inst = 32'hca00004;
      68112: inst = 32'h38632800;
      68113: inst = 32'h38842800;
      68114: inst = 32'h10a00001;
      68115: inst = 32'hca00a17;
      68116: inst = 32'h13e00001;
      68117: inst = 32'hfe0d96a;
      68118: inst = 32'h5be00000;
      68119: inst = 32'h8c50000;
      68120: inst = 32'h24612800;
      68121: inst = 32'h10a0ffff;
      68122: inst = 32'hca0fff8;
      68123: inst = 32'h24822800;
      68124: inst = 32'h10a00000;
      68125: inst = 32'hca00004;
      68126: inst = 32'h38632800;
      68127: inst = 32'h38842800;
      68128: inst = 32'h10a00001;
      68129: inst = 32'hca00a25;
      68130: inst = 32'h13e00001;
      68131: inst = 32'hfe0d96a;
      68132: inst = 32'h5be00000;
      68133: inst = 32'h8c50000;
      68134: inst = 32'h24612800;
      68135: inst = 32'h10a0ffff;
      68136: inst = 32'hca0fff8;
      68137: inst = 32'h24822800;
      68138: inst = 32'h10a00000;
      68139: inst = 32'hca00004;
      68140: inst = 32'h38632800;
      68141: inst = 32'h38842800;
      68142: inst = 32'h10a00001;
      68143: inst = 32'hca00a33;
      68144: inst = 32'h13e00001;
      68145: inst = 32'hfe0d96a;
      68146: inst = 32'h5be00000;
      68147: inst = 32'h8c50000;
      68148: inst = 32'h24612800;
      68149: inst = 32'h10a0ffff;
      68150: inst = 32'hca0fff8;
      68151: inst = 32'h24822800;
      68152: inst = 32'h10a00000;
      68153: inst = 32'hca00004;
      68154: inst = 32'h38632800;
      68155: inst = 32'h38842800;
      68156: inst = 32'h10a00001;
      68157: inst = 32'hca00a41;
      68158: inst = 32'h13e00001;
      68159: inst = 32'hfe0d96a;
      68160: inst = 32'h5be00000;
      68161: inst = 32'h8c50000;
      68162: inst = 32'h24612800;
      68163: inst = 32'h10a0ffff;
      68164: inst = 32'hca0fff8;
      68165: inst = 32'h24822800;
      68166: inst = 32'h10a00000;
      68167: inst = 32'hca00004;
      68168: inst = 32'h38632800;
      68169: inst = 32'h38842800;
      68170: inst = 32'h10a00001;
      68171: inst = 32'hca00a4f;
      68172: inst = 32'h13e00001;
      68173: inst = 32'hfe0d96a;
      68174: inst = 32'h5be00000;
      68175: inst = 32'h8c50000;
      68176: inst = 32'h24612800;
      68177: inst = 32'h10a0ffff;
      68178: inst = 32'hca0fff8;
      68179: inst = 32'h24822800;
      68180: inst = 32'h10a00000;
      68181: inst = 32'hca00004;
      68182: inst = 32'h38632800;
      68183: inst = 32'h38842800;
      68184: inst = 32'h10a00001;
      68185: inst = 32'hca00a5d;
      68186: inst = 32'h13e00001;
      68187: inst = 32'hfe0d96a;
      68188: inst = 32'h5be00000;
      68189: inst = 32'h8c50000;
      68190: inst = 32'h24612800;
      68191: inst = 32'h10a0ffff;
      68192: inst = 32'hca0fff8;
      68193: inst = 32'h24822800;
      68194: inst = 32'h10a00000;
      68195: inst = 32'hca00004;
      68196: inst = 32'h38632800;
      68197: inst = 32'h38842800;
      68198: inst = 32'h10a00001;
      68199: inst = 32'hca00a6b;
      68200: inst = 32'h13e00001;
      68201: inst = 32'hfe0d96a;
      68202: inst = 32'h5be00000;
      68203: inst = 32'h8c50000;
      68204: inst = 32'h24612800;
      68205: inst = 32'h10a0ffff;
      68206: inst = 32'hca0fff8;
      68207: inst = 32'h24822800;
      68208: inst = 32'h10a00000;
      68209: inst = 32'hca00004;
      68210: inst = 32'h38632800;
      68211: inst = 32'h38842800;
      68212: inst = 32'h10a00001;
      68213: inst = 32'hca00a79;
      68214: inst = 32'h13e00001;
      68215: inst = 32'hfe0d96a;
      68216: inst = 32'h5be00000;
      68217: inst = 32'h8c50000;
      68218: inst = 32'h24612800;
      68219: inst = 32'h10a0ffff;
      68220: inst = 32'hca0fff8;
      68221: inst = 32'h24822800;
      68222: inst = 32'h10a00000;
      68223: inst = 32'hca00004;
      68224: inst = 32'h38632800;
      68225: inst = 32'h38842800;
      68226: inst = 32'h10a00001;
      68227: inst = 32'hca00a87;
      68228: inst = 32'h13e00001;
      68229: inst = 32'hfe0d96a;
      68230: inst = 32'h5be00000;
      68231: inst = 32'h8c50000;
      68232: inst = 32'h24612800;
      68233: inst = 32'h10a0ffff;
      68234: inst = 32'hca0fff8;
      68235: inst = 32'h24822800;
      68236: inst = 32'h10a00000;
      68237: inst = 32'hca00004;
      68238: inst = 32'h38632800;
      68239: inst = 32'h38842800;
      68240: inst = 32'h10a00001;
      68241: inst = 32'hca00a95;
      68242: inst = 32'h13e00001;
      68243: inst = 32'hfe0d96a;
      68244: inst = 32'h5be00000;
      68245: inst = 32'h8c50000;
      68246: inst = 32'h24612800;
      68247: inst = 32'h10a0ffff;
      68248: inst = 32'hca0fff8;
      68249: inst = 32'h24822800;
      68250: inst = 32'h10a00000;
      68251: inst = 32'hca00004;
      68252: inst = 32'h38632800;
      68253: inst = 32'h38842800;
      68254: inst = 32'h10a00001;
      68255: inst = 32'hca00aa3;
      68256: inst = 32'h13e00001;
      68257: inst = 32'hfe0d96a;
      68258: inst = 32'h5be00000;
      68259: inst = 32'h8c50000;
      68260: inst = 32'h24612800;
      68261: inst = 32'h10a0ffff;
      68262: inst = 32'hca0fff8;
      68263: inst = 32'h24822800;
      68264: inst = 32'h10a00000;
      68265: inst = 32'hca00004;
      68266: inst = 32'h38632800;
      68267: inst = 32'h38842800;
      68268: inst = 32'h10a00001;
      68269: inst = 32'hca00ab1;
      68270: inst = 32'h13e00001;
      68271: inst = 32'hfe0d96a;
      68272: inst = 32'h5be00000;
      68273: inst = 32'h8c50000;
      68274: inst = 32'h24612800;
      68275: inst = 32'h10a0ffff;
      68276: inst = 32'hca0fff8;
      68277: inst = 32'h24822800;
      68278: inst = 32'h10a00000;
      68279: inst = 32'hca00004;
      68280: inst = 32'h38632800;
      68281: inst = 32'h38842800;
      68282: inst = 32'h10a00001;
      68283: inst = 32'hca00abf;
      68284: inst = 32'h13e00001;
      68285: inst = 32'hfe0d96a;
      68286: inst = 32'h5be00000;
      68287: inst = 32'h8c50000;
      68288: inst = 32'h24612800;
      68289: inst = 32'h10a0ffff;
      68290: inst = 32'hca0fff8;
      68291: inst = 32'h24822800;
      68292: inst = 32'h10a00000;
      68293: inst = 32'hca00004;
      68294: inst = 32'h38632800;
      68295: inst = 32'h38842800;
      68296: inst = 32'h10a00001;
      68297: inst = 32'hca00acd;
      68298: inst = 32'h13e00001;
      68299: inst = 32'hfe0d96a;
      68300: inst = 32'h5be00000;
      68301: inst = 32'h8c50000;
      68302: inst = 32'h24612800;
      68303: inst = 32'h10a0ffff;
      68304: inst = 32'hca0fff8;
      68305: inst = 32'h24822800;
      68306: inst = 32'h10a00000;
      68307: inst = 32'hca00004;
      68308: inst = 32'h38632800;
      68309: inst = 32'h38842800;
      68310: inst = 32'h10a00001;
      68311: inst = 32'hca00adb;
      68312: inst = 32'h13e00001;
      68313: inst = 32'hfe0d96a;
      68314: inst = 32'h5be00000;
      68315: inst = 32'h8c50000;
      68316: inst = 32'h24612800;
      68317: inst = 32'h10a0ffff;
      68318: inst = 32'hca0fff8;
      68319: inst = 32'h24822800;
      68320: inst = 32'h10a00000;
      68321: inst = 32'hca00004;
      68322: inst = 32'h38632800;
      68323: inst = 32'h38842800;
      68324: inst = 32'h10a00001;
      68325: inst = 32'hca00ae9;
      68326: inst = 32'h13e00001;
      68327: inst = 32'hfe0d96a;
      68328: inst = 32'h5be00000;
      68329: inst = 32'h8c50000;
      68330: inst = 32'h24612800;
      68331: inst = 32'h10a0ffff;
      68332: inst = 32'hca0fff8;
      68333: inst = 32'h24822800;
      68334: inst = 32'h10a00000;
      68335: inst = 32'hca00004;
      68336: inst = 32'h38632800;
      68337: inst = 32'h38842800;
      68338: inst = 32'h10a00001;
      68339: inst = 32'hca00af7;
      68340: inst = 32'h13e00001;
      68341: inst = 32'hfe0d96a;
      68342: inst = 32'h5be00000;
      68343: inst = 32'h8c50000;
      68344: inst = 32'h24612800;
      68345: inst = 32'h10a0ffff;
      68346: inst = 32'hca0fff8;
      68347: inst = 32'h24822800;
      68348: inst = 32'h10a00000;
      68349: inst = 32'hca00004;
      68350: inst = 32'h38632800;
      68351: inst = 32'h38842800;
      68352: inst = 32'h10a00001;
      68353: inst = 32'hca00b05;
      68354: inst = 32'h13e00001;
      68355: inst = 32'hfe0d96a;
      68356: inst = 32'h5be00000;
      68357: inst = 32'h8c50000;
      68358: inst = 32'h24612800;
      68359: inst = 32'h10a0ffff;
      68360: inst = 32'hca0fff8;
      68361: inst = 32'h24822800;
      68362: inst = 32'h10a00000;
      68363: inst = 32'hca00004;
      68364: inst = 32'h38632800;
      68365: inst = 32'h38842800;
      68366: inst = 32'h10a00001;
      68367: inst = 32'hca00b13;
      68368: inst = 32'h13e00001;
      68369: inst = 32'hfe0d96a;
      68370: inst = 32'h5be00000;
      68371: inst = 32'h8c50000;
      68372: inst = 32'h24612800;
      68373: inst = 32'h10a0ffff;
      68374: inst = 32'hca0fff8;
      68375: inst = 32'h24822800;
      68376: inst = 32'h10a00000;
      68377: inst = 32'hca00004;
      68378: inst = 32'h38632800;
      68379: inst = 32'h38842800;
      68380: inst = 32'h10a00001;
      68381: inst = 32'hca00b21;
      68382: inst = 32'h13e00001;
      68383: inst = 32'hfe0d96a;
      68384: inst = 32'h5be00000;
      68385: inst = 32'h8c50000;
      68386: inst = 32'h24612800;
      68387: inst = 32'h10a0ffff;
      68388: inst = 32'hca0fff8;
      68389: inst = 32'h24822800;
      68390: inst = 32'h10a00000;
      68391: inst = 32'hca00004;
      68392: inst = 32'h38632800;
      68393: inst = 32'h38842800;
      68394: inst = 32'h10a00001;
      68395: inst = 32'hca00b2f;
      68396: inst = 32'h13e00001;
      68397: inst = 32'hfe0d96a;
      68398: inst = 32'h5be00000;
      68399: inst = 32'h8c50000;
      68400: inst = 32'h24612800;
      68401: inst = 32'h10a0ffff;
      68402: inst = 32'hca0fff8;
      68403: inst = 32'h24822800;
      68404: inst = 32'h10a00000;
      68405: inst = 32'hca00004;
      68406: inst = 32'h38632800;
      68407: inst = 32'h38842800;
      68408: inst = 32'h10a00001;
      68409: inst = 32'hca00b3d;
      68410: inst = 32'h13e00001;
      68411: inst = 32'hfe0d96a;
      68412: inst = 32'h5be00000;
      68413: inst = 32'h8c50000;
      68414: inst = 32'h24612800;
      68415: inst = 32'h10a0ffff;
      68416: inst = 32'hca0fff8;
      68417: inst = 32'h24822800;
      68418: inst = 32'h10a00000;
      68419: inst = 32'hca00004;
      68420: inst = 32'h38632800;
      68421: inst = 32'h38842800;
      68422: inst = 32'h10a00001;
      68423: inst = 32'hca00b4b;
      68424: inst = 32'h13e00001;
      68425: inst = 32'hfe0d96a;
      68426: inst = 32'h5be00000;
      68427: inst = 32'h8c50000;
      68428: inst = 32'h24612800;
      68429: inst = 32'h10a0ffff;
      68430: inst = 32'hca0fff8;
      68431: inst = 32'h24822800;
      68432: inst = 32'h10a00000;
      68433: inst = 32'hca00004;
      68434: inst = 32'h38632800;
      68435: inst = 32'h38842800;
      68436: inst = 32'h10a00001;
      68437: inst = 32'hca00b59;
      68438: inst = 32'h13e00001;
      68439: inst = 32'hfe0d96a;
      68440: inst = 32'h5be00000;
      68441: inst = 32'h8c50000;
      68442: inst = 32'h24612800;
      68443: inst = 32'h10a0ffff;
      68444: inst = 32'hca0fff8;
      68445: inst = 32'h24822800;
      68446: inst = 32'h10a00000;
      68447: inst = 32'hca00004;
      68448: inst = 32'h38632800;
      68449: inst = 32'h38842800;
      68450: inst = 32'h10a00001;
      68451: inst = 32'hca00b67;
      68452: inst = 32'h13e00001;
      68453: inst = 32'hfe0d96a;
      68454: inst = 32'h5be00000;
      68455: inst = 32'h8c50000;
      68456: inst = 32'h24612800;
      68457: inst = 32'h10a0ffff;
      68458: inst = 32'hca0fff8;
      68459: inst = 32'h24822800;
      68460: inst = 32'h10a00000;
      68461: inst = 32'hca00004;
      68462: inst = 32'h38632800;
      68463: inst = 32'h38842800;
      68464: inst = 32'h10a00001;
      68465: inst = 32'hca00b75;
      68466: inst = 32'h13e00001;
      68467: inst = 32'hfe0d96a;
      68468: inst = 32'h5be00000;
      68469: inst = 32'h8c50000;
      68470: inst = 32'h24612800;
      68471: inst = 32'h10a0ffff;
      68472: inst = 32'hca0fff8;
      68473: inst = 32'h24822800;
      68474: inst = 32'h10a00000;
      68475: inst = 32'hca00004;
      68476: inst = 32'h38632800;
      68477: inst = 32'h38842800;
      68478: inst = 32'h10a00001;
      68479: inst = 32'hca00b83;
      68480: inst = 32'h13e00001;
      68481: inst = 32'hfe0d96a;
      68482: inst = 32'h5be00000;
      68483: inst = 32'h8c50000;
      68484: inst = 32'h24612800;
      68485: inst = 32'h10a0ffff;
      68486: inst = 32'hca0fff8;
      68487: inst = 32'h24822800;
      68488: inst = 32'h10a00000;
      68489: inst = 32'hca00004;
      68490: inst = 32'h38632800;
      68491: inst = 32'h38842800;
      68492: inst = 32'h10a00001;
      68493: inst = 32'hca00b91;
      68494: inst = 32'h13e00001;
      68495: inst = 32'hfe0d96a;
      68496: inst = 32'h5be00000;
      68497: inst = 32'h8c50000;
      68498: inst = 32'h24612800;
      68499: inst = 32'h10a0ffff;
      68500: inst = 32'hca0fff8;
      68501: inst = 32'h24822800;
      68502: inst = 32'h10a00000;
      68503: inst = 32'hca00004;
      68504: inst = 32'h38632800;
      68505: inst = 32'h38842800;
      68506: inst = 32'h10a00001;
      68507: inst = 32'hca00b9f;
      68508: inst = 32'h13e00001;
      68509: inst = 32'hfe0d96a;
      68510: inst = 32'h5be00000;
      68511: inst = 32'h8c50000;
      68512: inst = 32'h24612800;
      68513: inst = 32'h10a0ffff;
      68514: inst = 32'hca0fff8;
      68515: inst = 32'h24822800;
      68516: inst = 32'h10a00000;
      68517: inst = 32'hca00004;
      68518: inst = 32'h38632800;
      68519: inst = 32'h38842800;
      68520: inst = 32'h10a00001;
      68521: inst = 32'hca00bad;
      68522: inst = 32'h13e00001;
      68523: inst = 32'hfe0d96a;
      68524: inst = 32'h5be00000;
      68525: inst = 32'h8c50000;
      68526: inst = 32'h24612800;
      68527: inst = 32'h10a0ffff;
      68528: inst = 32'hca0fff8;
      68529: inst = 32'h24822800;
      68530: inst = 32'h10a00000;
      68531: inst = 32'hca00004;
      68532: inst = 32'h38632800;
      68533: inst = 32'h38842800;
      68534: inst = 32'h10a00001;
      68535: inst = 32'hca00bbb;
      68536: inst = 32'h13e00001;
      68537: inst = 32'hfe0d96a;
      68538: inst = 32'h5be00000;
      68539: inst = 32'h8c50000;
      68540: inst = 32'h24612800;
      68541: inst = 32'h10a0ffff;
      68542: inst = 32'hca0fff8;
      68543: inst = 32'h24822800;
      68544: inst = 32'h10a00000;
      68545: inst = 32'hca00004;
      68546: inst = 32'h38632800;
      68547: inst = 32'h38842800;
      68548: inst = 32'h10a00001;
      68549: inst = 32'hca00bc9;
      68550: inst = 32'h13e00001;
      68551: inst = 32'hfe0d96a;
      68552: inst = 32'h5be00000;
      68553: inst = 32'h8c50000;
      68554: inst = 32'h24612800;
      68555: inst = 32'h10a0ffff;
      68556: inst = 32'hca0fff8;
      68557: inst = 32'h24822800;
      68558: inst = 32'h10a00000;
      68559: inst = 32'hca00004;
      68560: inst = 32'h38632800;
      68561: inst = 32'h38842800;
      68562: inst = 32'h10a00001;
      68563: inst = 32'hca00bd7;
      68564: inst = 32'h13e00001;
      68565: inst = 32'hfe0d96a;
      68566: inst = 32'h5be00000;
      68567: inst = 32'h8c50000;
      68568: inst = 32'h24612800;
      68569: inst = 32'h10a0ffff;
      68570: inst = 32'hca0fff8;
      68571: inst = 32'h24822800;
      68572: inst = 32'h10a00000;
      68573: inst = 32'hca00004;
      68574: inst = 32'h38632800;
      68575: inst = 32'h38842800;
      68576: inst = 32'h10a00001;
      68577: inst = 32'hca00be5;
      68578: inst = 32'h13e00001;
      68579: inst = 32'hfe0d96a;
      68580: inst = 32'h5be00000;
      68581: inst = 32'h8c50000;
      68582: inst = 32'h24612800;
      68583: inst = 32'h10a0ffff;
      68584: inst = 32'hca0fff8;
      68585: inst = 32'h24822800;
      68586: inst = 32'h10a00000;
      68587: inst = 32'hca00004;
      68588: inst = 32'h38632800;
      68589: inst = 32'h38842800;
      68590: inst = 32'h10a00001;
      68591: inst = 32'hca00bf3;
      68592: inst = 32'h13e00001;
      68593: inst = 32'hfe0d96a;
      68594: inst = 32'h5be00000;
      68595: inst = 32'h8c50000;
      68596: inst = 32'h24612800;
      68597: inst = 32'h10a0ffff;
      68598: inst = 32'hca0fff8;
      68599: inst = 32'h24822800;
      68600: inst = 32'h10a00000;
      68601: inst = 32'hca00004;
      68602: inst = 32'h38632800;
      68603: inst = 32'h38842800;
      68604: inst = 32'h10a00001;
      68605: inst = 32'hca00c01;
      68606: inst = 32'h13e00001;
      68607: inst = 32'hfe0d96a;
      68608: inst = 32'h5be00000;
      68609: inst = 32'h8c50000;
      68610: inst = 32'h24612800;
      68611: inst = 32'h10a0ffff;
      68612: inst = 32'hca0fff8;
      68613: inst = 32'h24822800;
      68614: inst = 32'h10a00000;
      68615: inst = 32'hca00004;
      68616: inst = 32'h38632800;
      68617: inst = 32'h38842800;
      68618: inst = 32'h10a00001;
      68619: inst = 32'hca00c0f;
      68620: inst = 32'h13e00001;
      68621: inst = 32'hfe0d96a;
      68622: inst = 32'h5be00000;
      68623: inst = 32'h8c50000;
      68624: inst = 32'h24612800;
      68625: inst = 32'h10a0ffff;
      68626: inst = 32'hca0fff8;
      68627: inst = 32'h24822800;
      68628: inst = 32'h10a00000;
      68629: inst = 32'hca00004;
      68630: inst = 32'h38632800;
      68631: inst = 32'h38842800;
      68632: inst = 32'h10a00001;
      68633: inst = 32'hca00c1d;
      68634: inst = 32'h13e00001;
      68635: inst = 32'hfe0d96a;
      68636: inst = 32'h5be00000;
      68637: inst = 32'h8c50000;
      68638: inst = 32'h24612800;
      68639: inst = 32'h10a0ffff;
      68640: inst = 32'hca0fff8;
      68641: inst = 32'h24822800;
      68642: inst = 32'h10a00000;
      68643: inst = 32'hca00004;
      68644: inst = 32'h38632800;
      68645: inst = 32'h38842800;
      68646: inst = 32'h10a00001;
      68647: inst = 32'hca00c2b;
      68648: inst = 32'h13e00001;
      68649: inst = 32'hfe0d96a;
      68650: inst = 32'h5be00000;
      68651: inst = 32'h8c50000;
      68652: inst = 32'h24612800;
      68653: inst = 32'h10a0ffff;
      68654: inst = 32'hca0fff8;
      68655: inst = 32'h24822800;
      68656: inst = 32'h10a00000;
      68657: inst = 32'hca00004;
      68658: inst = 32'h38632800;
      68659: inst = 32'h38842800;
      68660: inst = 32'h10a00001;
      68661: inst = 32'hca00c39;
      68662: inst = 32'h13e00001;
      68663: inst = 32'hfe0d96a;
      68664: inst = 32'h5be00000;
      68665: inst = 32'h8c50000;
      68666: inst = 32'h24612800;
      68667: inst = 32'h10a0ffff;
      68668: inst = 32'hca0fff8;
      68669: inst = 32'h24822800;
      68670: inst = 32'h10a00000;
      68671: inst = 32'hca00004;
      68672: inst = 32'h38632800;
      68673: inst = 32'h38842800;
      68674: inst = 32'h10a00001;
      68675: inst = 32'hca00c47;
      68676: inst = 32'h13e00001;
      68677: inst = 32'hfe0d96a;
      68678: inst = 32'h5be00000;
      68679: inst = 32'h8c50000;
      68680: inst = 32'h24612800;
      68681: inst = 32'h10a0ffff;
      68682: inst = 32'hca0fff8;
      68683: inst = 32'h24822800;
      68684: inst = 32'h10a00000;
      68685: inst = 32'hca00004;
      68686: inst = 32'h38632800;
      68687: inst = 32'h38842800;
      68688: inst = 32'h10a00001;
      68689: inst = 32'hca00c55;
      68690: inst = 32'h13e00001;
      68691: inst = 32'hfe0d96a;
      68692: inst = 32'h5be00000;
      68693: inst = 32'h8c50000;
      68694: inst = 32'h24612800;
      68695: inst = 32'h10a0ffff;
      68696: inst = 32'hca0fff8;
      68697: inst = 32'h24822800;
      68698: inst = 32'h10a00000;
      68699: inst = 32'hca00004;
      68700: inst = 32'h38632800;
      68701: inst = 32'h38842800;
      68702: inst = 32'h10a00001;
      68703: inst = 32'hca00c63;
      68704: inst = 32'h13e00001;
      68705: inst = 32'hfe0d96a;
      68706: inst = 32'h5be00000;
      68707: inst = 32'h8c50000;
      68708: inst = 32'h24612800;
      68709: inst = 32'h10a0ffff;
      68710: inst = 32'hca0fff8;
      68711: inst = 32'h24822800;
      68712: inst = 32'h10a00000;
      68713: inst = 32'hca00004;
      68714: inst = 32'h38632800;
      68715: inst = 32'h38842800;
      68716: inst = 32'h10a00001;
      68717: inst = 32'hca00c71;
      68718: inst = 32'h13e00001;
      68719: inst = 32'hfe0d96a;
      68720: inst = 32'h5be00000;
      68721: inst = 32'h8c50000;
      68722: inst = 32'h24612800;
      68723: inst = 32'h10a0ffff;
      68724: inst = 32'hca0fff8;
      68725: inst = 32'h24822800;
      68726: inst = 32'h10a00000;
      68727: inst = 32'hca00004;
      68728: inst = 32'h38632800;
      68729: inst = 32'h38842800;
      68730: inst = 32'h10a00001;
      68731: inst = 32'hca00c7f;
      68732: inst = 32'h13e00001;
      68733: inst = 32'hfe0d96a;
      68734: inst = 32'h5be00000;
      68735: inst = 32'h8c50000;
      68736: inst = 32'h24612800;
      68737: inst = 32'h10a0ffff;
      68738: inst = 32'hca0fff8;
      68739: inst = 32'h24822800;
      68740: inst = 32'h10a00000;
      68741: inst = 32'hca00004;
      68742: inst = 32'h38632800;
      68743: inst = 32'h38842800;
      68744: inst = 32'h10a00001;
      68745: inst = 32'hca00c8d;
      68746: inst = 32'h13e00001;
      68747: inst = 32'hfe0d96a;
      68748: inst = 32'h5be00000;
      68749: inst = 32'h8c50000;
      68750: inst = 32'h24612800;
      68751: inst = 32'h10a0ffff;
      68752: inst = 32'hca0fff8;
      68753: inst = 32'h24822800;
      68754: inst = 32'h10a00000;
      68755: inst = 32'hca00004;
      68756: inst = 32'h38632800;
      68757: inst = 32'h38842800;
      68758: inst = 32'h10a00001;
      68759: inst = 32'hca00c9b;
      68760: inst = 32'h13e00001;
      68761: inst = 32'hfe0d96a;
      68762: inst = 32'h5be00000;
      68763: inst = 32'h8c50000;
      68764: inst = 32'h24612800;
      68765: inst = 32'h10a0ffff;
      68766: inst = 32'hca0fff8;
      68767: inst = 32'h24822800;
      68768: inst = 32'h10a00000;
      68769: inst = 32'hca00004;
      68770: inst = 32'h38632800;
      68771: inst = 32'h38842800;
      68772: inst = 32'h10a00001;
      68773: inst = 32'hca00ca9;
      68774: inst = 32'h13e00001;
      68775: inst = 32'hfe0d96a;
      68776: inst = 32'h5be00000;
      68777: inst = 32'h8c50000;
      68778: inst = 32'h24612800;
      68779: inst = 32'h10a0ffff;
      68780: inst = 32'hca0fff9;
      68781: inst = 32'h24822800;
      68782: inst = 32'h10a00000;
      68783: inst = 32'hca00004;
      68784: inst = 32'h38632800;
      68785: inst = 32'h38842800;
      68786: inst = 32'h10a00001;
      68787: inst = 32'hca00cb7;
      68788: inst = 32'h13e00001;
      68789: inst = 32'hfe0d96a;
      68790: inst = 32'h5be00000;
      68791: inst = 32'h8c50000;
      68792: inst = 32'h24612800;
      68793: inst = 32'h10a0ffff;
      68794: inst = 32'hca0fff9;
      68795: inst = 32'h24822800;
      68796: inst = 32'h10a00000;
      68797: inst = 32'hca00004;
      68798: inst = 32'h38632800;
      68799: inst = 32'h38842800;
      68800: inst = 32'h10a00001;
      68801: inst = 32'hca00cc5;
      68802: inst = 32'h13e00001;
      68803: inst = 32'hfe0d96a;
      68804: inst = 32'h5be00000;
      68805: inst = 32'h8c50000;
      68806: inst = 32'h24612800;
      68807: inst = 32'h10a0ffff;
      68808: inst = 32'hca0fff9;
      68809: inst = 32'h24822800;
      68810: inst = 32'h10a00000;
      68811: inst = 32'hca00004;
      68812: inst = 32'h38632800;
      68813: inst = 32'h38842800;
      68814: inst = 32'h10a00001;
      68815: inst = 32'hca00cd3;
      68816: inst = 32'h13e00001;
      68817: inst = 32'hfe0d96a;
      68818: inst = 32'h5be00000;
      68819: inst = 32'h8c50000;
      68820: inst = 32'h24612800;
      68821: inst = 32'h10a0ffff;
      68822: inst = 32'hca0fff9;
      68823: inst = 32'h24822800;
      68824: inst = 32'h10a00000;
      68825: inst = 32'hca00004;
      68826: inst = 32'h38632800;
      68827: inst = 32'h38842800;
      68828: inst = 32'h10a00001;
      68829: inst = 32'hca00ce1;
      68830: inst = 32'h13e00001;
      68831: inst = 32'hfe0d96a;
      68832: inst = 32'h5be00000;
      68833: inst = 32'h8c50000;
      68834: inst = 32'h24612800;
      68835: inst = 32'h10a0ffff;
      68836: inst = 32'hca0fff9;
      68837: inst = 32'h24822800;
      68838: inst = 32'h10a00000;
      68839: inst = 32'hca00004;
      68840: inst = 32'h38632800;
      68841: inst = 32'h38842800;
      68842: inst = 32'h10a00001;
      68843: inst = 32'hca00cef;
      68844: inst = 32'h13e00001;
      68845: inst = 32'hfe0d96a;
      68846: inst = 32'h5be00000;
      68847: inst = 32'h8c50000;
      68848: inst = 32'h24612800;
      68849: inst = 32'h10a0ffff;
      68850: inst = 32'hca0fff9;
      68851: inst = 32'h24822800;
      68852: inst = 32'h10a00000;
      68853: inst = 32'hca00004;
      68854: inst = 32'h38632800;
      68855: inst = 32'h38842800;
      68856: inst = 32'h10a00001;
      68857: inst = 32'hca00cfd;
      68858: inst = 32'h13e00001;
      68859: inst = 32'hfe0d96a;
      68860: inst = 32'h5be00000;
      68861: inst = 32'h8c50000;
      68862: inst = 32'h24612800;
      68863: inst = 32'h10a0ffff;
      68864: inst = 32'hca0fff9;
      68865: inst = 32'h24822800;
      68866: inst = 32'h10a00000;
      68867: inst = 32'hca00004;
      68868: inst = 32'h38632800;
      68869: inst = 32'h38842800;
      68870: inst = 32'h10a00001;
      68871: inst = 32'hca00d0b;
      68872: inst = 32'h13e00001;
      68873: inst = 32'hfe0d96a;
      68874: inst = 32'h5be00000;
      68875: inst = 32'h8c50000;
      68876: inst = 32'h24612800;
      68877: inst = 32'h10a0ffff;
      68878: inst = 32'hca0fff9;
      68879: inst = 32'h24822800;
      68880: inst = 32'h10a00000;
      68881: inst = 32'hca00004;
      68882: inst = 32'h38632800;
      68883: inst = 32'h38842800;
      68884: inst = 32'h10a00001;
      68885: inst = 32'hca00d19;
      68886: inst = 32'h13e00001;
      68887: inst = 32'hfe0d96a;
      68888: inst = 32'h5be00000;
      68889: inst = 32'h8c50000;
      68890: inst = 32'h24612800;
      68891: inst = 32'h10a0ffff;
      68892: inst = 32'hca0fff9;
      68893: inst = 32'h24822800;
      68894: inst = 32'h10a00000;
      68895: inst = 32'hca00004;
      68896: inst = 32'h38632800;
      68897: inst = 32'h38842800;
      68898: inst = 32'h10a00001;
      68899: inst = 32'hca00d27;
      68900: inst = 32'h13e00001;
      68901: inst = 32'hfe0d96a;
      68902: inst = 32'h5be00000;
      68903: inst = 32'h8c50000;
      68904: inst = 32'h24612800;
      68905: inst = 32'h10a0ffff;
      68906: inst = 32'hca0fff9;
      68907: inst = 32'h24822800;
      68908: inst = 32'h10a00000;
      68909: inst = 32'hca00004;
      68910: inst = 32'h38632800;
      68911: inst = 32'h38842800;
      68912: inst = 32'h10a00001;
      68913: inst = 32'hca00d35;
      68914: inst = 32'h13e00001;
      68915: inst = 32'hfe0d96a;
      68916: inst = 32'h5be00000;
      68917: inst = 32'h8c50000;
      68918: inst = 32'h24612800;
      68919: inst = 32'h10a0ffff;
      68920: inst = 32'hca0fff9;
      68921: inst = 32'h24822800;
      68922: inst = 32'h10a00000;
      68923: inst = 32'hca00004;
      68924: inst = 32'h38632800;
      68925: inst = 32'h38842800;
      68926: inst = 32'h10a00001;
      68927: inst = 32'hca00d43;
      68928: inst = 32'h13e00001;
      68929: inst = 32'hfe0d96a;
      68930: inst = 32'h5be00000;
      68931: inst = 32'h8c50000;
      68932: inst = 32'h24612800;
      68933: inst = 32'h10a0ffff;
      68934: inst = 32'hca0fff9;
      68935: inst = 32'h24822800;
      68936: inst = 32'h10a00000;
      68937: inst = 32'hca00004;
      68938: inst = 32'h38632800;
      68939: inst = 32'h38842800;
      68940: inst = 32'h10a00001;
      68941: inst = 32'hca00d51;
      68942: inst = 32'h13e00001;
      68943: inst = 32'hfe0d96a;
      68944: inst = 32'h5be00000;
      68945: inst = 32'h8c50000;
      68946: inst = 32'h24612800;
      68947: inst = 32'h10a0ffff;
      68948: inst = 32'hca0fff9;
      68949: inst = 32'h24822800;
      68950: inst = 32'h10a00000;
      68951: inst = 32'hca00004;
      68952: inst = 32'h38632800;
      68953: inst = 32'h38842800;
      68954: inst = 32'h10a00001;
      68955: inst = 32'hca00d5f;
      68956: inst = 32'h13e00001;
      68957: inst = 32'hfe0d96a;
      68958: inst = 32'h5be00000;
      68959: inst = 32'h8c50000;
      68960: inst = 32'h24612800;
      68961: inst = 32'h10a0ffff;
      68962: inst = 32'hca0fff9;
      68963: inst = 32'h24822800;
      68964: inst = 32'h10a00000;
      68965: inst = 32'hca00004;
      68966: inst = 32'h38632800;
      68967: inst = 32'h38842800;
      68968: inst = 32'h10a00001;
      68969: inst = 32'hca00d6d;
      68970: inst = 32'h13e00001;
      68971: inst = 32'hfe0d96a;
      68972: inst = 32'h5be00000;
      68973: inst = 32'h8c50000;
      68974: inst = 32'h24612800;
      68975: inst = 32'h10a0ffff;
      68976: inst = 32'hca0fff9;
      68977: inst = 32'h24822800;
      68978: inst = 32'h10a00000;
      68979: inst = 32'hca00004;
      68980: inst = 32'h38632800;
      68981: inst = 32'h38842800;
      68982: inst = 32'h10a00001;
      68983: inst = 32'hca00d7b;
      68984: inst = 32'h13e00001;
      68985: inst = 32'hfe0d96a;
      68986: inst = 32'h5be00000;
      68987: inst = 32'h8c50000;
      68988: inst = 32'h24612800;
      68989: inst = 32'h10a0ffff;
      68990: inst = 32'hca0fff9;
      68991: inst = 32'h24822800;
      68992: inst = 32'h10a00000;
      68993: inst = 32'hca00004;
      68994: inst = 32'h38632800;
      68995: inst = 32'h38842800;
      68996: inst = 32'h10a00001;
      68997: inst = 32'hca00d89;
      68998: inst = 32'h13e00001;
      68999: inst = 32'hfe0d96a;
      69000: inst = 32'h5be00000;
      69001: inst = 32'h8c50000;
      69002: inst = 32'h24612800;
      69003: inst = 32'h10a0ffff;
      69004: inst = 32'hca0fff9;
      69005: inst = 32'h24822800;
      69006: inst = 32'h10a00000;
      69007: inst = 32'hca00004;
      69008: inst = 32'h38632800;
      69009: inst = 32'h38842800;
      69010: inst = 32'h10a00001;
      69011: inst = 32'hca00d97;
      69012: inst = 32'h13e00001;
      69013: inst = 32'hfe0d96a;
      69014: inst = 32'h5be00000;
      69015: inst = 32'h8c50000;
      69016: inst = 32'h24612800;
      69017: inst = 32'h10a0ffff;
      69018: inst = 32'hca0fff9;
      69019: inst = 32'h24822800;
      69020: inst = 32'h10a00000;
      69021: inst = 32'hca00004;
      69022: inst = 32'h38632800;
      69023: inst = 32'h38842800;
      69024: inst = 32'h10a00001;
      69025: inst = 32'hca00da5;
      69026: inst = 32'h13e00001;
      69027: inst = 32'hfe0d96a;
      69028: inst = 32'h5be00000;
      69029: inst = 32'h8c50000;
      69030: inst = 32'h24612800;
      69031: inst = 32'h10a0ffff;
      69032: inst = 32'hca0fff9;
      69033: inst = 32'h24822800;
      69034: inst = 32'h10a00000;
      69035: inst = 32'hca00004;
      69036: inst = 32'h38632800;
      69037: inst = 32'h38842800;
      69038: inst = 32'h10a00001;
      69039: inst = 32'hca00db3;
      69040: inst = 32'h13e00001;
      69041: inst = 32'hfe0d96a;
      69042: inst = 32'h5be00000;
      69043: inst = 32'h8c50000;
      69044: inst = 32'h24612800;
      69045: inst = 32'h10a0ffff;
      69046: inst = 32'hca0fff9;
      69047: inst = 32'h24822800;
      69048: inst = 32'h10a00000;
      69049: inst = 32'hca00004;
      69050: inst = 32'h38632800;
      69051: inst = 32'h38842800;
      69052: inst = 32'h10a00001;
      69053: inst = 32'hca00dc1;
      69054: inst = 32'h13e00001;
      69055: inst = 32'hfe0d96a;
      69056: inst = 32'h5be00000;
      69057: inst = 32'h8c50000;
      69058: inst = 32'h24612800;
      69059: inst = 32'h10a0ffff;
      69060: inst = 32'hca0fff9;
      69061: inst = 32'h24822800;
      69062: inst = 32'h10a00000;
      69063: inst = 32'hca00004;
      69064: inst = 32'h38632800;
      69065: inst = 32'h38842800;
      69066: inst = 32'h10a00001;
      69067: inst = 32'hca00dcf;
      69068: inst = 32'h13e00001;
      69069: inst = 32'hfe0d96a;
      69070: inst = 32'h5be00000;
      69071: inst = 32'h8c50000;
      69072: inst = 32'h24612800;
      69073: inst = 32'h10a0ffff;
      69074: inst = 32'hca0fff9;
      69075: inst = 32'h24822800;
      69076: inst = 32'h10a00000;
      69077: inst = 32'hca00004;
      69078: inst = 32'h38632800;
      69079: inst = 32'h38842800;
      69080: inst = 32'h10a00001;
      69081: inst = 32'hca00ddd;
      69082: inst = 32'h13e00001;
      69083: inst = 32'hfe0d96a;
      69084: inst = 32'h5be00000;
      69085: inst = 32'h8c50000;
      69086: inst = 32'h24612800;
      69087: inst = 32'h10a0ffff;
      69088: inst = 32'hca0fff9;
      69089: inst = 32'h24822800;
      69090: inst = 32'h10a00000;
      69091: inst = 32'hca00004;
      69092: inst = 32'h38632800;
      69093: inst = 32'h38842800;
      69094: inst = 32'h10a00001;
      69095: inst = 32'hca00deb;
      69096: inst = 32'h13e00001;
      69097: inst = 32'hfe0d96a;
      69098: inst = 32'h5be00000;
      69099: inst = 32'h8c50000;
      69100: inst = 32'h24612800;
      69101: inst = 32'h10a0ffff;
      69102: inst = 32'hca0fff9;
      69103: inst = 32'h24822800;
      69104: inst = 32'h10a00000;
      69105: inst = 32'hca00004;
      69106: inst = 32'h38632800;
      69107: inst = 32'h38842800;
      69108: inst = 32'h10a00001;
      69109: inst = 32'hca00df9;
      69110: inst = 32'h13e00001;
      69111: inst = 32'hfe0d96a;
      69112: inst = 32'h5be00000;
      69113: inst = 32'h8c50000;
      69114: inst = 32'h24612800;
      69115: inst = 32'h10a0ffff;
      69116: inst = 32'hca0fff9;
      69117: inst = 32'h24822800;
      69118: inst = 32'h10a00000;
      69119: inst = 32'hca00004;
      69120: inst = 32'h38632800;
      69121: inst = 32'h38842800;
      69122: inst = 32'h10a00001;
      69123: inst = 32'hca00e07;
      69124: inst = 32'h13e00001;
      69125: inst = 32'hfe0d96a;
      69126: inst = 32'h5be00000;
      69127: inst = 32'h8c50000;
      69128: inst = 32'h24612800;
      69129: inst = 32'h10a0ffff;
      69130: inst = 32'hca0fff9;
      69131: inst = 32'h24822800;
      69132: inst = 32'h10a00000;
      69133: inst = 32'hca00004;
      69134: inst = 32'h38632800;
      69135: inst = 32'h38842800;
      69136: inst = 32'h10a00001;
      69137: inst = 32'hca00e15;
      69138: inst = 32'h13e00001;
      69139: inst = 32'hfe0d96a;
      69140: inst = 32'h5be00000;
      69141: inst = 32'h8c50000;
      69142: inst = 32'h24612800;
      69143: inst = 32'h10a0ffff;
      69144: inst = 32'hca0fff9;
      69145: inst = 32'h24822800;
      69146: inst = 32'h10a00000;
      69147: inst = 32'hca00004;
      69148: inst = 32'h38632800;
      69149: inst = 32'h38842800;
      69150: inst = 32'h10a00001;
      69151: inst = 32'hca00e23;
      69152: inst = 32'h13e00001;
      69153: inst = 32'hfe0d96a;
      69154: inst = 32'h5be00000;
      69155: inst = 32'h8c50000;
      69156: inst = 32'h24612800;
      69157: inst = 32'h10a0ffff;
      69158: inst = 32'hca0fff9;
      69159: inst = 32'h24822800;
      69160: inst = 32'h10a00000;
      69161: inst = 32'hca00004;
      69162: inst = 32'h38632800;
      69163: inst = 32'h38842800;
      69164: inst = 32'h10a00001;
      69165: inst = 32'hca00e31;
      69166: inst = 32'h13e00001;
      69167: inst = 32'hfe0d96a;
      69168: inst = 32'h5be00000;
      69169: inst = 32'h8c50000;
      69170: inst = 32'h24612800;
      69171: inst = 32'h10a0ffff;
      69172: inst = 32'hca0fff9;
      69173: inst = 32'h24822800;
      69174: inst = 32'h10a00000;
      69175: inst = 32'hca00004;
      69176: inst = 32'h38632800;
      69177: inst = 32'h38842800;
      69178: inst = 32'h10a00001;
      69179: inst = 32'hca00e3f;
      69180: inst = 32'h13e00001;
      69181: inst = 32'hfe0d96a;
      69182: inst = 32'h5be00000;
      69183: inst = 32'h8c50000;
      69184: inst = 32'h24612800;
      69185: inst = 32'h10a0ffff;
      69186: inst = 32'hca0fff9;
      69187: inst = 32'h24822800;
      69188: inst = 32'h10a00000;
      69189: inst = 32'hca00004;
      69190: inst = 32'h38632800;
      69191: inst = 32'h38842800;
      69192: inst = 32'h10a00001;
      69193: inst = 32'hca00e4d;
      69194: inst = 32'h13e00001;
      69195: inst = 32'hfe0d96a;
      69196: inst = 32'h5be00000;
      69197: inst = 32'h8c50000;
      69198: inst = 32'h24612800;
      69199: inst = 32'h10a0ffff;
      69200: inst = 32'hca0fff9;
      69201: inst = 32'h24822800;
      69202: inst = 32'h10a00000;
      69203: inst = 32'hca00004;
      69204: inst = 32'h38632800;
      69205: inst = 32'h38842800;
      69206: inst = 32'h10a00001;
      69207: inst = 32'hca00e5b;
      69208: inst = 32'h13e00001;
      69209: inst = 32'hfe0d96a;
      69210: inst = 32'h5be00000;
      69211: inst = 32'h8c50000;
      69212: inst = 32'h24612800;
      69213: inst = 32'h10a0ffff;
      69214: inst = 32'hca0fff9;
      69215: inst = 32'h24822800;
      69216: inst = 32'h10a00000;
      69217: inst = 32'hca00004;
      69218: inst = 32'h38632800;
      69219: inst = 32'h38842800;
      69220: inst = 32'h10a00001;
      69221: inst = 32'hca00e69;
      69222: inst = 32'h13e00001;
      69223: inst = 32'hfe0d96a;
      69224: inst = 32'h5be00000;
      69225: inst = 32'h8c50000;
      69226: inst = 32'h24612800;
      69227: inst = 32'h10a0ffff;
      69228: inst = 32'hca0fff9;
      69229: inst = 32'h24822800;
      69230: inst = 32'h10a00000;
      69231: inst = 32'hca00004;
      69232: inst = 32'h38632800;
      69233: inst = 32'h38842800;
      69234: inst = 32'h10a00001;
      69235: inst = 32'hca00e77;
      69236: inst = 32'h13e00001;
      69237: inst = 32'hfe0d96a;
      69238: inst = 32'h5be00000;
      69239: inst = 32'h8c50000;
      69240: inst = 32'h24612800;
      69241: inst = 32'h10a0ffff;
      69242: inst = 32'hca0fff9;
      69243: inst = 32'h24822800;
      69244: inst = 32'h10a00000;
      69245: inst = 32'hca00004;
      69246: inst = 32'h38632800;
      69247: inst = 32'h38842800;
      69248: inst = 32'h10a00001;
      69249: inst = 32'hca00e85;
      69250: inst = 32'h13e00001;
      69251: inst = 32'hfe0d96a;
      69252: inst = 32'h5be00000;
      69253: inst = 32'h8c50000;
      69254: inst = 32'h24612800;
      69255: inst = 32'h10a0ffff;
      69256: inst = 32'hca0fff9;
      69257: inst = 32'h24822800;
      69258: inst = 32'h10a00000;
      69259: inst = 32'hca00004;
      69260: inst = 32'h38632800;
      69261: inst = 32'h38842800;
      69262: inst = 32'h10a00001;
      69263: inst = 32'hca00e93;
      69264: inst = 32'h13e00001;
      69265: inst = 32'hfe0d96a;
      69266: inst = 32'h5be00000;
      69267: inst = 32'h8c50000;
      69268: inst = 32'h24612800;
      69269: inst = 32'h10a0ffff;
      69270: inst = 32'hca0fff9;
      69271: inst = 32'h24822800;
      69272: inst = 32'h10a00000;
      69273: inst = 32'hca00004;
      69274: inst = 32'h38632800;
      69275: inst = 32'h38842800;
      69276: inst = 32'h10a00001;
      69277: inst = 32'hca00ea1;
      69278: inst = 32'h13e00001;
      69279: inst = 32'hfe0d96a;
      69280: inst = 32'h5be00000;
      69281: inst = 32'h8c50000;
      69282: inst = 32'h24612800;
      69283: inst = 32'h10a0ffff;
      69284: inst = 32'hca0fff9;
      69285: inst = 32'h24822800;
      69286: inst = 32'h10a00000;
      69287: inst = 32'hca00004;
      69288: inst = 32'h38632800;
      69289: inst = 32'h38842800;
      69290: inst = 32'h10a00001;
      69291: inst = 32'hca00eaf;
      69292: inst = 32'h13e00001;
      69293: inst = 32'hfe0d96a;
      69294: inst = 32'h5be00000;
      69295: inst = 32'h8c50000;
      69296: inst = 32'h24612800;
      69297: inst = 32'h10a0ffff;
      69298: inst = 32'hca0fff9;
      69299: inst = 32'h24822800;
      69300: inst = 32'h10a00000;
      69301: inst = 32'hca00004;
      69302: inst = 32'h38632800;
      69303: inst = 32'h38842800;
      69304: inst = 32'h10a00001;
      69305: inst = 32'hca00ebd;
      69306: inst = 32'h13e00001;
      69307: inst = 32'hfe0d96a;
      69308: inst = 32'h5be00000;
      69309: inst = 32'h8c50000;
      69310: inst = 32'h24612800;
      69311: inst = 32'h10a0ffff;
      69312: inst = 32'hca0fff9;
      69313: inst = 32'h24822800;
      69314: inst = 32'h10a00000;
      69315: inst = 32'hca00004;
      69316: inst = 32'h38632800;
      69317: inst = 32'h38842800;
      69318: inst = 32'h10a00001;
      69319: inst = 32'hca00ecb;
      69320: inst = 32'h13e00001;
      69321: inst = 32'hfe0d96a;
      69322: inst = 32'h5be00000;
      69323: inst = 32'h8c50000;
      69324: inst = 32'h24612800;
      69325: inst = 32'h10a0ffff;
      69326: inst = 32'hca0fff9;
      69327: inst = 32'h24822800;
      69328: inst = 32'h10a00000;
      69329: inst = 32'hca00004;
      69330: inst = 32'h38632800;
      69331: inst = 32'h38842800;
      69332: inst = 32'h10a00001;
      69333: inst = 32'hca00ed9;
      69334: inst = 32'h13e00001;
      69335: inst = 32'hfe0d96a;
      69336: inst = 32'h5be00000;
      69337: inst = 32'h8c50000;
      69338: inst = 32'h24612800;
      69339: inst = 32'h10a0ffff;
      69340: inst = 32'hca0fff9;
      69341: inst = 32'h24822800;
      69342: inst = 32'h10a00000;
      69343: inst = 32'hca00004;
      69344: inst = 32'h38632800;
      69345: inst = 32'h38842800;
      69346: inst = 32'h10a00001;
      69347: inst = 32'hca00ee7;
      69348: inst = 32'h13e00001;
      69349: inst = 32'hfe0d96a;
      69350: inst = 32'h5be00000;
      69351: inst = 32'h8c50000;
      69352: inst = 32'h24612800;
      69353: inst = 32'h10a0ffff;
      69354: inst = 32'hca0fff9;
      69355: inst = 32'h24822800;
      69356: inst = 32'h10a00000;
      69357: inst = 32'hca00004;
      69358: inst = 32'h38632800;
      69359: inst = 32'h38842800;
      69360: inst = 32'h10a00001;
      69361: inst = 32'hca00ef5;
      69362: inst = 32'h13e00001;
      69363: inst = 32'hfe0d96a;
      69364: inst = 32'h5be00000;
      69365: inst = 32'h8c50000;
      69366: inst = 32'h24612800;
      69367: inst = 32'h10a0ffff;
      69368: inst = 32'hca0fff9;
      69369: inst = 32'h24822800;
      69370: inst = 32'h10a00000;
      69371: inst = 32'hca00004;
      69372: inst = 32'h38632800;
      69373: inst = 32'h38842800;
      69374: inst = 32'h10a00001;
      69375: inst = 32'hca00f03;
      69376: inst = 32'h13e00001;
      69377: inst = 32'hfe0d96a;
      69378: inst = 32'h5be00000;
      69379: inst = 32'h8c50000;
      69380: inst = 32'h24612800;
      69381: inst = 32'h10a0ffff;
      69382: inst = 32'hca0fff9;
      69383: inst = 32'h24822800;
      69384: inst = 32'h10a00000;
      69385: inst = 32'hca00004;
      69386: inst = 32'h38632800;
      69387: inst = 32'h38842800;
      69388: inst = 32'h10a00001;
      69389: inst = 32'hca00f11;
      69390: inst = 32'h13e00001;
      69391: inst = 32'hfe0d96a;
      69392: inst = 32'h5be00000;
      69393: inst = 32'h8c50000;
      69394: inst = 32'h24612800;
      69395: inst = 32'h10a0ffff;
      69396: inst = 32'hca0fff9;
      69397: inst = 32'h24822800;
      69398: inst = 32'h10a00000;
      69399: inst = 32'hca00004;
      69400: inst = 32'h38632800;
      69401: inst = 32'h38842800;
      69402: inst = 32'h10a00001;
      69403: inst = 32'hca00f1f;
      69404: inst = 32'h13e00001;
      69405: inst = 32'hfe0d96a;
      69406: inst = 32'h5be00000;
      69407: inst = 32'h8c50000;
      69408: inst = 32'h24612800;
      69409: inst = 32'h10a0ffff;
      69410: inst = 32'hca0fff9;
      69411: inst = 32'h24822800;
      69412: inst = 32'h10a00000;
      69413: inst = 32'hca00004;
      69414: inst = 32'h38632800;
      69415: inst = 32'h38842800;
      69416: inst = 32'h10a00001;
      69417: inst = 32'hca00f2d;
      69418: inst = 32'h13e00001;
      69419: inst = 32'hfe0d96a;
      69420: inst = 32'h5be00000;
      69421: inst = 32'h8c50000;
      69422: inst = 32'h24612800;
      69423: inst = 32'h10a0ffff;
      69424: inst = 32'hca0fff9;
      69425: inst = 32'h24822800;
      69426: inst = 32'h10a00000;
      69427: inst = 32'hca00004;
      69428: inst = 32'h38632800;
      69429: inst = 32'h38842800;
      69430: inst = 32'h10a00001;
      69431: inst = 32'hca00f3b;
      69432: inst = 32'h13e00001;
      69433: inst = 32'hfe0d96a;
      69434: inst = 32'h5be00000;
      69435: inst = 32'h8c50000;
      69436: inst = 32'h24612800;
      69437: inst = 32'h10a0ffff;
      69438: inst = 32'hca0fff9;
      69439: inst = 32'h24822800;
      69440: inst = 32'h10a00000;
      69441: inst = 32'hca00004;
      69442: inst = 32'h38632800;
      69443: inst = 32'h38842800;
      69444: inst = 32'h10a00001;
      69445: inst = 32'hca00f49;
      69446: inst = 32'h13e00001;
      69447: inst = 32'hfe0d96a;
      69448: inst = 32'h5be00000;
      69449: inst = 32'h8c50000;
      69450: inst = 32'h24612800;
      69451: inst = 32'h10a0ffff;
      69452: inst = 32'hca0fff9;
      69453: inst = 32'h24822800;
      69454: inst = 32'h10a00000;
      69455: inst = 32'hca00004;
      69456: inst = 32'h38632800;
      69457: inst = 32'h38842800;
      69458: inst = 32'h10a00001;
      69459: inst = 32'hca00f57;
      69460: inst = 32'h13e00001;
      69461: inst = 32'hfe0d96a;
      69462: inst = 32'h5be00000;
      69463: inst = 32'h8c50000;
      69464: inst = 32'h24612800;
      69465: inst = 32'h10a0ffff;
      69466: inst = 32'hca0fff9;
      69467: inst = 32'h24822800;
      69468: inst = 32'h10a00000;
      69469: inst = 32'hca00004;
      69470: inst = 32'h38632800;
      69471: inst = 32'h38842800;
      69472: inst = 32'h10a00001;
      69473: inst = 32'hca00f65;
      69474: inst = 32'h13e00001;
      69475: inst = 32'hfe0d96a;
      69476: inst = 32'h5be00000;
      69477: inst = 32'h8c50000;
      69478: inst = 32'h24612800;
      69479: inst = 32'h10a0ffff;
      69480: inst = 32'hca0fff9;
      69481: inst = 32'h24822800;
      69482: inst = 32'h10a00000;
      69483: inst = 32'hca00004;
      69484: inst = 32'h38632800;
      69485: inst = 32'h38842800;
      69486: inst = 32'h10a00001;
      69487: inst = 32'hca00f73;
      69488: inst = 32'h13e00001;
      69489: inst = 32'hfe0d96a;
      69490: inst = 32'h5be00000;
      69491: inst = 32'h8c50000;
      69492: inst = 32'h24612800;
      69493: inst = 32'h10a0ffff;
      69494: inst = 32'hca0fff9;
      69495: inst = 32'h24822800;
      69496: inst = 32'h10a00000;
      69497: inst = 32'hca00004;
      69498: inst = 32'h38632800;
      69499: inst = 32'h38842800;
      69500: inst = 32'h10a00001;
      69501: inst = 32'hca00f81;
      69502: inst = 32'h13e00001;
      69503: inst = 32'hfe0d96a;
      69504: inst = 32'h5be00000;
      69505: inst = 32'h8c50000;
      69506: inst = 32'h24612800;
      69507: inst = 32'h10a0ffff;
      69508: inst = 32'hca0fff9;
      69509: inst = 32'h24822800;
      69510: inst = 32'h10a00000;
      69511: inst = 32'hca00004;
      69512: inst = 32'h38632800;
      69513: inst = 32'h38842800;
      69514: inst = 32'h10a00001;
      69515: inst = 32'hca00f8f;
      69516: inst = 32'h13e00001;
      69517: inst = 32'hfe0d96a;
      69518: inst = 32'h5be00000;
      69519: inst = 32'h8c50000;
      69520: inst = 32'h24612800;
      69521: inst = 32'h10a0ffff;
      69522: inst = 32'hca0fff9;
      69523: inst = 32'h24822800;
      69524: inst = 32'h10a00000;
      69525: inst = 32'hca00004;
      69526: inst = 32'h38632800;
      69527: inst = 32'h38842800;
      69528: inst = 32'h10a00001;
      69529: inst = 32'hca00f9d;
      69530: inst = 32'h13e00001;
      69531: inst = 32'hfe0d96a;
      69532: inst = 32'h5be00000;
      69533: inst = 32'h8c50000;
      69534: inst = 32'h24612800;
      69535: inst = 32'h10a0ffff;
      69536: inst = 32'hca0fff9;
      69537: inst = 32'h24822800;
      69538: inst = 32'h10a00000;
      69539: inst = 32'hca00004;
      69540: inst = 32'h38632800;
      69541: inst = 32'h38842800;
      69542: inst = 32'h10a00001;
      69543: inst = 32'hca00fab;
      69544: inst = 32'h13e00001;
      69545: inst = 32'hfe0d96a;
      69546: inst = 32'h5be00000;
      69547: inst = 32'h8c50000;
      69548: inst = 32'h24612800;
      69549: inst = 32'h10a0ffff;
      69550: inst = 32'hca0fff9;
      69551: inst = 32'h24822800;
      69552: inst = 32'h10a00000;
      69553: inst = 32'hca00004;
      69554: inst = 32'h38632800;
      69555: inst = 32'h38842800;
      69556: inst = 32'h10a00001;
      69557: inst = 32'hca00fb9;
      69558: inst = 32'h13e00001;
      69559: inst = 32'hfe0d96a;
      69560: inst = 32'h5be00000;
      69561: inst = 32'h8c50000;
      69562: inst = 32'h24612800;
      69563: inst = 32'h10a0ffff;
      69564: inst = 32'hca0fff9;
      69565: inst = 32'h24822800;
      69566: inst = 32'h10a00000;
      69567: inst = 32'hca00004;
      69568: inst = 32'h38632800;
      69569: inst = 32'h38842800;
      69570: inst = 32'h10a00001;
      69571: inst = 32'hca00fc7;
      69572: inst = 32'h13e00001;
      69573: inst = 32'hfe0d96a;
      69574: inst = 32'h5be00000;
      69575: inst = 32'h8c50000;
      69576: inst = 32'h24612800;
      69577: inst = 32'h10a0ffff;
      69578: inst = 32'hca0fff9;
      69579: inst = 32'h24822800;
      69580: inst = 32'h10a00000;
      69581: inst = 32'hca00004;
      69582: inst = 32'h38632800;
      69583: inst = 32'h38842800;
      69584: inst = 32'h10a00001;
      69585: inst = 32'hca00fd5;
      69586: inst = 32'h13e00001;
      69587: inst = 32'hfe0d96a;
      69588: inst = 32'h5be00000;
      69589: inst = 32'h8c50000;
      69590: inst = 32'h24612800;
      69591: inst = 32'h10a0ffff;
      69592: inst = 32'hca0fff9;
      69593: inst = 32'h24822800;
      69594: inst = 32'h10a00000;
      69595: inst = 32'hca00004;
      69596: inst = 32'h38632800;
      69597: inst = 32'h38842800;
      69598: inst = 32'h10a00001;
      69599: inst = 32'hca00fe3;
      69600: inst = 32'h13e00001;
      69601: inst = 32'hfe0d96a;
      69602: inst = 32'h5be00000;
      69603: inst = 32'h8c50000;
      69604: inst = 32'h24612800;
      69605: inst = 32'h10a0ffff;
      69606: inst = 32'hca0fff9;
      69607: inst = 32'h24822800;
      69608: inst = 32'h10a00000;
      69609: inst = 32'hca00004;
      69610: inst = 32'h38632800;
      69611: inst = 32'h38842800;
      69612: inst = 32'h10a00001;
      69613: inst = 32'hca00ff1;
      69614: inst = 32'h13e00001;
      69615: inst = 32'hfe0d96a;
      69616: inst = 32'h5be00000;
      69617: inst = 32'h8c50000;
      69618: inst = 32'h24612800;
      69619: inst = 32'h10a0ffff;
      69620: inst = 32'hca0fff9;
      69621: inst = 32'h24822800;
      69622: inst = 32'h10a00000;
      69623: inst = 32'hca00004;
      69624: inst = 32'h38632800;
      69625: inst = 32'h38842800;
      69626: inst = 32'h10a00001;
      69627: inst = 32'hca00fff;
      69628: inst = 32'h13e00001;
      69629: inst = 32'hfe0d96a;
      69630: inst = 32'h5be00000;
      69631: inst = 32'h8c50000;
      69632: inst = 32'h24612800;
      69633: inst = 32'h10a0ffff;
      69634: inst = 32'hca0fff9;
      69635: inst = 32'h24822800;
      69636: inst = 32'h10a00000;
      69637: inst = 32'hca00004;
      69638: inst = 32'h38632800;
      69639: inst = 32'h38842800;
      69640: inst = 32'h10a00001;
      69641: inst = 32'hca0100d;
      69642: inst = 32'h13e00001;
      69643: inst = 32'hfe0d96a;
      69644: inst = 32'h5be00000;
      69645: inst = 32'h8c50000;
      69646: inst = 32'h24612800;
      69647: inst = 32'h10a0ffff;
      69648: inst = 32'hca0fff9;
      69649: inst = 32'h24822800;
      69650: inst = 32'h10a00000;
      69651: inst = 32'hca00004;
      69652: inst = 32'h38632800;
      69653: inst = 32'h38842800;
      69654: inst = 32'h10a00001;
      69655: inst = 32'hca0101b;
      69656: inst = 32'h13e00001;
      69657: inst = 32'hfe0d96a;
      69658: inst = 32'h5be00000;
      69659: inst = 32'h8c50000;
      69660: inst = 32'h24612800;
      69661: inst = 32'h10a0ffff;
      69662: inst = 32'hca0fff9;
      69663: inst = 32'h24822800;
      69664: inst = 32'h10a00000;
      69665: inst = 32'hca00004;
      69666: inst = 32'h38632800;
      69667: inst = 32'h38842800;
      69668: inst = 32'h10a00001;
      69669: inst = 32'hca01029;
      69670: inst = 32'h13e00001;
      69671: inst = 32'hfe0d96a;
      69672: inst = 32'h5be00000;
      69673: inst = 32'h8c50000;
      69674: inst = 32'h24612800;
      69675: inst = 32'h10a0ffff;
      69676: inst = 32'hca0fff9;
      69677: inst = 32'h24822800;
      69678: inst = 32'h10a00000;
      69679: inst = 32'hca00004;
      69680: inst = 32'h38632800;
      69681: inst = 32'h38842800;
      69682: inst = 32'h10a00001;
      69683: inst = 32'hca01037;
      69684: inst = 32'h13e00001;
      69685: inst = 32'hfe0d96a;
      69686: inst = 32'h5be00000;
      69687: inst = 32'h8c50000;
      69688: inst = 32'h24612800;
      69689: inst = 32'h10a0ffff;
      69690: inst = 32'hca0fff9;
      69691: inst = 32'h24822800;
      69692: inst = 32'h10a00000;
      69693: inst = 32'hca00004;
      69694: inst = 32'h38632800;
      69695: inst = 32'h38842800;
      69696: inst = 32'h10a00001;
      69697: inst = 32'hca01045;
      69698: inst = 32'h13e00001;
      69699: inst = 32'hfe0d96a;
      69700: inst = 32'h5be00000;
      69701: inst = 32'h8c50000;
      69702: inst = 32'h24612800;
      69703: inst = 32'h10a0ffff;
      69704: inst = 32'hca0fff9;
      69705: inst = 32'h24822800;
      69706: inst = 32'h10a00000;
      69707: inst = 32'hca00004;
      69708: inst = 32'h38632800;
      69709: inst = 32'h38842800;
      69710: inst = 32'h10a00001;
      69711: inst = 32'hca01053;
      69712: inst = 32'h13e00001;
      69713: inst = 32'hfe0d96a;
      69714: inst = 32'h5be00000;
      69715: inst = 32'h8c50000;
      69716: inst = 32'h24612800;
      69717: inst = 32'h10a0ffff;
      69718: inst = 32'hca0fff9;
      69719: inst = 32'h24822800;
      69720: inst = 32'h10a00000;
      69721: inst = 32'hca00004;
      69722: inst = 32'h38632800;
      69723: inst = 32'h38842800;
      69724: inst = 32'h10a00001;
      69725: inst = 32'hca01061;
      69726: inst = 32'h13e00001;
      69727: inst = 32'hfe0d96a;
      69728: inst = 32'h5be00000;
      69729: inst = 32'h8c50000;
      69730: inst = 32'h24612800;
      69731: inst = 32'h10a0ffff;
      69732: inst = 32'hca0fff9;
      69733: inst = 32'h24822800;
      69734: inst = 32'h10a00000;
      69735: inst = 32'hca00004;
      69736: inst = 32'h38632800;
      69737: inst = 32'h38842800;
      69738: inst = 32'h10a00001;
      69739: inst = 32'hca0106f;
      69740: inst = 32'h13e00001;
      69741: inst = 32'hfe0d96a;
      69742: inst = 32'h5be00000;
      69743: inst = 32'h8c50000;
      69744: inst = 32'h24612800;
      69745: inst = 32'h10a0ffff;
      69746: inst = 32'hca0fff9;
      69747: inst = 32'h24822800;
      69748: inst = 32'h10a00000;
      69749: inst = 32'hca00004;
      69750: inst = 32'h38632800;
      69751: inst = 32'h38842800;
      69752: inst = 32'h10a00001;
      69753: inst = 32'hca0107d;
      69754: inst = 32'h13e00001;
      69755: inst = 32'hfe0d96a;
      69756: inst = 32'h5be00000;
      69757: inst = 32'h8c50000;
      69758: inst = 32'h24612800;
      69759: inst = 32'h10a0ffff;
      69760: inst = 32'hca0fff9;
      69761: inst = 32'h24822800;
      69762: inst = 32'h10a00000;
      69763: inst = 32'hca00004;
      69764: inst = 32'h38632800;
      69765: inst = 32'h38842800;
      69766: inst = 32'h10a00001;
      69767: inst = 32'hca0108b;
      69768: inst = 32'h13e00001;
      69769: inst = 32'hfe0d96a;
      69770: inst = 32'h5be00000;
      69771: inst = 32'h8c50000;
      69772: inst = 32'h24612800;
      69773: inst = 32'h10a0ffff;
      69774: inst = 32'hca0fff9;
      69775: inst = 32'h24822800;
      69776: inst = 32'h10a00000;
      69777: inst = 32'hca00004;
      69778: inst = 32'h38632800;
      69779: inst = 32'h38842800;
      69780: inst = 32'h10a00001;
      69781: inst = 32'hca01099;
      69782: inst = 32'h13e00001;
      69783: inst = 32'hfe0d96a;
      69784: inst = 32'h5be00000;
      69785: inst = 32'h8c50000;
      69786: inst = 32'h24612800;
      69787: inst = 32'h10a0ffff;
      69788: inst = 32'hca0fff9;
      69789: inst = 32'h24822800;
      69790: inst = 32'h10a00000;
      69791: inst = 32'hca00004;
      69792: inst = 32'h38632800;
      69793: inst = 32'h38842800;
      69794: inst = 32'h10a00001;
      69795: inst = 32'hca010a7;
      69796: inst = 32'h13e00001;
      69797: inst = 32'hfe0d96a;
      69798: inst = 32'h5be00000;
      69799: inst = 32'h8c50000;
      69800: inst = 32'h24612800;
      69801: inst = 32'h10a0ffff;
      69802: inst = 32'hca0fff9;
      69803: inst = 32'h24822800;
      69804: inst = 32'h10a00000;
      69805: inst = 32'hca00004;
      69806: inst = 32'h38632800;
      69807: inst = 32'h38842800;
      69808: inst = 32'h10a00001;
      69809: inst = 32'hca010b5;
      69810: inst = 32'h13e00001;
      69811: inst = 32'hfe0d96a;
      69812: inst = 32'h5be00000;
      69813: inst = 32'h8c50000;
      69814: inst = 32'h24612800;
      69815: inst = 32'h10a0ffff;
      69816: inst = 32'hca0fff9;
      69817: inst = 32'h24822800;
      69818: inst = 32'h10a00000;
      69819: inst = 32'hca00004;
      69820: inst = 32'h38632800;
      69821: inst = 32'h38842800;
      69822: inst = 32'h10a00001;
      69823: inst = 32'hca010c3;
      69824: inst = 32'h13e00001;
      69825: inst = 32'hfe0d96a;
      69826: inst = 32'h5be00000;
      69827: inst = 32'h8c50000;
      69828: inst = 32'h24612800;
      69829: inst = 32'h10a0ffff;
      69830: inst = 32'hca0fff9;
      69831: inst = 32'h24822800;
      69832: inst = 32'h10a00000;
      69833: inst = 32'hca00004;
      69834: inst = 32'h38632800;
      69835: inst = 32'h38842800;
      69836: inst = 32'h10a00001;
      69837: inst = 32'hca010d1;
      69838: inst = 32'h13e00001;
      69839: inst = 32'hfe0d96a;
      69840: inst = 32'h5be00000;
      69841: inst = 32'h8c50000;
      69842: inst = 32'h24612800;
      69843: inst = 32'h10a0ffff;
      69844: inst = 32'hca0fff9;
      69845: inst = 32'h24822800;
      69846: inst = 32'h10a00000;
      69847: inst = 32'hca00004;
      69848: inst = 32'h38632800;
      69849: inst = 32'h38842800;
      69850: inst = 32'h10a00001;
      69851: inst = 32'hca010df;
      69852: inst = 32'h13e00001;
      69853: inst = 32'hfe0d96a;
      69854: inst = 32'h5be00000;
      69855: inst = 32'h8c50000;
      69856: inst = 32'h24612800;
      69857: inst = 32'h10a0ffff;
      69858: inst = 32'hca0fff9;
      69859: inst = 32'h24822800;
      69860: inst = 32'h10a00000;
      69861: inst = 32'hca00004;
      69862: inst = 32'h38632800;
      69863: inst = 32'h38842800;
      69864: inst = 32'h10a00001;
      69865: inst = 32'hca010ed;
      69866: inst = 32'h13e00001;
      69867: inst = 32'hfe0d96a;
      69868: inst = 32'h5be00000;
      69869: inst = 32'h8c50000;
      69870: inst = 32'h24612800;
      69871: inst = 32'h10a0ffff;
      69872: inst = 32'hca0fff9;
      69873: inst = 32'h24822800;
      69874: inst = 32'h10a00000;
      69875: inst = 32'hca00004;
      69876: inst = 32'h38632800;
      69877: inst = 32'h38842800;
      69878: inst = 32'h10a00001;
      69879: inst = 32'hca010fb;
      69880: inst = 32'h13e00001;
      69881: inst = 32'hfe0d96a;
      69882: inst = 32'h5be00000;
      69883: inst = 32'h8c50000;
      69884: inst = 32'h24612800;
      69885: inst = 32'h10a0ffff;
      69886: inst = 32'hca0fff9;
      69887: inst = 32'h24822800;
      69888: inst = 32'h10a00000;
      69889: inst = 32'hca00004;
      69890: inst = 32'h38632800;
      69891: inst = 32'h38842800;
      69892: inst = 32'h10a00001;
      69893: inst = 32'hca01109;
      69894: inst = 32'h13e00001;
      69895: inst = 32'hfe0d96a;
      69896: inst = 32'h5be00000;
      69897: inst = 32'h8c50000;
      69898: inst = 32'h24612800;
      69899: inst = 32'h10a0ffff;
      69900: inst = 32'hca0fff9;
      69901: inst = 32'h24822800;
      69902: inst = 32'h10a00000;
      69903: inst = 32'hca00004;
      69904: inst = 32'h38632800;
      69905: inst = 32'h38842800;
      69906: inst = 32'h10a00001;
      69907: inst = 32'hca01117;
      69908: inst = 32'h13e00001;
      69909: inst = 32'hfe0d96a;
      69910: inst = 32'h5be00000;
      69911: inst = 32'h8c50000;
      69912: inst = 32'h24612800;
      69913: inst = 32'h10a0ffff;
      69914: inst = 32'hca0fff9;
      69915: inst = 32'h24822800;
      69916: inst = 32'h10a00000;
      69917: inst = 32'hca00004;
      69918: inst = 32'h38632800;
      69919: inst = 32'h38842800;
      69920: inst = 32'h10a00001;
      69921: inst = 32'hca01125;
      69922: inst = 32'h13e00001;
      69923: inst = 32'hfe0d96a;
      69924: inst = 32'h5be00000;
      69925: inst = 32'h8c50000;
      69926: inst = 32'h24612800;
      69927: inst = 32'h10a0ffff;
      69928: inst = 32'hca0fff9;
      69929: inst = 32'h24822800;
      69930: inst = 32'h10a00000;
      69931: inst = 32'hca00004;
      69932: inst = 32'h38632800;
      69933: inst = 32'h38842800;
      69934: inst = 32'h10a00001;
      69935: inst = 32'hca01133;
      69936: inst = 32'h13e00001;
      69937: inst = 32'hfe0d96a;
      69938: inst = 32'h5be00000;
      69939: inst = 32'h8c50000;
      69940: inst = 32'h24612800;
      69941: inst = 32'h10a0ffff;
      69942: inst = 32'hca0fff9;
      69943: inst = 32'h24822800;
      69944: inst = 32'h10a00000;
      69945: inst = 32'hca00004;
      69946: inst = 32'h38632800;
      69947: inst = 32'h38842800;
      69948: inst = 32'h10a00001;
      69949: inst = 32'hca01141;
      69950: inst = 32'h13e00001;
      69951: inst = 32'hfe0d96a;
      69952: inst = 32'h5be00000;
      69953: inst = 32'h8c50000;
      69954: inst = 32'h24612800;
      69955: inst = 32'h10a0ffff;
      69956: inst = 32'hca0fff9;
      69957: inst = 32'h24822800;
      69958: inst = 32'h10a00000;
      69959: inst = 32'hca00004;
      69960: inst = 32'h38632800;
      69961: inst = 32'h38842800;
      69962: inst = 32'h10a00001;
      69963: inst = 32'hca0114f;
      69964: inst = 32'h13e00001;
      69965: inst = 32'hfe0d96a;
      69966: inst = 32'h5be00000;
      69967: inst = 32'h8c50000;
      69968: inst = 32'h24612800;
      69969: inst = 32'h10a0ffff;
      69970: inst = 32'hca0fff9;
      69971: inst = 32'h24822800;
      69972: inst = 32'h10a00000;
      69973: inst = 32'hca00004;
      69974: inst = 32'h38632800;
      69975: inst = 32'h38842800;
      69976: inst = 32'h10a00001;
      69977: inst = 32'hca0115d;
      69978: inst = 32'h13e00001;
      69979: inst = 32'hfe0d96a;
      69980: inst = 32'h5be00000;
      69981: inst = 32'h8c50000;
      69982: inst = 32'h24612800;
      69983: inst = 32'h10a0ffff;
      69984: inst = 32'hca0fff9;
      69985: inst = 32'h24822800;
      69986: inst = 32'h10a00000;
      69987: inst = 32'hca00004;
      69988: inst = 32'h38632800;
      69989: inst = 32'h38842800;
      69990: inst = 32'h10a00001;
      69991: inst = 32'hca0116b;
      69992: inst = 32'h13e00001;
      69993: inst = 32'hfe0d96a;
      69994: inst = 32'h5be00000;
      69995: inst = 32'h8c50000;
      69996: inst = 32'h24612800;
      69997: inst = 32'h10a0ffff;
      69998: inst = 32'hca0fff9;
      69999: inst = 32'h24822800;
      70000: inst = 32'h10a00000;
      70001: inst = 32'hca00004;
      70002: inst = 32'h38632800;
      70003: inst = 32'h38842800;
      70004: inst = 32'h10a00001;
      70005: inst = 32'hca01179;
      70006: inst = 32'h13e00001;
      70007: inst = 32'hfe0d96a;
      70008: inst = 32'h5be00000;
      70009: inst = 32'h8c50000;
      70010: inst = 32'h24612800;
      70011: inst = 32'h10a0ffff;
      70012: inst = 32'hca0fff9;
      70013: inst = 32'h24822800;
      70014: inst = 32'h10a00000;
      70015: inst = 32'hca00004;
      70016: inst = 32'h38632800;
      70017: inst = 32'h38842800;
      70018: inst = 32'h10a00001;
      70019: inst = 32'hca01187;
      70020: inst = 32'h13e00001;
      70021: inst = 32'hfe0d96a;
      70022: inst = 32'h5be00000;
      70023: inst = 32'h8c50000;
      70024: inst = 32'h24612800;
      70025: inst = 32'h10a0ffff;
      70026: inst = 32'hca0fff9;
      70027: inst = 32'h24822800;
      70028: inst = 32'h10a00000;
      70029: inst = 32'hca00004;
      70030: inst = 32'h38632800;
      70031: inst = 32'h38842800;
      70032: inst = 32'h10a00001;
      70033: inst = 32'hca01195;
      70034: inst = 32'h13e00001;
      70035: inst = 32'hfe0d96a;
      70036: inst = 32'h5be00000;
      70037: inst = 32'h8c50000;
      70038: inst = 32'h24612800;
      70039: inst = 32'h10a0ffff;
      70040: inst = 32'hca0fff9;
      70041: inst = 32'h24822800;
      70042: inst = 32'h10a00000;
      70043: inst = 32'hca00004;
      70044: inst = 32'h38632800;
      70045: inst = 32'h38842800;
      70046: inst = 32'h10a00001;
      70047: inst = 32'hca011a3;
      70048: inst = 32'h13e00001;
      70049: inst = 32'hfe0d96a;
      70050: inst = 32'h5be00000;
      70051: inst = 32'h8c50000;
      70052: inst = 32'h24612800;
      70053: inst = 32'h10a0ffff;
      70054: inst = 32'hca0fff9;
      70055: inst = 32'h24822800;
      70056: inst = 32'h10a00000;
      70057: inst = 32'hca00004;
      70058: inst = 32'h38632800;
      70059: inst = 32'h38842800;
      70060: inst = 32'h10a00001;
      70061: inst = 32'hca011b1;
      70062: inst = 32'h13e00001;
      70063: inst = 32'hfe0d96a;
      70064: inst = 32'h5be00000;
      70065: inst = 32'h8c50000;
      70066: inst = 32'h24612800;
      70067: inst = 32'h10a0ffff;
      70068: inst = 32'hca0fff9;
      70069: inst = 32'h24822800;
      70070: inst = 32'h10a00000;
      70071: inst = 32'hca00004;
      70072: inst = 32'h38632800;
      70073: inst = 32'h38842800;
      70074: inst = 32'h10a00001;
      70075: inst = 32'hca011bf;
      70076: inst = 32'h13e00001;
      70077: inst = 32'hfe0d96a;
      70078: inst = 32'h5be00000;
      70079: inst = 32'h8c50000;
      70080: inst = 32'h24612800;
      70081: inst = 32'h10a0ffff;
      70082: inst = 32'hca0fff9;
      70083: inst = 32'h24822800;
      70084: inst = 32'h10a00000;
      70085: inst = 32'hca00004;
      70086: inst = 32'h38632800;
      70087: inst = 32'h38842800;
      70088: inst = 32'h10a00001;
      70089: inst = 32'hca011cd;
      70090: inst = 32'h13e00001;
      70091: inst = 32'hfe0d96a;
      70092: inst = 32'h5be00000;
      70093: inst = 32'h8c50000;
      70094: inst = 32'h24612800;
      70095: inst = 32'h10a0ffff;
      70096: inst = 32'hca0fff9;
      70097: inst = 32'h24822800;
      70098: inst = 32'h10a00000;
      70099: inst = 32'hca00004;
      70100: inst = 32'h38632800;
      70101: inst = 32'h38842800;
      70102: inst = 32'h10a00001;
      70103: inst = 32'hca011db;
      70104: inst = 32'h13e00001;
      70105: inst = 32'hfe0d96a;
      70106: inst = 32'h5be00000;
      70107: inst = 32'h8c50000;
      70108: inst = 32'h24612800;
      70109: inst = 32'h10a0ffff;
      70110: inst = 32'hca0fff9;
      70111: inst = 32'h24822800;
      70112: inst = 32'h10a00000;
      70113: inst = 32'hca00004;
      70114: inst = 32'h38632800;
      70115: inst = 32'h38842800;
      70116: inst = 32'h10a00001;
      70117: inst = 32'hca011e9;
      70118: inst = 32'h13e00001;
      70119: inst = 32'hfe0d96a;
      70120: inst = 32'h5be00000;
      70121: inst = 32'h8c50000;
      70122: inst = 32'h24612800;
      70123: inst = 32'h10a0ffff;
      70124: inst = 32'hca0fffa;
      70125: inst = 32'h24822800;
      70126: inst = 32'h10a00000;
      70127: inst = 32'hca00004;
      70128: inst = 32'h38632800;
      70129: inst = 32'h38842800;
      70130: inst = 32'h10a00001;
      70131: inst = 32'hca011f7;
      70132: inst = 32'h13e00001;
      70133: inst = 32'hfe0d96a;
      70134: inst = 32'h5be00000;
      70135: inst = 32'h8c50000;
      70136: inst = 32'h24612800;
      70137: inst = 32'h10a0ffff;
      70138: inst = 32'hca0fffa;
      70139: inst = 32'h24822800;
      70140: inst = 32'h10a00000;
      70141: inst = 32'hca00004;
      70142: inst = 32'h38632800;
      70143: inst = 32'h38842800;
      70144: inst = 32'h10a00001;
      70145: inst = 32'hca01205;
      70146: inst = 32'h13e00001;
      70147: inst = 32'hfe0d96a;
      70148: inst = 32'h5be00000;
      70149: inst = 32'h8c50000;
      70150: inst = 32'h24612800;
      70151: inst = 32'h10a0ffff;
      70152: inst = 32'hca0fffa;
      70153: inst = 32'h24822800;
      70154: inst = 32'h10a00000;
      70155: inst = 32'hca00004;
      70156: inst = 32'h38632800;
      70157: inst = 32'h38842800;
      70158: inst = 32'h10a00001;
      70159: inst = 32'hca01213;
      70160: inst = 32'h13e00001;
      70161: inst = 32'hfe0d96a;
      70162: inst = 32'h5be00000;
      70163: inst = 32'h8c50000;
      70164: inst = 32'h24612800;
      70165: inst = 32'h10a0ffff;
      70166: inst = 32'hca0fffa;
      70167: inst = 32'h24822800;
      70168: inst = 32'h10a00000;
      70169: inst = 32'hca00004;
      70170: inst = 32'h38632800;
      70171: inst = 32'h38842800;
      70172: inst = 32'h10a00001;
      70173: inst = 32'hca01221;
      70174: inst = 32'h13e00001;
      70175: inst = 32'hfe0d96a;
      70176: inst = 32'h5be00000;
      70177: inst = 32'h8c50000;
      70178: inst = 32'h24612800;
      70179: inst = 32'h10a0ffff;
      70180: inst = 32'hca0fffa;
      70181: inst = 32'h24822800;
      70182: inst = 32'h10a00000;
      70183: inst = 32'hca00004;
      70184: inst = 32'h38632800;
      70185: inst = 32'h38842800;
      70186: inst = 32'h10a00001;
      70187: inst = 32'hca0122f;
      70188: inst = 32'h13e00001;
      70189: inst = 32'hfe0d96a;
      70190: inst = 32'h5be00000;
      70191: inst = 32'h8c50000;
      70192: inst = 32'h24612800;
      70193: inst = 32'h10a0ffff;
      70194: inst = 32'hca0fffa;
      70195: inst = 32'h24822800;
      70196: inst = 32'h10a00000;
      70197: inst = 32'hca00004;
      70198: inst = 32'h38632800;
      70199: inst = 32'h38842800;
      70200: inst = 32'h10a00001;
      70201: inst = 32'hca0123d;
      70202: inst = 32'h13e00001;
      70203: inst = 32'hfe0d96a;
      70204: inst = 32'h5be00000;
      70205: inst = 32'h8c50000;
      70206: inst = 32'h24612800;
      70207: inst = 32'h10a0ffff;
      70208: inst = 32'hca0fffa;
      70209: inst = 32'h24822800;
      70210: inst = 32'h10a00000;
      70211: inst = 32'hca00004;
      70212: inst = 32'h38632800;
      70213: inst = 32'h38842800;
      70214: inst = 32'h10a00001;
      70215: inst = 32'hca0124b;
      70216: inst = 32'h13e00001;
      70217: inst = 32'hfe0d96a;
      70218: inst = 32'h5be00000;
      70219: inst = 32'h8c50000;
      70220: inst = 32'h24612800;
      70221: inst = 32'h10a0ffff;
      70222: inst = 32'hca0fffa;
      70223: inst = 32'h24822800;
      70224: inst = 32'h10a00000;
      70225: inst = 32'hca00004;
      70226: inst = 32'h38632800;
      70227: inst = 32'h38842800;
      70228: inst = 32'h10a00001;
      70229: inst = 32'hca01259;
      70230: inst = 32'h13e00001;
      70231: inst = 32'hfe0d96a;
      70232: inst = 32'h5be00000;
      70233: inst = 32'h8c50000;
      70234: inst = 32'h24612800;
      70235: inst = 32'h10a0ffff;
      70236: inst = 32'hca0fffa;
      70237: inst = 32'h24822800;
      70238: inst = 32'h10a00000;
      70239: inst = 32'hca00004;
      70240: inst = 32'h38632800;
      70241: inst = 32'h38842800;
      70242: inst = 32'h10a00001;
      70243: inst = 32'hca01267;
      70244: inst = 32'h13e00001;
      70245: inst = 32'hfe0d96a;
      70246: inst = 32'h5be00000;
      70247: inst = 32'h8c50000;
      70248: inst = 32'h24612800;
      70249: inst = 32'h10a0ffff;
      70250: inst = 32'hca0fffa;
      70251: inst = 32'h24822800;
      70252: inst = 32'h10a00000;
      70253: inst = 32'hca00004;
      70254: inst = 32'h38632800;
      70255: inst = 32'h38842800;
      70256: inst = 32'h10a00001;
      70257: inst = 32'hca01275;
      70258: inst = 32'h13e00001;
      70259: inst = 32'hfe0d96a;
      70260: inst = 32'h5be00000;
      70261: inst = 32'h8c50000;
      70262: inst = 32'h24612800;
      70263: inst = 32'h10a0ffff;
      70264: inst = 32'hca0fffa;
      70265: inst = 32'h24822800;
      70266: inst = 32'h10a00000;
      70267: inst = 32'hca00004;
      70268: inst = 32'h38632800;
      70269: inst = 32'h38842800;
      70270: inst = 32'h10a00001;
      70271: inst = 32'hca01283;
      70272: inst = 32'h13e00001;
      70273: inst = 32'hfe0d96a;
      70274: inst = 32'h5be00000;
      70275: inst = 32'h8c50000;
      70276: inst = 32'h24612800;
      70277: inst = 32'h10a0ffff;
      70278: inst = 32'hca0fffa;
      70279: inst = 32'h24822800;
      70280: inst = 32'h10a00000;
      70281: inst = 32'hca00004;
      70282: inst = 32'h38632800;
      70283: inst = 32'h38842800;
      70284: inst = 32'h10a00001;
      70285: inst = 32'hca01291;
      70286: inst = 32'h13e00001;
      70287: inst = 32'hfe0d96a;
      70288: inst = 32'h5be00000;
      70289: inst = 32'h8c50000;
      70290: inst = 32'h24612800;
      70291: inst = 32'h10a0ffff;
      70292: inst = 32'hca0fffa;
      70293: inst = 32'h24822800;
      70294: inst = 32'h10a00000;
      70295: inst = 32'hca00004;
      70296: inst = 32'h38632800;
      70297: inst = 32'h38842800;
      70298: inst = 32'h10a00001;
      70299: inst = 32'hca0129f;
      70300: inst = 32'h13e00001;
      70301: inst = 32'hfe0d96a;
      70302: inst = 32'h5be00000;
      70303: inst = 32'h8c50000;
      70304: inst = 32'h24612800;
      70305: inst = 32'h10a0ffff;
      70306: inst = 32'hca0fffa;
      70307: inst = 32'h24822800;
      70308: inst = 32'h10a00000;
      70309: inst = 32'hca00004;
      70310: inst = 32'h38632800;
      70311: inst = 32'h38842800;
      70312: inst = 32'h10a00001;
      70313: inst = 32'hca012ad;
      70314: inst = 32'h13e00001;
      70315: inst = 32'hfe0d96a;
      70316: inst = 32'h5be00000;
      70317: inst = 32'h8c50000;
      70318: inst = 32'h24612800;
      70319: inst = 32'h10a0ffff;
      70320: inst = 32'hca0fffa;
      70321: inst = 32'h24822800;
      70322: inst = 32'h10a00000;
      70323: inst = 32'hca00004;
      70324: inst = 32'h38632800;
      70325: inst = 32'h38842800;
      70326: inst = 32'h10a00001;
      70327: inst = 32'hca012bb;
      70328: inst = 32'h13e00001;
      70329: inst = 32'hfe0d96a;
      70330: inst = 32'h5be00000;
      70331: inst = 32'h8c50000;
      70332: inst = 32'h24612800;
      70333: inst = 32'h10a0ffff;
      70334: inst = 32'hca0fffa;
      70335: inst = 32'h24822800;
      70336: inst = 32'h10a00000;
      70337: inst = 32'hca00004;
      70338: inst = 32'h38632800;
      70339: inst = 32'h38842800;
      70340: inst = 32'h10a00001;
      70341: inst = 32'hca012c9;
      70342: inst = 32'h13e00001;
      70343: inst = 32'hfe0d96a;
      70344: inst = 32'h5be00000;
      70345: inst = 32'h8c50000;
      70346: inst = 32'h24612800;
      70347: inst = 32'h10a0ffff;
      70348: inst = 32'hca0fffa;
      70349: inst = 32'h24822800;
      70350: inst = 32'h10a00000;
      70351: inst = 32'hca00004;
      70352: inst = 32'h38632800;
      70353: inst = 32'h38842800;
      70354: inst = 32'h10a00001;
      70355: inst = 32'hca012d7;
      70356: inst = 32'h13e00001;
      70357: inst = 32'hfe0d96a;
      70358: inst = 32'h5be00000;
      70359: inst = 32'h8c50000;
      70360: inst = 32'h24612800;
      70361: inst = 32'h10a0ffff;
      70362: inst = 32'hca0fffa;
      70363: inst = 32'h24822800;
      70364: inst = 32'h10a00000;
      70365: inst = 32'hca00004;
      70366: inst = 32'h38632800;
      70367: inst = 32'h38842800;
      70368: inst = 32'h10a00001;
      70369: inst = 32'hca012e5;
      70370: inst = 32'h13e00001;
      70371: inst = 32'hfe0d96a;
      70372: inst = 32'h5be00000;
      70373: inst = 32'h8c50000;
      70374: inst = 32'h24612800;
      70375: inst = 32'h10a0ffff;
      70376: inst = 32'hca0fffa;
      70377: inst = 32'h24822800;
      70378: inst = 32'h10a00000;
      70379: inst = 32'hca00004;
      70380: inst = 32'h38632800;
      70381: inst = 32'h38842800;
      70382: inst = 32'h10a00001;
      70383: inst = 32'hca012f3;
      70384: inst = 32'h13e00001;
      70385: inst = 32'hfe0d96a;
      70386: inst = 32'h5be00000;
      70387: inst = 32'h8c50000;
      70388: inst = 32'h24612800;
      70389: inst = 32'h10a0ffff;
      70390: inst = 32'hca0fffa;
      70391: inst = 32'h24822800;
      70392: inst = 32'h10a00000;
      70393: inst = 32'hca00004;
      70394: inst = 32'h38632800;
      70395: inst = 32'h38842800;
      70396: inst = 32'h10a00001;
      70397: inst = 32'hca01301;
      70398: inst = 32'h13e00001;
      70399: inst = 32'hfe0d96a;
      70400: inst = 32'h5be00000;
      70401: inst = 32'h8c50000;
      70402: inst = 32'h24612800;
      70403: inst = 32'h10a0ffff;
      70404: inst = 32'hca0fffa;
      70405: inst = 32'h24822800;
      70406: inst = 32'h10a00000;
      70407: inst = 32'hca00004;
      70408: inst = 32'h38632800;
      70409: inst = 32'h38842800;
      70410: inst = 32'h10a00001;
      70411: inst = 32'hca0130f;
      70412: inst = 32'h13e00001;
      70413: inst = 32'hfe0d96a;
      70414: inst = 32'h5be00000;
      70415: inst = 32'h8c50000;
      70416: inst = 32'h24612800;
      70417: inst = 32'h10a0ffff;
      70418: inst = 32'hca0fffa;
      70419: inst = 32'h24822800;
      70420: inst = 32'h10a00000;
      70421: inst = 32'hca00004;
      70422: inst = 32'h38632800;
      70423: inst = 32'h38842800;
      70424: inst = 32'h10a00001;
      70425: inst = 32'hca0131d;
      70426: inst = 32'h13e00001;
      70427: inst = 32'hfe0d96a;
      70428: inst = 32'h5be00000;
      70429: inst = 32'h8c50000;
      70430: inst = 32'h24612800;
      70431: inst = 32'h10a0ffff;
      70432: inst = 32'hca0fffa;
      70433: inst = 32'h24822800;
      70434: inst = 32'h10a00000;
      70435: inst = 32'hca00004;
      70436: inst = 32'h38632800;
      70437: inst = 32'h38842800;
      70438: inst = 32'h10a00001;
      70439: inst = 32'hca0132b;
      70440: inst = 32'h13e00001;
      70441: inst = 32'hfe0d96a;
      70442: inst = 32'h5be00000;
      70443: inst = 32'h8c50000;
      70444: inst = 32'h24612800;
      70445: inst = 32'h10a0ffff;
      70446: inst = 32'hca0fffa;
      70447: inst = 32'h24822800;
      70448: inst = 32'h10a00000;
      70449: inst = 32'hca00004;
      70450: inst = 32'h38632800;
      70451: inst = 32'h38842800;
      70452: inst = 32'h10a00001;
      70453: inst = 32'hca01339;
      70454: inst = 32'h13e00001;
      70455: inst = 32'hfe0d96a;
      70456: inst = 32'h5be00000;
      70457: inst = 32'h8c50000;
      70458: inst = 32'h24612800;
      70459: inst = 32'h10a0ffff;
      70460: inst = 32'hca0fffa;
      70461: inst = 32'h24822800;
      70462: inst = 32'h10a00000;
      70463: inst = 32'hca00004;
      70464: inst = 32'h38632800;
      70465: inst = 32'h38842800;
      70466: inst = 32'h10a00001;
      70467: inst = 32'hca01347;
      70468: inst = 32'h13e00001;
      70469: inst = 32'hfe0d96a;
      70470: inst = 32'h5be00000;
      70471: inst = 32'h8c50000;
      70472: inst = 32'h24612800;
      70473: inst = 32'h10a0ffff;
      70474: inst = 32'hca0fffa;
      70475: inst = 32'h24822800;
      70476: inst = 32'h10a00000;
      70477: inst = 32'hca00004;
      70478: inst = 32'h38632800;
      70479: inst = 32'h38842800;
      70480: inst = 32'h10a00001;
      70481: inst = 32'hca01355;
      70482: inst = 32'h13e00001;
      70483: inst = 32'hfe0d96a;
      70484: inst = 32'h5be00000;
      70485: inst = 32'h8c50000;
      70486: inst = 32'h24612800;
      70487: inst = 32'h10a0ffff;
      70488: inst = 32'hca0fffa;
      70489: inst = 32'h24822800;
      70490: inst = 32'h10a00000;
      70491: inst = 32'hca00004;
      70492: inst = 32'h38632800;
      70493: inst = 32'h38842800;
      70494: inst = 32'h10a00001;
      70495: inst = 32'hca01363;
      70496: inst = 32'h13e00001;
      70497: inst = 32'hfe0d96a;
      70498: inst = 32'h5be00000;
      70499: inst = 32'h8c50000;
      70500: inst = 32'h24612800;
      70501: inst = 32'h10a0ffff;
      70502: inst = 32'hca0fffa;
      70503: inst = 32'h24822800;
      70504: inst = 32'h10a00000;
      70505: inst = 32'hca00004;
      70506: inst = 32'h38632800;
      70507: inst = 32'h38842800;
      70508: inst = 32'h10a00001;
      70509: inst = 32'hca01371;
      70510: inst = 32'h13e00001;
      70511: inst = 32'hfe0d96a;
      70512: inst = 32'h5be00000;
      70513: inst = 32'h8c50000;
      70514: inst = 32'h24612800;
      70515: inst = 32'h10a0ffff;
      70516: inst = 32'hca0fffa;
      70517: inst = 32'h24822800;
      70518: inst = 32'h10a00000;
      70519: inst = 32'hca00004;
      70520: inst = 32'h38632800;
      70521: inst = 32'h38842800;
      70522: inst = 32'h10a00001;
      70523: inst = 32'hca0137f;
      70524: inst = 32'h13e00001;
      70525: inst = 32'hfe0d96a;
      70526: inst = 32'h5be00000;
      70527: inst = 32'h8c50000;
      70528: inst = 32'h24612800;
      70529: inst = 32'h10a0ffff;
      70530: inst = 32'hca0fffa;
      70531: inst = 32'h24822800;
      70532: inst = 32'h10a00000;
      70533: inst = 32'hca00004;
      70534: inst = 32'h38632800;
      70535: inst = 32'h38842800;
      70536: inst = 32'h10a00001;
      70537: inst = 32'hca0138d;
      70538: inst = 32'h13e00001;
      70539: inst = 32'hfe0d96a;
      70540: inst = 32'h5be00000;
      70541: inst = 32'h8c50000;
      70542: inst = 32'h24612800;
      70543: inst = 32'h10a0ffff;
      70544: inst = 32'hca0fffa;
      70545: inst = 32'h24822800;
      70546: inst = 32'h10a00000;
      70547: inst = 32'hca00004;
      70548: inst = 32'h38632800;
      70549: inst = 32'h38842800;
      70550: inst = 32'h10a00001;
      70551: inst = 32'hca0139b;
      70552: inst = 32'h13e00001;
      70553: inst = 32'hfe0d96a;
      70554: inst = 32'h5be00000;
      70555: inst = 32'h8c50000;
      70556: inst = 32'h24612800;
      70557: inst = 32'h10a0ffff;
      70558: inst = 32'hca0fffa;
      70559: inst = 32'h24822800;
      70560: inst = 32'h10a00000;
      70561: inst = 32'hca00004;
      70562: inst = 32'h38632800;
      70563: inst = 32'h38842800;
      70564: inst = 32'h10a00001;
      70565: inst = 32'hca013a9;
      70566: inst = 32'h13e00001;
      70567: inst = 32'hfe0d96a;
      70568: inst = 32'h5be00000;
      70569: inst = 32'h8c50000;
      70570: inst = 32'h24612800;
      70571: inst = 32'h10a0ffff;
      70572: inst = 32'hca0fffa;
      70573: inst = 32'h24822800;
      70574: inst = 32'h10a00000;
      70575: inst = 32'hca00004;
      70576: inst = 32'h38632800;
      70577: inst = 32'h38842800;
      70578: inst = 32'h10a00001;
      70579: inst = 32'hca013b7;
      70580: inst = 32'h13e00001;
      70581: inst = 32'hfe0d96a;
      70582: inst = 32'h5be00000;
      70583: inst = 32'h8c50000;
      70584: inst = 32'h24612800;
      70585: inst = 32'h10a0ffff;
      70586: inst = 32'hca0fffa;
      70587: inst = 32'h24822800;
      70588: inst = 32'h10a00000;
      70589: inst = 32'hca00004;
      70590: inst = 32'h38632800;
      70591: inst = 32'h38842800;
      70592: inst = 32'h10a00001;
      70593: inst = 32'hca013c5;
      70594: inst = 32'h13e00001;
      70595: inst = 32'hfe0d96a;
      70596: inst = 32'h5be00000;
      70597: inst = 32'h8c50000;
      70598: inst = 32'h24612800;
      70599: inst = 32'h10a0ffff;
      70600: inst = 32'hca0fffa;
      70601: inst = 32'h24822800;
      70602: inst = 32'h10a00000;
      70603: inst = 32'hca00004;
      70604: inst = 32'h38632800;
      70605: inst = 32'h38842800;
      70606: inst = 32'h10a00001;
      70607: inst = 32'hca013d3;
      70608: inst = 32'h13e00001;
      70609: inst = 32'hfe0d96a;
      70610: inst = 32'h5be00000;
      70611: inst = 32'h8c50000;
      70612: inst = 32'h24612800;
      70613: inst = 32'h10a0ffff;
      70614: inst = 32'hca0fffa;
      70615: inst = 32'h24822800;
      70616: inst = 32'h10a00000;
      70617: inst = 32'hca00004;
      70618: inst = 32'h38632800;
      70619: inst = 32'h38842800;
      70620: inst = 32'h10a00001;
      70621: inst = 32'hca013e1;
      70622: inst = 32'h13e00001;
      70623: inst = 32'hfe0d96a;
      70624: inst = 32'h5be00000;
      70625: inst = 32'h8c50000;
      70626: inst = 32'h24612800;
      70627: inst = 32'h10a0ffff;
      70628: inst = 32'hca0fffa;
      70629: inst = 32'h24822800;
      70630: inst = 32'h10a00000;
      70631: inst = 32'hca00004;
      70632: inst = 32'h38632800;
      70633: inst = 32'h38842800;
      70634: inst = 32'h10a00001;
      70635: inst = 32'hca013ef;
      70636: inst = 32'h13e00001;
      70637: inst = 32'hfe0d96a;
      70638: inst = 32'h5be00000;
      70639: inst = 32'h8c50000;
      70640: inst = 32'h24612800;
      70641: inst = 32'h10a0ffff;
      70642: inst = 32'hca0fffa;
      70643: inst = 32'h24822800;
      70644: inst = 32'h10a00000;
      70645: inst = 32'hca00004;
      70646: inst = 32'h38632800;
      70647: inst = 32'h38842800;
      70648: inst = 32'h10a00001;
      70649: inst = 32'hca013fd;
      70650: inst = 32'h13e00001;
      70651: inst = 32'hfe0d96a;
      70652: inst = 32'h5be00000;
      70653: inst = 32'h8c50000;
      70654: inst = 32'h24612800;
      70655: inst = 32'h10a0ffff;
      70656: inst = 32'hca0fffa;
      70657: inst = 32'h24822800;
      70658: inst = 32'h10a00000;
      70659: inst = 32'hca00004;
      70660: inst = 32'h38632800;
      70661: inst = 32'h38842800;
      70662: inst = 32'h10a00001;
      70663: inst = 32'hca0140b;
      70664: inst = 32'h13e00001;
      70665: inst = 32'hfe0d96a;
      70666: inst = 32'h5be00000;
      70667: inst = 32'h8c50000;
      70668: inst = 32'h24612800;
      70669: inst = 32'h10a0ffff;
      70670: inst = 32'hca0fffa;
      70671: inst = 32'h24822800;
      70672: inst = 32'h10a00000;
      70673: inst = 32'hca00004;
      70674: inst = 32'h38632800;
      70675: inst = 32'h38842800;
      70676: inst = 32'h10a00001;
      70677: inst = 32'hca01419;
      70678: inst = 32'h13e00001;
      70679: inst = 32'hfe0d96a;
      70680: inst = 32'h5be00000;
      70681: inst = 32'h8c50000;
      70682: inst = 32'h24612800;
      70683: inst = 32'h10a0ffff;
      70684: inst = 32'hca0fffa;
      70685: inst = 32'h24822800;
      70686: inst = 32'h10a00000;
      70687: inst = 32'hca00004;
      70688: inst = 32'h38632800;
      70689: inst = 32'h38842800;
      70690: inst = 32'h10a00001;
      70691: inst = 32'hca01427;
      70692: inst = 32'h13e00001;
      70693: inst = 32'hfe0d96a;
      70694: inst = 32'h5be00000;
      70695: inst = 32'h8c50000;
      70696: inst = 32'h24612800;
      70697: inst = 32'h10a0ffff;
      70698: inst = 32'hca0fffa;
      70699: inst = 32'h24822800;
      70700: inst = 32'h10a00000;
      70701: inst = 32'hca00004;
      70702: inst = 32'h38632800;
      70703: inst = 32'h38842800;
      70704: inst = 32'h10a00001;
      70705: inst = 32'hca01435;
      70706: inst = 32'h13e00001;
      70707: inst = 32'hfe0d96a;
      70708: inst = 32'h5be00000;
      70709: inst = 32'h8c50000;
      70710: inst = 32'h24612800;
      70711: inst = 32'h10a0ffff;
      70712: inst = 32'hca0fffa;
      70713: inst = 32'h24822800;
      70714: inst = 32'h10a00000;
      70715: inst = 32'hca00004;
      70716: inst = 32'h38632800;
      70717: inst = 32'h38842800;
      70718: inst = 32'h10a00001;
      70719: inst = 32'hca01443;
      70720: inst = 32'h13e00001;
      70721: inst = 32'hfe0d96a;
      70722: inst = 32'h5be00000;
      70723: inst = 32'h8c50000;
      70724: inst = 32'h24612800;
      70725: inst = 32'h10a0ffff;
      70726: inst = 32'hca0fffa;
      70727: inst = 32'h24822800;
      70728: inst = 32'h10a00000;
      70729: inst = 32'hca00004;
      70730: inst = 32'h38632800;
      70731: inst = 32'h38842800;
      70732: inst = 32'h10a00001;
      70733: inst = 32'hca01451;
      70734: inst = 32'h13e00001;
      70735: inst = 32'hfe0d96a;
      70736: inst = 32'h5be00000;
      70737: inst = 32'h8c50000;
      70738: inst = 32'h24612800;
      70739: inst = 32'h10a0ffff;
      70740: inst = 32'hca0fffa;
      70741: inst = 32'h24822800;
      70742: inst = 32'h10a00000;
      70743: inst = 32'hca00004;
      70744: inst = 32'h38632800;
      70745: inst = 32'h38842800;
      70746: inst = 32'h10a00001;
      70747: inst = 32'hca0145f;
      70748: inst = 32'h13e00001;
      70749: inst = 32'hfe0d96a;
      70750: inst = 32'h5be00000;
      70751: inst = 32'h8c50000;
      70752: inst = 32'h24612800;
      70753: inst = 32'h10a0ffff;
      70754: inst = 32'hca0fffa;
      70755: inst = 32'h24822800;
      70756: inst = 32'h10a00000;
      70757: inst = 32'hca00004;
      70758: inst = 32'h38632800;
      70759: inst = 32'h38842800;
      70760: inst = 32'h10a00001;
      70761: inst = 32'hca0146d;
      70762: inst = 32'h13e00001;
      70763: inst = 32'hfe0d96a;
      70764: inst = 32'h5be00000;
      70765: inst = 32'h8c50000;
      70766: inst = 32'h24612800;
      70767: inst = 32'h10a0ffff;
      70768: inst = 32'hca0fffa;
      70769: inst = 32'h24822800;
      70770: inst = 32'h10a00000;
      70771: inst = 32'hca00004;
      70772: inst = 32'h38632800;
      70773: inst = 32'h38842800;
      70774: inst = 32'h10a00001;
      70775: inst = 32'hca0147b;
      70776: inst = 32'h13e00001;
      70777: inst = 32'hfe0d96a;
      70778: inst = 32'h5be00000;
      70779: inst = 32'h8c50000;
      70780: inst = 32'h24612800;
      70781: inst = 32'h10a0ffff;
      70782: inst = 32'hca0fffa;
      70783: inst = 32'h24822800;
      70784: inst = 32'h10a00000;
      70785: inst = 32'hca00004;
      70786: inst = 32'h38632800;
      70787: inst = 32'h38842800;
      70788: inst = 32'h10a00001;
      70789: inst = 32'hca01489;
      70790: inst = 32'h13e00001;
      70791: inst = 32'hfe0d96a;
      70792: inst = 32'h5be00000;
      70793: inst = 32'h8c50000;
      70794: inst = 32'h24612800;
      70795: inst = 32'h10a0ffff;
      70796: inst = 32'hca0fffa;
      70797: inst = 32'h24822800;
      70798: inst = 32'h10a00000;
      70799: inst = 32'hca00004;
      70800: inst = 32'h38632800;
      70801: inst = 32'h38842800;
      70802: inst = 32'h10a00001;
      70803: inst = 32'hca01497;
      70804: inst = 32'h13e00001;
      70805: inst = 32'hfe0d96a;
      70806: inst = 32'h5be00000;
      70807: inst = 32'h8c50000;
      70808: inst = 32'h24612800;
      70809: inst = 32'h10a0ffff;
      70810: inst = 32'hca0fffa;
      70811: inst = 32'h24822800;
      70812: inst = 32'h10a00000;
      70813: inst = 32'hca00004;
      70814: inst = 32'h38632800;
      70815: inst = 32'h38842800;
      70816: inst = 32'h10a00001;
      70817: inst = 32'hca014a5;
      70818: inst = 32'h13e00001;
      70819: inst = 32'hfe0d96a;
      70820: inst = 32'h5be00000;
      70821: inst = 32'h8c50000;
      70822: inst = 32'h24612800;
      70823: inst = 32'h10a0ffff;
      70824: inst = 32'hca0fffa;
      70825: inst = 32'h24822800;
      70826: inst = 32'h10a00000;
      70827: inst = 32'hca00004;
      70828: inst = 32'h38632800;
      70829: inst = 32'h38842800;
      70830: inst = 32'h10a00001;
      70831: inst = 32'hca014b3;
      70832: inst = 32'h13e00001;
      70833: inst = 32'hfe0d96a;
      70834: inst = 32'h5be00000;
      70835: inst = 32'h8c50000;
      70836: inst = 32'h24612800;
      70837: inst = 32'h10a0ffff;
      70838: inst = 32'hca0fffa;
      70839: inst = 32'h24822800;
      70840: inst = 32'h10a00000;
      70841: inst = 32'hca00004;
      70842: inst = 32'h38632800;
      70843: inst = 32'h38842800;
      70844: inst = 32'h10a00001;
      70845: inst = 32'hca014c1;
      70846: inst = 32'h13e00001;
      70847: inst = 32'hfe0d96a;
      70848: inst = 32'h5be00000;
      70849: inst = 32'h8c50000;
      70850: inst = 32'h24612800;
      70851: inst = 32'h10a0ffff;
      70852: inst = 32'hca0fffa;
      70853: inst = 32'h24822800;
      70854: inst = 32'h10a00000;
      70855: inst = 32'hca00004;
      70856: inst = 32'h38632800;
      70857: inst = 32'h38842800;
      70858: inst = 32'h10a00001;
      70859: inst = 32'hca014cf;
      70860: inst = 32'h13e00001;
      70861: inst = 32'hfe0d96a;
      70862: inst = 32'h5be00000;
      70863: inst = 32'h8c50000;
      70864: inst = 32'h24612800;
      70865: inst = 32'h10a0ffff;
      70866: inst = 32'hca0fffa;
      70867: inst = 32'h24822800;
      70868: inst = 32'h10a00000;
      70869: inst = 32'hca00004;
      70870: inst = 32'h38632800;
      70871: inst = 32'h38842800;
      70872: inst = 32'h10a00001;
      70873: inst = 32'hca014dd;
      70874: inst = 32'h13e00001;
      70875: inst = 32'hfe0d96a;
      70876: inst = 32'h5be00000;
      70877: inst = 32'h8c50000;
      70878: inst = 32'h24612800;
      70879: inst = 32'h10a0ffff;
      70880: inst = 32'hca0fffa;
      70881: inst = 32'h24822800;
      70882: inst = 32'h10a00000;
      70883: inst = 32'hca00004;
      70884: inst = 32'h38632800;
      70885: inst = 32'h38842800;
      70886: inst = 32'h10a00001;
      70887: inst = 32'hca014eb;
      70888: inst = 32'h13e00001;
      70889: inst = 32'hfe0d96a;
      70890: inst = 32'h5be00000;
      70891: inst = 32'h8c50000;
      70892: inst = 32'h24612800;
      70893: inst = 32'h10a0ffff;
      70894: inst = 32'hca0fffa;
      70895: inst = 32'h24822800;
      70896: inst = 32'h10a00000;
      70897: inst = 32'hca00004;
      70898: inst = 32'h38632800;
      70899: inst = 32'h38842800;
      70900: inst = 32'h10a00001;
      70901: inst = 32'hca014f9;
      70902: inst = 32'h13e00001;
      70903: inst = 32'hfe0d96a;
      70904: inst = 32'h5be00000;
      70905: inst = 32'h8c50000;
      70906: inst = 32'h24612800;
      70907: inst = 32'h10a0ffff;
      70908: inst = 32'hca0fffa;
      70909: inst = 32'h24822800;
      70910: inst = 32'h10a00000;
      70911: inst = 32'hca00004;
      70912: inst = 32'h38632800;
      70913: inst = 32'h38842800;
      70914: inst = 32'h10a00001;
      70915: inst = 32'hca01507;
      70916: inst = 32'h13e00001;
      70917: inst = 32'hfe0d96a;
      70918: inst = 32'h5be00000;
      70919: inst = 32'h8c50000;
      70920: inst = 32'h24612800;
      70921: inst = 32'h10a0ffff;
      70922: inst = 32'hca0fffa;
      70923: inst = 32'h24822800;
      70924: inst = 32'h10a00000;
      70925: inst = 32'hca00004;
      70926: inst = 32'h38632800;
      70927: inst = 32'h38842800;
      70928: inst = 32'h10a00001;
      70929: inst = 32'hca01515;
      70930: inst = 32'h13e00001;
      70931: inst = 32'hfe0d96a;
      70932: inst = 32'h5be00000;
      70933: inst = 32'h8c50000;
      70934: inst = 32'h24612800;
      70935: inst = 32'h10a0ffff;
      70936: inst = 32'hca0fffa;
      70937: inst = 32'h24822800;
      70938: inst = 32'h10a00000;
      70939: inst = 32'hca00004;
      70940: inst = 32'h38632800;
      70941: inst = 32'h38842800;
      70942: inst = 32'h10a00001;
      70943: inst = 32'hca01523;
      70944: inst = 32'h13e00001;
      70945: inst = 32'hfe0d96a;
      70946: inst = 32'h5be00000;
      70947: inst = 32'h8c50000;
      70948: inst = 32'h24612800;
      70949: inst = 32'h10a0ffff;
      70950: inst = 32'hca0fffa;
      70951: inst = 32'h24822800;
      70952: inst = 32'h10a00000;
      70953: inst = 32'hca00004;
      70954: inst = 32'h38632800;
      70955: inst = 32'h38842800;
      70956: inst = 32'h10a00001;
      70957: inst = 32'hca01531;
      70958: inst = 32'h13e00001;
      70959: inst = 32'hfe0d96a;
      70960: inst = 32'h5be00000;
      70961: inst = 32'h8c50000;
      70962: inst = 32'h24612800;
      70963: inst = 32'h10a0ffff;
      70964: inst = 32'hca0fffa;
      70965: inst = 32'h24822800;
      70966: inst = 32'h10a00000;
      70967: inst = 32'hca00004;
      70968: inst = 32'h38632800;
      70969: inst = 32'h38842800;
      70970: inst = 32'h10a00001;
      70971: inst = 32'hca0153f;
      70972: inst = 32'h13e00001;
      70973: inst = 32'hfe0d96a;
      70974: inst = 32'h5be00000;
      70975: inst = 32'h8c50000;
      70976: inst = 32'h24612800;
      70977: inst = 32'h10a0ffff;
      70978: inst = 32'hca0fffa;
      70979: inst = 32'h24822800;
      70980: inst = 32'h10a00000;
      70981: inst = 32'hca00004;
      70982: inst = 32'h38632800;
      70983: inst = 32'h38842800;
      70984: inst = 32'h10a00001;
      70985: inst = 32'hca0154d;
      70986: inst = 32'h13e00001;
      70987: inst = 32'hfe0d96a;
      70988: inst = 32'h5be00000;
      70989: inst = 32'h8c50000;
      70990: inst = 32'h24612800;
      70991: inst = 32'h10a0ffff;
      70992: inst = 32'hca0fffa;
      70993: inst = 32'h24822800;
      70994: inst = 32'h10a00000;
      70995: inst = 32'hca00004;
      70996: inst = 32'h38632800;
      70997: inst = 32'h38842800;
      70998: inst = 32'h10a00001;
      70999: inst = 32'hca0155b;
      71000: inst = 32'h13e00001;
      71001: inst = 32'hfe0d96a;
      71002: inst = 32'h5be00000;
      71003: inst = 32'h8c50000;
      71004: inst = 32'h24612800;
      71005: inst = 32'h10a0ffff;
      71006: inst = 32'hca0fffa;
      71007: inst = 32'h24822800;
      71008: inst = 32'h10a00000;
      71009: inst = 32'hca00004;
      71010: inst = 32'h38632800;
      71011: inst = 32'h38842800;
      71012: inst = 32'h10a00001;
      71013: inst = 32'hca01569;
      71014: inst = 32'h13e00001;
      71015: inst = 32'hfe0d96a;
      71016: inst = 32'h5be00000;
      71017: inst = 32'h8c50000;
      71018: inst = 32'h24612800;
      71019: inst = 32'h10a0ffff;
      71020: inst = 32'hca0fffa;
      71021: inst = 32'h24822800;
      71022: inst = 32'h10a00000;
      71023: inst = 32'hca00004;
      71024: inst = 32'h38632800;
      71025: inst = 32'h38842800;
      71026: inst = 32'h10a00001;
      71027: inst = 32'hca01577;
      71028: inst = 32'h13e00001;
      71029: inst = 32'hfe0d96a;
      71030: inst = 32'h5be00000;
      71031: inst = 32'h8c50000;
      71032: inst = 32'h24612800;
      71033: inst = 32'h10a0ffff;
      71034: inst = 32'hca0fffa;
      71035: inst = 32'h24822800;
      71036: inst = 32'h10a00000;
      71037: inst = 32'hca00004;
      71038: inst = 32'h38632800;
      71039: inst = 32'h38842800;
      71040: inst = 32'h10a00001;
      71041: inst = 32'hca01585;
      71042: inst = 32'h13e00001;
      71043: inst = 32'hfe0d96a;
      71044: inst = 32'h5be00000;
      71045: inst = 32'h8c50000;
      71046: inst = 32'h24612800;
      71047: inst = 32'h10a0ffff;
      71048: inst = 32'hca0fffa;
      71049: inst = 32'h24822800;
      71050: inst = 32'h10a00000;
      71051: inst = 32'hca00004;
      71052: inst = 32'h38632800;
      71053: inst = 32'h38842800;
      71054: inst = 32'h10a00001;
      71055: inst = 32'hca01593;
      71056: inst = 32'h13e00001;
      71057: inst = 32'hfe0d96a;
      71058: inst = 32'h5be00000;
      71059: inst = 32'h8c50000;
      71060: inst = 32'h24612800;
      71061: inst = 32'h10a0ffff;
      71062: inst = 32'hca0fffa;
      71063: inst = 32'h24822800;
      71064: inst = 32'h10a00000;
      71065: inst = 32'hca00004;
      71066: inst = 32'h38632800;
      71067: inst = 32'h38842800;
      71068: inst = 32'h10a00001;
      71069: inst = 32'hca015a1;
      71070: inst = 32'h13e00001;
      71071: inst = 32'hfe0d96a;
      71072: inst = 32'h5be00000;
      71073: inst = 32'h8c50000;
      71074: inst = 32'h24612800;
      71075: inst = 32'h10a0ffff;
      71076: inst = 32'hca0fffa;
      71077: inst = 32'h24822800;
      71078: inst = 32'h10a00000;
      71079: inst = 32'hca00004;
      71080: inst = 32'h38632800;
      71081: inst = 32'h38842800;
      71082: inst = 32'h10a00001;
      71083: inst = 32'hca015af;
      71084: inst = 32'h13e00001;
      71085: inst = 32'hfe0d96a;
      71086: inst = 32'h5be00000;
      71087: inst = 32'h8c50000;
      71088: inst = 32'h24612800;
      71089: inst = 32'h10a0ffff;
      71090: inst = 32'hca0fffa;
      71091: inst = 32'h24822800;
      71092: inst = 32'h10a00000;
      71093: inst = 32'hca00004;
      71094: inst = 32'h38632800;
      71095: inst = 32'h38842800;
      71096: inst = 32'h10a00001;
      71097: inst = 32'hca015bd;
      71098: inst = 32'h13e00001;
      71099: inst = 32'hfe0d96a;
      71100: inst = 32'h5be00000;
      71101: inst = 32'h8c50000;
      71102: inst = 32'h24612800;
      71103: inst = 32'h10a0ffff;
      71104: inst = 32'hca0fffa;
      71105: inst = 32'h24822800;
      71106: inst = 32'h10a00000;
      71107: inst = 32'hca00004;
      71108: inst = 32'h38632800;
      71109: inst = 32'h38842800;
      71110: inst = 32'h10a00001;
      71111: inst = 32'hca015cb;
      71112: inst = 32'h13e00001;
      71113: inst = 32'hfe0d96a;
      71114: inst = 32'h5be00000;
      71115: inst = 32'h8c50000;
      71116: inst = 32'h24612800;
      71117: inst = 32'h10a0ffff;
      71118: inst = 32'hca0fffa;
      71119: inst = 32'h24822800;
      71120: inst = 32'h10a00000;
      71121: inst = 32'hca00004;
      71122: inst = 32'h38632800;
      71123: inst = 32'h38842800;
      71124: inst = 32'h10a00001;
      71125: inst = 32'hca015d9;
      71126: inst = 32'h13e00001;
      71127: inst = 32'hfe0d96a;
      71128: inst = 32'h5be00000;
      71129: inst = 32'h8c50000;
      71130: inst = 32'h24612800;
      71131: inst = 32'h10a0ffff;
      71132: inst = 32'hca0fffa;
      71133: inst = 32'h24822800;
      71134: inst = 32'h10a00000;
      71135: inst = 32'hca00004;
      71136: inst = 32'h38632800;
      71137: inst = 32'h38842800;
      71138: inst = 32'h10a00001;
      71139: inst = 32'hca015e7;
      71140: inst = 32'h13e00001;
      71141: inst = 32'hfe0d96a;
      71142: inst = 32'h5be00000;
      71143: inst = 32'h8c50000;
      71144: inst = 32'h24612800;
      71145: inst = 32'h10a0ffff;
      71146: inst = 32'hca0fffa;
      71147: inst = 32'h24822800;
      71148: inst = 32'h10a00000;
      71149: inst = 32'hca00004;
      71150: inst = 32'h38632800;
      71151: inst = 32'h38842800;
      71152: inst = 32'h10a00001;
      71153: inst = 32'hca015f5;
      71154: inst = 32'h13e00001;
      71155: inst = 32'hfe0d96a;
      71156: inst = 32'h5be00000;
      71157: inst = 32'h8c50000;
      71158: inst = 32'h24612800;
      71159: inst = 32'h10a0ffff;
      71160: inst = 32'hca0fffa;
      71161: inst = 32'h24822800;
      71162: inst = 32'h10a00000;
      71163: inst = 32'hca00004;
      71164: inst = 32'h38632800;
      71165: inst = 32'h38842800;
      71166: inst = 32'h10a00001;
      71167: inst = 32'hca01603;
      71168: inst = 32'h13e00001;
      71169: inst = 32'hfe0d96a;
      71170: inst = 32'h5be00000;
      71171: inst = 32'h8c50000;
      71172: inst = 32'h24612800;
      71173: inst = 32'h10a0ffff;
      71174: inst = 32'hca0fffa;
      71175: inst = 32'h24822800;
      71176: inst = 32'h10a00000;
      71177: inst = 32'hca00004;
      71178: inst = 32'h38632800;
      71179: inst = 32'h38842800;
      71180: inst = 32'h10a00001;
      71181: inst = 32'hca01611;
      71182: inst = 32'h13e00001;
      71183: inst = 32'hfe0d96a;
      71184: inst = 32'h5be00000;
      71185: inst = 32'h8c50000;
      71186: inst = 32'h24612800;
      71187: inst = 32'h10a0ffff;
      71188: inst = 32'hca0fffa;
      71189: inst = 32'h24822800;
      71190: inst = 32'h10a00000;
      71191: inst = 32'hca00004;
      71192: inst = 32'h38632800;
      71193: inst = 32'h38842800;
      71194: inst = 32'h10a00001;
      71195: inst = 32'hca0161f;
      71196: inst = 32'h13e00001;
      71197: inst = 32'hfe0d96a;
      71198: inst = 32'h5be00000;
      71199: inst = 32'h8c50000;
      71200: inst = 32'h24612800;
      71201: inst = 32'h10a0ffff;
      71202: inst = 32'hca0fffa;
      71203: inst = 32'h24822800;
      71204: inst = 32'h10a00000;
      71205: inst = 32'hca00004;
      71206: inst = 32'h38632800;
      71207: inst = 32'h38842800;
      71208: inst = 32'h10a00001;
      71209: inst = 32'hca0162d;
      71210: inst = 32'h13e00001;
      71211: inst = 32'hfe0d96a;
      71212: inst = 32'h5be00000;
      71213: inst = 32'h8c50000;
      71214: inst = 32'h24612800;
      71215: inst = 32'h10a0ffff;
      71216: inst = 32'hca0fffa;
      71217: inst = 32'h24822800;
      71218: inst = 32'h10a00000;
      71219: inst = 32'hca00004;
      71220: inst = 32'h38632800;
      71221: inst = 32'h38842800;
      71222: inst = 32'h10a00001;
      71223: inst = 32'hca0163b;
      71224: inst = 32'h13e00001;
      71225: inst = 32'hfe0d96a;
      71226: inst = 32'h5be00000;
      71227: inst = 32'h8c50000;
      71228: inst = 32'h24612800;
      71229: inst = 32'h10a0ffff;
      71230: inst = 32'hca0fffa;
      71231: inst = 32'h24822800;
      71232: inst = 32'h10a00000;
      71233: inst = 32'hca00004;
      71234: inst = 32'h38632800;
      71235: inst = 32'h38842800;
      71236: inst = 32'h10a00001;
      71237: inst = 32'hca01649;
      71238: inst = 32'h13e00001;
      71239: inst = 32'hfe0d96a;
      71240: inst = 32'h5be00000;
      71241: inst = 32'h8c50000;
      71242: inst = 32'h24612800;
      71243: inst = 32'h10a0ffff;
      71244: inst = 32'hca0fffa;
      71245: inst = 32'h24822800;
      71246: inst = 32'h10a00000;
      71247: inst = 32'hca00004;
      71248: inst = 32'h38632800;
      71249: inst = 32'h38842800;
      71250: inst = 32'h10a00001;
      71251: inst = 32'hca01657;
      71252: inst = 32'h13e00001;
      71253: inst = 32'hfe0d96a;
      71254: inst = 32'h5be00000;
      71255: inst = 32'h8c50000;
      71256: inst = 32'h24612800;
      71257: inst = 32'h10a0ffff;
      71258: inst = 32'hca0fffa;
      71259: inst = 32'h24822800;
      71260: inst = 32'h10a00000;
      71261: inst = 32'hca00004;
      71262: inst = 32'h38632800;
      71263: inst = 32'h38842800;
      71264: inst = 32'h10a00001;
      71265: inst = 32'hca01665;
      71266: inst = 32'h13e00001;
      71267: inst = 32'hfe0d96a;
      71268: inst = 32'h5be00000;
      71269: inst = 32'h8c50000;
      71270: inst = 32'h24612800;
      71271: inst = 32'h10a0ffff;
      71272: inst = 32'hca0fffa;
      71273: inst = 32'h24822800;
      71274: inst = 32'h10a00000;
      71275: inst = 32'hca00004;
      71276: inst = 32'h38632800;
      71277: inst = 32'h38842800;
      71278: inst = 32'h10a00001;
      71279: inst = 32'hca01673;
      71280: inst = 32'h13e00001;
      71281: inst = 32'hfe0d96a;
      71282: inst = 32'h5be00000;
      71283: inst = 32'h8c50000;
      71284: inst = 32'h24612800;
      71285: inst = 32'h10a0ffff;
      71286: inst = 32'hca0fffa;
      71287: inst = 32'h24822800;
      71288: inst = 32'h10a00000;
      71289: inst = 32'hca00004;
      71290: inst = 32'h38632800;
      71291: inst = 32'h38842800;
      71292: inst = 32'h10a00001;
      71293: inst = 32'hca01681;
      71294: inst = 32'h13e00001;
      71295: inst = 32'hfe0d96a;
      71296: inst = 32'h5be00000;
      71297: inst = 32'h8c50000;
      71298: inst = 32'h24612800;
      71299: inst = 32'h10a0ffff;
      71300: inst = 32'hca0fffa;
      71301: inst = 32'h24822800;
      71302: inst = 32'h10a00000;
      71303: inst = 32'hca00004;
      71304: inst = 32'h38632800;
      71305: inst = 32'h38842800;
      71306: inst = 32'h10a00001;
      71307: inst = 32'hca0168f;
      71308: inst = 32'h13e00001;
      71309: inst = 32'hfe0d96a;
      71310: inst = 32'h5be00000;
      71311: inst = 32'h8c50000;
      71312: inst = 32'h24612800;
      71313: inst = 32'h10a0ffff;
      71314: inst = 32'hca0fffa;
      71315: inst = 32'h24822800;
      71316: inst = 32'h10a00000;
      71317: inst = 32'hca00004;
      71318: inst = 32'h38632800;
      71319: inst = 32'h38842800;
      71320: inst = 32'h10a00001;
      71321: inst = 32'hca0169d;
      71322: inst = 32'h13e00001;
      71323: inst = 32'hfe0d96a;
      71324: inst = 32'h5be00000;
      71325: inst = 32'h8c50000;
      71326: inst = 32'h24612800;
      71327: inst = 32'h10a0ffff;
      71328: inst = 32'hca0fffa;
      71329: inst = 32'h24822800;
      71330: inst = 32'h10a00000;
      71331: inst = 32'hca00004;
      71332: inst = 32'h38632800;
      71333: inst = 32'h38842800;
      71334: inst = 32'h10a00001;
      71335: inst = 32'hca016ab;
      71336: inst = 32'h13e00001;
      71337: inst = 32'hfe0d96a;
      71338: inst = 32'h5be00000;
      71339: inst = 32'h8c50000;
      71340: inst = 32'h24612800;
      71341: inst = 32'h10a0ffff;
      71342: inst = 32'hca0fffa;
      71343: inst = 32'h24822800;
      71344: inst = 32'h10a00000;
      71345: inst = 32'hca00004;
      71346: inst = 32'h38632800;
      71347: inst = 32'h38842800;
      71348: inst = 32'h10a00001;
      71349: inst = 32'hca016b9;
      71350: inst = 32'h13e00001;
      71351: inst = 32'hfe0d96a;
      71352: inst = 32'h5be00000;
      71353: inst = 32'h8c50000;
      71354: inst = 32'h24612800;
      71355: inst = 32'h10a0ffff;
      71356: inst = 32'hca0fffa;
      71357: inst = 32'h24822800;
      71358: inst = 32'h10a00000;
      71359: inst = 32'hca00004;
      71360: inst = 32'h38632800;
      71361: inst = 32'h38842800;
      71362: inst = 32'h10a00001;
      71363: inst = 32'hca016c7;
      71364: inst = 32'h13e00001;
      71365: inst = 32'hfe0d96a;
      71366: inst = 32'h5be00000;
      71367: inst = 32'h8c50000;
      71368: inst = 32'h24612800;
      71369: inst = 32'h10a0ffff;
      71370: inst = 32'hca0fffa;
      71371: inst = 32'h24822800;
      71372: inst = 32'h10a00000;
      71373: inst = 32'hca00004;
      71374: inst = 32'h38632800;
      71375: inst = 32'h38842800;
      71376: inst = 32'h10a00001;
      71377: inst = 32'hca016d5;
      71378: inst = 32'h13e00001;
      71379: inst = 32'hfe0d96a;
      71380: inst = 32'h5be00000;
      71381: inst = 32'h8c50000;
      71382: inst = 32'h24612800;
      71383: inst = 32'h10a0ffff;
      71384: inst = 32'hca0fffa;
      71385: inst = 32'h24822800;
      71386: inst = 32'h10a00000;
      71387: inst = 32'hca00004;
      71388: inst = 32'h38632800;
      71389: inst = 32'h38842800;
      71390: inst = 32'h10a00001;
      71391: inst = 32'hca016e3;
      71392: inst = 32'h13e00001;
      71393: inst = 32'hfe0d96a;
      71394: inst = 32'h5be00000;
      71395: inst = 32'h8c50000;
      71396: inst = 32'h24612800;
      71397: inst = 32'h10a0ffff;
      71398: inst = 32'hca0fffa;
      71399: inst = 32'h24822800;
      71400: inst = 32'h10a00000;
      71401: inst = 32'hca00004;
      71402: inst = 32'h38632800;
      71403: inst = 32'h38842800;
      71404: inst = 32'h10a00001;
      71405: inst = 32'hca016f1;
      71406: inst = 32'h13e00001;
      71407: inst = 32'hfe0d96a;
      71408: inst = 32'h5be00000;
      71409: inst = 32'h8c50000;
      71410: inst = 32'h24612800;
      71411: inst = 32'h10a0ffff;
      71412: inst = 32'hca0fffa;
      71413: inst = 32'h24822800;
      71414: inst = 32'h10a00000;
      71415: inst = 32'hca00004;
      71416: inst = 32'h38632800;
      71417: inst = 32'h38842800;
      71418: inst = 32'h10a00001;
      71419: inst = 32'hca016ff;
      71420: inst = 32'h13e00001;
      71421: inst = 32'hfe0d96a;
      71422: inst = 32'h5be00000;
      71423: inst = 32'h8c50000;
      71424: inst = 32'h24612800;
      71425: inst = 32'h10a0ffff;
      71426: inst = 32'hca0fffa;
      71427: inst = 32'h24822800;
      71428: inst = 32'h10a00000;
      71429: inst = 32'hca00004;
      71430: inst = 32'h38632800;
      71431: inst = 32'h38842800;
      71432: inst = 32'h10a00001;
      71433: inst = 32'hca0170d;
      71434: inst = 32'h13e00001;
      71435: inst = 32'hfe0d96a;
      71436: inst = 32'h5be00000;
      71437: inst = 32'h8c50000;
      71438: inst = 32'h24612800;
      71439: inst = 32'h10a0ffff;
      71440: inst = 32'hca0fffa;
      71441: inst = 32'h24822800;
      71442: inst = 32'h10a00000;
      71443: inst = 32'hca00004;
      71444: inst = 32'h38632800;
      71445: inst = 32'h38842800;
      71446: inst = 32'h10a00001;
      71447: inst = 32'hca0171b;
      71448: inst = 32'h13e00001;
      71449: inst = 32'hfe0d96a;
      71450: inst = 32'h5be00000;
      71451: inst = 32'h8c50000;
      71452: inst = 32'h24612800;
      71453: inst = 32'h10a0ffff;
      71454: inst = 32'hca0fffa;
      71455: inst = 32'h24822800;
      71456: inst = 32'h10a00000;
      71457: inst = 32'hca00004;
      71458: inst = 32'h38632800;
      71459: inst = 32'h38842800;
      71460: inst = 32'h10a00001;
      71461: inst = 32'hca01729;
      71462: inst = 32'h13e00001;
      71463: inst = 32'hfe0d96a;
      71464: inst = 32'h5be00000;
      71465: inst = 32'h8c50000;
      71466: inst = 32'h24612800;
      71467: inst = 32'h10a0ffff;
      71468: inst = 32'hca0fffb;
      71469: inst = 32'h24822800;
      71470: inst = 32'h10a00000;
      71471: inst = 32'hca00004;
      71472: inst = 32'h38632800;
      71473: inst = 32'h38842800;
      71474: inst = 32'h10a00001;
      71475: inst = 32'hca01737;
      71476: inst = 32'h13e00001;
      71477: inst = 32'hfe0d96a;
      71478: inst = 32'h5be00000;
      71479: inst = 32'h8c50000;
      71480: inst = 32'h24612800;
      71481: inst = 32'h10a0ffff;
      71482: inst = 32'hca0fffb;
      71483: inst = 32'h24822800;
      71484: inst = 32'h10a00000;
      71485: inst = 32'hca00004;
      71486: inst = 32'h38632800;
      71487: inst = 32'h38842800;
      71488: inst = 32'h10a00001;
      71489: inst = 32'hca01745;
      71490: inst = 32'h13e00001;
      71491: inst = 32'hfe0d96a;
      71492: inst = 32'h5be00000;
      71493: inst = 32'h8c50000;
      71494: inst = 32'h24612800;
      71495: inst = 32'h10a0ffff;
      71496: inst = 32'hca0fffb;
      71497: inst = 32'h24822800;
      71498: inst = 32'h10a00000;
      71499: inst = 32'hca00004;
      71500: inst = 32'h38632800;
      71501: inst = 32'h38842800;
      71502: inst = 32'h10a00001;
      71503: inst = 32'hca01753;
      71504: inst = 32'h13e00001;
      71505: inst = 32'hfe0d96a;
      71506: inst = 32'h5be00000;
      71507: inst = 32'h8c50000;
      71508: inst = 32'h24612800;
      71509: inst = 32'h10a0ffff;
      71510: inst = 32'hca0fffb;
      71511: inst = 32'h24822800;
      71512: inst = 32'h10a00000;
      71513: inst = 32'hca00004;
      71514: inst = 32'h38632800;
      71515: inst = 32'h38842800;
      71516: inst = 32'h10a00001;
      71517: inst = 32'hca01761;
      71518: inst = 32'h13e00001;
      71519: inst = 32'hfe0d96a;
      71520: inst = 32'h5be00000;
      71521: inst = 32'h8c50000;
      71522: inst = 32'h24612800;
      71523: inst = 32'h10a0ffff;
      71524: inst = 32'hca0fffb;
      71525: inst = 32'h24822800;
      71526: inst = 32'h10a00000;
      71527: inst = 32'hca00004;
      71528: inst = 32'h38632800;
      71529: inst = 32'h38842800;
      71530: inst = 32'h10a00001;
      71531: inst = 32'hca0176f;
      71532: inst = 32'h13e00001;
      71533: inst = 32'hfe0d96a;
      71534: inst = 32'h5be00000;
      71535: inst = 32'h8c50000;
      71536: inst = 32'h24612800;
      71537: inst = 32'h10a0ffff;
      71538: inst = 32'hca0fffb;
      71539: inst = 32'h24822800;
      71540: inst = 32'h10a00000;
      71541: inst = 32'hca00004;
      71542: inst = 32'h38632800;
      71543: inst = 32'h38842800;
      71544: inst = 32'h10a00001;
      71545: inst = 32'hca0177d;
      71546: inst = 32'h13e00001;
      71547: inst = 32'hfe0d96a;
      71548: inst = 32'h5be00000;
      71549: inst = 32'h8c50000;
      71550: inst = 32'h24612800;
      71551: inst = 32'h10a0ffff;
      71552: inst = 32'hca0fffb;
      71553: inst = 32'h24822800;
      71554: inst = 32'h10a00000;
      71555: inst = 32'hca00004;
      71556: inst = 32'h38632800;
      71557: inst = 32'h38842800;
      71558: inst = 32'h10a00001;
      71559: inst = 32'hca0178b;
      71560: inst = 32'h13e00001;
      71561: inst = 32'hfe0d96a;
      71562: inst = 32'h5be00000;
      71563: inst = 32'h8c50000;
      71564: inst = 32'h24612800;
      71565: inst = 32'h10a0ffff;
      71566: inst = 32'hca0fffb;
      71567: inst = 32'h24822800;
      71568: inst = 32'h10a00000;
      71569: inst = 32'hca00004;
      71570: inst = 32'h38632800;
      71571: inst = 32'h38842800;
      71572: inst = 32'h10a00001;
      71573: inst = 32'hca01799;
      71574: inst = 32'h13e00001;
      71575: inst = 32'hfe0d96a;
      71576: inst = 32'h5be00000;
      71577: inst = 32'h8c50000;
      71578: inst = 32'h24612800;
      71579: inst = 32'h10a0ffff;
      71580: inst = 32'hca0fffb;
      71581: inst = 32'h24822800;
      71582: inst = 32'h10a00000;
      71583: inst = 32'hca00004;
      71584: inst = 32'h38632800;
      71585: inst = 32'h38842800;
      71586: inst = 32'h10a00001;
      71587: inst = 32'hca017a7;
      71588: inst = 32'h13e00001;
      71589: inst = 32'hfe0d96a;
      71590: inst = 32'h5be00000;
      71591: inst = 32'h8c50000;
      71592: inst = 32'h24612800;
      71593: inst = 32'h10a0ffff;
      71594: inst = 32'hca0fffb;
      71595: inst = 32'h24822800;
      71596: inst = 32'h10a00000;
      71597: inst = 32'hca00004;
      71598: inst = 32'h38632800;
      71599: inst = 32'h38842800;
      71600: inst = 32'h10a00001;
      71601: inst = 32'hca017b5;
      71602: inst = 32'h13e00001;
      71603: inst = 32'hfe0d96a;
      71604: inst = 32'h5be00000;
      71605: inst = 32'h8c50000;
      71606: inst = 32'h24612800;
      71607: inst = 32'h10a0ffff;
      71608: inst = 32'hca0fffb;
      71609: inst = 32'h24822800;
      71610: inst = 32'h10a00000;
      71611: inst = 32'hca00004;
      71612: inst = 32'h38632800;
      71613: inst = 32'h38842800;
      71614: inst = 32'h10a00001;
      71615: inst = 32'hca017c3;
      71616: inst = 32'h13e00001;
      71617: inst = 32'hfe0d96a;
      71618: inst = 32'h5be00000;
      71619: inst = 32'h8c50000;
      71620: inst = 32'h24612800;
      71621: inst = 32'h10a0ffff;
      71622: inst = 32'hca0fffb;
      71623: inst = 32'h24822800;
      71624: inst = 32'h10a00000;
      71625: inst = 32'hca00004;
      71626: inst = 32'h38632800;
      71627: inst = 32'h38842800;
      71628: inst = 32'h10a00001;
      71629: inst = 32'hca017d1;
      71630: inst = 32'h13e00001;
      71631: inst = 32'hfe0d96a;
      71632: inst = 32'h5be00000;
      71633: inst = 32'h8c50000;
      71634: inst = 32'h24612800;
      71635: inst = 32'h10a0ffff;
      71636: inst = 32'hca0fffb;
      71637: inst = 32'h24822800;
      71638: inst = 32'h10a00000;
      71639: inst = 32'hca00004;
      71640: inst = 32'h38632800;
      71641: inst = 32'h38842800;
      71642: inst = 32'h10a00001;
      71643: inst = 32'hca017df;
      71644: inst = 32'h13e00001;
      71645: inst = 32'hfe0d96a;
      71646: inst = 32'h5be00000;
      71647: inst = 32'h8c50000;
      71648: inst = 32'h24612800;
      71649: inst = 32'h10a0ffff;
      71650: inst = 32'hca0fffb;
      71651: inst = 32'h24822800;
      71652: inst = 32'h10a00000;
      71653: inst = 32'hca00004;
      71654: inst = 32'h38632800;
      71655: inst = 32'h38842800;
      71656: inst = 32'h10a00001;
      71657: inst = 32'hca017ed;
      71658: inst = 32'h13e00001;
      71659: inst = 32'hfe0d96a;
      71660: inst = 32'h5be00000;
      71661: inst = 32'h8c50000;
      71662: inst = 32'h24612800;
      71663: inst = 32'h10a0ffff;
      71664: inst = 32'hca0fffb;
      71665: inst = 32'h24822800;
      71666: inst = 32'h10a00000;
      71667: inst = 32'hca00004;
      71668: inst = 32'h38632800;
      71669: inst = 32'h38842800;
      71670: inst = 32'h10a00001;
      71671: inst = 32'hca017fb;
      71672: inst = 32'h13e00001;
      71673: inst = 32'hfe0d96a;
      71674: inst = 32'h5be00000;
      71675: inst = 32'h8c50000;
      71676: inst = 32'h24612800;
      71677: inst = 32'h10a0ffff;
      71678: inst = 32'hca0fffb;
      71679: inst = 32'h24822800;
      71680: inst = 32'h10a00000;
      71681: inst = 32'hca00004;
      71682: inst = 32'h38632800;
      71683: inst = 32'h38842800;
      71684: inst = 32'h10a00001;
      71685: inst = 32'hca01809;
      71686: inst = 32'h13e00001;
      71687: inst = 32'hfe0d96a;
      71688: inst = 32'h5be00000;
      71689: inst = 32'h8c50000;
      71690: inst = 32'h24612800;
      71691: inst = 32'h10a0ffff;
      71692: inst = 32'hca0fffb;
      71693: inst = 32'h24822800;
      71694: inst = 32'h10a00000;
      71695: inst = 32'hca00004;
      71696: inst = 32'h38632800;
      71697: inst = 32'h38842800;
      71698: inst = 32'h10a00001;
      71699: inst = 32'hca01817;
      71700: inst = 32'h13e00001;
      71701: inst = 32'hfe0d96a;
      71702: inst = 32'h5be00000;
      71703: inst = 32'h8c50000;
      71704: inst = 32'h24612800;
      71705: inst = 32'h10a0ffff;
      71706: inst = 32'hca0fffb;
      71707: inst = 32'h24822800;
      71708: inst = 32'h10a00000;
      71709: inst = 32'hca00004;
      71710: inst = 32'h38632800;
      71711: inst = 32'h38842800;
      71712: inst = 32'h10a00001;
      71713: inst = 32'hca01825;
      71714: inst = 32'h13e00001;
      71715: inst = 32'hfe0d96a;
      71716: inst = 32'h5be00000;
      71717: inst = 32'h8c50000;
      71718: inst = 32'h24612800;
      71719: inst = 32'h10a0ffff;
      71720: inst = 32'hca0fffb;
      71721: inst = 32'h24822800;
      71722: inst = 32'h10a00000;
      71723: inst = 32'hca00004;
      71724: inst = 32'h38632800;
      71725: inst = 32'h38842800;
      71726: inst = 32'h10a00001;
      71727: inst = 32'hca01833;
      71728: inst = 32'h13e00001;
      71729: inst = 32'hfe0d96a;
      71730: inst = 32'h5be00000;
      71731: inst = 32'h8c50000;
      71732: inst = 32'h24612800;
      71733: inst = 32'h10a0ffff;
      71734: inst = 32'hca0fffb;
      71735: inst = 32'h24822800;
      71736: inst = 32'h10a00000;
      71737: inst = 32'hca00004;
      71738: inst = 32'h38632800;
      71739: inst = 32'h38842800;
      71740: inst = 32'h10a00001;
      71741: inst = 32'hca01841;
      71742: inst = 32'h13e00001;
      71743: inst = 32'hfe0d96a;
      71744: inst = 32'h5be00000;
      71745: inst = 32'h8c50000;
      71746: inst = 32'h24612800;
      71747: inst = 32'h10a0ffff;
      71748: inst = 32'hca0fffb;
      71749: inst = 32'h24822800;
      71750: inst = 32'h10a00000;
      71751: inst = 32'hca00004;
      71752: inst = 32'h38632800;
      71753: inst = 32'h38842800;
      71754: inst = 32'h10a00001;
      71755: inst = 32'hca0184f;
      71756: inst = 32'h13e00001;
      71757: inst = 32'hfe0d96a;
      71758: inst = 32'h5be00000;
      71759: inst = 32'h8c50000;
      71760: inst = 32'h24612800;
      71761: inst = 32'h10a0ffff;
      71762: inst = 32'hca0fffb;
      71763: inst = 32'h24822800;
      71764: inst = 32'h10a00000;
      71765: inst = 32'hca00004;
      71766: inst = 32'h38632800;
      71767: inst = 32'h38842800;
      71768: inst = 32'h10a00001;
      71769: inst = 32'hca0185d;
      71770: inst = 32'h13e00001;
      71771: inst = 32'hfe0d96a;
      71772: inst = 32'h5be00000;
      71773: inst = 32'h8c50000;
      71774: inst = 32'h24612800;
      71775: inst = 32'h10a0ffff;
      71776: inst = 32'hca0fffb;
      71777: inst = 32'h24822800;
      71778: inst = 32'h10a00000;
      71779: inst = 32'hca00004;
      71780: inst = 32'h38632800;
      71781: inst = 32'h38842800;
      71782: inst = 32'h10a00001;
      71783: inst = 32'hca0186b;
      71784: inst = 32'h13e00001;
      71785: inst = 32'hfe0d96a;
      71786: inst = 32'h5be00000;
      71787: inst = 32'h8c50000;
      71788: inst = 32'h24612800;
      71789: inst = 32'h10a0ffff;
      71790: inst = 32'hca0fffb;
      71791: inst = 32'h24822800;
      71792: inst = 32'h10a00000;
      71793: inst = 32'hca00004;
      71794: inst = 32'h38632800;
      71795: inst = 32'h38842800;
      71796: inst = 32'h10a00001;
      71797: inst = 32'hca01879;
      71798: inst = 32'h13e00001;
      71799: inst = 32'hfe0d96a;
      71800: inst = 32'h5be00000;
      71801: inst = 32'h8c50000;
      71802: inst = 32'h24612800;
      71803: inst = 32'h10a0ffff;
      71804: inst = 32'hca0fffb;
      71805: inst = 32'h24822800;
      71806: inst = 32'h10a00000;
      71807: inst = 32'hca00004;
      71808: inst = 32'h38632800;
      71809: inst = 32'h38842800;
      71810: inst = 32'h10a00001;
      71811: inst = 32'hca01887;
      71812: inst = 32'h13e00001;
      71813: inst = 32'hfe0d96a;
      71814: inst = 32'h5be00000;
      71815: inst = 32'h8c50000;
      71816: inst = 32'h24612800;
      71817: inst = 32'h10a0ffff;
      71818: inst = 32'hca0fffb;
      71819: inst = 32'h24822800;
      71820: inst = 32'h10a00000;
      71821: inst = 32'hca00004;
      71822: inst = 32'h38632800;
      71823: inst = 32'h38842800;
      71824: inst = 32'h10a00001;
      71825: inst = 32'hca01895;
      71826: inst = 32'h13e00001;
      71827: inst = 32'hfe0d96a;
      71828: inst = 32'h5be00000;
      71829: inst = 32'h8c50000;
      71830: inst = 32'h24612800;
      71831: inst = 32'h10a0ffff;
      71832: inst = 32'hca0fffb;
      71833: inst = 32'h24822800;
      71834: inst = 32'h10a00000;
      71835: inst = 32'hca00004;
      71836: inst = 32'h38632800;
      71837: inst = 32'h38842800;
      71838: inst = 32'h10a00001;
      71839: inst = 32'hca018a3;
      71840: inst = 32'h13e00001;
      71841: inst = 32'hfe0d96a;
      71842: inst = 32'h5be00000;
      71843: inst = 32'h8c50000;
      71844: inst = 32'h24612800;
      71845: inst = 32'h10a0ffff;
      71846: inst = 32'hca0fffb;
      71847: inst = 32'h24822800;
      71848: inst = 32'h10a00000;
      71849: inst = 32'hca00004;
      71850: inst = 32'h38632800;
      71851: inst = 32'h38842800;
      71852: inst = 32'h10a00001;
      71853: inst = 32'hca018b1;
      71854: inst = 32'h13e00001;
      71855: inst = 32'hfe0d96a;
      71856: inst = 32'h5be00000;
      71857: inst = 32'h8c50000;
      71858: inst = 32'h24612800;
      71859: inst = 32'h10a0ffff;
      71860: inst = 32'hca0fffb;
      71861: inst = 32'h24822800;
      71862: inst = 32'h10a00000;
      71863: inst = 32'hca00004;
      71864: inst = 32'h38632800;
      71865: inst = 32'h38842800;
      71866: inst = 32'h10a00001;
      71867: inst = 32'hca018bf;
      71868: inst = 32'h13e00001;
      71869: inst = 32'hfe0d96a;
      71870: inst = 32'h5be00000;
      71871: inst = 32'h8c50000;
      71872: inst = 32'h24612800;
      71873: inst = 32'h10a0ffff;
      71874: inst = 32'hca0fffb;
      71875: inst = 32'h24822800;
      71876: inst = 32'h10a00000;
      71877: inst = 32'hca00004;
      71878: inst = 32'h38632800;
      71879: inst = 32'h38842800;
      71880: inst = 32'h10a00001;
      71881: inst = 32'hca018cd;
      71882: inst = 32'h13e00001;
      71883: inst = 32'hfe0d96a;
      71884: inst = 32'h5be00000;
      71885: inst = 32'h8c50000;
      71886: inst = 32'h24612800;
      71887: inst = 32'h10a0ffff;
      71888: inst = 32'hca0fffb;
      71889: inst = 32'h24822800;
      71890: inst = 32'h10a00000;
      71891: inst = 32'hca00004;
      71892: inst = 32'h38632800;
      71893: inst = 32'h38842800;
      71894: inst = 32'h10a00001;
      71895: inst = 32'hca018db;
      71896: inst = 32'h13e00001;
      71897: inst = 32'hfe0d96a;
      71898: inst = 32'h5be00000;
      71899: inst = 32'h8c50000;
      71900: inst = 32'h24612800;
      71901: inst = 32'h10a0ffff;
      71902: inst = 32'hca0fffb;
      71903: inst = 32'h24822800;
      71904: inst = 32'h10a00000;
      71905: inst = 32'hca00004;
      71906: inst = 32'h38632800;
      71907: inst = 32'h38842800;
      71908: inst = 32'h10a00001;
      71909: inst = 32'hca018e9;
      71910: inst = 32'h13e00001;
      71911: inst = 32'hfe0d96a;
      71912: inst = 32'h5be00000;
      71913: inst = 32'h8c50000;
      71914: inst = 32'h24612800;
      71915: inst = 32'h10a0ffff;
      71916: inst = 32'hca0fffb;
      71917: inst = 32'h24822800;
      71918: inst = 32'h10a00000;
      71919: inst = 32'hca00004;
      71920: inst = 32'h38632800;
      71921: inst = 32'h38842800;
      71922: inst = 32'h10a00001;
      71923: inst = 32'hca018f7;
      71924: inst = 32'h13e00001;
      71925: inst = 32'hfe0d96a;
      71926: inst = 32'h5be00000;
      71927: inst = 32'h8c50000;
      71928: inst = 32'h24612800;
      71929: inst = 32'h10a0ffff;
      71930: inst = 32'hca0fffb;
      71931: inst = 32'h24822800;
      71932: inst = 32'h10a00000;
      71933: inst = 32'hca00004;
      71934: inst = 32'h38632800;
      71935: inst = 32'h38842800;
      71936: inst = 32'h10a00001;
      71937: inst = 32'hca01905;
      71938: inst = 32'h13e00001;
      71939: inst = 32'hfe0d96a;
      71940: inst = 32'h5be00000;
      71941: inst = 32'h8c50000;
      71942: inst = 32'h24612800;
      71943: inst = 32'h10a0ffff;
      71944: inst = 32'hca0fffb;
      71945: inst = 32'h24822800;
      71946: inst = 32'h10a00000;
      71947: inst = 32'hca00004;
      71948: inst = 32'h38632800;
      71949: inst = 32'h38842800;
      71950: inst = 32'h10a00001;
      71951: inst = 32'hca01913;
      71952: inst = 32'h13e00001;
      71953: inst = 32'hfe0d96a;
      71954: inst = 32'h5be00000;
      71955: inst = 32'h8c50000;
      71956: inst = 32'h24612800;
      71957: inst = 32'h10a0ffff;
      71958: inst = 32'hca0fffb;
      71959: inst = 32'h24822800;
      71960: inst = 32'h10a00000;
      71961: inst = 32'hca00004;
      71962: inst = 32'h38632800;
      71963: inst = 32'h38842800;
      71964: inst = 32'h10a00001;
      71965: inst = 32'hca01921;
      71966: inst = 32'h13e00001;
      71967: inst = 32'hfe0d96a;
      71968: inst = 32'h5be00000;
      71969: inst = 32'h8c50000;
      71970: inst = 32'h24612800;
      71971: inst = 32'h10a0ffff;
      71972: inst = 32'hca0fffb;
      71973: inst = 32'h24822800;
      71974: inst = 32'h10a00000;
      71975: inst = 32'hca00004;
      71976: inst = 32'h38632800;
      71977: inst = 32'h38842800;
      71978: inst = 32'h10a00001;
      71979: inst = 32'hca0192f;
      71980: inst = 32'h13e00001;
      71981: inst = 32'hfe0d96a;
      71982: inst = 32'h5be00000;
      71983: inst = 32'h8c50000;
      71984: inst = 32'h24612800;
      71985: inst = 32'h10a0ffff;
      71986: inst = 32'hca0fffb;
      71987: inst = 32'h24822800;
      71988: inst = 32'h10a00000;
      71989: inst = 32'hca00004;
      71990: inst = 32'h38632800;
      71991: inst = 32'h38842800;
      71992: inst = 32'h10a00001;
      71993: inst = 32'hca0193d;
      71994: inst = 32'h13e00001;
      71995: inst = 32'hfe0d96a;
      71996: inst = 32'h5be00000;
      71997: inst = 32'h8c50000;
      71998: inst = 32'h24612800;
      71999: inst = 32'h10a0ffff;
      72000: inst = 32'hca0fffb;
      72001: inst = 32'h24822800;
      72002: inst = 32'h10a00000;
      72003: inst = 32'hca00004;
      72004: inst = 32'h38632800;
      72005: inst = 32'h38842800;
      72006: inst = 32'h10a00001;
      72007: inst = 32'hca0194b;
      72008: inst = 32'h13e00001;
      72009: inst = 32'hfe0d96a;
      72010: inst = 32'h5be00000;
      72011: inst = 32'h8c50000;
      72012: inst = 32'h24612800;
      72013: inst = 32'h10a0ffff;
      72014: inst = 32'hca0fffb;
      72015: inst = 32'h24822800;
      72016: inst = 32'h10a00000;
      72017: inst = 32'hca00004;
      72018: inst = 32'h38632800;
      72019: inst = 32'h38842800;
      72020: inst = 32'h10a00001;
      72021: inst = 32'hca01959;
      72022: inst = 32'h13e00001;
      72023: inst = 32'hfe0d96a;
      72024: inst = 32'h5be00000;
      72025: inst = 32'h8c50000;
      72026: inst = 32'h24612800;
      72027: inst = 32'h10a0ffff;
      72028: inst = 32'hca0fffb;
      72029: inst = 32'h24822800;
      72030: inst = 32'h10a00000;
      72031: inst = 32'hca00004;
      72032: inst = 32'h38632800;
      72033: inst = 32'h38842800;
      72034: inst = 32'h10a00001;
      72035: inst = 32'hca01967;
      72036: inst = 32'h13e00001;
      72037: inst = 32'hfe0d96a;
      72038: inst = 32'h5be00000;
      72039: inst = 32'h8c50000;
      72040: inst = 32'h24612800;
      72041: inst = 32'h10a0ffff;
      72042: inst = 32'hca0fffb;
      72043: inst = 32'h24822800;
      72044: inst = 32'h10a00000;
      72045: inst = 32'hca00004;
      72046: inst = 32'h38632800;
      72047: inst = 32'h38842800;
      72048: inst = 32'h10a00001;
      72049: inst = 32'hca01975;
      72050: inst = 32'h13e00001;
      72051: inst = 32'hfe0d96a;
      72052: inst = 32'h5be00000;
      72053: inst = 32'h8c50000;
      72054: inst = 32'h24612800;
      72055: inst = 32'h10a0ffff;
      72056: inst = 32'hca0fffb;
      72057: inst = 32'h24822800;
      72058: inst = 32'h10a00000;
      72059: inst = 32'hca00004;
      72060: inst = 32'h38632800;
      72061: inst = 32'h38842800;
      72062: inst = 32'h10a00001;
      72063: inst = 32'hca01983;
      72064: inst = 32'h13e00001;
      72065: inst = 32'hfe0d96a;
      72066: inst = 32'h5be00000;
      72067: inst = 32'h8c50000;
      72068: inst = 32'h24612800;
      72069: inst = 32'h10a0ffff;
      72070: inst = 32'hca0fffb;
      72071: inst = 32'h24822800;
      72072: inst = 32'h10a00000;
      72073: inst = 32'hca00004;
      72074: inst = 32'h38632800;
      72075: inst = 32'h38842800;
      72076: inst = 32'h10a00001;
      72077: inst = 32'hca01991;
      72078: inst = 32'h13e00001;
      72079: inst = 32'hfe0d96a;
      72080: inst = 32'h5be00000;
      72081: inst = 32'h8c50000;
      72082: inst = 32'h24612800;
      72083: inst = 32'h10a0ffff;
      72084: inst = 32'hca0fffb;
      72085: inst = 32'h24822800;
      72086: inst = 32'h10a00000;
      72087: inst = 32'hca00004;
      72088: inst = 32'h38632800;
      72089: inst = 32'h38842800;
      72090: inst = 32'h10a00001;
      72091: inst = 32'hca0199f;
      72092: inst = 32'h13e00001;
      72093: inst = 32'hfe0d96a;
      72094: inst = 32'h5be00000;
      72095: inst = 32'h8c50000;
      72096: inst = 32'h24612800;
      72097: inst = 32'h10a0ffff;
      72098: inst = 32'hca0fffb;
      72099: inst = 32'h24822800;
      72100: inst = 32'h10a00000;
      72101: inst = 32'hca00004;
      72102: inst = 32'h38632800;
      72103: inst = 32'h38842800;
      72104: inst = 32'h10a00001;
      72105: inst = 32'hca019ad;
      72106: inst = 32'h13e00001;
      72107: inst = 32'hfe0d96a;
      72108: inst = 32'h5be00000;
      72109: inst = 32'h8c50000;
      72110: inst = 32'h24612800;
      72111: inst = 32'h10a0ffff;
      72112: inst = 32'hca0fffb;
      72113: inst = 32'h24822800;
      72114: inst = 32'h10a00000;
      72115: inst = 32'hca00004;
      72116: inst = 32'h38632800;
      72117: inst = 32'h38842800;
      72118: inst = 32'h10a00001;
      72119: inst = 32'hca019bb;
      72120: inst = 32'h13e00001;
      72121: inst = 32'hfe0d96a;
      72122: inst = 32'h5be00000;
      72123: inst = 32'h8c50000;
      72124: inst = 32'h24612800;
      72125: inst = 32'h10a0ffff;
      72126: inst = 32'hca0fffb;
      72127: inst = 32'h24822800;
      72128: inst = 32'h10a00000;
      72129: inst = 32'hca00004;
      72130: inst = 32'h38632800;
      72131: inst = 32'h38842800;
      72132: inst = 32'h10a00001;
      72133: inst = 32'hca019c9;
      72134: inst = 32'h13e00001;
      72135: inst = 32'hfe0d96a;
      72136: inst = 32'h5be00000;
      72137: inst = 32'h8c50000;
      72138: inst = 32'h24612800;
      72139: inst = 32'h10a0ffff;
      72140: inst = 32'hca0fffb;
      72141: inst = 32'h24822800;
      72142: inst = 32'h10a00000;
      72143: inst = 32'hca00004;
      72144: inst = 32'h38632800;
      72145: inst = 32'h38842800;
      72146: inst = 32'h10a00001;
      72147: inst = 32'hca019d7;
      72148: inst = 32'h13e00001;
      72149: inst = 32'hfe0d96a;
      72150: inst = 32'h5be00000;
      72151: inst = 32'h8c50000;
      72152: inst = 32'h24612800;
      72153: inst = 32'h10a0ffff;
      72154: inst = 32'hca0fffb;
      72155: inst = 32'h24822800;
      72156: inst = 32'h10a00000;
      72157: inst = 32'hca00004;
      72158: inst = 32'h38632800;
      72159: inst = 32'h38842800;
      72160: inst = 32'h10a00001;
      72161: inst = 32'hca019e5;
      72162: inst = 32'h13e00001;
      72163: inst = 32'hfe0d96a;
      72164: inst = 32'h5be00000;
      72165: inst = 32'h8c50000;
      72166: inst = 32'h24612800;
      72167: inst = 32'h10a0ffff;
      72168: inst = 32'hca0fffb;
      72169: inst = 32'h24822800;
      72170: inst = 32'h10a00000;
      72171: inst = 32'hca00004;
      72172: inst = 32'h38632800;
      72173: inst = 32'h38842800;
      72174: inst = 32'h10a00001;
      72175: inst = 32'hca019f3;
      72176: inst = 32'h13e00001;
      72177: inst = 32'hfe0d96a;
      72178: inst = 32'h5be00000;
      72179: inst = 32'h8c50000;
      72180: inst = 32'h24612800;
      72181: inst = 32'h10a0ffff;
      72182: inst = 32'hca0fffb;
      72183: inst = 32'h24822800;
      72184: inst = 32'h10a00000;
      72185: inst = 32'hca00004;
      72186: inst = 32'h38632800;
      72187: inst = 32'h38842800;
      72188: inst = 32'h10a00001;
      72189: inst = 32'hca01a01;
      72190: inst = 32'h13e00001;
      72191: inst = 32'hfe0d96a;
      72192: inst = 32'h5be00000;
      72193: inst = 32'h8c50000;
      72194: inst = 32'h24612800;
      72195: inst = 32'h10a0ffff;
      72196: inst = 32'hca0fffb;
      72197: inst = 32'h24822800;
      72198: inst = 32'h10a00000;
      72199: inst = 32'hca00004;
      72200: inst = 32'h38632800;
      72201: inst = 32'h38842800;
      72202: inst = 32'h10a00001;
      72203: inst = 32'hca01a0f;
      72204: inst = 32'h13e00001;
      72205: inst = 32'hfe0d96a;
      72206: inst = 32'h5be00000;
      72207: inst = 32'h8c50000;
      72208: inst = 32'h24612800;
      72209: inst = 32'h10a0ffff;
      72210: inst = 32'hca0fffb;
      72211: inst = 32'h24822800;
      72212: inst = 32'h10a00000;
      72213: inst = 32'hca00004;
      72214: inst = 32'h38632800;
      72215: inst = 32'h38842800;
      72216: inst = 32'h10a00001;
      72217: inst = 32'hca01a1d;
      72218: inst = 32'h13e00001;
      72219: inst = 32'hfe0d96a;
      72220: inst = 32'h5be00000;
      72221: inst = 32'h8c50000;
      72222: inst = 32'h24612800;
      72223: inst = 32'h10a0ffff;
      72224: inst = 32'hca0fffb;
      72225: inst = 32'h24822800;
      72226: inst = 32'h10a00000;
      72227: inst = 32'hca00004;
      72228: inst = 32'h38632800;
      72229: inst = 32'h38842800;
      72230: inst = 32'h10a00001;
      72231: inst = 32'hca01a2b;
      72232: inst = 32'h13e00001;
      72233: inst = 32'hfe0d96a;
      72234: inst = 32'h5be00000;
      72235: inst = 32'h8c50000;
      72236: inst = 32'h24612800;
      72237: inst = 32'h10a0ffff;
      72238: inst = 32'hca0fffb;
      72239: inst = 32'h24822800;
      72240: inst = 32'h10a00000;
      72241: inst = 32'hca00004;
      72242: inst = 32'h38632800;
      72243: inst = 32'h38842800;
      72244: inst = 32'h10a00001;
      72245: inst = 32'hca01a39;
      72246: inst = 32'h13e00001;
      72247: inst = 32'hfe0d96a;
      72248: inst = 32'h5be00000;
      72249: inst = 32'h8c50000;
      72250: inst = 32'h24612800;
      72251: inst = 32'h10a0ffff;
      72252: inst = 32'hca0fffb;
      72253: inst = 32'h24822800;
      72254: inst = 32'h10a00000;
      72255: inst = 32'hca00004;
      72256: inst = 32'h38632800;
      72257: inst = 32'h38842800;
      72258: inst = 32'h10a00001;
      72259: inst = 32'hca01a47;
      72260: inst = 32'h13e00001;
      72261: inst = 32'hfe0d96a;
      72262: inst = 32'h5be00000;
      72263: inst = 32'h8c50000;
      72264: inst = 32'h24612800;
      72265: inst = 32'h10a0ffff;
      72266: inst = 32'hca0fffb;
      72267: inst = 32'h24822800;
      72268: inst = 32'h10a00000;
      72269: inst = 32'hca00004;
      72270: inst = 32'h38632800;
      72271: inst = 32'h38842800;
      72272: inst = 32'h10a00001;
      72273: inst = 32'hca01a55;
      72274: inst = 32'h13e00001;
      72275: inst = 32'hfe0d96a;
      72276: inst = 32'h5be00000;
      72277: inst = 32'h8c50000;
      72278: inst = 32'h24612800;
      72279: inst = 32'h10a0ffff;
      72280: inst = 32'hca0fffb;
      72281: inst = 32'h24822800;
      72282: inst = 32'h10a00000;
      72283: inst = 32'hca00004;
      72284: inst = 32'h38632800;
      72285: inst = 32'h38842800;
      72286: inst = 32'h10a00001;
      72287: inst = 32'hca01a63;
      72288: inst = 32'h13e00001;
      72289: inst = 32'hfe0d96a;
      72290: inst = 32'h5be00000;
      72291: inst = 32'h8c50000;
      72292: inst = 32'h24612800;
      72293: inst = 32'h10a0ffff;
      72294: inst = 32'hca0fffb;
      72295: inst = 32'h24822800;
      72296: inst = 32'h10a00000;
      72297: inst = 32'hca00004;
      72298: inst = 32'h38632800;
      72299: inst = 32'h38842800;
      72300: inst = 32'h10a00001;
      72301: inst = 32'hca01a71;
      72302: inst = 32'h13e00001;
      72303: inst = 32'hfe0d96a;
      72304: inst = 32'h5be00000;
      72305: inst = 32'h8c50000;
      72306: inst = 32'h24612800;
      72307: inst = 32'h10a0ffff;
      72308: inst = 32'hca0fffb;
      72309: inst = 32'h24822800;
      72310: inst = 32'h10a00000;
      72311: inst = 32'hca00004;
      72312: inst = 32'h38632800;
      72313: inst = 32'h38842800;
      72314: inst = 32'h10a00001;
      72315: inst = 32'hca01a7f;
      72316: inst = 32'h13e00001;
      72317: inst = 32'hfe0d96a;
      72318: inst = 32'h5be00000;
      72319: inst = 32'h8c50000;
      72320: inst = 32'h24612800;
      72321: inst = 32'h10a0ffff;
      72322: inst = 32'hca0fffb;
      72323: inst = 32'h24822800;
      72324: inst = 32'h10a00000;
      72325: inst = 32'hca00004;
      72326: inst = 32'h38632800;
      72327: inst = 32'h38842800;
      72328: inst = 32'h10a00001;
      72329: inst = 32'hca01a8d;
      72330: inst = 32'h13e00001;
      72331: inst = 32'hfe0d96a;
      72332: inst = 32'h5be00000;
      72333: inst = 32'h8c50000;
      72334: inst = 32'h24612800;
      72335: inst = 32'h10a0ffff;
      72336: inst = 32'hca0fffb;
      72337: inst = 32'h24822800;
      72338: inst = 32'h10a00000;
      72339: inst = 32'hca00004;
      72340: inst = 32'h38632800;
      72341: inst = 32'h38842800;
      72342: inst = 32'h10a00001;
      72343: inst = 32'hca01a9b;
      72344: inst = 32'h13e00001;
      72345: inst = 32'hfe0d96a;
      72346: inst = 32'h5be00000;
      72347: inst = 32'h8c50000;
      72348: inst = 32'h24612800;
      72349: inst = 32'h10a0ffff;
      72350: inst = 32'hca0fffb;
      72351: inst = 32'h24822800;
      72352: inst = 32'h10a00000;
      72353: inst = 32'hca00004;
      72354: inst = 32'h38632800;
      72355: inst = 32'h38842800;
      72356: inst = 32'h10a00001;
      72357: inst = 32'hca01aa9;
      72358: inst = 32'h13e00001;
      72359: inst = 32'hfe0d96a;
      72360: inst = 32'h5be00000;
      72361: inst = 32'h8c50000;
      72362: inst = 32'h24612800;
      72363: inst = 32'h10a0ffff;
      72364: inst = 32'hca0fffb;
      72365: inst = 32'h24822800;
      72366: inst = 32'h10a00000;
      72367: inst = 32'hca00004;
      72368: inst = 32'h38632800;
      72369: inst = 32'h38842800;
      72370: inst = 32'h10a00001;
      72371: inst = 32'hca01ab7;
      72372: inst = 32'h13e00001;
      72373: inst = 32'hfe0d96a;
      72374: inst = 32'h5be00000;
      72375: inst = 32'h8c50000;
      72376: inst = 32'h24612800;
      72377: inst = 32'h10a0ffff;
      72378: inst = 32'hca0fffb;
      72379: inst = 32'h24822800;
      72380: inst = 32'h10a00000;
      72381: inst = 32'hca00004;
      72382: inst = 32'h38632800;
      72383: inst = 32'h38842800;
      72384: inst = 32'h10a00001;
      72385: inst = 32'hca01ac5;
      72386: inst = 32'h13e00001;
      72387: inst = 32'hfe0d96a;
      72388: inst = 32'h5be00000;
      72389: inst = 32'h8c50000;
      72390: inst = 32'h24612800;
      72391: inst = 32'h10a0ffff;
      72392: inst = 32'hca0fffb;
      72393: inst = 32'h24822800;
      72394: inst = 32'h10a00000;
      72395: inst = 32'hca00004;
      72396: inst = 32'h38632800;
      72397: inst = 32'h38842800;
      72398: inst = 32'h10a00001;
      72399: inst = 32'hca01ad3;
      72400: inst = 32'h13e00001;
      72401: inst = 32'hfe0d96a;
      72402: inst = 32'h5be00000;
      72403: inst = 32'h8c50000;
      72404: inst = 32'h24612800;
      72405: inst = 32'h10a0ffff;
      72406: inst = 32'hca0fffb;
      72407: inst = 32'h24822800;
      72408: inst = 32'h10a00000;
      72409: inst = 32'hca00004;
      72410: inst = 32'h38632800;
      72411: inst = 32'h38842800;
      72412: inst = 32'h10a00001;
      72413: inst = 32'hca01ae1;
      72414: inst = 32'h13e00001;
      72415: inst = 32'hfe0d96a;
      72416: inst = 32'h5be00000;
      72417: inst = 32'h8c50000;
      72418: inst = 32'h24612800;
      72419: inst = 32'h10a0ffff;
      72420: inst = 32'hca0fffb;
      72421: inst = 32'h24822800;
      72422: inst = 32'h10a00000;
      72423: inst = 32'hca00004;
      72424: inst = 32'h38632800;
      72425: inst = 32'h38842800;
      72426: inst = 32'h10a00001;
      72427: inst = 32'hca01aef;
      72428: inst = 32'h13e00001;
      72429: inst = 32'hfe0d96a;
      72430: inst = 32'h5be00000;
      72431: inst = 32'h8c50000;
      72432: inst = 32'h24612800;
      72433: inst = 32'h10a0ffff;
      72434: inst = 32'hca0fffb;
      72435: inst = 32'h24822800;
      72436: inst = 32'h10a00000;
      72437: inst = 32'hca00004;
      72438: inst = 32'h38632800;
      72439: inst = 32'h38842800;
      72440: inst = 32'h10a00001;
      72441: inst = 32'hca01afd;
      72442: inst = 32'h13e00001;
      72443: inst = 32'hfe0d96a;
      72444: inst = 32'h5be00000;
      72445: inst = 32'h8c50000;
      72446: inst = 32'h24612800;
      72447: inst = 32'h10a0ffff;
      72448: inst = 32'hca0fffb;
      72449: inst = 32'h24822800;
      72450: inst = 32'h10a00000;
      72451: inst = 32'hca00004;
      72452: inst = 32'h38632800;
      72453: inst = 32'h38842800;
      72454: inst = 32'h10a00001;
      72455: inst = 32'hca01b0b;
      72456: inst = 32'h13e00001;
      72457: inst = 32'hfe0d96a;
      72458: inst = 32'h5be00000;
      72459: inst = 32'h8c50000;
      72460: inst = 32'h24612800;
      72461: inst = 32'h10a0ffff;
      72462: inst = 32'hca0fffb;
      72463: inst = 32'h24822800;
      72464: inst = 32'h10a00000;
      72465: inst = 32'hca00004;
      72466: inst = 32'h38632800;
      72467: inst = 32'h38842800;
      72468: inst = 32'h10a00001;
      72469: inst = 32'hca01b19;
      72470: inst = 32'h13e00001;
      72471: inst = 32'hfe0d96a;
      72472: inst = 32'h5be00000;
      72473: inst = 32'h8c50000;
      72474: inst = 32'h24612800;
      72475: inst = 32'h10a0ffff;
      72476: inst = 32'hca0fffb;
      72477: inst = 32'h24822800;
      72478: inst = 32'h10a00000;
      72479: inst = 32'hca00004;
      72480: inst = 32'h38632800;
      72481: inst = 32'h38842800;
      72482: inst = 32'h10a00001;
      72483: inst = 32'hca01b27;
      72484: inst = 32'h13e00001;
      72485: inst = 32'hfe0d96a;
      72486: inst = 32'h5be00000;
      72487: inst = 32'h8c50000;
      72488: inst = 32'h24612800;
      72489: inst = 32'h10a0ffff;
      72490: inst = 32'hca0fffb;
      72491: inst = 32'h24822800;
      72492: inst = 32'h10a00000;
      72493: inst = 32'hca00004;
      72494: inst = 32'h38632800;
      72495: inst = 32'h38842800;
      72496: inst = 32'h10a00001;
      72497: inst = 32'hca01b35;
      72498: inst = 32'h13e00001;
      72499: inst = 32'hfe0d96a;
      72500: inst = 32'h5be00000;
      72501: inst = 32'h8c50000;
      72502: inst = 32'h24612800;
      72503: inst = 32'h10a0ffff;
      72504: inst = 32'hca0fffb;
      72505: inst = 32'h24822800;
      72506: inst = 32'h10a00000;
      72507: inst = 32'hca00004;
      72508: inst = 32'h38632800;
      72509: inst = 32'h38842800;
      72510: inst = 32'h10a00001;
      72511: inst = 32'hca01b43;
      72512: inst = 32'h13e00001;
      72513: inst = 32'hfe0d96a;
      72514: inst = 32'h5be00000;
      72515: inst = 32'h8c50000;
      72516: inst = 32'h24612800;
      72517: inst = 32'h10a0ffff;
      72518: inst = 32'hca0fffb;
      72519: inst = 32'h24822800;
      72520: inst = 32'h10a00000;
      72521: inst = 32'hca00004;
      72522: inst = 32'h38632800;
      72523: inst = 32'h38842800;
      72524: inst = 32'h10a00001;
      72525: inst = 32'hca01b51;
      72526: inst = 32'h13e00001;
      72527: inst = 32'hfe0d96a;
      72528: inst = 32'h5be00000;
      72529: inst = 32'h8c50000;
      72530: inst = 32'h24612800;
      72531: inst = 32'h10a0ffff;
      72532: inst = 32'hca0fffb;
      72533: inst = 32'h24822800;
      72534: inst = 32'h10a00000;
      72535: inst = 32'hca00004;
      72536: inst = 32'h38632800;
      72537: inst = 32'h38842800;
      72538: inst = 32'h10a00001;
      72539: inst = 32'hca01b5f;
      72540: inst = 32'h13e00001;
      72541: inst = 32'hfe0d96a;
      72542: inst = 32'h5be00000;
      72543: inst = 32'h8c50000;
      72544: inst = 32'h24612800;
      72545: inst = 32'h10a0ffff;
      72546: inst = 32'hca0fffb;
      72547: inst = 32'h24822800;
      72548: inst = 32'h10a00000;
      72549: inst = 32'hca00004;
      72550: inst = 32'h38632800;
      72551: inst = 32'h38842800;
      72552: inst = 32'h10a00001;
      72553: inst = 32'hca01b6d;
      72554: inst = 32'h13e00001;
      72555: inst = 32'hfe0d96a;
      72556: inst = 32'h5be00000;
      72557: inst = 32'h8c50000;
      72558: inst = 32'h24612800;
      72559: inst = 32'h10a0ffff;
      72560: inst = 32'hca0fffb;
      72561: inst = 32'h24822800;
      72562: inst = 32'h10a00000;
      72563: inst = 32'hca00004;
      72564: inst = 32'h38632800;
      72565: inst = 32'h38842800;
      72566: inst = 32'h10a00001;
      72567: inst = 32'hca01b7b;
      72568: inst = 32'h13e00001;
      72569: inst = 32'hfe0d96a;
      72570: inst = 32'h5be00000;
      72571: inst = 32'h8c50000;
      72572: inst = 32'h24612800;
      72573: inst = 32'h10a0ffff;
      72574: inst = 32'hca0fffb;
      72575: inst = 32'h24822800;
      72576: inst = 32'h10a00000;
      72577: inst = 32'hca00004;
      72578: inst = 32'h38632800;
      72579: inst = 32'h38842800;
      72580: inst = 32'h10a00001;
      72581: inst = 32'hca01b89;
      72582: inst = 32'h13e00001;
      72583: inst = 32'hfe0d96a;
      72584: inst = 32'h5be00000;
      72585: inst = 32'h8c50000;
      72586: inst = 32'h24612800;
      72587: inst = 32'h10a0ffff;
      72588: inst = 32'hca0fffb;
      72589: inst = 32'h24822800;
      72590: inst = 32'h10a00000;
      72591: inst = 32'hca00004;
      72592: inst = 32'h38632800;
      72593: inst = 32'h38842800;
      72594: inst = 32'h10a00001;
      72595: inst = 32'hca01b97;
      72596: inst = 32'h13e00001;
      72597: inst = 32'hfe0d96a;
      72598: inst = 32'h5be00000;
      72599: inst = 32'h8c50000;
      72600: inst = 32'h24612800;
      72601: inst = 32'h10a0ffff;
      72602: inst = 32'hca0fffb;
      72603: inst = 32'h24822800;
      72604: inst = 32'h10a00000;
      72605: inst = 32'hca00004;
      72606: inst = 32'h38632800;
      72607: inst = 32'h38842800;
      72608: inst = 32'h10a00001;
      72609: inst = 32'hca01ba5;
      72610: inst = 32'h13e00001;
      72611: inst = 32'hfe0d96a;
      72612: inst = 32'h5be00000;
      72613: inst = 32'h8c50000;
      72614: inst = 32'h24612800;
      72615: inst = 32'h10a0ffff;
      72616: inst = 32'hca0fffb;
      72617: inst = 32'h24822800;
      72618: inst = 32'h10a00000;
      72619: inst = 32'hca00004;
      72620: inst = 32'h38632800;
      72621: inst = 32'h38842800;
      72622: inst = 32'h10a00001;
      72623: inst = 32'hca01bb3;
      72624: inst = 32'h13e00001;
      72625: inst = 32'hfe0d96a;
      72626: inst = 32'h5be00000;
      72627: inst = 32'h8c50000;
      72628: inst = 32'h24612800;
      72629: inst = 32'h10a0ffff;
      72630: inst = 32'hca0fffb;
      72631: inst = 32'h24822800;
      72632: inst = 32'h10a00000;
      72633: inst = 32'hca00004;
      72634: inst = 32'h38632800;
      72635: inst = 32'h38842800;
      72636: inst = 32'h10a00001;
      72637: inst = 32'hca01bc1;
      72638: inst = 32'h13e00001;
      72639: inst = 32'hfe0d96a;
      72640: inst = 32'h5be00000;
      72641: inst = 32'h8c50000;
      72642: inst = 32'h24612800;
      72643: inst = 32'h10a0ffff;
      72644: inst = 32'hca0fffb;
      72645: inst = 32'h24822800;
      72646: inst = 32'h10a00000;
      72647: inst = 32'hca00004;
      72648: inst = 32'h38632800;
      72649: inst = 32'h38842800;
      72650: inst = 32'h10a00001;
      72651: inst = 32'hca01bcf;
      72652: inst = 32'h13e00001;
      72653: inst = 32'hfe0d96a;
      72654: inst = 32'h5be00000;
      72655: inst = 32'h8c50000;
      72656: inst = 32'h24612800;
      72657: inst = 32'h10a0ffff;
      72658: inst = 32'hca0fffb;
      72659: inst = 32'h24822800;
      72660: inst = 32'h10a00000;
      72661: inst = 32'hca00004;
      72662: inst = 32'h38632800;
      72663: inst = 32'h38842800;
      72664: inst = 32'h10a00001;
      72665: inst = 32'hca01bdd;
      72666: inst = 32'h13e00001;
      72667: inst = 32'hfe0d96a;
      72668: inst = 32'h5be00000;
      72669: inst = 32'h8c50000;
      72670: inst = 32'h24612800;
      72671: inst = 32'h10a0ffff;
      72672: inst = 32'hca0fffb;
      72673: inst = 32'h24822800;
      72674: inst = 32'h10a00000;
      72675: inst = 32'hca00004;
      72676: inst = 32'h38632800;
      72677: inst = 32'h38842800;
      72678: inst = 32'h10a00001;
      72679: inst = 32'hca01beb;
      72680: inst = 32'h13e00001;
      72681: inst = 32'hfe0d96a;
      72682: inst = 32'h5be00000;
      72683: inst = 32'h8c50000;
      72684: inst = 32'h24612800;
      72685: inst = 32'h10a0ffff;
      72686: inst = 32'hca0fffb;
      72687: inst = 32'h24822800;
      72688: inst = 32'h10a00000;
      72689: inst = 32'hca00004;
      72690: inst = 32'h38632800;
      72691: inst = 32'h38842800;
      72692: inst = 32'h10a00001;
      72693: inst = 32'hca01bf9;
      72694: inst = 32'h13e00001;
      72695: inst = 32'hfe0d96a;
      72696: inst = 32'h5be00000;
      72697: inst = 32'h8c50000;
      72698: inst = 32'h24612800;
      72699: inst = 32'h10a0ffff;
      72700: inst = 32'hca0fffb;
      72701: inst = 32'h24822800;
      72702: inst = 32'h10a00000;
      72703: inst = 32'hca00004;
      72704: inst = 32'h38632800;
      72705: inst = 32'h38842800;
      72706: inst = 32'h10a00001;
      72707: inst = 32'hca01c07;
      72708: inst = 32'h13e00001;
      72709: inst = 32'hfe0d96a;
      72710: inst = 32'h5be00000;
      72711: inst = 32'h8c50000;
      72712: inst = 32'h24612800;
      72713: inst = 32'h10a0ffff;
      72714: inst = 32'hca0fffb;
      72715: inst = 32'h24822800;
      72716: inst = 32'h10a00000;
      72717: inst = 32'hca00004;
      72718: inst = 32'h38632800;
      72719: inst = 32'h38842800;
      72720: inst = 32'h10a00001;
      72721: inst = 32'hca01c15;
      72722: inst = 32'h13e00001;
      72723: inst = 32'hfe0d96a;
      72724: inst = 32'h5be00000;
      72725: inst = 32'h8c50000;
      72726: inst = 32'h24612800;
      72727: inst = 32'h10a0ffff;
      72728: inst = 32'hca0fffb;
      72729: inst = 32'h24822800;
      72730: inst = 32'h10a00000;
      72731: inst = 32'hca00004;
      72732: inst = 32'h38632800;
      72733: inst = 32'h38842800;
      72734: inst = 32'h10a00001;
      72735: inst = 32'hca01c23;
      72736: inst = 32'h13e00001;
      72737: inst = 32'hfe0d96a;
      72738: inst = 32'h5be00000;
      72739: inst = 32'h8c50000;
      72740: inst = 32'h24612800;
      72741: inst = 32'h10a0ffff;
      72742: inst = 32'hca0fffb;
      72743: inst = 32'h24822800;
      72744: inst = 32'h10a00000;
      72745: inst = 32'hca00004;
      72746: inst = 32'h38632800;
      72747: inst = 32'h38842800;
      72748: inst = 32'h10a00001;
      72749: inst = 32'hca01c31;
      72750: inst = 32'h13e00001;
      72751: inst = 32'hfe0d96a;
      72752: inst = 32'h5be00000;
      72753: inst = 32'h8c50000;
      72754: inst = 32'h24612800;
      72755: inst = 32'h10a0ffff;
      72756: inst = 32'hca0fffb;
      72757: inst = 32'h24822800;
      72758: inst = 32'h10a00000;
      72759: inst = 32'hca00004;
      72760: inst = 32'h38632800;
      72761: inst = 32'h38842800;
      72762: inst = 32'h10a00001;
      72763: inst = 32'hca01c3f;
      72764: inst = 32'h13e00001;
      72765: inst = 32'hfe0d96a;
      72766: inst = 32'h5be00000;
      72767: inst = 32'h8c50000;
      72768: inst = 32'h24612800;
      72769: inst = 32'h10a0ffff;
      72770: inst = 32'hca0fffb;
      72771: inst = 32'h24822800;
      72772: inst = 32'h10a00000;
      72773: inst = 32'hca00004;
      72774: inst = 32'h38632800;
      72775: inst = 32'h38842800;
      72776: inst = 32'h10a00001;
      72777: inst = 32'hca01c4d;
      72778: inst = 32'h13e00001;
      72779: inst = 32'hfe0d96a;
      72780: inst = 32'h5be00000;
      72781: inst = 32'h8c50000;
      72782: inst = 32'h24612800;
      72783: inst = 32'h10a0ffff;
      72784: inst = 32'hca0fffb;
      72785: inst = 32'h24822800;
      72786: inst = 32'h10a00000;
      72787: inst = 32'hca00004;
      72788: inst = 32'h38632800;
      72789: inst = 32'h38842800;
      72790: inst = 32'h10a00001;
      72791: inst = 32'hca01c5b;
      72792: inst = 32'h13e00001;
      72793: inst = 32'hfe0d96a;
      72794: inst = 32'h5be00000;
      72795: inst = 32'h8c50000;
      72796: inst = 32'h24612800;
      72797: inst = 32'h10a0ffff;
      72798: inst = 32'hca0fffb;
      72799: inst = 32'h24822800;
      72800: inst = 32'h10a00000;
      72801: inst = 32'hca00004;
      72802: inst = 32'h38632800;
      72803: inst = 32'h38842800;
      72804: inst = 32'h10a00001;
      72805: inst = 32'hca01c69;
      72806: inst = 32'h13e00001;
      72807: inst = 32'hfe0d96a;
      72808: inst = 32'h5be00000;
      72809: inst = 32'h8c50000;
      72810: inst = 32'h24612800;
      72811: inst = 32'h10a0ffff;
      72812: inst = 32'hca0fffc;
      72813: inst = 32'h24822800;
      72814: inst = 32'h10a00000;
      72815: inst = 32'hca00004;
      72816: inst = 32'h38632800;
      72817: inst = 32'h38842800;
      72818: inst = 32'h10a00001;
      72819: inst = 32'hca01c77;
      72820: inst = 32'h13e00001;
      72821: inst = 32'hfe0d96a;
      72822: inst = 32'h5be00000;
      72823: inst = 32'h8c50000;
      72824: inst = 32'h24612800;
      72825: inst = 32'h10a0ffff;
      72826: inst = 32'hca0fffc;
      72827: inst = 32'h24822800;
      72828: inst = 32'h10a00000;
      72829: inst = 32'hca00004;
      72830: inst = 32'h38632800;
      72831: inst = 32'h38842800;
      72832: inst = 32'h10a00001;
      72833: inst = 32'hca01c85;
      72834: inst = 32'h13e00001;
      72835: inst = 32'hfe0d96a;
      72836: inst = 32'h5be00000;
      72837: inst = 32'h8c50000;
      72838: inst = 32'h24612800;
      72839: inst = 32'h10a0ffff;
      72840: inst = 32'hca0fffc;
      72841: inst = 32'h24822800;
      72842: inst = 32'h10a00000;
      72843: inst = 32'hca00004;
      72844: inst = 32'h38632800;
      72845: inst = 32'h38842800;
      72846: inst = 32'h10a00001;
      72847: inst = 32'hca01c93;
      72848: inst = 32'h13e00001;
      72849: inst = 32'hfe0d96a;
      72850: inst = 32'h5be00000;
      72851: inst = 32'h8c50000;
      72852: inst = 32'h24612800;
      72853: inst = 32'h10a0ffff;
      72854: inst = 32'hca0fffc;
      72855: inst = 32'h24822800;
      72856: inst = 32'h10a00000;
      72857: inst = 32'hca00004;
      72858: inst = 32'h38632800;
      72859: inst = 32'h38842800;
      72860: inst = 32'h10a00001;
      72861: inst = 32'hca01ca1;
      72862: inst = 32'h13e00001;
      72863: inst = 32'hfe0d96a;
      72864: inst = 32'h5be00000;
      72865: inst = 32'h8c50000;
      72866: inst = 32'h24612800;
      72867: inst = 32'h10a0ffff;
      72868: inst = 32'hca0fffc;
      72869: inst = 32'h24822800;
      72870: inst = 32'h10a00000;
      72871: inst = 32'hca00004;
      72872: inst = 32'h38632800;
      72873: inst = 32'h38842800;
      72874: inst = 32'h10a00001;
      72875: inst = 32'hca01caf;
      72876: inst = 32'h13e00001;
      72877: inst = 32'hfe0d96a;
      72878: inst = 32'h5be00000;
      72879: inst = 32'h8c50000;
      72880: inst = 32'h24612800;
      72881: inst = 32'h10a0ffff;
      72882: inst = 32'hca0fffc;
      72883: inst = 32'h24822800;
      72884: inst = 32'h10a00000;
      72885: inst = 32'hca00004;
      72886: inst = 32'h38632800;
      72887: inst = 32'h38842800;
      72888: inst = 32'h10a00001;
      72889: inst = 32'hca01cbd;
      72890: inst = 32'h13e00001;
      72891: inst = 32'hfe0d96a;
      72892: inst = 32'h5be00000;
      72893: inst = 32'h8c50000;
      72894: inst = 32'h24612800;
      72895: inst = 32'h10a0ffff;
      72896: inst = 32'hca0fffc;
      72897: inst = 32'h24822800;
      72898: inst = 32'h10a00000;
      72899: inst = 32'hca00004;
      72900: inst = 32'h38632800;
      72901: inst = 32'h38842800;
      72902: inst = 32'h10a00001;
      72903: inst = 32'hca01ccb;
      72904: inst = 32'h13e00001;
      72905: inst = 32'hfe0d96a;
      72906: inst = 32'h5be00000;
      72907: inst = 32'h8c50000;
      72908: inst = 32'h24612800;
      72909: inst = 32'h10a0ffff;
      72910: inst = 32'hca0fffc;
      72911: inst = 32'h24822800;
      72912: inst = 32'h10a00000;
      72913: inst = 32'hca00004;
      72914: inst = 32'h38632800;
      72915: inst = 32'h38842800;
      72916: inst = 32'h10a00001;
      72917: inst = 32'hca01cd9;
      72918: inst = 32'h13e00001;
      72919: inst = 32'hfe0d96a;
      72920: inst = 32'h5be00000;
      72921: inst = 32'h8c50000;
      72922: inst = 32'h24612800;
      72923: inst = 32'h10a0ffff;
      72924: inst = 32'hca0fffc;
      72925: inst = 32'h24822800;
      72926: inst = 32'h10a00000;
      72927: inst = 32'hca00004;
      72928: inst = 32'h38632800;
      72929: inst = 32'h38842800;
      72930: inst = 32'h10a00001;
      72931: inst = 32'hca01ce7;
      72932: inst = 32'h13e00001;
      72933: inst = 32'hfe0d96a;
      72934: inst = 32'h5be00000;
      72935: inst = 32'h8c50000;
      72936: inst = 32'h24612800;
      72937: inst = 32'h10a0ffff;
      72938: inst = 32'hca0fffc;
      72939: inst = 32'h24822800;
      72940: inst = 32'h10a00000;
      72941: inst = 32'hca00004;
      72942: inst = 32'h38632800;
      72943: inst = 32'h38842800;
      72944: inst = 32'h10a00001;
      72945: inst = 32'hca01cf5;
      72946: inst = 32'h13e00001;
      72947: inst = 32'hfe0d96a;
      72948: inst = 32'h5be00000;
      72949: inst = 32'h8c50000;
      72950: inst = 32'h24612800;
      72951: inst = 32'h10a0ffff;
      72952: inst = 32'hca0fffc;
      72953: inst = 32'h24822800;
      72954: inst = 32'h10a00000;
      72955: inst = 32'hca00004;
      72956: inst = 32'h38632800;
      72957: inst = 32'h38842800;
      72958: inst = 32'h10a00001;
      72959: inst = 32'hca01d03;
      72960: inst = 32'h13e00001;
      72961: inst = 32'hfe0d96a;
      72962: inst = 32'h5be00000;
      72963: inst = 32'h8c50000;
      72964: inst = 32'h24612800;
      72965: inst = 32'h10a0ffff;
      72966: inst = 32'hca0fffc;
      72967: inst = 32'h24822800;
      72968: inst = 32'h10a00000;
      72969: inst = 32'hca00004;
      72970: inst = 32'h38632800;
      72971: inst = 32'h38842800;
      72972: inst = 32'h10a00001;
      72973: inst = 32'hca01d11;
      72974: inst = 32'h13e00001;
      72975: inst = 32'hfe0d96a;
      72976: inst = 32'h5be00000;
      72977: inst = 32'h8c50000;
      72978: inst = 32'h24612800;
      72979: inst = 32'h10a0ffff;
      72980: inst = 32'hca0fffc;
      72981: inst = 32'h24822800;
      72982: inst = 32'h10a00000;
      72983: inst = 32'hca00004;
      72984: inst = 32'h38632800;
      72985: inst = 32'h38842800;
      72986: inst = 32'h10a00001;
      72987: inst = 32'hca01d1f;
      72988: inst = 32'h13e00001;
      72989: inst = 32'hfe0d96a;
      72990: inst = 32'h5be00000;
      72991: inst = 32'h8c50000;
      72992: inst = 32'h24612800;
      72993: inst = 32'h10a0ffff;
      72994: inst = 32'hca0fffc;
      72995: inst = 32'h24822800;
      72996: inst = 32'h10a00000;
      72997: inst = 32'hca00004;
      72998: inst = 32'h38632800;
      72999: inst = 32'h38842800;
      73000: inst = 32'h10a00001;
      73001: inst = 32'hca01d2d;
      73002: inst = 32'h13e00001;
      73003: inst = 32'hfe0d96a;
      73004: inst = 32'h5be00000;
      73005: inst = 32'h8c50000;
      73006: inst = 32'h24612800;
      73007: inst = 32'h10a0ffff;
      73008: inst = 32'hca0fffc;
      73009: inst = 32'h24822800;
      73010: inst = 32'h10a00000;
      73011: inst = 32'hca00004;
      73012: inst = 32'h38632800;
      73013: inst = 32'h38842800;
      73014: inst = 32'h10a00001;
      73015: inst = 32'hca01d3b;
      73016: inst = 32'h13e00001;
      73017: inst = 32'hfe0d96a;
      73018: inst = 32'h5be00000;
      73019: inst = 32'h8c50000;
      73020: inst = 32'h24612800;
      73021: inst = 32'h10a0ffff;
      73022: inst = 32'hca0fffc;
      73023: inst = 32'h24822800;
      73024: inst = 32'h10a00000;
      73025: inst = 32'hca00004;
      73026: inst = 32'h38632800;
      73027: inst = 32'h38842800;
      73028: inst = 32'h10a00001;
      73029: inst = 32'hca01d49;
      73030: inst = 32'h13e00001;
      73031: inst = 32'hfe0d96a;
      73032: inst = 32'h5be00000;
      73033: inst = 32'h8c50000;
      73034: inst = 32'h24612800;
      73035: inst = 32'h10a0ffff;
      73036: inst = 32'hca0fffc;
      73037: inst = 32'h24822800;
      73038: inst = 32'h10a00000;
      73039: inst = 32'hca00004;
      73040: inst = 32'h38632800;
      73041: inst = 32'h38842800;
      73042: inst = 32'h10a00001;
      73043: inst = 32'hca01d57;
      73044: inst = 32'h13e00001;
      73045: inst = 32'hfe0d96a;
      73046: inst = 32'h5be00000;
      73047: inst = 32'h8c50000;
      73048: inst = 32'h24612800;
      73049: inst = 32'h10a0ffff;
      73050: inst = 32'hca0fffc;
      73051: inst = 32'h24822800;
      73052: inst = 32'h10a00000;
      73053: inst = 32'hca00004;
      73054: inst = 32'h38632800;
      73055: inst = 32'h38842800;
      73056: inst = 32'h10a00001;
      73057: inst = 32'hca01d65;
      73058: inst = 32'h13e00001;
      73059: inst = 32'hfe0d96a;
      73060: inst = 32'h5be00000;
      73061: inst = 32'h8c50000;
      73062: inst = 32'h24612800;
      73063: inst = 32'h10a0ffff;
      73064: inst = 32'hca0fffc;
      73065: inst = 32'h24822800;
      73066: inst = 32'h10a00000;
      73067: inst = 32'hca00004;
      73068: inst = 32'h38632800;
      73069: inst = 32'h38842800;
      73070: inst = 32'h10a00001;
      73071: inst = 32'hca01d73;
      73072: inst = 32'h13e00001;
      73073: inst = 32'hfe0d96a;
      73074: inst = 32'h5be00000;
      73075: inst = 32'h8c50000;
      73076: inst = 32'h24612800;
      73077: inst = 32'h10a0ffff;
      73078: inst = 32'hca0fffc;
      73079: inst = 32'h24822800;
      73080: inst = 32'h10a00000;
      73081: inst = 32'hca00004;
      73082: inst = 32'h38632800;
      73083: inst = 32'h38842800;
      73084: inst = 32'h10a00001;
      73085: inst = 32'hca01d81;
      73086: inst = 32'h13e00001;
      73087: inst = 32'hfe0d96a;
      73088: inst = 32'h5be00000;
      73089: inst = 32'h8c50000;
      73090: inst = 32'h24612800;
      73091: inst = 32'h10a0ffff;
      73092: inst = 32'hca0fffc;
      73093: inst = 32'h24822800;
      73094: inst = 32'h10a00000;
      73095: inst = 32'hca00004;
      73096: inst = 32'h38632800;
      73097: inst = 32'h38842800;
      73098: inst = 32'h10a00001;
      73099: inst = 32'hca01d8f;
      73100: inst = 32'h13e00001;
      73101: inst = 32'hfe0d96a;
      73102: inst = 32'h5be00000;
      73103: inst = 32'h8c50000;
      73104: inst = 32'h24612800;
      73105: inst = 32'h10a0ffff;
      73106: inst = 32'hca0fffc;
      73107: inst = 32'h24822800;
      73108: inst = 32'h10a00000;
      73109: inst = 32'hca00004;
      73110: inst = 32'h38632800;
      73111: inst = 32'h38842800;
      73112: inst = 32'h10a00001;
      73113: inst = 32'hca01d9d;
      73114: inst = 32'h13e00001;
      73115: inst = 32'hfe0d96a;
      73116: inst = 32'h5be00000;
      73117: inst = 32'h8c50000;
      73118: inst = 32'h24612800;
      73119: inst = 32'h10a0ffff;
      73120: inst = 32'hca0fffc;
      73121: inst = 32'h24822800;
      73122: inst = 32'h10a00000;
      73123: inst = 32'hca00004;
      73124: inst = 32'h38632800;
      73125: inst = 32'h38842800;
      73126: inst = 32'h10a00001;
      73127: inst = 32'hca01dab;
      73128: inst = 32'h13e00001;
      73129: inst = 32'hfe0d96a;
      73130: inst = 32'h5be00000;
      73131: inst = 32'h8c50000;
      73132: inst = 32'h24612800;
      73133: inst = 32'h10a0ffff;
      73134: inst = 32'hca0fffc;
      73135: inst = 32'h24822800;
      73136: inst = 32'h10a00000;
      73137: inst = 32'hca00004;
      73138: inst = 32'h38632800;
      73139: inst = 32'h38842800;
      73140: inst = 32'h10a00001;
      73141: inst = 32'hca01db9;
      73142: inst = 32'h13e00001;
      73143: inst = 32'hfe0d96a;
      73144: inst = 32'h5be00000;
      73145: inst = 32'h8c50000;
      73146: inst = 32'h24612800;
      73147: inst = 32'h10a0ffff;
      73148: inst = 32'hca0fffc;
      73149: inst = 32'h24822800;
      73150: inst = 32'h10a00000;
      73151: inst = 32'hca00004;
      73152: inst = 32'h38632800;
      73153: inst = 32'h38842800;
      73154: inst = 32'h10a00001;
      73155: inst = 32'hca01dc7;
      73156: inst = 32'h13e00001;
      73157: inst = 32'hfe0d96a;
      73158: inst = 32'h5be00000;
      73159: inst = 32'h8c50000;
      73160: inst = 32'h24612800;
      73161: inst = 32'h10a0ffff;
      73162: inst = 32'hca0fffc;
      73163: inst = 32'h24822800;
      73164: inst = 32'h10a00000;
      73165: inst = 32'hca00004;
      73166: inst = 32'h38632800;
      73167: inst = 32'h38842800;
      73168: inst = 32'h10a00001;
      73169: inst = 32'hca01dd5;
      73170: inst = 32'h13e00001;
      73171: inst = 32'hfe0d96a;
      73172: inst = 32'h5be00000;
      73173: inst = 32'h8c50000;
      73174: inst = 32'h24612800;
      73175: inst = 32'h10a0ffff;
      73176: inst = 32'hca0fffc;
      73177: inst = 32'h24822800;
      73178: inst = 32'h10a00000;
      73179: inst = 32'hca00004;
      73180: inst = 32'h38632800;
      73181: inst = 32'h38842800;
      73182: inst = 32'h10a00001;
      73183: inst = 32'hca01de3;
      73184: inst = 32'h13e00001;
      73185: inst = 32'hfe0d96a;
      73186: inst = 32'h5be00000;
      73187: inst = 32'h8c50000;
      73188: inst = 32'h24612800;
      73189: inst = 32'h10a0ffff;
      73190: inst = 32'hca0fffc;
      73191: inst = 32'h24822800;
      73192: inst = 32'h10a00000;
      73193: inst = 32'hca00004;
      73194: inst = 32'h38632800;
      73195: inst = 32'h38842800;
      73196: inst = 32'h10a00001;
      73197: inst = 32'hca01df1;
      73198: inst = 32'h13e00001;
      73199: inst = 32'hfe0d96a;
      73200: inst = 32'h5be00000;
      73201: inst = 32'h8c50000;
      73202: inst = 32'h24612800;
      73203: inst = 32'h10a0ffff;
      73204: inst = 32'hca0fffc;
      73205: inst = 32'h24822800;
      73206: inst = 32'h10a00000;
      73207: inst = 32'hca00004;
      73208: inst = 32'h38632800;
      73209: inst = 32'h38842800;
      73210: inst = 32'h10a00001;
      73211: inst = 32'hca01dff;
      73212: inst = 32'h13e00001;
      73213: inst = 32'hfe0d96a;
      73214: inst = 32'h5be00000;
      73215: inst = 32'h8c50000;
      73216: inst = 32'h24612800;
      73217: inst = 32'h10a0ffff;
      73218: inst = 32'hca0fffc;
      73219: inst = 32'h24822800;
      73220: inst = 32'h10a00000;
      73221: inst = 32'hca00004;
      73222: inst = 32'h38632800;
      73223: inst = 32'h38842800;
      73224: inst = 32'h10a00001;
      73225: inst = 32'hca01e0d;
      73226: inst = 32'h13e00001;
      73227: inst = 32'hfe0d96a;
      73228: inst = 32'h5be00000;
      73229: inst = 32'h8c50000;
      73230: inst = 32'h24612800;
      73231: inst = 32'h10a0ffff;
      73232: inst = 32'hca0fffc;
      73233: inst = 32'h24822800;
      73234: inst = 32'h10a00000;
      73235: inst = 32'hca00004;
      73236: inst = 32'h38632800;
      73237: inst = 32'h38842800;
      73238: inst = 32'h10a00001;
      73239: inst = 32'hca01e1b;
      73240: inst = 32'h13e00001;
      73241: inst = 32'hfe0d96a;
      73242: inst = 32'h5be00000;
      73243: inst = 32'h8c50000;
      73244: inst = 32'h24612800;
      73245: inst = 32'h10a0ffff;
      73246: inst = 32'hca0fffc;
      73247: inst = 32'h24822800;
      73248: inst = 32'h10a00000;
      73249: inst = 32'hca00004;
      73250: inst = 32'h38632800;
      73251: inst = 32'h38842800;
      73252: inst = 32'h10a00001;
      73253: inst = 32'hca01e29;
      73254: inst = 32'h13e00001;
      73255: inst = 32'hfe0d96a;
      73256: inst = 32'h5be00000;
      73257: inst = 32'h8c50000;
      73258: inst = 32'h24612800;
      73259: inst = 32'h10a0ffff;
      73260: inst = 32'hca0fffc;
      73261: inst = 32'h24822800;
      73262: inst = 32'h10a00000;
      73263: inst = 32'hca00004;
      73264: inst = 32'h38632800;
      73265: inst = 32'h38842800;
      73266: inst = 32'h10a00001;
      73267: inst = 32'hca01e37;
      73268: inst = 32'h13e00001;
      73269: inst = 32'hfe0d96a;
      73270: inst = 32'h5be00000;
      73271: inst = 32'h8c50000;
      73272: inst = 32'h24612800;
      73273: inst = 32'h10a0ffff;
      73274: inst = 32'hca0fffc;
      73275: inst = 32'h24822800;
      73276: inst = 32'h10a00000;
      73277: inst = 32'hca00004;
      73278: inst = 32'h38632800;
      73279: inst = 32'h38842800;
      73280: inst = 32'h10a00001;
      73281: inst = 32'hca01e45;
      73282: inst = 32'h13e00001;
      73283: inst = 32'hfe0d96a;
      73284: inst = 32'h5be00000;
      73285: inst = 32'h8c50000;
      73286: inst = 32'h24612800;
      73287: inst = 32'h10a0ffff;
      73288: inst = 32'hca0fffc;
      73289: inst = 32'h24822800;
      73290: inst = 32'h10a00000;
      73291: inst = 32'hca00004;
      73292: inst = 32'h38632800;
      73293: inst = 32'h38842800;
      73294: inst = 32'h10a00001;
      73295: inst = 32'hca01e53;
      73296: inst = 32'h13e00001;
      73297: inst = 32'hfe0d96a;
      73298: inst = 32'h5be00000;
      73299: inst = 32'h8c50000;
      73300: inst = 32'h24612800;
      73301: inst = 32'h10a0ffff;
      73302: inst = 32'hca0fffc;
      73303: inst = 32'h24822800;
      73304: inst = 32'h10a00000;
      73305: inst = 32'hca00004;
      73306: inst = 32'h38632800;
      73307: inst = 32'h38842800;
      73308: inst = 32'h10a00001;
      73309: inst = 32'hca01e61;
      73310: inst = 32'h13e00001;
      73311: inst = 32'hfe0d96a;
      73312: inst = 32'h5be00000;
      73313: inst = 32'h8c50000;
      73314: inst = 32'h24612800;
      73315: inst = 32'h10a0ffff;
      73316: inst = 32'hca0fffc;
      73317: inst = 32'h24822800;
      73318: inst = 32'h10a00000;
      73319: inst = 32'hca00004;
      73320: inst = 32'h38632800;
      73321: inst = 32'h38842800;
      73322: inst = 32'h10a00001;
      73323: inst = 32'hca01e6f;
      73324: inst = 32'h13e00001;
      73325: inst = 32'hfe0d96a;
      73326: inst = 32'h5be00000;
      73327: inst = 32'h8c50000;
      73328: inst = 32'h24612800;
      73329: inst = 32'h10a0ffff;
      73330: inst = 32'hca0fffc;
      73331: inst = 32'h24822800;
      73332: inst = 32'h10a00000;
      73333: inst = 32'hca00004;
      73334: inst = 32'h38632800;
      73335: inst = 32'h38842800;
      73336: inst = 32'h10a00001;
      73337: inst = 32'hca01e7d;
      73338: inst = 32'h13e00001;
      73339: inst = 32'hfe0d96a;
      73340: inst = 32'h5be00000;
      73341: inst = 32'h8c50000;
      73342: inst = 32'h24612800;
      73343: inst = 32'h10a0ffff;
      73344: inst = 32'hca0fffc;
      73345: inst = 32'h24822800;
      73346: inst = 32'h10a00000;
      73347: inst = 32'hca00004;
      73348: inst = 32'h38632800;
      73349: inst = 32'h38842800;
      73350: inst = 32'h10a00001;
      73351: inst = 32'hca01e8b;
      73352: inst = 32'h13e00001;
      73353: inst = 32'hfe0d96a;
      73354: inst = 32'h5be00000;
      73355: inst = 32'h8c50000;
      73356: inst = 32'h24612800;
      73357: inst = 32'h10a0ffff;
      73358: inst = 32'hca0fffc;
      73359: inst = 32'h24822800;
      73360: inst = 32'h10a00000;
      73361: inst = 32'hca00004;
      73362: inst = 32'h38632800;
      73363: inst = 32'h38842800;
      73364: inst = 32'h10a00001;
      73365: inst = 32'hca01e99;
      73366: inst = 32'h13e00001;
      73367: inst = 32'hfe0d96a;
      73368: inst = 32'h5be00000;
      73369: inst = 32'h8c50000;
      73370: inst = 32'h24612800;
      73371: inst = 32'h10a0ffff;
      73372: inst = 32'hca0fffc;
      73373: inst = 32'h24822800;
      73374: inst = 32'h10a00000;
      73375: inst = 32'hca00004;
      73376: inst = 32'h38632800;
      73377: inst = 32'h38842800;
      73378: inst = 32'h10a00001;
      73379: inst = 32'hca01ea7;
      73380: inst = 32'h13e00001;
      73381: inst = 32'hfe0d96a;
      73382: inst = 32'h5be00000;
      73383: inst = 32'h8c50000;
      73384: inst = 32'h24612800;
      73385: inst = 32'h10a0ffff;
      73386: inst = 32'hca0fffc;
      73387: inst = 32'h24822800;
      73388: inst = 32'h10a00000;
      73389: inst = 32'hca00004;
      73390: inst = 32'h38632800;
      73391: inst = 32'h38842800;
      73392: inst = 32'h10a00001;
      73393: inst = 32'hca01eb5;
      73394: inst = 32'h13e00001;
      73395: inst = 32'hfe0d96a;
      73396: inst = 32'h5be00000;
      73397: inst = 32'h8c50000;
      73398: inst = 32'h24612800;
      73399: inst = 32'h10a0ffff;
      73400: inst = 32'hca0fffc;
      73401: inst = 32'h24822800;
      73402: inst = 32'h10a00000;
      73403: inst = 32'hca00004;
      73404: inst = 32'h38632800;
      73405: inst = 32'h38842800;
      73406: inst = 32'h10a00001;
      73407: inst = 32'hca01ec3;
      73408: inst = 32'h13e00001;
      73409: inst = 32'hfe0d96a;
      73410: inst = 32'h5be00000;
      73411: inst = 32'h8c50000;
      73412: inst = 32'h24612800;
      73413: inst = 32'h10a0ffff;
      73414: inst = 32'hca0fffc;
      73415: inst = 32'h24822800;
      73416: inst = 32'h10a00000;
      73417: inst = 32'hca00004;
      73418: inst = 32'h38632800;
      73419: inst = 32'h38842800;
      73420: inst = 32'h10a00001;
      73421: inst = 32'hca01ed1;
      73422: inst = 32'h13e00001;
      73423: inst = 32'hfe0d96a;
      73424: inst = 32'h5be00000;
      73425: inst = 32'h8c50000;
      73426: inst = 32'h24612800;
      73427: inst = 32'h10a0ffff;
      73428: inst = 32'hca0fffc;
      73429: inst = 32'h24822800;
      73430: inst = 32'h10a00000;
      73431: inst = 32'hca00004;
      73432: inst = 32'h38632800;
      73433: inst = 32'h38842800;
      73434: inst = 32'h10a00001;
      73435: inst = 32'hca01edf;
      73436: inst = 32'h13e00001;
      73437: inst = 32'hfe0d96a;
      73438: inst = 32'h5be00000;
      73439: inst = 32'h8c50000;
      73440: inst = 32'h24612800;
      73441: inst = 32'h10a0ffff;
      73442: inst = 32'hca0fffc;
      73443: inst = 32'h24822800;
      73444: inst = 32'h10a00000;
      73445: inst = 32'hca00004;
      73446: inst = 32'h38632800;
      73447: inst = 32'h38842800;
      73448: inst = 32'h10a00001;
      73449: inst = 32'hca01eed;
      73450: inst = 32'h13e00001;
      73451: inst = 32'hfe0d96a;
      73452: inst = 32'h5be00000;
      73453: inst = 32'h8c50000;
      73454: inst = 32'h24612800;
      73455: inst = 32'h10a0ffff;
      73456: inst = 32'hca0fffc;
      73457: inst = 32'h24822800;
      73458: inst = 32'h10a00000;
      73459: inst = 32'hca00004;
      73460: inst = 32'h38632800;
      73461: inst = 32'h38842800;
      73462: inst = 32'h10a00001;
      73463: inst = 32'hca01efb;
      73464: inst = 32'h13e00001;
      73465: inst = 32'hfe0d96a;
      73466: inst = 32'h5be00000;
      73467: inst = 32'h8c50000;
      73468: inst = 32'h24612800;
      73469: inst = 32'h10a0ffff;
      73470: inst = 32'hca0fffc;
      73471: inst = 32'h24822800;
      73472: inst = 32'h10a00000;
      73473: inst = 32'hca00004;
      73474: inst = 32'h38632800;
      73475: inst = 32'h38842800;
      73476: inst = 32'h10a00001;
      73477: inst = 32'hca01f09;
      73478: inst = 32'h13e00001;
      73479: inst = 32'hfe0d96a;
      73480: inst = 32'h5be00000;
      73481: inst = 32'h8c50000;
      73482: inst = 32'h24612800;
      73483: inst = 32'h10a0ffff;
      73484: inst = 32'hca0fffc;
      73485: inst = 32'h24822800;
      73486: inst = 32'h10a00000;
      73487: inst = 32'hca00004;
      73488: inst = 32'h38632800;
      73489: inst = 32'h38842800;
      73490: inst = 32'h10a00001;
      73491: inst = 32'hca01f17;
      73492: inst = 32'h13e00001;
      73493: inst = 32'hfe0d96a;
      73494: inst = 32'h5be00000;
      73495: inst = 32'h8c50000;
      73496: inst = 32'h24612800;
      73497: inst = 32'h10a0ffff;
      73498: inst = 32'hca0fffc;
      73499: inst = 32'h24822800;
      73500: inst = 32'h10a00000;
      73501: inst = 32'hca00004;
      73502: inst = 32'h38632800;
      73503: inst = 32'h38842800;
      73504: inst = 32'h10a00001;
      73505: inst = 32'hca01f25;
      73506: inst = 32'h13e00001;
      73507: inst = 32'hfe0d96a;
      73508: inst = 32'h5be00000;
      73509: inst = 32'h8c50000;
      73510: inst = 32'h24612800;
      73511: inst = 32'h10a0ffff;
      73512: inst = 32'hca0fffc;
      73513: inst = 32'h24822800;
      73514: inst = 32'h10a00000;
      73515: inst = 32'hca00004;
      73516: inst = 32'h38632800;
      73517: inst = 32'h38842800;
      73518: inst = 32'h10a00001;
      73519: inst = 32'hca01f33;
      73520: inst = 32'h13e00001;
      73521: inst = 32'hfe0d96a;
      73522: inst = 32'h5be00000;
      73523: inst = 32'h8c50000;
      73524: inst = 32'h24612800;
      73525: inst = 32'h10a0ffff;
      73526: inst = 32'hca0fffc;
      73527: inst = 32'h24822800;
      73528: inst = 32'h10a00000;
      73529: inst = 32'hca00004;
      73530: inst = 32'h38632800;
      73531: inst = 32'h38842800;
      73532: inst = 32'h10a00001;
      73533: inst = 32'hca01f41;
      73534: inst = 32'h13e00001;
      73535: inst = 32'hfe0d96a;
      73536: inst = 32'h5be00000;
      73537: inst = 32'h8c50000;
      73538: inst = 32'h24612800;
      73539: inst = 32'h10a0ffff;
      73540: inst = 32'hca0fffc;
      73541: inst = 32'h24822800;
      73542: inst = 32'h10a00000;
      73543: inst = 32'hca00004;
      73544: inst = 32'h38632800;
      73545: inst = 32'h38842800;
      73546: inst = 32'h10a00001;
      73547: inst = 32'hca01f4f;
      73548: inst = 32'h13e00001;
      73549: inst = 32'hfe0d96a;
      73550: inst = 32'h5be00000;
      73551: inst = 32'h8c50000;
      73552: inst = 32'h24612800;
      73553: inst = 32'h10a0ffff;
      73554: inst = 32'hca0fffc;
      73555: inst = 32'h24822800;
      73556: inst = 32'h10a00000;
      73557: inst = 32'hca00004;
      73558: inst = 32'h38632800;
      73559: inst = 32'h38842800;
      73560: inst = 32'h10a00001;
      73561: inst = 32'hca01f5d;
      73562: inst = 32'h13e00001;
      73563: inst = 32'hfe0d96a;
      73564: inst = 32'h5be00000;
      73565: inst = 32'h8c50000;
      73566: inst = 32'h24612800;
      73567: inst = 32'h10a0ffff;
      73568: inst = 32'hca0fffc;
      73569: inst = 32'h24822800;
      73570: inst = 32'h10a00000;
      73571: inst = 32'hca00004;
      73572: inst = 32'h38632800;
      73573: inst = 32'h38842800;
      73574: inst = 32'h10a00001;
      73575: inst = 32'hca01f6b;
      73576: inst = 32'h13e00001;
      73577: inst = 32'hfe0d96a;
      73578: inst = 32'h5be00000;
      73579: inst = 32'h8c50000;
      73580: inst = 32'h24612800;
      73581: inst = 32'h10a0ffff;
      73582: inst = 32'hca0fffc;
      73583: inst = 32'h24822800;
      73584: inst = 32'h10a00000;
      73585: inst = 32'hca00004;
      73586: inst = 32'h38632800;
      73587: inst = 32'h38842800;
      73588: inst = 32'h10a00001;
      73589: inst = 32'hca01f79;
      73590: inst = 32'h13e00001;
      73591: inst = 32'hfe0d96a;
      73592: inst = 32'h5be00000;
      73593: inst = 32'h8c50000;
      73594: inst = 32'h24612800;
      73595: inst = 32'h10a0ffff;
      73596: inst = 32'hca0fffc;
      73597: inst = 32'h24822800;
      73598: inst = 32'h10a00000;
      73599: inst = 32'hca00004;
      73600: inst = 32'h38632800;
      73601: inst = 32'h38842800;
      73602: inst = 32'h10a00001;
      73603: inst = 32'hca01f87;
      73604: inst = 32'h13e00001;
      73605: inst = 32'hfe0d96a;
      73606: inst = 32'h5be00000;
      73607: inst = 32'h8c50000;
      73608: inst = 32'h24612800;
      73609: inst = 32'h10a0ffff;
      73610: inst = 32'hca0fffc;
      73611: inst = 32'h24822800;
      73612: inst = 32'h10a00000;
      73613: inst = 32'hca00004;
      73614: inst = 32'h38632800;
      73615: inst = 32'h38842800;
      73616: inst = 32'h10a00001;
      73617: inst = 32'hca01f95;
      73618: inst = 32'h13e00001;
      73619: inst = 32'hfe0d96a;
      73620: inst = 32'h5be00000;
      73621: inst = 32'h8c50000;
      73622: inst = 32'h24612800;
      73623: inst = 32'h10a0ffff;
      73624: inst = 32'hca0fffc;
      73625: inst = 32'h24822800;
      73626: inst = 32'h10a00000;
      73627: inst = 32'hca00004;
      73628: inst = 32'h38632800;
      73629: inst = 32'h38842800;
      73630: inst = 32'h10a00001;
      73631: inst = 32'hca01fa3;
      73632: inst = 32'h13e00001;
      73633: inst = 32'hfe0d96a;
      73634: inst = 32'h5be00000;
      73635: inst = 32'h8c50000;
      73636: inst = 32'h24612800;
      73637: inst = 32'h10a0ffff;
      73638: inst = 32'hca0fffc;
      73639: inst = 32'h24822800;
      73640: inst = 32'h10a00000;
      73641: inst = 32'hca00004;
      73642: inst = 32'h38632800;
      73643: inst = 32'h38842800;
      73644: inst = 32'h10a00001;
      73645: inst = 32'hca01fb1;
      73646: inst = 32'h13e00001;
      73647: inst = 32'hfe0d96a;
      73648: inst = 32'h5be00000;
      73649: inst = 32'h8c50000;
      73650: inst = 32'h24612800;
      73651: inst = 32'h10a0ffff;
      73652: inst = 32'hca0fffc;
      73653: inst = 32'h24822800;
      73654: inst = 32'h10a00000;
      73655: inst = 32'hca00004;
      73656: inst = 32'h38632800;
      73657: inst = 32'h38842800;
      73658: inst = 32'h10a00001;
      73659: inst = 32'hca01fbf;
      73660: inst = 32'h13e00001;
      73661: inst = 32'hfe0d96a;
      73662: inst = 32'h5be00000;
      73663: inst = 32'h8c50000;
      73664: inst = 32'h24612800;
      73665: inst = 32'h10a0ffff;
      73666: inst = 32'hca0fffc;
      73667: inst = 32'h24822800;
      73668: inst = 32'h10a00000;
      73669: inst = 32'hca00004;
      73670: inst = 32'h38632800;
      73671: inst = 32'h38842800;
      73672: inst = 32'h10a00001;
      73673: inst = 32'hca01fcd;
      73674: inst = 32'h13e00001;
      73675: inst = 32'hfe0d96a;
      73676: inst = 32'h5be00000;
      73677: inst = 32'h8c50000;
      73678: inst = 32'h24612800;
      73679: inst = 32'h10a0ffff;
      73680: inst = 32'hca0fffc;
      73681: inst = 32'h24822800;
      73682: inst = 32'h10a00000;
      73683: inst = 32'hca00004;
      73684: inst = 32'h38632800;
      73685: inst = 32'h38842800;
      73686: inst = 32'h10a00001;
      73687: inst = 32'hca01fdb;
      73688: inst = 32'h13e00001;
      73689: inst = 32'hfe0d96a;
      73690: inst = 32'h5be00000;
      73691: inst = 32'h8c50000;
      73692: inst = 32'h24612800;
      73693: inst = 32'h10a0ffff;
      73694: inst = 32'hca0fffc;
      73695: inst = 32'h24822800;
      73696: inst = 32'h10a00000;
      73697: inst = 32'hca00004;
      73698: inst = 32'h38632800;
      73699: inst = 32'h38842800;
      73700: inst = 32'h10a00001;
      73701: inst = 32'hca01fe9;
      73702: inst = 32'h13e00001;
      73703: inst = 32'hfe0d96a;
      73704: inst = 32'h5be00000;
      73705: inst = 32'h8c50000;
      73706: inst = 32'h24612800;
      73707: inst = 32'h10a0ffff;
      73708: inst = 32'hca0fffc;
      73709: inst = 32'h24822800;
      73710: inst = 32'h10a00000;
      73711: inst = 32'hca00004;
      73712: inst = 32'h38632800;
      73713: inst = 32'h38842800;
      73714: inst = 32'h10a00001;
      73715: inst = 32'hca01ff7;
      73716: inst = 32'h13e00001;
      73717: inst = 32'hfe0d96a;
      73718: inst = 32'h5be00000;
      73719: inst = 32'h8c50000;
      73720: inst = 32'h24612800;
      73721: inst = 32'h10a0ffff;
      73722: inst = 32'hca0fffc;
      73723: inst = 32'h24822800;
      73724: inst = 32'h10a00000;
      73725: inst = 32'hca00004;
      73726: inst = 32'h38632800;
      73727: inst = 32'h38842800;
      73728: inst = 32'h10a00001;
      73729: inst = 32'hca02005;
      73730: inst = 32'h13e00001;
      73731: inst = 32'hfe0d96a;
      73732: inst = 32'h5be00000;
      73733: inst = 32'h8c50000;
      73734: inst = 32'h24612800;
      73735: inst = 32'h10a0ffff;
      73736: inst = 32'hca0fffc;
      73737: inst = 32'h24822800;
      73738: inst = 32'h10a00000;
      73739: inst = 32'hca00004;
      73740: inst = 32'h38632800;
      73741: inst = 32'h38842800;
      73742: inst = 32'h10a00001;
      73743: inst = 32'hca02013;
      73744: inst = 32'h13e00001;
      73745: inst = 32'hfe0d96a;
      73746: inst = 32'h5be00000;
      73747: inst = 32'h8c50000;
      73748: inst = 32'h24612800;
      73749: inst = 32'h10a0ffff;
      73750: inst = 32'hca0fffc;
      73751: inst = 32'h24822800;
      73752: inst = 32'h10a00000;
      73753: inst = 32'hca00004;
      73754: inst = 32'h38632800;
      73755: inst = 32'h38842800;
      73756: inst = 32'h10a00001;
      73757: inst = 32'hca02021;
      73758: inst = 32'h13e00001;
      73759: inst = 32'hfe0d96a;
      73760: inst = 32'h5be00000;
      73761: inst = 32'h8c50000;
      73762: inst = 32'h24612800;
      73763: inst = 32'h10a0ffff;
      73764: inst = 32'hca0fffc;
      73765: inst = 32'h24822800;
      73766: inst = 32'h10a00000;
      73767: inst = 32'hca00004;
      73768: inst = 32'h38632800;
      73769: inst = 32'h38842800;
      73770: inst = 32'h10a00001;
      73771: inst = 32'hca0202f;
      73772: inst = 32'h13e00001;
      73773: inst = 32'hfe0d96a;
      73774: inst = 32'h5be00000;
      73775: inst = 32'h8c50000;
      73776: inst = 32'h24612800;
      73777: inst = 32'h10a0ffff;
      73778: inst = 32'hca0fffc;
      73779: inst = 32'h24822800;
      73780: inst = 32'h10a00000;
      73781: inst = 32'hca00004;
      73782: inst = 32'h38632800;
      73783: inst = 32'h38842800;
      73784: inst = 32'h10a00001;
      73785: inst = 32'hca0203d;
      73786: inst = 32'h13e00001;
      73787: inst = 32'hfe0d96a;
      73788: inst = 32'h5be00000;
      73789: inst = 32'h8c50000;
      73790: inst = 32'h24612800;
      73791: inst = 32'h10a0ffff;
      73792: inst = 32'hca0fffc;
      73793: inst = 32'h24822800;
      73794: inst = 32'h10a00000;
      73795: inst = 32'hca00004;
      73796: inst = 32'h38632800;
      73797: inst = 32'h38842800;
      73798: inst = 32'h10a00001;
      73799: inst = 32'hca0204b;
      73800: inst = 32'h13e00001;
      73801: inst = 32'hfe0d96a;
      73802: inst = 32'h5be00000;
      73803: inst = 32'h8c50000;
      73804: inst = 32'h24612800;
      73805: inst = 32'h10a0ffff;
      73806: inst = 32'hca0fffc;
      73807: inst = 32'h24822800;
      73808: inst = 32'h10a00000;
      73809: inst = 32'hca00004;
      73810: inst = 32'h38632800;
      73811: inst = 32'h38842800;
      73812: inst = 32'h10a00001;
      73813: inst = 32'hca02059;
      73814: inst = 32'h13e00001;
      73815: inst = 32'hfe0d96a;
      73816: inst = 32'h5be00000;
      73817: inst = 32'h8c50000;
      73818: inst = 32'h24612800;
      73819: inst = 32'h10a0ffff;
      73820: inst = 32'hca0fffc;
      73821: inst = 32'h24822800;
      73822: inst = 32'h10a00000;
      73823: inst = 32'hca00004;
      73824: inst = 32'h38632800;
      73825: inst = 32'h38842800;
      73826: inst = 32'h10a00001;
      73827: inst = 32'hca02067;
      73828: inst = 32'h13e00001;
      73829: inst = 32'hfe0d96a;
      73830: inst = 32'h5be00000;
      73831: inst = 32'h8c50000;
      73832: inst = 32'h24612800;
      73833: inst = 32'h10a0ffff;
      73834: inst = 32'hca0fffc;
      73835: inst = 32'h24822800;
      73836: inst = 32'h10a00000;
      73837: inst = 32'hca00004;
      73838: inst = 32'h38632800;
      73839: inst = 32'h38842800;
      73840: inst = 32'h10a00001;
      73841: inst = 32'hca02075;
      73842: inst = 32'h13e00001;
      73843: inst = 32'hfe0d96a;
      73844: inst = 32'h5be00000;
      73845: inst = 32'h8c50000;
      73846: inst = 32'h24612800;
      73847: inst = 32'h10a0ffff;
      73848: inst = 32'hca0fffc;
      73849: inst = 32'h24822800;
      73850: inst = 32'h10a00000;
      73851: inst = 32'hca00004;
      73852: inst = 32'h38632800;
      73853: inst = 32'h38842800;
      73854: inst = 32'h10a00001;
      73855: inst = 32'hca02083;
      73856: inst = 32'h13e00001;
      73857: inst = 32'hfe0d96a;
      73858: inst = 32'h5be00000;
      73859: inst = 32'h8c50000;
      73860: inst = 32'h24612800;
      73861: inst = 32'h10a0ffff;
      73862: inst = 32'hca0fffc;
      73863: inst = 32'h24822800;
      73864: inst = 32'h10a00000;
      73865: inst = 32'hca00004;
      73866: inst = 32'h38632800;
      73867: inst = 32'h38842800;
      73868: inst = 32'h10a00001;
      73869: inst = 32'hca02091;
      73870: inst = 32'h13e00001;
      73871: inst = 32'hfe0d96a;
      73872: inst = 32'h5be00000;
      73873: inst = 32'h8c50000;
      73874: inst = 32'h24612800;
      73875: inst = 32'h10a0ffff;
      73876: inst = 32'hca0fffc;
      73877: inst = 32'h24822800;
      73878: inst = 32'h10a00000;
      73879: inst = 32'hca00004;
      73880: inst = 32'h38632800;
      73881: inst = 32'h38842800;
      73882: inst = 32'h10a00001;
      73883: inst = 32'hca0209f;
      73884: inst = 32'h13e00001;
      73885: inst = 32'hfe0d96a;
      73886: inst = 32'h5be00000;
      73887: inst = 32'h8c50000;
      73888: inst = 32'h24612800;
      73889: inst = 32'h10a0ffff;
      73890: inst = 32'hca0fffc;
      73891: inst = 32'h24822800;
      73892: inst = 32'h10a00000;
      73893: inst = 32'hca00004;
      73894: inst = 32'h38632800;
      73895: inst = 32'h38842800;
      73896: inst = 32'h10a00001;
      73897: inst = 32'hca020ad;
      73898: inst = 32'h13e00001;
      73899: inst = 32'hfe0d96a;
      73900: inst = 32'h5be00000;
      73901: inst = 32'h8c50000;
      73902: inst = 32'h24612800;
      73903: inst = 32'h10a0ffff;
      73904: inst = 32'hca0fffc;
      73905: inst = 32'h24822800;
      73906: inst = 32'h10a00000;
      73907: inst = 32'hca00004;
      73908: inst = 32'h38632800;
      73909: inst = 32'h38842800;
      73910: inst = 32'h10a00001;
      73911: inst = 32'hca020bb;
      73912: inst = 32'h13e00001;
      73913: inst = 32'hfe0d96a;
      73914: inst = 32'h5be00000;
      73915: inst = 32'h8c50000;
      73916: inst = 32'h24612800;
      73917: inst = 32'h10a0ffff;
      73918: inst = 32'hca0fffc;
      73919: inst = 32'h24822800;
      73920: inst = 32'h10a00000;
      73921: inst = 32'hca00004;
      73922: inst = 32'h38632800;
      73923: inst = 32'h38842800;
      73924: inst = 32'h10a00001;
      73925: inst = 32'hca020c9;
      73926: inst = 32'h13e00001;
      73927: inst = 32'hfe0d96a;
      73928: inst = 32'h5be00000;
      73929: inst = 32'h8c50000;
      73930: inst = 32'h24612800;
      73931: inst = 32'h10a0ffff;
      73932: inst = 32'hca0fffc;
      73933: inst = 32'h24822800;
      73934: inst = 32'h10a00000;
      73935: inst = 32'hca00004;
      73936: inst = 32'h38632800;
      73937: inst = 32'h38842800;
      73938: inst = 32'h10a00001;
      73939: inst = 32'hca020d7;
      73940: inst = 32'h13e00001;
      73941: inst = 32'hfe0d96a;
      73942: inst = 32'h5be00000;
      73943: inst = 32'h8c50000;
      73944: inst = 32'h24612800;
      73945: inst = 32'h10a0ffff;
      73946: inst = 32'hca0fffc;
      73947: inst = 32'h24822800;
      73948: inst = 32'h10a00000;
      73949: inst = 32'hca00004;
      73950: inst = 32'h38632800;
      73951: inst = 32'h38842800;
      73952: inst = 32'h10a00001;
      73953: inst = 32'hca020e5;
      73954: inst = 32'h13e00001;
      73955: inst = 32'hfe0d96a;
      73956: inst = 32'h5be00000;
      73957: inst = 32'h8c50000;
      73958: inst = 32'h24612800;
      73959: inst = 32'h10a0ffff;
      73960: inst = 32'hca0fffc;
      73961: inst = 32'h24822800;
      73962: inst = 32'h10a00000;
      73963: inst = 32'hca00004;
      73964: inst = 32'h38632800;
      73965: inst = 32'h38842800;
      73966: inst = 32'h10a00001;
      73967: inst = 32'hca020f3;
      73968: inst = 32'h13e00001;
      73969: inst = 32'hfe0d96a;
      73970: inst = 32'h5be00000;
      73971: inst = 32'h8c50000;
      73972: inst = 32'h24612800;
      73973: inst = 32'h10a0ffff;
      73974: inst = 32'hca0fffc;
      73975: inst = 32'h24822800;
      73976: inst = 32'h10a00000;
      73977: inst = 32'hca00004;
      73978: inst = 32'h38632800;
      73979: inst = 32'h38842800;
      73980: inst = 32'h10a00001;
      73981: inst = 32'hca02101;
      73982: inst = 32'h13e00001;
      73983: inst = 32'hfe0d96a;
      73984: inst = 32'h5be00000;
      73985: inst = 32'h8c50000;
      73986: inst = 32'h24612800;
      73987: inst = 32'h10a0ffff;
      73988: inst = 32'hca0fffc;
      73989: inst = 32'h24822800;
      73990: inst = 32'h10a00000;
      73991: inst = 32'hca00004;
      73992: inst = 32'h38632800;
      73993: inst = 32'h38842800;
      73994: inst = 32'h10a00001;
      73995: inst = 32'hca0210f;
      73996: inst = 32'h13e00001;
      73997: inst = 32'hfe0d96a;
      73998: inst = 32'h5be00000;
      73999: inst = 32'h8c50000;
      74000: inst = 32'h24612800;
      74001: inst = 32'h10a0ffff;
      74002: inst = 32'hca0fffc;
      74003: inst = 32'h24822800;
      74004: inst = 32'h10a00000;
      74005: inst = 32'hca00004;
      74006: inst = 32'h38632800;
      74007: inst = 32'h38842800;
      74008: inst = 32'h10a00001;
      74009: inst = 32'hca0211d;
      74010: inst = 32'h13e00001;
      74011: inst = 32'hfe0d96a;
      74012: inst = 32'h5be00000;
      74013: inst = 32'h8c50000;
      74014: inst = 32'h24612800;
      74015: inst = 32'h10a0ffff;
      74016: inst = 32'hca0fffc;
      74017: inst = 32'h24822800;
      74018: inst = 32'h10a00000;
      74019: inst = 32'hca00004;
      74020: inst = 32'h38632800;
      74021: inst = 32'h38842800;
      74022: inst = 32'h10a00001;
      74023: inst = 32'hca0212b;
      74024: inst = 32'h13e00001;
      74025: inst = 32'hfe0d96a;
      74026: inst = 32'h5be00000;
      74027: inst = 32'h8c50000;
      74028: inst = 32'h24612800;
      74029: inst = 32'h10a0ffff;
      74030: inst = 32'hca0fffc;
      74031: inst = 32'h24822800;
      74032: inst = 32'h10a00000;
      74033: inst = 32'hca00004;
      74034: inst = 32'h38632800;
      74035: inst = 32'h38842800;
      74036: inst = 32'h10a00001;
      74037: inst = 32'hca02139;
      74038: inst = 32'h13e00001;
      74039: inst = 32'hfe0d96a;
      74040: inst = 32'h5be00000;
      74041: inst = 32'h8c50000;
      74042: inst = 32'h24612800;
      74043: inst = 32'h10a0ffff;
      74044: inst = 32'hca0fffc;
      74045: inst = 32'h24822800;
      74046: inst = 32'h10a00000;
      74047: inst = 32'hca00004;
      74048: inst = 32'h38632800;
      74049: inst = 32'h38842800;
      74050: inst = 32'h10a00001;
      74051: inst = 32'hca02147;
      74052: inst = 32'h13e00001;
      74053: inst = 32'hfe0d96a;
      74054: inst = 32'h5be00000;
      74055: inst = 32'h8c50000;
      74056: inst = 32'h24612800;
      74057: inst = 32'h10a0ffff;
      74058: inst = 32'hca0fffc;
      74059: inst = 32'h24822800;
      74060: inst = 32'h10a00000;
      74061: inst = 32'hca00004;
      74062: inst = 32'h38632800;
      74063: inst = 32'h38842800;
      74064: inst = 32'h10a00001;
      74065: inst = 32'hca02155;
      74066: inst = 32'h13e00001;
      74067: inst = 32'hfe0d96a;
      74068: inst = 32'h5be00000;
      74069: inst = 32'h8c50000;
      74070: inst = 32'h24612800;
      74071: inst = 32'h10a0ffff;
      74072: inst = 32'hca0fffc;
      74073: inst = 32'h24822800;
      74074: inst = 32'h10a00000;
      74075: inst = 32'hca00004;
      74076: inst = 32'h38632800;
      74077: inst = 32'h38842800;
      74078: inst = 32'h10a00001;
      74079: inst = 32'hca02163;
      74080: inst = 32'h13e00001;
      74081: inst = 32'hfe0d96a;
      74082: inst = 32'h5be00000;
      74083: inst = 32'h8c50000;
      74084: inst = 32'h24612800;
      74085: inst = 32'h10a0ffff;
      74086: inst = 32'hca0fffc;
      74087: inst = 32'h24822800;
      74088: inst = 32'h10a00000;
      74089: inst = 32'hca00004;
      74090: inst = 32'h38632800;
      74091: inst = 32'h38842800;
      74092: inst = 32'h10a00001;
      74093: inst = 32'hca02171;
      74094: inst = 32'h13e00001;
      74095: inst = 32'hfe0d96a;
      74096: inst = 32'h5be00000;
      74097: inst = 32'h8c50000;
      74098: inst = 32'h24612800;
      74099: inst = 32'h10a0ffff;
      74100: inst = 32'hca0fffc;
      74101: inst = 32'h24822800;
      74102: inst = 32'h10a00000;
      74103: inst = 32'hca00004;
      74104: inst = 32'h38632800;
      74105: inst = 32'h38842800;
      74106: inst = 32'h10a00001;
      74107: inst = 32'hca0217f;
      74108: inst = 32'h13e00001;
      74109: inst = 32'hfe0d96a;
      74110: inst = 32'h5be00000;
      74111: inst = 32'h8c50000;
      74112: inst = 32'h24612800;
      74113: inst = 32'h10a0ffff;
      74114: inst = 32'hca0fffc;
      74115: inst = 32'h24822800;
      74116: inst = 32'h10a00000;
      74117: inst = 32'hca00004;
      74118: inst = 32'h38632800;
      74119: inst = 32'h38842800;
      74120: inst = 32'h10a00001;
      74121: inst = 32'hca0218d;
      74122: inst = 32'h13e00001;
      74123: inst = 32'hfe0d96a;
      74124: inst = 32'h5be00000;
      74125: inst = 32'h8c50000;
      74126: inst = 32'h24612800;
      74127: inst = 32'h10a0ffff;
      74128: inst = 32'hca0fffc;
      74129: inst = 32'h24822800;
      74130: inst = 32'h10a00000;
      74131: inst = 32'hca00004;
      74132: inst = 32'h38632800;
      74133: inst = 32'h38842800;
      74134: inst = 32'h10a00001;
      74135: inst = 32'hca0219b;
      74136: inst = 32'h13e00001;
      74137: inst = 32'hfe0d96a;
      74138: inst = 32'h5be00000;
      74139: inst = 32'h8c50000;
      74140: inst = 32'h24612800;
      74141: inst = 32'h10a0ffff;
      74142: inst = 32'hca0fffc;
      74143: inst = 32'h24822800;
      74144: inst = 32'h10a00000;
      74145: inst = 32'hca00004;
      74146: inst = 32'h38632800;
      74147: inst = 32'h38842800;
      74148: inst = 32'h10a00001;
      74149: inst = 32'hca021a9;
      74150: inst = 32'h13e00001;
      74151: inst = 32'hfe0d96a;
      74152: inst = 32'h5be00000;
      74153: inst = 32'h8c50000;
      74154: inst = 32'h24612800;
      74155: inst = 32'h10a0ffff;
      74156: inst = 32'hca0fffd;
      74157: inst = 32'h24822800;
      74158: inst = 32'h10a00000;
      74159: inst = 32'hca00004;
      74160: inst = 32'h38632800;
      74161: inst = 32'h38842800;
      74162: inst = 32'h10a00001;
      74163: inst = 32'hca021b7;
      74164: inst = 32'h13e00001;
      74165: inst = 32'hfe0d96a;
      74166: inst = 32'h5be00000;
      74167: inst = 32'h8c50000;
      74168: inst = 32'h24612800;
      74169: inst = 32'h10a0ffff;
      74170: inst = 32'hca0fffd;
      74171: inst = 32'h24822800;
      74172: inst = 32'h10a00000;
      74173: inst = 32'hca00004;
      74174: inst = 32'h38632800;
      74175: inst = 32'h38842800;
      74176: inst = 32'h10a00001;
      74177: inst = 32'hca021c5;
      74178: inst = 32'h13e00001;
      74179: inst = 32'hfe0d96a;
      74180: inst = 32'h5be00000;
      74181: inst = 32'h8c50000;
      74182: inst = 32'h24612800;
      74183: inst = 32'h10a0ffff;
      74184: inst = 32'hca0fffd;
      74185: inst = 32'h24822800;
      74186: inst = 32'h10a00000;
      74187: inst = 32'hca00004;
      74188: inst = 32'h38632800;
      74189: inst = 32'h38842800;
      74190: inst = 32'h10a00001;
      74191: inst = 32'hca021d3;
      74192: inst = 32'h13e00001;
      74193: inst = 32'hfe0d96a;
      74194: inst = 32'h5be00000;
      74195: inst = 32'h8c50000;
      74196: inst = 32'h24612800;
      74197: inst = 32'h10a0ffff;
      74198: inst = 32'hca0fffd;
      74199: inst = 32'h24822800;
      74200: inst = 32'h10a00000;
      74201: inst = 32'hca00004;
      74202: inst = 32'h38632800;
      74203: inst = 32'h38842800;
      74204: inst = 32'h10a00001;
      74205: inst = 32'hca021e1;
      74206: inst = 32'h13e00001;
      74207: inst = 32'hfe0d96a;
      74208: inst = 32'h5be00000;
      74209: inst = 32'h8c50000;
      74210: inst = 32'h24612800;
      74211: inst = 32'h10a0ffff;
      74212: inst = 32'hca0fffd;
      74213: inst = 32'h24822800;
      74214: inst = 32'h10a00000;
      74215: inst = 32'hca00004;
      74216: inst = 32'h38632800;
      74217: inst = 32'h38842800;
      74218: inst = 32'h10a00001;
      74219: inst = 32'hca021ef;
      74220: inst = 32'h13e00001;
      74221: inst = 32'hfe0d96a;
      74222: inst = 32'h5be00000;
      74223: inst = 32'h8c50000;
      74224: inst = 32'h24612800;
      74225: inst = 32'h10a0ffff;
      74226: inst = 32'hca0fffd;
      74227: inst = 32'h24822800;
      74228: inst = 32'h10a00000;
      74229: inst = 32'hca00004;
      74230: inst = 32'h38632800;
      74231: inst = 32'h38842800;
      74232: inst = 32'h10a00001;
      74233: inst = 32'hca021fd;
      74234: inst = 32'h13e00001;
      74235: inst = 32'hfe0d96a;
      74236: inst = 32'h5be00000;
      74237: inst = 32'h8c50000;
      74238: inst = 32'h24612800;
      74239: inst = 32'h10a0ffff;
      74240: inst = 32'hca0fffd;
      74241: inst = 32'h24822800;
      74242: inst = 32'h10a00000;
      74243: inst = 32'hca00004;
      74244: inst = 32'h38632800;
      74245: inst = 32'h38842800;
      74246: inst = 32'h10a00001;
      74247: inst = 32'hca0220b;
      74248: inst = 32'h13e00001;
      74249: inst = 32'hfe0d96a;
      74250: inst = 32'h5be00000;
      74251: inst = 32'h8c50000;
      74252: inst = 32'h24612800;
      74253: inst = 32'h10a0ffff;
      74254: inst = 32'hca0fffd;
      74255: inst = 32'h24822800;
      74256: inst = 32'h10a00000;
      74257: inst = 32'hca00004;
      74258: inst = 32'h38632800;
      74259: inst = 32'h38842800;
      74260: inst = 32'h10a00001;
      74261: inst = 32'hca02219;
      74262: inst = 32'h13e00001;
      74263: inst = 32'hfe0d96a;
      74264: inst = 32'h5be00000;
      74265: inst = 32'h8c50000;
      74266: inst = 32'h24612800;
      74267: inst = 32'h10a0ffff;
      74268: inst = 32'hca0fffd;
      74269: inst = 32'h24822800;
      74270: inst = 32'h10a00000;
      74271: inst = 32'hca00004;
      74272: inst = 32'h38632800;
      74273: inst = 32'h38842800;
      74274: inst = 32'h10a00001;
      74275: inst = 32'hca02227;
      74276: inst = 32'h13e00001;
      74277: inst = 32'hfe0d96a;
      74278: inst = 32'h5be00000;
      74279: inst = 32'h8c50000;
      74280: inst = 32'h24612800;
      74281: inst = 32'h10a0ffff;
      74282: inst = 32'hca0fffd;
      74283: inst = 32'h24822800;
      74284: inst = 32'h10a00000;
      74285: inst = 32'hca00004;
      74286: inst = 32'h38632800;
      74287: inst = 32'h38842800;
      74288: inst = 32'h10a00001;
      74289: inst = 32'hca02235;
      74290: inst = 32'h13e00001;
      74291: inst = 32'hfe0d96a;
      74292: inst = 32'h5be00000;
      74293: inst = 32'h8c50000;
      74294: inst = 32'h24612800;
      74295: inst = 32'h10a0ffff;
      74296: inst = 32'hca0fffd;
      74297: inst = 32'h24822800;
      74298: inst = 32'h10a00000;
      74299: inst = 32'hca00004;
      74300: inst = 32'h38632800;
      74301: inst = 32'h38842800;
      74302: inst = 32'h10a00001;
      74303: inst = 32'hca02243;
      74304: inst = 32'h13e00001;
      74305: inst = 32'hfe0d96a;
      74306: inst = 32'h5be00000;
      74307: inst = 32'h8c50000;
      74308: inst = 32'h24612800;
      74309: inst = 32'h10a0ffff;
      74310: inst = 32'hca0fffd;
      74311: inst = 32'h24822800;
      74312: inst = 32'h10a00000;
      74313: inst = 32'hca00004;
      74314: inst = 32'h38632800;
      74315: inst = 32'h38842800;
      74316: inst = 32'h10a00001;
      74317: inst = 32'hca02251;
      74318: inst = 32'h13e00001;
      74319: inst = 32'hfe0d96a;
      74320: inst = 32'h5be00000;
      74321: inst = 32'h8c50000;
      74322: inst = 32'h24612800;
      74323: inst = 32'h10a0ffff;
      74324: inst = 32'hca0fffd;
      74325: inst = 32'h24822800;
      74326: inst = 32'h10a00000;
      74327: inst = 32'hca00004;
      74328: inst = 32'h38632800;
      74329: inst = 32'h38842800;
      74330: inst = 32'h10a00001;
      74331: inst = 32'hca0225f;
      74332: inst = 32'h13e00001;
      74333: inst = 32'hfe0d96a;
      74334: inst = 32'h5be00000;
      74335: inst = 32'h8c50000;
      74336: inst = 32'h24612800;
      74337: inst = 32'h10a0ffff;
      74338: inst = 32'hca0fffd;
      74339: inst = 32'h24822800;
      74340: inst = 32'h10a00000;
      74341: inst = 32'hca00004;
      74342: inst = 32'h38632800;
      74343: inst = 32'h38842800;
      74344: inst = 32'h10a00001;
      74345: inst = 32'hca0226d;
      74346: inst = 32'h13e00001;
      74347: inst = 32'hfe0d96a;
      74348: inst = 32'h5be00000;
      74349: inst = 32'h8c50000;
      74350: inst = 32'h24612800;
      74351: inst = 32'h10a0ffff;
      74352: inst = 32'hca0fffd;
      74353: inst = 32'h24822800;
      74354: inst = 32'h10a00000;
      74355: inst = 32'hca00004;
      74356: inst = 32'h38632800;
      74357: inst = 32'h38842800;
      74358: inst = 32'h10a00001;
      74359: inst = 32'hca0227b;
      74360: inst = 32'h13e00001;
      74361: inst = 32'hfe0d96a;
      74362: inst = 32'h5be00000;
      74363: inst = 32'h8c50000;
      74364: inst = 32'h24612800;
      74365: inst = 32'h10a0ffff;
      74366: inst = 32'hca0fffd;
      74367: inst = 32'h24822800;
      74368: inst = 32'h10a00000;
      74369: inst = 32'hca00004;
      74370: inst = 32'h38632800;
      74371: inst = 32'h38842800;
      74372: inst = 32'h10a00001;
      74373: inst = 32'hca02289;
      74374: inst = 32'h13e00001;
      74375: inst = 32'hfe0d96a;
      74376: inst = 32'h5be00000;
      74377: inst = 32'h8c50000;
      74378: inst = 32'h24612800;
      74379: inst = 32'h10a0ffff;
      74380: inst = 32'hca0fffd;
      74381: inst = 32'h24822800;
      74382: inst = 32'h10a00000;
      74383: inst = 32'hca00004;
      74384: inst = 32'h38632800;
      74385: inst = 32'h38842800;
      74386: inst = 32'h10a00001;
      74387: inst = 32'hca02297;
      74388: inst = 32'h13e00001;
      74389: inst = 32'hfe0d96a;
      74390: inst = 32'h5be00000;
      74391: inst = 32'h8c50000;
      74392: inst = 32'h24612800;
      74393: inst = 32'h10a0ffff;
      74394: inst = 32'hca0fffd;
      74395: inst = 32'h24822800;
      74396: inst = 32'h10a00000;
      74397: inst = 32'hca00004;
      74398: inst = 32'h38632800;
      74399: inst = 32'h38842800;
      74400: inst = 32'h10a00001;
      74401: inst = 32'hca022a5;
      74402: inst = 32'h13e00001;
      74403: inst = 32'hfe0d96a;
      74404: inst = 32'h5be00000;
      74405: inst = 32'h8c50000;
      74406: inst = 32'h24612800;
      74407: inst = 32'h10a0ffff;
      74408: inst = 32'hca0fffd;
      74409: inst = 32'h24822800;
      74410: inst = 32'h10a00000;
      74411: inst = 32'hca00004;
      74412: inst = 32'h38632800;
      74413: inst = 32'h38842800;
      74414: inst = 32'h10a00001;
      74415: inst = 32'hca022b3;
      74416: inst = 32'h13e00001;
      74417: inst = 32'hfe0d96a;
      74418: inst = 32'h5be00000;
      74419: inst = 32'h8c50000;
      74420: inst = 32'h24612800;
      74421: inst = 32'h10a0ffff;
      74422: inst = 32'hca0fffd;
      74423: inst = 32'h24822800;
      74424: inst = 32'h10a00000;
      74425: inst = 32'hca00004;
      74426: inst = 32'h38632800;
      74427: inst = 32'h38842800;
      74428: inst = 32'h10a00001;
      74429: inst = 32'hca022c1;
      74430: inst = 32'h13e00001;
      74431: inst = 32'hfe0d96a;
      74432: inst = 32'h5be00000;
      74433: inst = 32'h8c50000;
      74434: inst = 32'h24612800;
      74435: inst = 32'h10a0ffff;
      74436: inst = 32'hca0fffd;
      74437: inst = 32'h24822800;
      74438: inst = 32'h10a00000;
      74439: inst = 32'hca00004;
      74440: inst = 32'h38632800;
      74441: inst = 32'h38842800;
      74442: inst = 32'h10a00001;
      74443: inst = 32'hca022cf;
      74444: inst = 32'h13e00001;
      74445: inst = 32'hfe0d96a;
      74446: inst = 32'h5be00000;
      74447: inst = 32'h8c50000;
      74448: inst = 32'h24612800;
      74449: inst = 32'h10a0ffff;
      74450: inst = 32'hca0fffd;
      74451: inst = 32'h24822800;
      74452: inst = 32'h10a00000;
      74453: inst = 32'hca00004;
      74454: inst = 32'h38632800;
      74455: inst = 32'h38842800;
      74456: inst = 32'h10a00001;
      74457: inst = 32'hca022dd;
      74458: inst = 32'h13e00001;
      74459: inst = 32'hfe0d96a;
      74460: inst = 32'h5be00000;
      74461: inst = 32'h8c50000;
      74462: inst = 32'h24612800;
      74463: inst = 32'h10a0ffff;
      74464: inst = 32'hca0fffd;
      74465: inst = 32'h24822800;
      74466: inst = 32'h10a00000;
      74467: inst = 32'hca00004;
      74468: inst = 32'h38632800;
      74469: inst = 32'h38842800;
      74470: inst = 32'h10a00001;
      74471: inst = 32'hca022eb;
      74472: inst = 32'h13e00001;
      74473: inst = 32'hfe0d96a;
      74474: inst = 32'h5be00000;
      74475: inst = 32'h8c50000;
      74476: inst = 32'h24612800;
      74477: inst = 32'h10a0ffff;
      74478: inst = 32'hca0fffd;
      74479: inst = 32'h24822800;
      74480: inst = 32'h10a00000;
      74481: inst = 32'hca00004;
      74482: inst = 32'h38632800;
      74483: inst = 32'h38842800;
      74484: inst = 32'h10a00001;
      74485: inst = 32'hca022f9;
      74486: inst = 32'h13e00001;
      74487: inst = 32'hfe0d96a;
      74488: inst = 32'h5be00000;
      74489: inst = 32'h8c50000;
      74490: inst = 32'h24612800;
      74491: inst = 32'h10a0ffff;
      74492: inst = 32'hca0fffd;
      74493: inst = 32'h24822800;
      74494: inst = 32'h10a00000;
      74495: inst = 32'hca00004;
      74496: inst = 32'h38632800;
      74497: inst = 32'h38842800;
      74498: inst = 32'h10a00001;
      74499: inst = 32'hca02307;
      74500: inst = 32'h13e00001;
      74501: inst = 32'hfe0d96a;
      74502: inst = 32'h5be00000;
      74503: inst = 32'h8c50000;
      74504: inst = 32'h24612800;
      74505: inst = 32'h10a0ffff;
      74506: inst = 32'hca0fffd;
      74507: inst = 32'h24822800;
      74508: inst = 32'h10a00000;
      74509: inst = 32'hca00004;
      74510: inst = 32'h38632800;
      74511: inst = 32'h38842800;
      74512: inst = 32'h10a00001;
      74513: inst = 32'hca02315;
      74514: inst = 32'h13e00001;
      74515: inst = 32'hfe0d96a;
      74516: inst = 32'h5be00000;
      74517: inst = 32'h8c50000;
      74518: inst = 32'h24612800;
      74519: inst = 32'h10a0ffff;
      74520: inst = 32'hca0fffd;
      74521: inst = 32'h24822800;
      74522: inst = 32'h10a00000;
      74523: inst = 32'hca00004;
      74524: inst = 32'h38632800;
      74525: inst = 32'h38842800;
      74526: inst = 32'h10a00001;
      74527: inst = 32'hca02323;
      74528: inst = 32'h13e00001;
      74529: inst = 32'hfe0d96a;
      74530: inst = 32'h5be00000;
      74531: inst = 32'h8c50000;
      74532: inst = 32'h24612800;
      74533: inst = 32'h10a0ffff;
      74534: inst = 32'hca0fffd;
      74535: inst = 32'h24822800;
      74536: inst = 32'h10a00000;
      74537: inst = 32'hca00004;
      74538: inst = 32'h38632800;
      74539: inst = 32'h38842800;
      74540: inst = 32'h10a00001;
      74541: inst = 32'hca02331;
      74542: inst = 32'h13e00001;
      74543: inst = 32'hfe0d96a;
      74544: inst = 32'h5be00000;
      74545: inst = 32'h8c50000;
      74546: inst = 32'h24612800;
      74547: inst = 32'h10a0ffff;
      74548: inst = 32'hca0fffd;
      74549: inst = 32'h24822800;
      74550: inst = 32'h10a00000;
      74551: inst = 32'hca00004;
      74552: inst = 32'h38632800;
      74553: inst = 32'h38842800;
      74554: inst = 32'h10a00001;
      74555: inst = 32'hca0233f;
      74556: inst = 32'h13e00001;
      74557: inst = 32'hfe0d96a;
      74558: inst = 32'h5be00000;
      74559: inst = 32'h8c50000;
      74560: inst = 32'h24612800;
      74561: inst = 32'h10a0ffff;
      74562: inst = 32'hca0fffd;
      74563: inst = 32'h24822800;
      74564: inst = 32'h10a00000;
      74565: inst = 32'hca00004;
      74566: inst = 32'h38632800;
      74567: inst = 32'h38842800;
      74568: inst = 32'h10a00001;
      74569: inst = 32'hca0234d;
      74570: inst = 32'h13e00001;
      74571: inst = 32'hfe0d96a;
      74572: inst = 32'h5be00000;
      74573: inst = 32'h8c50000;
      74574: inst = 32'h24612800;
      74575: inst = 32'h10a0ffff;
      74576: inst = 32'hca0fffd;
      74577: inst = 32'h24822800;
      74578: inst = 32'h10a00000;
      74579: inst = 32'hca00004;
      74580: inst = 32'h38632800;
      74581: inst = 32'h38842800;
      74582: inst = 32'h10a00001;
      74583: inst = 32'hca0235b;
      74584: inst = 32'h13e00001;
      74585: inst = 32'hfe0d96a;
      74586: inst = 32'h5be00000;
      74587: inst = 32'h8c50000;
      74588: inst = 32'h24612800;
      74589: inst = 32'h10a0ffff;
      74590: inst = 32'hca0fffd;
      74591: inst = 32'h24822800;
      74592: inst = 32'h10a00000;
      74593: inst = 32'hca00004;
      74594: inst = 32'h38632800;
      74595: inst = 32'h38842800;
      74596: inst = 32'h10a00001;
      74597: inst = 32'hca02369;
      74598: inst = 32'h13e00001;
      74599: inst = 32'hfe0d96a;
      74600: inst = 32'h5be00000;
      74601: inst = 32'h8c50000;
      74602: inst = 32'h24612800;
      74603: inst = 32'h10a0ffff;
      74604: inst = 32'hca0fffd;
      74605: inst = 32'h24822800;
      74606: inst = 32'h10a00000;
      74607: inst = 32'hca00004;
      74608: inst = 32'h38632800;
      74609: inst = 32'h38842800;
      74610: inst = 32'h10a00001;
      74611: inst = 32'hca02377;
      74612: inst = 32'h13e00001;
      74613: inst = 32'hfe0d96a;
      74614: inst = 32'h5be00000;
      74615: inst = 32'h8c50000;
      74616: inst = 32'h24612800;
      74617: inst = 32'h10a0ffff;
      74618: inst = 32'hca0fffd;
      74619: inst = 32'h24822800;
      74620: inst = 32'h10a00000;
      74621: inst = 32'hca00004;
      74622: inst = 32'h38632800;
      74623: inst = 32'h38842800;
      74624: inst = 32'h10a00001;
      74625: inst = 32'hca02385;
      74626: inst = 32'h13e00001;
      74627: inst = 32'hfe0d96a;
      74628: inst = 32'h5be00000;
      74629: inst = 32'h8c50000;
      74630: inst = 32'h24612800;
      74631: inst = 32'h10a0ffff;
      74632: inst = 32'hca0fffd;
      74633: inst = 32'h24822800;
      74634: inst = 32'h10a00000;
      74635: inst = 32'hca00004;
      74636: inst = 32'h38632800;
      74637: inst = 32'h38842800;
      74638: inst = 32'h10a00001;
      74639: inst = 32'hca02393;
      74640: inst = 32'h13e00001;
      74641: inst = 32'hfe0d96a;
      74642: inst = 32'h5be00000;
      74643: inst = 32'h8c50000;
      74644: inst = 32'h24612800;
      74645: inst = 32'h10a0ffff;
      74646: inst = 32'hca0fffd;
      74647: inst = 32'h24822800;
      74648: inst = 32'h10a00000;
      74649: inst = 32'hca00004;
      74650: inst = 32'h38632800;
      74651: inst = 32'h38842800;
      74652: inst = 32'h10a00001;
      74653: inst = 32'hca023a1;
      74654: inst = 32'h13e00001;
      74655: inst = 32'hfe0d96a;
      74656: inst = 32'h5be00000;
      74657: inst = 32'h8c50000;
      74658: inst = 32'h24612800;
      74659: inst = 32'h10a0ffff;
      74660: inst = 32'hca0fffd;
      74661: inst = 32'h24822800;
      74662: inst = 32'h10a00000;
      74663: inst = 32'hca00004;
      74664: inst = 32'h38632800;
      74665: inst = 32'h38842800;
      74666: inst = 32'h10a00001;
      74667: inst = 32'hca023af;
      74668: inst = 32'h13e00001;
      74669: inst = 32'hfe0d96a;
      74670: inst = 32'h5be00000;
      74671: inst = 32'h8c50000;
      74672: inst = 32'h24612800;
      74673: inst = 32'h10a0ffff;
      74674: inst = 32'hca0fffd;
      74675: inst = 32'h24822800;
      74676: inst = 32'h10a00000;
      74677: inst = 32'hca00004;
      74678: inst = 32'h38632800;
      74679: inst = 32'h38842800;
      74680: inst = 32'h10a00001;
      74681: inst = 32'hca023bd;
      74682: inst = 32'h13e00001;
      74683: inst = 32'hfe0d96a;
      74684: inst = 32'h5be00000;
      74685: inst = 32'h8c50000;
      74686: inst = 32'h24612800;
      74687: inst = 32'h10a0ffff;
      74688: inst = 32'hca0fffd;
      74689: inst = 32'h24822800;
      74690: inst = 32'h10a00000;
      74691: inst = 32'hca00004;
      74692: inst = 32'h38632800;
      74693: inst = 32'h38842800;
      74694: inst = 32'h10a00001;
      74695: inst = 32'hca023cb;
      74696: inst = 32'h13e00001;
      74697: inst = 32'hfe0d96a;
      74698: inst = 32'h5be00000;
      74699: inst = 32'h8c50000;
      74700: inst = 32'h24612800;
      74701: inst = 32'h10a0ffff;
      74702: inst = 32'hca0fffd;
      74703: inst = 32'h24822800;
      74704: inst = 32'h10a00000;
      74705: inst = 32'hca00004;
      74706: inst = 32'h38632800;
      74707: inst = 32'h38842800;
      74708: inst = 32'h10a00001;
      74709: inst = 32'hca023d9;
      74710: inst = 32'h13e00001;
      74711: inst = 32'hfe0d96a;
      74712: inst = 32'h5be00000;
      74713: inst = 32'h8c50000;
      74714: inst = 32'h24612800;
      74715: inst = 32'h10a0ffff;
      74716: inst = 32'hca0fffd;
      74717: inst = 32'h24822800;
      74718: inst = 32'h10a00000;
      74719: inst = 32'hca00004;
      74720: inst = 32'h38632800;
      74721: inst = 32'h38842800;
      74722: inst = 32'h10a00001;
      74723: inst = 32'hca023e7;
      74724: inst = 32'h13e00001;
      74725: inst = 32'hfe0d96a;
      74726: inst = 32'h5be00000;
      74727: inst = 32'h8c50000;
      74728: inst = 32'h24612800;
      74729: inst = 32'h10a0ffff;
      74730: inst = 32'hca0fffd;
      74731: inst = 32'h24822800;
      74732: inst = 32'h10a00000;
      74733: inst = 32'hca00004;
      74734: inst = 32'h38632800;
      74735: inst = 32'h38842800;
      74736: inst = 32'h10a00001;
      74737: inst = 32'hca023f5;
      74738: inst = 32'h13e00001;
      74739: inst = 32'hfe0d96a;
      74740: inst = 32'h5be00000;
      74741: inst = 32'h8c50000;
      74742: inst = 32'h24612800;
      74743: inst = 32'h10a0ffff;
      74744: inst = 32'hca0fffd;
      74745: inst = 32'h24822800;
      74746: inst = 32'h10a00000;
      74747: inst = 32'hca00004;
      74748: inst = 32'h38632800;
      74749: inst = 32'h38842800;
      74750: inst = 32'h10a00001;
      74751: inst = 32'hca02403;
      74752: inst = 32'h13e00001;
      74753: inst = 32'hfe0d96a;
      74754: inst = 32'h5be00000;
      74755: inst = 32'h8c50000;
      74756: inst = 32'h24612800;
      74757: inst = 32'h10a0ffff;
      74758: inst = 32'hca0fffd;
      74759: inst = 32'h24822800;
      74760: inst = 32'h10a00000;
      74761: inst = 32'hca00004;
      74762: inst = 32'h38632800;
      74763: inst = 32'h38842800;
      74764: inst = 32'h10a00001;
      74765: inst = 32'hca02411;
      74766: inst = 32'h13e00001;
      74767: inst = 32'hfe0d96a;
      74768: inst = 32'h5be00000;
      74769: inst = 32'h8c50000;
      74770: inst = 32'h24612800;
      74771: inst = 32'h10a0ffff;
      74772: inst = 32'hca0fffd;
      74773: inst = 32'h24822800;
      74774: inst = 32'h10a00000;
      74775: inst = 32'hca00004;
      74776: inst = 32'h38632800;
      74777: inst = 32'h38842800;
      74778: inst = 32'h10a00001;
      74779: inst = 32'hca0241f;
      74780: inst = 32'h13e00001;
      74781: inst = 32'hfe0d96a;
      74782: inst = 32'h5be00000;
      74783: inst = 32'h8c50000;
      74784: inst = 32'h24612800;
      74785: inst = 32'h10a0ffff;
      74786: inst = 32'hca0fffd;
      74787: inst = 32'h24822800;
      74788: inst = 32'h10a00000;
      74789: inst = 32'hca00004;
      74790: inst = 32'h38632800;
      74791: inst = 32'h38842800;
      74792: inst = 32'h10a00001;
      74793: inst = 32'hca0242d;
      74794: inst = 32'h13e00001;
      74795: inst = 32'hfe0d96a;
      74796: inst = 32'h5be00000;
      74797: inst = 32'h8c50000;
      74798: inst = 32'h24612800;
      74799: inst = 32'h10a0ffff;
      74800: inst = 32'hca0fffd;
      74801: inst = 32'h24822800;
      74802: inst = 32'h10a00000;
      74803: inst = 32'hca00004;
      74804: inst = 32'h38632800;
      74805: inst = 32'h38842800;
      74806: inst = 32'h10a00001;
      74807: inst = 32'hca0243b;
      74808: inst = 32'h13e00001;
      74809: inst = 32'hfe0d96a;
      74810: inst = 32'h5be00000;
      74811: inst = 32'h8c50000;
      74812: inst = 32'h24612800;
      74813: inst = 32'h10a0ffff;
      74814: inst = 32'hca0fffd;
      74815: inst = 32'h24822800;
      74816: inst = 32'h10a00000;
      74817: inst = 32'hca00004;
      74818: inst = 32'h38632800;
      74819: inst = 32'h38842800;
      74820: inst = 32'h10a00001;
      74821: inst = 32'hca02449;
      74822: inst = 32'h13e00001;
      74823: inst = 32'hfe0d96a;
      74824: inst = 32'h5be00000;
      74825: inst = 32'h8c50000;
      74826: inst = 32'h24612800;
      74827: inst = 32'h10a0ffff;
      74828: inst = 32'hca0fffd;
      74829: inst = 32'h24822800;
      74830: inst = 32'h10a00000;
      74831: inst = 32'hca00004;
      74832: inst = 32'h38632800;
      74833: inst = 32'h38842800;
      74834: inst = 32'h10a00001;
      74835: inst = 32'hca02457;
      74836: inst = 32'h13e00001;
      74837: inst = 32'hfe0d96a;
      74838: inst = 32'h5be00000;
      74839: inst = 32'h8c50000;
      74840: inst = 32'h24612800;
      74841: inst = 32'h10a0ffff;
      74842: inst = 32'hca0fffd;
      74843: inst = 32'h24822800;
      74844: inst = 32'h10a00000;
      74845: inst = 32'hca00004;
      74846: inst = 32'h38632800;
      74847: inst = 32'h38842800;
      74848: inst = 32'h10a00001;
      74849: inst = 32'hca02465;
      74850: inst = 32'h13e00001;
      74851: inst = 32'hfe0d96a;
      74852: inst = 32'h5be00000;
      74853: inst = 32'h8c50000;
      74854: inst = 32'h24612800;
      74855: inst = 32'h10a0ffff;
      74856: inst = 32'hca0fffd;
      74857: inst = 32'h24822800;
      74858: inst = 32'h10a00000;
      74859: inst = 32'hca00004;
      74860: inst = 32'h38632800;
      74861: inst = 32'h38842800;
      74862: inst = 32'h10a00001;
      74863: inst = 32'hca02473;
      74864: inst = 32'h13e00001;
      74865: inst = 32'hfe0d96a;
      74866: inst = 32'h5be00000;
      74867: inst = 32'h8c50000;
      74868: inst = 32'h24612800;
      74869: inst = 32'h10a0ffff;
      74870: inst = 32'hca0fffd;
      74871: inst = 32'h24822800;
      74872: inst = 32'h10a00000;
      74873: inst = 32'hca00004;
      74874: inst = 32'h38632800;
      74875: inst = 32'h38842800;
      74876: inst = 32'h10a00001;
      74877: inst = 32'hca02481;
      74878: inst = 32'h13e00001;
      74879: inst = 32'hfe0d96a;
      74880: inst = 32'h5be00000;
      74881: inst = 32'h8c50000;
      74882: inst = 32'h24612800;
      74883: inst = 32'h10a0ffff;
      74884: inst = 32'hca0fffd;
      74885: inst = 32'h24822800;
      74886: inst = 32'h10a00000;
      74887: inst = 32'hca00004;
      74888: inst = 32'h38632800;
      74889: inst = 32'h38842800;
      74890: inst = 32'h10a00001;
      74891: inst = 32'hca0248f;
      74892: inst = 32'h13e00001;
      74893: inst = 32'hfe0d96a;
      74894: inst = 32'h5be00000;
      74895: inst = 32'h8c50000;
      74896: inst = 32'h24612800;
      74897: inst = 32'h10a0ffff;
      74898: inst = 32'hca0fffd;
      74899: inst = 32'h24822800;
      74900: inst = 32'h10a00000;
      74901: inst = 32'hca00004;
      74902: inst = 32'h38632800;
      74903: inst = 32'h38842800;
      74904: inst = 32'h10a00001;
      74905: inst = 32'hca0249d;
      74906: inst = 32'h13e00001;
      74907: inst = 32'hfe0d96a;
      74908: inst = 32'h5be00000;
      74909: inst = 32'h8c50000;
      74910: inst = 32'h24612800;
      74911: inst = 32'h10a0ffff;
      74912: inst = 32'hca0fffd;
      74913: inst = 32'h24822800;
      74914: inst = 32'h10a00000;
      74915: inst = 32'hca00004;
      74916: inst = 32'h38632800;
      74917: inst = 32'h38842800;
      74918: inst = 32'h10a00001;
      74919: inst = 32'hca024ab;
      74920: inst = 32'h13e00001;
      74921: inst = 32'hfe0d96a;
      74922: inst = 32'h5be00000;
      74923: inst = 32'h8c50000;
      74924: inst = 32'h24612800;
      74925: inst = 32'h10a0ffff;
      74926: inst = 32'hca0fffd;
      74927: inst = 32'h24822800;
      74928: inst = 32'h10a00000;
      74929: inst = 32'hca00004;
      74930: inst = 32'h38632800;
      74931: inst = 32'h38842800;
      74932: inst = 32'h10a00001;
      74933: inst = 32'hca024b9;
      74934: inst = 32'h13e00001;
      74935: inst = 32'hfe0d96a;
      74936: inst = 32'h5be00000;
      74937: inst = 32'h8c50000;
      74938: inst = 32'h24612800;
      74939: inst = 32'h10a0ffff;
      74940: inst = 32'hca0fffd;
      74941: inst = 32'h24822800;
      74942: inst = 32'h10a00000;
      74943: inst = 32'hca00004;
      74944: inst = 32'h38632800;
      74945: inst = 32'h38842800;
      74946: inst = 32'h10a00001;
      74947: inst = 32'hca024c7;
      74948: inst = 32'h13e00001;
      74949: inst = 32'hfe0d96a;
      74950: inst = 32'h5be00000;
      74951: inst = 32'h8c50000;
      74952: inst = 32'h24612800;
      74953: inst = 32'h10a0ffff;
      74954: inst = 32'hca0fffd;
      74955: inst = 32'h24822800;
      74956: inst = 32'h10a00000;
      74957: inst = 32'hca00004;
      74958: inst = 32'h38632800;
      74959: inst = 32'h38842800;
      74960: inst = 32'h10a00001;
      74961: inst = 32'hca024d5;
      74962: inst = 32'h13e00001;
      74963: inst = 32'hfe0d96a;
      74964: inst = 32'h5be00000;
      74965: inst = 32'h8c50000;
      74966: inst = 32'h24612800;
      74967: inst = 32'h10a0ffff;
      74968: inst = 32'hca0fffd;
      74969: inst = 32'h24822800;
      74970: inst = 32'h10a00000;
      74971: inst = 32'hca00004;
      74972: inst = 32'h38632800;
      74973: inst = 32'h38842800;
      74974: inst = 32'h10a00001;
      74975: inst = 32'hca024e3;
      74976: inst = 32'h13e00001;
      74977: inst = 32'hfe0d96a;
      74978: inst = 32'h5be00000;
      74979: inst = 32'h8c50000;
      74980: inst = 32'h24612800;
      74981: inst = 32'h10a0ffff;
      74982: inst = 32'hca0fffd;
      74983: inst = 32'h24822800;
      74984: inst = 32'h10a00000;
      74985: inst = 32'hca00004;
      74986: inst = 32'h38632800;
      74987: inst = 32'h38842800;
      74988: inst = 32'h10a00001;
      74989: inst = 32'hca024f1;
      74990: inst = 32'h13e00001;
      74991: inst = 32'hfe0d96a;
      74992: inst = 32'h5be00000;
      74993: inst = 32'h8c50000;
      74994: inst = 32'h24612800;
      74995: inst = 32'h10a0ffff;
      74996: inst = 32'hca0fffd;
      74997: inst = 32'h24822800;
      74998: inst = 32'h10a00000;
      74999: inst = 32'hca00004;
      75000: inst = 32'h38632800;
      75001: inst = 32'h38842800;
      75002: inst = 32'h10a00001;
      75003: inst = 32'hca024ff;
      75004: inst = 32'h13e00001;
      75005: inst = 32'hfe0d96a;
      75006: inst = 32'h5be00000;
      75007: inst = 32'h8c50000;
      75008: inst = 32'h24612800;
      75009: inst = 32'h10a0ffff;
      75010: inst = 32'hca0fffd;
      75011: inst = 32'h24822800;
      75012: inst = 32'h10a00000;
      75013: inst = 32'hca00004;
      75014: inst = 32'h38632800;
      75015: inst = 32'h38842800;
      75016: inst = 32'h10a00001;
      75017: inst = 32'hca0250d;
      75018: inst = 32'h13e00001;
      75019: inst = 32'hfe0d96a;
      75020: inst = 32'h5be00000;
      75021: inst = 32'h8c50000;
      75022: inst = 32'h24612800;
      75023: inst = 32'h10a0ffff;
      75024: inst = 32'hca0fffd;
      75025: inst = 32'h24822800;
      75026: inst = 32'h10a00000;
      75027: inst = 32'hca00004;
      75028: inst = 32'h38632800;
      75029: inst = 32'h38842800;
      75030: inst = 32'h10a00001;
      75031: inst = 32'hca0251b;
      75032: inst = 32'h13e00001;
      75033: inst = 32'hfe0d96a;
      75034: inst = 32'h5be00000;
      75035: inst = 32'h8c50000;
      75036: inst = 32'h24612800;
      75037: inst = 32'h10a0ffff;
      75038: inst = 32'hca0fffd;
      75039: inst = 32'h24822800;
      75040: inst = 32'h10a00000;
      75041: inst = 32'hca00004;
      75042: inst = 32'h38632800;
      75043: inst = 32'h38842800;
      75044: inst = 32'h10a00001;
      75045: inst = 32'hca02529;
      75046: inst = 32'h13e00001;
      75047: inst = 32'hfe0d96a;
      75048: inst = 32'h5be00000;
      75049: inst = 32'h8c50000;
      75050: inst = 32'h24612800;
      75051: inst = 32'h10a0ffff;
      75052: inst = 32'hca0fffd;
      75053: inst = 32'h24822800;
      75054: inst = 32'h10a00000;
      75055: inst = 32'hca00004;
      75056: inst = 32'h38632800;
      75057: inst = 32'h38842800;
      75058: inst = 32'h10a00001;
      75059: inst = 32'hca02537;
      75060: inst = 32'h13e00001;
      75061: inst = 32'hfe0d96a;
      75062: inst = 32'h5be00000;
      75063: inst = 32'h8c50000;
      75064: inst = 32'h24612800;
      75065: inst = 32'h10a0ffff;
      75066: inst = 32'hca0fffd;
      75067: inst = 32'h24822800;
      75068: inst = 32'h10a00000;
      75069: inst = 32'hca00004;
      75070: inst = 32'h38632800;
      75071: inst = 32'h38842800;
      75072: inst = 32'h10a00001;
      75073: inst = 32'hca02545;
      75074: inst = 32'h13e00001;
      75075: inst = 32'hfe0d96a;
      75076: inst = 32'h5be00000;
      75077: inst = 32'h8c50000;
      75078: inst = 32'h24612800;
      75079: inst = 32'h10a0ffff;
      75080: inst = 32'hca0fffd;
      75081: inst = 32'h24822800;
      75082: inst = 32'h10a00000;
      75083: inst = 32'hca00004;
      75084: inst = 32'h38632800;
      75085: inst = 32'h38842800;
      75086: inst = 32'h10a00001;
      75087: inst = 32'hca02553;
      75088: inst = 32'h13e00001;
      75089: inst = 32'hfe0d96a;
      75090: inst = 32'h5be00000;
      75091: inst = 32'h8c50000;
      75092: inst = 32'h24612800;
      75093: inst = 32'h10a0ffff;
      75094: inst = 32'hca0fffd;
      75095: inst = 32'h24822800;
      75096: inst = 32'h10a00000;
      75097: inst = 32'hca00004;
      75098: inst = 32'h38632800;
      75099: inst = 32'h38842800;
      75100: inst = 32'h10a00001;
      75101: inst = 32'hca02561;
      75102: inst = 32'h13e00001;
      75103: inst = 32'hfe0d96a;
      75104: inst = 32'h5be00000;
      75105: inst = 32'h8c50000;
      75106: inst = 32'h24612800;
      75107: inst = 32'h10a0ffff;
      75108: inst = 32'hca0fffd;
      75109: inst = 32'h24822800;
      75110: inst = 32'h10a00000;
      75111: inst = 32'hca00004;
      75112: inst = 32'h38632800;
      75113: inst = 32'h38842800;
      75114: inst = 32'h10a00001;
      75115: inst = 32'hca0256f;
      75116: inst = 32'h13e00001;
      75117: inst = 32'hfe0d96a;
      75118: inst = 32'h5be00000;
      75119: inst = 32'h8c50000;
      75120: inst = 32'h24612800;
      75121: inst = 32'h10a0ffff;
      75122: inst = 32'hca0fffd;
      75123: inst = 32'h24822800;
      75124: inst = 32'h10a00000;
      75125: inst = 32'hca00004;
      75126: inst = 32'h38632800;
      75127: inst = 32'h38842800;
      75128: inst = 32'h10a00001;
      75129: inst = 32'hca0257d;
      75130: inst = 32'h13e00001;
      75131: inst = 32'hfe0d96a;
      75132: inst = 32'h5be00000;
      75133: inst = 32'h8c50000;
      75134: inst = 32'h24612800;
      75135: inst = 32'h10a0ffff;
      75136: inst = 32'hca0fffd;
      75137: inst = 32'h24822800;
      75138: inst = 32'h10a00000;
      75139: inst = 32'hca00004;
      75140: inst = 32'h38632800;
      75141: inst = 32'h38842800;
      75142: inst = 32'h10a00001;
      75143: inst = 32'hca0258b;
      75144: inst = 32'h13e00001;
      75145: inst = 32'hfe0d96a;
      75146: inst = 32'h5be00000;
      75147: inst = 32'h8c50000;
      75148: inst = 32'h24612800;
      75149: inst = 32'h10a0ffff;
      75150: inst = 32'hca0fffd;
      75151: inst = 32'h24822800;
      75152: inst = 32'h10a00000;
      75153: inst = 32'hca00004;
      75154: inst = 32'h38632800;
      75155: inst = 32'h38842800;
      75156: inst = 32'h10a00001;
      75157: inst = 32'hca02599;
      75158: inst = 32'h13e00001;
      75159: inst = 32'hfe0d96a;
      75160: inst = 32'h5be00000;
      75161: inst = 32'h8c50000;
      75162: inst = 32'h24612800;
      75163: inst = 32'h10a0ffff;
      75164: inst = 32'hca0fffd;
      75165: inst = 32'h24822800;
      75166: inst = 32'h10a00000;
      75167: inst = 32'hca00004;
      75168: inst = 32'h38632800;
      75169: inst = 32'h38842800;
      75170: inst = 32'h10a00001;
      75171: inst = 32'hca025a7;
      75172: inst = 32'h13e00001;
      75173: inst = 32'hfe0d96a;
      75174: inst = 32'h5be00000;
      75175: inst = 32'h8c50000;
      75176: inst = 32'h24612800;
      75177: inst = 32'h10a0ffff;
      75178: inst = 32'hca0fffd;
      75179: inst = 32'h24822800;
      75180: inst = 32'h10a00000;
      75181: inst = 32'hca00004;
      75182: inst = 32'h38632800;
      75183: inst = 32'h38842800;
      75184: inst = 32'h10a00001;
      75185: inst = 32'hca025b5;
      75186: inst = 32'h13e00001;
      75187: inst = 32'hfe0d96a;
      75188: inst = 32'h5be00000;
      75189: inst = 32'h8c50000;
      75190: inst = 32'h24612800;
      75191: inst = 32'h10a0ffff;
      75192: inst = 32'hca0fffd;
      75193: inst = 32'h24822800;
      75194: inst = 32'h10a00000;
      75195: inst = 32'hca00004;
      75196: inst = 32'h38632800;
      75197: inst = 32'h38842800;
      75198: inst = 32'h10a00001;
      75199: inst = 32'hca025c3;
      75200: inst = 32'h13e00001;
      75201: inst = 32'hfe0d96a;
      75202: inst = 32'h5be00000;
      75203: inst = 32'h8c50000;
      75204: inst = 32'h24612800;
      75205: inst = 32'h10a0ffff;
      75206: inst = 32'hca0fffd;
      75207: inst = 32'h24822800;
      75208: inst = 32'h10a00000;
      75209: inst = 32'hca00004;
      75210: inst = 32'h38632800;
      75211: inst = 32'h38842800;
      75212: inst = 32'h10a00001;
      75213: inst = 32'hca025d1;
      75214: inst = 32'h13e00001;
      75215: inst = 32'hfe0d96a;
      75216: inst = 32'h5be00000;
      75217: inst = 32'h8c50000;
      75218: inst = 32'h24612800;
      75219: inst = 32'h10a0ffff;
      75220: inst = 32'hca0fffd;
      75221: inst = 32'h24822800;
      75222: inst = 32'h10a00000;
      75223: inst = 32'hca00004;
      75224: inst = 32'h38632800;
      75225: inst = 32'h38842800;
      75226: inst = 32'h10a00001;
      75227: inst = 32'hca025df;
      75228: inst = 32'h13e00001;
      75229: inst = 32'hfe0d96a;
      75230: inst = 32'h5be00000;
      75231: inst = 32'h8c50000;
      75232: inst = 32'h24612800;
      75233: inst = 32'h10a0ffff;
      75234: inst = 32'hca0fffd;
      75235: inst = 32'h24822800;
      75236: inst = 32'h10a00000;
      75237: inst = 32'hca00004;
      75238: inst = 32'h38632800;
      75239: inst = 32'h38842800;
      75240: inst = 32'h10a00001;
      75241: inst = 32'hca025ed;
      75242: inst = 32'h13e00001;
      75243: inst = 32'hfe0d96a;
      75244: inst = 32'h5be00000;
      75245: inst = 32'h8c50000;
      75246: inst = 32'h24612800;
      75247: inst = 32'h10a0ffff;
      75248: inst = 32'hca0fffd;
      75249: inst = 32'h24822800;
      75250: inst = 32'h10a00000;
      75251: inst = 32'hca00004;
      75252: inst = 32'h38632800;
      75253: inst = 32'h38842800;
      75254: inst = 32'h10a00001;
      75255: inst = 32'hca025fb;
      75256: inst = 32'h13e00001;
      75257: inst = 32'hfe0d96a;
      75258: inst = 32'h5be00000;
      75259: inst = 32'h8c50000;
      75260: inst = 32'h24612800;
      75261: inst = 32'h10a0ffff;
      75262: inst = 32'hca0fffd;
      75263: inst = 32'h24822800;
      75264: inst = 32'h10a00000;
      75265: inst = 32'hca00004;
      75266: inst = 32'h38632800;
      75267: inst = 32'h38842800;
      75268: inst = 32'h10a00001;
      75269: inst = 32'hca02609;
      75270: inst = 32'h13e00001;
      75271: inst = 32'hfe0d96a;
      75272: inst = 32'h5be00000;
      75273: inst = 32'h8c50000;
      75274: inst = 32'h24612800;
      75275: inst = 32'h10a0ffff;
      75276: inst = 32'hca0fffd;
      75277: inst = 32'h24822800;
      75278: inst = 32'h10a00000;
      75279: inst = 32'hca00004;
      75280: inst = 32'h38632800;
      75281: inst = 32'h38842800;
      75282: inst = 32'h10a00001;
      75283: inst = 32'hca02617;
      75284: inst = 32'h13e00001;
      75285: inst = 32'hfe0d96a;
      75286: inst = 32'h5be00000;
      75287: inst = 32'h8c50000;
      75288: inst = 32'h24612800;
      75289: inst = 32'h10a0ffff;
      75290: inst = 32'hca0fffd;
      75291: inst = 32'h24822800;
      75292: inst = 32'h10a00000;
      75293: inst = 32'hca00004;
      75294: inst = 32'h38632800;
      75295: inst = 32'h38842800;
      75296: inst = 32'h10a00001;
      75297: inst = 32'hca02625;
      75298: inst = 32'h13e00001;
      75299: inst = 32'hfe0d96a;
      75300: inst = 32'h5be00000;
      75301: inst = 32'h8c50000;
      75302: inst = 32'h24612800;
      75303: inst = 32'h10a0ffff;
      75304: inst = 32'hca0fffd;
      75305: inst = 32'h24822800;
      75306: inst = 32'h10a00000;
      75307: inst = 32'hca00004;
      75308: inst = 32'h38632800;
      75309: inst = 32'h38842800;
      75310: inst = 32'h10a00001;
      75311: inst = 32'hca02633;
      75312: inst = 32'h13e00001;
      75313: inst = 32'hfe0d96a;
      75314: inst = 32'h5be00000;
      75315: inst = 32'h8c50000;
      75316: inst = 32'h24612800;
      75317: inst = 32'h10a0ffff;
      75318: inst = 32'hca0fffd;
      75319: inst = 32'h24822800;
      75320: inst = 32'h10a00000;
      75321: inst = 32'hca00004;
      75322: inst = 32'h38632800;
      75323: inst = 32'h38842800;
      75324: inst = 32'h10a00001;
      75325: inst = 32'hca02641;
      75326: inst = 32'h13e00001;
      75327: inst = 32'hfe0d96a;
      75328: inst = 32'h5be00000;
      75329: inst = 32'h8c50000;
      75330: inst = 32'h24612800;
      75331: inst = 32'h10a0ffff;
      75332: inst = 32'hca0fffd;
      75333: inst = 32'h24822800;
      75334: inst = 32'h10a00000;
      75335: inst = 32'hca00004;
      75336: inst = 32'h38632800;
      75337: inst = 32'h38842800;
      75338: inst = 32'h10a00001;
      75339: inst = 32'hca0264f;
      75340: inst = 32'h13e00001;
      75341: inst = 32'hfe0d96a;
      75342: inst = 32'h5be00000;
      75343: inst = 32'h8c50000;
      75344: inst = 32'h24612800;
      75345: inst = 32'h10a0ffff;
      75346: inst = 32'hca0fffd;
      75347: inst = 32'h24822800;
      75348: inst = 32'h10a00000;
      75349: inst = 32'hca00004;
      75350: inst = 32'h38632800;
      75351: inst = 32'h38842800;
      75352: inst = 32'h10a00001;
      75353: inst = 32'hca0265d;
      75354: inst = 32'h13e00001;
      75355: inst = 32'hfe0d96a;
      75356: inst = 32'h5be00000;
      75357: inst = 32'h8c50000;
      75358: inst = 32'h24612800;
      75359: inst = 32'h10a0ffff;
      75360: inst = 32'hca0fffd;
      75361: inst = 32'h24822800;
      75362: inst = 32'h10a00000;
      75363: inst = 32'hca00004;
      75364: inst = 32'h38632800;
      75365: inst = 32'h38842800;
      75366: inst = 32'h10a00001;
      75367: inst = 32'hca0266b;
      75368: inst = 32'h13e00001;
      75369: inst = 32'hfe0d96a;
      75370: inst = 32'h5be00000;
      75371: inst = 32'h8c50000;
      75372: inst = 32'h24612800;
      75373: inst = 32'h10a0ffff;
      75374: inst = 32'hca0fffd;
      75375: inst = 32'h24822800;
      75376: inst = 32'h10a00000;
      75377: inst = 32'hca00004;
      75378: inst = 32'h38632800;
      75379: inst = 32'h38842800;
      75380: inst = 32'h10a00001;
      75381: inst = 32'hca02679;
      75382: inst = 32'h13e00001;
      75383: inst = 32'hfe0d96a;
      75384: inst = 32'h5be00000;
      75385: inst = 32'h8c50000;
      75386: inst = 32'h24612800;
      75387: inst = 32'h10a0ffff;
      75388: inst = 32'hca0fffd;
      75389: inst = 32'h24822800;
      75390: inst = 32'h10a00000;
      75391: inst = 32'hca00004;
      75392: inst = 32'h38632800;
      75393: inst = 32'h38842800;
      75394: inst = 32'h10a00001;
      75395: inst = 32'hca02687;
      75396: inst = 32'h13e00001;
      75397: inst = 32'hfe0d96a;
      75398: inst = 32'h5be00000;
      75399: inst = 32'h8c50000;
      75400: inst = 32'h24612800;
      75401: inst = 32'h10a0ffff;
      75402: inst = 32'hca0fffd;
      75403: inst = 32'h24822800;
      75404: inst = 32'h10a00000;
      75405: inst = 32'hca00004;
      75406: inst = 32'h38632800;
      75407: inst = 32'h38842800;
      75408: inst = 32'h10a00001;
      75409: inst = 32'hca02695;
      75410: inst = 32'h13e00001;
      75411: inst = 32'hfe0d96a;
      75412: inst = 32'h5be00000;
      75413: inst = 32'h8c50000;
      75414: inst = 32'h24612800;
      75415: inst = 32'h10a0ffff;
      75416: inst = 32'hca0fffd;
      75417: inst = 32'h24822800;
      75418: inst = 32'h10a00000;
      75419: inst = 32'hca00004;
      75420: inst = 32'h38632800;
      75421: inst = 32'h38842800;
      75422: inst = 32'h10a00001;
      75423: inst = 32'hca026a3;
      75424: inst = 32'h13e00001;
      75425: inst = 32'hfe0d96a;
      75426: inst = 32'h5be00000;
      75427: inst = 32'h8c50000;
      75428: inst = 32'h24612800;
      75429: inst = 32'h10a0ffff;
      75430: inst = 32'hca0fffd;
      75431: inst = 32'h24822800;
      75432: inst = 32'h10a00000;
      75433: inst = 32'hca00004;
      75434: inst = 32'h38632800;
      75435: inst = 32'h38842800;
      75436: inst = 32'h10a00001;
      75437: inst = 32'hca026b1;
      75438: inst = 32'h13e00001;
      75439: inst = 32'hfe0d96a;
      75440: inst = 32'h5be00000;
      75441: inst = 32'h8c50000;
      75442: inst = 32'h24612800;
      75443: inst = 32'h10a0ffff;
      75444: inst = 32'hca0fffd;
      75445: inst = 32'h24822800;
      75446: inst = 32'h10a00000;
      75447: inst = 32'hca00004;
      75448: inst = 32'h38632800;
      75449: inst = 32'h38842800;
      75450: inst = 32'h10a00001;
      75451: inst = 32'hca026bf;
      75452: inst = 32'h13e00001;
      75453: inst = 32'hfe0d96a;
      75454: inst = 32'h5be00000;
      75455: inst = 32'h8c50000;
      75456: inst = 32'h24612800;
      75457: inst = 32'h10a0ffff;
      75458: inst = 32'hca0fffd;
      75459: inst = 32'h24822800;
      75460: inst = 32'h10a00000;
      75461: inst = 32'hca00004;
      75462: inst = 32'h38632800;
      75463: inst = 32'h38842800;
      75464: inst = 32'h10a00001;
      75465: inst = 32'hca026cd;
      75466: inst = 32'h13e00001;
      75467: inst = 32'hfe0d96a;
      75468: inst = 32'h5be00000;
      75469: inst = 32'h8c50000;
      75470: inst = 32'h24612800;
      75471: inst = 32'h10a0ffff;
      75472: inst = 32'hca0fffd;
      75473: inst = 32'h24822800;
      75474: inst = 32'h10a00000;
      75475: inst = 32'hca00004;
      75476: inst = 32'h38632800;
      75477: inst = 32'h38842800;
      75478: inst = 32'h10a00001;
      75479: inst = 32'hca026db;
      75480: inst = 32'h13e00001;
      75481: inst = 32'hfe0d96a;
      75482: inst = 32'h5be00000;
      75483: inst = 32'h8c50000;
      75484: inst = 32'h24612800;
      75485: inst = 32'h10a0ffff;
      75486: inst = 32'hca0fffd;
      75487: inst = 32'h24822800;
      75488: inst = 32'h10a00000;
      75489: inst = 32'hca00004;
      75490: inst = 32'h38632800;
      75491: inst = 32'h38842800;
      75492: inst = 32'h10a00001;
      75493: inst = 32'hca026e9;
      75494: inst = 32'h13e00001;
      75495: inst = 32'hfe0d96a;
      75496: inst = 32'h5be00000;
      75497: inst = 32'h8c50000;
      75498: inst = 32'h24612800;
      75499: inst = 32'h10a0ffff;
      75500: inst = 32'hca0fffe;
      75501: inst = 32'h24822800;
      75502: inst = 32'h10a00000;
      75503: inst = 32'hca00004;
      75504: inst = 32'h38632800;
      75505: inst = 32'h38842800;
      75506: inst = 32'h10a00001;
      75507: inst = 32'hca026f7;
      75508: inst = 32'h13e00001;
      75509: inst = 32'hfe0d96a;
      75510: inst = 32'h5be00000;
      75511: inst = 32'h8c50000;
      75512: inst = 32'h24612800;
      75513: inst = 32'h10a0ffff;
      75514: inst = 32'hca0fffe;
      75515: inst = 32'h24822800;
      75516: inst = 32'h10a00000;
      75517: inst = 32'hca00004;
      75518: inst = 32'h38632800;
      75519: inst = 32'h38842800;
      75520: inst = 32'h10a00001;
      75521: inst = 32'hca02705;
      75522: inst = 32'h13e00001;
      75523: inst = 32'hfe0d96a;
      75524: inst = 32'h5be00000;
      75525: inst = 32'h8c50000;
      75526: inst = 32'h24612800;
      75527: inst = 32'h10a0ffff;
      75528: inst = 32'hca0fffe;
      75529: inst = 32'h24822800;
      75530: inst = 32'h10a00000;
      75531: inst = 32'hca00004;
      75532: inst = 32'h38632800;
      75533: inst = 32'h38842800;
      75534: inst = 32'h10a00001;
      75535: inst = 32'hca02713;
      75536: inst = 32'h13e00001;
      75537: inst = 32'hfe0d96a;
      75538: inst = 32'h5be00000;
      75539: inst = 32'h8c50000;
      75540: inst = 32'h24612800;
      75541: inst = 32'h10a0ffff;
      75542: inst = 32'hca0fffe;
      75543: inst = 32'h24822800;
      75544: inst = 32'h10a00000;
      75545: inst = 32'hca00004;
      75546: inst = 32'h38632800;
      75547: inst = 32'h38842800;
      75548: inst = 32'h10a00001;
      75549: inst = 32'hca02721;
      75550: inst = 32'h13e00001;
      75551: inst = 32'hfe0d96a;
      75552: inst = 32'h5be00000;
      75553: inst = 32'h8c50000;
      75554: inst = 32'h24612800;
      75555: inst = 32'h10a0ffff;
      75556: inst = 32'hca0fffe;
      75557: inst = 32'h24822800;
      75558: inst = 32'h10a00000;
      75559: inst = 32'hca00004;
      75560: inst = 32'h38632800;
      75561: inst = 32'h38842800;
      75562: inst = 32'h10a00001;
      75563: inst = 32'hca0272f;
      75564: inst = 32'h13e00001;
      75565: inst = 32'hfe0d96a;
      75566: inst = 32'h5be00000;
      75567: inst = 32'h8c50000;
      75568: inst = 32'h24612800;
      75569: inst = 32'h10a0ffff;
      75570: inst = 32'hca0fffe;
      75571: inst = 32'h24822800;
      75572: inst = 32'h10a00000;
      75573: inst = 32'hca00004;
      75574: inst = 32'h38632800;
      75575: inst = 32'h38842800;
      75576: inst = 32'h10a00001;
      75577: inst = 32'hca0273d;
      75578: inst = 32'h13e00001;
      75579: inst = 32'hfe0d96a;
      75580: inst = 32'h5be00000;
      75581: inst = 32'h8c50000;
      75582: inst = 32'h24612800;
      75583: inst = 32'h10a0ffff;
      75584: inst = 32'hca0fffe;
      75585: inst = 32'h24822800;
      75586: inst = 32'h10a00000;
      75587: inst = 32'hca00004;
      75588: inst = 32'h38632800;
      75589: inst = 32'h38842800;
      75590: inst = 32'h10a00001;
      75591: inst = 32'hca0274b;
      75592: inst = 32'h13e00001;
      75593: inst = 32'hfe0d96a;
      75594: inst = 32'h5be00000;
      75595: inst = 32'h8c50000;
      75596: inst = 32'h24612800;
      75597: inst = 32'h10a0ffff;
      75598: inst = 32'hca0fffe;
      75599: inst = 32'h24822800;
      75600: inst = 32'h10a00000;
      75601: inst = 32'hca00004;
      75602: inst = 32'h38632800;
      75603: inst = 32'h38842800;
      75604: inst = 32'h10a00001;
      75605: inst = 32'hca02759;
      75606: inst = 32'h13e00001;
      75607: inst = 32'hfe0d96a;
      75608: inst = 32'h5be00000;
      75609: inst = 32'h8c50000;
      75610: inst = 32'h24612800;
      75611: inst = 32'h10a0ffff;
      75612: inst = 32'hca0fffe;
      75613: inst = 32'h24822800;
      75614: inst = 32'h10a00000;
      75615: inst = 32'hca00004;
      75616: inst = 32'h38632800;
      75617: inst = 32'h38842800;
      75618: inst = 32'h10a00001;
      75619: inst = 32'hca02767;
      75620: inst = 32'h13e00001;
      75621: inst = 32'hfe0d96a;
      75622: inst = 32'h5be00000;
      75623: inst = 32'h8c50000;
      75624: inst = 32'h24612800;
      75625: inst = 32'h10a0ffff;
      75626: inst = 32'hca0fffe;
      75627: inst = 32'h24822800;
      75628: inst = 32'h10a00000;
      75629: inst = 32'hca00004;
      75630: inst = 32'h38632800;
      75631: inst = 32'h38842800;
      75632: inst = 32'h10a00001;
      75633: inst = 32'hca02775;
      75634: inst = 32'h13e00001;
      75635: inst = 32'hfe0d96a;
      75636: inst = 32'h5be00000;
      75637: inst = 32'h8c50000;
      75638: inst = 32'h24612800;
      75639: inst = 32'h10a0ffff;
      75640: inst = 32'hca0fffe;
      75641: inst = 32'h24822800;
      75642: inst = 32'h10a00000;
      75643: inst = 32'hca00004;
      75644: inst = 32'h38632800;
      75645: inst = 32'h38842800;
      75646: inst = 32'h10a00001;
      75647: inst = 32'hca02783;
      75648: inst = 32'h13e00001;
      75649: inst = 32'hfe0d96a;
      75650: inst = 32'h5be00000;
      75651: inst = 32'h8c50000;
      75652: inst = 32'h24612800;
      75653: inst = 32'h10a0ffff;
      75654: inst = 32'hca0fffe;
      75655: inst = 32'h24822800;
      75656: inst = 32'h10a00000;
      75657: inst = 32'hca00004;
      75658: inst = 32'h38632800;
      75659: inst = 32'h38842800;
      75660: inst = 32'h10a00001;
      75661: inst = 32'hca02791;
      75662: inst = 32'h13e00001;
      75663: inst = 32'hfe0d96a;
      75664: inst = 32'h5be00000;
      75665: inst = 32'h8c50000;
      75666: inst = 32'h24612800;
      75667: inst = 32'h10a0ffff;
      75668: inst = 32'hca0fffe;
      75669: inst = 32'h24822800;
      75670: inst = 32'h10a00000;
      75671: inst = 32'hca00004;
      75672: inst = 32'h38632800;
      75673: inst = 32'h38842800;
      75674: inst = 32'h10a00001;
      75675: inst = 32'hca0279f;
      75676: inst = 32'h13e00001;
      75677: inst = 32'hfe0d96a;
      75678: inst = 32'h5be00000;
      75679: inst = 32'h8c50000;
      75680: inst = 32'h24612800;
      75681: inst = 32'h10a0ffff;
      75682: inst = 32'hca0fffe;
      75683: inst = 32'h24822800;
      75684: inst = 32'h10a00000;
      75685: inst = 32'hca00004;
      75686: inst = 32'h38632800;
      75687: inst = 32'h38842800;
      75688: inst = 32'h10a00001;
      75689: inst = 32'hca027ad;
      75690: inst = 32'h13e00001;
      75691: inst = 32'hfe0d96a;
      75692: inst = 32'h5be00000;
      75693: inst = 32'h8c50000;
      75694: inst = 32'h24612800;
      75695: inst = 32'h10a0ffff;
      75696: inst = 32'hca0fffe;
      75697: inst = 32'h24822800;
      75698: inst = 32'h10a00000;
      75699: inst = 32'hca00004;
      75700: inst = 32'h38632800;
      75701: inst = 32'h38842800;
      75702: inst = 32'h10a00001;
      75703: inst = 32'hca027bb;
      75704: inst = 32'h13e00001;
      75705: inst = 32'hfe0d96a;
      75706: inst = 32'h5be00000;
      75707: inst = 32'h8c50000;
      75708: inst = 32'h24612800;
      75709: inst = 32'h10a0ffff;
      75710: inst = 32'hca0fffe;
      75711: inst = 32'h24822800;
      75712: inst = 32'h10a00000;
      75713: inst = 32'hca00004;
      75714: inst = 32'h38632800;
      75715: inst = 32'h38842800;
      75716: inst = 32'h10a00001;
      75717: inst = 32'hca027c9;
      75718: inst = 32'h13e00001;
      75719: inst = 32'hfe0d96a;
      75720: inst = 32'h5be00000;
      75721: inst = 32'h8c50000;
      75722: inst = 32'h24612800;
      75723: inst = 32'h10a0ffff;
      75724: inst = 32'hca0fffe;
      75725: inst = 32'h24822800;
      75726: inst = 32'h10a00000;
      75727: inst = 32'hca00004;
      75728: inst = 32'h38632800;
      75729: inst = 32'h38842800;
      75730: inst = 32'h10a00001;
      75731: inst = 32'hca027d7;
      75732: inst = 32'h13e00001;
      75733: inst = 32'hfe0d96a;
      75734: inst = 32'h5be00000;
      75735: inst = 32'h8c50000;
      75736: inst = 32'h24612800;
      75737: inst = 32'h10a0ffff;
      75738: inst = 32'hca0fffe;
      75739: inst = 32'h24822800;
      75740: inst = 32'h10a00000;
      75741: inst = 32'hca00004;
      75742: inst = 32'h38632800;
      75743: inst = 32'h38842800;
      75744: inst = 32'h10a00001;
      75745: inst = 32'hca027e5;
      75746: inst = 32'h13e00001;
      75747: inst = 32'hfe0d96a;
      75748: inst = 32'h5be00000;
      75749: inst = 32'h8c50000;
      75750: inst = 32'h24612800;
      75751: inst = 32'h10a0ffff;
      75752: inst = 32'hca0fffe;
      75753: inst = 32'h24822800;
      75754: inst = 32'h10a00000;
      75755: inst = 32'hca00004;
      75756: inst = 32'h38632800;
      75757: inst = 32'h38842800;
      75758: inst = 32'h10a00001;
      75759: inst = 32'hca027f3;
      75760: inst = 32'h13e00001;
      75761: inst = 32'hfe0d96a;
      75762: inst = 32'h5be00000;
      75763: inst = 32'h8c50000;
      75764: inst = 32'h24612800;
      75765: inst = 32'h10a0ffff;
      75766: inst = 32'hca0fffe;
      75767: inst = 32'h24822800;
      75768: inst = 32'h10a00000;
      75769: inst = 32'hca00004;
      75770: inst = 32'h38632800;
      75771: inst = 32'h38842800;
      75772: inst = 32'h10a00001;
      75773: inst = 32'hca02801;
      75774: inst = 32'h13e00001;
      75775: inst = 32'hfe0d96a;
      75776: inst = 32'h5be00000;
      75777: inst = 32'h8c50000;
      75778: inst = 32'h24612800;
      75779: inst = 32'h10a0ffff;
      75780: inst = 32'hca0fffe;
      75781: inst = 32'h24822800;
      75782: inst = 32'h10a00000;
      75783: inst = 32'hca00004;
      75784: inst = 32'h38632800;
      75785: inst = 32'h38842800;
      75786: inst = 32'h10a00001;
      75787: inst = 32'hca0280f;
      75788: inst = 32'h13e00001;
      75789: inst = 32'hfe0d96a;
      75790: inst = 32'h5be00000;
      75791: inst = 32'h8c50000;
      75792: inst = 32'h24612800;
      75793: inst = 32'h10a0ffff;
      75794: inst = 32'hca0fffe;
      75795: inst = 32'h24822800;
      75796: inst = 32'h10a00000;
      75797: inst = 32'hca00004;
      75798: inst = 32'h38632800;
      75799: inst = 32'h38842800;
      75800: inst = 32'h10a00001;
      75801: inst = 32'hca0281d;
      75802: inst = 32'h13e00001;
      75803: inst = 32'hfe0d96a;
      75804: inst = 32'h5be00000;
      75805: inst = 32'h8c50000;
      75806: inst = 32'h24612800;
      75807: inst = 32'h10a0ffff;
      75808: inst = 32'hca0fffe;
      75809: inst = 32'h24822800;
      75810: inst = 32'h10a00000;
      75811: inst = 32'hca00004;
      75812: inst = 32'h38632800;
      75813: inst = 32'h38842800;
      75814: inst = 32'h10a00001;
      75815: inst = 32'hca0282b;
      75816: inst = 32'h13e00001;
      75817: inst = 32'hfe0d96a;
      75818: inst = 32'h5be00000;
      75819: inst = 32'h8c50000;
      75820: inst = 32'h24612800;
      75821: inst = 32'h10a0ffff;
      75822: inst = 32'hca0fffe;
      75823: inst = 32'h24822800;
      75824: inst = 32'h10a00000;
      75825: inst = 32'hca00004;
      75826: inst = 32'h38632800;
      75827: inst = 32'h38842800;
      75828: inst = 32'h10a00001;
      75829: inst = 32'hca02839;
      75830: inst = 32'h13e00001;
      75831: inst = 32'hfe0d96a;
      75832: inst = 32'h5be00000;
      75833: inst = 32'h8c50000;
      75834: inst = 32'h24612800;
      75835: inst = 32'h10a0ffff;
      75836: inst = 32'hca0fffe;
      75837: inst = 32'h24822800;
      75838: inst = 32'h10a00000;
      75839: inst = 32'hca00004;
      75840: inst = 32'h38632800;
      75841: inst = 32'h38842800;
      75842: inst = 32'h10a00001;
      75843: inst = 32'hca02847;
      75844: inst = 32'h13e00001;
      75845: inst = 32'hfe0d96a;
      75846: inst = 32'h5be00000;
      75847: inst = 32'h8c50000;
      75848: inst = 32'h24612800;
      75849: inst = 32'h10a0ffff;
      75850: inst = 32'hca0fffe;
      75851: inst = 32'h24822800;
      75852: inst = 32'h10a00000;
      75853: inst = 32'hca00004;
      75854: inst = 32'h38632800;
      75855: inst = 32'h38842800;
      75856: inst = 32'h10a00001;
      75857: inst = 32'hca02855;
      75858: inst = 32'h13e00001;
      75859: inst = 32'hfe0d96a;
      75860: inst = 32'h5be00000;
      75861: inst = 32'h8c50000;
      75862: inst = 32'h24612800;
      75863: inst = 32'h10a0ffff;
      75864: inst = 32'hca0fffe;
      75865: inst = 32'h24822800;
      75866: inst = 32'h10a00000;
      75867: inst = 32'hca00004;
      75868: inst = 32'h38632800;
      75869: inst = 32'h38842800;
      75870: inst = 32'h10a00001;
      75871: inst = 32'hca02863;
      75872: inst = 32'h13e00001;
      75873: inst = 32'hfe0d96a;
      75874: inst = 32'h5be00000;
      75875: inst = 32'h8c50000;
      75876: inst = 32'h24612800;
      75877: inst = 32'h10a0ffff;
      75878: inst = 32'hca0fffe;
      75879: inst = 32'h24822800;
      75880: inst = 32'h10a00000;
      75881: inst = 32'hca00004;
      75882: inst = 32'h38632800;
      75883: inst = 32'h38842800;
      75884: inst = 32'h10a00001;
      75885: inst = 32'hca02871;
      75886: inst = 32'h13e00001;
      75887: inst = 32'hfe0d96a;
      75888: inst = 32'h5be00000;
      75889: inst = 32'h8c50000;
      75890: inst = 32'h24612800;
      75891: inst = 32'h10a0ffff;
      75892: inst = 32'hca0fffe;
      75893: inst = 32'h24822800;
      75894: inst = 32'h10a00000;
      75895: inst = 32'hca00004;
      75896: inst = 32'h38632800;
      75897: inst = 32'h38842800;
      75898: inst = 32'h10a00001;
      75899: inst = 32'hca0287f;
      75900: inst = 32'h13e00001;
      75901: inst = 32'hfe0d96a;
      75902: inst = 32'h5be00000;
      75903: inst = 32'h8c50000;
      75904: inst = 32'h24612800;
      75905: inst = 32'h10a0ffff;
      75906: inst = 32'hca0fffe;
      75907: inst = 32'h24822800;
      75908: inst = 32'h10a00000;
      75909: inst = 32'hca00004;
      75910: inst = 32'h38632800;
      75911: inst = 32'h38842800;
      75912: inst = 32'h10a00001;
      75913: inst = 32'hca0288d;
      75914: inst = 32'h13e00001;
      75915: inst = 32'hfe0d96a;
      75916: inst = 32'h5be00000;
      75917: inst = 32'h8c50000;
      75918: inst = 32'h24612800;
      75919: inst = 32'h10a0ffff;
      75920: inst = 32'hca0fffe;
      75921: inst = 32'h24822800;
      75922: inst = 32'h10a00000;
      75923: inst = 32'hca00004;
      75924: inst = 32'h38632800;
      75925: inst = 32'h38842800;
      75926: inst = 32'h10a00001;
      75927: inst = 32'hca0289b;
      75928: inst = 32'h13e00001;
      75929: inst = 32'hfe0d96a;
      75930: inst = 32'h5be00000;
      75931: inst = 32'h8c50000;
      75932: inst = 32'h24612800;
      75933: inst = 32'h10a0ffff;
      75934: inst = 32'hca0fffe;
      75935: inst = 32'h24822800;
      75936: inst = 32'h10a00000;
      75937: inst = 32'hca00004;
      75938: inst = 32'h38632800;
      75939: inst = 32'h38842800;
      75940: inst = 32'h10a00001;
      75941: inst = 32'hca028a9;
      75942: inst = 32'h13e00001;
      75943: inst = 32'hfe0d96a;
      75944: inst = 32'h5be00000;
      75945: inst = 32'h8c50000;
      75946: inst = 32'h24612800;
      75947: inst = 32'h10a0ffff;
      75948: inst = 32'hca0fffe;
      75949: inst = 32'h24822800;
      75950: inst = 32'h10a00000;
      75951: inst = 32'hca00004;
      75952: inst = 32'h38632800;
      75953: inst = 32'h38842800;
      75954: inst = 32'h10a00001;
      75955: inst = 32'hca028b7;
      75956: inst = 32'h13e00001;
      75957: inst = 32'hfe0d96a;
      75958: inst = 32'h5be00000;
      75959: inst = 32'h8c50000;
      75960: inst = 32'h24612800;
      75961: inst = 32'h10a0ffff;
      75962: inst = 32'hca0fffe;
      75963: inst = 32'h24822800;
      75964: inst = 32'h10a00000;
      75965: inst = 32'hca00004;
      75966: inst = 32'h38632800;
      75967: inst = 32'h38842800;
      75968: inst = 32'h10a00001;
      75969: inst = 32'hca028c5;
      75970: inst = 32'h13e00001;
      75971: inst = 32'hfe0d96a;
      75972: inst = 32'h5be00000;
      75973: inst = 32'h8c50000;
      75974: inst = 32'h24612800;
      75975: inst = 32'h10a0ffff;
      75976: inst = 32'hca0fffe;
      75977: inst = 32'h24822800;
      75978: inst = 32'h10a00000;
      75979: inst = 32'hca00004;
      75980: inst = 32'h38632800;
      75981: inst = 32'h38842800;
      75982: inst = 32'h10a00001;
      75983: inst = 32'hca028d3;
      75984: inst = 32'h13e00001;
      75985: inst = 32'hfe0d96a;
      75986: inst = 32'h5be00000;
      75987: inst = 32'h8c50000;
      75988: inst = 32'h24612800;
      75989: inst = 32'h10a0ffff;
      75990: inst = 32'hca0fffe;
      75991: inst = 32'h24822800;
      75992: inst = 32'h10a00000;
      75993: inst = 32'hca00004;
      75994: inst = 32'h38632800;
      75995: inst = 32'h38842800;
      75996: inst = 32'h10a00001;
      75997: inst = 32'hca028e1;
      75998: inst = 32'h13e00001;
      75999: inst = 32'hfe0d96a;
      76000: inst = 32'h5be00000;
      76001: inst = 32'h8c50000;
      76002: inst = 32'h24612800;
      76003: inst = 32'h10a0ffff;
      76004: inst = 32'hca0fffe;
      76005: inst = 32'h24822800;
      76006: inst = 32'h10a00000;
      76007: inst = 32'hca00004;
      76008: inst = 32'h38632800;
      76009: inst = 32'h38842800;
      76010: inst = 32'h10a00001;
      76011: inst = 32'hca028ef;
      76012: inst = 32'h13e00001;
      76013: inst = 32'hfe0d96a;
      76014: inst = 32'h5be00000;
      76015: inst = 32'h8c50000;
      76016: inst = 32'h24612800;
      76017: inst = 32'h10a0ffff;
      76018: inst = 32'hca0fffe;
      76019: inst = 32'h24822800;
      76020: inst = 32'h10a00000;
      76021: inst = 32'hca00004;
      76022: inst = 32'h38632800;
      76023: inst = 32'h38842800;
      76024: inst = 32'h10a00001;
      76025: inst = 32'hca028fd;
      76026: inst = 32'h13e00001;
      76027: inst = 32'hfe0d96a;
      76028: inst = 32'h5be00000;
      76029: inst = 32'h8c50000;
      76030: inst = 32'h24612800;
      76031: inst = 32'h10a0ffff;
      76032: inst = 32'hca0fffe;
      76033: inst = 32'h24822800;
      76034: inst = 32'h10a00000;
      76035: inst = 32'hca00004;
      76036: inst = 32'h38632800;
      76037: inst = 32'h38842800;
      76038: inst = 32'h10a00001;
      76039: inst = 32'hca0290b;
      76040: inst = 32'h13e00001;
      76041: inst = 32'hfe0d96a;
      76042: inst = 32'h5be00000;
      76043: inst = 32'h8c50000;
      76044: inst = 32'h24612800;
      76045: inst = 32'h10a0ffff;
      76046: inst = 32'hca0fffe;
      76047: inst = 32'h24822800;
      76048: inst = 32'h10a00000;
      76049: inst = 32'hca00004;
      76050: inst = 32'h38632800;
      76051: inst = 32'h38842800;
      76052: inst = 32'h10a00001;
      76053: inst = 32'hca02919;
      76054: inst = 32'h13e00001;
      76055: inst = 32'hfe0d96a;
      76056: inst = 32'h5be00000;
      76057: inst = 32'h8c50000;
      76058: inst = 32'h24612800;
      76059: inst = 32'h10a0ffff;
      76060: inst = 32'hca0fffe;
      76061: inst = 32'h24822800;
      76062: inst = 32'h10a00000;
      76063: inst = 32'hca00004;
      76064: inst = 32'h38632800;
      76065: inst = 32'h38842800;
      76066: inst = 32'h10a00001;
      76067: inst = 32'hca02927;
      76068: inst = 32'h13e00001;
      76069: inst = 32'hfe0d96a;
      76070: inst = 32'h5be00000;
      76071: inst = 32'h8c50000;
      76072: inst = 32'h24612800;
      76073: inst = 32'h10a0ffff;
      76074: inst = 32'hca0fffe;
      76075: inst = 32'h24822800;
      76076: inst = 32'h10a00000;
      76077: inst = 32'hca00004;
      76078: inst = 32'h38632800;
      76079: inst = 32'h38842800;
      76080: inst = 32'h10a00001;
      76081: inst = 32'hca02935;
      76082: inst = 32'h13e00001;
      76083: inst = 32'hfe0d96a;
      76084: inst = 32'h5be00000;
      76085: inst = 32'h8c50000;
      76086: inst = 32'h24612800;
      76087: inst = 32'h10a0ffff;
      76088: inst = 32'hca0fffe;
      76089: inst = 32'h24822800;
      76090: inst = 32'h10a00000;
      76091: inst = 32'hca00004;
      76092: inst = 32'h38632800;
      76093: inst = 32'h38842800;
      76094: inst = 32'h10a00001;
      76095: inst = 32'hca02943;
      76096: inst = 32'h13e00001;
      76097: inst = 32'hfe0d96a;
      76098: inst = 32'h5be00000;
      76099: inst = 32'h8c50000;
      76100: inst = 32'h24612800;
      76101: inst = 32'h10a0ffff;
      76102: inst = 32'hca0fffe;
      76103: inst = 32'h24822800;
      76104: inst = 32'h10a00000;
      76105: inst = 32'hca00004;
      76106: inst = 32'h38632800;
      76107: inst = 32'h38842800;
      76108: inst = 32'h10a00001;
      76109: inst = 32'hca02951;
      76110: inst = 32'h13e00001;
      76111: inst = 32'hfe0d96a;
      76112: inst = 32'h5be00000;
      76113: inst = 32'h8c50000;
      76114: inst = 32'h24612800;
      76115: inst = 32'h10a0ffff;
      76116: inst = 32'hca0fffe;
      76117: inst = 32'h24822800;
      76118: inst = 32'h10a00000;
      76119: inst = 32'hca00004;
      76120: inst = 32'h38632800;
      76121: inst = 32'h38842800;
      76122: inst = 32'h10a00001;
      76123: inst = 32'hca0295f;
      76124: inst = 32'h13e00001;
      76125: inst = 32'hfe0d96a;
      76126: inst = 32'h5be00000;
      76127: inst = 32'h8c50000;
      76128: inst = 32'h24612800;
      76129: inst = 32'h10a0ffff;
      76130: inst = 32'hca0fffe;
      76131: inst = 32'h24822800;
      76132: inst = 32'h10a00000;
      76133: inst = 32'hca00004;
      76134: inst = 32'h38632800;
      76135: inst = 32'h38842800;
      76136: inst = 32'h10a00001;
      76137: inst = 32'hca0296d;
      76138: inst = 32'h13e00001;
      76139: inst = 32'hfe0d96a;
      76140: inst = 32'h5be00000;
      76141: inst = 32'h8c50000;
      76142: inst = 32'h24612800;
      76143: inst = 32'h10a0ffff;
      76144: inst = 32'hca0fffe;
      76145: inst = 32'h24822800;
      76146: inst = 32'h10a00000;
      76147: inst = 32'hca00004;
      76148: inst = 32'h38632800;
      76149: inst = 32'h38842800;
      76150: inst = 32'h10a00001;
      76151: inst = 32'hca0297b;
      76152: inst = 32'h13e00001;
      76153: inst = 32'hfe0d96a;
      76154: inst = 32'h5be00000;
      76155: inst = 32'h8c50000;
      76156: inst = 32'h24612800;
      76157: inst = 32'h10a0ffff;
      76158: inst = 32'hca0fffe;
      76159: inst = 32'h24822800;
      76160: inst = 32'h10a00000;
      76161: inst = 32'hca00004;
      76162: inst = 32'h38632800;
      76163: inst = 32'h38842800;
      76164: inst = 32'h10a00001;
      76165: inst = 32'hca02989;
      76166: inst = 32'h13e00001;
      76167: inst = 32'hfe0d96a;
      76168: inst = 32'h5be00000;
      76169: inst = 32'h8c50000;
      76170: inst = 32'h24612800;
      76171: inst = 32'h10a0ffff;
      76172: inst = 32'hca0fffe;
      76173: inst = 32'h24822800;
      76174: inst = 32'h10a00000;
      76175: inst = 32'hca00004;
      76176: inst = 32'h38632800;
      76177: inst = 32'h38842800;
      76178: inst = 32'h10a00001;
      76179: inst = 32'hca02997;
      76180: inst = 32'h13e00001;
      76181: inst = 32'hfe0d96a;
      76182: inst = 32'h5be00000;
      76183: inst = 32'h8c50000;
      76184: inst = 32'h24612800;
      76185: inst = 32'h10a0ffff;
      76186: inst = 32'hca0fffe;
      76187: inst = 32'h24822800;
      76188: inst = 32'h10a00000;
      76189: inst = 32'hca00004;
      76190: inst = 32'h38632800;
      76191: inst = 32'h38842800;
      76192: inst = 32'h10a00001;
      76193: inst = 32'hca029a5;
      76194: inst = 32'h13e00001;
      76195: inst = 32'hfe0d96a;
      76196: inst = 32'h5be00000;
      76197: inst = 32'h8c50000;
      76198: inst = 32'h24612800;
      76199: inst = 32'h10a0ffff;
      76200: inst = 32'hca0fffe;
      76201: inst = 32'h24822800;
      76202: inst = 32'h10a00000;
      76203: inst = 32'hca00004;
      76204: inst = 32'h38632800;
      76205: inst = 32'h38842800;
      76206: inst = 32'h10a00001;
      76207: inst = 32'hca029b3;
      76208: inst = 32'h13e00001;
      76209: inst = 32'hfe0d96a;
      76210: inst = 32'h5be00000;
      76211: inst = 32'h8c50000;
      76212: inst = 32'h24612800;
      76213: inst = 32'h10a0ffff;
      76214: inst = 32'hca0fffe;
      76215: inst = 32'h24822800;
      76216: inst = 32'h10a00000;
      76217: inst = 32'hca00004;
      76218: inst = 32'h38632800;
      76219: inst = 32'h38842800;
      76220: inst = 32'h10a00001;
      76221: inst = 32'hca029c1;
      76222: inst = 32'h13e00001;
      76223: inst = 32'hfe0d96a;
      76224: inst = 32'h5be00000;
      76225: inst = 32'h8c50000;
      76226: inst = 32'h24612800;
      76227: inst = 32'h10a0ffff;
      76228: inst = 32'hca0fffe;
      76229: inst = 32'h24822800;
      76230: inst = 32'h10a00000;
      76231: inst = 32'hca00004;
      76232: inst = 32'h38632800;
      76233: inst = 32'h38842800;
      76234: inst = 32'h10a00001;
      76235: inst = 32'hca029cf;
      76236: inst = 32'h13e00001;
      76237: inst = 32'hfe0d96a;
      76238: inst = 32'h5be00000;
      76239: inst = 32'h8c50000;
      76240: inst = 32'h24612800;
      76241: inst = 32'h10a0ffff;
      76242: inst = 32'hca0fffe;
      76243: inst = 32'h24822800;
      76244: inst = 32'h10a00000;
      76245: inst = 32'hca00004;
      76246: inst = 32'h38632800;
      76247: inst = 32'h38842800;
      76248: inst = 32'h10a00001;
      76249: inst = 32'hca029dd;
      76250: inst = 32'h13e00001;
      76251: inst = 32'hfe0d96a;
      76252: inst = 32'h5be00000;
      76253: inst = 32'h8c50000;
      76254: inst = 32'h24612800;
      76255: inst = 32'h10a0ffff;
      76256: inst = 32'hca0fffe;
      76257: inst = 32'h24822800;
      76258: inst = 32'h10a00000;
      76259: inst = 32'hca00004;
      76260: inst = 32'h38632800;
      76261: inst = 32'h38842800;
      76262: inst = 32'h10a00001;
      76263: inst = 32'hca029eb;
      76264: inst = 32'h13e00001;
      76265: inst = 32'hfe0d96a;
      76266: inst = 32'h5be00000;
      76267: inst = 32'h8c50000;
      76268: inst = 32'h24612800;
      76269: inst = 32'h10a0ffff;
      76270: inst = 32'hca0fffe;
      76271: inst = 32'h24822800;
      76272: inst = 32'h10a00000;
      76273: inst = 32'hca00004;
      76274: inst = 32'h38632800;
      76275: inst = 32'h38842800;
      76276: inst = 32'h10a00001;
      76277: inst = 32'hca029f9;
      76278: inst = 32'h13e00001;
      76279: inst = 32'hfe0d96a;
      76280: inst = 32'h5be00000;
      76281: inst = 32'h8c50000;
      76282: inst = 32'h24612800;
      76283: inst = 32'h10a0ffff;
      76284: inst = 32'hca0fffe;
      76285: inst = 32'h24822800;
      76286: inst = 32'h10a00000;
      76287: inst = 32'hca00004;
      76288: inst = 32'h38632800;
      76289: inst = 32'h38842800;
      76290: inst = 32'h10a00001;
      76291: inst = 32'hca02a07;
      76292: inst = 32'h13e00001;
      76293: inst = 32'hfe0d96a;
      76294: inst = 32'h5be00000;
      76295: inst = 32'h8c50000;
      76296: inst = 32'h24612800;
      76297: inst = 32'h10a0ffff;
      76298: inst = 32'hca0fffe;
      76299: inst = 32'h24822800;
      76300: inst = 32'h10a00000;
      76301: inst = 32'hca00004;
      76302: inst = 32'h38632800;
      76303: inst = 32'h38842800;
      76304: inst = 32'h10a00001;
      76305: inst = 32'hca02a15;
      76306: inst = 32'h13e00001;
      76307: inst = 32'hfe0d96a;
      76308: inst = 32'h5be00000;
      76309: inst = 32'h8c50000;
      76310: inst = 32'h24612800;
      76311: inst = 32'h10a0ffff;
      76312: inst = 32'hca0fffe;
      76313: inst = 32'h24822800;
      76314: inst = 32'h10a00000;
      76315: inst = 32'hca00004;
      76316: inst = 32'h38632800;
      76317: inst = 32'h38842800;
      76318: inst = 32'h10a00001;
      76319: inst = 32'hca02a23;
      76320: inst = 32'h13e00001;
      76321: inst = 32'hfe0d96a;
      76322: inst = 32'h5be00000;
      76323: inst = 32'h8c50000;
      76324: inst = 32'h24612800;
      76325: inst = 32'h10a0ffff;
      76326: inst = 32'hca0fffe;
      76327: inst = 32'h24822800;
      76328: inst = 32'h10a00000;
      76329: inst = 32'hca00004;
      76330: inst = 32'h38632800;
      76331: inst = 32'h38842800;
      76332: inst = 32'h10a00001;
      76333: inst = 32'hca02a31;
      76334: inst = 32'h13e00001;
      76335: inst = 32'hfe0d96a;
      76336: inst = 32'h5be00000;
      76337: inst = 32'h8c50000;
      76338: inst = 32'h24612800;
      76339: inst = 32'h10a0ffff;
      76340: inst = 32'hca0fffe;
      76341: inst = 32'h24822800;
      76342: inst = 32'h10a00000;
      76343: inst = 32'hca00004;
      76344: inst = 32'h38632800;
      76345: inst = 32'h38842800;
      76346: inst = 32'h10a00001;
      76347: inst = 32'hca02a3f;
      76348: inst = 32'h13e00001;
      76349: inst = 32'hfe0d96a;
      76350: inst = 32'h5be00000;
      76351: inst = 32'h8c50000;
      76352: inst = 32'h24612800;
      76353: inst = 32'h10a0ffff;
      76354: inst = 32'hca0fffe;
      76355: inst = 32'h24822800;
      76356: inst = 32'h10a00000;
      76357: inst = 32'hca00004;
      76358: inst = 32'h38632800;
      76359: inst = 32'h38842800;
      76360: inst = 32'h10a00001;
      76361: inst = 32'hca02a4d;
      76362: inst = 32'h13e00001;
      76363: inst = 32'hfe0d96a;
      76364: inst = 32'h5be00000;
      76365: inst = 32'h8c50000;
      76366: inst = 32'h24612800;
      76367: inst = 32'h10a0ffff;
      76368: inst = 32'hca0fffe;
      76369: inst = 32'h24822800;
      76370: inst = 32'h10a00000;
      76371: inst = 32'hca00004;
      76372: inst = 32'h38632800;
      76373: inst = 32'h38842800;
      76374: inst = 32'h10a00001;
      76375: inst = 32'hca02a5b;
      76376: inst = 32'h13e00001;
      76377: inst = 32'hfe0d96a;
      76378: inst = 32'h5be00000;
      76379: inst = 32'h8c50000;
      76380: inst = 32'h24612800;
      76381: inst = 32'h10a0ffff;
      76382: inst = 32'hca0fffe;
      76383: inst = 32'h24822800;
      76384: inst = 32'h10a00000;
      76385: inst = 32'hca00004;
      76386: inst = 32'h38632800;
      76387: inst = 32'h38842800;
      76388: inst = 32'h10a00001;
      76389: inst = 32'hca02a69;
      76390: inst = 32'h13e00001;
      76391: inst = 32'hfe0d96a;
      76392: inst = 32'h5be00000;
      76393: inst = 32'h8c50000;
      76394: inst = 32'h24612800;
      76395: inst = 32'h10a0ffff;
      76396: inst = 32'hca0fffe;
      76397: inst = 32'h24822800;
      76398: inst = 32'h10a00000;
      76399: inst = 32'hca00004;
      76400: inst = 32'h38632800;
      76401: inst = 32'h38842800;
      76402: inst = 32'h10a00001;
      76403: inst = 32'hca02a77;
      76404: inst = 32'h13e00001;
      76405: inst = 32'hfe0d96a;
      76406: inst = 32'h5be00000;
      76407: inst = 32'h8c50000;
      76408: inst = 32'h24612800;
      76409: inst = 32'h10a0ffff;
      76410: inst = 32'hca0fffe;
      76411: inst = 32'h24822800;
      76412: inst = 32'h10a00000;
      76413: inst = 32'hca00004;
      76414: inst = 32'h38632800;
      76415: inst = 32'h38842800;
      76416: inst = 32'h10a00001;
      76417: inst = 32'hca02a85;
      76418: inst = 32'h13e00001;
      76419: inst = 32'hfe0d96a;
      76420: inst = 32'h5be00000;
      76421: inst = 32'h8c50000;
      76422: inst = 32'h24612800;
      76423: inst = 32'h10a0ffff;
      76424: inst = 32'hca0fffe;
      76425: inst = 32'h24822800;
      76426: inst = 32'h10a00000;
      76427: inst = 32'hca00004;
      76428: inst = 32'h38632800;
      76429: inst = 32'h38842800;
      76430: inst = 32'h10a00001;
      76431: inst = 32'hca02a93;
      76432: inst = 32'h13e00001;
      76433: inst = 32'hfe0d96a;
      76434: inst = 32'h5be00000;
      76435: inst = 32'h8c50000;
      76436: inst = 32'h24612800;
      76437: inst = 32'h10a0ffff;
      76438: inst = 32'hca0fffe;
      76439: inst = 32'h24822800;
      76440: inst = 32'h10a00000;
      76441: inst = 32'hca00004;
      76442: inst = 32'h38632800;
      76443: inst = 32'h38842800;
      76444: inst = 32'h10a00001;
      76445: inst = 32'hca02aa1;
      76446: inst = 32'h13e00001;
      76447: inst = 32'hfe0d96a;
      76448: inst = 32'h5be00000;
      76449: inst = 32'h8c50000;
      76450: inst = 32'h24612800;
      76451: inst = 32'h10a0ffff;
      76452: inst = 32'hca0fffe;
      76453: inst = 32'h24822800;
      76454: inst = 32'h10a00000;
      76455: inst = 32'hca00004;
      76456: inst = 32'h38632800;
      76457: inst = 32'h38842800;
      76458: inst = 32'h10a00001;
      76459: inst = 32'hca02aaf;
      76460: inst = 32'h13e00001;
      76461: inst = 32'hfe0d96a;
      76462: inst = 32'h5be00000;
      76463: inst = 32'h8c50000;
      76464: inst = 32'h24612800;
      76465: inst = 32'h10a0ffff;
      76466: inst = 32'hca0fffe;
      76467: inst = 32'h24822800;
      76468: inst = 32'h10a00000;
      76469: inst = 32'hca00004;
      76470: inst = 32'h38632800;
      76471: inst = 32'h38842800;
      76472: inst = 32'h10a00001;
      76473: inst = 32'hca02abd;
      76474: inst = 32'h13e00001;
      76475: inst = 32'hfe0d96a;
      76476: inst = 32'h5be00000;
      76477: inst = 32'h8c50000;
      76478: inst = 32'h24612800;
      76479: inst = 32'h10a0ffff;
      76480: inst = 32'hca0fffe;
      76481: inst = 32'h24822800;
      76482: inst = 32'h10a00000;
      76483: inst = 32'hca00004;
      76484: inst = 32'h38632800;
      76485: inst = 32'h38842800;
      76486: inst = 32'h10a00001;
      76487: inst = 32'hca02acb;
      76488: inst = 32'h13e00001;
      76489: inst = 32'hfe0d96a;
      76490: inst = 32'h5be00000;
      76491: inst = 32'h8c50000;
      76492: inst = 32'h24612800;
      76493: inst = 32'h10a0ffff;
      76494: inst = 32'hca0fffe;
      76495: inst = 32'h24822800;
      76496: inst = 32'h10a00000;
      76497: inst = 32'hca00004;
      76498: inst = 32'h38632800;
      76499: inst = 32'h38842800;
      76500: inst = 32'h10a00001;
      76501: inst = 32'hca02ad9;
      76502: inst = 32'h13e00001;
      76503: inst = 32'hfe0d96a;
      76504: inst = 32'h5be00000;
      76505: inst = 32'h8c50000;
      76506: inst = 32'h24612800;
      76507: inst = 32'h10a0ffff;
      76508: inst = 32'hca0fffe;
      76509: inst = 32'h24822800;
      76510: inst = 32'h10a00000;
      76511: inst = 32'hca00004;
      76512: inst = 32'h38632800;
      76513: inst = 32'h38842800;
      76514: inst = 32'h10a00001;
      76515: inst = 32'hca02ae7;
      76516: inst = 32'h13e00001;
      76517: inst = 32'hfe0d96a;
      76518: inst = 32'h5be00000;
      76519: inst = 32'h8c50000;
      76520: inst = 32'h24612800;
      76521: inst = 32'h10a0ffff;
      76522: inst = 32'hca0fffe;
      76523: inst = 32'h24822800;
      76524: inst = 32'h10a00000;
      76525: inst = 32'hca00004;
      76526: inst = 32'h38632800;
      76527: inst = 32'h38842800;
      76528: inst = 32'h10a00001;
      76529: inst = 32'hca02af5;
      76530: inst = 32'h13e00001;
      76531: inst = 32'hfe0d96a;
      76532: inst = 32'h5be00000;
      76533: inst = 32'h8c50000;
      76534: inst = 32'h24612800;
      76535: inst = 32'h10a0ffff;
      76536: inst = 32'hca0fffe;
      76537: inst = 32'h24822800;
      76538: inst = 32'h10a00000;
      76539: inst = 32'hca00004;
      76540: inst = 32'h38632800;
      76541: inst = 32'h38842800;
      76542: inst = 32'h10a00001;
      76543: inst = 32'hca02b03;
      76544: inst = 32'h13e00001;
      76545: inst = 32'hfe0d96a;
      76546: inst = 32'h5be00000;
      76547: inst = 32'h8c50000;
      76548: inst = 32'h24612800;
      76549: inst = 32'h10a0ffff;
      76550: inst = 32'hca0fffe;
      76551: inst = 32'h24822800;
      76552: inst = 32'h10a00000;
      76553: inst = 32'hca00004;
      76554: inst = 32'h38632800;
      76555: inst = 32'h38842800;
      76556: inst = 32'h10a00001;
      76557: inst = 32'hca02b11;
      76558: inst = 32'h13e00001;
      76559: inst = 32'hfe0d96a;
      76560: inst = 32'h5be00000;
      76561: inst = 32'h8c50000;
      76562: inst = 32'h24612800;
      76563: inst = 32'h10a0ffff;
      76564: inst = 32'hca0fffe;
      76565: inst = 32'h24822800;
      76566: inst = 32'h10a00000;
      76567: inst = 32'hca00004;
      76568: inst = 32'h38632800;
      76569: inst = 32'h38842800;
      76570: inst = 32'h10a00001;
      76571: inst = 32'hca02b1f;
      76572: inst = 32'h13e00001;
      76573: inst = 32'hfe0d96a;
      76574: inst = 32'h5be00000;
      76575: inst = 32'h8c50000;
      76576: inst = 32'h24612800;
      76577: inst = 32'h10a0ffff;
      76578: inst = 32'hca0fffe;
      76579: inst = 32'h24822800;
      76580: inst = 32'h10a00000;
      76581: inst = 32'hca00004;
      76582: inst = 32'h38632800;
      76583: inst = 32'h38842800;
      76584: inst = 32'h10a00001;
      76585: inst = 32'hca02b2d;
      76586: inst = 32'h13e00001;
      76587: inst = 32'hfe0d96a;
      76588: inst = 32'h5be00000;
      76589: inst = 32'h8c50000;
      76590: inst = 32'h24612800;
      76591: inst = 32'h10a0ffff;
      76592: inst = 32'hca0fffe;
      76593: inst = 32'h24822800;
      76594: inst = 32'h10a00000;
      76595: inst = 32'hca00004;
      76596: inst = 32'h38632800;
      76597: inst = 32'h38842800;
      76598: inst = 32'h10a00001;
      76599: inst = 32'hca02b3b;
      76600: inst = 32'h13e00001;
      76601: inst = 32'hfe0d96a;
      76602: inst = 32'h5be00000;
      76603: inst = 32'h8c50000;
      76604: inst = 32'h24612800;
      76605: inst = 32'h10a0ffff;
      76606: inst = 32'hca0fffe;
      76607: inst = 32'h24822800;
      76608: inst = 32'h10a00000;
      76609: inst = 32'hca00004;
      76610: inst = 32'h38632800;
      76611: inst = 32'h38842800;
      76612: inst = 32'h10a00001;
      76613: inst = 32'hca02b49;
      76614: inst = 32'h13e00001;
      76615: inst = 32'hfe0d96a;
      76616: inst = 32'h5be00000;
      76617: inst = 32'h8c50000;
      76618: inst = 32'h24612800;
      76619: inst = 32'h10a0ffff;
      76620: inst = 32'hca0fffe;
      76621: inst = 32'h24822800;
      76622: inst = 32'h10a00000;
      76623: inst = 32'hca00004;
      76624: inst = 32'h38632800;
      76625: inst = 32'h38842800;
      76626: inst = 32'h10a00001;
      76627: inst = 32'hca02b57;
      76628: inst = 32'h13e00001;
      76629: inst = 32'hfe0d96a;
      76630: inst = 32'h5be00000;
      76631: inst = 32'h8c50000;
      76632: inst = 32'h24612800;
      76633: inst = 32'h10a0ffff;
      76634: inst = 32'hca0fffe;
      76635: inst = 32'h24822800;
      76636: inst = 32'h10a00000;
      76637: inst = 32'hca00004;
      76638: inst = 32'h38632800;
      76639: inst = 32'h38842800;
      76640: inst = 32'h10a00001;
      76641: inst = 32'hca02b65;
      76642: inst = 32'h13e00001;
      76643: inst = 32'hfe0d96a;
      76644: inst = 32'h5be00000;
      76645: inst = 32'h8c50000;
      76646: inst = 32'h24612800;
      76647: inst = 32'h10a0ffff;
      76648: inst = 32'hca0fffe;
      76649: inst = 32'h24822800;
      76650: inst = 32'h10a00000;
      76651: inst = 32'hca00004;
      76652: inst = 32'h38632800;
      76653: inst = 32'h38842800;
      76654: inst = 32'h10a00001;
      76655: inst = 32'hca02b73;
      76656: inst = 32'h13e00001;
      76657: inst = 32'hfe0d96a;
      76658: inst = 32'h5be00000;
      76659: inst = 32'h8c50000;
      76660: inst = 32'h24612800;
      76661: inst = 32'h10a0ffff;
      76662: inst = 32'hca0fffe;
      76663: inst = 32'h24822800;
      76664: inst = 32'h10a00000;
      76665: inst = 32'hca00004;
      76666: inst = 32'h38632800;
      76667: inst = 32'h38842800;
      76668: inst = 32'h10a00001;
      76669: inst = 32'hca02b81;
      76670: inst = 32'h13e00001;
      76671: inst = 32'hfe0d96a;
      76672: inst = 32'h5be00000;
      76673: inst = 32'h8c50000;
      76674: inst = 32'h24612800;
      76675: inst = 32'h10a0ffff;
      76676: inst = 32'hca0fffe;
      76677: inst = 32'h24822800;
      76678: inst = 32'h10a00000;
      76679: inst = 32'hca00004;
      76680: inst = 32'h38632800;
      76681: inst = 32'h38842800;
      76682: inst = 32'h10a00001;
      76683: inst = 32'hca02b8f;
      76684: inst = 32'h13e00001;
      76685: inst = 32'hfe0d96a;
      76686: inst = 32'h5be00000;
      76687: inst = 32'h8c50000;
      76688: inst = 32'h24612800;
      76689: inst = 32'h10a0ffff;
      76690: inst = 32'hca0fffe;
      76691: inst = 32'h24822800;
      76692: inst = 32'h10a00000;
      76693: inst = 32'hca00004;
      76694: inst = 32'h38632800;
      76695: inst = 32'h38842800;
      76696: inst = 32'h10a00001;
      76697: inst = 32'hca02b9d;
      76698: inst = 32'h13e00001;
      76699: inst = 32'hfe0d96a;
      76700: inst = 32'h5be00000;
      76701: inst = 32'h8c50000;
      76702: inst = 32'h24612800;
      76703: inst = 32'h10a0ffff;
      76704: inst = 32'hca0fffe;
      76705: inst = 32'h24822800;
      76706: inst = 32'h10a00000;
      76707: inst = 32'hca00004;
      76708: inst = 32'h38632800;
      76709: inst = 32'h38842800;
      76710: inst = 32'h10a00001;
      76711: inst = 32'hca02bab;
      76712: inst = 32'h13e00001;
      76713: inst = 32'hfe0d96a;
      76714: inst = 32'h5be00000;
      76715: inst = 32'h8c50000;
      76716: inst = 32'h24612800;
      76717: inst = 32'h10a0ffff;
      76718: inst = 32'hca0fffe;
      76719: inst = 32'h24822800;
      76720: inst = 32'h10a00000;
      76721: inst = 32'hca00004;
      76722: inst = 32'h38632800;
      76723: inst = 32'h38842800;
      76724: inst = 32'h10a00001;
      76725: inst = 32'hca02bb9;
      76726: inst = 32'h13e00001;
      76727: inst = 32'hfe0d96a;
      76728: inst = 32'h5be00000;
      76729: inst = 32'h8c50000;
      76730: inst = 32'h24612800;
      76731: inst = 32'h10a0ffff;
      76732: inst = 32'hca0fffe;
      76733: inst = 32'h24822800;
      76734: inst = 32'h10a00000;
      76735: inst = 32'hca00004;
      76736: inst = 32'h38632800;
      76737: inst = 32'h38842800;
      76738: inst = 32'h10a00001;
      76739: inst = 32'hca02bc7;
      76740: inst = 32'h13e00001;
      76741: inst = 32'hfe0d96a;
      76742: inst = 32'h5be00000;
      76743: inst = 32'h8c50000;
      76744: inst = 32'h24612800;
      76745: inst = 32'h10a0ffff;
      76746: inst = 32'hca0fffe;
      76747: inst = 32'h24822800;
      76748: inst = 32'h10a00000;
      76749: inst = 32'hca00004;
      76750: inst = 32'h38632800;
      76751: inst = 32'h38842800;
      76752: inst = 32'h10a00001;
      76753: inst = 32'hca02bd5;
      76754: inst = 32'h13e00001;
      76755: inst = 32'hfe0d96a;
      76756: inst = 32'h5be00000;
      76757: inst = 32'h8c50000;
      76758: inst = 32'h24612800;
      76759: inst = 32'h10a0ffff;
      76760: inst = 32'hca0fffe;
      76761: inst = 32'h24822800;
      76762: inst = 32'h10a00000;
      76763: inst = 32'hca00004;
      76764: inst = 32'h38632800;
      76765: inst = 32'h38842800;
      76766: inst = 32'h10a00001;
      76767: inst = 32'hca02be3;
      76768: inst = 32'h13e00001;
      76769: inst = 32'hfe0d96a;
      76770: inst = 32'h5be00000;
      76771: inst = 32'h8c50000;
      76772: inst = 32'h24612800;
      76773: inst = 32'h10a0ffff;
      76774: inst = 32'hca0fffe;
      76775: inst = 32'h24822800;
      76776: inst = 32'h10a00000;
      76777: inst = 32'hca00004;
      76778: inst = 32'h38632800;
      76779: inst = 32'h38842800;
      76780: inst = 32'h10a00001;
      76781: inst = 32'hca02bf1;
      76782: inst = 32'h13e00001;
      76783: inst = 32'hfe0d96a;
      76784: inst = 32'h5be00000;
      76785: inst = 32'h8c50000;
      76786: inst = 32'h24612800;
      76787: inst = 32'h10a0ffff;
      76788: inst = 32'hca0fffe;
      76789: inst = 32'h24822800;
      76790: inst = 32'h10a00000;
      76791: inst = 32'hca00004;
      76792: inst = 32'h38632800;
      76793: inst = 32'h38842800;
      76794: inst = 32'h10a00001;
      76795: inst = 32'hca02bff;
      76796: inst = 32'h13e00001;
      76797: inst = 32'hfe0d96a;
      76798: inst = 32'h5be00000;
      76799: inst = 32'h8c50000;
      76800: inst = 32'h24612800;
      76801: inst = 32'h10a0ffff;
      76802: inst = 32'hca0fffe;
      76803: inst = 32'h24822800;
      76804: inst = 32'h10a00000;
      76805: inst = 32'hca00004;
      76806: inst = 32'h38632800;
      76807: inst = 32'h38842800;
      76808: inst = 32'h10a00001;
      76809: inst = 32'hca02c0d;
      76810: inst = 32'h13e00001;
      76811: inst = 32'hfe0d96a;
      76812: inst = 32'h5be00000;
      76813: inst = 32'h8c50000;
      76814: inst = 32'h24612800;
      76815: inst = 32'h10a0ffff;
      76816: inst = 32'hca0fffe;
      76817: inst = 32'h24822800;
      76818: inst = 32'h10a00000;
      76819: inst = 32'hca00004;
      76820: inst = 32'h38632800;
      76821: inst = 32'h38842800;
      76822: inst = 32'h10a00001;
      76823: inst = 32'hca02c1b;
      76824: inst = 32'h13e00001;
      76825: inst = 32'hfe0d96a;
      76826: inst = 32'h5be00000;
      76827: inst = 32'h8c50000;
      76828: inst = 32'h24612800;
      76829: inst = 32'h10a0ffff;
      76830: inst = 32'hca0fffe;
      76831: inst = 32'h24822800;
      76832: inst = 32'h10a00000;
      76833: inst = 32'hca00004;
      76834: inst = 32'h38632800;
      76835: inst = 32'h38842800;
      76836: inst = 32'h10a00001;
      76837: inst = 32'hca02c29;
      76838: inst = 32'h13e00001;
      76839: inst = 32'hfe0d96a;
      76840: inst = 32'h5be00000;
      76841: inst = 32'h8c50000;
      76842: inst = 32'h24612800;
      76843: inst = 32'h10a0ffff;
      76844: inst = 32'hca0ffff;
      76845: inst = 32'h24822800;
      76846: inst = 32'h10a00000;
      76847: inst = 32'hca00004;
      76848: inst = 32'h38632800;
      76849: inst = 32'h38842800;
      76850: inst = 32'h10a00001;
      76851: inst = 32'hca02c37;
      76852: inst = 32'h13e00001;
      76853: inst = 32'hfe0d96a;
      76854: inst = 32'h5be00000;
      76855: inst = 32'h8c50000;
      76856: inst = 32'h24612800;
      76857: inst = 32'h10a0ffff;
      76858: inst = 32'hca0ffff;
      76859: inst = 32'h24822800;
      76860: inst = 32'h10a00000;
      76861: inst = 32'hca00004;
      76862: inst = 32'h38632800;
      76863: inst = 32'h38842800;
      76864: inst = 32'h10a00001;
      76865: inst = 32'hca02c45;
      76866: inst = 32'h13e00001;
      76867: inst = 32'hfe0d96a;
      76868: inst = 32'h5be00000;
      76869: inst = 32'h8c50000;
      76870: inst = 32'h24612800;
      76871: inst = 32'h10a0ffff;
      76872: inst = 32'hca0ffff;
      76873: inst = 32'h24822800;
      76874: inst = 32'h10a00000;
      76875: inst = 32'hca00004;
      76876: inst = 32'h38632800;
      76877: inst = 32'h38842800;
      76878: inst = 32'h10a00001;
      76879: inst = 32'hca02c53;
      76880: inst = 32'h13e00001;
      76881: inst = 32'hfe0d96a;
      76882: inst = 32'h5be00000;
      76883: inst = 32'h8c50000;
      76884: inst = 32'h24612800;
      76885: inst = 32'h10a0ffff;
      76886: inst = 32'hca0ffff;
      76887: inst = 32'h24822800;
      76888: inst = 32'h10a00000;
      76889: inst = 32'hca00004;
      76890: inst = 32'h38632800;
      76891: inst = 32'h38842800;
      76892: inst = 32'h10a00001;
      76893: inst = 32'hca02c61;
      76894: inst = 32'h13e00001;
      76895: inst = 32'hfe0d96a;
      76896: inst = 32'h5be00000;
      76897: inst = 32'h8c50000;
      76898: inst = 32'h24612800;
      76899: inst = 32'h10a0ffff;
      76900: inst = 32'hca0ffff;
      76901: inst = 32'h24822800;
      76902: inst = 32'h10a00000;
      76903: inst = 32'hca00004;
      76904: inst = 32'h38632800;
      76905: inst = 32'h38842800;
      76906: inst = 32'h10a00001;
      76907: inst = 32'hca02c6f;
      76908: inst = 32'h13e00001;
      76909: inst = 32'hfe0d96a;
      76910: inst = 32'h5be00000;
      76911: inst = 32'h8c50000;
      76912: inst = 32'h24612800;
      76913: inst = 32'h10a0ffff;
      76914: inst = 32'hca0ffff;
      76915: inst = 32'h24822800;
      76916: inst = 32'h10a00000;
      76917: inst = 32'hca00004;
      76918: inst = 32'h38632800;
      76919: inst = 32'h38842800;
      76920: inst = 32'h10a00001;
      76921: inst = 32'hca02c7d;
      76922: inst = 32'h13e00001;
      76923: inst = 32'hfe0d96a;
      76924: inst = 32'h5be00000;
      76925: inst = 32'h8c50000;
      76926: inst = 32'h24612800;
      76927: inst = 32'h10a0ffff;
      76928: inst = 32'hca0ffff;
      76929: inst = 32'h24822800;
      76930: inst = 32'h10a00000;
      76931: inst = 32'hca00004;
      76932: inst = 32'h38632800;
      76933: inst = 32'h38842800;
      76934: inst = 32'h10a00001;
      76935: inst = 32'hca02c8b;
      76936: inst = 32'h13e00001;
      76937: inst = 32'hfe0d96a;
      76938: inst = 32'h5be00000;
      76939: inst = 32'h8c50000;
      76940: inst = 32'h24612800;
      76941: inst = 32'h10a0ffff;
      76942: inst = 32'hca0ffff;
      76943: inst = 32'h24822800;
      76944: inst = 32'h10a00000;
      76945: inst = 32'hca00004;
      76946: inst = 32'h38632800;
      76947: inst = 32'h38842800;
      76948: inst = 32'h10a00001;
      76949: inst = 32'hca02c99;
      76950: inst = 32'h13e00001;
      76951: inst = 32'hfe0d96a;
      76952: inst = 32'h5be00000;
      76953: inst = 32'h8c50000;
      76954: inst = 32'h24612800;
      76955: inst = 32'h10a0ffff;
      76956: inst = 32'hca0ffff;
      76957: inst = 32'h24822800;
      76958: inst = 32'h10a00000;
      76959: inst = 32'hca00004;
      76960: inst = 32'h38632800;
      76961: inst = 32'h38842800;
      76962: inst = 32'h10a00001;
      76963: inst = 32'hca02ca7;
      76964: inst = 32'h13e00001;
      76965: inst = 32'hfe0d96a;
      76966: inst = 32'h5be00000;
      76967: inst = 32'h8c50000;
      76968: inst = 32'h24612800;
      76969: inst = 32'h10a0ffff;
      76970: inst = 32'hca0ffff;
      76971: inst = 32'h24822800;
      76972: inst = 32'h10a00000;
      76973: inst = 32'hca00004;
      76974: inst = 32'h38632800;
      76975: inst = 32'h38842800;
      76976: inst = 32'h10a00001;
      76977: inst = 32'hca02cb5;
      76978: inst = 32'h13e00001;
      76979: inst = 32'hfe0d96a;
      76980: inst = 32'h5be00000;
      76981: inst = 32'h8c50000;
      76982: inst = 32'h24612800;
      76983: inst = 32'h10a0ffff;
      76984: inst = 32'hca0ffff;
      76985: inst = 32'h24822800;
      76986: inst = 32'h10a00000;
      76987: inst = 32'hca00004;
      76988: inst = 32'h38632800;
      76989: inst = 32'h38842800;
      76990: inst = 32'h10a00001;
      76991: inst = 32'hca02cc3;
      76992: inst = 32'h13e00001;
      76993: inst = 32'hfe0d96a;
      76994: inst = 32'h5be00000;
      76995: inst = 32'h8c50000;
      76996: inst = 32'h24612800;
      76997: inst = 32'h10a0ffff;
      76998: inst = 32'hca0ffff;
      76999: inst = 32'h24822800;
      77000: inst = 32'h10a00000;
      77001: inst = 32'hca00004;
      77002: inst = 32'h38632800;
      77003: inst = 32'h38842800;
      77004: inst = 32'h10a00001;
      77005: inst = 32'hca02cd1;
      77006: inst = 32'h13e00001;
      77007: inst = 32'hfe0d96a;
      77008: inst = 32'h5be00000;
      77009: inst = 32'h8c50000;
      77010: inst = 32'h24612800;
      77011: inst = 32'h10a0ffff;
      77012: inst = 32'hca0ffff;
      77013: inst = 32'h24822800;
      77014: inst = 32'h10a00000;
      77015: inst = 32'hca00004;
      77016: inst = 32'h38632800;
      77017: inst = 32'h38842800;
      77018: inst = 32'h10a00001;
      77019: inst = 32'hca02cdf;
      77020: inst = 32'h13e00001;
      77021: inst = 32'hfe0d96a;
      77022: inst = 32'h5be00000;
      77023: inst = 32'h8c50000;
      77024: inst = 32'h24612800;
      77025: inst = 32'h10a0ffff;
      77026: inst = 32'hca0ffff;
      77027: inst = 32'h24822800;
      77028: inst = 32'h10a00000;
      77029: inst = 32'hca00004;
      77030: inst = 32'h38632800;
      77031: inst = 32'h38842800;
      77032: inst = 32'h10a00001;
      77033: inst = 32'hca02ced;
      77034: inst = 32'h13e00001;
      77035: inst = 32'hfe0d96a;
      77036: inst = 32'h5be00000;
      77037: inst = 32'h8c50000;
      77038: inst = 32'h24612800;
      77039: inst = 32'h10a0ffff;
      77040: inst = 32'hca0ffff;
      77041: inst = 32'h24822800;
      77042: inst = 32'h10a00000;
      77043: inst = 32'hca00004;
      77044: inst = 32'h38632800;
      77045: inst = 32'h38842800;
      77046: inst = 32'h10a00001;
      77047: inst = 32'hca02cfb;
      77048: inst = 32'h13e00001;
      77049: inst = 32'hfe0d96a;
      77050: inst = 32'h5be00000;
      77051: inst = 32'h8c50000;
      77052: inst = 32'h24612800;
      77053: inst = 32'h10a0ffff;
      77054: inst = 32'hca0ffff;
      77055: inst = 32'h24822800;
      77056: inst = 32'h10a00000;
      77057: inst = 32'hca00004;
      77058: inst = 32'h38632800;
      77059: inst = 32'h38842800;
      77060: inst = 32'h10a00001;
      77061: inst = 32'hca02d09;
      77062: inst = 32'h13e00001;
      77063: inst = 32'hfe0d96a;
      77064: inst = 32'h5be00000;
      77065: inst = 32'h8c50000;
      77066: inst = 32'h24612800;
      77067: inst = 32'h10a0ffff;
      77068: inst = 32'hca0ffff;
      77069: inst = 32'h24822800;
      77070: inst = 32'h10a00000;
      77071: inst = 32'hca00004;
      77072: inst = 32'h38632800;
      77073: inst = 32'h38842800;
      77074: inst = 32'h10a00001;
      77075: inst = 32'hca02d17;
      77076: inst = 32'h13e00001;
      77077: inst = 32'hfe0d96a;
      77078: inst = 32'h5be00000;
      77079: inst = 32'h8c50000;
      77080: inst = 32'h24612800;
      77081: inst = 32'h10a0ffff;
      77082: inst = 32'hca0ffff;
      77083: inst = 32'h24822800;
      77084: inst = 32'h10a00000;
      77085: inst = 32'hca00004;
      77086: inst = 32'h38632800;
      77087: inst = 32'h38842800;
      77088: inst = 32'h10a00001;
      77089: inst = 32'hca02d25;
      77090: inst = 32'h13e00001;
      77091: inst = 32'hfe0d96a;
      77092: inst = 32'h5be00000;
      77093: inst = 32'h8c50000;
      77094: inst = 32'h24612800;
      77095: inst = 32'h10a0ffff;
      77096: inst = 32'hca0ffff;
      77097: inst = 32'h24822800;
      77098: inst = 32'h10a00000;
      77099: inst = 32'hca00004;
      77100: inst = 32'h38632800;
      77101: inst = 32'h38842800;
      77102: inst = 32'h10a00001;
      77103: inst = 32'hca02d33;
      77104: inst = 32'h13e00001;
      77105: inst = 32'hfe0d96a;
      77106: inst = 32'h5be00000;
      77107: inst = 32'h8c50000;
      77108: inst = 32'h24612800;
      77109: inst = 32'h10a0ffff;
      77110: inst = 32'hca0ffff;
      77111: inst = 32'h24822800;
      77112: inst = 32'h10a00000;
      77113: inst = 32'hca00004;
      77114: inst = 32'h38632800;
      77115: inst = 32'h38842800;
      77116: inst = 32'h10a00001;
      77117: inst = 32'hca02d41;
      77118: inst = 32'h13e00001;
      77119: inst = 32'hfe0d96a;
      77120: inst = 32'h5be00000;
      77121: inst = 32'h8c50000;
      77122: inst = 32'h24612800;
      77123: inst = 32'h10a0ffff;
      77124: inst = 32'hca0ffff;
      77125: inst = 32'h24822800;
      77126: inst = 32'h10a00000;
      77127: inst = 32'hca00004;
      77128: inst = 32'h38632800;
      77129: inst = 32'h38842800;
      77130: inst = 32'h10a00001;
      77131: inst = 32'hca02d4f;
      77132: inst = 32'h13e00001;
      77133: inst = 32'hfe0d96a;
      77134: inst = 32'h5be00000;
      77135: inst = 32'h8c50000;
      77136: inst = 32'h24612800;
      77137: inst = 32'h10a0ffff;
      77138: inst = 32'hca0ffff;
      77139: inst = 32'h24822800;
      77140: inst = 32'h10a00000;
      77141: inst = 32'hca00004;
      77142: inst = 32'h38632800;
      77143: inst = 32'h38842800;
      77144: inst = 32'h10a00001;
      77145: inst = 32'hca02d5d;
      77146: inst = 32'h13e00001;
      77147: inst = 32'hfe0d96a;
      77148: inst = 32'h5be00000;
      77149: inst = 32'h8c50000;
      77150: inst = 32'h24612800;
      77151: inst = 32'h10a0ffff;
      77152: inst = 32'hca0ffff;
      77153: inst = 32'h24822800;
      77154: inst = 32'h10a00000;
      77155: inst = 32'hca00004;
      77156: inst = 32'h38632800;
      77157: inst = 32'h38842800;
      77158: inst = 32'h10a00001;
      77159: inst = 32'hca02d6b;
      77160: inst = 32'h13e00001;
      77161: inst = 32'hfe0d96a;
      77162: inst = 32'h5be00000;
      77163: inst = 32'h8c50000;
      77164: inst = 32'h24612800;
      77165: inst = 32'h10a0ffff;
      77166: inst = 32'hca0ffff;
      77167: inst = 32'h24822800;
      77168: inst = 32'h10a00000;
      77169: inst = 32'hca00004;
      77170: inst = 32'h38632800;
      77171: inst = 32'h38842800;
      77172: inst = 32'h10a00001;
      77173: inst = 32'hca02d79;
      77174: inst = 32'h13e00001;
      77175: inst = 32'hfe0d96a;
      77176: inst = 32'h5be00000;
      77177: inst = 32'h8c50000;
      77178: inst = 32'h24612800;
      77179: inst = 32'h10a0ffff;
      77180: inst = 32'hca0ffff;
      77181: inst = 32'h24822800;
      77182: inst = 32'h10a00000;
      77183: inst = 32'hca00004;
      77184: inst = 32'h38632800;
      77185: inst = 32'h38842800;
      77186: inst = 32'h10a00001;
      77187: inst = 32'hca02d87;
      77188: inst = 32'h13e00001;
      77189: inst = 32'hfe0d96a;
      77190: inst = 32'h5be00000;
      77191: inst = 32'h8c50000;
      77192: inst = 32'h24612800;
      77193: inst = 32'h10a0ffff;
      77194: inst = 32'hca0ffff;
      77195: inst = 32'h24822800;
      77196: inst = 32'h10a00000;
      77197: inst = 32'hca00004;
      77198: inst = 32'h38632800;
      77199: inst = 32'h38842800;
      77200: inst = 32'h10a00001;
      77201: inst = 32'hca02d95;
      77202: inst = 32'h13e00001;
      77203: inst = 32'hfe0d96a;
      77204: inst = 32'h5be00000;
      77205: inst = 32'h8c50000;
      77206: inst = 32'h24612800;
      77207: inst = 32'h10a0ffff;
      77208: inst = 32'hca0ffff;
      77209: inst = 32'h24822800;
      77210: inst = 32'h10a00000;
      77211: inst = 32'hca00004;
      77212: inst = 32'h38632800;
      77213: inst = 32'h38842800;
      77214: inst = 32'h10a00001;
      77215: inst = 32'hca02da3;
      77216: inst = 32'h13e00001;
      77217: inst = 32'hfe0d96a;
      77218: inst = 32'h5be00000;
      77219: inst = 32'h8c50000;
      77220: inst = 32'h24612800;
      77221: inst = 32'h10a0ffff;
      77222: inst = 32'hca0ffff;
      77223: inst = 32'h24822800;
      77224: inst = 32'h10a00000;
      77225: inst = 32'hca00004;
      77226: inst = 32'h38632800;
      77227: inst = 32'h38842800;
      77228: inst = 32'h10a00001;
      77229: inst = 32'hca02db1;
      77230: inst = 32'h13e00001;
      77231: inst = 32'hfe0d96a;
      77232: inst = 32'h5be00000;
      77233: inst = 32'h8c50000;
      77234: inst = 32'h24612800;
      77235: inst = 32'h10a0ffff;
      77236: inst = 32'hca0ffff;
      77237: inst = 32'h24822800;
      77238: inst = 32'h10a00000;
      77239: inst = 32'hca00004;
      77240: inst = 32'h38632800;
      77241: inst = 32'h38842800;
      77242: inst = 32'h10a00001;
      77243: inst = 32'hca02dbf;
      77244: inst = 32'h13e00001;
      77245: inst = 32'hfe0d96a;
      77246: inst = 32'h5be00000;
      77247: inst = 32'h8c50000;
      77248: inst = 32'h24612800;
      77249: inst = 32'h10a0ffff;
      77250: inst = 32'hca0ffff;
      77251: inst = 32'h24822800;
      77252: inst = 32'h10a00000;
      77253: inst = 32'hca00004;
      77254: inst = 32'h38632800;
      77255: inst = 32'h38842800;
      77256: inst = 32'h10a00001;
      77257: inst = 32'hca02dcd;
      77258: inst = 32'h13e00001;
      77259: inst = 32'hfe0d96a;
      77260: inst = 32'h5be00000;
      77261: inst = 32'h8c50000;
      77262: inst = 32'h24612800;
      77263: inst = 32'h10a0ffff;
      77264: inst = 32'hca0ffff;
      77265: inst = 32'h24822800;
      77266: inst = 32'h10a00000;
      77267: inst = 32'hca00004;
      77268: inst = 32'h38632800;
      77269: inst = 32'h38842800;
      77270: inst = 32'h10a00001;
      77271: inst = 32'hca02ddb;
      77272: inst = 32'h13e00001;
      77273: inst = 32'hfe0d96a;
      77274: inst = 32'h5be00000;
      77275: inst = 32'h8c50000;
      77276: inst = 32'h24612800;
      77277: inst = 32'h10a0ffff;
      77278: inst = 32'hca0ffff;
      77279: inst = 32'h24822800;
      77280: inst = 32'h10a00000;
      77281: inst = 32'hca00004;
      77282: inst = 32'h38632800;
      77283: inst = 32'h38842800;
      77284: inst = 32'h10a00001;
      77285: inst = 32'hca02de9;
      77286: inst = 32'h13e00001;
      77287: inst = 32'hfe0d96a;
      77288: inst = 32'h5be00000;
      77289: inst = 32'h8c50000;
      77290: inst = 32'h24612800;
      77291: inst = 32'h10a0ffff;
      77292: inst = 32'hca0ffff;
      77293: inst = 32'h24822800;
      77294: inst = 32'h10a00000;
      77295: inst = 32'hca00004;
      77296: inst = 32'h38632800;
      77297: inst = 32'h38842800;
      77298: inst = 32'h10a00001;
      77299: inst = 32'hca02df7;
      77300: inst = 32'h13e00001;
      77301: inst = 32'hfe0d96a;
      77302: inst = 32'h5be00000;
      77303: inst = 32'h8c50000;
      77304: inst = 32'h24612800;
      77305: inst = 32'h10a0ffff;
      77306: inst = 32'hca0ffff;
      77307: inst = 32'h24822800;
      77308: inst = 32'h10a00000;
      77309: inst = 32'hca00004;
      77310: inst = 32'h38632800;
      77311: inst = 32'h38842800;
      77312: inst = 32'h10a00001;
      77313: inst = 32'hca02e05;
      77314: inst = 32'h13e00001;
      77315: inst = 32'hfe0d96a;
      77316: inst = 32'h5be00000;
      77317: inst = 32'h8c50000;
      77318: inst = 32'h24612800;
      77319: inst = 32'h10a0ffff;
      77320: inst = 32'hca0ffff;
      77321: inst = 32'h24822800;
      77322: inst = 32'h10a00000;
      77323: inst = 32'hca00004;
      77324: inst = 32'h38632800;
      77325: inst = 32'h38842800;
      77326: inst = 32'h10a00001;
      77327: inst = 32'hca02e13;
      77328: inst = 32'h13e00001;
      77329: inst = 32'hfe0d96a;
      77330: inst = 32'h5be00000;
      77331: inst = 32'h8c50000;
      77332: inst = 32'h24612800;
      77333: inst = 32'h10a0ffff;
      77334: inst = 32'hca0ffff;
      77335: inst = 32'h24822800;
      77336: inst = 32'h10a00000;
      77337: inst = 32'hca00004;
      77338: inst = 32'h38632800;
      77339: inst = 32'h38842800;
      77340: inst = 32'h10a00001;
      77341: inst = 32'hca02e21;
      77342: inst = 32'h13e00001;
      77343: inst = 32'hfe0d96a;
      77344: inst = 32'h5be00000;
      77345: inst = 32'h8c50000;
      77346: inst = 32'h24612800;
      77347: inst = 32'h10a0ffff;
      77348: inst = 32'hca0ffff;
      77349: inst = 32'h24822800;
      77350: inst = 32'h10a00000;
      77351: inst = 32'hca00004;
      77352: inst = 32'h38632800;
      77353: inst = 32'h38842800;
      77354: inst = 32'h10a00001;
      77355: inst = 32'hca02e2f;
      77356: inst = 32'h13e00001;
      77357: inst = 32'hfe0d96a;
      77358: inst = 32'h5be00000;
      77359: inst = 32'h8c50000;
      77360: inst = 32'h24612800;
      77361: inst = 32'h10a0ffff;
      77362: inst = 32'hca0ffff;
      77363: inst = 32'h24822800;
      77364: inst = 32'h10a00000;
      77365: inst = 32'hca00004;
      77366: inst = 32'h38632800;
      77367: inst = 32'h38842800;
      77368: inst = 32'h10a00001;
      77369: inst = 32'hca02e3d;
      77370: inst = 32'h13e00001;
      77371: inst = 32'hfe0d96a;
      77372: inst = 32'h5be00000;
      77373: inst = 32'h8c50000;
      77374: inst = 32'h24612800;
      77375: inst = 32'h10a0ffff;
      77376: inst = 32'hca0ffff;
      77377: inst = 32'h24822800;
      77378: inst = 32'h10a00000;
      77379: inst = 32'hca00004;
      77380: inst = 32'h38632800;
      77381: inst = 32'h38842800;
      77382: inst = 32'h10a00001;
      77383: inst = 32'hca02e4b;
      77384: inst = 32'h13e00001;
      77385: inst = 32'hfe0d96a;
      77386: inst = 32'h5be00000;
      77387: inst = 32'h8c50000;
      77388: inst = 32'h24612800;
      77389: inst = 32'h10a0ffff;
      77390: inst = 32'hca0ffff;
      77391: inst = 32'h24822800;
      77392: inst = 32'h10a00000;
      77393: inst = 32'hca00004;
      77394: inst = 32'h38632800;
      77395: inst = 32'h38842800;
      77396: inst = 32'h10a00001;
      77397: inst = 32'hca02e59;
      77398: inst = 32'h13e00001;
      77399: inst = 32'hfe0d96a;
      77400: inst = 32'h5be00000;
      77401: inst = 32'h8c50000;
      77402: inst = 32'h24612800;
      77403: inst = 32'h10a0ffff;
      77404: inst = 32'hca0ffff;
      77405: inst = 32'h24822800;
      77406: inst = 32'h10a00000;
      77407: inst = 32'hca00004;
      77408: inst = 32'h38632800;
      77409: inst = 32'h38842800;
      77410: inst = 32'h10a00001;
      77411: inst = 32'hca02e67;
      77412: inst = 32'h13e00001;
      77413: inst = 32'hfe0d96a;
      77414: inst = 32'h5be00000;
      77415: inst = 32'h8c50000;
      77416: inst = 32'h24612800;
      77417: inst = 32'h10a0ffff;
      77418: inst = 32'hca0ffff;
      77419: inst = 32'h24822800;
      77420: inst = 32'h10a00000;
      77421: inst = 32'hca00004;
      77422: inst = 32'h38632800;
      77423: inst = 32'h38842800;
      77424: inst = 32'h10a00001;
      77425: inst = 32'hca02e75;
      77426: inst = 32'h13e00001;
      77427: inst = 32'hfe0d96a;
      77428: inst = 32'h5be00000;
      77429: inst = 32'h8c50000;
      77430: inst = 32'h24612800;
      77431: inst = 32'h10a0ffff;
      77432: inst = 32'hca0ffff;
      77433: inst = 32'h24822800;
      77434: inst = 32'h10a00000;
      77435: inst = 32'hca00004;
      77436: inst = 32'h38632800;
      77437: inst = 32'h38842800;
      77438: inst = 32'h10a00001;
      77439: inst = 32'hca02e83;
      77440: inst = 32'h13e00001;
      77441: inst = 32'hfe0d96a;
      77442: inst = 32'h5be00000;
      77443: inst = 32'h8c50000;
      77444: inst = 32'h24612800;
      77445: inst = 32'h10a0ffff;
      77446: inst = 32'hca0ffff;
      77447: inst = 32'h24822800;
      77448: inst = 32'h10a00000;
      77449: inst = 32'hca00004;
      77450: inst = 32'h38632800;
      77451: inst = 32'h38842800;
      77452: inst = 32'h10a00001;
      77453: inst = 32'hca02e91;
      77454: inst = 32'h13e00001;
      77455: inst = 32'hfe0d96a;
      77456: inst = 32'h5be00000;
      77457: inst = 32'h8c50000;
      77458: inst = 32'h24612800;
      77459: inst = 32'h10a0ffff;
      77460: inst = 32'hca0ffff;
      77461: inst = 32'h24822800;
      77462: inst = 32'h10a00000;
      77463: inst = 32'hca00004;
      77464: inst = 32'h38632800;
      77465: inst = 32'h38842800;
      77466: inst = 32'h10a00001;
      77467: inst = 32'hca02e9f;
      77468: inst = 32'h13e00001;
      77469: inst = 32'hfe0d96a;
      77470: inst = 32'h5be00000;
      77471: inst = 32'h8c50000;
      77472: inst = 32'h24612800;
      77473: inst = 32'h10a0ffff;
      77474: inst = 32'hca0ffff;
      77475: inst = 32'h24822800;
      77476: inst = 32'h10a00000;
      77477: inst = 32'hca00004;
      77478: inst = 32'h38632800;
      77479: inst = 32'h38842800;
      77480: inst = 32'h10a00001;
      77481: inst = 32'hca02ead;
      77482: inst = 32'h13e00001;
      77483: inst = 32'hfe0d96a;
      77484: inst = 32'h5be00000;
      77485: inst = 32'h8c50000;
      77486: inst = 32'h24612800;
      77487: inst = 32'h10a0ffff;
      77488: inst = 32'hca0ffff;
      77489: inst = 32'h24822800;
      77490: inst = 32'h10a00000;
      77491: inst = 32'hca00004;
      77492: inst = 32'h38632800;
      77493: inst = 32'h38842800;
      77494: inst = 32'h10a00001;
      77495: inst = 32'hca02ebb;
      77496: inst = 32'h13e00001;
      77497: inst = 32'hfe0d96a;
      77498: inst = 32'h5be00000;
      77499: inst = 32'h8c50000;
      77500: inst = 32'h24612800;
      77501: inst = 32'h10a0ffff;
      77502: inst = 32'hca0ffff;
      77503: inst = 32'h24822800;
      77504: inst = 32'h10a00000;
      77505: inst = 32'hca00004;
      77506: inst = 32'h38632800;
      77507: inst = 32'h38842800;
      77508: inst = 32'h10a00001;
      77509: inst = 32'hca02ec9;
      77510: inst = 32'h13e00001;
      77511: inst = 32'hfe0d96a;
      77512: inst = 32'h5be00000;
      77513: inst = 32'h8c50000;
      77514: inst = 32'h24612800;
      77515: inst = 32'h10a0ffff;
      77516: inst = 32'hca0ffff;
      77517: inst = 32'h24822800;
      77518: inst = 32'h10a00000;
      77519: inst = 32'hca00004;
      77520: inst = 32'h38632800;
      77521: inst = 32'h38842800;
      77522: inst = 32'h10a00001;
      77523: inst = 32'hca02ed7;
      77524: inst = 32'h13e00001;
      77525: inst = 32'hfe0d96a;
      77526: inst = 32'h5be00000;
      77527: inst = 32'h8c50000;
      77528: inst = 32'h24612800;
      77529: inst = 32'h10a0ffff;
      77530: inst = 32'hca0ffff;
      77531: inst = 32'h24822800;
      77532: inst = 32'h10a00000;
      77533: inst = 32'hca00004;
      77534: inst = 32'h38632800;
      77535: inst = 32'h38842800;
      77536: inst = 32'h10a00001;
      77537: inst = 32'hca02ee5;
      77538: inst = 32'h13e00001;
      77539: inst = 32'hfe0d96a;
      77540: inst = 32'h5be00000;
      77541: inst = 32'h8c50000;
      77542: inst = 32'h24612800;
      77543: inst = 32'h10a0ffff;
      77544: inst = 32'hca0ffff;
      77545: inst = 32'h24822800;
      77546: inst = 32'h10a00000;
      77547: inst = 32'hca00004;
      77548: inst = 32'h38632800;
      77549: inst = 32'h38842800;
      77550: inst = 32'h10a00001;
      77551: inst = 32'hca02ef3;
      77552: inst = 32'h13e00001;
      77553: inst = 32'hfe0d96a;
      77554: inst = 32'h5be00000;
      77555: inst = 32'h8c50000;
      77556: inst = 32'h24612800;
      77557: inst = 32'h10a0ffff;
      77558: inst = 32'hca0ffff;
      77559: inst = 32'h24822800;
      77560: inst = 32'h10a00000;
      77561: inst = 32'hca00004;
      77562: inst = 32'h38632800;
      77563: inst = 32'h38842800;
      77564: inst = 32'h10a00001;
      77565: inst = 32'hca02f01;
      77566: inst = 32'h13e00001;
      77567: inst = 32'hfe0d96a;
      77568: inst = 32'h5be00000;
      77569: inst = 32'h8c50000;
      77570: inst = 32'h24612800;
      77571: inst = 32'h10a0ffff;
      77572: inst = 32'hca0ffff;
      77573: inst = 32'h24822800;
      77574: inst = 32'h10a00000;
      77575: inst = 32'hca00004;
      77576: inst = 32'h38632800;
      77577: inst = 32'h38842800;
      77578: inst = 32'h10a00001;
      77579: inst = 32'hca02f0f;
      77580: inst = 32'h13e00001;
      77581: inst = 32'hfe0d96a;
      77582: inst = 32'h5be00000;
      77583: inst = 32'h8c50000;
      77584: inst = 32'h24612800;
      77585: inst = 32'h10a0ffff;
      77586: inst = 32'hca0ffff;
      77587: inst = 32'h24822800;
      77588: inst = 32'h10a00000;
      77589: inst = 32'hca00004;
      77590: inst = 32'h38632800;
      77591: inst = 32'h38842800;
      77592: inst = 32'h10a00001;
      77593: inst = 32'hca02f1d;
      77594: inst = 32'h13e00001;
      77595: inst = 32'hfe0d96a;
      77596: inst = 32'h5be00000;
      77597: inst = 32'h8c50000;
      77598: inst = 32'h24612800;
      77599: inst = 32'h10a0ffff;
      77600: inst = 32'hca0ffff;
      77601: inst = 32'h24822800;
      77602: inst = 32'h10a00000;
      77603: inst = 32'hca00004;
      77604: inst = 32'h38632800;
      77605: inst = 32'h38842800;
      77606: inst = 32'h10a00001;
      77607: inst = 32'hca02f2b;
      77608: inst = 32'h13e00001;
      77609: inst = 32'hfe0d96a;
      77610: inst = 32'h5be00000;
      77611: inst = 32'h8c50000;
      77612: inst = 32'h24612800;
      77613: inst = 32'h10a0ffff;
      77614: inst = 32'hca0ffff;
      77615: inst = 32'h24822800;
      77616: inst = 32'h10a00000;
      77617: inst = 32'hca00004;
      77618: inst = 32'h38632800;
      77619: inst = 32'h38842800;
      77620: inst = 32'h10a00001;
      77621: inst = 32'hca02f39;
      77622: inst = 32'h13e00001;
      77623: inst = 32'hfe0d96a;
      77624: inst = 32'h5be00000;
      77625: inst = 32'h8c50000;
      77626: inst = 32'h24612800;
      77627: inst = 32'h10a0ffff;
      77628: inst = 32'hca0ffff;
      77629: inst = 32'h24822800;
      77630: inst = 32'h10a00000;
      77631: inst = 32'hca00004;
      77632: inst = 32'h38632800;
      77633: inst = 32'h38842800;
      77634: inst = 32'h10a00001;
      77635: inst = 32'hca02f47;
      77636: inst = 32'h13e00001;
      77637: inst = 32'hfe0d96a;
      77638: inst = 32'h5be00000;
      77639: inst = 32'h8c50000;
      77640: inst = 32'h24612800;
      77641: inst = 32'h10a0ffff;
      77642: inst = 32'hca0ffff;
      77643: inst = 32'h24822800;
      77644: inst = 32'h10a00000;
      77645: inst = 32'hca00004;
      77646: inst = 32'h38632800;
      77647: inst = 32'h38842800;
      77648: inst = 32'h10a00001;
      77649: inst = 32'hca02f55;
      77650: inst = 32'h13e00001;
      77651: inst = 32'hfe0d96a;
      77652: inst = 32'h5be00000;
      77653: inst = 32'h8c50000;
      77654: inst = 32'h24612800;
      77655: inst = 32'h10a0ffff;
      77656: inst = 32'hca0ffff;
      77657: inst = 32'h24822800;
      77658: inst = 32'h10a00000;
      77659: inst = 32'hca00004;
      77660: inst = 32'h38632800;
      77661: inst = 32'h38842800;
      77662: inst = 32'h10a00001;
      77663: inst = 32'hca02f63;
      77664: inst = 32'h13e00001;
      77665: inst = 32'hfe0d96a;
      77666: inst = 32'h5be00000;
      77667: inst = 32'h8c50000;
      77668: inst = 32'h24612800;
      77669: inst = 32'h10a0ffff;
      77670: inst = 32'hca0ffff;
      77671: inst = 32'h24822800;
      77672: inst = 32'h10a00000;
      77673: inst = 32'hca00004;
      77674: inst = 32'h38632800;
      77675: inst = 32'h38842800;
      77676: inst = 32'h10a00001;
      77677: inst = 32'hca02f71;
      77678: inst = 32'h13e00001;
      77679: inst = 32'hfe0d96a;
      77680: inst = 32'h5be00000;
      77681: inst = 32'h8c50000;
      77682: inst = 32'h24612800;
      77683: inst = 32'h10a0ffff;
      77684: inst = 32'hca0ffff;
      77685: inst = 32'h24822800;
      77686: inst = 32'h10a00000;
      77687: inst = 32'hca00004;
      77688: inst = 32'h38632800;
      77689: inst = 32'h38842800;
      77690: inst = 32'h10a00001;
      77691: inst = 32'hca02f7f;
      77692: inst = 32'h13e00001;
      77693: inst = 32'hfe0d96a;
      77694: inst = 32'h5be00000;
      77695: inst = 32'h8c50000;
      77696: inst = 32'h24612800;
      77697: inst = 32'h10a0ffff;
      77698: inst = 32'hca0ffff;
      77699: inst = 32'h24822800;
      77700: inst = 32'h10a00000;
      77701: inst = 32'hca00004;
      77702: inst = 32'h38632800;
      77703: inst = 32'h38842800;
      77704: inst = 32'h10a00001;
      77705: inst = 32'hca02f8d;
      77706: inst = 32'h13e00001;
      77707: inst = 32'hfe0d96a;
      77708: inst = 32'h5be00000;
      77709: inst = 32'h8c50000;
      77710: inst = 32'h24612800;
      77711: inst = 32'h10a0ffff;
      77712: inst = 32'hca0ffff;
      77713: inst = 32'h24822800;
      77714: inst = 32'h10a00000;
      77715: inst = 32'hca00004;
      77716: inst = 32'h38632800;
      77717: inst = 32'h38842800;
      77718: inst = 32'h10a00001;
      77719: inst = 32'hca02f9b;
      77720: inst = 32'h13e00001;
      77721: inst = 32'hfe0d96a;
      77722: inst = 32'h5be00000;
      77723: inst = 32'h8c50000;
      77724: inst = 32'h24612800;
      77725: inst = 32'h10a0ffff;
      77726: inst = 32'hca0ffff;
      77727: inst = 32'h24822800;
      77728: inst = 32'h10a00000;
      77729: inst = 32'hca00004;
      77730: inst = 32'h38632800;
      77731: inst = 32'h38842800;
      77732: inst = 32'h10a00001;
      77733: inst = 32'hca02fa9;
      77734: inst = 32'h13e00001;
      77735: inst = 32'hfe0d96a;
      77736: inst = 32'h5be00000;
      77737: inst = 32'h8c50000;
      77738: inst = 32'h24612800;
      77739: inst = 32'h10a0ffff;
      77740: inst = 32'hca0ffff;
      77741: inst = 32'h24822800;
      77742: inst = 32'h10a00000;
      77743: inst = 32'hca00004;
      77744: inst = 32'h38632800;
      77745: inst = 32'h38842800;
      77746: inst = 32'h10a00001;
      77747: inst = 32'hca02fb7;
      77748: inst = 32'h13e00001;
      77749: inst = 32'hfe0d96a;
      77750: inst = 32'h5be00000;
      77751: inst = 32'h8c50000;
      77752: inst = 32'h24612800;
      77753: inst = 32'h10a0ffff;
      77754: inst = 32'hca0ffff;
      77755: inst = 32'h24822800;
      77756: inst = 32'h10a00000;
      77757: inst = 32'hca00004;
      77758: inst = 32'h38632800;
      77759: inst = 32'h38842800;
      77760: inst = 32'h10a00001;
      77761: inst = 32'hca02fc5;
      77762: inst = 32'h13e00001;
      77763: inst = 32'hfe0d96a;
      77764: inst = 32'h5be00000;
      77765: inst = 32'h8c50000;
      77766: inst = 32'h24612800;
      77767: inst = 32'h10a0ffff;
      77768: inst = 32'hca0ffff;
      77769: inst = 32'h24822800;
      77770: inst = 32'h10a00000;
      77771: inst = 32'hca00004;
      77772: inst = 32'h38632800;
      77773: inst = 32'h38842800;
      77774: inst = 32'h10a00001;
      77775: inst = 32'hca02fd3;
      77776: inst = 32'h13e00001;
      77777: inst = 32'hfe0d96a;
      77778: inst = 32'h5be00000;
      77779: inst = 32'h8c50000;
      77780: inst = 32'h24612800;
      77781: inst = 32'h10a0ffff;
      77782: inst = 32'hca0ffff;
      77783: inst = 32'h24822800;
      77784: inst = 32'h10a00000;
      77785: inst = 32'hca00004;
      77786: inst = 32'h38632800;
      77787: inst = 32'h38842800;
      77788: inst = 32'h10a00001;
      77789: inst = 32'hca02fe1;
      77790: inst = 32'h13e00001;
      77791: inst = 32'hfe0d96a;
      77792: inst = 32'h5be00000;
      77793: inst = 32'h8c50000;
      77794: inst = 32'h24612800;
      77795: inst = 32'h10a0ffff;
      77796: inst = 32'hca0ffff;
      77797: inst = 32'h24822800;
      77798: inst = 32'h10a00000;
      77799: inst = 32'hca00004;
      77800: inst = 32'h38632800;
      77801: inst = 32'h38842800;
      77802: inst = 32'h10a00001;
      77803: inst = 32'hca02fef;
      77804: inst = 32'h13e00001;
      77805: inst = 32'hfe0d96a;
      77806: inst = 32'h5be00000;
      77807: inst = 32'h8c50000;
      77808: inst = 32'h24612800;
      77809: inst = 32'h10a0ffff;
      77810: inst = 32'hca0ffff;
      77811: inst = 32'h24822800;
      77812: inst = 32'h10a00000;
      77813: inst = 32'hca00004;
      77814: inst = 32'h38632800;
      77815: inst = 32'h38842800;
      77816: inst = 32'h10a00001;
      77817: inst = 32'hca02ffd;
      77818: inst = 32'h13e00001;
      77819: inst = 32'hfe0d96a;
      77820: inst = 32'h5be00000;
      77821: inst = 32'h8c50000;
      77822: inst = 32'h24612800;
      77823: inst = 32'h10a0ffff;
      77824: inst = 32'hca0ffff;
      77825: inst = 32'h24822800;
      77826: inst = 32'h10a00000;
      77827: inst = 32'hca00004;
      77828: inst = 32'h38632800;
      77829: inst = 32'h38842800;
      77830: inst = 32'h10a00001;
      77831: inst = 32'hca0300b;
      77832: inst = 32'h13e00001;
      77833: inst = 32'hfe0d96a;
      77834: inst = 32'h5be00000;
      77835: inst = 32'h8c50000;
      77836: inst = 32'h24612800;
      77837: inst = 32'h10a0ffff;
      77838: inst = 32'hca0ffff;
      77839: inst = 32'h24822800;
      77840: inst = 32'h10a00000;
      77841: inst = 32'hca00004;
      77842: inst = 32'h38632800;
      77843: inst = 32'h38842800;
      77844: inst = 32'h10a00001;
      77845: inst = 32'hca03019;
      77846: inst = 32'h13e00001;
      77847: inst = 32'hfe0d96a;
      77848: inst = 32'h5be00000;
      77849: inst = 32'h8c50000;
      77850: inst = 32'h24612800;
      77851: inst = 32'h10a0ffff;
      77852: inst = 32'hca0ffff;
      77853: inst = 32'h24822800;
      77854: inst = 32'h10a00000;
      77855: inst = 32'hca00004;
      77856: inst = 32'h38632800;
      77857: inst = 32'h38842800;
      77858: inst = 32'h10a00001;
      77859: inst = 32'hca03027;
      77860: inst = 32'h13e00001;
      77861: inst = 32'hfe0d96a;
      77862: inst = 32'h5be00000;
      77863: inst = 32'h8c50000;
      77864: inst = 32'h24612800;
      77865: inst = 32'h10a0ffff;
      77866: inst = 32'hca0ffff;
      77867: inst = 32'h24822800;
      77868: inst = 32'h10a00000;
      77869: inst = 32'hca00004;
      77870: inst = 32'h38632800;
      77871: inst = 32'h38842800;
      77872: inst = 32'h10a00001;
      77873: inst = 32'hca03035;
      77874: inst = 32'h13e00001;
      77875: inst = 32'hfe0d96a;
      77876: inst = 32'h5be00000;
      77877: inst = 32'h8c50000;
      77878: inst = 32'h24612800;
      77879: inst = 32'h10a0ffff;
      77880: inst = 32'hca0ffff;
      77881: inst = 32'h24822800;
      77882: inst = 32'h10a00000;
      77883: inst = 32'hca00004;
      77884: inst = 32'h38632800;
      77885: inst = 32'h38842800;
      77886: inst = 32'h10a00001;
      77887: inst = 32'hca03043;
      77888: inst = 32'h13e00001;
      77889: inst = 32'hfe0d96a;
      77890: inst = 32'h5be00000;
      77891: inst = 32'h8c50000;
      77892: inst = 32'h24612800;
      77893: inst = 32'h10a0ffff;
      77894: inst = 32'hca0ffff;
      77895: inst = 32'h24822800;
      77896: inst = 32'h10a00000;
      77897: inst = 32'hca00004;
      77898: inst = 32'h38632800;
      77899: inst = 32'h38842800;
      77900: inst = 32'h10a00001;
      77901: inst = 32'hca03051;
      77902: inst = 32'h13e00001;
      77903: inst = 32'hfe0d96a;
      77904: inst = 32'h5be00000;
      77905: inst = 32'h8c50000;
      77906: inst = 32'h24612800;
      77907: inst = 32'h10a0ffff;
      77908: inst = 32'hca0ffff;
      77909: inst = 32'h24822800;
      77910: inst = 32'h10a00000;
      77911: inst = 32'hca00004;
      77912: inst = 32'h38632800;
      77913: inst = 32'h38842800;
      77914: inst = 32'h10a00001;
      77915: inst = 32'hca0305f;
      77916: inst = 32'h13e00001;
      77917: inst = 32'hfe0d96a;
      77918: inst = 32'h5be00000;
      77919: inst = 32'h8c50000;
      77920: inst = 32'h24612800;
      77921: inst = 32'h10a0ffff;
      77922: inst = 32'hca0ffff;
      77923: inst = 32'h24822800;
      77924: inst = 32'h10a00000;
      77925: inst = 32'hca00004;
      77926: inst = 32'h38632800;
      77927: inst = 32'h38842800;
      77928: inst = 32'h10a00001;
      77929: inst = 32'hca0306d;
      77930: inst = 32'h13e00001;
      77931: inst = 32'hfe0d96a;
      77932: inst = 32'h5be00000;
      77933: inst = 32'h8c50000;
      77934: inst = 32'h24612800;
      77935: inst = 32'h10a0ffff;
      77936: inst = 32'hca0ffff;
      77937: inst = 32'h24822800;
      77938: inst = 32'h10a00000;
      77939: inst = 32'hca00004;
      77940: inst = 32'h38632800;
      77941: inst = 32'h38842800;
      77942: inst = 32'h10a00001;
      77943: inst = 32'hca0307b;
      77944: inst = 32'h13e00001;
      77945: inst = 32'hfe0d96a;
      77946: inst = 32'h5be00000;
      77947: inst = 32'h8c50000;
      77948: inst = 32'h24612800;
      77949: inst = 32'h10a0ffff;
      77950: inst = 32'hca0ffff;
      77951: inst = 32'h24822800;
      77952: inst = 32'h10a00000;
      77953: inst = 32'hca00004;
      77954: inst = 32'h38632800;
      77955: inst = 32'h38842800;
      77956: inst = 32'h10a00001;
      77957: inst = 32'hca03089;
      77958: inst = 32'h13e00001;
      77959: inst = 32'hfe0d96a;
      77960: inst = 32'h5be00000;
      77961: inst = 32'h8c50000;
      77962: inst = 32'h24612800;
      77963: inst = 32'h10a0ffff;
      77964: inst = 32'hca0ffff;
      77965: inst = 32'h24822800;
      77966: inst = 32'h10a00000;
      77967: inst = 32'hca00004;
      77968: inst = 32'h38632800;
      77969: inst = 32'h38842800;
      77970: inst = 32'h10a00001;
      77971: inst = 32'hca03097;
      77972: inst = 32'h13e00001;
      77973: inst = 32'hfe0d96a;
      77974: inst = 32'h5be00000;
      77975: inst = 32'h8c50000;
      77976: inst = 32'h24612800;
      77977: inst = 32'h10a0ffff;
      77978: inst = 32'hca0ffff;
      77979: inst = 32'h24822800;
      77980: inst = 32'h10a00000;
      77981: inst = 32'hca00004;
      77982: inst = 32'h38632800;
      77983: inst = 32'h38842800;
      77984: inst = 32'h10a00001;
      77985: inst = 32'hca030a5;
      77986: inst = 32'h13e00001;
      77987: inst = 32'hfe0d96a;
      77988: inst = 32'h5be00000;
      77989: inst = 32'h8c50000;
      77990: inst = 32'h24612800;
      77991: inst = 32'h10a0ffff;
      77992: inst = 32'hca0ffff;
      77993: inst = 32'h24822800;
      77994: inst = 32'h10a00000;
      77995: inst = 32'hca00004;
      77996: inst = 32'h38632800;
      77997: inst = 32'h38842800;
      77998: inst = 32'h10a00001;
      77999: inst = 32'hca030b3;
      78000: inst = 32'h13e00001;
      78001: inst = 32'hfe0d96a;
      78002: inst = 32'h5be00000;
      78003: inst = 32'h8c50000;
      78004: inst = 32'h24612800;
      78005: inst = 32'h10a0ffff;
      78006: inst = 32'hca0ffff;
      78007: inst = 32'h24822800;
      78008: inst = 32'h10a00000;
      78009: inst = 32'hca00004;
      78010: inst = 32'h38632800;
      78011: inst = 32'h38842800;
      78012: inst = 32'h10a00001;
      78013: inst = 32'hca030c1;
      78014: inst = 32'h13e00001;
      78015: inst = 32'hfe0d96a;
      78016: inst = 32'h5be00000;
      78017: inst = 32'h8c50000;
      78018: inst = 32'h24612800;
      78019: inst = 32'h10a0ffff;
      78020: inst = 32'hca0ffff;
      78021: inst = 32'h24822800;
      78022: inst = 32'h10a00000;
      78023: inst = 32'hca00004;
      78024: inst = 32'h38632800;
      78025: inst = 32'h38842800;
      78026: inst = 32'h10a00001;
      78027: inst = 32'hca030cf;
      78028: inst = 32'h13e00001;
      78029: inst = 32'hfe0d96a;
      78030: inst = 32'h5be00000;
      78031: inst = 32'h8c50000;
      78032: inst = 32'h24612800;
      78033: inst = 32'h10a0ffff;
      78034: inst = 32'hca0ffff;
      78035: inst = 32'h24822800;
      78036: inst = 32'h10a00000;
      78037: inst = 32'hca00004;
      78038: inst = 32'h38632800;
      78039: inst = 32'h38842800;
      78040: inst = 32'h10a00001;
      78041: inst = 32'hca030dd;
      78042: inst = 32'h13e00001;
      78043: inst = 32'hfe0d96a;
      78044: inst = 32'h5be00000;
      78045: inst = 32'h8c50000;
      78046: inst = 32'h24612800;
      78047: inst = 32'h10a0ffff;
      78048: inst = 32'hca0ffff;
      78049: inst = 32'h24822800;
      78050: inst = 32'h10a00000;
      78051: inst = 32'hca00004;
      78052: inst = 32'h38632800;
      78053: inst = 32'h38842800;
      78054: inst = 32'h10a00001;
      78055: inst = 32'hca030eb;
      78056: inst = 32'h13e00001;
      78057: inst = 32'hfe0d96a;
      78058: inst = 32'h5be00000;
      78059: inst = 32'h8c50000;
      78060: inst = 32'h24612800;
      78061: inst = 32'h10a0ffff;
      78062: inst = 32'hca0ffff;
      78063: inst = 32'h24822800;
      78064: inst = 32'h10a00000;
      78065: inst = 32'hca00004;
      78066: inst = 32'h38632800;
      78067: inst = 32'h38842800;
      78068: inst = 32'h10a00001;
      78069: inst = 32'hca030f9;
      78070: inst = 32'h13e00001;
      78071: inst = 32'hfe0d96a;
      78072: inst = 32'h5be00000;
      78073: inst = 32'h8c50000;
      78074: inst = 32'h24612800;
      78075: inst = 32'h10a0ffff;
      78076: inst = 32'hca0ffff;
      78077: inst = 32'h24822800;
      78078: inst = 32'h10a00000;
      78079: inst = 32'hca00004;
      78080: inst = 32'h38632800;
      78081: inst = 32'h38842800;
      78082: inst = 32'h10a00001;
      78083: inst = 32'hca03107;
      78084: inst = 32'h13e00001;
      78085: inst = 32'hfe0d96a;
      78086: inst = 32'h5be00000;
      78087: inst = 32'h8c50000;
      78088: inst = 32'h24612800;
      78089: inst = 32'h10a0ffff;
      78090: inst = 32'hca0ffff;
      78091: inst = 32'h24822800;
      78092: inst = 32'h10a00000;
      78093: inst = 32'hca00004;
      78094: inst = 32'h38632800;
      78095: inst = 32'h38842800;
      78096: inst = 32'h10a00001;
      78097: inst = 32'hca03115;
      78098: inst = 32'h13e00001;
      78099: inst = 32'hfe0d96a;
      78100: inst = 32'h5be00000;
      78101: inst = 32'h8c50000;
      78102: inst = 32'h24612800;
      78103: inst = 32'h10a0ffff;
      78104: inst = 32'hca0ffff;
      78105: inst = 32'h24822800;
      78106: inst = 32'h10a00000;
      78107: inst = 32'hca00004;
      78108: inst = 32'h38632800;
      78109: inst = 32'h38842800;
      78110: inst = 32'h10a00001;
      78111: inst = 32'hca03123;
      78112: inst = 32'h13e00001;
      78113: inst = 32'hfe0d96a;
      78114: inst = 32'h5be00000;
      78115: inst = 32'h8c50000;
      78116: inst = 32'h24612800;
      78117: inst = 32'h10a0ffff;
      78118: inst = 32'hca0ffff;
      78119: inst = 32'h24822800;
      78120: inst = 32'h10a00000;
      78121: inst = 32'hca00004;
      78122: inst = 32'h38632800;
      78123: inst = 32'h38842800;
      78124: inst = 32'h10a00001;
      78125: inst = 32'hca03131;
      78126: inst = 32'h13e00001;
      78127: inst = 32'hfe0d96a;
      78128: inst = 32'h5be00000;
      78129: inst = 32'h8c50000;
      78130: inst = 32'h24612800;
      78131: inst = 32'h10a0ffff;
      78132: inst = 32'hca0ffff;
      78133: inst = 32'h24822800;
      78134: inst = 32'h10a00000;
      78135: inst = 32'hca00004;
      78136: inst = 32'h38632800;
      78137: inst = 32'h38842800;
      78138: inst = 32'h10a00001;
      78139: inst = 32'hca0313f;
      78140: inst = 32'h13e00001;
      78141: inst = 32'hfe0d96a;
      78142: inst = 32'h5be00000;
      78143: inst = 32'h8c50000;
      78144: inst = 32'h24612800;
      78145: inst = 32'h10a0ffff;
      78146: inst = 32'hca0ffff;
      78147: inst = 32'h24822800;
      78148: inst = 32'h10a00000;
      78149: inst = 32'hca00004;
      78150: inst = 32'h38632800;
      78151: inst = 32'h38842800;
      78152: inst = 32'h10a00001;
      78153: inst = 32'hca0314d;
      78154: inst = 32'h13e00001;
      78155: inst = 32'hfe0d96a;
      78156: inst = 32'h5be00000;
      78157: inst = 32'h8c50000;
      78158: inst = 32'h24612800;
      78159: inst = 32'h10a0ffff;
      78160: inst = 32'hca0ffff;
      78161: inst = 32'h24822800;
      78162: inst = 32'h10a00000;
      78163: inst = 32'hca00004;
      78164: inst = 32'h38632800;
      78165: inst = 32'h38842800;
      78166: inst = 32'h10a00001;
      78167: inst = 32'hca0315b;
      78168: inst = 32'h13e00001;
      78169: inst = 32'hfe0d96a;
      78170: inst = 32'h5be00000;
      78171: inst = 32'h8c50000;
      78172: inst = 32'h24612800;
      78173: inst = 32'h10a0ffff;
      78174: inst = 32'hca0ffff;
      78175: inst = 32'h24822800;
      78176: inst = 32'h10a00000;
      78177: inst = 32'hca00004;
      78178: inst = 32'h38632800;
      78179: inst = 32'h38842800;
      78180: inst = 32'h10a00001;
      78181: inst = 32'hca03169;
      78182: inst = 32'h13e00001;
      78183: inst = 32'hfe0d96a;
      78184: inst = 32'h5be00000;
      78185: inst = 32'h8c50000;
      78186: inst = 32'h24612800;
      78187: inst = 32'h10a00000;
      78188: inst = 32'hca00000;
      78189: inst = 32'h24822800;
      78190: inst = 32'h10a00000;
      78191: inst = 32'hca00004;
      78192: inst = 32'h38632800;
      78193: inst = 32'h38842800;
      78194: inst = 32'h10a00001;
      78195: inst = 32'hca03177;
      78196: inst = 32'h13e00001;
      78197: inst = 32'hfe0d96a;
      78198: inst = 32'h5be00000;
      78199: inst = 32'h8c50000;
      78200: inst = 32'h24612800;
      78201: inst = 32'h10a00000;
      78202: inst = 32'hca00000;
      78203: inst = 32'h24822800;
      78204: inst = 32'h10a00000;
      78205: inst = 32'hca00004;
      78206: inst = 32'h38632800;
      78207: inst = 32'h38842800;
      78208: inst = 32'h10a00001;
      78209: inst = 32'hca03185;
      78210: inst = 32'h13e00001;
      78211: inst = 32'hfe0d96a;
      78212: inst = 32'h5be00000;
      78213: inst = 32'h8c50000;
      78214: inst = 32'h24612800;
      78215: inst = 32'h10a00000;
      78216: inst = 32'hca00000;
      78217: inst = 32'h24822800;
      78218: inst = 32'h10a00000;
      78219: inst = 32'hca00004;
      78220: inst = 32'h38632800;
      78221: inst = 32'h38842800;
      78222: inst = 32'h10a00001;
      78223: inst = 32'hca03193;
      78224: inst = 32'h13e00001;
      78225: inst = 32'hfe0d96a;
      78226: inst = 32'h5be00000;
      78227: inst = 32'h8c50000;
      78228: inst = 32'h24612800;
      78229: inst = 32'h10a00000;
      78230: inst = 32'hca00000;
      78231: inst = 32'h24822800;
      78232: inst = 32'h10a00000;
      78233: inst = 32'hca00004;
      78234: inst = 32'h38632800;
      78235: inst = 32'h38842800;
      78236: inst = 32'h10a00001;
      78237: inst = 32'hca031a1;
      78238: inst = 32'h13e00001;
      78239: inst = 32'hfe0d96a;
      78240: inst = 32'h5be00000;
      78241: inst = 32'h8c50000;
      78242: inst = 32'h24612800;
      78243: inst = 32'h10a00000;
      78244: inst = 32'hca00000;
      78245: inst = 32'h24822800;
      78246: inst = 32'h10a00000;
      78247: inst = 32'hca00004;
      78248: inst = 32'h38632800;
      78249: inst = 32'h38842800;
      78250: inst = 32'h10a00001;
      78251: inst = 32'hca031af;
      78252: inst = 32'h13e00001;
      78253: inst = 32'hfe0d96a;
      78254: inst = 32'h5be00000;
      78255: inst = 32'h8c50000;
      78256: inst = 32'h24612800;
      78257: inst = 32'h10a00000;
      78258: inst = 32'hca00000;
      78259: inst = 32'h24822800;
      78260: inst = 32'h10a00000;
      78261: inst = 32'hca00004;
      78262: inst = 32'h38632800;
      78263: inst = 32'h38842800;
      78264: inst = 32'h10a00001;
      78265: inst = 32'hca031bd;
      78266: inst = 32'h13e00001;
      78267: inst = 32'hfe0d96a;
      78268: inst = 32'h5be00000;
      78269: inst = 32'h8c50000;
      78270: inst = 32'h24612800;
      78271: inst = 32'h10a00000;
      78272: inst = 32'hca00000;
      78273: inst = 32'h24822800;
      78274: inst = 32'h10a00000;
      78275: inst = 32'hca00004;
      78276: inst = 32'h38632800;
      78277: inst = 32'h38842800;
      78278: inst = 32'h10a00001;
      78279: inst = 32'hca031cb;
      78280: inst = 32'h13e00001;
      78281: inst = 32'hfe0d96a;
      78282: inst = 32'h5be00000;
      78283: inst = 32'h8c50000;
      78284: inst = 32'h24612800;
      78285: inst = 32'h10a00000;
      78286: inst = 32'hca00000;
      78287: inst = 32'h24822800;
      78288: inst = 32'h10a00000;
      78289: inst = 32'hca00004;
      78290: inst = 32'h38632800;
      78291: inst = 32'h38842800;
      78292: inst = 32'h10a00001;
      78293: inst = 32'hca031d9;
      78294: inst = 32'h13e00001;
      78295: inst = 32'hfe0d96a;
      78296: inst = 32'h5be00000;
      78297: inst = 32'h8c50000;
      78298: inst = 32'h24612800;
      78299: inst = 32'h10a00000;
      78300: inst = 32'hca00000;
      78301: inst = 32'h24822800;
      78302: inst = 32'h10a00000;
      78303: inst = 32'hca00004;
      78304: inst = 32'h38632800;
      78305: inst = 32'h38842800;
      78306: inst = 32'h10a00001;
      78307: inst = 32'hca031e7;
      78308: inst = 32'h13e00001;
      78309: inst = 32'hfe0d96a;
      78310: inst = 32'h5be00000;
      78311: inst = 32'h8c50000;
      78312: inst = 32'h24612800;
      78313: inst = 32'h10a00000;
      78314: inst = 32'hca00000;
      78315: inst = 32'h24822800;
      78316: inst = 32'h10a00000;
      78317: inst = 32'hca00004;
      78318: inst = 32'h38632800;
      78319: inst = 32'h38842800;
      78320: inst = 32'h10a00001;
      78321: inst = 32'hca031f5;
      78322: inst = 32'h13e00001;
      78323: inst = 32'hfe0d96a;
      78324: inst = 32'h5be00000;
      78325: inst = 32'h8c50000;
      78326: inst = 32'h24612800;
      78327: inst = 32'h10a00000;
      78328: inst = 32'hca00000;
      78329: inst = 32'h24822800;
      78330: inst = 32'h10a00000;
      78331: inst = 32'hca00004;
      78332: inst = 32'h38632800;
      78333: inst = 32'h38842800;
      78334: inst = 32'h10a00001;
      78335: inst = 32'hca03203;
      78336: inst = 32'h13e00001;
      78337: inst = 32'hfe0d96a;
      78338: inst = 32'h5be00000;
      78339: inst = 32'h8c50000;
      78340: inst = 32'h24612800;
      78341: inst = 32'h10a00000;
      78342: inst = 32'hca00000;
      78343: inst = 32'h24822800;
      78344: inst = 32'h10a00000;
      78345: inst = 32'hca00004;
      78346: inst = 32'h38632800;
      78347: inst = 32'h38842800;
      78348: inst = 32'h10a00001;
      78349: inst = 32'hca03211;
      78350: inst = 32'h13e00001;
      78351: inst = 32'hfe0d96a;
      78352: inst = 32'h5be00000;
      78353: inst = 32'h8c50000;
      78354: inst = 32'h24612800;
      78355: inst = 32'h10a00000;
      78356: inst = 32'hca00000;
      78357: inst = 32'h24822800;
      78358: inst = 32'h10a00000;
      78359: inst = 32'hca00004;
      78360: inst = 32'h38632800;
      78361: inst = 32'h38842800;
      78362: inst = 32'h10a00001;
      78363: inst = 32'hca0321f;
      78364: inst = 32'h13e00001;
      78365: inst = 32'hfe0d96a;
      78366: inst = 32'h5be00000;
      78367: inst = 32'h8c50000;
      78368: inst = 32'h24612800;
      78369: inst = 32'h10a00000;
      78370: inst = 32'hca00000;
      78371: inst = 32'h24822800;
      78372: inst = 32'h10a00000;
      78373: inst = 32'hca00004;
      78374: inst = 32'h38632800;
      78375: inst = 32'h38842800;
      78376: inst = 32'h10a00001;
      78377: inst = 32'hca0322d;
      78378: inst = 32'h13e00001;
      78379: inst = 32'hfe0d96a;
      78380: inst = 32'h5be00000;
      78381: inst = 32'h8c50000;
      78382: inst = 32'h24612800;
      78383: inst = 32'h10a00000;
      78384: inst = 32'hca00000;
      78385: inst = 32'h24822800;
      78386: inst = 32'h10a00000;
      78387: inst = 32'hca00004;
      78388: inst = 32'h38632800;
      78389: inst = 32'h38842800;
      78390: inst = 32'h10a00001;
      78391: inst = 32'hca0323b;
      78392: inst = 32'h13e00001;
      78393: inst = 32'hfe0d96a;
      78394: inst = 32'h5be00000;
      78395: inst = 32'h8c50000;
      78396: inst = 32'h24612800;
      78397: inst = 32'h10a00000;
      78398: inst = 32'hca00000;
      78399: inst = 32'h24822800;
      78400: inst = 32'h10a00000;
      78401: inst = 32'hca00004;
      78402: inst = 32'h38632800;
      78403: inst = 32'h38842800;
      78404: inst = 32'h10a00001;
      78405: inst = 32'hca03249;
      78406: inst = 32'h13e00001;
      78407: inst = 32'hfe0d96a;
      78408: inst = 32'h5be00000;
      78409: inst = 32'h8c50000;
      78410: inst = 32'h24612800;
      78411: inst = 32'h10a00000;
      78412: inst = 32'hca00000;
      78413: inst = 32'h24822800;
      78414: inst = 32'h10a00000;
      78415: inst = 32'hca00004;
      78416: inst = 32'h38632800;
      78417: inst = 32'h38842800;
      78418: inst = 32'h10a00001;
      78419: inst = 32'hca03257;
      78420: inst = 32'h13e00001;
      78421: inst = 32'hfe0d96a;
      78422: inst = 32'h5be00000;
      78423: inst = 32'h8c50000;
      78424: inst = 32'h24612800;
      78425: inst = 32'h10a00000;
      78426: inst = 32'hca00000;
      78427: inst = 32'h24822800;
      78428: inst = 32'h10a00000;
      78429: inst = 32'hca00004;
      78430: inst = 32'h38632800;
      78431: inst = 32'h38842800;
      78432: inst = 32'h10a00001;
      78433: inst = 32'hca03265;
      78434: inst = 32'h13e00001;
      78435: inst = 32'hfe0d96a;
      78436: inst = 32'h5be00000;
      78437: inst = 32'h8c50000;
      78438: inst = 32'h24612800;
      78439: inst = 32'h10a00000;
      78440: inst = 32'hca00000;
      78441: inst = 32'h24822800;
      78442: inst = 32'h10a00000;
      78443: inst = 32'hca00004;
      78444: inst = 32'h38632800;
      78445: inst = 32'h38842800;
      78446: inst = 32'h10a00001;
      78447: inst = 32'hca03273;
      78448: inst = 32'h13e00001;
      78449: inst = 32'hfe0d96a;
      78450: inst = 32'h5be00000;
      78451: inst = 32'h8c50000;
      78452: inst = 32'h24612800;
      78453: inst = 32'h10a00000;
      78454: inst = 32'hca00000;
      78455: inst = 32'h24822800;
      78456: inst = 32'h10a00000;
      78457: inst = 32'hca00004;
      78458: inst = 32'h38632800;
      78459: inst = 32'h38842800;
      78460: inst = 32'h10a00001;
      78461: inst = 32'hca03281;
      78462: inst = 32'h13e00001;
      78463: inst = 32'hfe0d96a;
      78464: inst = 32'h5be00000;
      78465: inst = 32'h8c50000;
      78466: inst = 32'h24612800;
      78467: inst = 32'h10a00000;
      78468: inst = 32'hca00000;
      78469: inst = 32'h24822800;
      78470: inst = 32'h10a00000;
      78471: inst = 32'hca00004;
      78472: inst = 32'h38632800;
      78473: inst = 32'h38842800;
      78474: inst = 32'h10a00001;
      78475: inst = 32'hca0328f;
      78476: inst = 32'h13e00001;
      78477: inst = 32'hfe0d96a;
      78478: inst = 32'h5be00000;
      78479: inst = 32'h8c50000;
      78480: inst = 32'h24612800;
      78481: inst = 32'h10a00000;
      78482: inst = 32'hca00000;
      78483: inst = 32'h24822800;
      78484: inst = 32'h10a00000;
      78485: inst = 32'hca00004;
      78486: inst = 32'h38632800;
      78487: inst = 32'h38842800;
      78488: inst = 32'h10a00001;
      78489: inst = 32'hca0329d;
      78490: inst = 32'h13e00001;
      78491: inst = 32'hfe0d96a;
      78492: inst = 32'h5be00000;
      78493: inst = 32'h8c50000;
      78494: inst = 32'h24612800;
      78495: inst = 32'h10a00000;
      78496: inst = 32'hca00000;
      78497: inst = 32'h24822800;
      78498: inst = 32'h10a00000;
      78499: inst = 32'hca00004;
      78500: inst = 32'h38632800;
      78501: inst = 32'h38842800;
      78502: inst = 32'h10a00001;
      78503: inst = 32'hca032ab;
      78504: inst = 32'h13e00001;
      78505: inst = 32'hfe0d96a;
      78506: inst = 32'h5be00000;
      78507: inst = 32'h8c50000;
      78508: inst = 32'h24612800;
      78509: inst = 32'h10a00000;
      78510: inst = 32'hca00000;
      78511: inst = 32'h24822800;
      78512: inst = 32'h10a00000;
      78513: inst = 32'hca00004;
      78514: inst = 32'h38632800;
      78515: inst = 32'h38842800;
      78516: inst = 32'h10a00001;
      78517: inst = 32'hca032b9;
      78518: inst = 32'h13e00001;
      78519: inst = 32'hfe0d96a;
      78520: inst = 32'h5be00000;
      78521: inst = 32'h8c50000;
      78522: inst = 32'h24612800;
      78523: inst = 32'h10a00000;
      78524: inst = 32'hca00000;
      78525: inst = 32'h24822800;
      78526: inst = 32'h10a00000;
      78527: inst = 32'hca00004;
      78528: inst = 32'h38632800;
      78529: inst = 32'h38842800;
      78530: inst = 32'h10a00001;
      78531: inst = 32'hca032c7;
      78532: inst = 32'h13e00001;
      78533: inst = 32'hfe0d96a;
      78534: inst = 32'h5be00000;
      78535: inst = 32'h8c50000;
      78536: inst = 32'h24612800;
      78537: inst = 32'h10a00000;
      78538: inst = 32'hca00000;
      78539: inst = 32'h24822800;
      78540: inst = 32'h10a00000;
      78541: inst = 32'hca00004;
      78542: inst = 32'h38632800;
      78543: inst = 32'h38842800;
      78544: inst = 32'h10a00001;
      78545: inst = 32'hca032d5;
      78546: inst = 32'h13e00001;
      78547: inst = 32'hfe0d96a;
      78548: inst = 32'h5be00000;
      78549: inst = 32'h8c50000;
      78550: inst = 32'h24612800;
      78551: inst = 32'h10a00000;
      78552: inst = 32'hca00000;
      78553: inst = 32'h24822800;
      78554: inst = 32'h10a00000;
      78555: inst = 32'hca00004;
      78556: inst = 32'h38632800;
      78557: inst = 32'h38842800;
      78558: inst = 32'h10a00001;
      78559: inst = 32'hca032e3;
      78560: inst = 32'h13e00001;
      78561: inst = 32'hfe0d96a;
      78562: inst = 32'h5be00000;
      78563: inst = 32'h8c50000;
      78564: inst = 32'h24612800;
      78565: inst = 32'h10a00000;
      78566: inst = 32'hca00000;
      78567: inst = 32'h24822800;
      78568: inst = 32'h10a00000;
      78569: inst = 32'hca00004;
      78570: inst = 32'h38632800;
      78571: inst = 32'h38842800;
      78572: inst = 32'h10a00001;
      78573: inst = 32'hca032f1;
      78574: inst = 32'h13e00001;
      78575: inst = 32'hfe0d96a;
      78576: inst = 32'h5be00000;
      78577: inst = 32'h8c50000;
      78578: inst = 32'h24612800;
      78579: inst = 32'h10a00000;
      78580: inst = 32'hca00000;
      78581: inst = 32'h24822800;
      78582: inst = 32'h10a00000;
      78583: inst = 32'hca00004;
      78584: inst = 32'h38632800;
      78585: inst = 32'h38842800;
      78586: inst = 32'h10a00001;
      78587: inst = 32'hca032ff;
      78588: inst = 32'h13e00001;
      78589: inst = 32'hfe0d96a;
      78590: inst = 32'h5be00000;
      78591: inst = 32'h8c50000;
      78592: inst = 32'h24612800;
      78593: inst = 32'h10a00000;
      78594: inst = 32'hca00000;
      78595: inst = 32'h24822800;
      78596: inst = 32'h10a00000;
      78597: inst = 32'hca00004;
      78598: inst = 32'h38632800;
      78599: inst = 32'h38842800;
      78600: inst = 32'h10a00001;
      78601: inst = 32'hca0330d;
      78602: inst = 32'h13e00001;
      78603: inst = 32'hfe0d96a;
      78604: inst = 32'h5be00000;
      78605: inst = 32'h8c50000;
      78606: inst = 32'h24612800;
      78607: inst = 32'h10a00000;
      78608: inst = 32'hca00000;
      78609: inst = 32'h24822800;
      78610: inst = 32'h10a00000;
      78611: inst = 32'hca00004;
      78612: inst = 32'h38632800;
      78613: inst = 32'h38842800;
      78614: inst = 32'h10a00001;
      78615: inst = 32'hca0331b;
      78616: inst = 32'h13e00001;
      78617: inst = 32'hfe0d96a;
      78618: inst = 32'h5be00000;
      78619: inst = 32'h8c50000;
      78620: inst = 32'h24612800;
      78621: inst = 32'h10a00000;
      78622: inst = 32'hca00000;
      78623: inst = 32'h24822800;
      78624: inst = 32'h10a00000;
      78625: inst = 32'hca00004;
      78626: inst = 32'h38632800;
      78627: inst = 32'h38842800;
      78628: inst = 32'h10a00001;
      78629: inst = 32'hca03329;
      78630: inst = 32'h13e00001;
      78631: inst = 32'hfe0d96a;
      78632: inst = 32'h5be00000;
      78633: inst = 32'h8c50000;
      78634: inst = 32'h24612800;
      78635: inst = 32'h10a00000;
      78636: inst = 32'hca00000;
      78637: inst = 32'h24822800;
      78638: inst = 32'h10a00000;
      78639: inst = 32'hca00004;
      78640: inst = 32'h38632800;
      78641: inst = 32'h38842800;
      78642: inst = 32'h10a00001;
      78643: inst = 32'hca03337;
      78644: inst = 32'h13e00001;
      78645: inst = 32'hfe0d96a;
      78646: inst = 32'h5be00000;
      78647: inst = 32'h8c50000;
      78648: inst = 32'h24612800;
      78649: inst = 32'h10a00000;
      78650: inst = 32'hca00000;
      78651: inst = 32'h24822800;
      78652: inst = 32'h10a00000;
      78653: inst = 32'hca00004;
      78654: inst = 32'h38632800;
      78655: inst = 32'h38842800;
      78656: inst = 32'h10a00001;
      78657: inst = 32'hca03345;
      78658: inst = 32'h13e00001;
      78659: inst = 32'hfe0d96a;
      78660: inst = 32'h5be00000;
      78661: inst = 32'h8c50000;
      78662: inst = 32'h24612800;
      78663: inst = 32'h10a00000;
      78664: inst = 32'hca00000;
      78665: inst = 32'h24822800;
      78666: inst = 32'h10a00000;
      78667: inst = 32'hca00004;
      78668: inst = 32'h38632800;
      78669: inst = 32'h38842800;
      78670: inst = 32'h10a00001;
      78671: inst = 32'hca03353;
      78672: inst = 32'h13e00001;
      78673: inst = 32'hfe0d96a;
      78674: inst = 32'h5be00000;
      78675: inst = 32'h8c50000;
      78676: inst = 32'h24612800;
      78677: inst = 32'h10a00000;
      78678: inst = 32'hca00000;
      78679: inst = 32'h24822800;
      78680: inst = 32'h10a00000;
      78681: inst = 32'hca00004;
      78682: inst = 32'h38632800;
      78683: inst = 32'h38842800;
      78684: inst = 32'h10a00001;
      78685: inst = 32'hca03361;
      78686: inst = 32'h13e00001;
      78687: inst = 32'hfe0d96a;
      78688: inst = 32'h5be00000;
      78689: inst = 32'h8c50000;
      78690: inst = 32'h24612800;
      78691: inst = 32'h10a00000;
      78692: inst = 32'hca00000;
      78693: inst = 32'h24822800;
      78694: inst = 32'h10a00000;
      78695: inst = 32'hca00004;
      78696: inst = 32'h38632800;
      78697: inst = 32'h38842800;
      78698: inst = 32'h10a00001;
      78699: inst = 32'hca0336f;
      78700: inst = 32'h13e00001;
      78701: inst = 32'hfe0d96a;
      78702: inst = 32'h5be00000;
      78703: inst = 32'h8c50000;
      78704: inst = 32'h24612800;
      78705: inst = 32'h10a00000;
      78706: inst = 32'hca00000;
      78707: inst = 32'h24822800;
      78708: inst = 32'h10a00000;
      78709: inst = 32'hca00004;
      78710: inst = 32'h38632800;
      78711: inst = 32'h38842800;
      78712: inst = 32'h10a00001;
      78713: inst = 32'hca0337d;
      78714: inst = 32'h13e00001;
      78715: inst = 32'hfe0d96a;
      78716: inst = 32'h5be00000;
      78717: inst = 32'h8c50000;
      78718: inst = 32'h24612800;
      78719: inst = 32'h10a00000;
      78720: inst = 32'hca00000;
      78721: inst = 32'h24822800;
      78722: inst = 32'h10a00000;
      78723: inst = 32'hca00004;
      78724: inst = 32'h38632800;
      78725: inst = 32'h38842800;
      78726: inst = 32'h10a00001;
      78727: inst = 32'hca0338b;
      78728: inst = 32'h13e00001;
      78729: inst = 32'hfe0d96a;
      78730: inst = 32'h5be00000;
      78731: inst = 32'h8c50000;
      78732: inst = 32'h24612800;
      78733: inst = 32'h10a00000;
      78734: inst = 32'hca00000;
      78735: inst = 32'h24822800;
      78736: inst = 32'h10a00000;
      78737: inst = 32'hca00004;
      78738: inst = 32'h38632800;
      78739: inst = 32'h38842800;
      78740: inst = 32'h10a00001;
      78741: inst = 32'hca03399;
      78742: inst = 32'h13e00001;
      78743: inst = 32'hfe0d96a;
      78744: inst = 32'h5be00000;
      78745: inst = 32'h8c50000;
      78746: inst = 32'h24612800;
      78747: inst = 32'h10a00000;
      78748: inst = 32'hca00000;
      78749: inst = 32'h24822800;
      78750: inst = 32'h10a00000;
      78751: inst = 32'hca00004;
      78752: inst = 32'h38632800;
      78753: inst = 32'h38842800;
      78754: inst = 32'h10a00001;
      78755: inst = 32'hca033a7;
      78756: inst = 32'h13e00001;
      78757: inst = 32'hfe0d96a;
      78758: inst = 32'h5be00000;
      78759: inst = 32'h8c50000;
      78760: inst = 32'h24612800;
      78761: inst = 32'h10a00000;
      78762: inst = 32'hca00000;
      78763: inst = 32'h24822800;
      78764: inst = 32'h10a00000;
      78765: inst = 32'hca00004;
      78766: inst = 32'h38632800;
      78767: inst = 32'h38842800;
      78768: inst = 32'h10a00001;
      78769: inst = 32'hca033b5;
      78770: inst = 32'h13e00001;
      78771: inst = 32'hfe0d96a;
      78772: inst = 32'h5be00000;
      78773: inst = 32'h8c50000;
      78774: inst = 32'h24612800;
      78775: inst = 32'h10a00000;
      78776: inst = 32'hca00000;
      78777: inst = 32'h24822800;
      78778: inst = 32'h10a00000;
      78779: inst = 32'hca00004;
      78780: inst = 32'h38632800;
      78781: inst = 32'h38842800;
      78782: inst = 32'h10a00001;
      78783: inst = 32'hca033c3;
      78784: inst = 32'h13e00001;
      78785: inst = 32'hfe0d96a;
      78786: inst = 32'h5be00000;
      78787: inst = 32'h8c50000;
      78788: inst = 32'h24612800;
      78789: inst = 32'h10a00000;
      78790: inst = 32'hca00000;
      78791: inst = 32'h24822800;
      78792: inst = 32'h10a00000;
      78793: inst = 32'hca00004;
      78794: inst = 32'h38632800;
      78795: inst = 32'h38842800;
      78796: inst = 32'h10a00001;
      78797: inst = 32'hca033d1;
      78798: inst = 32'h13e00001;
      78799: inst = 32'hfe0d96a;
      78800: inst = 32'h5be00000;
      78801: inst = 32'h8c50000;
      78802: inst = 32'h24612800;
      78803: inst = 32'h10a00000;
      78804: inst = 32'hca00000;
      78805: inst = 32'h24822800;
      78806: inst = 32'h10a00000;
      78807: inst = 32'hca00004;
      78808: inst = 32'h38632800;
      78809: inst = 32'h38842800;
      78810: inst = 32'h10a00001;
      78811: inst = 32'hca033df;
      78812: inst = 32'h13e00001;
      78813: inst = 32'hfe0d96a;
      78814: inst = 32'h5be00000;
      78815: inst = 32'h8c50000;
      78816: inst = 32'h24612800;
      78817: inst = 32'h10a00000;
      78818: inst = 32'hca00000;
      78819: inst = 32'h24822800;
      78820: inst = 32'h10a00000;
      78821: inst = 32'hca00004;
      78822: inst = 32'h38632800;
      78823: inst = 32'h38842800;
      78824: inst = 32'h10a00001;
      78825: inst = 32'hca033ed;
      78826: inst = 32'h13e00001;
      78827: inst = 32'hfe0d96a;
      78828: inst = 32'h5be00000;
      78829: inst = 32'h8c50000;
      78830: inst = 32'h24612800;
      78831: inst = 32'h10a00000;
      78832: inst = 32'hca00000;
      78833: inst = 32'h24822800;
      78834: inst = 32'h10a00000;
      78835: inst = 32'hca00004;
      78836: inst = 32'h38632800;
      78837: inst = 32'h38842800;
      78838: inst = 32'h10a00001;
      78839: inst = 32'hca033fb;
      78840: inst = 32'h13e00001;
      78841: inst = 32'hfe0d96a;
      78842: inst = 32'h5be00000;
      78843: inst = 32'h8c50000;
      78844: inst = 32'h24612800;
      78845: inst = 32'h10a00000;
      78846: inst = 32'hca00000;
      78847: inst = 32'h24822800;
      78848: inst = 32'h10a00000;
      78849: inst = 32'hca00004;
      78850: inst = 32'h38632800;
      78851: inst = 32'h38842800;
      78852: inst = 32'h10a00001;
      78853: inst = 32'hca03409;
      78854: inst = 32'h13e00001;
      78855: inst = 32'hfe0d96a;
      78856: inst = 32'h5be00000;
      78857: inst = 32'h8c50000;
      78858: inst = 32'h24612800;
      78859: inst = 32'h10a00000;
      78860: inst = 32'hca00000;
      78861: inst = 32'h24822800;
      78862: inst = 32'h10a00000;
      78863: inst = 32'hca00004;
      78864: inst = 32'h38632800;
      78865: inst = 32'h38842800;
      78866: inst = 32'h10a00001;
      78867: inst = 32'hca03417;
      78868: inst = 32'h13e00001;
      78869: inst = 32'hfe0d96a;
      78870: inst = 32'h5be00000;
      78871: inst = 32'h8c50000;
      78872: inst = 32'h24612800;
      78873: inst = 32'h10a00000;
      78874: inst = 32'hca00000;
      78875: inst = 32'h24822800;
      78876: inst = 32'h10a00000;
      78877: inst = 32'hca00004;
      78878: inst = 32'h38632800;
      78879: inst = 32'h38842800;
      78880: inst = 32'h10a00001;
      78881: inst = 32'hca03425;
      78882: inst = 32'h13e00001;
      78883: inst = 32'hfe0d96a;
      78884: inst = 32'h5be00000;
      78885: inst = 32'h8c50000;
      78886: inst = 32'h24612800;
      78887: inst = 32'h10a00000;
      78888: inst = 32'hca00000;
      78889: inst = 32'h24822800;
      78890: inst = 32'h10a00000;
      78891: inst = 32'hca00004;
      78892: inst = 32'h38632800;
      78893: inst = 32'h38842800;
      78894: inst = 32'h10a00001;
      78895: inst = 32'hca03433;
      78896: inst = 32'h13e00001;
      78897: inst = 32'hfe0d96a;
      78898: inst = 32'h5be00000;
      78899: inst = 32'h8c50000;
      78900: inst = 32'h24612800;
      78901: inst = 32'h10a00000;
      78902: inst = 32'hca00000;
      78903: inst = 32'h24822800;
      78904: inst = 32'h10a00000;
      78905: inst = 32'hca00004;
      78906: inst = 32'h38632800;
      78907: inst = 32'h38842800;
      78908: inst = 32'h10a00001;
      78909: inst = 32'hca03441;
      78910: inst = 32'h13e00001;
      78911: inst = 32'hfe0d96a;
      78912: inst = 32'h5be00000;
      78913: inst = 32'h8c50000;
      78914: inst = 32'h24612800;
      78915: inst = 32'h10a00000;
      78916: inst = 32'hca00000;
      78917: inst = 32'h24822800;
      78918: inst = 32'h10a00000;
      78919: inst = 32'hca00004;
      78920: inst = 32'h38632800;
      78921: inst = 32'h38842800;
      78922: inst = 32'h10a00001;
      78923: inst = 32'hca0344f;
      78924: inst = 32'h13e00001;
      78925: inst = 32'hfe0d96a;
      78926: inst = 32'h5be00000;
      78927: inst = 32'h8c50000;
      78928: inst = 32'h24612800;
      78929: inst = 32'h10a00000;
      78930: inst = 32'hca00000;
      78931: inst = 32'h24822800;
      78932: inst = 32'h10a00000;
      78933: inst = 32'hca00004;
      78934: inst = 32'h38632800;
      78935: inst = 32'h38842800;
      78936: inst = 32'h10a00001;
      78937: inst = 32'hca0345d;
      78938: inst = 32'h13e00001;
      78939: inst = 32'hfe0d96a;
      78940: inst = 32'h5be00000;
      78941: inst = 32'h8c50000;
      78942: inst = 32'h24612800;
      78943: inst = 32'h10a00000;
      78944: inst = 32'hca00000;
      78945: inst = 32'h24822800;
      78946: inst = 32'h10a00000;
      78947: inst = 32'hca00004;
      78948: inst = 32'h38632800;
      78949: inst = 32'h38842800;
      78950: inst = 32'h10a00001;
      78951: inst = 32'hca0346b;
      78952: inst = 32'h13e00001;
      78953: inst = 32'hfe0d96a;
      78954: inst = 32'h5be00000;
      78955: inst = 32'h8c50000;
      78956: inst = 32'h24612800;
      78957: inst = 32'h10a00000;
      78958: inst = 32'hca00000;
      78959: inst = 32'h24822800;
      78960: inst = 32'h10a00000;
      78961: inst = 32'hca00004;
      78962: inst = 32'h38632800;
      78963: inst = 32'h38842800;
      78964: inst = 32'h10a00001;
      78965: inst = 32'hca03479;
      78966: inst = 32'h13e00001;
      78967: inst = 32'hfe0d96a;
      78968: inst = 32'h5be00000;
      78969: inst = 32'h8c50000;
      78970: inst = 32'h24612800;
      78971: inst = 32'h10a00000;
      78972: inst = 32'hca00000;
      78973: inst = 32'h24822800;
      78974: inst = 32'h10a00000;
      78975: inst = 32'hca00004;
      78976: inst = 32'h38632800;
      78977: inst = 32'h38842800;
      78978: inst = 32'h10a00001;
      78979: inst = 32'hca03487;
      78980: inst = 32'h13e00001;
      78981: inst = 32'hfe0d96a;
      78982: inst = 32'h5be00000;
      78983: inst = 32'h8c50000;
      78984: inst = 32'h24612800;
      78985: inst = 32'h10a00000;
      78986: inst = 32'hca00000;
      78987: inst = 32'h24822800;
      78988: inst = 32'h10a00000;
      78989: inst = 32'hca00004;
      78990: inst = 32'h38632800;
      78991: inst = 32'h38842800;
      78992: inst = 32'h10a00001;
      78993: inst = 32'hca03495;
      78994: inst = 32'h13e00001;
      78995: inst = 32'hfe0d96a;
      78996: inst = 32'h5be00000;
      78997: inst = 32'h8c50000;
      78998: inst = 32'h24612800;
      78999: inst = 32'h10a00000;
      79000: inst = 32'hca00000;
      79001: inst = 32'h24822800;
      79002: inst = 32'h10a00000;
      79003: inst = 32'hca00004;
      79004: inst = 32'h38632800;
      79005: inst = 32'h38842800;
      79006: inst = 32'h10a00001;
      79007: inst = 32'hca034a3;
      79008: inst = 32'h13e00001;
      79009: inst = 32'hfe0d96a;
      79010: inst = 32'h5be00000;
      79011: inst = 32'h8c50000;
      79012: inst = 32'h24612800;
      79013: inst = 32'h10a00000;
      79014: inst = 32'hca00000;
      79015: inst = 32'h24822800;
      79016: inst = 32'h10a00000;
      79017: inst = 32'hca00004;
      79018: inst = 32'h38632800;
      79019: inst = 32'h38842800;
      79020: inst = 32'h10a00001;
      79021: inst = 32'hca034b1;
      79022: inst = 32'h13e00001;
      79023: inst = 32'hfe0d96a;
      79024: inst = 32'h5be00000;
      79025: inst = 32'h8c50000;
      79026: inst = 32'h24612800;
      79027: inst = 32'h10a00000;
      79028: inst = 32'hca00000;
      79029: inst = 32'h24822800;
      79030: inst = 32'h10a00000;
      79031: inst = 32'hca00004;
      79032: inst = 32'h38632800;
      79033: inst = 32'h38842800;
      79034: inst = 32'h10a00001;
      79035: inst = 32'hca034bf;
      79036: inst = 32'h13e00001;
      79037: inst = 32'hfe0d96a;
      79038: inst = 32'h5be00000;
      79039: inst = 32'h8c50000;
      79040: inst = 32'h24612800;
      79041: inst = 32'h10a00000;
      79042: inst = 32'hca00000;
      79043: inst = 32'h24822800;
      79044: inst = 32'h10a00000;
      79045: inst = 32'hca00004;
      79046: inst = 32'h38632800;
      79047: inst = 32'h38842800;
      79048: inst = 32'h10a00001;
      79049: inst = 32'hca034cd;
      79050: inst = 32'h13e00001;
      79051: inst = 32'hfe0d96a;
      79052: inst = 32'h5be00000;
      79053: inst = 32'h8c50000;
      79054: inst = 32'h24612800;
      79055: inst = 32'h10a00000;
      79056: inst = 32'hca00000;
      79057: inst = 32'h24822800;
      79058: inst = 32'h10a00000;
      79059: inst = 32'hca00004;
      79060: inst = 32'h38632800;
      79061: inst = 32'h38842800;
      79062: inst = 32'h10a00001;
      79063: inst = 32'hca034db;
      79064: inst = 32'h13e00001;
      79065: inst = 32'hfe0d96a;
      79066: inst = 32'h5be00000;
      79067: inst = 32'h8c50000;
      79068: inst = 32'h24612800;
      79069: inst = 32'h10a00000;
      79070: inst = 32'hca00000;
      79071: inst = 32'h24822800;
      79072: inst = 32'h10a00000;
      79073: inst = 32'hca00004;
      79074: inst = 32'h38632800;
      79075: inst = 32'h38842800;
      79076: inst = 32'h10a00001;
      79077: inst = 32'hca034e9;
      79078: inst = 32'h13e00001;
      79079: inst = 32'hfe0d96a;
      79080: inst = 32'h5be00000;
      79081: inst = 32'h8c50000;
      79082: inst = 32'h24612800;
      79083: inst = 32'h10a00000;
      79084: inst = 32'hca00000;
      79085: inst = 32'h24822800;
      79086: inst = 32'h10a00000;
      79087: inst = 32'hca00004;
      79088: inst = 32'h38632800;
      79089: inst = 32'h38842800;
      79090: inst = 32'h10a00001;
      79091: inst = 32'hca034f7;
      79092: inst = 32'h13e00001;
      79093: inst = 32'hfe0d96a;
      79094: inst = 32'h5be00000;
      79095: inst = 32'h8c50000;
      79096: inst = 32'h24612800;
      79097: inst = 32'h10a00000;
      79098: inst = 32'hca00000;
      79099: inst = 32'h24822800;
      79100: inst = 32'h10a00000;
      79101: inst = 32'hca00004;
      79102: inst = 32'h38632800;
      79103: inst = 32'h38842800;
      79104: inst = 32'h10a00001;
      79105: inst = 32'hca03505;
      79106: inst = 32'h13e00001;
      79107: inst = 32'hfe0d96a;
      79108: inst = 32'h5be00000;
      79109: inst = 32'h8c50000;
      79110: inst = 32'h24612800;
      79111: inst = 32'h10a00000;
      79112: inst = 32'hca00000;
      79113: inst = 32'h24822800;
      79114: inst = 32'h10a00000;
      79115: inst = 32'hca00004;
      79116: inst = 32'h38632800;
      79117: inst = 32'h38842800;
      79118: inst = 32'h10a00001;
      79119: inst = 32'hca03513;
      79120: inst = 32'h13e00001;
      79121: inst = 32'hfe0d96a;
      79122: inst = 32'h5be00000;
      79123: inst = 32'h8c50000;
      79124: inst = 32'h24612800;
      79125: inst = 32'h10a00000;
      79126: inst = 32'hca00000;
      79127: inst = 32'h24822800;
      79128: inst = 32'h10a00000;
      79129: inst = 32'hca00004;
      79130: inst = 32'h38632800;
      79131: inst = 32'h38842800;
      79132: inst = 32'h10a00001;
      79133: inst = 32'hca03521;
      79134: inst = 32'h13e00001;
      79135: inst = 32'hfe0d96a;
      79136: inst = 32'h5be00000;
      79137: inst = 32'h8c50000;
      79138: inst = 32'h24612800;
      79139: inst = 32'h10a00000;
      79140: inst = 32'hca00000;
      79141: inst = 32'h24822800;
      79142: inst = 32'h10a00000;
      79143: inst = 32'hca00004;
      79144: inst = 32'h38632800;
      79145: inst = 32'h38842800;
      79146: inst = 32'h10a00001;
      79147: inst = 32'hca0352f;
      79148: inst = 32'h13e00001;
      79149: inst = 32'hfe0d96a;
      79150: inst = 32'h5be00000;
      79151: inst = 32'h8c50000;
      79152: inst = 32'h24612800;
      79153: inst = 32'h10a00000;
      79154: inst = 32'hca00000;
      79155: inst = 32'h24822800;
      79156: inst = 32'h10a00000;
      79157: inst = 32'hca00004;
      79158: inst = 32'h38632800;
      79159: inst = 32'h38842800;
      79160: inst = 32'h10a00001;
      79161: inst = 32'hca0353d;
      79162: inst = 32'h13e00001;
      79163: inst = 32'hfe0d96a;
      79164: inst = 32'h5be00000;
      79165: inst = 32'h8c50000;
      79166: inst = 32'h24612800;
      79167: inst = 32'h10a00000;
      79168: inst = 32'hca00000;
      79169: inst = 32'h24822800;
      79170: inst = 32'h10a00000;
      79171: inst = 32'hca00004;
      79172: inst = 32'h38632800;
      79173: inst = 32'h38842800;
      79174: inst = 32'h10a00001;
      79175: inst = 32'hca0354b;
      79176: inst = 32'h13e00001;
      79177: inst = 32'hfe0d96a;
      79178: inst = 32'h5be00000;
      79179: inst = 32'h8c50000;
      79180: inst = 32'h24612800;
      79181: inst = 32'h10a00000;
      79182: inst = 32'hca00000;
      79183: inst = 32'h24822800;
      79184: inst = 32'h10a00000;
      79185: inst = 32'hca00004;
      79186: inst = 32'h38632800;
      79187: inst = 32'h38842800;
      79188: inst = 32'h10a00001;
      79189: inst = 32'hca03559;
      79190: inst = 32'h13e00001;
      79191: inst = 32'hfe0d96a;
      79192: inst = 32'h5be00000;
      79193: inst = 32'h8c50000;
      79194: inst = 32'h24612800;
      79195: inst = 32'h10a00000;
      79196: inst = 32'hca00000;
      79197: inst = 32'h24822800;
      79198: inst = 32'h10a00000;
      79199: inst = 32'hca00004;
      79200: inst = 32'h38632800;
      79201: inst = 32'h38842800;
      79202: inst = 32'h10a00001;
      79203: inst = 32'hca03567;
      79204: inst = 32'h13e00001;
      79205: inst = 32'hfe0d96a;
      79206: inst = 32'h5be00000;
      79207: inst = 32'h8c50000;
      79208: inst = 32'h24612800;
      79209: inst = 32'h10a00000;
      79210: inst = 32'hca00000;
      79211: inst = 32'h24822800;
      79212: inst = 32'h10a00000;
      79213: inst = 32'hca00004;
      79214: inst = 32'h38632800;
      79215: inst = 32'h38842800;
      79216: inst = 32'h10a00001;
      79217: inst = 32'hca03575;
      79218: inst = 32'h13e00001;
      79219: inst = 32'hfe0d96a;
      79220: inst = 32'h5be00000;
      79221: inst = 32'h8c50000;
      79222: inst = 32'h24612800;
      79223: inst = 32'h10a00000;
      79224: inst = 32'hca00000;
      79225: inst = 32'h24822800;
      79226: inst = 32'h10a00000;
      79227: inst = 32'hca00004;
      79228: inst = 32'h38632800;
      79229: inst = 32'h38842800;
      79230: inst = 32'h10a00001;
      79231: inst = 32'hca03583;
      79232: inst = 32'h13e00001;
      79233: inst = 32'hfe0d96a;
      79234: inst = 32'h5be00000;
      79235: inst = 32'h8c50000;
      79236: inst = 32'h24612800;
      79237: inst = 32'h10a00000;
      79238: inst = 32'hca00000;
      79239: inst = 32'h24822800;
      79240: inst = 32'h10a00000;
      79241: inst = 32'hca00004;
      79242: inst = 32'h38632800;
      79243: inst = 32'h38842800;
      79244: inst = 32'h10a00001;
      79245: inst = 32'hca03591;
      79246: inst = 32'h13e00001;
      79247: inst = 32'hfe0d96a;
      79248: inst = 32'h5be00000;
      79249: inst = 32'h8c50000;
      79250: inst = 32'h24612800;
      79251: inst = 32'h10a00000;
      79252: inst = 32'hca00000;
      79253: inst = 32'h24822800;
      79254: inst = 32'h10a00000;
      79255: inst = 32'hca00004;
      79256: inst = 32'h38632800;
      79257: inst = 32'h38842800;
      79258: inst = 32'h10a00001;
      79259: inst = 32'hca0359f;
      79260: inst = 32'h13e00001;
      79261: inst = 32'hfe0d96a;
      79262: inst = 32'h5be00000;
      79263: inst = 32'h8c50000;
      79264: inst = 32'h24612800;
      79265: inst = 32'h10a00000;
      79266: inst = 32'hca00000;
      79267: inst = 32'h24822800;
      79268: inst = 32'h10a00000;
      79269: inst = 32'hca00004;
      79270: inst = 32'h38632800;
      79271: inst = 32'h38842800;
      79272: inst = 32'h10a00001;
      79273: inst = 32'hca035ad;
      79274: inst = 32'h13e00001;
      79275: inst = 32'hfe0d96a;
      79276: inst = 32'h5be00000;
      79277: inst = 32'h8c50000;
      79278: inst = 32'h24612800;
      79279: inst = 32'h10a00000;
      79280: inst = 32'hca00000;
      79281: inst = 32'h24822800;
      79282: inst = 32'h10a00000;
      79283: inst = 32'hca00004;
      79284: inst = 32'h38632800;
      79285: inst = 32'h38842800;
      79286: inst = 32'h10a00001;
      79287: inst = 32'hca035bb;
      79288: inst = 32'h13e00001;
      79289: inst = 32'hfe0d96a;
      79290: inst = 32'h5be00000;
      79291: inst = 32'h8c50000;
      79292: inst = 32'h24612800;
      79293: inst = 32'h10a00000;
      79294: inst = 32'hca00000;
      79295: inst = 32'h24822800;
      79296: inst = 32'h10a00000;
      79297: inst = 32'hca00004;
      79298: inst = 32'h38632800;
      79299: inst = 32'h38842800;
      79300: inst = 32'h10a00001;
      79301: inst = 32'hca035c9;
      79302: inst = 32'h13e00001;
      79303: inst = 32'hfe0d96a;
      79304: inst = 32'h5be00000;
      79305: inst = 32'h8c50000;
      79306: inst = 32'h24612800;
      79307: inst = 32'h10a00000;
      79308: inst = 32'hca00000;
      79309: inst = 32'h24822800;
      79310: inst = 32'h10a00000;
      79311: inst = 32'hca00004;
      79312: inst = 32'h38632800;
      79313: inst = 32'h38842800;
      79314: inst = 32'h10a00001;
      79315: inst = 32'hca035d7;
      79316: inst = 32'h13e00001;
      79317: inst = 32'hfe0d96a;
      79318: inst = 32'h5be00000;
      79319: inst = 32'h8c50000;
      79320: inst = 32'h24612800;
      79321: inst = 32'h10a00000;
      79322: inst = 32'hca00000;
      79323: inst = 32'h24822800;
      79324: inst = 32'h10a00000;
      79325: inst = 32'hca00004;
      79326: inst = 32'h38632800;
      79327: inst = 32'h38842800;
      79328: inst = 32'h10a00001;
      79329: inst = 32'hca035e5;
      79330: inst = 32'h13e00001;
      79331: inst = 32'hfe0d96a;
      79332: inst = 32'h5be00000;
      79333: inst = 32'h8c50000;
      79334: inst = 32'h24612800;
      79335: inst = 32'h10a00000;
      79336: inst = 32'hca00000;
      79337: inst = 32'h24822800;
      79338: inst = 32'h10a00000;
      79339: inst = 32'hca00004;
      79340: inst = 32'h38632800;
      79341: inst = 32'h38842800;
      79342: inst = 32'h10a00001;
      79343: inst = 32'hca035f3;
      79344: inst = 32'h13e00001;
      79345: inst = 32'hfe0d96a;
      79346: inst = 32'h5be00000;
      79347: inst = 32'h8c50000;
      79348: inst = 32'h24612800;
      79349: inst = 32'h10a00000;
      79350: inst = 32'hca00000;
      79351: inst = 32'h24822800;
      79352: inst = 32'h10a00000;
      79353: inst = 32'hca00004;
      79354: inst = 32'h38632800;
      79355: inst = 32'h38842800;
      79356: inst = 32'h10a00001;
      79357: inst = 32'hca03601;
      79358: inst = 32'h13e00001;
      79359: inst = 32'hfe0d96a;
      79360: inst = 32'h5be00000;
      79361: inst = 32'h8c50000;
      79362: inst = 32'h24612800;
      79363: inst = 32'h10a00000;
      79364: inst = 32'hca00000;
      79365: inst = 32'h24822800;
      79366: inst = 32'h10a00000;
      79367: inst = 32'hca00004;
      79368: inst = 32'h38632800;
      79369: inst = 32'h38842800;
      79370: inst = 32'h10a00001;
      79371: inst = 32'hca0360f;
      79372: inst = 32'h13e00001;
      79373: inst = 32'hfe0d96a;
      79374: inst = 32'h5be00000;
      79375: inst = 32'h8c50000;
      79376: inst = 32'h24612800;
      79377: inst = 32'h10a00000;
      79378: inst = 32'hca00000;
      79379: inst = 32'h24822800;
      79380: inst = 32'h10a00000;
      79381: inst = 32'hca00004;
      79382: inst = 32'h38632800;
      79383: inst = 32'h38842800;
      79384: inst = 32'h10a00001;
      79385: inst = 32'hca0361d;
      79386: inst = 32'h13e00001;
      79387: inst = 32'hfe0d96a;
      79388: inst = 32'h5be00000;
      79389: inst = 32'h8c50000;
      79390: inst = 32'h24612800;
      79391: inst = 32'h10a00000;
      79392: inst = 32'hca00000;
      79393: inst = 32'h24822800;
      79394: inst = 32'h10a00000;
      79395: inst = 32'hca00004;
      79396: inst = 32'h38632800;
      79397: inst = 32'h38842800;
      79398: inst = 32'h10a00001;
      79399: inst = 32'hca0362b;
      79400: inst = 32'h13e00001;
      79401: inst = 32'hfe0d96a;
      79402: inst = 32'h5be00000;
      79403: inst = 32'h8c50000;
      79404: inst = 32'h24612800;
      79405: inst = 32'h10a00000;
      79406: inst = 32'hca00000;
      79407: inst = 32'h24822800;
      79408: inst = 32'h10a00000;
      79409: inst = 32'hca00004;
      79410: inst = 32'h38632800;
      79411: inst = 32'h38842800;
      79412: inst = 32'h10a00001;
      79413: inst = 32'hca03639;
      79414: inst = 32'h13e00001;
      79415: inst = 32'hfe0d96a;
      79416: inst = 32'h5be00000;
      79417: inst = 32'h8c50000;
      79418: inst = 32'h24612800;
      79419: inst = 32'h10a00000;
      79420: inst = 32'hca00000;
      79421: inst = 32'h24822800;
      79422: inst = 32'h10a00000;
      79423: inst = 32'hca00004;
      79424: inst = 32'h38632800;
      79425: inst = 32'h38842800;
      79426: inst = 32'h10a00001;
      79427: inst = 32'hca03647;
      79428: inst = 32'h13e00001;
      79429: inst = 32'hfe0d96a;
      79430: inst = 32'h5be00000;
      79431: inst = 32'h8c50000;
      79432: inst = 32'h24612800;
      79433: inst = 32'h10a00000;
      79434: inst = 32'hca00000;
      79435: inst = 32'h24822800;
      79436: inst = 32'h10a00000;
      79437: inst = 32'hca00004;
      79438: inst = 32'h38632800;
      79439: inst = 32'h38842800;
      79440: inst = 32'h10a00001;
      79441: inst = 32'hca03655;
      79442: inst = 32'h13e00001;
      79443: inst = 32'hfe0d96a;
      79444: inst = 32'h5be00000;
      79445: inst = 32'h8c50000;
      79446: inst = 32'h24612800;
      79447: inst = 32'h10a00000;
      79448: inst = 32'hca00000;
      79449: inst = 32'h24822800;
      79450: inst = 32'h10a00000;
      79451: inst = 32'hca00004;
      79452: inst = 32'h38632800;
      79453: inst = 32'h38842800;
      79454: inst = 32'h10a00001;
      79455: inst = 32'hca03663;
      79456: inst = 32'h13e00001;
      79457: inst = 32'hfe0d96a;
      79458: inst = 32'h5be00000;
      79459: inst = 32'h8c50000;
      79460: inst = 32'h24612800;
      79461: inst = 32'h10a00000;
      79462: inst = 32'hca00000;
      79463: inst = 32'h24822800;
      79464: inst = 32'h10a00000;
      79465: inst = 32'hca00004;
      79466: inst = 32'h38632800;
      79467: inst = 32'h38842800;
      79468: inst = 32'h10a00001;
      79469: inst = 32'hca03671;
      79470: inst = 32'h13e00001;
      79471: inst = 32'hfe0d96a;
      79472: inst = 32'h5be00000;
      79473: inst = 32'h8c50000;
      79474: inst = 32'h24612800;
      79475: inst = 32'h10a00000;
      79476: inst = 32'hca00000;
      79477: inst = 32'h24822800;
      79478: inst = 32'h10a00000;
      79479: inst = 32'hca00004;
      79480: inst = 32'h38632800;
      79481: inst = 32'h38842800;
      79482: inst = 32'h10a00001;
      79483: inst = 32'hca0367f;
      79484: inst = 32'h13e00001;
      79485: inst = 32'hfe0d96a;
      79486: inst = 32'h5be00000;
      79487: inst = 32'h8c50000;
      79488: inst = 32'h24612800;
      79489: inst = 32'h10a00000;
      79490: inst = 32'hca00000;
      79491: inst = 32'h24822800;
      79492: inst = 32'h10a00000;
      79493: inst = 32'hca00004;
      79494: inst = 32'h38632800;
      79495: inst = 32'h38842800;
      79496: inst = 32'h10a00001;
      79497: inst = 32'hca0368d;
      79498: inst = 32'h13e00001;
      79499: inst = 32'hfe0d96a;
      79500: inst = 32'h5be00000;
      79501: inst = 32'h8c50000;
      79502: inst = 32'h24612800;
      79503: inst = 32'h10a00000;
      79504: inst = 32'hca00000;
      79505: inst = 32'h24822800;
      79506: inst = 32'h10a00000;
      79507: inst = 32'hca00004;
      79508: inst = 32'h38632800;
      79509: inst = 32'h38842800;
      79510: inst = 32'h10a00001;
      79511: inst = 32'hca0369b;
      79512: inst = 32'h13e00001;
      79513: inst = 32'hfe0d96a;
      79514: inst = 32'h5be00000;
      79515: inst = 32'h8c50000;
      79516: inst = 32'h24612800;
      79517: inst = 32'h10a00000;
      79518: inst = 32'hca00000;
      79519: inst = 32'h24822800;
      79520: inst = 32'h10a00000;
      79521: inst = 32'hca00004;
      79522: inst = 32'h38632800;
      79523: inst = 32'h38842800;
      79524: inst = 32'h10a00001;
      79525: inst = 32'hca036a9;
      79526: inst = 32'h13e00001;
      79527: inst = 32'hfe0d96a;
      79528: inst = 32'h5be00000;
      79529: inst = 32'h8c50000;
      79530: inst = 32'h24612800;
      79531: inst = 32'h10a00000;
      79532: inst = 32'hca00001;
      79533: inst = 32'h24822800;
      79534: inst = 32'h10a00000;
      79535: inst = 32'hca00004;
      79536: inst = 32'h38632800;
      79537: inst = 32'h38842800;
      79538: inst = 32'h10a00001;
      79539: inst = 32'hca036b7;
      79540: inst = 32'h13e00001;
      79541: inst = 32'hfe0d96a;
      79542: inst = 32'h5be00000;
      79543: inst = 32'h8c50000;
      79544: inst = 32'h24612800;
      79545: inst = 32'h10a00000;
      79546: inst = 32'hca00001;
      79547: inst = 32'h24822800;
      79548: inst = 32'h10a00000;
      79549: inst = 32'hca00004;
      79550: inst = 32'h38632800;
      79551: inst = 32'h38842800;
      79552: inst = 32'h10a00001;
      79553: inst = 32'hca036c5;
      79554: inst = 32'h13e00001;
      79555: inst = 32'hfe0d96a;
      79556: inst = 32'h5be00000;
      79557: inst = 32'h8c50000;
      79558: inst = 32'h24612800;
      79559: inst = 32'h10a00000;
      79560: inst = 32'hca00001;
      79561: inst = 32'h24822800;
      79562: inst = 32'h10a00000;
      79563: inst = 32'hca00004;
      79564: inst = 32'h38632800;
      79565: inst = 32'h38842800;
      79566: inst = 32'h10a00001;
      79567: inst = 32'hca036d3;
      79568: inst = 32'h13e00001;
      79569: inst = 32'hfe0d96a;
      79570: inst = 32'h5be00000;
      79571: inst = 32'h8c50000;
      79572: inst = 32'h24612800;
      79573: inst = 32'h10a00000;
      79574: inst = 32'hca00001;
      79575: inst = 32'h24822800;
      79576: inst = 32'h10a00000;
      79577: inst = 32'hca00004;
      79578: inst = 32'h38632800;
      79579: inst = 32'h38842800;
      79580: inst = 32'h10a00001;
      79581: inst = 32'hca036e1;
      79582: inst = 32'h13e00001;
      79583: inst = 32'hfe0d96a;
      79584: inst = 32'h5be00000;
      79585: inst = 32'h8c50000;
      79586: inst = 32'h24612800;
      79587: inst = 32'h10a00000;
      79588: inst = 32'hca00001;
      79589: inst = 32'h24822800;
      79590: inst = 32'h10a00000;
      79591: inst = 32'hca00004;
      79592: inst = 32'h38632800;
      79593: inst = 32'h38842800;
      79594: inst = 32'h10a00001;
      79595: inst = 32'hca036ef;
      79596: inst = 32'h13e00001;
      79597: inst = 32'hfe0d96a;
      79598: inst = 32'h5be00000;
      79599: inst = 32'h8c50000;
      79600: inst = 32'h24612800;
      79601: inst = 32'h10a00000;
      79602: inst = 32'hca00001;
      79603: inst = 32'h24822800;
      79604: inst = 32'h10a00000;
      79605: inst = 32'hca00004;
      79606: inst = 32'h38632800;
      79607: inst = 32'h38842800;
      79608: inst = 32'h10a00001;
      79609: inst = 32'hca036fd;
      79610: inst = 32'h13e00001;
      79611: inst = 32'hfe0d96a;
      79612: inst = 32'h5be00000;
      79613: inst = 32'h8c50000;
      79614: inst = 32'h24612800;
      79615: inst = 32'h10a00000;
      79616: inst = 32'hca00001;
      79617: inst = 32'h24822800;
      79618: inst = 32'h10a00000;
      79619: inst = 32'hca00004;
      79620: inst = 32'h38632800;
      79621: inst = 32'h38842800;
      79622: inst = 32'h10a00001;
      79623: inst = 32'hca0370b;
      79624: inst = 32'h13e00001;
      79625: inst = 32'hfe0d96a;
      79626: inst = 32'h5be00000;
      79627: inst = 32'h8c50000;
      79628: inst = 32'h24612800;
      79629: inst = 32'h10a00000;
      79630: inst = 32'hca00001;
      79631: inst = 32'h24822800;
      79632: inst = 32'h10a00000;
      79633: inst = 32'hca00004;
      79634: inst = 32'h38632800;
      79635: inst = 32'h38842800;
      79636: inst = 32'h10a00001;
      79637: inst = 32'hca03719;
      79638: inst = 32'h13e00001;
      79639: inst = 32'hfe0d96a;
      79640: inst = 32'h5be00000;
      79641: inst = 32'h8c50000;
      79642: inst = 32'h24612800;
      79643: inst = 32'h10a00000;
      79644: inst = 32'hca00001;
      79645: inst = 32'h24822800;
      79646: inst = 32'h10a00000;
      79647: inst = 32'hca00004;
      79648: inst = 32'h38632800;
      79649: inst = 32'h38842800;
      79650: inst = 32'h10a00001;
      79651: inst = 32'hca03727;
      79652: inst = 32'h13e00001;
      79653: inst = 32'hfe0d96a;
      79654: inst = 32'h5be00000;
      79655: inst = 32'h8c50000;
      79656: inst = 32'h24612800;
      79657: inst = 32'h10a00000;
      79658: inst = 32'hca00001;
      79659: inst = 32'h24822800;
      79660: inst = 32'h10a00000;
      79661: inst = 32'hca00004;
      79662: inst = 32'h38632800;
      79663: inst = 32'h38842800;
      79664: inst = 32'h10a00001;
      79665: inst = 32'hca03735;
      79666: inst = 32'h13e00001;
      79667: inst = 32'hfe0d96a;
      79668: inst = 32'h5be00000;
      79669: inst = 32'h8c50000;
      79670: inst = 32'h24612800;
      79671: inst = 32'h10a00000;
      79672: inst = 32'hca00001;
      79673: inst = 32'h24822800;
      79674: inst = 32'h10a00000;
      79675: inst = 32'hca00004;
      79676: inst = 32'h38632800;
      79677: inst = 32'h38842800;
      79678: inst = 32'h10a00001;
      79679: inst = 32'hca03743;
      79680: inst = 32'h13e00001;
      79681: inst = 32'hfe0d96a;
      79682: inst = 32'h5be00000;
      79683: inst = 32'h8c50000;
      79684: inst = 32'h24612800;
      79685: inst = 32'h10a00000;
      79686: inst = 32'hca00001;
      79687: inst = 32'h24822800;
      79688: inst = 32'h10a00000;
      79689: inst = 32'hca00004;
      79690: inst = 32'h38632800;
      79691: inst = 32'h38842800;
      79692: inst = 32'h10a00001;
      79693: inst = 32'hca03751;
      79694: inst = 32'h13e00001;
      79695: inst = 32'hfe0d96a;
      79696: inst = 32'h5be00000;
      79697: inst = 32'h8c50000;
      79698: inst = 32'h24612800;
      79699: inst = 32'h10a00000;
      79700: inst = 32'hca00001;
      79701: inst = 32'h24822800;
      79702: inst = 32'h10a00000;
      79703: inst = 32'hca00004;
      79704: inst = 32'h38632800;
      79705: inst = 32'h38842800;
      79706: inst = 32'h10a00001;
      79707: inst = 32'hca0375f;
      79708: inst = 32'h13e00001;
      79709: inst = 32'hfe0d96a;
      79710: inst = 32'h5be00000;
      79711: inst = 32'h8c50000;
      79712: inst = 32'h24612800;
      79713: inst = 32'h10a00000;
      79714: inst = 32'hca00001;
      79715: inst = 32'h24822800;
      79716: inst = 32'h10a00000;
      79717: inst = 32'hca00004;
      79718: inst = 32'h38632800;
      79719: inst = 32'h38842800;
      79720: inst = 32'h10a00001;
      79721: inst = 32'hca0376d;
      79722: inst = 32'h13e00001;
      79723: inst = 32'hfe0d96a;
      79724: inst = 32'h5be00000;
      79725: inst = 32'h8c50000;
      79726: inst = 32'h24612800;
      79727: inst = 32'h10a00000;
      79728: inst = 32'hca00001;
      79729: inst = 32'h24822800;
      79730: inst = 32'h10a00000;
      79731: inst = 32'hca00004;
      79732: inst = 32'h38632800;
      79733: inst = 32'h38842800;
      79734: inst = 32'h10a00001;
      79735: inst = 32'hca0377b;
      79736: inst = 32'h13e00001;
      79737: inst = 32'hfe0d96a;
      79738: inst = 32'h5be00000;
      79739: inst = 32'h8c50000;
      79740: inst = 32'h24612800;
      79741: inst = 32'h10a00000;
      79742: inst = 32'hca00001;
      79743: inst = 32'h24822800;
      79744: inst = 32'h10a00000;
      79745: inst = 32'hca00004;
      79746: inst = 32'h38632800;
      79747: inst = 32'h38842800;
      79748: inst = 32'h10a00001;
      79749: inst = 32'hca03789;
      79750: inst = 32'h13e00001;
      79751: inst = 32'hfe0d96a;
      79752: inst = 32'h5be00000;
      79753: inst = 32'h8c50000;
      79754: inst = 32'h24612800;
      79755: inst = 32'h10a00000;
      79756: inst = 32'hca00001;
      79757: inst = 32'h24822800;
      79758: inst = 32'h10a00000;
      79759: inst = 32'hca00004;
      79760: inst = 32'h38632800;
      79761: inst = 32'h38842800;
      79762: inst = 32'h10a00001;
      79763: inst = 32'hca03797;
      79764: inst = 32'h13e00001;
      79765: inst = 32'hfe0d96a;
      79766: inst = 32'h5be00000;
      79767: inst = 32'h8c50000;
      79768: inst = 32'h24612800;
      79769: inst = 32'h10a00000;
      79770: inst = 32'hca00001;
      79771: inst = 32'h24822800;
      79772: inst = 32'h10a00000;
      79773: inst = 32'hca00004;
      79774: inst = 32'h38632800;
      79775: inst = 32'h38842800;
      79776: inst = 32'h10a00001;
      79777: inst = 32'hca037a5;
      79778: inst = 32'h13e00001;
      79779: inst = 32'hfe0d96a;
      79780: inst = 32'h5be00000;
      79781: inst = 32'h8c50000;
      79782: inst = 32'h24612800;
      79783: inst = 32'h10a00000;
      79784: inst = 32'hca00001;
      79785: inst = 32'h24822800;
      79786: inst = 32'h10a00000;
      79787: inst = 32'hca00004;
      79788: inst = 32'h38632800;
      79789: inst = 32'h38842800;
      79790: inst = 32'h10a00001;
      79791: inst = 32'hca037b3;
      79792: inst = 32'h13e00001;
      79793: inst = 32'hfe0d96a;
      79794: inst = 32'h5be00000;
      79795: inst = 32'h8c50000;
      79796: inst = 32'h24612800;
      79797: inst = 32'h10a00000;
      79798: inst = 32'hca00001;
      79799: inst = 32'h24822800;
      79800: inst = 32'h10a00000;
      79801: inst = 32'hca00004;
      79802: inst = 32'h38632800;
      79803: inst = 32'h38842800;
      79804: inst = 32'h10a00001;
      79805: inst = 32'hca037c1;
      79806: inst = 32'h13e00001;
      79807: inst = 32'hfe0d96a;
      79808: inst = 32'h5be00000;
      79809: inst = 32'h8c50000;
      79810: inst = 32'h24612800;
      79811: inst = 32'h10a00000;
      79812: inst = 32'hca00001;
      79813: inst = 32'h24822800;
      79814: inst = 32'h10a00000;
      79815: inst = 32'hca00004;
      79816: inst = 32'h38632800;
      79817: inst = 32'h38842800;
      79818: inst = 32'h10a00001;
      79819: inst = 32'hca037cf;
      79820: inst = 32'h13e00001;
      79821: inst = 32'hfe0d96a;
      79822: inst = 32'h5be00000;
      79823: inst = 32'h8c50000;
      79824: inst = 32'h24612800;
      79825: inst = 32'h10a00000;
      79826: inst = 32'hca00001;
      79827: inst = 32'h24822800;
      79828: inst = 32'h10a00000;
      79829: inst = 32'hca00004;
      79830: inst = 32'h38632800;
      79831: inst = 32'h38842800;
      79832: inst = 32'h10a00001;
      79833: inst = 32'hca037dd;
      79834: inst = 32'h13e00001;
      79835: inst = 32'hfe0d96a;
      79836: inst = 32'h5be00000;
      79837: inst = 32'h8c50000;
      79838: inst = 32'h24612800;
      79839: inst = 32'h10a00000;
      79840: inst = 32'hca00001;
      79841: inst = 32'h24822800;
      79842: inst = 32'h10a00000;
      79843: inst = 32'hca00004;
      79844: inst = 32'h38632800;
      79845: inst = 32'h38842800;
      79846: inst = 32'h10a00001;
      79847: inst = 32'hca037eb;
      79848: inst = 32'h13e00001;
      79849: inst = 32'hfe0d96a;
      79850: inst = 32'h5be00000;
      79851: inst = 32'h8c50000;
      79852: inst = 32'h24612800;
      79853: inst = 32'h10a00000;
      79854: inst = 32'hca00001;
      79855: inst = 32'h24822800;
      79856: inst = 32'h10a00000;
      79857: inst = 32'hca00004;
      79858: inst = 32'h38632800;
      79859: inst = 32'h38842800;
      79860: inst = 32'h10a00001;
      79861: inst = 32'hca037f9;
      79862: inst = 32'h13e00001;
      79863: inst = 32'hfe0d96a;
      79864: inst = 32'h5be00000;
      79865: inst = 32'h8c50000;
      79866: inst = 32'h24612800;
      79867: inst = 32'h10a00000;
      79868: inst = 32'hca00001;
      79869: inst = 32'h24822800;
      79870: inst = 32'h10a00000;
      79871: inst = 32'hca00004;
      79872: inst = 32'h38632800;
      79873: inst = 32'h38842800;
      79874: inst = 32'h10a00001;
      79875: inst = 32'hca03807;
      79876: inst = 32'h13e00001;
      79877: inst = 32'hfe0d96a;
      79878: inst = 32'h5be00000;
      79879: inst = 32'h8c50000;
      79880: inst = 32'h24612800;
      79881: inst = 32'h10a00000;
      79882: inst = 32'hca00001;
      79883: inst = 32'h24822800;
      79884: inst = 32'h10a00000;
      79885: inst = 32'hca00004;
      79886: inst = 32'h38632800;
      79887: inst = 32'h38842800;
      79888: inst = 32'h10a00001;
      79889: inst = 32'hca03815;
      79890: inst = 32'h13e00001;
      79891: inst = 32'hfe0d96a;
      79892: inst = 32'h5be00000;
      79893: inst = 32'h8c50000;
      79894: inst = 32'h24612800;
      79895: inst = 32'h10a00000;
      79896: inst = 32'hca00001;
      79897: inst = 32'h24822800;
      79898: inst = 32'h10a00000;
      79899: inst = 32'hca00004;
      79900: inst = 32'h38632800;
      79901: inst = 32'h38842800;
      79902: inst = 32'h10a00001;
      79903: inst = 32'hca03823;
      79904: inst = 32'h13e00001;
      79905: inst = 32'hfe0d96a;
      79906: inst = 32'h5be00000;
      79907: inst = 32'h8c50000;
      79908: inst = 32'h24612800;
      79909: inst = 32'h10a00000;
      79910: inst = 32'hca00001;
      79911: inst = 32'h24822800;
      79912: inst = 32'h10a00000;
      79913: inst = 32'hca00004;
      79914: inst = 32'h38632800;
      79915: inst = 32'h38842800;
      79916: inst = 32'h10a00001;
      79917: inst = 32'hca03831;
      79918: inst = 32'h13e00001;
      79919: inst = 32'hfe0d96a;
      79920: inst = 32'h5be00000;
      79921: inst = 32'h8c50000;
      79922: inst = 32'h24612800;
      79923: inst = 32'h10a00000;
      79924: inst = 32'hca00001;
      79925: inst = 32'h24822800;
      79926: inst = 32'h10a00000;
      79927: inst = 32'hca00004;
      79928: inst = 32'h38632800;
      79929: inst = 32'h38842800;
      79930: inst = 32'h10a00001;
      79931: inst = 32'hca0383f;
      79932: inst = 32'h13e00001;
      79933: inst = 32'hfe0d96a;
      79934: inst = 32'h5be00000;
      79935: inst = 32'h8c50000;
      79936: inst = 32'h24612800;
      79937: inst = 32'h10a00000;
      79938: inst = 32'hca00001;
      79939: inst = 32'h24822800;
      79940: inst = 32'h10a00000;
      79941: inst = 32'hca00004;
      79942: inst = 32'h38632800;
      79943: inst = 32'h38842800;
      79944: inst = 32'h10a00001;
      79945: inst = 32'hca0384d;
      79946: inst = 32'h13e00001;
      79947: inst = 32'hfe0d96a;
      79948: inst = 32'h5be00000;
      79949: inst = 32'h8c50000;
      79950: inst = 32'h24612800;
      79951: inst = 32'h10a00000;
      79952: inst = 32'hca00001;
      79953: inst = 32'h24822800;
      79954: inst = 32'h10a00000;
      79955: inst = 32'hca00004;
      79956: inst = 32'h38632800;
      79957: inst = 32'h38842800;
      79958: inst = 32'h10a00001;
      79959: inst = 32'hca0385b;
      79960: inst = 32'h13e00001;
      79961: inst = 32'hfe0d96a;
      79962: inst = 32'h5be00000;
      79963: inst = 32'h8c50000;
      79964: inst = 32'h24612800;
      79965: inst = 32'h10a00000;
      79966: inst = 32'hca00001;
      79967: inst = 32'h24822800;
      79968: inst = 32'h10a00000;
      79969: inst = 32'hca00004;
      79970: inst = 32'h38632800;
      79971: inst = 32'h38842800;
      79972: inst = 32'h10a00001;
      79973: inst = 32'hca03869;
      79974: inst = 32'h13e00001;
      79975: inst = 32'hfe0d96a;
      79976: inst = 32'h5be00000;
      79977: inst = 32'h8c50000;
      79978: inst = 32'h24612800;
      79979: inst = 32'h10a00000;
      79980: inst = 32'hca00001;
      79981: inst = 32'h24822800;
      79982: inst = 32'h10a00000;
      79983: inst = 32'hca00004;
      79984: inst = 32'h38632800;
      79985: inst = 32'h38842800;
      79986: inst = 32'h10a00001;
      79987: inst = 32'hca03877;
      79988: inst = 32'h13e00001;
      79989: inst = 32'hfe0d96a;
      79990: inst = 32'h5be00000;
      79991: inst = 32'h8c50000;
      79992: inst = 32'h24612800;
      79993: inst = 32'h10a00000;
      79994: inst = 32'hca00001;
      79995: inst = 32'h24822800;
      79996: inst = 32'h10a00000;
      79997: inst = 32'hca00004;
      79998: inst = 32'h38632800;
      79999: inst = 32'h38842800;
      80000: inst = 32'h10a00001;
      80001: inst = 32'hca03885;
      80002: inst = 32'h13e00001;
      80003: inst = 32'hfe0d96a;
      80004: inst = 32'h5be00000;
      80005: inst = 32'h8c50000;
      80006: inst = 32'h24612800;
      80007: inst = 32'h10a00000;
      80008: inst = 32'hca00001;
      80009: inst = 32'h24822800;
      80010: inst = 32'h10a00000;
      80011: inst = 32'hca00004;
      80012: inst = 32'h38632800;
      80013: inst = 32'h38842800;
      80014: inst = 32'h10a00001;
      80015: inst = 32'hca03893;
      80016: inst = 32'h13e00001;
      80017: inst = 32'hfe0d96a;
      80018: inst = 32'h5be00000;
      80019: inst = 32'h8c50000;
      80020: inst = 32'h24612800;
      80021: inst = 32'h10a00000;
      80022: inst = 32'hca00001;
      80023: inst = 32'h24822800;
      80024: inst = 32'h10a00000;
      80025: inst = 32'hca00004;
      80026: inst = 32'h38632800;
      80027: inst = 32'h38842800;
      80028: inst = 32'h10a00001;
      80029: inst = 32'hca038a1;
      80030: inst = 32'h13e00001;
      80031: inst = 32'hfe0d96a;
      80032: inst = 32'h5be00000;
      80033: inst = 32'h8c50000;
      80034: inst = 32'h24612800;
      80035: inst = 32'h10a00000;
      80036: inst = 32'hca00001;
      80037: inst = 32'h24822800;
      80038: inst = 32'h10a00000;
      80039: inst = 32'hca00004;
      80040: inst = 32'h38632800;
      80041: inst = 32'h38842800;
      80042: inst = 32'h10a00001;
      80043: inst = 32'hca038af;
      80044: inst = 32'h13e00001;
      80045: inst = 32'hfe0d96a;
      80046: inst = 32'h5be00000;
      80047: inst = 32'h8c50000;
      80048: inst = 32'h24612800;
      80049: inst = 32'h10a00000;
      80050: inst = 32'hca00001;
      80051: inst = 32'h24822800;
      80052: inst = 32'h10a00000;
      80053: inst = 32'hca00004;
      80054: inst = 32'h38632800;
      80055: inst = 32'h38842800;
      80056: inst = 32'h10a00001;
      80057: inst = 32'hca038bd;
      80058: inst = 32'h13e00001;
      80059: inst = 32'hfe0d96a;
      80060: inst = 32'h5be00000;
      80061: inst = 32'h8c50000;
      80062: inst = 32'h24612800;
      80063: inst = 32'h10a00000;
      80064: inst = 32'hca00001;
      80065: inst = 32'h24822800;
      80066: inst = 32'h10a00000;
      80067: inst = 32'hca00004;
      80068: inst = 32'h38632800;
      80069: inst = 32'h38842800;
      80070: inst = 32'h10a00001;
      80071: inst = 32'hca038cb;
      80072: inst = 32'h13e00001;
      80073: inst = 32'hfe0d96a;
      80074: inst = 32'h5be00000;
      80075: inst = 32'h8c50000;
      80076: inst = 32'h24612800;
      80077: inst = 32'h10a00000;
      80078: inst = 32'hca00001;
      80079: inst = 32'h24822800;
      80080: inst = 32'h10a00000;
      80081: inst = 32'hca00004;
      80082: inst = 32'h38632800;
      80083: inst = 32'h38842800;
      80084: inst = 32'h10a00001;
      80085: inst = 32'hca038d9;
      80086: inst = 32'h13e00001;
      80087: inst = 32'hfe0d96a;
      80088: inst = 32'h5be00000;
      80089: inst = 32'h8c50000;
      80090: inst = 32'h24612800;
      80091: inst = 32'h10a00000;
      80092: inst = 32'hca00001;
      80093: inst = 32'h24822800;
      80094: inst = 32'h10a00000;
      80095: inst = 32'hca00004;
      80096: inst = 32'h38632800;
      80097: inst = 32'h38842800;
      80098: inst = 32'h10a00001;
      80099: inst = 32'hca038e7;
      80100: inst = 32'h13e00001;
      80101: inst = 32'hfe0d96a;
      80102: inst = 32'h5be00000;
      80103: inst = 32'h8c50000;
      80104: inst = 32'h24612800;
      80105: inst = 32'h10a00000;
      80106: inst = 32'hca00001;
      80107: inst = 32'h24822800;
      80108: inst = 32'h10a00000;
      80109: inst = 32'hca00004;
      80110: inst = 32'h38632800;
      80111: inst = 32'h38842800;
      80112: inst = 32'h10a00001;
      80113: inst = 32'hca038f5;
      80114: inst = 32'h13e00001;
      80115: inst = 32'hfe0d96a;
      80116: inst = 32'h5be00000;
      80117: inst = 32'h8c50000;
      80118: inst = 32'h24612800;
      80119: inst = 32'h10a00000;
      80120: inst = 32'hca00001;
      80121: inst = 32'h24822800;
      80122: inst = 32'h10a00000;
      80123: inst = 32'hca00004;
      80124: inst = 32'h38632800;
      80125: inst = 32'h38842800;
      80126: inst = 32'h10a00001;
      80127: inst = 32'hca03903;
      80128: inst = 32'h13e00001;
      80129: inst = 32'hfe0d96a;
      80130: inst = 32'h5be00000;
      80131: inst = 32'h8c50000;
      80132: inst = 32'h24612800;
      80133: inst = 32'h10a00000;
      80134: inst = 32'hca00001;
      80135: inst = 32'h24822800;
      80136: inst = 32'h10a00000;
      80137: inst = 32'hca00004;
      80138: inst = 32'h38632800;
      80139: inst = 32'h38842800;
      80140: inst = 32'h10a00001;
      80141: inst = 32'hca03911;
      80142: inst = 32'h13e00001;
      80143: inst = 32'hfe0d96a;
      80144: inst = 32'h5be00000;
      80145: inst = 32'h8c50000;
      80146: inst = 32'h24612800;
      80147: inst = 32'h10a00000;
      80148: inst = 32'hca00001;
      80149: inst = 32'h24822800;
      80150: inst = 32'h10a00000;
      80151: inst = 32'hca00004;
      80152: inst = 32'h38632800;
      80153: inst = 32'h38842800;
      80154: inst = 32'h10a00001;
      80155: inst = 32'hca0391f;
      80156: inst = 32'h13e00001;
      80157: inst = 32'hfe0d96a;
      80158: inst = 32'h5be00000;
      80159: inst = 32'h8c50000;
      80160: inst = 32'h24612800;
      80161: inst = 32'h10a00000;
      80162: inst = 32'hca00001;
      80163: inst = 32'h24822800;
      80164: inst = 32'h10a00000;
      80165: inst = 32'hca00004;
      80166: inst = 32'h38632800;
      80167: inst = 32'h38842800;
      80168: inst = 32'h10a00001;
      80169: inst = 32'hca0392d;
      80170: inst = 32'h13e00001;
      80171: inst = 32'hfe0d96a;
      80172: inst = 32'h5be00000;
      80173: inst = 32'h8c50000;
      80174: inst = 32'h24612800;
      80175: inst = 32'h10a00000;
      80176: inst = 32'hca00001;
      80177: inst = 32'h24822800;
      80178: inst = 32'h10a00000;
      80179: inst = 32'hca00004;
      80180: inst = 32'h38632800;
      80181: inst = 32'h38842800;
      80182: inst = 32'h10a00001;
      80183: inst = 32'hca0393b;
      80184: inst = 32'h13e00001;
      80185: inst = 32'hfe0d96a;
      80186: inst = 32'h5be00000;
      80187: inst = 32'h8c50000;
      80188: inst = 32'h24612800;
      80189: inst = 32'h10a00000;
      80190: inst = 32'hca00001;
      80191: inst = 32'h24822800;
      80192: inst = 32'h10a00000;
      80193: inst = 32'hca00004;
      80194: inst = 32'h38632800;
      80195: inst = 32'h38842800;
      80196: inst = 32'h10a00001;
      80197: inst = 32'hca03949;
      80198: inst = 32'h13e00001;
      80199: inst = 32'hfe0d96a;
      80200: inst = 32'h5be00000;
      80201: inst = 32'h8c50000;
      80202: inst = 32'h24612800;
      80203: inst = 32'h10a00000;
      80204: inst = 32'hca00001;
      80205: inst = 32'h24822800;
      80206: inst = 32'h10a00000;
      80207: inst = 32'hca00004;
      80208: inst = 32'h38632800;
      80209: inst = 32'h38842800;
      80210: inst = 32'h10a00001;
      80211: inst = 32'hca03957;
      80212: inst = 32'h13e00001;
      80213: inst = 32'hfe0d96a;
      80214: inst = 32'h5be00000;
      80215: inst = 32'h8c50000;
      80216: inst = 32'h24612800;
      80217: inst = 32'h10a00000;
      80218: inst = 32'hca00001;
      80219: inst = 32'h24822800;
      80220: inst = 32'h10a00000;
      80221: inst = 32'hca00004;
      80222: inst = 32'h38632800;
      80223: inst = 32'h38842800;
      80224: inst = 32'h10a00001;
      80225: inst = 32'hca03965;
      80226: inst = 32'h13e00001;
      80227: inst = 32'hfe0d96a;
      80228: inst = 32'h5be00000;
      80229: inst = 32'h8c50000;
      80230: inst = 32'h24612800;
      80231: inst = 32'h10a00000;
      80232: inst = 32'hca00001;
      80233: inst = 32'h24822800;
      80234: inst = 32'h10a00000;
      80235: inst = 32'hca00004;
      80236: inst = 32'h38632800;
      80237: inst = 32'h38842800;
      80238: inst = 32'h10a00001;
      80239: inst = 32'hca03973;
      80240: inst = 32'h13e00001;
      80241: inst = 32'hfe0d96a;
      80242: inst = 32'h5be00000;
      80243: inst = 32'h8c50000;
      80244: inst = 32'h24612800;
      80245: inst = 32'h10a00000;
      80246: inst = 32'hca00001;
      80247: inst = 32'h24822800;
      80248: inst = 32'h10a00000;
      80249: inst = 32'hca00004;
      80250: inst = 32'h38632800;
      80251: inst = 32'h38842800;
      80252: inst = 32'h10a00001;
      80253: inst = 32'hca03981;
      80254: inst = 32'h13e00001;
      80255: inst = 32'hfe0d96a;
      80256: inst = 32'h5be00000;
      80257: inst = 32'h8c50000;
      80258: inst = 32'h24612800;
      80259: inst = 32'h10a00000;
      80260: inst = 32'hca00001;
      80261: inst = 32'h24822800;
      80262: inst = 32'h10a00000;
      80263: inst = 32'hca00004;
      80264: inst = 32'h38632800;
      80265: inst = 32'h38842800;
      80266: inst = 32'h10a00001;
      80267: inst = 32'hca0398f;
      80268: inst = 32'h13e00001;
      80269: inst = 32'hfe0d96a;
      80270: inst = 32'h5be00000;
      80271: inst = 32'h8c50000;
      80272: inst = 32'h24612800;
      80273: inst = 32'h10a00000;
      80274: inst = 32'hca00001;
      80275: inst = 32'h24822800;
      80276: inst = 32'h10a00000;
      80277: inst = 32'hca00004;
      80278: inst = 32'h38632800;
      80279: inst = 32'h38842800;
      80280: inst = 32'h10a00001;
      80281: inst = 32'hca0399d;
      80282: inst = 32'h13e00001;
      80283: inst = 32'hfe0d96a;
      80284: inst = 32'h5be00000;
      80285: inst = 32'h8c50000;
      80286: inst = 32'h24612800;
      80287: inst = 32'h10a00000;
      80288: inst = 32'hca00001;
      80289: inst = 32'h24822800;
      80290: inst = 32'h10a00000;
      80291: inst = 32'hca00004;
      80292: inst = 32'h38632800;
      80293: inst = 32'h38842800;
      80294: inst = 32'h10a00001;
      80295: inst = 32'hca039ab;
      80296: inst = 32'h13e00001;
      80297: inst = 32'hfe0d96a;
      80298: inst = 32'h5be00000;
      80299: inst = 32'h8c50000;
      80300: inst = 32'h24612800;
      80301: inst = 32'h10a00000;
      80302: inst = 32'hca00001;
      80303: inst = 32'h24822800;
      80304: inst = 32'h10a00000;
      80305: inst = 32'hca00004;
      80306: inst = 32'h38632800;
      80307: inst = 32'h38842800;
      80308: inst = 32'h10a00001;
      80309: inst = 32'hca039b9;
      80310: inst = 32'h13e00001;
      80311: inst = 32'hfe0d96a;
      80312: inst = 32'h5be00000;
      80313: inst = 32'h8c50000;
      80314: inst = 32'h24612800;
      80315: inst = 32'h10a00000;
      80316: inst = 32'hca00001;
      80317: inst = 32'h24822800;
      80318: inst = 32'h10a00000;
      80319: inst = 32'hca00004;
      80320: inst = 32'h38632800;
      80321: inst = 32'h38842800;
      80322: inst = 32'h10a00001;
      80323: inst = 32'hca039c7;
      80324: inst = 32'h13e00001;
      80325: inst = 32'hfe0d96a;
      80326: inst = 32'h5be00000;
      80327: inst = 32'h8c50000;
      80328: inst = 32'h24612800;
      80329: inst = 32'h10a00000;
      80330: inst = 32'hca00001;
      80331: inst = 32'h24822800;
      80332: inst = 32'h10a00000;
      80333: inst = 32'hca00004;
      80334: inst = 32'h38632800;
      80335: inst = 32'h38842800;
      80336: inst = 32'h10a00001;
      80337: inst = 32'hca039d5;
      80338: inst = 32'h13e00001;
      80339: inst = 32'hfe0d96a;
      80340: inst = 32'h5be00000;
      80341: inst = 32'h8c50000;
      80342: inst = 32'h24612800;
      80343: inst = 32'h10a00000;
      80344: inst = 32'hca00001;
      80345: inst = 32'h24822800;
      80346: inst = 32'h10a00000;
      80347: inst = 32'hca00004;
      80348: inst = 32'h38632800;
      80349: inst = 32'h38842800;
      80350: inst = 32'h10a00001;
      80351: inst = 32'hca039e3;
      80352: inst = 32'h13e00001;
      80353: inst = 32'hfe0d96a;
      80354: inst = 32'h5be00000;
      80355: inst = 32'h8c50000;
      80356: inst = 32'h24612800;
      80357: inst = 32'h10a00000;
      80358: inst = 32'hca00001;
      80359: inst = 32'h24822800;
      80360: inst = 32'h10a00000;
      80361: inst = 32'hca00004;
      80362: inst = 32'h38632800;
      80363: inst = 32'h38842800;
      80364: inst = 32'h10a00001;
      80365: inst = 32'hca039f1;
      80366: inst = 32'h13e00001;
      80367: inst = 32'hfe0d96a;
      80368: inst = 32'h5be00000;
      80369: inst = 32'h8c50000;
      80370: inst = 32'h24612800;
      80371: inst = 32'h10a00000;
      80372: inst = 32'hca00001;
      80373: inst = 32'h24822800;
      80374: inst = 32'h10a00000;
      80375: inst = 32'hca00004;
      80376: inst = 32'h38632800;
      80377: inst = 32'h38842800;
      80378: inst = 32'h10a00001;
      80379: inst = 32'hca039ff;
      80380: inst = 32'h13e00001;
      80381: inst = 32'hfe0d96a;
      80382: inst = 32'h5be00000;
      80383: inst = 32'h8c50000;
      80384: inst = 32'h24612800;
      80385: inst = 32'h10a00000;
      80386: inst = 32'hca00001;
      80387: inst = 32'h24822800;
      80388: inst = 32'h10a00000;
      80389: inst = 32'hca00004;
      80390: inst = 32'h38632800;
      80391: inst = 32'h38842800;
      80392: inst = 32'h10a00001;
      80393: inst = 32'hca03a0d;
      80394: inst = 32'h13e00001;
      80395: inst = 32'hfe0d96a;
      80396: inst = 32'h5be00000;
      80397: inst = 32'h8c50000;
      80398: inst = 32'h24612800;
      80399: inst = 32'h10a00000;
      80400: inst = 32'hca00001;
      80401: inst = 32'h24822800;
      80402: inst = 32'h10a00000;
      80403: inst = 32'hca00004;
      80404: inst = 32'h38632800;
      80405: inst = 32'h38842800;
      80406: inst = 32'h10a00001;
      80407: inst = 32'hca03a1b;
      80408: inst = 32'h13e00001;
      80409: inst = 32'hfe0d96a;
      80410: inst = 32'h5be00000;
      80411: inst = 32'h8c50000;
      80412: inst = 32'h24612800;
      80413: inst = 32'h10a00000;
      80414: inst = 32'hca00001;
      80415: inst = 32'h24822800;
      80416: inst = 32'h10a00000;
      80417: inst = 32'hca00004;
      80418: inst = 32'h38632800;
      80419: inst = 32'h38842800;
      80420: inst = 32'h10a00001;
      80421: inst = 32'hca03a29;
      80422: inst = 32'h13e00001;
      80423: inst = 32'hfe0d96a;
      80424: inst = 32'h5be00000;
      80425: inst = 32'h8c50000;
      80426: inst = 32'h24612800;
      80427: inst = 32'h10a00000;
      80428: inst = 32'hca00001;
      80429: inst = 32'h24822800;
      80430: inst = 32'h10a00000;
      80431: inst = 32'hca00004;
      80432: inst = 32'h38632800;
      80433: inst = 32'h38842800;
      80434: inst = 32'h10a00001;
      80435: inst = 32'hca03a37;
      80436: inst = 32'h13e00001;
      80437: inst = 32'hfe0d96a;
      80438: inst = 32'h5be00000;
      80439: inst = 32'h8c50000;
      80440: inst = 32'h24612800;
      80441: inst = 32'h10a00000;
      80442: inst = 32'hca00001;
      80443: inst = 32'h24822800;
      80444: inst = 32'h10a00000;
      80445: inst = 32'hca00004;
      80446: inst = 32'h38632800;
      80447: inst = 32'h38842800;
      80448: inst = 32'h10a00001;
      80449: inst = 32'hca03a45;
      80450: inst = 32'h13e00001;
      80451: inst = 32'hfe0d96a;
      80452: inst = 32'h5be00000;
      80453: inst = 32'h8c50000;
      80454: inst = 32'h24612800;
      80455: inst = 32'h10a00000;
      80456: inst = 32'hca00001;
      80457: inst = 32'h24822800;
      80458: inst = 32'h10a00000;
      80459: inst = 32'hca00004;
      80460: inst = 32'h38632800;
      80461: inst = 32'h38842800;
      80462: inst = 32'h10a00001;
      80463: inst = 32'hca03a53;
      80464: inst = 32'h13e00001;
      80465: inst = 32'hfe0d96a;
      80466: inst = 32'h5be00000;
      80467: inst = 32'h8c50000;
      80468: inst = 32'h24612800;
      80469: inst = 32'h10a00000;
      80470: inst = 32'hca00001;
      80471: inst = 32'h24822800;
      80472: inst = 32'h10a00000;
      80473: inst = 32'hca00004;
      80474: inst = 32'h38632800;
      80475: inst = 32'h38842800;
      80476: inst = 32'h10a00001;
      80477: inst = 32'hca03a61;
      80478: inst = 32'h13e00001;
      80479: inst = 32'hfe0d96a;
      80480: inst = 32'h5be00000;
      80481: inst = 32'h8c50000;
      80482: inst = 32'h24612800;
      80483: inst = 32'h10a00000;
      80484: inst = 32'hca00001;
      80485: inst = 32'h24822800;
      80486: inst = 32'h10a00000;
      80487: inst = 32'hca00004;
      80488: inst = 32'h38632800;
      80489: inst = 32'h38842800;
      80490: inst = 32'h10a00001;
      80491: inst = 32'hca03a6f;
      80492: inst = 32'h13e00001;
      80493: inst = 32'hfe0d96a;
      80494: inst = 32'h5be00000;
      80495: inst = 32'h8c50000;
      80496: inst = 32'h24612800;
      80497: inst = 32'h10a00000;
      80498: inst = 32'hca00001;
      80499: inst = 32'h24822800;
      80500: inst = 32'h10a00000;
      80501: inst = 32'hca00004;
      80502: inst = 32'h38632800;
      80503: inst = 32'h38842800;
      80504: inst = 32'h10a00001;
      80505: inst = 32'hca03a7d;
      80506: inst = 32'h13e00001;
      80507: inst = 32'hfe0d96a;
      80508: inst = 32'h5be00000;
      80509: inst = 32'h8c50000;
      80510: inst = 32'h24612800;
      80511: inst = 32'h10a00000;
      80512: inst = 32'hca00001;
      80513: inst = 32'h24822800;
      80514: inst = 32'h10a00000;
      80515: inst = 32'hca00004;
      80516: inst = 32'h38632800;
      80517: inst = 32'h38842800;
      80518: inst = 32'h10a00001;
      80519: inst = 32'hca03a8b;
      80520: inst = 32'h13e00001;
      80521: inst = 32'hfe0d96a;
      80522: inst = 32'h5be00000;
      80523: inst = 32'h8c50000;
      80524: inst = 32'h24612800;
      80525: inst = 32'h10a00000;
      80526: inst = 32'hca00001;
      80527: inst = 32'h24822800;
      80528: inst = 32'h10a00000;
      80529: inst = 32'hca00004;
      80530: inst = 32'h38632800;
      80531: inst = 32'h38842800;
      80532: inst = 32'h10a00001;
      80533: inst = 32'hca03a99;
      80534: inst = 32'h13e00001;
      80535: inst = 32'hfe0d96a;
      80536: inst = 32'h5be00000;
      80537: inst = 32'h8c50000;
      80538: inst = 32'h24612800;
      80539: inst = 32'h10a00000;
      80540: inst = 32'hca00001;
      80541: inst = 32'h24822800;
      80542: inst = 32'h10a00000;
      80543: inst = 32'hca00004;
      80544: inst = 32'h38632800;
      80545: inst = 32'h38842800;
      80546: inst = 32'h10a00001;
      80547: inst = 32'hca03aa7;
      80548: inst = 32'h13e00001;
      80549: inst = 32'hfe0d96a;
      80550: inst = 32'h5be00000;
      80551: inst = 32'h8c50000;
      80552: inst = 32'h24612800;
      80553: inst = 32'h10a00000;
      80554: inst = 32'hca00001;
      80555: inst = 32'h24822800;
      80556: inst = 32'h10a00000;
      80557: inst = 32'hca00004;
      80558: inst = 32'h38632800;
      80559: inst = 32'h38842800;
      80560: inst = 32'h10a00001;
      80561: inst = 32'hca03ab5;
      80562: inst = 32'h13e00001;
      80563: inst = 32'hfe0d96a;
      80564: inst = 32'h5be00000;
      80565: inst = 32'h8c50000;
      80566: inst = 32'h24612800;
      80567: inst = 32'h10a00000;
      80568: inst = 32'hca00001;
      80569: inst = 32'h24822800;
      80570: inst = 32'h10a00000;
      80571: inst = 32'hca00004;
      80572: inst = 32'h38632800;
      80573: inst = 32'h38842800;
      80574: inst = 32'h10a00001;
      80575: inst = 32'hca03ac3;
      80576: inst = 32'h13e00001;
      80577: inst = 32'hfe0d96a;
      80578: inst = 32'h5be00000;
      80579: inst = 32'h8c50000;
      80580: inst = 32'h24612800;
      80581: inst = 32'h10a00000;
      80582: inst = 32'hca00001;
      80583: inst = 32'h24822800;
      80584: inst = 32'h10a00000;
      80585: inst = 32'hca00004;
      80586: inst = 32'h38632800;
      80587: inst = 32'h38842800;
      80588: inst = 32'h10a00001;
      80589: inst = 32'hca03ad1;
      80590: inst = 32'h13e00001;
      80591: inst = 32'hfe0d96a;
      80592: inst = 32'h5be00000;
      80593: inst = 32'h8c50000;
      80594: inst = 32'h24612800;
      80595: inst = 32'h10a00000;
      80596: inst = 32'hca00001;
      80597: inst = 32'h24822800;
      80598: inst = 32'h10a00000;
      80599: inst = 32'hca00004;
      80600: inst = 32'h38632800;
      80601: inst = 32'h38842800;
      80602: inst = 32'h10a00001;
      80603: inst = 32'hca03adf;
      80604: inst = 32'h13e00001;
      80605: inst = 32'hfe0d96a;
      80606: inst = 32'h5be00000;
      80607: inst = 32'h8c50000;
      80608: inst = 32'h24612800;
      80609: inst = 32'h10a00000;
      80610: inst = 32'hca00001;
      80611: inst = 32'h24822800;
      80612: inst = 32'h10a00000;
      80613: inst = 32'hca00004;
      80614: inst = 32'h38632800;
      80615: inst = 32'h38842800;
      80616: inst = 32'h10a00001;
      80617: inst = 32'hca03aed;
      80618: inst = 32'h13e00001;
      80619: inst = 32'hfe0d96a;
      80620: inst = 32'h5be00000;
      80621: inst = 32'h8c50000;
      80622: inst = 32'h24612800;
      80623: inst = 32'h10a00000;
      80624: inst = 32'hca00001;
      80625: inst = 32'h24822800;
      80626: inst = 32'h10a00000;
      80627: inst = 32'hca00004;
      80628: inst = 32'h38632800;
      80629: inst = 32'h38842800;
      80630: inst = 32'h10a00001;
      80631: inst = 32'hca03afb;
      80632: inst = 32'h13e00001;
      80633: inst = 32'hfe0d96a;
      80634: inst = 32'h5be00000;
      80635: inst = 32'h8c50000;
      80636: inst = 32'h24612800;
      80637: inst = 32'h10a00000;
      80638: inst = 32'hca00001;
      80639: inst = 32'h24822800;
      80640: inst = 32'h10a00000;
      80641: inst = 32'hca00004;
      80642: inst = 32'h38632800;
      80643: inst = 32'h38842800;
      80644: inst = 32'h10a00001;
      80645: inst = 32'hca03b09;
      80646: inst = 32'h13e00001;
      80647: inst = 32'hfe0d96a;
      80648: inst = 32'h5be00000;
      80649: inst = 32'h8c50000;
      80650: inst = 32'h24612800;
      80651: inst = 32'h10a00000;
      80652: inst = 32'hca00001;
      80653: inst = 32'h24822800;
      80654: inst = 32'h10a00000;
      80655: inst = 32'hca00004;
      80656: inst = 32'h38632800;
      80657: inst = 32'h38842800;
      80658: inst = 32'h10a00001;
      80659: inst = 32'hca03b17;
      80660: inst = 32'h13e00001;
      80661: inst = 32'hfe0d96a;
      80662: inst = 32'h5be00000;
      80663: inst = 32'h8c50000;
      80664: inst = 32'h24612800;
      80665: inst = 32'h10a00000;
      80666: inst = 32'hca00001;
      80667: inst = 32'h24822800;
      80668: inst = 32'h10a00000;
      80669: inst = 32'hca00004;
      80670: inst = 32'h38632800;
      80671: inst = 32'h38842800;
      80672: inst = 32'h10a00001;
      80673: inst = 32'hca03b25;
      80674: inst = 32'h13e00001;
      80675: inst = 32'hfe0d96a;
      80676: inst = 32'h5be00000;
      80677: inst = 32'h8c50000;
      80678: inst = 32'h24612800;
      80679: inst = 32'h10a00000;
      80680: inst = 32'hca00001;
      80681: inst = 32'h24822800;
      80682: inst = 32'h10a00000;
      80683: inst = 32'hca00004;
      80684: inst = 32'h38632800;
      80685: inst = 32'h38842800;
      80686: inst = 32'h10a00001;
      80687: inst = 32'hca03b33;
      80688: inst = 32'h13e00001;
      80689: inst = 32'hfe0d96a;
      80690: inst = 32'h5be00000;
      80691: inst = 32'h8c50000;
      80692: inst = 32'h24612800;
      80693: inst = 32'h10a00000;
      80694: inst = 32'hca00001;
      80695: inst = 32'h24822800;
      80696: inst = 32'h10a00000;
      80697: inst = 32'hca00004;
      80698: inst = 32'h38632800;
      80699: inst = 32'h38842800;
      80700: inst = 32'h10a00001;
      80701: inst = 32'hca03b41;
      80702: inst = 32'h13e00001;
      80703: inst = 32'hfe0d96a;
      80704: inst = 32'h5be00000;
      80705: inst = 32'h8c50000;
      80706: inst = 32'h24612800;
      80707: inst = 32'h10a00000;
      80708: inst = 32'hca00001;
      80709: inst = 32'h24822800;
      80710: inst = 32'h10a00000;
      80711: inst = 32'hca00004;
      80712: inst = 32'h38632800;
      80713: inst = 32'h38842800;
      80714: inst = 32'h10a00001;
      80715: inst = 32'hca03b4f;
      80716: inst = 32'h13e00001;
      80717: inst = 32'hfe0d96a;
      80718: inst = 32'h5be00000;
      80719: inst = 32'h8c50000;
      80720: inst = 32'h24612800;
      80721: inst = 32'h10a00000;
      80722: inst = 32'hca00001;
      80723: inst = 32'h24822800;
      80724: inst = 32'h10a00000;
      80725: inst = 32'hca00004;
      80726: inst = 32'h38632800;
      80727: inst = 32'h38842800;
      80728: inst = 32'h10a00001;
      80729: inst = 32'hca03b5d;
      80730: inst = 32'h13e00001;
      80731: inst = 32'hfe0d96a;
      80732: inst = 32'h5be00000;
      80733: inst = 32'h8c50000;
      80734: inst = 32'h24612800;
      80735: inst = 32'h10a00000;
      80736: inst = 32'hca00001;
      80737: inst = 32'h24822800;
      80738: inst = 32'h10a00000;
      80739: inst = 32'hca00004;
      80740: inst = 32'h38632800;
      80741: inst = 32'h38842800;
      80742: inst = 32'h10a00001;
      80743: inst = 32'hca03b6b;
      80744: inst = 32'h13e00001;
      80745: inst = 32'hfe0d96a;
      80746: inst = 32'h5be00000;
      80747: inst = 32'h8c50000;
      80748: inst = 32'h24612800;
      80749: inst = 32'h10a00000;
      80750: inst = 32'hca00001;
      80751: inst = 32'h24822800;
      80752: inst = 32'h10a00000;
      80753: inst = 32'hca00004;
      80754: inst = 32'h38632800;
      80755: inst = 32'h38842800;
      80756: inst = 32'h10a00001;
      80757: inst = 32'hca03b79;
      80758: inst = 32'h13e00001;
      80759: inst = 32'hfe0d96a;
      80760: inst = 32'h5be00000;
      80761: inst = 32'h8c50000;
      80762: inst = 32'h24612800;
      80763: inst = 32'h10a00000;
      80764: inst = 32'hca00001;
      80765: inst = 32'h24822800;
      80766: inst = 32'h10a00000;
      80767: inst = 32'hca00004;
      80768: inst = 32'h38632800;
      80769: inst = 32'h38842800;
      80770: inst = 32'h10a00001;
      80771: inst = 32'hca03b87;
      80772: inst = 32'h13e00001;
      80773: inst = 32'hfe0d96a;
      80774: inst = 32'h5be00000;
      80775: inst = 32'h8c50000;
      80776: inst = 32'h24612800;
      80777: inst = 32'h10a00000;
      80778: inst = 32'hca00001;
      80779: inst = 32'h24822800;
      80780: inst = 32'h10a00000;
      80781: inst = 32'hca00004;
      80782: inst = 32'h38632800;
      80783: inst = 32'h38842800;
      80784: inst = 32'h10a00001;
      80785: inst = 32'hca03b95;
      80786: inst = 32'h13e00001;
      80787: inst = 32'hfe0d96a;
      80788: inst = 32'h5be00000;
      80789: inst = 32'h8c50000;
      80790: inst = 32'h24612800;
      80791: inst = 32'h10a00000;
      80792: inst = 32'hca00001;
      80793: inst = 32'h24822800;
      80794: inst = 32'h10a00000;
      80795: inst = 32'hca00004;
      80796: inst = 32'h38632800;
      80797: inst = 32'h38842800;
      80798: inst = 32'h10a00001;
      80799: inst = 32'hca03ba3;
      80800: inst = 32'h13e00001;
      80801: inst = 32'hfe0d96a;
      80802: inst = 32'h5be00000;
      80803: inst = 32'h8c50000;
      80804: inst = 32'h24612800;
      80805: inst = 32'h10a00000;
      80806: inst = 32'hca00001;
      80807: inst = 32'h24822800;
      80808: inst = 32'h10a00000;
      80809: inst = 32'hca00004;
      80810: inst = 32'h38632800;
      80811: inst = 32'h38842800;
      80812: inst = 32'h10a00001;
      80813: inst = 32'hca03bb1;
      80814: inst = 32'h13e00001;
      80815: inst = 32'hfe0d96a;
      80816: inst = 32'h5be00000;
      80817: inst = 32'h8c50000;
      80818: inst = 32'h24612800;
      80819: inst = 32'h10a00000;
      80820: inst = 32'hca00001;
      80821: inst = 32'h24822800;
      80822: inst = 32'h10a00000;
      80823: inst = 32'hca00004;
      80824: inst = 32'h38632800;
      80825: inst = 32'h38842800;
      80826: inst = 32'h10a00001;
      80827: inst = 32'hca03bbf;
      80828: inst = 32'h13e00001;
      80829: inst = 32'hfe0d96a;
      80830: inst = 32'h5be00000;
      80831: inst = 32'h8c50000;
      80832: inst = 32'h24612800;
      80833: inst = 32'h10a00000;
      80834: inst = 32'hca00001;
      80835: inst = 32'h24822800;
      80836: inst = 32'h10a00000;
      80837: inst = 32'hca00004;
      80838: inst = 32'h38632800;
      80839: inst = 32'h38842800;
      80840: inst = 32'h10a00001;
      80841: inst = 32'hca03bcd;
      80842: inst = 32'h13e00001;
      80843: inst = 32'hfe0d96a;
      80844: inst = 32'h5be00000;
      80845: inst = 32'h8c50000;
      80846: inst = 32'h24612800;
      80847: inst = 32'h10a00000;
      80848: inst = 32'hca00001;
      80849: inst = 32'h24822800;
      80850: inst = 32'h10a00000;
      80851: inst = 32'hca00004;
      80852: inst = 32'h38632800;
      80853: inst = 32'h38842800;
      80854: inst = 32'h10a00001;
      80855: inst = 32'hca03bdb;
      80856: inst = 32'h13e00001;
      80857: inst = 32'hfe0d96a;
      80858: inst = 32'h5be00000;
      80859: inst = 32'h8c50000;
      80860: inst = 32'h24612800;
      80861: inst = 32'h10a00000;
      80862: inst = 32'hca00001;
      80863: inst = 32'h24822800;
      80864: inst = 32'h10a00000;
      80865: inst = 32'hca00004;
      80866: inst = 32'h38632800;
      80867: inst = 32'h38842800;
      80868: inst = 32'h10a00001;
      80869: inst = 32'hca03be9;
      80870: inst = 32'h13e00001;
      80871: inst = 32'hfe0d96a;
      80872: inst = 32'h5be00000;
      80873: inst = 32'h8c50000;
      80874: inst = 32'h24612800;
      80875: inst = 32'h10a00000;
      80876: inst = 32'hca00002;
      80877: inst = 32'h24822800;
      80878: inst = 32'h10a00000;
      80879: inst = 32'hca00004;
      80880: inst = 32'h38632800;
      80881: inst = 32'h38842800;
      80882: inst = 32'h10a00001;
      80883: inst = 32'hca03bf7;
      80884: inst = 32'h13e00001;
      80885: inst = 32'hfe0d96a;
      80886: inst = 32'h5be00000;
      80887: inst = 32'h8c50000;
      80888: inst = 32'h24612800;
      80889: inst = 32'h10a00000;
      80890: inst = 32'hca00002;
      80891: inst = 32'h24822800;
      80892: inst = 32'h10a00000;
      80893: inst = 32'hca00004;
      80894: inst = 32'h38632800;
      80895: inst = 32'h38842800;
      80896: inst = 32'h10a00001;
      80897: inst = 32'hca03c05;
      80898: inst = 32'h13e00001;
      80899: inst = 32'hfe0d96a;
      80900: inst = 32'h5be00000;
      80901: inst = 32'h8c50000;
      80902: inst = 32'h24612800;
      80903: inst = 32'h10a00000;
      80904: inst = 32'hca00002;
      80905: inst = 32'h24822800;
      80906: inst = 32'h10a00000;
      80907: inst = 32'hca00004;
      80908: inst = 32'h38632800;
      80909: inst = 32'h38842800;
      80910: inst = 32'h10a00001;
      80911: inst = 32'hca03c13;
      80912: inst = 32'h13e00001;
      80913: inst = 32'hfe0d96a;
      80914: inst = 32'h5be00000;
      80915: inst = 32'h8c50000;
      80916: inst = 32'h24612800;
      80917: inst = 32'h10a00000;
      80918: inst = 32'hca00002;
      80919: inst = 32'h24822800;
      80920: inst = 32'h10a00000;
      80921: inst = 32'hca00004;
      80922: inst = 32'h38632800;
      80923: inst = 32'h38842800;
      80924: inst = 32'h10a00001;
      80925: inst = 32'hca03c21;
      80926: inst = 32'h13e00001;
      80927: inst = 32'hfe0d96a;
      80928: inst = 32'h5be00000;
      80929: inst = 32'h8c50000;
      80930: inst = 32'h24612800;
      80931: inst = 32'h10a00000;
      80932: inst = 32'hca00002;
      80933: inst = 32'h24822800;
      80934: inst = 32'h10a00000;
      80935: inst = 32'hca00004;
      80936: inst = 32'h38632800;
      80937: inst = 32'h38842800;
      80938: inst = 32'h10a00001;
      80939: inst = 32'hca03c2f;
      80940: inst = 32'h13e00001;
      80941: inst = 32'hfe0d96a;
      80942: inst = 32'h5be00000;
      80943: inst = 32'h8c50000;
      80944: inst = 32'h24612800;
      80945: inst = 32'h10a00000;
      80946: inst = 32'hca00002;
      80947: inst = 32'h24822800;
      80948: inst = 32'h10a00000;
      80949: inst = 32'hca00004;
      80950: inst = 32'h38632800;
      80951: inst = 32'h38842800;
      80952: inst = 32'h10a00001;
      80953: inst = 32'hca03c3d;
      80954: inst = 32'h13e00001;
      80955: inst = 32'hfe0d96a;
      80956: inst = 32'h5be00000;
      80957: inst = 32'h8c50000;
      80958: inst = 32'h24612800;
      80959: inst = 32'h10a00000;
      80960: inst = 32'hca00002;
      80961: inst = 32'h24822800;
      80962: inst = 32'h10a00000;
      80963: inst = 32'hca00004;
      80964: inst = 32'h38632800;
      80965: inst = 32'h38842800;
      80966: inst = 32'h10a00001;
      80967: inst = 32'hca03c4b;
      80968: inst = 32'h13e00001;
      80969: inst = 32'hfe0d96a;
      80970: inst = 32'h5be00000;
      80971: inst = 32'h8c50000;
      80972: inst = 32'h24612800;
      80973: inst = 32'h10a00000;
      80974: inst = 32'hca00002;
      80975: inst = 32'h24822800;
      80976: inst = 32'h10a00000;
      80977: inst = 32'hca00004;
      80978: inst = 32'h38632800;
      80979: inst = 32'h38842800;
      80980: inst = 32'h10a00001;
      80981: inst = 32'hca03c59;
      80982: inst = 32'h13e00001;
      80983: inst = 32'hfe0d96a;
      80984: inst = 32'h5be00000;
      80985: inst = 32'h8c50000;
      80986: inst = 32'h24612800;
      80987: inst = 32'h10a00000;
      80988: inst = 32'hca00002;
      80989: inst = 32'h24822800;
      80990: inst = 32'h10a00000;
      80991: inst = 32'hca00004;
      80992: inst = 32'h38632800;
      80993: inst = 32'h38842800;
      80994: inst = 32'h10a00001;
      80995: inst = 32'hca03c67;
      80996: inst = 32'h13e00001;
      80997: inst = 32'hfe0d96a;
      80998: inst = 32'h5be00000;
      80999: inst = 32'h8c50000;
      81000: inst = 32'h24612800;
      81001: inst = 32'h10a00000;
      81002: inst = 32'hca00002;
      81003: inst = 32'h24822800;
      81004: inst = 32'h10a00000;
      81005: inst = 32'hca00004;
      81006: inst = 32'h38632800;
      81007: inst = 32'h38842800;
      81008: inst = 32'h10a00001;
      81009: inst = 32'hca03c75;
      81010: inst = 32'h13e00001;
      81011: inst = 32'hfe0d96a;
      81012: inst = 32'h5be00000;
      81013: inst = 32'h8c50000;
      81014: inst = 32'h24612800;
      81015: inst = 32'h10a00000;
      81016: inst = 32'hca00002;
      81017: inst = 32'h24822800;
      81018: inst = 32'h10a00000;
      81019: inst = 32'hca00004;
      81020: inst = 32'h38632800;
      81021: inst = 32'h38842800;
      81022: inst = 32'h10a00001;
      81023: inst = 32'hca03c83;
      81024: inst = 32'h13e00001;
      81025: inst = 32'hfe0d96a;
      81026: inst = 32'h5be00000;
      81027: inst = 32'h8c50000;
      81028: inst = 32'h24612800;
      81029: inst = 32'h10a00000;
      81030: inst = 32'hca00002;
      81031: inst = 32'h24822800;
      81032: inst = 32'h10a00000;
      81033: inst = 32'hca00004;
      81034: inst = 32'h38632800;
      81035: inst = 32'h38842800;
      81036: inst = 32'h10a00001;
      81037: inst = 32'hca03c91;
      81038: inst = 32'h13e00001;
      81039: inst = 32'hfe0d96a;
      81040: inst = 32'h5be00000;
      81041: inst = 32'h8c50000;
      81042: inst = 32'h24612800;
      81043: inst = 32'h10a00000;
      81044: inst = 32'hca00002;
      81045: inst = 32'h24822800;
      81046: inst = 32'h10a00000;
      81047: inst = 32'hca00004;
      81048: inst = 32'h38632800;
      81049: inst = 32'h38842800;
      81050: inst = 32'h10a00001;
      81051: inst = 32'hca03c9f;
      81052: inst = 32'h13e00001;
      81053: inst = 32'hfe0d96a;
      81054: inst = 32'h5be00000;
      81055: inst = 32'h8c50000;
      81056: inst = 32'h24612800;
      81057: inst = 32'h10a00000;
      81058: inst = 32'hca00002;
      81059: inst = 32'h24822800;
      81060: inst = 32'h10a00000;
      81061: inst = 32'hca00004;
      81062: inst = 32'h38632800;
      81063: inst = 32'h38842800;
      81064: inst = 32'h10a00001;
      81065: inst = 32'hca03cad;
      81066: inst = 32'h13e00001;
      81067: inst = 32'hfe0d96a;
      81068: inst = 32'h5be00000;
      81069: inst = 32'h8c50000;
      81070: inst = 32'h24612800;
      81071: inst = 32'h10a00000;
      81072: inst = 32'hca00002;
      81073: inst = 32'h24822800;
      81074: inst = 32'h10a00000;
      81075: inst = 32'hca00004;
      81076: inst = 32'h38632800;
      81077: inst = 32'h38842800;
      81078: inst = 32'h10a00001;
      81079: inst = 32'hca03cbb;
      81080: inst = 32'h13e00001;
      81081: inst = 32'hfe0d96a;
      81082: inst = 32'h5be00000;
      81083: inst = 32'h8c50000;
      81084: inst = 32'h24612800;
      81085: inst = 32'h10a00000;
      81086: inst = 32'hca00002;
      81087: inst = 32'h24822800;
      81088: inst = 32'h10a00000;
      81089: inst = 32'hca00004;
      81090: inst = 32'h38632800;
      81091: inst = 32'h38842800;
      81092: inst = 32'h10a00001;
      81093: inst = 32'hca03cc9;
      81094: inst = 32'h13e00001;
      81095: inst = 32'hfe0d96a;
      81096: inst = 32'h5be00000;
      81097: inst = 32'h8c50000;
      81098: inst = 32'h24612800;
      81099: inst = 32'h10a00000;
      81100: inst = 32'hca00002;
      81101: inst = 32'h24822800;
      81102: inst = 32'h10a00000;
      81103: inst = 32'hca00004;
      81104: inst = 32'h38632800;
      81105: inst = 32'h38842800;
      81106: inst = 32'h10a00001;
      81107: inst = 32'hca03cd7;
      81108: inst = 32'h13e00001;
      81109: inst = 32'hfe0d96a;
      81110: inst = 32'h5be00000;
      81111: inst = 32'h8c50000;
      81112: inst = 32'h24612800;
      81113: inst = 32'h10a00000;
      81114: inst = 32'hca00002;
      81115: inst = 32'h24822800;
      81116: inst = 32'h10a00000;
      81117: inst = 32'hca00004;
      81118: inst = 32'h38632800;
      81119: inst = 32'h38842800;
      81120: inst = 32'h10a00001;
      81121: inst = 32'hca03ce5;
      81122: inst = 32'h13e00001;
      81123: inst = 32'hfe0d96a;
      81124: inst = 32'h5be00000;
      81125: inst = 32'h8c50000;
      81126: inst = 32'h24612800;
      81127: inst = 32'h10a00000;
      81128: inst = 32'hca00002;
      81129: inst = 32'h24822800;
      81130: inst = 32'h10a00000;
      81131: inst = 32'hca00004;
      81132: inst = 32'h38632800;
      81133: inst = 32'h38842800;
      81134: inst = 32'h10a00001;
      81135: inst = 32'hca03cf3;
      81136: inst = 32'h13e00001;
      81137: inst = 32'hfe0d96a;
      81138: inst = 32'h5be00000;
      81139: inst = 32'h8c50000;
      81140: inst = 32'h24612800;
      81141: inst = 32'h10a00000;
      81142: inst = 32'hca00002;
      81143: inst = 32'h24822800;
      81144: inst = 32'h10a00000;
      81145: inst = 32'hca00004;
      81146: inst = 32'h38632800;
      81147: inst = 32'h38842800;
      81148: inst = 32'h10a00001;
      81149: inst = 32'hca03d01;
      81150: inst = 32'h13e00001;
      81151: inst = 32'hfe0d96a;
      81152: inst = 32'h5be00000;
      81153: inst = 32'h8c50000;
      81154: inst = 32'h24612800;
      81155: inst = 32'h10a00000;
      81156: inst = 32'hca00002;
      81157: inst = 32'h24822800;
      81158: inst = 32'h10a00000;
      81159: inst = 32'hca00004;
      81160: inst = 32'h38632800;
      81161: inst = 32'h38842800;
      81162: inst = 32'h10a00001;
      81163: inst = 32'hca03d0f;
      81164: inst = 32'h13e00001;
      81165: inst = 32'hfe0d96a;
      81166: inst = 32'h5be00000;
      81167: inst = 32'h8c50000;
      81168: inst = 32'h24612800;
      81169: inst = 32'h10a00000;
      81170: inst = 32'hca00002;
      81171: inst = 32'h24822800;
      81172: inst = 32'h10a00000;
      81173: inst = 32'hca00004;
      81174: inst = 32'h38632800;
      81175: inst = 32'h38842800;
      81176: inst = 32'h10a00001;
      81177: inst = 32'hca03d1d;
      81178: inst = 32'h13e00001;
      81179: inst = 32'hfe0d96a;
      81180: inst = 32'h5be00000;
      81181: inst = 32'h8c50000;
      81182: inst = 32'h24612800;
      81183: inst = 32'h10a00000;
      81184: inst = 32'hca00002;
      81185: inst = 32'h24822800;
      81186: inst = 32'h10a00000;
      81187: inst = 32'hca00004;
      81188: inst = 32'h38632800;
      81189: inst = 32'h38842800;
      81190: inst = 32'h10a00001;
      81191: inst = 32'hca03d2b;
      81192: inst = 32'h13e00001;
      81193: inst = 32'hfe0d96a;
      81194: inst = 32'h5be00000;
      81195: inst = 32'h8c50000;
      81196: inst = 32'h24612800;
      81197: inst = 32'h10a00000;
      81198: inst = 32'hca00002;
      81199: inst = 32'h24822800;
      81200: inst = 32'h10a00000;
      81201: inst = 32'hca00004;
      81202: inst = 32'h38632800;
      81203: inst = 32'h38842800;
      81204: inst = 32'h10a00001;
      81205: inst = 32'hca03d39;
      81206: inst = 32'h13e00001;
      81207: inst = 32'hfe0d96a;
      81208: inst = 32'h5be00000;
      81209: inst = 32'h8c50000;
      81210: inst = 32'h24612800;
      81211: inst = 32'h10a00000;
      81212: inst = 32'hca00002;
      81213: inst = 32'h24822800;
      81214: inst = 32'h10a00000;
      81215: inst = 32'hca00004;
      81216: inst = 32'h38632800;
      81217: inst = 32'h38842800;
      81218: inst = 32'h10a00001;
      81219: inst = 32'hca03d47;
      81220: inst = 32'h13e00001;
      81221: inst = 32'hfe0d96a;
      81222: inst = 32'h5be00000;
      81223: inst = 32'h8c50000;
      81224: inst = 32'h24612800;
      81225: inst = 32'h10a00000;
      81226: inst = 32'hca00002;
      81227: inst = 32'h24822800;
      81228: inst = 32'h10a00000;
      81229: inst = 32'hca00004;
      81230: inst = 32'h38632800;
      81231: inst = 32'h38842800;
      81232: inst = 32'h10a00001;
      81233: inst = 32'hca03d55;
      81234: inst = 32'h13e00001;
      81235: inst = 32'hfe0d96a;
      81236: inst = 32'h5be00000;
      81237: inst = 32'h8c50000;
      81238: inst = 32'h24612800;
      81239: inst = 32'h10a00000;
      81240: inst = 32'hca00002;
      81241: inst = 32'h24822800;
      81242: inst = 32'h10a00000;
      81243: inst = 32'hca00004;
      81244: inst = 32'h38632800;
      81245: inst = 32'h38842800;
      81246: inst = 32'h10a00001;
      81247: inst = 32'hca03d63;
      81248: inst = 32'h13e00001;
      81249: inst = 32'hfe0d96a;
      81250: inst = 32'h5be00000;
      81251: inst = 32'h8c50000;
      81252: inst = 32'h24612800;
      81253: inst = 32'h10a00000;
      81254: inst = 32'hca00002;
      81255: inst = 32'h24822800;
      81256: inst = 32'h10a00000;
      81257: inst = 32'hca00004;
      81258: inst = 32'h38632800;
      81259: inst = 32'h38842800;
      81260: inst = 32'h10a00001;
      81261: inst = 32'hca03d71;
      81262: inst = 32'h13e00001;
      81263: inst = 32'hfe0d96a;
      81264: inst = 32'h5be00000;
      81265: inst = 32'h8c50000;
      81266: inst = 32'h24612800;
      81267: inst = 32'h10a00000;
      81268: inst = 32'hca00002;
      81269: inst = 32'h24822800;
      81270: inst = 32'h10a00000;
      81271: inst = 32'hca00004;
      81272: inst = 32'h38632800;
      81273: inst = 32'h38842800;
      81274: inst = 32'h10a00001;
      81275: inst = 32'hca03d7f;
      81276: inst = 32'h13e00001;
      81277: inst = 32'hfe0d96a;
      81278: inst = 32'h5be00000;
      81279: inst = 32'h8c50000;
      81280: inst = 32'h24612800;
      81281: inst = 32'h10a00000;
      81282: inst = 32'hca00002;
      81283: inst = 32'h24822800;
      81284: inst = 32'h10a00000;
      81285: inst = 32'hca00004;
      81286: inst = 32'h38632800;
      81287: inst = 32'h38842800;
      81288: inst = 32'h10a00001;
      81289: inst = 32'hca03d8d;
      81290: inst = 32'h13e00001;
      81291: inst = 32'hfe0d96a;
      81292: inst = 32'h5be00000;
      81293: inst = 32'h8c50000;
      81294: inst = 32'h24612800;
      81295: inst = 32'h10a00000;
      81296: inst = 32'hca00002;
      81297: inst = 32'h24822800;
      81298: inst = 32'h10a00000;
      81299: inst = 32'hca00004;
      81300: inst = 32'h38632800;
      81301: inst = 32'h38842800;
      81302: inst = 32'h10a00001;
      81303: inst = 32'hca03d9b;
      81304: inst = 32'h13e00001;
      81305: inst = 32'hfe0d96a;
      81306: inst = 32'h5be00000;
      81307: inst = 32'h8c50000;
      81308: inst = 32'h24612800;
      81309: inst = 32'h10a00000;
      81310: inst = 32'hca00002;
      81311: inst = 32'h24822800;
      81312: inst = 32'h10a00000;
      81313: inst = 32'hca00004;
      81314: inst = 32'h38632800;
      81315: inst = 32'h38842800;
      81316: inst = 32'h10a00001;
      81317: inst = 32'hca03da9;
      81318: inst = 32'h13e00001;
      81319: inst = 32'hfe0d96a;
      81320: inst = 32'h5be00000;
      81321: inst = 32'h8c50000;
      81322: inst = 32'h24612800;
      81323: inst = 32'h10a00000;
      81324: inst = 32'hca00002;
      81325: inst = 32'h24822800;
      81326: inst = 32'h10a00000;
      81327: inst = 32'hca00004;
      81328: inst = 32'h38632800;
      81329: inst = 32'h38842800;
      81330: inst = 32'h10a00001;
      81331: inst = 32'hca03db7;
      81332: inst = 32'h13e00001;
      81333: inst = 32'hfe0d96a;
      81334: inst = 32'h5be00000;
      81335: inst = 32'h8c50000;
      81336: inst = 32'h24612800;
      81337: inst = 32'h10a00000;
      81338: inst = 32'hca00002;
      81339: inst = 32'h24822800;
      81340: inst = 32'h10a00000;
      81341: inst = 32'hca00004;
      81342: inst = 32'h38632800;
      81343: inst = 32'h38842800;
      81344: inst = 32'h10a00001;
      81345: inst = 32'hca03dc5;
      81346: inst = 32'h13e00001;
      81347: inst = 32'hfe0d96a;
      81348: inst = 32'h5be00000;
      81349: inst = 32'h8c50000;
      81350: inst = 32'h24612800;
      81351: inst = 32'h10a00000;
      81352: inst = 32'hca00002;
      81353: inst = 32'h24822800;
      81354: inst = 32'h10a00000;
      81355: inst = 32'hca00004;
      81356: inst = 32'h38632800;
      81357: inst = 32'h38842800;
      81358: inst = 32'h10a00001;
      81359: inst = 32'hca03dd3;
      81360: inst = 32'h13e00001;
      81361: inst = 32'hfe0d96a;
      81362: inst = 32'h5be00000;
      81363: inst = 32'h8c50000;
      81364: inst = 32'h24612800;
      81365: inst = 32'h10a00000;
      81366: inst = 32'hca00002;
      81367: inst = 32'h24822800;
      81368: inst = 32'h10a00000;
      81369: inst = 32'hca00004;
      81370: inst = 32'h38632800;
      81371: inst = 32'h38842800;
      81372: inst = 32'h10a00001;
      81373: inst = 32'hca03de1;
      81374: inst = 32'h13e00001;
      81375: inst = 32'hfe0d96a;
      81376: inst = 32'h5be00000;
      81377: inst = 32'h8c50000;
      81378: inst = 32'h24612800;
      81379: inst = 32'h10a00000;
      81380: inst = 32'hca00002;
      81381: inst = 32'h24822800;
      81382: inst = 32'h10a00000;
      81383: inst = 32'hca00004;
      81384: inst = 32'h38632800;
      81385: inst = 32'h38842800;
      81386: inst = 32'h10a00001;
      81387: inst = 32'hca03def;
      81388: inst = 32'h13e00001;
      81389: inst = 32'hfe0d96a;
      81390: inst = 32'h5be00000;
      81391: inst = 32'h8c50000;
      81392: inst = 32'h24612800;
      81393: inst = 32'h10a00000;
      81394: inst = 32'hca00002;
      81395: inst = 32'h24822800;
      81396: inst = 32'h10a00000;
      81397: inst = 32'hca00004;
      81398: inst = 32'h38632800;
      81399: inst = 32'h38842800;
      81400: inst = 32'h10a00001;
      81401: inst = 32'hca03dfd;
      81402: inst = 32'h13e00001;
      81403: inst = 32'hfe0d96a;
      81404: inst = 32'h5be00000;
      81405: inst = 32'h8c50000;
      81406: inst = 32'h24612800;
      81407: inst = 32'h10a00000;
      81408: inst = 32'hca00002;
      81409: inst = 32'h24822800;
      81410: inst = 32'h10a00000;
      81411: inst = 32'hca00004;
      81412: inst = 32'h38632800;
      81413: inst = 32'h38842800;
      81414: inst = 32'h10a00001;
      81415: inst = 32'hca03e0b;
      81416: inst = 32'h13e00001;
      81417: inst = 32'hfe0d96a;
      81418: inst = 32'h5be00000;
      81419: inst = 32'h8c50000;
      81420: inst = 32'h24612800;
      81421: inst = 32'h10a00000;
      81422: inst = 32'hca00002;
      81423: inst = 32'h24822800;
      81424: inst = 32'h10a00000;
      81425: inst = 32'hca00004;
      81426: inst = 32'h38632800;
      81427: inst = 32'h38842800;
      81428: inst = 32'h10a00001;
      81429: inst = 32'hca03e19;
      81430: inst = 32'h13e00001;
      81431: inst = 32'hfe0d96a;
      81432: inst = 32'h5be00000;
      81433: inst = 32'h8c50000;
      81434: inst = 32'h24612800;
      81435: inst = 32'h10a00000;
      81436: inst = 32'hca00002;
      81437: inst = 32'h24822800;
      81438: inst = 32'h10a00000;
      81439: inst = 32'hca00004;
      81440: inst = 32'h38632800;
      81441: inst = 32'h38842800;
      81442: inst = 32'h10a00001;
      81443: inst = 32'hca03e27;
      81444: inst = 32'h13e00001;
      81445: inst = 32'hfe0d96a;
      81446: inst = 32'h5be00000;
      81447: inst = 32'h8c50000;
      81448: inst = 32'h24612800;
      81449: inst = 32'h10a00000;
      81450: inst = 32'hca00002;
      81451: inst = 32'h24822800;
      81452: inst = 32'h10a00000;
      81453: inst = 32'hca00004;
      81454: inst = 32'h38632800;
      81455: inst = 32'h38842800;
      81456: inst = 32'h10a00001;
      81457: inst = 32'hca03e35;
      81458: inst = 32'h13e00001;
      81459: inst = 32'hfe0d96a;
      81460: inst = 32'h5be00000;
      81461: inst = 32'h8c50000;
      81462: inst = 32'h24612800;
      81463: inst = 32'h10a00000;
      81464: inst = 32'hca00002;
      81465: inst = 32'h24822800;
      81466: inst = 32'h10a00000;
      81467: inst = 32'hca00004;
      81468: inst = 32'h38632800;
      81469: inst = 32'h38842800;
      81470: inst = 32'h10a00001;
      81471: inst = 32'hca03e43;
      81472: inst = 32'h13e00001;
      81473: inst = 32'hfe0d96a;
      81474: inst = 32'h5be00000;
      81475: inst = 32'h8c50000;
      81476: inst = 32'h24612800;
      81477: inst = 32'h10a00000;
      81478: inst = 32'hca00002;
      81479: inst = 32'h24822800;
      81480: inst = 32'h10a00000;
      81481: inst = 32'hca00004;
      81482: inst = 32'h38632800;
      81483: inst = 32'h38842800;
      81484: inst = 32'h10a00001;
      81485: inst = 32'hca03e51;
      81486: inst = 32'h13e00001;
      81487: inst = 32'hfe0d96a;
      81488: inst = 32'h5be00000;
      81489: inst = 32'h8c50000;
      81490: inst = 32'h24612800;
      81491: inst = 32'h10a00000;
      81492: inst = 32'hca00002;
      81493: inst = 32'h24822800;
      81494: inst = 32'h10a00000;
      81495: inst = 32'hca00004;
      81496: inst = 32'h38632800;
      81497: inst = 32'h38842800;
      81498: inst = 32'h10a00001;
      81499: inst = 32'hca03e5f;
      81500: inst = 32'h13e00001;
      81501: inst = 32'hfe0d96a;
      81502: inst = 32'h5be00000;
      81503: inst = 32'h8c50000;
      81504: inst = 32'h24612800;
      81505: inst = 32'h10a00000;
      81506: inst = 32'hca00002;
      81507: inst = 32'h24822800;
      81508: inst = 32'h10a00000;
      81509: inst = 32'hca00004;
      81510: inst = 32'h38632800;
      81511: inst = 32'h38842800;
      81512: inst = 32'h10a00001;
      81513: inst = 32'hca03e6d;
      81514: inst = 32'h13e00001;
      81515: inst = 32'hfe0d96a;
      81516: inst = 32'h5be00000;
      81517: inst = 32'h8c50000;
      81518: inst = 32'h24612800;
      81519: inst = 32'h10a00000;
      81520: inst = 32'hca00002;
      81521: inst = 32'h24822800;
      81522: inst = 32'h10a00000;
      81523: inst = 32'hca00004;
      81524: inst = 32'h38632800;
      81525: inst = 32'h38842800;
      81526: inst = 32'h10a00001;
      81527: inst = 32'hca03e7b;
      81528: inst = 32'h13e00001;
      81529: inst = 32'hfe0d96a;
      81530: inst = 32'h5be00000;
      81531: inst = 32'h8c50000;
      81532: inst = 32'h24612800;
      81533: inst = 32'h10a00000;
      81534: inst = 32'hca00002;
      81535: inst = 32'h24822800;
      81536: inst = 32'h10a00000;
      81537: inst = 32'hca00004;
      81538: inst = 32'h38632800;
      81539: inst = 32'h38842800;
      81540: inst = 32'h10a00001;
      81541: inst = 32'hca03e89;
      81542: inst = 32'h13e00001;
      81543: inst = 32'hfe0d96a;
      81544: inst = 32'h5be00000;
      81545: inst = 32'h8c50000;
      81546: inst = 32'h24612800;
      81547: inst = 32'h10a00000;
      81548: inst = 32'hca00002;
      81549: inst = 32'h24822800;
      81550: inst = 32'h10a00000;
      81551: inst = 32'hca00004;
      81552: inst = 32'h38632800;
      81553: inst = 32'h38842800;
      81554: inst = 32'h10a00001;
      81555: inst = 32'hca03e97;
      81556: inst = 32'h13e00001;
      81557: inst = 32'hfe0d96a;
      81558: inst = 32'h5be00000;
      81559: inst = 32'h8c50000;
      81560: inst = 32'h24612800;
      81561: inst = 32'h10a00000;
      81562: inst = 32'hca00002;
      81563: inst = 32'h24822800;
      81564: inst = 32'h10a00000;
      81565: inst = 32'hca00004;
      81566: inst = 32'h38632800;
      81567: inst = 32'h38842800;
      81568: inst = 32'h10a00001;
      81569: inst = 32'hca03ea5;
      81570: inst = 32'h13e00001;
      81571: inst = 32'hfe0d96a;
      81572: inst = 32'h5be00000;
      81573: inst = 32'h8c50000;
      81574: inst = 32'h24612800;
      81575: inst = 32'h10a00000;
      81576: inst = 32'hca00002;
      81577: inst = 32'h24822800;
      81578: inst = 32'h10a00000;
      81579: inst = 32'hca00004;
      81580: inst = 32'h38632800;
      81581: inst = 32'h38842800;
      81582: inst = 32'h10a00001;
      81583: inst = 32'hca03eb3;
      81584: inst = 32'h13e00001;
      81585: inst = 32'hfe0d96a;
      81586: inst = 32'h5be00000;
      81587: inst = 32'h8c50000;
      81588: inst = 32'h24612800;
      81589: inst = 32'h10a00000;
      81590: inst = 32'hca00002;
      81591: inst = 32'h24822800;
      81592: inst = 32'h10a00000;
      81593: inst = 32'hca00004;
      81594: inst = 32'h38632800;
      81595: inst = 32'h38842800;
      81596: inst = 32'h10a00001;
      81597: inst = 32'hca03ec1;
      81598: inst = 32'h13e00001;
      81599: inst = 32'hfe0d96a;
      81600: inst = 32'h5be00000;
      81601: inst = 32'h8c50000;
      81602: inst = 32'h24612800;
      81603: inst = 32'h10a00000;
      81604: inst = 32'hca00002;
      81605: inst = 32'h24822800;
      81606: inst = 32'h10a00000;
      81607: inst = 32'hca00004;
      81608: inst = 32'h38632800;
      81609: inst = 32'h38842800;
      81610: inst = 32'h10a00001;
      81611: inst = 32'hca03ecf;
      81612: inst = 32'h13e00001;
      81613: inst = 32'hfe0d96a;
      81614: inst = 32'h5be00000;
      81615: inst = 32'h8c50000;
      81616: inst = 32'h24612800;
      81617: inst = 32'h10a00000;
      81618: inst = 32'hca00002;
      81619: inst = 32'h24822800;
      81620: inst = 32'h10a00000;
      81621: inst = 32'hca00004;
      81622: inst = 32'h38632800;
      81623: inst = 32'h38842800;
      81624: inst = 32'h10a00001;
      81625: inst = 32'hca03edd;
      81626: inst = 32'h13e00001;
      81627: inst = 32'hfe0d96a;
      81628: inst = 32'h5be00000;
      81629: inst = 32'h8c50000;
      81630: inst = 32'h24612800;
      81631: inst = 32'h10a00000;
      81632: inst = 32'hca00002;
      81633: inst = 32'h24822800;
      81634: inst = 32'h10a00000;
      81635: inst = 32'hca00004;
      81636: inst = 32'h38632800;
      81637: inst = 32'h38842800;
      81638: inst = 32'h10a00001;
      81639: inst = 32'hca03eeb;
      81640: inst = 32'h13e00001;
      81641: inst = 32'hfe0d96a;
      81642: inst = 32'h5be00000;
      81643: inst = 32'h8c50000;
      81644: inst = 32'h24612800;
      81645: inst = 32'h10a00000;
      81646: inst = 32'hca00002;
      81647: inst = 32'h24822800;
      81648: inst = 32'h10a00000;
      81649: inst = 32'hca00004;
      81650: inst = 32'h38632800;
      81651: inst = 32'h38842800;
      81652: inst = 32'h10a00001;
      81653: inst = 32'hca03ef9;
      81654: inst = 32'h13e00001;
      81655: inst = 32'hfe0d96a;
      81656: inst = 32'h5be00000;
      81657: inst = 32'h8c50000;
      81658: inst = 32'h24612800;
      81659: inst = 32'h10a00000;
      81660: inst = 32'hca00002;
      81661: inst = 32'h24822800;
      81662: inst = 32'h10a00000;
      81663: inst = 32'hca00004;
      81664: inst = 32'h38632800;
      81665: inst = 32'h38842800;
      81666: inst = 32'h10a00001;
      81667: inst = 32'hca03f07;
      81668: inst = 32'h13e00001;
      81669: inst = 32'hfe0d96a;
      81670: inst = 32'h5be00000;
      81671: inst = 32'h8c50000;
      81672: inst = 32'h24612800;
      81673: inst = 32'h10a00000;
      81674: inst = 32'hca00002;
      81675: inst = 32'h24822800;
      81676: inst = 32'h10a00000;
      81677: inst = 32'hca00004;
      81678: inst = 32'h38632800;
      81679: inst = 32'h38842800;
      81680: inst = 32'h10a00001;
      81681: inst = 32'hca03f15;
      81682: inst = 32'h13e00001;
      81683: inst = 32'hfe0d96a;
      81684: inst = 32'h5be00000;
      81685: inst = 32'h8c50000;
      81686: inst = 32'h24612800;
      81687: inst = 32'h10a00000;
      81688: inst = 32'hca00002;
      81689: inst = 32'h24822800;
      81690: inst = 32'h10a00000;
      81691: inst = 32'hca00004;
      81692: inst = 32'h38632800;
      81693: inst = 32'h38842800;
      81694: inst = 32'h10a00001;
      81695: inst = 32'hca03f23;
      81696: inst = 32'h13e00001;
      81697: inst = 32'hfe0d96a;
      81698: inst = 32'h5be00000;
      81699: inst = 32'h8c50000;
      81700: inst = 32'h24612800;
      81701: inst = 32'h10a00000;
      81702: inst = 32'hca00002;
      81703: inst = 32'h24822800;
      81704: inst = 32'h10a00000;
      81705: inst = 32'hca00004;
      81706: inst = 32'h38632800;
      81707: inst = 32'h38842800;
      81708: inst = 32'h10a00001;
      81709: inst = 32'hca03f31;
      81710: inst = 32'h13e00001;
      81711: inst = 32'hfe0d96a;
      81712: inst = 32'h5be00000;
      81713: inst = 32'h8c50000;
      81714: inst = 32'h24612800;
      81715: inst = 32'h10a00000;
      81716: inst = 32'hca00002;
      81717: inst = 32'h24822800;
      81718: inst = 32'h10a00000;
      81719: inst = 32'hca00004;
      81720: inst = 32'h38632800;
      81721: inst = 32'h38842800;
      81722: inst = 32'h10a00001;
      81723: inst = 32'hca03f3f;
      81724: inst = 32'h13e00001;
      81725: inst = 32'hfe0d96a;
      81726: inst = 32'h5be00000;
      81727: inst = 32'h8c50000;
      81728: inst = 32'h24612800;
      81729: inst = 32'h10a00000;
      81730: inst = 32'hca00002;
      81731: inst = 32'h24822800;
      81732: inst = 32'h10a00000;
      81733: inst = 32'hca00004;
      81734: inst = 32'h38632800;
      81735: inst = 32'h38842800;
      81736: inst = 32'h10a00001;
      81737: inst = 32'hca03f4d;
      81738: inst = 32'h13e00001;
      81739: inst = 32'hfe0d96a;
      81740: inst = 32'h5be00000;
      81741: inst = 32'h8c50000;
      81742: inst = 32'h24612800;
      81743: inst = 32'h10a00000;
      81744: inst = 32'hca00002;
      81745: inst = 32'h24822800;
      81746: inst = 32'h10a00000;
      81747: inst = 32'hca00004;
      81748: inst = 32'h38632800;
      81749: inst = 32'h38842800;
      81750: inst = 32'h10a00001;
      81751: inst = 32'hca03f5b;
      81752: inst = 32'h13e00001;
      81753: inst = 32'hfe0d96a;
      81754: inst = 32'h5be00000;
      81755: inst = 32'h8c50000;
      81756: inst = 32'h24612800;
      81757: inst = 32'h10a00000;
      81758: inst = 32'hca00002;
      81759: inst = 32'h24822800;
      81760: inst = 32'h10a00000;
      81761: inst = 32'hca00004;
      81762: inst = 32'h38632800;
      81763: inst = 32'h38842800;
      81764: inst = 32'h10a00001;
      81765: inst = 32'hca03f69;
      81766: inst = 32'h13e00001;
      81767: inst = 32'hfe0d96a;
      81768: inst = 32'h5be00000;
      81769: inst = 32'h8c50000;
      81770: inst = 32'h24612800;
      81771: inst = 32'h10a00000;
      81772: inst = 32'hca00002;
      81773: inst = 32'h24822800;
      81774: inst = 32'h10a00000;
      81775: inst = 32'hca00004;
      81776: inst = 32'h38632800;
      81777: inst = 32'h38842800;
      81778: inst = 32'h10a00001;
      81779: inst = 32'hca03f77;
      81780: inst = 32'h13e00001;
      81781: inst = 32'hfe0d96a;
      81782: inst = 32'h5be00000;
      81783: inst = 32'h8c50000;
      81784: inst = 32'h24612800;
      81785: inst = 32'h10a00000;
      81786: inst = 32'hca00002;
      81787: inst = 32'h24822800;
      81788: inst = 32'h10a00000;
      81789: inst = 32'hca00004;
      81790: inst = 32'h38632800;
      81791: inst = 32'h38842800;
      81792: inst = 32'h10a00001;
      81793: inst = 32'hca03f85;
      81794: inst = 32'h13e00001;
      81795: inst = 32'hfe0d96a;
      81796: inst = 32'h5be00000;
      81797: inst = 32'h8c50000;
      81798: inst = 32'h24612800;
      81799: inst = 32'h10a00000;
      81800: inst = 32'hca00002;
      81801: inst = 32'h24822800;
      81802: inst = 32'h10a00000;
      81803: inst = 32'hca00004;
      81804: inst = 32'h38632800;
      81805: inst = 32'h38842800;
      81806: inst = 32'h10a00001;
      81807: inst = 32'hca03f93;
      81808: inst = 32'h13e00001;
      81809: inst = 32'hfe0d96a;
      81810: inst = 32'h5be00000;
      81811: inst = 32'h8c50000;
      81812: inst = 32'h24612800;
      81813: inst = 32'h10a00000;
      81814: inst = 32'hca00002;
      81815: inst = 32'h24822800;
      81816: inst = 32'h10a00000;
      81817: inst = 32'hca00004;
      81818: inst = 32'h38632800;
      81819: inst = 32'h38842800;
      81820: inst = 32'h10a00001;
      81821: inst = 32'hca03fa1;
      81822: inst = 32'h13e00001;
      81823: inst = 32'hfe0d96a;
      81824: inst = 32'h5be00000;
      81825: inst = 32'h8c50000;
      81826: inst = 32'h24612800;
      81827: inst = 32'h10a00000;
      81828: inst = 32'hca00002;
      81829: inst = 32'h24822800;
      81830: inst = 32'h10a00000;
      81831: inst = 32'hca00004;
      81832: inst = 32'h38632800;
      81833: inst = 32'h38842800;
      81834: inst = 32'h10a00001;
      81835: inst = 32'hca03faf;
      81836: inst = 32'h13e00001;
      81837: inst = 32'hfe0d96a;
      81838: inst = 32'h5be00000;
      81839: inst = 32'h8c50000;
      81840: inst = 32'h24612800;
      81841: inst = 32'h10a00000;
      81842: inst = 32'hca00002;
      81843: inst = 32'h24822800;
      81844: inst = 32'h10a00000;
      81845: inst = 32'hca00004;
      81846: inst = 32'h38632800;
      81847: inst = 32'h38842800;
      81848: inst = 32'h10a00001;
      81849: inst = 32'hca03fbd;
      81850: inst = 32'h13e00001;
      81851: inst = 32'hfe0d96a;
      81852: inst = 32'h5be00000;
      81853: inst = 32'h8c50000;
      81854: inst = 32'h24612800;
      81855: inst = 32'h10a00000;
      81856: inst = 32'hca00002;
      81857: inst = 32'h24822800;
      81858: inst = 32'h10a00000;
      81859: inst = 32'hca00004;
      81860: inst = 32'h38632800;
      81861: inst = 32'h38842800;
      81862: inst = 32'h10a00001;
      81863: inst = 32'hca03fcb;
      81864: inst = 32'h13e00001;
      81865: inst = 32'hfe0d96a;
      81866: inst = 32'h5be00000;
      81867: inst = 32'h8c50000;
      81868: inst = 32'h24612800;
      81869: inst = 32'h10a00000;
      81870: inst = 32'hca00002;
      81871: inst = 32'h24822800;
      81872: inst = 32'h10a00000;
      81873: inst = 32'hca00004;
      81874: inst = 32'h38632800;
      81875: inst = 32'h38842800;
      81876: inst = 32'h10a00001;
      81877: inst = 32'hca03fd9;
      81878: inst = 32'h13e00001;
      81879: inst = 32'hfe0d96a;
      81880: inst = 32'h5be00000;
      81881: inst = 32'h8c50000;
      81882: inst = 32'h24612800;
      81883: inst = 32'h10a00000;
      81884: inst = 32'hca00002;
      81885: inst = 32'h24822800;
      81886: inst = 32'h10a00000;
      81887: inst = 32'hca00004;
      81888: inst = 32'h38632800;
      81889: inst = 32'h38842800;
      81890: inst = 32'h10a00001;
      81891: inst = 32'hca03fe7;
      81892: inst = 32'h13e00001;
      81893: inst = 32'hfe0d96a;
      81894: inst = 32'h5be00000;
      81895: inst = 32'h8c50000;
      81896: inst = 32'h24612800;
      81897: inst = 32'h10a00000;
      81898: inst = 32'hca00002;
      81899: inst = 32'h24822800;
      81900: inst = 32'h10a00000;
      81901: inst = 32'hca00004;
      81902: inst = 32'h38632800;
      81903: inst = 32'h38842800;
      81904: inst = 32'h10a00001;
      81905: inst = 32'hca03ff5;
      81906: inst = 32'h13e00001;
      81907: inst = 32'hfe0d96a;
      81908: inst = 32'h5be00000;
      81909: inst = 32'h8c50000;
      81910: inst = 32'h24612800;
      81911: inst = 32'h10a00000;
      81912: inst = 32'hca00002;
      81913: inst = 32'h24822800;
      81914: inst = 32'h10a00000;
      81915: inst = 32'hca00004;
      81916: inst = 32'h38632800;
      81917: inst = 32'h38842800;
      81918: inst = 32'h10a00001;
      81919: inst = 32'hca04003;
      81920: inst = 32'h13e00001;
      81921: inst = 32'hfe0d96a;
      81922: inst = 32'h5be00000;
      81923: inst = 32'h8c50000;
      81924: inst = 32'h24612800;
      81925: inst = 32'h10a00000;
      81926: inst = 32'hca00002;
      81927: inst = 32'h24822800;
      81928: inst = 32'h10a00000;
      81929: inst = 32'hca00004;
      81930: inst = 32'h38632800;
      81931: inst = 32'h38842800;
      81932: inst = 32'h10a00001;
      81933: inst = 32'hca04011;
      81934: inst = 32'h13e00001;
      81935: inst = 32'hfe0d96a;
      81936: inst = 32'h5be00000;
      81937: inst = 32'h8c50000;
      81938: inst = 32'h24612800;
      81939: inst = 32'h10a00000;
      81940: inst = 32'hca00002;
      81941: inst = 32'h24822800;
      81942: inst = 32'h10a00000;
      81943: inst = 32'hca00004;
      81944: inst = 32'h38632800;
      81945: inst = 32'h38842800;
      81946: inst = 32'h10a00001;
      81947: inst = 32'hca0401f;
      81948: inst = 32'h13e00001;
      81949: inst = 32'hfe0d96a;
      81950: inst = 32'h5be00000;
      81951: inst = 32'h8c50000;
      81952: inst = 32'h24612800;
      81953: inst = 32'h10a00000;
      81954: inst = 32'hca00002;
      81955: inst = 32'h24822800;
      81956: inst = 32'h10a00000;
      81957: inst = 32'hca00004;
      81958: inst = 32'h38632800;
      81959: inst = 32'h38842800;
      81960: inst = 32'h10a00001;
      81961: inst = 32'hca0402d;
      81962: inst = 32'h13e00001;
      81963: inst = 32'hfe0d96a;
      81964: inst = 32'h5be00000;
      81965: inst = 32'h8c50000;
      81966: inst = 32'h24612800;
      81967: inst = 32'h10a00000;
      81968: inst = 32'hca00002;
      81969: inst = 32'h24822800;
      81970: inst = 32'h10a00000;
      81971: inst = 32'hca00004;
      81972: inst = 32'h38632800;
      81973: inst = 32'h38842800;
      81974: inst = 32'h10a00001;
      81975: inst = 32'hca0403b;
      81976: inst = 32'h13e00001;
      81977: inst = 32'hfe0d96a;
      81978: inst = 32'h5be00000;
      81979: inst = 32'h8c50000;
      81980: inst = 32'h24612800;
      81981: inst = 32'h10a00000;
      81982: inst = 32'hca00002;
      81983: inst = 32'h24822800;
      81984: inst = 32'h10a00000;
      81985: inst = 32'hca00004;
      81986: inst = 32'h38632800;
      81987: inst = 32'h38842800;
      81988: inst = 32'h10a00001;
      81989: inst = 32'hca04049;
      81990: inst = 32'h13e00001;
      81991: inst = 32'hfe0d96a;
      81992: inst = 32'h5be00000;
      81993: inst = 32'h8c50000;
      81994: inst = 32'h24612800;
      81995: inst = 32'h10a00000;
      81996: inst = 32'hca00002;
      81997: inst = 32'h24822800;
      81998: inst = 32'h10a00000;
      81999: inst = 32'hca00004;
      82000: inst = 32'h38632800;
      82001: inst = 32'h38842800;
      82002: inst = 32'h10a00001;
      82003: inst = 32'hca04057;
      82004: inst = 32'h13e00001;
      82005: inst = 32'hfe0d96a;
      82006: inst = 32'h5be00000;
      82007: inst = 32'h8c50000;
      82008: inst = 32'h24612800;
      82009: inst = 32'h10a00000;
      82010: inst = 32'hca00002;
      82011: inst = 32'h24822800;
      82012: inst = 32'h10a00000;
      82013: inst = 32'hca00004;
      82014: inst = 32'h38632800;
      82015: inst = 32'h38842800;
      82016: inst = 32'h10a00001;
      82017: inst = 32'hca04065;
      82018: inst = 32'h13e00001;
      82019: inst = 32'hfe0d96a;
      82020: inst = 32'h5be00000;
      82021: inst = 32'h8c50000;
      82022: inst = 32'h24612800;
      82023: inst = 32'h10a00000;
      82024: inst = 32'hca00002;
      82025: inst = 32'h24822800;
      82026: inst = 32'h10a00000;
      82027: inst = 32'hca00004;
      82028: inst = 32'h38632800;
      82029: inst = 32'h38842800;
      82030: inst = 32'h10a00001;
      82031: inst = 32'hca04073;
      82032: inst = 32'h13e00001;
      82033: inst = 32'hfe0d96a;
      82034: inst = 32'h5be00000;
      82035: inst = 32'h8c50000;
      82036: inst = 32'h24612800;
      82037: inst = 32'h10a00000;
      82038: inst = 32'hca00002;
      82039: inst = 32'h24822800;
      82040: inst = 32'h10a00000;
      82041: inst = 32'hca00004;
      82042: inst = 32'h38632800;
      82043: inst = 32'h38842800;
      82044: inst = 32'h10a00001;
      82045: inst = 32'hca04081;
      82046: inst = 32'h13e00001;
      82047: inst = 32'hfe0d96a;
      82048: inst = 32'h5be00000;
      82049: inst = 32'h8c50000;
      82050: inst = 32'h24612800;
      82051: inst = 32'h10a00000;
      82052: inst = 32'hca00002;
      82053: inst = 32'h24822800;
      82054: inst = 32'h10a00000;
      82055: inst = 32'hca00004;
      82056: inst = 32'h38632800;
      82057: inst = 32'h38842800;
      82058: inst = 32'h10a00001;
      82059: inst = 32'hca0408f;
      82060: inst = 32'h13e00001;
      82061: inst = 32'hfe0d96a;
      82062: inst = 32'h5be00000;
      82063: inst = 32'h8c50000;
      82064: inst = 32'h24612800;
      82065: inst = 32'h10a00000;
      82066: inst = 32'hca00002;
      82067: inst = 32'h24822800;
      82068: inst = 32'h10a00000;
      82069: inst = 32'hca00004;
      82070: inst = 32'h38632800;
      82071: inst = 32'h38842800;
      82072: inst = 32'h10a00001;
      82073: inst = 32'hca0409d;
      82074: inst = 32'h13e00001;
      82075: inst = 32'hfe0d96a;
      82076: inst = 32'h5be00000;
      82077: inst = 32'h8c50000;
      82078: inst = 32'h24612800;
      82079: inst = 32'h10a00000;
      82080: inst = 32'hca00002;
      82081: inst = 32'h24822800;
      82082: inst = 32'h10a00000;
      82083: inst = 32'hca00004;
      82084: inst = 32'h38632800;
      82085: inst = 32'h38842800;
      82086: inst = 32'h10a00001;
      82087: inst = 32'hca040ab;
      82088: inst = 32'h13e00001;
      82089: inst = 32'hfe0d96a;
      82090: inst = 32'h5be00000;
      82091: inst = 32'h8c50000;
      82092: inst = 32'h24612800;
      82093: inst = 32'h10a00000;
      82094: inst = 32'hca00002;
      82095: inst = 32'h24822800;
      82096: inst = 32'h10a00000;
      82097: inst = 32'hca00004;
      82098: inst = 32'h38632800;
      82099: inst = 32'h38842800;
      82100: inst = 32'h10a00001;
      82101: inst = 32'hca040b9;
      82102: inst = 32'h13e00001;
      82103: inst = 32'hfe0d96a;
      82104: inst = 32'h5be00000;
      82105: inst = 32'h8c50000;
      82106: inst = 32'h24612800;
      82107: inst = 32'h10a00000;
      82108: inst = 32'hca00002;
      82109: inst = 32'h24822800;
      82110: inst = 32'h10a00000;
      82111: inst = 32'hca00004;
      82112: inst = 32'h38632800;
      82113: inst = 32'h38842800;
      82114: inst = 32'h10a00001;
      82115: inst = 32'hca040c7;
      82116: inst = 32'h13e00001;
      82117: inst = 32'hfe0d96a;
      82118: inst = 32'h5be00000;
      82119: inst = 32'h8c50000;
      82120: inst = 32'h24612800;
      82121: inst = 32'h10a00000;
      82122: inst = 32'hca00002;
      82123: inst = 32'h24822800;
      82124: inst = 32'h10a00000;
      82125: inst = 32'hca00004;
      82126: inst = 32'h38632800;
      82127: inst = 32'h38842800;
      82128: inst = 32'h10a00001;
      82129: inst = 32'hca040d5;
      82130: inst = 32'h13e00001;
      82131: inst = 32'hfe0d96a;
      82132: inst = 32'h5be00000;
      82133: inst = 32'h8c50000;
      82134: inst = 32'h24612800;
      82135: inst = 32'h10a00000;
      82136: inst = 32'hca00002;
      82137: inst = 32'h24822800;
      82138: inst = 32'h10a00000;
      82139: inst = 32'hca00004;
      82140: inst = 32'h38632800;
      82141: inst = 32'h38842800;
      82142: inst = 32'h10a00001;
      82143: inst = 32'hca040e3;
      82144: inst = 32'h13e00001;
      82145: inst = 32'hfe0d96a;
      82146: inst = 32'h5be00000;
      82147: inst = 32'h8c50000;
      82148: inst = 32'h24612800;
      82149: inst = 32'h10a00000;
      82150: inst = 32'hca00002;
      82151: inst = 32'h24822800;
      82152: inst = 32'h10a00000;
      82153: inst = 32'hca00004;
      82154: inst = 32'h38632800;
      82155: inst = 32'h38842800;
      82156: inst = 32'h10a00001;
      82157: inst = 32'hca040f1;
      82158: inst = 32'h13e00001;
      82159: inst = 32'hfe0d96a;
      82160: inst = 32'h5be00000;
      82161: inst = 32'h8c50000;
      82162: inst = 32'h24612800;
      82163: inst = 32'h10a00000;
      82164: inst = 32'hca00002;
      82165: inst = 32'h24822800;
      82166: inst = 32'h10a00000;
      82167: inst = 32'hca00004;
      82168: inst = 32'h38632800;
      82169: inst = 32'h38842800;
      82170: inst = 32'h10a00001;
      82171: inst = 32'hca040ff;
      82172: inst = 32'h13e00001;
      82173: inst = 32'hfe0d96a;
      82174: inst = 32'h5be00000;
      82175: inst = 32'h8c50000;
      82176: inst = 32'h24612800;
      82177: inst = 32'h10a00000;
      82178: inst = 32'hca00002;
      82179: inst = 32'h24822800;
      82180: inst = 32'h10a00000;
      82181: inst = 32'hca00004;
      82182: inst = 32'h38632800;
      82183: inst = 32'h38842800;
      82184: inst = 32'h10a00001;
      82185: inst = 32'hca0410d;
      82186: inst = 32'h13e00001;
      82187: inst = 32'hfe0d96a;
      82188: inst = 32'h5be00000;
      82189: inst = 32'h8c50000;
      82190: inst = 32'h24612800;
      82191: inst = 32'h10a00000;
      82192: inst = 32'hca00002;
      82193: inst = 32'h24822800;
      82194: inst = 32'h10a00000;
      82195: inst = 32'hca00004;
      82196: inst = 32'h38632800;
      82197: inst = 32'h38842800;
      82198: inst = 32'h10a00001;
      82199: inst = 32'hca0411b;
      82200: inst = 32'h13e00001;
      82201: inst = 32'hfe0d96a;
      82202: inst = 32'h5be00000;
      82203: inst = 32'h8c50000;
      82204: inst = 32'h24612800;
      82205: inst = 32'h10a00000;
      82206: inst = 32'hca00002;
      82207: inst = 32'h24822800;
      82208: inst = 32'h10a00000;
      82209: inst = 32'hca00004;
      82210: inst = 32'h38632800;
      82211: inst = 32'h38842800;
      82212: inst = 32'h10a00001;
      82213: inst = 32'hca04129;
      82214: inst = 32'h13e00001;
      82215: inst = 32'hfe0d96a;
      82216: inst = 32'h5be00000;
      82217: inst = 32'h8c50000;
      82218: inst = 32'h24612800;
      82219: inst = 32'h10a00000;
      82220: inst = 32'hca00003;
      82221: inst = 32'h24822800;
      82222: inst = 32'h10a00000;
      82223: inst = 32'hca00004;
      82224: inst = 32'h38632800;
      82225: inst = 32'h38842800;
      82226: inst = 32'h10a00001;
      82227: inst = 32'hca04137;
      82228: inst = 32'h13e00001;
      82229: inst = 32'hfe0d96a;
      82230: inst = 32'h5be00000;
      82231: inst = 32'h8c50000;
      82232: inst = 32'h24612800;
      82233: inst = 32'h10a00000;
      82234: inst = 32'hca00003;
      82235: inst = 32'h24822800;
      82236: inst = 32'h10a00000;
      82237: inst = 32'hca00004;
      82238: inst = 32'h38632800;
      82239: inst = 32'h38842800;
      82240: inst = 32'h10a00001;
      82241: inst = 32'hca04145;
      82242: inst = 32'h13e00001;
      82243: inst = 32'hfe0d96a;
      82244: inst = 32'h5be00000;
      82245: inst = 32'h8c50000;
      82246: inst = 32'h24612800;
      82247: inst = 32'h10a00000;
      82248: inst = 32'hca00003;
      82249: inst = 32'h24822800;
      82250: inst = 32'h10a00000;
      82251: inst = 32'hca00004;
      82252: inst = 32'h38632800;
      82253: inst = 32'h38842800;
      82254: inst = 32'h10a00001;
      82255: inst = 32'hca04153;
      82256: inst = 32'h13e00001;
      82257: inst = 32'hfe0d96a;
      82258: inst = 32'h5be00000;
      82259: inst = 32'h8c50000;
      82260: inst = 32'h24612800;
      82261: inst = 32'h10a00000;
      82262: inst = 32'hca00003;
      82263: inst = 32'h24822800;
      82264: inst = 32'h10a00000;
      82265: inst = 32'hca00004;
      82266: inst = 32'h38632800;
      82267: inst = 32'h38842800;
      82268: inst = 32'h10a00001;
      82269: inst = 32'hca04161;
      82270: inst = 32'h13e00001;
      82271: inst = 32'hfe0d96a;
      82272: inst = 32'h5be00000;
      82273: inst = 32'h8c50000;
      82274: inst = 32'h24612800;
      82275: inst = 32'h10a00000;
      82276: inst = 32'hca00003;
      82277: inst = 32'h24822800;
      82278: inst = 32'h10a00000;
      82279: inst = 32'hca00004;
      82280: inst = 32'h38632800;
      82281: inst = 32'h38842800;
      82282: inst = 32'h10a00001;
      82283: inst = 32'hca0416f;
      82284: inst = 32'h13e00001;
      82285: inst = 32'hfe0d96a;
      82286: inst = 32'h5be00000;
      82287: inst = 32'h8c50000;
      82288: inst = 32'h24612800;
      82289: inst = 32'h10a00000;
      82290: inst = 32'hca00003;
      82291: inst = 32'h24822800;
      82292: inst = 32'h10a00000;
      82293: inst = 32'hca00004;
      82294: inst = 32'h38632800;
      82295: inst = 32'h38842800;
      82296: inst = 32'h10a00001;
      82297: inst = 32'hca0417d;
      82298: inst = 32'h13e00001;
      82299: inst = 32'hfe0d96a;
      82300: inst = 32'h5be00000;
      82301: inst = 32'h8c50000;
      82302: inst = 32'h24612800;
      82303: inst = 32'h10a00000;
      82304: inst = 32'hca00003;
      82305: inst = 32'h24822800;
      82306: inst = 32'h10a00000;
      82307: inst = 32'hca00004;
      82308: inst = 32'h38632800;
      82309: inst = 32'h38842800;
      82310: inst = 32'h10a00001;
      82311: inst = 32'hca0418b;
      82312: inst = 32'h13e00001;
      82313: inst = 32'hfe0d96a;
      82314: inst = 32'h5be00000;
      82315: inst = 32'h8c50000;
      82316: inst = 32'h24612800;
      82317: inst = 32'h10a00000;
      82318: inst = 32'hca00003;
      82319: inst = 32'h24822800;
      82320: inst = 32'h10a00000;
      82321: inst = 32'hca00004;
      82322: inst = 32'h38632800;
      82323: inst = 32'h38842800;
      82324: inst = 32'h10a00001;
      82325: inst = 32'hca04199;
      82326: inst = 32'h13e00001;
      82327: inst = 32'hfe0d96a;
      82328: inst = 32'h5be00000;
      82329: inst = 32'h8c50000;
      82330: inst = 32'h24612800;
      82331: inst = 32'h10a00000;
      82332: inst = 32'hca00003;
      82333: inst = 32'h24822800;
      82334: inst = 32'h10a00000;
      82335: inst = 32'hca00004;
      82336: inst = 32'h38632800;
      82337: inst = 32'h38842800;
      82338: inst = 32'h10a00001;
      82339: inst = 32'hca041a7;
      82340: inst = 32'h13e00001;
      82341: inst = 32'hfe0d96a;
      82342: inst = 32'h5be00000;
      82343: inst = 32'h8c50000;
      82344: inst = 32'h24612800;
      82345: inst = 32'h10a00000;
      82346: inst = 32'hca00003;
      82347: inst = 32'h24822800;
      82348: inst = 32'h10a00000;
      82349: inst = 32'hca00004;
      82350: inst = 32'h38632800;
      82351: inst = 32'h38842800;
      82352: inst = 32'h10a00001;
      82353: inst = 32'hca041b5;
      82354: inst = 32'h13e00001;
      82355: inst = 32'hfe0d96a;
      82356: inst = 32'h5be00000;
      82357: inst = 32'h8c50000;
      82358: inst = 32'h24612800;
      82359: inst = 32'h10a00000;
      82360: inst = 32'hca00003;
      82361: inst = 32'h24822800;
      82362: inst = 32'h10a00000;
      82363: inst = 32'hca00004;
      82364: inst = 32'h38632800;
      82365: inst = 32'h38842800;
      82366: inst = 32'h10a00001;
      82367: inst = 32'hca041c3;
      82368: inst = 32'h13e00001;
      82369: inst = 32'hfe0d96a;
      82370: inst = 32'h5be00000;
      82371: inst = 32'h8c50000;
      82372: inst = 32'h24612800;
      82373: inst = 32'h10a00000;
      82374: inst = 32'hca00003;
      82375: inst = 32'h24822800;
      82376: inst = 32'h10a00000;
      82377: inst = 32'hca00004;
      82378: inst = 32'h38632800;
      82379: inst = 32'h38842800;
      82380: inst = 32'h10a00001;
      82381: inst = 32'hca041d1;
      82382: inst = 32'h13e00001;
      82383: inst = 32'hfe0d96a;
      82384: inst = 32'h5be00000;
      82385: inst = 32'h8c50000;
      82386: inst = 32'h24612800;
      82387: inst = 32'h10a00000;
      82388: inst = 32'hca00003;
      82389: inst = 32'h24822800;
      82390: inst = 32'h10a00000;
      82391: inst = 32'hca00004;
      82392: inst = 32'h38632800;
      82393: inst = 32'h38842800;
      82394: inst = 32'h10a00001;
      82395: inst = 32'hca041df;
      82396: inst = 32'h13e00001;
      82397: inst = 32'hfe0d96a;
      82398: inst = 32'h5be00000;
      82399: inst = 32'h8c50000;
      82400: inst = 32'h24612800;
      82401: inst = 32'h10a00000;
      82402: inst = 32'hca00003;
      82403: inst = 32'h24822800;
      82404: inst = 32'h10a00000;
      82405: inst = 32'hca00004;
      82406: inst = 32'h38632800;
      82407: inst = 32'h38842800;
      82408: inst = 32'h10a00001;
      82409: inst = 32'hca041ed;
      82410: inst = 32'h13e00001;
      82411: inst = 32'hfe0d96a;
      82412: inst = 32'h5be00000;
      82413: inst = 32'h8c50000;
      82414: inst = 32'h24612800;
      82415: inst = 32'h10a00000;
      82416: inst = 32'hca00003;
      82417: inst = 32'h24822800;
      82418: inst = 32'h10a00000;
      82419: inst = 32'hca00004;
      82420: inst = 32'h38632800;
      82421: inst = 32'h38842800;
      82422: inst = 32'h10a00001;
      82423: inst = 32'hca041fb;
      82424: inst = 32'h13e00001;
      82425: inst = 32'hfe0d96a;
      82426: inst = 32'h5be00000;
      82427: inst = 32'h8c50000;
      82428: inst = 32'h24612800;
      82429: inst = 32'h10a00000;
      82430: inst = 32'hca00003;
      82431: inst = 32'h24822800;
      82432: inst = 32'h10a00000;
      82433: inst = 32'hca00004;
      82434: inst = 32'h38632800;
      82435: inst = 32'h38842800;
      82436: inst = 32'h10a00001;
      82437: inst = 32'hca04209;
      82438: inst = 32'h13e00001;
      82439: inst = 32'hfe0d96a;
      82440: inst = 32'h5be00000;
      82441: inst = 32'h8c50000;
      82442: inst = 32'h24612800;
      82443: inst = 32'h10a00000;
      82444: inst = 32'hca00003;
      82445: inst = 32'h24822800;
      82446: inst = 32'h10a00000;
      82447: inst = 32'hca00004;
      82448: inst = 32'h38632800;
      82449: inst = 32'h38842800;
      82450: inst = 32'h10a00001;
      82451: inst = 32'hca04217;
      82452: inst = 32'h13e00001;
      82453: inst = 32'hfe0d96a;
      82454: inst = 32'h5be00000;
      82455: inst = 32'h8c50000;
      82456: inst = 32'h24612800;
      82457: inst = 32'h10a00000;
      82458: inst = 32'hca00003;
      82459: inst = 32'h24822800;
      82460: inst = 32'h10a00000;
      82461: inst = 32'hca00004;
      82462: inst = 32'h38632800;
      82463: inst = 32'h38842800;
      82464: inst = 32'h10a00001;
      82465: inst = 32'hca04225;
      82466: inst = 32'h13e00001;
      82467: inst = 32'hfe0d96a;
      82468: inst = 32'h5be00000;
      82469: inst = 32'h8c50000;
      82470: inst = 32'h24612800;
      82471: inst = 32'h10a00000;
      82472: inst = 32'hca00003;
      82473: inst = 32'h24822800;
      82474: inst = 32'h10a00000;
      82475: inst = 32'hca00004;
      82476: inst = 32'h38632800;
      82477: inst = 32'h38842800;
      82478: inst = 32'h10a00001;
      82479: inst = 32'hca04233;
      82480: inst = 32'h13e00001;
      82481: inst = 32'hfe0d96a;
      82482: inst = 32'h5be00000;
      82483: inst = 32'h8c50000;
      82484: inst = 32'h24612800;
      82485: inst = 32'h10a00000;
      82486: inst = 32'hca00003;
      82487: inst = 32'h24822800;
      82488: inst = 32'h10a00000;
      82489: inst = 32'hca00004;
      82490: inst = 32'h38632800;
      82491: inst = 32'h38842800;
      82492: inst = 32'h10a00001;
      82493: inst = 32'hca04241;
      82494: inst = 32'h13e00001;
      82495: inst = 32'hfe0d96a;
      82496: inst = 32'h5be00000;
      82497: inst = 32'h8c50000;
      82498: inst = 32'h24612800;
      82499: inst = 32'h10a00000;
      82500: inst = 32'hca00003;
      82501: inst = 32'h24822800;
      82502: inst = 32'h10a00000;
      82503: inst = 32'hca00004;
      82504: inst = 32'h38632800;
      82505: inst = 32'h38842800;
      82506: inst = 32'h10a00001;
      82507: inst = 32'hca0424f;
      82508: inst = 32'h13e00001;
      82509: inst = 32'hfe0d96a;
      82510: inst = 32'h5be00000;
      82511: inst = 32'h8c50000;
      82512: inst = 32'h24612800;
      82513: inst = 32'h10a00000;
      82514: inst = 32'hca00003;
      82515: inst = 32'h24822800;
      82516: inst = 32'h10a00000;
      82517: inst = 32'hca00004;
      82518: inst = 32'h38632800;
      82519: inst = 32'h38842800;
      82520: inst = 32'h10a00001;
      82521: inst = 32'hca0425d;
      82522: inst = 32'h13e00001;
      82523: inst = 32'hfe0d96a;
      82524: inst = 32'h5be00000;
      82525: inst = 32'h8c50000;
      82526: inst = 32'h24612800;
      82527: inst = 32'h10a00000;
      82528: inst = 32'hca00003;
      82529: inst = 32'h24822800;
      82530: inst = 32'h10a00000;
      82531: inst = 32'hca00004;
      82532: inst = 32'h38632800;
      82533: inst = 32'h38842800;
      82534: inst = 32'h10a00001;
      82535: inst = 32'hca0426b;
      82536: inst = 32'h13e00001;
      82537: inst = 32'hfe0d96a;
      82538: inst = 32'h5be00000;
      82539: inst = 32'h8c50000;
      82540: inst = 32'h24612800;
      82541: inst = 32'h10a00000;
      82542: inst = 32'hca00003;
      82543: inst = 32'h24822800;
      82544: inst = 32'h10a00000;
      82545: inst = 32'hca00004;
      82546: inst = 32'h38632800;
      82547: inst = 32'h38842800;
      82548: inst = 32'h10a00001;
      82549: inst = 32'hca04279;
      82550: inst = 32'h13e00001;
      82551: inst = 32'hfe0d96a;
      82552: inst = 32'h5be00000;
      82553: inst = 32'h8c50000;
      82554: inst = 32'h24612800;
      82555: inst = 32'h10a00000;
      82556: inst = 32'hca00003;
      82557: inst = 32'h24822800;
      82558: inst = 32'h10a00000;
      82559: inst = 32'hca00004;
      82560: inst = 32'h38632800;
      82561: inst = 32'h38842800;
      82562: inst = 32'h10a00001;
      82563: inst = 32'hca04287;
      82564: inst = 32'h13e00001;
      82565: inst = 32'hfe0d96a;
      82566: inst = 32'h5be00000;
      82567: inst = 32'h8c50000;
      82568: inst = 32'h24612800;
      82569: inst = 32'h10a00000;
      82570: inst = 32'hca00003;
      82571: inst = 32'h24822800;
      82572: inst = 32'h10a00000;
      82573: inst = 32'hca00004;
      82574: inst = 32'h38632800;
      82575: inst = 32'h38842800;
      82576: inst = 32'h10a00001;
      82577: inst = 32'hca04295;
      82578: inst = 32'h13e00001;
      82579: inst = 32'hfe0d96a;
      82580: inst = 32'h5be00000;
      82581: inst = 32'h8c50000;
      82582: inst = 32'h24612800;
      82583: inst = 32'h10a00000;
      82584: inst = 32'hca00003;
      82585: inst = 32'h24822800;
      82586: inst = 32'h10a00000;
      82587: inst = 32'hca00004;
      82588: inst = 32'h38632800;
      82589: inst = 32'h38842800;
      82590: inst = 32'h10a00001;
      82591: inst = 32'hca042a3;
      82592: inst = 32'h13e00001;
      82593: inst = 32'hfe0d96a;
      82594: inst = 32'h5be00000;
      82595: inst = 32'h8c50000;
      82596: inst = 32'h24612800;
      82597: inst = 32'h10a00000;
      82598: inst = 32'hca00003;
      82599: inst = 32'h24822800;
      82600: inst = 32'h10a00000;
      82601: inst = 32'hca00004;
      82602: inst = 32'h38632800;
      82603: inst = 32'h38842800;
      82604: inst = 32'h10a00001;
      82605: inst = 32'hca042b1;
      82606: inst = 32'h13e00001;
      82607: inst = 32'hfe0d96a;
      82608: inst = 32'h5be00000;
      82609: inst = 32'h8c50000;
      82610: inst = 32'h24612800;
      82611: inst = 32'h10a00000;
      82612: inst = 32'hca00003;
      82613: inst = 32'h24822800;
      82614: inst = 32'h10a00000;
      82615: inst = 32'hca00004;
      82616: inst = 32'h38632800;
      82617: inst = 32'h38842800;
      82618: inst = 32'h10a00001;
      82619: inst = 32'hca042bf;
      82620: inst = 32'h13e00001;
      82621: inst = 32'hfe0d96a;
      82622: inst = 32'h5be00000;
      82623: inst = 32'h8c50000;
      82624: inst = 32'h24612800;
      82625: inst = 32'h10a00000;
      82626: inst = 32'hca00003;
      82627: inst = 32'h24822800;
      82628: inst = 32'h10a00000;
      82629: inst = 32'hca00004;
      82630: inst = 32'h38632800;
      82631: inst = 32'h38842800;
      82632: inst = 32'h10a00001;
      82633: inst = 32'hca042cd;
      82634: inst = 32'h13e00001;
      82635: inst = 32'hfe0d96a;
      82636: inst = 32'h5be00000;
      82637: inst = 32'h8c50000;
      82638: inst = 32'h24612800;
      82639: inst = 32'h10a00000;
      82640: inst = 32'hca00003;
      82641: inst = 32'h24822800;
      82642: inst = 32'h10a00000;
      82643: inst = 32'hca00004;
      82644: inst = 32'h38632800;
      82645: inst = 32'h38842800;
      82646: inst = 32'h10a00001;
      82647: inst = 32'hca042db;
      82648: inst = 32'h13e00001;
      82649: inst = 32'hfe0d96a;
      82650: inst = 32'h5be00000;
      82651: inst = 32'h8c50000;
      82652: inst = 32'h24612800;
      82653: inst = 32'h10a00000;
      82654: inst = 32'hca00003;
      82655: inst = 32'h24822800;
      82656: inst = 32'h10a00000;
      82657: inst = 32'hca00004;
      82658: inst = 32'h38632800;
      82659: inst = 32'h38842800;
      82660: inst = 32'h10a00001;
      82661: inst = 32'hca042e9;
      82662: inst = 32'h13e00001;
      82663: inst = 32'hfe0d96a;
      82664: inst = 32'h5be00000;
      82665: inst = 32'h8c50000;
      82666: inst = 32'h24612800;
      82667: inst = 32'h10a00000;
      82668: inst = 32'hca00003;
      82669: inst = 32'h24822800;
      82670: inst = 32'h10a00000;
      82671: inst = 32'hca00004;
      82672: inst = 32'h38632800;
      82673: inst = 32'h38842800;
      82674: inst = 32'h10a00001;
      82675: inst = 32'hca042f7;
      82676: inst = 32'h13e00001;
      82677: inst = 32'hfe0d96a;
      82678: inst = 32'h5be00000;
      82679: inst = 32'h8c50000;
      82680: inst = 32'h24612800;
      82681: inst = 32'h10a00000;
      82682: inst = 32'hca00003;
      82683: inst = 32'h24822800;
      82684: inst = 32'h10a00000;
      82685: inst = 32'hca00004;
      82686: inst = 32'h38632800;
      82687: inst = 32'h38842800;
      82688: inst = 32'h10a00001;
      82689: inst = 32'hca04305;
      82690: inst = 32'h13e00001;
      82691: inst = 32'hfe0d96a;
      82692: inst = 32'h5be00000;
      82693: inst = 32'h8c50000;
      82694: inst = 32'h24612800;
      82695: inst = 32'h10a00000;
      82696: inst = 32'hca00003;
      82697: inst = 32'h24822800;
      82698: inst = 32'h10a00000;
      82699: inst = 32'hca00004;
      82700: inst = 32'h38632800;
      82701: inst = 32'h38842800;
      82702: inst = 32'h10a00001;
      82703: inst = 32'hca04313;
      82704: inst = 32'h13e00001;
      82705: inst = 32'hfe0d96a;
      82706: inst = 32'h5be00000;
      82707: inst = 32'h8c50000;
      82708: inst = 32'h24612800;
      82709: inst = 32'h10a00000;
      82710: inst = 32'hca00003;
      82711: inst = 32'h24822800;
      82712: inst = 32'h10a00000;
      82713: inst = 32'hca00004;
      82714: inst = 32'h38632800;
      82715: inst = 32'h38842800;
      82716: inst = 32'h10a00001;
      82717: inst = 32'hca04321;
      82718: inst = 32'h13e00001;
      82719: inst = 32'hfe0d96a;
      82720: inst = 32'h5be00000;
      82721: inst = 32'h8c50000;
      82722: inst = 32'h24612800;
      82723: inst = 32'h10a00000;
      82724: inst = 32'hca00003;
      82725: inst = 32'h24822800;
      82726: inst = 32'h10a00000;
      82727: inst = 32'hca00004;
      82728: inst = 32'h38632800;
      82729: inst = 32'h38842800;
      82730: inst = 32'h10a00001;
      82731: inst = 32'hca0432f;
      82732: inst = 32'h13e00001;
      82733: inst = 32'hfe0d96a;
      82734: inst = 32'h5be00000;
      82735: inst = 32'h8c50000;
      82736: inst = 32'h24612800;
      82737: inst = 32'h10a00000;
      82738: inst = 32'hca00003;
      82739: inst = 32'h24822800;
      82740: inst = 32'h10a00000;
      82741: inst = 32'hca00004;
      82742: inst = 32'h38632800;
      82743: inst = 32'h38842800;
      82744: inst = 32'h10a00001;
      82745: inst = 32'hca0433d;
      82746: inst = 32'h13e00001;
      82747: inst = 32'hfe0d96a;
      82748: inst = 32'h5be00000;
      82749: inst = 32'h8c50000;
      82750: inst = 32'h24612800;
      82751: inst = 32'h10a00000;
      82752: inst = 32'hca00003;
      82753: inst = 32'h24822800;
      82754: inst = 32'h10a00000;
      82755: inst = 32'hca00004;
      82756: inst = 32'h38632800;
      82757: inst = 32'h38842800;
      82758: inst = 32'h10a00001;
      82759: inst = 32'hca0434b;
      82760: inst = 32'h13e00001;
      82761: inst = 32'hfe0d96a;
      82762: inst = 32'h5be00000;
      82763: inst = 32'h8c50000;
      82764: inst = 32'h24612800;
      82765: inst = 32'h10a00000;
      82766: inst = 32'hca00003;
      82767: inst = 32'h24822800;
      82768: inst = 32'h10a00000;
      82769: inst = 32'hca00004;
      82770: inst = 32'h38632800;
      82771: inst = 32'h38842800;
      82772: inst = 32'h10a00001;
      82773: inst = 32'hca04359;
      82774: inst = 32'h13e00001;
      82775: inst = 32'hfe0d96a;
      82776: inst = 32'h5be00000;
      82777: inst = 32'h8c50000;
      82778: inst = 32'h24612800;
      82779: inst = 32'h10a00000;
      82780: inst = 32'hca00003;
      82781: inst = 32'h24822800;
      82782: inst = 32'h10a00000;
      82783: inst = 32'hca00004;
      82784: inst = 32'h38632800;
      82785: inst = 32'h38842800;
      82786: inst = 32'h10a00001;
      82787: inst = 32'hca04367;
      82788: inst = 32'h13e00001;
      82789: inst = 32'hfe0d96a;
      82790: inst = 32'h5be00000;
      82791: inst = 32'h8c50000;
      82792: inst = 32'h24612800;
      82793: inst = 32'h10a00000;
      82794: inst = 32'hca00003;
      82795: inst = 32'h24822800;
      82796: inst = 32'h10a00000;
      82797: inst = 32'hca00004;
      82798: inst = 32'h38632800;
      82799: inst = 32'h38842800;
      82800: inst = 32'h10a00001;
      82801: inst = 32'hca04375;
      82802: inst = 32'h13e00001;
      82803: inst = 32'hfe0d96a;
      82804: inst = 32'h5be00000;
      82805: inst = 32'h8c50000;
      82806: inst = 32'h24612800;
      82807: inst = 32'h10a00000;
      82808: inst = 32'hca00003;
      82809: inst = 32'h24822800;
      82810: inst = 32'h10a00000;
      82811: inst = 32'hca00004;
      82812: inst = 32'h38632800;
      82813: inst = 32'h38842800;
      82814: inst = 32'h10a00001;
      82815: inst = 32'hca04383;
      82816: inst = 32'h13e00001;
      82817: inst = 32'hfe0d96a;
      82818: inst = 32'h5be00000;
      82819: inst = 32'h8c50000;
      82820: inst = 32'h24612800;
      82821: inst = 32'h10a00000;
      82822: inst = 32'hca00003;
      82823: inst = 32'h24822800;
      82824: inst = 32'h10a00000;
      82825: inst = 32'hca00004;
      82826: inst = 32'h38632800;
      82827: inst = 32'h38842800;
      82828: inst = 32'h10a00001;
      82829: inst = 32'hca04391;
      82830: inst = 32'h13e00001;
      82831: inst = 32'hfe0d96a;
      82832: inst = 32'h5be00000;
      82833: inst = 32'h8c50000;
      82834: inst = 32'h24612800;
      82835: inst = 32'h10a00000;
      82836: inst = 32'hca00003;
      82837: inst = 32'h24822800;
      82838: inst = 32'h10a00000;
      82839: inst = 32'hca00004;
      82840: inst = 32'h38632800;
      82841: inst = 32'h38842800;
      82842: inst = 32'h10a00001;
      82843: inst = 32'hca0439f;
      82844: inst = 32'h13e00001;
      82845: inst = 32'hfe0d96a;
      82846: inst = 32'h5be00000;
      82847: inst = 32'h8c50000;
      82848: inst = 32'h24612800;
      82849: inst = 32'h10a00000;
      82850: inst = 32'hca00003;
      82851: inst = 32'h24822800;
      82852: inst = 32'h10a00000;
      82853: inst = 32'hca00004;
      82854: inst = 32'h38632800;
      82855: inst = 32'h38842800;
      82856: inst = 32'h10a00001;
      82857: inst = 32'hca043ad;
      82858: inst = 32'h13e00001;
      82859: inst = 32'hfe0d96a;
      82860: inst = 32'h5be00000;
      82861: inst = 32'h8c50000;
      82862: inst = 32'h24612800;
      82863: inst = 32'h10a00000;
      82864: inst = 32'hca00003;
      82865: inst = 32'h24822800;
      82866: inst = 32'h10a00000;
      82867: inst = 32'hca00004;
      82868: inst = 32'h38632800;
      82869: inst = 32'h38842800;
      82870: inst = 32'h10a00001;
      82871: inst = 32'hca043bb;
      82872: inst = 32'h13e00001;
      82873: inst = 32'hfe0d96a;
      82874: inst = 32'h5be00000;
      82875: inst = 32'h8c50000;
      82876: inst = 32'h24612800;
      82877: inst = 32'h10a00000;
      82878: inst = 32'hca00003;
      82879: inst = 32'h24822800;
      82880: inst = 32'h10a00000;
      82881: inst = 32'hca00004;
      82882: inst = 32'h38632800;
      82883: inst = 32'h38842800;
      82884: inst = 32'h10a00001;
      82885: inst = 32'hca043c9;
      82886: inst = 32'h13e00001;
      82887: inst = 32'hfe0d96a;
      82888: inst = 32'h5be00000;
      82889: inst = 32'h8c50000;
      82890: inst = 32'h24612800;
      82891: inst = 32'h10a00000;
      82892: inst = 32'hca00003;
      82893: inst = 32'h24822800;
      82894: inst = 32'h10a00000;
      82895: inst = 32'hca00004;
      82896: inst = 32'h38632800;
      82897: inst = 32'h38842800;
      82898: inst = 32'h10a00001;
      82899: inst = 32'hca043d7;
      82900: inst = 32'h13e00001;
      82901: inst = 32'hfe0d96a;
      82902: inst = 32'h5be00000;
      82903: inst = 32'h8c50000;
      82904: inst = 32'h24612800;
      82905: inst = 32'h10a00000;
      82906: inst = 32'hca00003;
      82907: inst = 32'h24822800;
      82908: inst = 32'h10a00000;
      82909: inst = 32'hca00004;
      82910: inst = 32'h38632800;
      82911: inst = 32'h38842800;
      82912: inst = 32'h10a00001;
      82913: inst = 32'hca043e5;
      82914: inst = 32'h13e00001;
      82915: inst = 32'hfe0d96a;
      82916: inst = 32'h5be00000;
      82917: inst = 32'h8c50000;
      82918: inst = 32'h24612800;
      82919: inst = 32'h10a00000;
      82920: inst = 32'hca00003;
      82921: inst = 32'h24822800;
      82922: inst = 32'h10a00000;
      82923: inst = 32'hca00004;
      82924: inst = 32'h38632800;
      82925: inst = 32'h38842800;
      82926: inst = 32'h10a00001;
      82927: inst = 32'hca043f3;
      82928: inst = 32'h13e00001;
      82929: inst = 32'hfe0d96a;
      82930: inst = 32'h5be00000;
      82931: inst = 32'h8c50000;
      82932: inst = 32'h24612800;
      82933: inst = 32'h10a00000;
      82934: inst = 32'hca00003;
      82935: inst = 32'h24822800;
      82936: inst = 32'h10a00000;
      82937: inst = 32'hca00004;
      82938: inst = 32'h38632800;
      82939: inst = 32'h38842800;
      82940: inst = 32'h10a00001;
      82941: inst = 32'hca04401;
      82942: inst = 32'h13e00001;
      82943: inst = 32'hfe0d96a;
      82944: inst = 32'h5be00000;
      82945: inst = 32'h8c50000;
      82946: inst = 32'h24612800;
      82947: inst = 32'h10a00000;
      82948: inst = 32'hca00003;
      82949: inst = 32'h24822800;
      82950: inst = 32'h10a00000;
      82951: inst = 32'hca00004;
      82952: inst = 32'h38632800;
      82953: inst = 32'h38842800;
      82954: inst = 32'h10a00001;
      82955: inst = 32'hca0440f;
      82956: inst = 32'h13e00001;
      82957: inst = 32'hfe0d96a;
      82958: inst = 32'h5be00000;
      82959: inst = 32'h8c50000;
      82960: inst = 32'h24612800;
      82961: inst = 32'h10a00000;
      82962: inst = 32'hca00003;
      82963: inst = 32'h24822800;
      82964: inst = 32'h10a00000;
      82965: inst = 32'hca00004;
      82966: inst = 32'h38632800;
      82967: inst = 32'h38842800;
      82968: inst = 32'h10a00001;
      82969: inst = 32'hca0441d;
      82970: inst = 32'h13e00001;
      82971: inst = 32'hfe0d96a;
      82972: inst = 32'h5be00000;
      82973: inst = 32'h8c50000;
      82974: inst = 32'h24612800;
      82975: inst = 32'h10a00000;
      82976: inst = 32'hca00003;
      82977: inst = 32'h24822800;
      82978: inst = 32'h10a00000;
      82979: inst = 32'hca00004;
      82980: inst = 32'h38632800;
      82981: inst = 32'h38842800;
      82982: inst = 32'h10a00001;
      82983: inst = 32'hca0442b;
      82984: inst = 32'h13e00001;
      82985: inst = 32'hfe0d96a;
      82986: inst = 32'h5be00000;
      82987: inst = 32'h8c50000;
      82988: inst = 32'h24612800;
      82989: inst = 32'h10a00000;
      82990: inst = 32'hca00003;
      82991: inst = 32'h24822800;
      82992: inst = 32'h10a00000;
      82993: inst = 32'hca00004;
      82994: inst = 32'h38632800;
      82995: inst = 32'h38842800;
      82996: inst = 32'h10a00001;
      82997: inst = 32'hca04439;
      82998: inst = 32'h13e00001;
      82999: inst = 32'hfe0d96a;
      83000: inst = 32'h5be00000;
      83001: inst = 32'h8c50000;
      83002: inst = 32'h24612800;
      83003: inst = 32'h10a00000;
      83004: inst = 32'hca00003;
      83005: inst = 32'h24822800;
      83006: inst = 32'h10a00000;
      83007: inst = 32'hca00004;
      83008: inst = 32'h38632800;
      83009: inst = 32'h38842800;
      83010: inst = 32'h10a00001;
      83011: inst = 32'hca04447;
      83012: inst = 32'h13e00001;
      83013: inst = 32'hfe0d96a;
      83014: inst = 32'h5be00000;
      83015: inst = 32'h8c50000;
      83016: inst = 32'h24612800;
      83017: inst = 32'h10a00000;
      83018: inst = 32'hca00003;
      83019: inst = 32'h24822800;
      83020: inst = 32'h10a00000;
      83021: inst = 32'hca00004;
      83022: inst = 32'h38632800;
      83023: inst = 32'h38842800;
      83024: inst = 32'h10a00001;
      83025: inst = 32'hca04455;
      83026: inst = 32'h13e00001;
      83027: inst = 32'hfe0d96a;
      83028: inst = 32'h5be00000;
      83029: inst = 32'h8c50000;
      83030: inst = 32'h24612800;
      83031: inst = 32'h10a00000;
      83032: inst = 32'hca00003;
      83033: inst = 32'h24822800;
      83034: inst = 32'h10a00000;
      83035: inst = 32'hca00004;
      83036: inst = 32'h38632800;
      83037: inst = 32'h38842800;
      83038: inst = 32'h10a00001;
      83039: inst = 32'hca04463;
      83040: inst = 32'h13e00001;
      83041: inst = 32'hfe0d96a;
      83042: inst = 32'h5be00000;
      83043: inst = 32'h8c50000;
      83044: inst = 32'h24612800;
      83045: inst = 32'h10a00000;
      83046: inst = 32'hca00003;
      83047: inst = 32'h24822800;
      83048: inst = 32'h10a00000;
      83049: inst = 32'hca00004;
      83050: inst = 32'h38632800;
      83051: inst = 32'h38842800;
      83052: inst = 32'h10a00001;
      83053: inst = 32'hca04471;
      83054: inst = 32'h13e00001;
      83055: inst = 32'hfe0d96a;
      83056: inst = 32'h5be00000;
      83057: inst = 32'h8c50000;
      83058: inst = 32'h24612800;
      83059: inst = 32'h10a00000;
      83060: inst = 32'hca00003;
      83061: inst = 32'h24822800;
      83062: inst = 32'h10a00000;
      83063: inst = 32'hca00004;
      83064: inst = 32'h38632800;
      83065: inst = 32'h38842800;
      83066: inst = 32'h10a00001;
      83067: inst = 32'hca0447f;
      83068: inst = 32'h13e00001;
      83069: inst = 32'hfe0d96a;
      83070: inst = 32'h5be00000;
      83071: inst = 32'h8c50000;
      83072: inst = 32'h24612800;
      83073: inst = 32'h10a00000;
      83074: inst = 32'hca00003;
      83075: inst = 32'h24822800;
      83076: inst = 32'h10a00000;
      83077: inst = 32'hca00004;
      83078: inst = 32'h38632800;
      83079: inst = 32'h38842800;
      83080: inst = 32'h10a00001;
      83081: inst = 32'hca0448d;
      83082: inst = 32'h13e00001;
      83083: inst = 32'hfe0d96a;
      83084: inst = 32'h5be00000;
      83085: inst = 32'h8c50000;
      83086: inst = 32'h24612800;
      83087: inst = 32'h10a00000;
      83088: inst = 32'hca00003;
      83089: inst = 32'h24822800;
      83090: inst = 32'h10a00000;
      83091: inst = 32'hca00004;
      83092: inst = 32'h38632800;
      83093: inst = 32'h38842800;
      83094: inst = 32'h10a00001;
      83095: inst = 32'hca0449b;
      83096: inst = 32'h13e00001;
      83097: inst = 32'hfe0d96a;
      83098: inst = 32'h5be00000;
      83099: inst = 32'h8c50000;
      83100: inst = 32'h24612800;
      83101: inst = 32'h10a00000;
      83102: inst = 32'hca00003;
      83103: inst = 32'h24822800;
      83104: inst = 32'h10a00000;
      83105: inst = 32'hca00004;
      83106: inst = 32'h38632800;
      83107: inst = 32'h38842800;
      83108: inst = 32'h10a00001;
      83109: inst = 32'hca044a9;
      83110: inst = 32'h13e00001;
      83111: inst = 32'hfe0d96a;
      83112: inst = 32'h5be00000;
      83113: inst = 32'h8c50000;
      83114: inst = 32'h24612800;
      83115: inst = 32'h10a00000;
      83116: inst = 32'hca00003;
      83117: inst = 32'h24822800;
      83118: inst = 32'h10a00000;
      83119: inst = 32'hca00004;
      83120: inst = 32'h38632800;
      83121: inst = 32'h38842800;
      83122: inst = 32'h10a00001;
      83123: inst = 32'hca044b7;
      83124: inst = 32'h13e00001;
      83125: inst = 32'hfe0d96a;
      83126: inst = 32'h5be00000;
      83127: inst = 32'h8c50000;
      83128: inst = 32'h24612800;
      83129: inst = 32'h10a00000;
      83130: inst = 32'hca00003;
      83131: inst = 32'h24822800;
      83132: inst = 32'h10a00000;
      83133: inst = 32'hca00004;
      83134: inst = 32'h38632800;
      83135: inst = 32'h38842800;
      83136: inst = 32'h10a00001;
      83137: inst = 32'hca044c5;
      83138: inst = 32'h13e00001;
      83139: inst = 32'hfe0d96a;
      83140: inst = 32'h5be00000;
      83141: inst = 32'h8c50000;
      83142: inst = 32'h24612800;
      83143: inst = 32'h10a00000;
      83144: inst = 32'hca00003;
      83145: inst = 32'h24822800;
      83146: inst = 32'h10a00000;
      83147: inst = 32'hca00004;
      83148: inst = 32'h38632800;
      83149: inst = 32'h38842800;
      83150: inst = 32'h10a00001;
      83151: inst = 32'hca044d3;
      83152: inst = 32'h13e00001;
      83153: inst = 32'hfe0d96a;
      83154: inst = 32'h5be00000;
      83155: inst = 32'h8c50000;
      83156: inst = 32'h24612800;
      83157: inst = 32'h10a00000;
      83158: inst = 32'hca00003;
      83159: inst = 32'h24822800;
      83160: inst = 32'h10a00000;
      83161: inst = 32'hca00004;
      83162: inst = 32'h38632800;
      83163: inst = 32'h38842800;
      83164: inst = 32'h10a00001;
      83165: inst = 32'hca044e1;
      83166: inst = 32'h13e00001;
      83167: inst = 32'hfe0d96a;
      83168: inst = 32'h5be00000;
      83169: inst = 32'h8c50000;
      83170: inst = 32'h24612800;
      83171: inst = 32'h10a00000;
      83172: inst = 32'hca00003;
      83173: inst = 32'h24822800;
      83174: inst = 32'h10a00000;
      83175: inst = 32'hca00004;
      83176: inst = 32'h38632800;
      83177: inst = 32'h38842800;
      83178: inst = 32'h10a00001;
      83179: inst = 32'hca044ef;
      83180: inst = 32'h13e00001;
      83181: inst = 32'hfe0d96a;
      83182: inst = 32'h5be00000;
      83183: inst = 32'h8c50000;
      83184: inst = 32'h24612800;
      83185: inst = 32'h10a00000;
      83186: inst = 32'hca00003;
      83187: inst = 32'h24822800;
      83188: inst = 32'h10a00000;
      83189: inst = 32'hca00004;
      83190: inst = 32'h38632800;
      83191: inst = 32'h38842800;
      83192: inst = 32'h10a00001;
      83193: inst = 32'hca044fd;
      83194: inst = 32'h13e00001;
      83195: inst = 32'hfe0d96a;
      83196: inst = 32'h5be00000;
      83197: inst = 32'h8c50000;
      83198: inst = 32'h24612800;
      83199: inst = 32'h10a00000;
      83200: inst = 32'hca00003;
      83201: inst = 32'h24822800;
      83202: inst = 32'h10a00000;
      83203: inst = 32'hca00004;
      83204: inst = 32'h38632800;
      83205: inst = 32'h38842800;
      83206: inst = 32'h10a00001;
      83207: inst = 32'hca0450b;
      83208: inst = 32'h13e00001;
      83209: inst = 32'hfe0d96a;
      83210: inst = 32'h5be00000;
      83211: inst = 32'h8c50000;
      83212: inst = 32'h24612800;
      83213: inst = 32'h10a00000;
      83214: inst = 32'hca00003;
      83215: inst = 32'h24822800;
      83216: inst = 32'h10a00000;
      83217: inst = 32'hca00004;
      83218: inst = 32'h38632800;
      83219: inst = 32'h38842800;
      83220: inst = 32'h10a00001;
      83221: inst = 32'hca04519;
      83222: inst = 32'h13e00001;
      83223: inst = 32'hfe0d96a;
      83224: inst = 32'h5be00000;
      83225: inst = 32'h8c50000;
      83226: inst = 32'h24612800;
      83227: inst = 32'h10a00000;
      83228: inst = 32'hca00003;
      83229: inst = 32'h24822800;
      83230: inst = 32'h10a00000;
      83231: inst = 32'hca00004;
      83232: inst = 32'h38632800;
      83233: inst = 32'h38842800;
      83234: inst = 32'h10a00001;
      83235: inst = 32'hca04527;
      83236: inst = 32'h13e00001;
      83237: inst = 32'hfe0d96a;
      83238: inst = 32'h5be00000;
      83239: inst = 32'h8c50000;
      83240: inst = 32'h24612800;
      83241: inst = 32'h10a00000;
      83242: inst = 32'hca00003;
      83243: inst = 32'h24822800;
      83244: inst = 32'h10a00000;
      83245: inst = 32'hca00004;
      83246: inst = 32'h38632800;
      83247: inst = 32'h38842800;
      83248: inst = 32'h10a00001;
      83249: inst = 32'hca04535;
      83250: inst = 32'h13e00001;
      83251: inst = 32'hfe0d96a;
      83252: inst = 32'h5be00000;
      83253: inst = 32'h8c50000;
      83254: inst = 32'h24612800;
      83255: inst = 32'h10a00000;
      83256: inst = 32'hca00003;
      83257: inst = 32'h24822800;
      83258: inst = 32'h10a00000;
      83259: inst = 32'hca00004;
      83260: inst = 32'h38632800;
      83261: inst = 32'h38842800;
      83262: inst = 32'h10a00001;
      83263: inst = 32'hca04543;
      83264: inst = 32'h13e00001;
      83265: inst = 32'hfe0d96a;
      83266: inst = 32'h5be00000;
      83267: inst = 32'h8c50000;
      83268: inst = 32'h24612800;
      83269: inst = 32'h10a00000;
      83270: inst = 32'hca00003;
      83271: inst = 32'h24822800;
      83272: inst = 32'h10a00000;
      83273: inst = 32'hca00004;
      83274: inst = 32'h38632800;
      83275: inst = 32'h38842800;
      83276: inst = 32'h10a00001;
      83277: inst = 32'hca04551;
      83278: inst = 32'h13e00001;
      83279: inst = 32'hfe0d96a;
      83280: inst = 32'h5be00000;
      83281: inst = 32'h8c50000;
      83282: inst = 32'h24612800;
      83283: inst = 32'h10a00000;
      83284: inst = 32'hca00003;
      83285: inst = 32'h24822800;
      83286: inst = 32'h10a00000;
      83287: inst = 32'hca00004;
      83288: inst = 32'h38632800;
      83289: inst = 32'h38842800;
      83290: inst = 32'h10a00001;
      83291: inst = 32'hca0455f;
      83292: inst = 32'h13e00001;
      83293: inst = 32'hfe0d96a;
      83294: inst = 32'h5be00000;
      83295: inst = 32'h8c50000;
      83296: inst = 32'h24612800;
      83297: inst = 32'h10a00000;
      83298: inst = 32'hca00003;
      83299: inst = 32'h24822800;
      83300: inst = 32'h10a00000;
      83301: inst = 32'hca00004;
      83302: inst = 32'h38632800;
      83303: inst = 32'h38842800;
      83304: inst = 32'h10a00001;
      83305: inst = 32'hca0456d;
      83306: inst = 32'h13e00001;
      83307: inst = 32'hfe0d96a;
      83308: inst = 32'h5be00000;
      83309: inst = 32'h8c50000;
      83310: inst = 32'h24612800;
      83311: inst = 32'h10a00000;
      83312: inst = 32'hca00003;
      83313: inst = 32'h24822800;
      83314: inst = 32'h10a00000;
      83315: inst = 32'hca00004;
      83316: inst = 32'h38632800;
      83317: inst = 32'h38842800;
      83318: inst = 32'h10a00001;
      83319: inst = 32'hca0457b;
      83320: inst = 32'h13e00001;
      83321: inst = 32'hfe0d96a;
      83322: inst = 32'h5be00000;
      83323: inst = 32'h8c50000;
      83324: inst = 32'h24612800;
      83325: inst = 32'h10a00000;
      83326: inst = 32'hca00003;
      83327: inst = 32'h24822800;
      83328: inst = 32'h10a00000;
      83329: inst = 32'hca00004;
      83330: inst = 32'h38632800;
      83331: inst = 32'h38842800;
      83332: inst = 32'h10a00001;
      83333: inst = 32'hca04589;
      83334: inst = 32'h13e00001;
      83335: inst = 32'hfe0d96a;
      83336: inst = 32'h5be00000;
      83337: inst = 32'h8c50000;
      83338: inst = 32'h24612800;
      83339: inst = 32'h10a00000;
      83340: inst = 32'hca00003;
      83341: inst = 32'h24822800;
      83342: inst = 32'h10a00000;
      83343: inst = 32'hca00004;
      83344: inst = 32'h38632800;
      83345: inst = 32'h38842800;
      83346: inst = 32'h10a00001;
      83347: inst = 32'hca04597;
      83348: inst = 32'h13e00001;
      83349: inst = 32'hfe0d96a;
      83350: inst = 32'h5be00000;
      83351: inst = 32'h8c50000;
      83352: inst = 32'h24612800;
      83353: inst = 32'h10a00000;
      83354: inst = 32'hca00003;
      83355: inst = 32'h24822800;
      83356: inst = 32'h10a00000;
      83357: inst = 32'hca00004;
      83358: inst = 32'h38632800;
      83359: inst = 32'h38842800;
      83360: inst = 32'h10a00001;
      83361: inst = 32'hca045a5;
      83362: inst = 32'h13e00001;
      83363: inst = 32'hfe0d96a;
      83364: inst = 32'h5be00000;
      83365: inst = 32'h8c50000;
      83366: inst = 32'h24612800;
      83367: inst = 32'h10a00000;
      83368: inst = 32'hca00003;
      83369: inst = 32'h24822800;
      83370: inst = 32'h10a00000;
      83371: inst = 32'hca00004;
      83372: inst = 32'h38632800;
      83373: inst = 32'h38842800;
      83374: inst = 32'h10a00001;
      83375: inst = 32'hca045b3;
      83376: inst = 32'h13e00001;
      83377: inst = 32'hfe0d96a;
      83378: inst = 32'h5be00000;
      83379: inst = 32'h8c50000;
      83380: inst = 32'h24612800;
      83381: inst = 32'h10a00000;
      83382: inst = 32'hca00003;
      83383: inst = 32'h24822800;
      83384: inst = 32'h10a00000;
      83385: inst = 32'hca00004;
      83386: inst = 32'h38632800;
      83387: inst = 32'h38842800;
      83388: inst = 32'h10a00001;
      83389: inst = 32'hca045c1;
      83390: inst = 32'h13e00001;
      83391: inst = 32'hfe0d96a;
      83392: inst = 32'h5be00000;
      83393: inst = 32'h8c50000;
      83394: inst = 32'h24612800;
      83395: inst = 32'h10a00000;
      83396: inst = 32'hca00003;
      83397: inst = 32'h24822800;
      83398: inst = 32'h10a00000;
      83399: inst = 32'hca00004;
      83400: inst = 32'h38632800;
      83401: inst = 32'h38842800;
      83402: inst = 32'h10a00001;
      83403: inst = 32'hca045cf;
      83404: inst = 32'h13e00001;
      83405: inst = 32'hfe0d96a;
      83406: inst = 32'h5be00000;
      83407: inst = 32'h8c50000;
      83408: inst = 32'h24612800;
      83409: inst = 32'h10a00000;
      83410: inst = 32'hca00003;
      83411: inst = 32'h24822800;
      83412: inst = 32'h10a00000;
      83413: inst = 32'hca00004;
      83414: inst = 32'h38632800;
      83415: inst = 32'h38842800;
      83416: inst = 32'h10a00001;
      83417: inst = 32'hca045dd;
      83418: inst = 32'h13e00001;
      83419: inst = 32'hfe0d96a;
      83420: inst = 32'h5be00000;
      83421: inst = 32'h8c50000;
      83422: inst = 32'h24612800;
      83423: inst = 32'h10a00000;
      83424: inst = 32'hca00003;
      83425: inst = 32'h24822800;
      83426: inst = 32'h10a00000;
      83427: inst = 32'hca00004;
      83428: inst = 32'h38632800;
      83429: inst = 32'h38842800;
      83430: inst = 32'h10a00001;
      83431: inst = 32'hca045eb;
      83432: inst = 32'h13e00001;
      83433: inst = 32'hfe0d96a;
      83434: inst = 32'h5be00000;
      83435: inst = 32'h8c50000;
      83436: inst = 32'h24612800;
      83437: inst = 32'h10a00000;
      83438: inst = 32'hca00003;
      83439: inst = 32'h24822800;
      83440: inst = 32'h10a00000;
      83441: inst = 32'hca00004;
      83442: inst = 32'h38632800;
      83443: inst = 32'h38842800;
      83444: inst = 32'h10a00001;
      83445: inst = 32'hca045f9;
      83446: inst = 32'h13e00001;
      83447: inst = 32'hfe0d96a;
      83448: inst = 32'h5be00000;
      83449: inst = 32'h8c50000;
      83450: inst = 32'h24612800;
      83451: inst = 32'h10a00000;
      83452: inst = 32'hca00003;
      83453: inst = 32'h24822800;
      83454: inst = 32'h10a00000;
      83455: inst = 32'hca00004;
      83456: inst = 32'h38632800;
      83457: inst = 32'h38842800;
      83458: inst = 32'h10a00001;
      83459: inst = 32'hca04607;
      83460: inst = 32'h13e00001;
      83461: inst = 32'hfe0d96a;
      83462: inst = 32'h5be00000;
      83463: inst = 32'h8c50000;
      83464: inst = 32'h24612800;
      83465: inst = 32'h10a00000;
      83466: inst = 32'hca00003;
      83467: inst = 32'h24822800;
      83468: inst = 32'h10a00000;
      83469: inst = 32'hca00004;
      83470: inst = 32'h38632800;
      83471: inst = 32'h38842800;
      83472: inst = 32'h10a00001;
      83473: inst = 32'hca04615;
      83474: inst = 32'h13e00001;
      83475: inst = 32'hfe0d96a;
      83476: inst = 32'h5be00000;
      83477: inst = 32'h8c50000;
      83478: inst = 32'h24612800;
      83479: inst = 32'h10a00000;
      83480: inst = 32'hca00003;
      83481: inst = 32'h24822800;
      83482: inst = 32'h10a00000;
      83483: inst = 32'hca00004;
      83484: inst = 32'h38632800;
      83485: inst = 32'h38842800;
      83486: inst = 32'h10a00001;
      83487: inst = 32'hca04623;
      83488: inst = 32'h13e00001;
      83489: inst = 32'hfe0d96a;
      83490: inst = 32'h5be00000;
      83491: inst = 32'h8c50000;
      83492: inst = 32'h24612800;
      83493: inst = 32'h10a00000;
      83494: inst = 32'hca00003;
      83495: inst = 32'h24822800;
      83496: inst = 32'h10a00000;
      83497: inst = 32'hca00004;
      83498: inst = 32'h38632800;
      83499: inst = 32'h38842800;
      83500: inst = 32'h10a00001;
      83501: inst = 32'hca04631;
      83502: inst = 32'h13e00001;
      83503: inst = 32'hfe0d96a;
      83504: inst = 32'h5be00000;
      83505: inst = 32'h8c50000;
      83506: inst = 32'h24612800;
      83507: inst = 32'h10a00000;
      83508: inst = 32'hca00003;
      83509: inst = 32'h24822800;
      83510: inst = 32'h10a00000;
      83511: inst = 32'hca00004;
      83512: inst = 32'h38632800;
      83513: inst = 32'h38842800;
      83514: inst = 32'h10a00001;
      83515: inst = 32'hca0463f;
      83516: inst = 32'h13e00001;
      83517: inst = 32'hfe0d96a;
      83518: inst = 32'h5be00000;
      83519: inst = 32'h8c50000;
      83520: inst = 32'h24612800;
      83521: inst = 32'h10a00000;
      83522: inst = 32'hca00003;
      83523: inst = 32'h24822800;
      83524: inst = 32'h10a00000;
      83525: inst = 32'hca00004;
      83526: inst = 32'h38632800;
      83527: inst = 32'h38842800;
      83528: inst = 32'h10a00001;
      83529: inst = 32'hca0464d;
      83530: inst = 32'h13e00001;
      83531: inst = 32'hfe0d96a;
      83532: inst = 32'h5be00000;
      83533: inst = 32'h8c50000;
      83534: inst = 32'h24612800;
      83535: inst = 32'h10a00000;
      83536: inst = 32'hca00003;
      83537: inst = 32'h24822800;
      83538: inst = 32'h10a00000;
      83539: inst = 32'hca00004;
      83540: inst = 32'h38632800;
      83541: inst = 32'h38842800;
      83542: inst = 32'h10a00001;
      83543: inst = 32'hca0465b;
      83544: inst = 32'h13e00001;
      83545: inst = 32'hfe0d96a;
      83546: inst = 32'h5be00000;
      83547: inst = 32'h8c50000;
      83548: inst = 32'h24612800;
      83549: inst = 32'h10a00000;
      83550: inst = 32'hca00003;
      83551: inst = 32'h24822800;
      83552: inst = 32'h10a00000;
      83553: inst = 32'hca00004;
      83554: inst = 32'h38632800;
      83555: inst = 32'h38842800;
      83556: inst = 32'h10a00001;
      83557: inst = 32'hca04669;
      83558: inst = 32'h13e00001;
      83559: inst = 32'hfe0d96a;
      83560: inst = 32'h5be00000;
      83561: inst = 32'h8c50000;
      83562: inst = 32'h24612800;
      83563: inst = 32'h10a00000;
      83564: inst = 32'hca00004;
      83565: inst = 32'h24822800;
      83566: inst = 32'h10a00000;
      83567: inst = 32'hca00004;
      83568: inst = 32'h38632800;
      83569: inst = 32'h38842800;
      83570: inst = 32'h10a00001;
      83571: inst = 32'hca04677;
      83572: inst = 32'h13e00001;
      83573: inst = 32'hfe0d96a;
      83574: inst = 32'h5be00000;
      83575: inst = 32'h8c50000;
      83576: inst = 32'h24612800;
      83577: inst = 32'h10a00000;
      83578: inst = 32'hca00004;
      83579: inst = 32'h24822800;
      83580: inst = 32'h10a00000;
      83581: inst = 32'hca00004;
      83582: inst = 32'h38632800;
      83583: inst = 32'h38842800;
      83584: inst = 32'h10a00001;
      83585: inst = 32'hca04685;
      83586: inst = 32'h13e00001;
      83587: inst = 32'hfe0d96a;
      83588: inst = 32'h5be00000;
      83589: inst = 32'h8c50000;
      83590: inst = 32'h24612800;
      83591: inst = 32'h10a00000;
      83592: inst = 32'hca00004;
      83593: inst = 32'h24822800;
      83594: inst = 32'h10a00000;
      83595: inst = 32'hca00004;
      83596: inst = 32'h38632800;
      83597: inst = 32'h38842800;
      83598: inst = 32'h10a00001;
      83599: inst = 32'hca04693;
      83600: inst = 32'h13e00001;
      83601: inst = 32'hfe0d96a;
      83602: inst = 32'h5be00000;
      83603: inst = 32'h8c50000;
      83604: inst = 32'h24612800;
      83605: inst = 32'h10a00000;
      83606: inst = 32'hca00004;
      83607: inst = 32'h24822800;
      83608: inst = 32'h10a00000;
      83609: inst = 32'hca00004;
      83610: inst = 32'h38632800;
      83611: inst = 32'h38842800;
      83612: inst = 32'h10a00001;
      83613: inst = 32'hca046a1;
      83614: inst = 32'h13e00001;
      83615: inst = 32'hfe0d96a;
      83616: inst = 32'h5be00000;
      83617: inst = 32'h8c50000;
      83618: inst = 32'h24612800;
      83619: inst = 32'h10a00000;
      83620: inst = 32'hca00004;
      83621: inst = 32'h24822800;
      83622: inst = 32'h10a00000;
      83623: inst = 32'hca00004;
      83624: inst = 32'h38632800;
      83625: inst = 32'h38842800;
      83626: inst = 32'h10a00001;
      83627: inst = 32'hca046af;
      83628: inst = 32'h13e00001;
      83629: inst = 32'hfe0d96a;
      83630: inst = 32'h5be00000;
      83631: inst = 32'h8c50000;
      83632: inst = 32'h24612800;
      83633: inst = 32'h10a00000;
      83634: inst = 32'hca00004;
      83635: inst = 32'h24822800;
      83636: inst = 32'h10a00000;
      83637: inst = 32'hca00004;
      83638: inst = 32'h38632800;
      83639: inst = 32'h38842800;
      83640: inst = 32'h10a00001;
      83641: inst = 32'hca046bd;
      83642: inst = 32'h13e00001;
      83643: inst = 32'hfe0d96a;
      83644: inst = 32'h5be00000;
      83645: inst = 32'h8c50000;
      83646: inst = 32'h24612800;
      83647: inst = 32'h10a00000;
      83648: inst = 32'hca00004;
      83649: inst = 32'h24822800;
      83650: inst = 32'h10a00000;
      83651: inst = 32'hca00004;
      83652: inst = 32'h38632800;
      83653: inst = 32'h38842800;
      83654: inst = 32'h10a00001;
      83655: inst = 32'hca046cb;
      83656: inst = 32'h13e00001;
      83657: inst = 32'hfe0d96a;
      83658: inst = 32'h5be00000;
      83659: inst = 32'h8c50000;
      83660: inst = 32'h24612800;
      83661: inst = 32'h10a00000;
      83662: inst = 32'hca00004;
      83663: inst = 32'h24822800;
      83664: inst = 32'h10a00000;
      83665: inst = 32'hca00004;
      83666: inst = 32'h38632800;
      83667: inst = 32'h38842800;
      83668: inst = 32'h10a00001;
      83669: inst = 32'hca046d9;
      83670: inst = 32'h13e00001;
      83671: inst = 32'hfe0d96a;
      83672: inst = 32'h5be00000;
      83673: inst = 32'h8c50000;
      83674: inst = 32'h24612800;
      83675: inst = 32'h10a00000;
      83676: inst = 32'hca00004;
      83677: inst = 32'h24822800;
      83678: inst = 32'h10a00000;
      83679: inst = 32'hca00004;
      83680: inst = 32'h38632800;
      83681: inst = 32'h38842800;
      83682: inst = 32'h10a00001;
      83683: inst = 32'hca046e7;
      83684: inst = 32'h13e00001;
      83685: inst = 32'hfe0d96a;
      83686: inst = 32'h5be00000;
      83687: inst = 32'h8c50000;
      83688: inst = 32'h24612800;
      83689: inst = 32'h10a00000;
      83690: inst = 32'hca00004;
      83691: inst = 32'h24822800;
      83692: inst = 32'h10a00000;
      83693: inst = 32'hca00004;
      83694: inst = 32'h38632800;
      83695: inst = 32'h38842800;
      83696: inst = 32'h10a00001;
      83697: inst = 32'hca046f5;
      83698: inst = 32'h13e00001;
      83699: inst = 32'hfe0d96a;
      83700: inst = 32'h5be00000;
      83701: inst = 32'h8c50000;
      83702: inst = 32'h24612800;
      83703: inst = 32'h10a00000;
      83704: inst = 32'hca00004;
      83705: inst = 32'h24822800;
      83706: inst = 32'h10a00000;
      83707: inst = 32'hca00004;
      83708: inst = 32'h38632800;
      83709: inst = 32'h38842800;
      83710: inst = 32'h10a00001;
      83711: inst = 32'hca04703;
      83712: inst = 32'h13e00001;
      83713: inst = 32'hfe0d96a;
      83714: inst = 32'h5be00000;
      83715: inst = 32'h8c50000;
      83716: inst = 32'h24612800;
      83717: inst = 32'h10a00000;
      83718: inst = 32'hca00004;
      83719: inst = 32'h24822800;
      83720: inst = 32'h10a00000;
      83721: inst = 32'hca00004;
      83722: inst = 32'h38632800;
      83723: inst = 32'h38842800;
      83724: inst = 32'h10a00001;
      83725: inst = 32'hca04711;
      83726: inst = 32'h13e00001;
      83727: inst = 32'hfe0d96a;
      83728: inst = 32'h5be00000;
      83729: inst = 32'h8c50000;
      83730: inst = 32'h24612800;
      83731: inst = 32'h10a00000;
      83732: inst = 32'hca00004;
      83733: inst = 32'h24822800;
      83734: inst = 32'h10a00000;
      83735: inst = 32'hca00004;
      83736: inst = 32'h38632800;
      83737: inst = 32'h38842800;
      83738: inst = 32'h10a00001;
      83739: inst = 32'hca0471f;
      83740: inst = 32'h13e00001;
      83741: inst = 32'hfe0d96a;
      83742: inst = 32'h5be00000;
      83743: inst = 32'h8c50000;
      83744: inst = 32'h24612800;
      83745: inst = 32'h10a00000;
      83746: inst = 32'hca00004;
      83747: inst = 32'h24822800;
      83748: inst = 32'h10a00000;
      83749: inst = 32'hca00004;
      83750: inst = 32'h38632800;
      83751: inst = 32'h38842800;
      83752: inst = 32'h10a00001;
      83753: inst = 32'hca0472d;
      83754: inst = 32'h13e00001;
      83755: inst = 32'hfe0d96a;
      83756: inst = 32'h5be00000;
      83757: inst = 32'h8c50000;
      83758: inst = 32'h24612800;
      83759: inst = 32'h10a00000;
      83760: inst = 32'hca00004;
      83761: inst = 32'h24822800;
      83762: inst = 32'h10a00000;
      83763: inst = 32'hca00004;
      83764: inst = 32'h38632800;
      83765: inst = 32'h38842800;
      83766: inst = 32'h10a00001;
      83767: inst = 32'hca0473b;
      83768: inst = 32'h13e00001;
      83769: inst = 32'hfe0d96a;
      83770: inst = 32'h5be00000;
      83771: inst = 32'h8c50000;
      83772: inst = 32'h24612800;
      83773: inst = 32'h10a00000;
      83774: inst = 32'hca00004;
      83775: inst = 32'h24822800;
      83776: inst = 32'h10a00000;
      83777: inst = 32'hca00004;
      83778: inst = 32'h38632800;
      83779: inst = 32'h38842800;
      83780: inst = 32'h10a00001;
      83781: inst = 32'hca04749;
      83782: inst = 32'h13e00001;
      83783: inst = 32'hfe0d96a;
      83784: inst = 32'h5be00000;
      83785: inst = 32'h8c50000;
      83786: inst = 32'h24612800;
      83787: inst = 32'h10a00000;
      83788: inst = 32'hca00004;
      83789: inst = 32'h24822800;
      83790: inst = 32'h10a00000;
      83791: inst = 32'hca00004;
      83792: inst = 32'h38632800;
      83793: inst = 32'h38842800;
      83794: inst = 32'h10a00001;
      83795: inst = 32'hca04757;
      83796: inst = 32'h13e00001;
      83797: inst = 32'hfe0d96a;
      83798: inst = 32'h5be00000;
      83799: inst = 32'h8c50000;
      83800: inst = 32'h24612800;
      83801: inst = 32'h10a00000;
      83802: inst = 32'hca00004;
      83803: inst = 32'h24822800;
      83804: inst = 32'h10a00000;
      83805: inst = 32'hca00004;
      83806: inst = 32'h38632800;
      83807: inst = 32'h38842800;
      83808: inst = 32'h10a00001;
      83809: inst = 32'hca04765;
      83810: inst = 32'h13e00001;
      83811: inst = 32'hfe0d96a;
      83812: inst = 32'h5be00000;
      83813: inst = 32'h8c50000;
      83814: inst = 32'h24612800;
      83815: inst = 32'h10a00000;
      83816: inst = 32'hca00004;
      83817: inst = 32'h24822800;
      83818: inst = 32'h10a00000;
      83819: inst = 32'hca00004;
      83820: inst = 32'h38632800;
      83821: inst = 32'h38842800;
      83822: inst = 32'h10a00001;
      83823: inst = 32'hca04773;
      83824: inst = 32'h13e00001;
      83825: inst = 32'hfe0d96a;
      83826: inst = 32'h5be00000;
      83827: inst = 32'h8c50000;
      83828: inst = 32'h24612800;
      83829: inst = 32'h10a00000;
      83830: inst = 32'hca00004;
      83831: inst = 32'h24822800;
      83832: inst = 32'h10a00000;
      83833: inst = 32'hca00004;
      83834: inst = 32'h38632800;
      83835: inst = 32'h38842800;
      83836: inst = 32'h10a00001;
      83837: inst = 32'hca04781;
      83838: inst = 32'h13e00001;
      83839: inst = 32'hfe0d96a;
      83840: inst = 32'h5be00000;
      83841: inst = 32'h8c50000;
      83842: inst = 32'h24612800;
      83843: inst = 32'h10a00000;
      83844: inst = 32'hca00004;
      83845: inst = 32'h24822800;
      83846: inst = 32'h10a00000;
      83847: inst = 32'hca00004;
      83848: inst = 32'h38632800;
      83849: inst = 32'h38842800;
      83850: inst = 32'h10a00001;
      83851: inst = 32'hca0478f;
      83852: inst = 32'h13e00001;
      83853: inst = 32'hfe0d96a;
      83854: inst = 32'h5be00000;
      83855: inst = 32'h8c50000;
      83856: inst = 32'h24612800;
      83857: inst = 32'h10a00000;
      83858: inst = 32'hca00004;
      83859: inst = 32'h24822800;
      83860: inst = 32'h10a00000;
      83861: inst = 32'hca00004;
      83862: inst = 32'h38632800;
      83863: inst = 32'h38842800;
      83864: inst = 32'h10a00001;
      83865: inst = 32'hca0479d;
      83866: inst = 32'h13e00001;
      83867: inst = 32'hfe0d96a;
      83868: inst = 32'h5be00000;
      83869: inst = 32'h8c50000;
      83870: inst = 32'h24612800;
      83871: inst = 32'h10a00000;
      83872: inst = 32'hca00004;
      83873: inst = 32'h24822800;
      83874: inst = 32'h10a00000;
      83875: inst = 32'hca00004;
      83876: inst = 32'h38632800;
      83877: inst = 32'h38842800;
      83878: inst = 32'h10a00001;
      83879: inst = 32'hca047ab;
      83880: inst = 32'h13e00001;
      83881: inst = 32'hfe0d96a;
      83882: inst = 32'h5be00000;
      83883: inst = 32'h8c50000;
      83884: inst = 32'h24612800;
      83885: inst = 32'h10a00000;
      83886: inst = 32'hca00004;
      83887: inst = 32'h24822800;
      83888: inst = 32'h10a00000;
      83889: inst = 32'hca00004;
      83890: inst = 32'h38632800;
      83891: inst = 32'h38842800;
      83892: inst = 32'h10a00001;
      83893: inst = 32'hca047b9;
      83894: inst = 32'h13e00001;
      83895: inst = 32'hfe0d96a;
      83896: inst = 32'h5be00000;
      83897: inst = 32'h8c50000;
      83898: inst = 32'h24612800;
      83899: inst = 32'h10a00000;
      83900: inst = 32'hca00004;
      83901: inst = 32'h24822800;
      83902: inst = 32'h10a00000;
      83903: inst = 32'hca00004;
      83904: inst = 32'h38632800;
      83905: inst = 32'h38842800;
      83906: inst = 32'h10a00001;
      83907: inst = 32'hca047c7;
      83908: inst = 32'h13e00001;
      83909: inst = 32'hfe0d96a;
      83910: inst = 32'h5be00000;
      83911: inst = 32'h8c50000;
      83912: inst = 32'h24612800;
      83913: inst = 32'h10a00000;
      83914: inst = 32'hca00004;
      83915: inst = 32'h24822800;
      83916: inst = 32'h10a00000;
      83917: inst = 32'hca00004;
      83918: inst = 32'h38632800;
      83919: inst = 32'h38842800;
      83920: inst = 32'h10a00001;
      83921: inst = 32'hca047d5;
      83922: inst = 32'h13e00001;
      83923: inst = 32'hfe0d96a;
      83924: inst = 32'h5be00000;
      83925: inst = 32'h8c50000;
      83926: inst = 32'h24612800;
      83927: inst = 32'h10a00000;
      83928: inst = 32'hca00004;
      83929: inst = 32'h24822800;
      83930: inst = 32'h10a00000;
      83931: inst = 32'hca00004;
      83932: inst = 32'h38632800;
      83933: inst = 32'h38842800;
      83934: inst = 32'h10a00001;
      83935: inst = 32'hca047e3;
      83936: inst = 32'h13e00001;
      83937: inst = 32'hfe0d96a;
      83938: inst = 32'h5be00000;
      83939: inst = 32'h8c50000;
      83940: inst = 32'h24612800;
      83941: inst = 32'h10a00000;
      83942: inst = 32'hca00004;
      83943: inst = 32'h24822800;
      83944: inst = 32'h10a00000;
      83945: inst = 32'hca00004;
      83946: inst = 32'h38632800;
      83947: inst = 32'h38842800;
      83948: inst = 32'h10a00001;
      83949: inst = 32'hca047f1;
      83950: inst = 32'h13e00001;
      83951: inst = 32'hfe0d96a;
      83952: inst = 32'h5be00000;
      83953: inst = 32'h8c50000;
      83954: inst = 32'h24612800;
      83955: inst = 32'h10a00000;
      83956: inst = 32'hca00004;
      83957: inst = 32'h24822800;
      83958: inst = 32'h10a00000;
      83959: inst = 32'hca00004;
      83960: inst = 32'h38632800;
      83961: inst = 32'h38842800;
      83962: inst = 32'h10a00001;
      83963: inst = 32'hca047ff;
      83964: inst = 32'h13e00001;
      83965: inst = 32'hfe0d96a;
      83966: inst = 32'h5be00000;
      83967: inst = 32'h8c50000;
      83968: inst = 32'h24612800;
      83969: inst = 32'h10a00000;
      83970: inst = 32'hca00004;
      83971: inst = 32'h24822800;
      83972: inst = 32'h10a00000;
      83973: inst = 32'hca00004;
      83974: inst = 32'h38632800;
      83975: inst = 32'h38842800;
      83976: inst = 32'h10a00001;
      83977: inst = 32'hca0480d;
      83978: inst = 32'h13e00001;
      83979: inst = 32'hfe0d96a;
      83980: inst = 32'h5be00000;
      83981: inst = 32'h8c50000;
      83982: inst = 32'h24612800;
      83983: inst = 32'h10a00000;
      83984: inst = 32'hca00004;
      83985: inst = 32'h24822800;
      83986: inst = 32'h10a00000;
      83987: inst = 32'hca00004;
      83988: inst = 32'h38632800;
      83989: inst = 32'h38842800;
      83990: inst = 32'h10a00001;
      83991: inst = 32'hca0481b;
      83992: inst = 32'h13e00001;
      83993: inst = 32'hfe0d96a;
      83994: inst = 32'h5be00000;
      83995: inst = 32'h8c50000;
      83996: inst = 32'h24612800;
      83997: inst = 32'h10a00000;
      83998: inst = 32'hca00004;
      83999: inst = 32'h24822800;
      84000: inst = 32'h10a00000;
      84001: inst = 32'hca00004;
      84002: inst = 32'h38632800;
      84003: inst = 32'h38842800;
      84004: inst = 32'h10a00001;
      84005: inst = 32'hca04829;
      84006: inst = 32'h13e00001;
      84007: inst = 32'hfe0d96a;
      84008: inst = 32'h5be00000;
      84009: inst = 32'h8c50000;
      84010: inst = 32'h24612800;
      84011: inst = 32'h10a00000;
      84012: inst = 32'hca00004;
      84013: inst = 32'h24822800;
      84014: inst = 32'h10a00000;
      84015: inst = 32'hca00004;
      84016: inst = 32'h38632800;
      84017: inst = 32'h38842800;
      84018: inst = 32'h10a00001;
      84019: inst = 32'hca04837;
      84020: inst = 32'h13e00001;
      84021: inst = 32'hfe0d96a;
      84022: inst = 32'h5be00000;
      84023: inst = 32'h8c50000;
      84024: inst = 32'h24612800;
      84025: inst = 32'h10a00000;
      84026: inst = 32'hca00004;
      84027: inst = 32'h24822800;
      84028: inst = 32'h10a00000;
      84029: inst = 32'hca00004;
      84030: inst = 32'h38632800;
      84031: inst = 32'h38842800;
      84032: inst = 32'h10a00001;
      84033: inst = 32'hca04845;
      84034: inst = 32'h13e00001;
      84035: inst = 32'hfe0d96a;
      84036: inst = 32'h5be00000;
      84037: inst = 32'h8c50000;
      84038: inst = 32'h24612800;
      84039: inst = 32'h10a00000;
      84040: inst = 32'hca00004;
      84041: inst = 32'h24822800;
      84042: inst = 32'h10a00000;
      84043: inst = 32'hca00004;
      84044: inst = 32'h38632800;
      84045: inst = 32'h38842800;
      84046: inst = 32'h10a00001;
      84047: inst = 32'hca04853;
      84048: inst = 32'h13e00001;
      84049: inst = 32'hfe0d96a;
      84050: inst = 32'h5be00000;
      84051: inst = 32'h8c50000;
      84052: inst = 32'h24612800;
      84053: inst = 32'h10a00000;
      84054: inst = 32'hca00004;
      84055: inst = 32'h24822800;
      84056: inst = 32'h10a00000;
      84057: inst = 32'hca00004;
      84058: inst = 32'h38632800;
      84059: inst = 32'h38842800;
      84060: inst = 32'h10a00001;
      84061: inst = 32'hca04861;
      84062: inst = 32'h13e00001;
      84063: inst = 32'hfe0d96a;
      84064: inst = 32'h5be00000;
      84065: inst = 32'h8c50000;
      84066: inst = 32'h24612800;
      84067: inst = 32'h10a00000;
      84068: inst = 32'hca00004;
      84069: inst = 32'h24822800;
      84070: inst = 32'h10a00000;
      84071: inst = 32'hca00004;
      84072: inst = 32'h38632800;
      84073: inst = 32'h38842800;
      84074: inst = 32'h10a00001;
      84075: inst = 32'hca0486f;
      84076: inst = 32'h13e00001;
      84077: inst = 32'hfe0d96a;
      84078: inst = 32'h5be00000;
      84079: inst = 32'h8c50000;
      84080: inst = 32'h24612800;
      84081: inst = 32'h10a00000;
      84082: inst = 32'hca00004;
      84083: inst = 32'h24822800;
      84084: inst = 32'h10a00000;
      84085: inst = 32'hca00004;
      84086: inst = 32'h38632800;
      84087: inst = 32'h38842800;
      84088: inst = 32'h10a00001;
      84089: inst = 32'hca0487d;
      84090: inst = 32'h13e00001;
      84091: inst = 32'hfe0d96a;
      84092: inst = 32'h5be00000;
      84093: inst = 32'h8c50000;
      84094: inst = 32'h24612800;
      84095: inst = 32'h10a00000;
      84096: inst = 32'hca00004;
      84097: inst = 32'h24822800;
      84098: inst = 32'h10a00000;
      84099: inst = 32'hca00004;
      84100: inst = 32'h38632800;
      84101: inst = 32'h38842800;
      84102: inst = 32'h10a00001;
      84103: inst = 32'hca0488b;
      84104: inst = 32'h13e00001;
      84105: inst = 32'hfe0d96a;
      84106: inst = 32'h5be00000;
      84107: inst = 32'h8c50000;
      84108: inst = 32'h24612800;
      84109: inst = 32'h10a00000;
      84110: inst = 32'hca00004;
      84111: inst = 32'h24822800;
      84112: inst = 32'h10a00000;
      84113: inst = 32'hca00004;
      84114: inst = 32'h38632800;
      84115: inst = 32'h38842800;
      84116: inst = 32'h10a00001;
      84117: inst = 32'hca04899;
      84118: inst = 32'h13e00001;
      84119: inst = 32'hfe0d96a;
      84120: inst = 32'h5be00000;
      84121: inst = 32'h8c50000;
      84122: inst = 32'h24612800;
      84123: inst = 32'h10a00000;
      84124: inst = 32'hca00004;
      84125: inst = 32'h24822800;
      84126: inst = 32'h10a00000;
      84127: inst = 32'hca00004;
      84128: inst = 32'h38632800;
      84129: inst = 32'h38842800;
      84130: inst = 32'h10a00001;
      84131: inst = 32'hca048a7;
      84132: inst = 32'h13e00001;
      84133: inst = 32'hfe0d96a;
      84134: inst = 32'h5be00000;
      84135: inst = 32'h8c50000;
      84136: inst = 32'h24612800;
      84137: inst = 32'h10a00000;
      84138: inst = 32'hca00004;
      84139: inst = 32'h24822800;
      84140: inst = 32'h10a00000;
      84141: inst = 32'hca00004;
      84142: inst = 32'h38632800;
      84143: inst = 32'h38842800;
      84144: inst = 32'h10a00001;
      84145: inst = 32'hca048b5;
      84146: inst = 32'h13e00001;
      84147: inst = 32'hfe0d96a;
      84148: inst = 32'h5be00000;
      84149: inst = 32'h8c50000;
      84150: inst = 32'h24612800;
      84151: inst = 32'h10a00000;
      84152: inst = 32'hca00004;
      84153: inst = 32'h24822800;
      84154: inst = 32'h10a00000;
      84155: inst = 32'hca00004;
      84156: inst = 32'h38632800;
      84157: inst = 32'h38842800;
      84158: inst = 32'h10a00001;
      84159: inst = 32'hca048c3;
      84160: inst = 32'h13e00001;
      84161: inst = 32'hfe0d96a;
      84162: inst = 32'h5be00000;
      84163: inst = 32'h8c50000;
      84164: inst = 32'h24612800;
      84165: inst = 32'h10a00000;
      84166: inst = 32'hca00004;
      84167: inst = 32'h24822800;
      84168: inst = 32'h10a00000;
      84169: inst = 32'hca00004;
      84170: inst = 32'h38632800;
      84171: inst = 32'h38842800;
      84172: inst = 32'h10a00001;
      84173: inst = 32'hca048d1;
      84174: inst = 32'h13e00001;
      84175: inst = 32'hfe0d96a;
      84176: inst = 32'h5be00000;
      84177: inst = 32'h8c50000;
      84178: inst = 32'h24612800;
      84179: inst = 32'h10a00000;
      84180: inst = 32'hca00004;
      84181: inst = 32'h24822800;
      84182: inst = 32'h10a00000;
      84183: inst = 32'hca00004;
      84184: inst = 32'h38632800;
      84185: inst = 32'h38842800;
      84186: inst = 32'h10a00001;
      84187: inst = 32'hca048df;
      84188: inst = 32'h13e00001;
      84189: inst = 32'hfe0d96a;
      84190: inst = 32'h5be00000;
      84191: inst = 32'h8c50000;
      84192: inst = 32'h24612800;
      84193: inst = 32'h10a00000;
      84194: inst = 32'hca00004;
      84195: inst = 32'h24822800;
      84196: inst = 32'h10a00000;
      84197: inst = 32'hca00004;
      84198: inst = 32'h38632800;
      84199: inst = 32'h38842800;
      84200: inst = 32'h10a00001;
      84201: inst = 32'hca048ed;
      84202: inst = 32'h13e00001;
      84203: inst = 32'hfe0d96a;
      84204: inst = 32'h5be00000;
      84205: inst = 32'h8c50000;
      84206: inst = 32'h24612800;
      84207: inst = 32'h10a00000;
      84208: inst = 32'hca00004;
      84209: inst = 32'h24822800;
      84210: inst = 32'h10a00000;
      84211: inst = 32'hca00004;
      84212: inst = 32'h38632800;
      84213: inst = 32'h38842800;
      84214: inst = 32'h10a00001;
      84215: inst = 32'hca048fb;
      84216: inst = 32'h13e00001;
      84217: inst = 32'hfe0d96a;
      84218: inst = 32'h5be00000;
      84219: inst = 32'h8c50000;
      84220: inst = 32'h24612800;
      84221: inst = 32'h10a00000;
      84222: inst = 32'hca00004;
      84223: inst = 32'h24822800;
      84224: inst = 32'h10a00000;
      84225: inst = 32'hca00004;
      84226: inst = 32'h38632800;
      84227: inst = 32'h38842800;
      84228: inst = 32'h10a00001;
      84229: inst = 32'hca04909;
      84230: inst = 32'h13e00001;
      84231: inst = 32'hfe0d96a;
      84232: inst = 32'h5be00000;
      84233: inst = 32'h8c50000;
      84234: inst = 32'h24612800;
      84235: inst = 32'h10a00000;
      84236: inst = 32'hca00004;
      84237: inst = 32'h24822800;
      84238: inst = 32'h10a00000;
      84239: inst = 32'hca00004;
      84240: inst = 32'h38632800;
      84241: inst = 32'h38842800;
      84242: inst = 32'h10a00001;
      84243: inst = 32'hca04917;
      84244: inst = 32'h13e00001;
      84245: inst = 32'hfe0d96a;
      84246: inst = 32'h5be00000;
      84247: inst = 32'h8c50000;
      84248: inst = 32'h24612800;
      84249: inst = 32'h10a00000;
      84250: inst = 32'hca00004;
      84251: inst = 32'h24822800;
      84252: inst = 32'h10a00000;
      84253: inst = 32'hca00004;
      84254: inst = 32'h38632800;
      84255: inst = 32'h38842800;
      84256: inst = 32'h10a00001;
      84257: inst = 32'hca04925;
      84258: inst = 32'h13e00001;
      84259: inst = 32'hfe0d96a;
      84260: inst = 32'h5be00000;
      84261: inst = 32'h8c50000;
      84262: inst = 32'h24612800;
      84263: inst = 32'h10a00000;
      84264: inst = 32'hca00004;
      84265: inst = 32'h24822800;
      84266: inst = 32'h10a00000;
      84267: inst = 32'hca00004;
      84268: inst = 32'h38632800;
      84269: inst = 32'h38842800;
      84270: inst = 32'h10a00001;
      84271: inst = 32'hca04933;
      84272: inst = 32'h13e00001;
      84273: inst = 32'hfe0d96a;
      84274: inst = 32'h5be00000;
      84275: inst = 32'h8c50000;
      84276: inst = 32'h24612800;
      84277: inst = 32'h10a00000;
      84278: inst = 32'hca00004;
      84279: inst = 32'h24822800;
      84280: inst = 32'h10a00000;
      84281: inst = 32'hca00004;
      84282: inst = 32'h38632800;
      84283: inst = 32'h38842800;
      84284: inst = 32'h10a00001;
      84285: inst = 32'hca04941;
      84286: inst = 32'h13e00001;
      84287: inst = 32'hfe0d96a;
      84288: inst = 32'h5be00000;
      84289: inst = 32'h8c50000;
      84290: inst = 32'h24612800;
      84291: inst = 32'h10a00000;
      84292: inst = 32'hca00004;
      84293: inst = 32'h24822800;
      84294: inst = 32'h10a00000;
      84295: inst = 32'hca00004;
      84296: inst = 32'h38632800;
      84297: inst = 32'h38842800;
      84298: inst = 32'h10a00001;
      84299: inst = 32'hca0494f;
      84300: inst = 32'h13e00001;
      84301: inst = 32'hfe0d96a;
      84302: inst = 32'h5be00000;
      84303: inst = 32'h8c50000;
      84304: inst = 32'h24612800;
      84305: inst = 32'h10a00000;
      84306: inst = 32'hca00004;
      84307: inst = 32'h24822800;
      84308: inst = 32'h10a00000;
      84309: inst = 32'hca00004;
      84310: inst = 32'h38632800;
      84311: inst = 32'h38842800;
      84312: inst = 32'h10a00001;
      84313: inst = 32'hca0495d;
      84314: inst = 32'h13e00001;
      84315: inst = 32'hfe0d96a;
      84316: inst = 32'h5be00000;
      84317: inst = 32'h8c50000;
      84318: inst = 32'h24612800;
      84319: inst = 32'h10a00000;
      84320: inst = 32'hca00004;
      84321: inst = 32'h24822800;
      84322: inst = 32'h10a00000;
      84323: inst = 32'hca00004;
      84324: inst = 32'h38632800;
      84325: inst = 32'h38842800;
      84326: inst = 32'h10a00001;
      84327: inst = 32'hca0496b;
      84328: inst = 32'h13e00001;
      84329: inst = 32'hfe0d96a;
      84330: inst = 32'h5be00000;
      84331: inst = 32'h8c50000;
      84332: inst = 32'h24612800;
      84333: inst = 32'h10a00000;
      84334: inst = 32'hca00004;
      84335: inst = 32'h24822800;
      84336: inst = 32'h10a00000;
      84337: inst = 32'hca00004;
      84338: inst = 32'h38632800;
      84339: inst = 32'h38842800;
      84340: inst = 32'h10a00001;
      84341: inst = 32'hca04979;
      84342: inst = 32'h13e00001;
      84343: inst = 32'hfe0d96a;
      84344: inst = 32'h5be00000;
      84345: inst = 32'h8c50000;
      84346: inst = 32'h24612800;
      84347: inst = 32'h10a00000;
      84348: inst = 32'hca00004;
      84349: inst = 32'h24822800;
      84350: inst = 32'h10a00000;
      84351: inst = 32'hca00004;
      84352: inst = 32'h38632800;
      84353: inst = 32'h38842800;
      84354: inst = 32'h10a00001;
      84355: inst = 32'hca04987;
      84356: inst = 32'h13e00001;
      84357: inst = 32'hfe0d96a;
      84358: inst = 32'h5be00000;
      84359: inst = 32'h8c50000;
      84360: inst = 32'h24612800;
      84361: inst = 32'h10a00000;
      84362: inst = 32'hca00004;
      84363: inst = 32'h24822800;
      84364: inst = 32'h10a00000;
      84365: inst = 32'hca00004;
      84366: inst = 32'h38632800;
      84367: inst = 32'h38842800;
      84368: inst = 32'h10a00001;
      84369: inst = 32'hca04995;
      84370: inst = 32'h13e00001;
      84371: inst = 32'hfe0d96a;
      84372: inst = 32'h5be00000;
      84373: inst = 32'h8c50000;
      84374: inst = 32'h24612800;
      84375: inst = 32'h10a00000;
      84376: inst = 32'hca00004;
      84377: inst = 32'h24822800;
      84378: inst = 32'h10a00000;
      84379: inst = 32'hca00004;
      84380: inst = 32'h38632800;
      84381: inst = 32'h38842800;
      84382: inst = 32'h10a00001;
      84383: inst = 32'hca049a3;
      84384: inst = 32'h13e00001;
      84385: inst = 32'hfe0d96a;
      84386: inst = 32'h5be00000;
      84387: inst = 32'h8c50000;
      84388: inst = 32'h24612800;
      84389: inst = 32'h10a00000;
      84390: inst = 32'hca00004;
      84391: inst = 32'h24822800;
      84392: inst = 32'h10a00000;
      84393: inst = 32'hca00004;
      84394: inst = 32'h38632800;
      84395: inst = 32'h38842800;
      84396: inst = 32'h10a00001;
      84397: inst = 32'hca049b1;
      84398: inst = 32'h13e00001;
      84399: inst = 32'hfe0d96a;
      84400: inst = 32'h5be00000;
      84401: inst = 32'h8c50000;
      84402: inst = 32'h24612800;
      84403: inst = 32'h10a00000;
      84404: inst = 32'hca00004;
      84405: inst = 32'h24822800;
      84406: inst = 32'h10a00000;
      84407: inst = 32'hca00004;
      84408: inst = 32'h38632800;
      84409: inst = 32'h38842800;
      84410: inst = 32'h10a00001;
      84411: inst = 32'hca049bf;
      84412: inst = 32'h13e00001;
      84413: inst = 32'hfe0d96a;
      84414: inst = 32'h5be00000;
      84415: inst = 32'h8c50000;
      84416: inst = 32'h24612800;
      84417: inst = 32'h10a00000;
      84418: inst = 32'hca00004;
      84419: inst = 32'h24822800;
      84420: inst = 32'h10a00000;
      84421: inst = 32'hca00004;
      84422: inst = 32'h38632800;
      84423: inst = 32'h38842800;
      84424: inst = 32'h10a00001;
      84425: inst = 32'hca049cd;
      84426: inst = 32'h13e00001;
      84427: inst = 32'hfe0d96a;
      84428: inst = 32'h5be00000;
      84429: inst = 32'h8c50000;
      84430: inst = 32'h24612800;
      84431: inst = 32'h10a00000;
      84432: inst = 32'hca00004;
      84433: inst = 32'h24822800;
      84434: inst = 32'h10a00000;
      84435: inst = 32'hca00004;
      84436: inst = 32'h38632800;
      84437: inst = 32'h38842800;
      84438: inst = 32'h10a00001;
      84439: inst = 32'hca049db;
      84440: inst = 32'h13e00001;
      84441: inst = 32'hfe0d96a;
      84442: inst = 32'h5be00000;
      84443: inst = 32'h8c50000;
      84444: inst = 32'h24612800;
      84445: inst = 32'h10a00000;
      84446: inst = 32'hca00004;
      84447: inst = 32'h24822800;
      84448: inst = 32'h10a00000;
      84449: inst = 32'hca00004;
      84450: inst = 32'h38632800;
      84451: inst = 32'h38842800;
      84452: inst = 32'h10a00001;
      84453: inst = 32'hca049e9;
      84454: inst = 32'h13e00001;
      84455: inst = 32'hfe0d96a;
      84456: inst = 32'h5be00000;
      84457: inst = 32'h8c50000;
      84458: inst = 32'h24612800;
      84459: inst = 32'h10a00000;
      84460: inst = 32'hca00004;
      84461: inst = 32'h24822800;
      84462: inst = 32'h10a00000;
      84463: inst = 32'hca00004;
      84464: inst = 32'h38632800;
      84465: inst = 32'h38842800;
      84466: inst = 32'h10a00001;
      84467: inst = 32'hca049f7;
      84468: inst = 32'h13e00001;
      84469: inst = 32'hfe0d96a;
      84470: inst = 32'h5be00000;
      84471: inst = 32'h8c50000;
      84472: inst = 32'h24612800;
      84473: inst = 32'h10a00000;
      84474: inst = 32'hca00004;
      84475: inst = 32'h24822800;
      84476: inst = 32'h10a00000;
      84477: inst = 32'hca00004;
      84478: inst = 32'h38632800;
      84479: inst = 32'h38842800;
      84480: inst = 32'h10a00001;
      84481: inst = 32'hca04a05;
      84482: inst = 32'h13e00001;
      84483: inst = 32'hfe0d96a;
      84484: inst = 32'h5be00000;
      84485: inst = 32'h8c50000;
      84486: inst = 32'h24612800;
      84487: inst = 32'h10a00000;
      84488: inst = 32'hca00004;
      84489: inst = 32'h24822800;
      84490: inst = 32'h10a00000;
      84491: inst = 32'hca00004;
      84492: inst = 32'h38632800;
      84493: inst = 32'h38842800;
      84494: inst = 32'h10a00001;
      84495: inst = 32'hca04a13;
      84496: inst = 32'h13e00001;
      84497: inst = 32'hfe0d96a;
      84498: inst = 32'h5be00000;
      84499: inst = 32'h8c50000;
      84500: inst = 32'h24612800;
      84501: inst = 32'h10a00000;
      84502: inst = 32'hca00004;
      84503: inst = 32'h24822800;
      84504: inst = 32'h10a00000;
      84505: inst = 32'hca00004;
      84506: inst = 32'h38632800;
      84507: inst = 32'h38842800;
      84508: inst = 32'h10a00001;
      84509: inst = 32'hca04a21;
      84510: inst = 32'h13e00001;
      84511: inst = 32'hfe0d96a;
      84512: inst = 32'h5be00000;
      84513: inst = 32'h8c50000;
      84514: inst = 32'h24612800;
      84515: inst = 32'h10a00000;
      84516: inst = 32'hca00004;
      84517: inst = 32'h24822800;
      84518: inst = 32'h10a00000;
      84519: inst = 32'hca00004;
      84520: inst = 32'h38632800;
      84521: inst = 32'h38842800;
      84522: inst = 32'h10a00001;
      84523: inst = 32'hca04a2f;
      84524: inst = 32'h13e00001;
      84525: inst = 32'hfe0d96a;
      84526: inst = 32'h5be00000;
      84527: inst = 32'h8c50000;
      84528: inst = 32'h24612800;
      84529: inst = 32'h10a00000;
      84530: inst = 32'hca00004;
      84531: inst = 32'h24822800;
      84532: inst = 32'h10a00000;
      84533: inst = 32'hca00004;
      84534: inst = 32'h38632800;
      84535: inst = 32'h38842800;
      84536: inst = 32'h10a00001;
      84537: inst = 32'hca04a3d;
      84538: inst = 32'h13e00001;
      84539: inst = 32'hfe0d96a;
      84540: inst = 32'h5be00000;
      84541: inst = 32'h8c50000;
      84542: inst = 32'h24612800;
      84543: inst = 32'h10a00000;
      84544: inst = 32'hca00004;
      84545: inst = 32'h24822800;
      84546: inst = 32'h10a00000;
      84547: inst = 32'hca00004;
      84548: inst = 32'h38632800;
      84549: inst = 32'h38842800;
      84550: inst = 32'h10a00001;
      84551: inst = 32'hca04a4b;
      84552: inst = 32'h13e00001;
      84553: inst = 32'hfe0d96a;
      84554: inst = 32'h5be00000;
      84555: inst = 32'h8c50000;
      84556: inst = 32'h24612800;
      84557: inst = 32'h10a00000;
      84558: inst = 32'hca00004;
      84559: inst = 32'h24822800;
      84560: inst = 32'h10a00000;
      84561: inst = 32'hca00004;
      84562: inst = 32'h38632800;
      84563: inst = 32'h38842800;
      84564: inst = 32'h10a00001;
      84565: inst = 32'hca04a59;
      84566: inst = 32'h13e00001;
      84567: inst = 32'hfe0d96a;
      84568: inst = 32'h5be00000;
      84569: inst = 32'h8c50000;
      84570: inst = 32'h24612800;
      84571: inst = 32'h10a00000;
      84572: inst = 32'hca00004;
      84573: inst = 32'h24822800;
      84574: inst = 32'h10a00000;
      84575: inst = 32'hca00004;
      84576: inst = 32'h38632800;
      84577: inst = 32'h38842800;
      84578: inst = 32'h10a00001;
      84579: inst = 32'hca04a67;
      84580: inst = 32'h13e00001;
      84581: inst = 32'hfe0d96a;
      84582: inst = 32'h5be00000;
      84583: inst = 32'h8c50000;
      84584: inst = 32'h24612800;
      84585: inst = 32'h10a00000;
      84586: inst = 32'hca00004;
      84587: inst = 32'h24822800;
      84588: inst = 32'h10a00000;
      84589: inst = 32'hca00004;
      84590: inst = 32'h38632800;
      84591: inst = 32'h38842800;
      84592: inst = 32'h10a00001;
      84593: inst = 32'hca04a75;
      84594: inst = 32'h13e00001;
      84595: inst = 32'hfe0d96a;
      84596: inst = 32'h5be00000;
      84597: inst = 32'h8c50000;
      84598: inst = 32'h24612800;
      84599: inst = 32'h10a00000;
      84600: inst = 32'hca00004;
      84601: inst = 32'h24822800;
      84602: inst = 32'h10a00000;
      84603: inst = 32'hca00004;
      84604: inst = 32'h38632800;
      84605: inst = 32'h38842800;
      84606: inst = 32'h10a00001;
      84607: inst = 32'hca04a83;
      84608: inst = 32'h13e00001;
      84609: inst = 32'hfe0d96a;
      84610: inst = 32'h5be00000;
      84611: inst = 32'h8c50000;
      84612: inst = 32'h24612800;
      84613: inst = 32'h10a00000;
      84614: inst = 32'hca00004;
      84615: inst = 32'h24822800;
      84616: inst = 32'h10a00000;
      84617: inst = 32'hca00004;
      84618: inst = 32'h38632800;
      84619: inst = 32'h38842800;
      84620: inst = 32'h10a00001;
      84621: inst = 32'hca04a91;
      84622: inst = 32'h13e00001;
      84623: inst = 32'hfe0d96a;
      84624: inst = 32'h5be00000;
      84625: inst = 32'h8c50000;
      84626: inst = 32'h24612800;
      84627: inst = 32'h10a00000;
      84628: inst = 32'hca00004;
      84629: inst = 32'h24822800;
      84630: inst = 32'h10a00000;
      84631: inst = 32'hca00004;
      84632: inst = 32'h38632800;
      84633: inst = 32'h38842800;
      84634: inst = 32'h10a00001;
      84635: inst = 32'hca04a9f;
      84636: inst = 32'h13e00001;
      84637: inst = 32'hfe0d96a;
      84638: inst = 32'h5be00000;
      84639: inst = 32'h8c50000;
      84640: inst = 32'h24612800;
      84641: inst = 32'h10a00000;
      84642: inst = 32'hca00004;
      84643: inst = 32'h24822800;
      84644: inst = 32'h10a00000;
      84645: inst = 32'hca00004;
      84646: inst = 32'h38632800;
      84647: inst = 32'h38842800;
      84648: inst = 32'h10a00001;
      84649: inst = 32'hca04aad;
      84650: inst = 32'h13e00001;
      84651: inst = 32'hfe0d96a;
      84652: inst = 32'h5be00000;
      84653: inst = 32'h8c50000;
      84654: inst = 32'h24612800;
      84655: inst = 32'h10a00000;
      84656: inst = 32'hca00004;
      84657: inst = 32'h24822800;
      84658: inst = 32'h10a00000;
      84659: inst = 32'hca00004;
      84660: inst = 32'h38632800;
      84661: inst = 32'h38842800;
      84662: inst = 32'h10a00001;
      84663: inst = 32'hca04abb;
      84664: inst = 32'h13e00001;
      84665: inst = 32'hfe0d96a;
      84666: inst = 32'h5be00000;
      84667: inst = 32'h8c50000;
      84668: inst = 32'h24612800;
      84669: inst = 32'h10a00000;
      84670: inst = 32'hca00004;
      84671: inst = 32'h24822800;
      84672: inst = 32'h10a00000;
      84673: inst = 32'hca00004;
      84674: inst = 32'h38632800;
      84675: inst = 32'h38842800;
      84676: inst = 32'h10a00001;
      84677: inst = 32'hca04ac9;
      84678: inst = 32'h13e00001;
      84679: inst = 32'hfe0d96a;
      84680: inst = 32'h5be00000;
      84681: inst = 32'h8c50000;
      84682: inst = 32'h24612800;
      84683: inst = 32'h10a00000;
      84684: inst = 32'hca00004;
      84685: inst = 32'h24822800;
      84686: inst = 32'h10a00000;
      84687: inst = 32'hca00004;
      84688: inst = 32'h38632800;
      84689: inst = 32'h38842800;
      84690: inst = 32'h10a00001;
      84691: inst = 32'hca04ad7;
      84692: inst = 32'h13e00001;
      84693: inst = 32'hfe0d96a;
      84694: inst = 32'h5be00000;
      84695: inst = 32'h8c50000;
      84696: inst = 32'h24612800;
      84697: inst = 32'h10a00000;
      84698: inst = 32'hca00004;
      84699: inst = 32'h24822800;
      84700: inst = 32'h10a00000;
      84701: inst = 32'hca00004;
      84702: inst = 32'h38632800;
      84703: inst = 32'h38842800;
      84704: inst = 32'h10a00001;
      84705: inst = 32'hca04ae5;
      84706: inst = 32'h13e00001;
      84707: inst = 32'hfe0d96a;
      84708: inst = 32'h5be00000;
      84709: inst = 32'h8c50000;
      84710: inst = 32'h24612800;
      84711: inst = 32'h10a00000;
      84712: inst = 32'hca00004;
      84713: inst = 32'h24822800;
      84714: inst = 32'h10a00000;
      84715: inst = 32'hca00004;
      84716: inst = 32'h38632800;
      84717: inst = 32'h38842800;
      84718: inst = 32'h10a00001;
      84719: inst = 32'hca04af3;
      84720: inst = 32'h13e00001;
      84721: inst = 32'hfe0d96a;
      84722: inst = 32'h5be00000;
      84723: inst = 32'h8c50000;
      84724: inst = 32'h24612800;
      84725: inst = 32'h10a00000;
      84726: inst = 32'hca00004;
      84727: inst = 32'h24822800;
      84728: inst = 32'h10a00000;
      84729: inst = 32'hca00004;
      84730: inst = 32'h38632800;
      84731: inst = 32'h38842800;
      84732: inst = 32'h10a00001;
      84733: inst = 32'hca04b01;
      84734: inst = 32'h13e00001;
      84735: inst = 32'hfe0d96a;
      84736: inst = 32'h5be00000;
      84737: inst = 32'h8c50000;
      84738: inst = 32'h24612800;
      84739: inst = 32'h10a00000;
      84740: inst = 32'hca00004;
      84741: inst = 32'h24822800;
      84742: inst = 32'h10a00000;
      84743: inst = 32'hca00004;
      84744: inst = 32'h38632800;
      84745: inst = 32'h38842800;
      84746: inst = 32'h10a00001;
      84747: inst = 32'hca04b0f;
      84748: inst = 32'h13e00001;
      84749: inst = 32'hfe0d96a;
      84750: inst = 32'h5be00000;
      84751: inst = 32'h8c50000;
      84752: inst = 32'h24612800;
      84753: inst = 32'h10a00000;
      84754: inst = 32'hca00004;
      84755: inst = 32'h24822800;
      84756: inst = 32'h10a00000;
      84757: inst = 32'hca00004;
      84758: inst = 32'h38632800;
      84759: inst = 32'h38842800;
      84760: inst = 32'h10a00001;
      84761: inst = 32'hca04b1d;
      84762: inst = 32'h13e00001;
      84763: inst = 32'hfe0d96a;
      84764: inst = 32'h5be00000;
      84765: inst = 32'h8c50000;
      84766: inst = 32'h24612800;
      84767: inst = 32'h10a00000;
      84768: inst = 32'hca00004;
      84769: inst = 32'h24822800;
      84770: inst = 32'h10a00000;
      84771: inst = 32'hca00004;
      84772: inst = 32'h38632800;
      84773: inst = 32'h38842800;
      84774: inst = 32'h10a00001;
      84775: inst = 32'hca04b2b;
      84776: inst = 32'h13e00001;
      84777: inst = 32'hfe0d96a;
      84778: inst = 32'h5be00000;
      84779: inst = 32'h8c50000;
      84780: inst = 32'h24612800;
      84781: inst = 32'h10a00000;
      84782: inst = 32'hca00004;
      84783: inst = 32'h24822800;
      84784: inst = 32'h10a00000;
      84785: inst = 32'hca00004;
      84786: inst = 32'h38632800;
      84787: inst = 32'h38842800;
      84788: inst = 32'h10a00001;
      84789: inst = 32'hca04b39;
      84790: inst = 32'h13e00001;
      84791: inst = 32'hfe0d96a;
      84792: inst = 32'h5be00000;
      84793: inst = 32'h8c50000;
      84794: inst = 32'h24612800;
      84795: inst = 32'h10a00000;
      84796: inst = 32'hca00004;
      84797: inst = 32'h24822800;
      84798: inst = 32'h10a00000;
      84799: inst = 32'hca00004;
      84800: inst = 32'h38632800;
      84801: inst = 32'h38842800;
      84802: inst = 32'h10a00001;
      84803: inst = 32'hca04b47;
      84804: inst = 32'h13e00001;
      84805: inst = 32'hfe0d96a;
      84806: inst = 32'h5be00000;
      84807: inst = 32'h8c50000;
      84808: inst = 32'h24612800;
      84809: inst = 32'h10a00000;
      84810: inst = 32'hca00004;
      84811: inst = 32'h24822800;
      84812: inst = 32'h10a00000;
      84813: inst = 32'hca00004;
      84814: inst = 32'h38632800;
      84815: inst = 32'h38842800;
      84816: inst = 32'h10a00001;
      84817: inst = 32'hca04b55;
      84818: inst = 32'h13e00001;
      84819: inst = 32'hfe0d96a;
      84820: inst = 32'h5be00000;
      84821: inst = 32'h8c50000;
      84822: inst = 32'h24612800;
      84823: inst = 32'h10a00000;
      84824: inst = 32'hca00004;
      84825: inst = 32'h24822800;
      84826: inst = 32'h10a00000;
      84827: inst = 32'hca00004;
      84828: inst = 32'h38632800;
      84829: inst = 32'h38842800;
      84830: inst = 32'h10a00001;
      84831: inst = 32'hca04b63;
      84832: inst = 32'h13e00001;
      84833: inst = 32'hfe0d96a;
      84834: inst = 32'h5be00000;
      84835: inst = 32'h8c50000;
      84836: inst = 32'h24612800;
      84837: inst = 32'h10a00000;
      84838: inst = 32'hca00004;
      84839: inst = 32'h24822800;
      84840: inst = 32'h10a00000;
      84841: inst = 32'hca00004;
      84842: inst = 32'h38632800;
      84843: inst = 32'h38842800;
      84844: inst = 32'h10a00001;
      84845: inst = 32'hca04b71;
      84846: inst = 32'h13e00001;
      84847: inst = 32'hfe0d96a;
      84848: inst = 32'h5be00000;
      84849: inst = 32'h8c50000;
      84850: inst = 32'h24612800;
      84851: inst = 32'h10a00000;
      84852: inst = 32'hca00004;
      84853: inst = 32'h24822800;
      84854: inst = 32'h10a00000;
      84855: inst = 32'hca00004;
      84856: inst = 32'h38632800;
      84857: inst = 32'h38842800;
      84858: inst = 32'h10a00001;
      84859: inst = 32'hca04b7f;
      84860: inst = 32'h13e00001;
      84861: inst = 32'hfe0d96a;
      84862: inst = 32'h5be00000;
      84863: inst = 32'h8c50000;
      84864: inst = 32'h24612800;
      84865: inst = 32'h10a00000;
      84866: inst = 32'hca00004;
      84867: inst = 32'h24822800;
      84868: inst = 32'h10a00000;
      84869: inst = 32'hca00004;
      84870: inst = 32'h38632800;
      84871: inst = 32'h38842800;
      84872: inst = 32'h10a00001;
      84873: inst = 32'hca04b8d;
      84874: inst = 32'h13e00001;
      84875: inst = 32'hfe0d96a;
      84876: inst = 32'h5be00000;
      84877: inst = 32'h8c50000;
      84878: inst = 32'h24612800;
      84879: inst = 32'h10a00000;
      84880: inst = 32'hca00004;
      84881: inst = 32'h24822800;
      84882: inst = 32'h10a00000;
      84883: inst = 32'hca00004;
      84884: inst = 32'h38632800;
      84885: inst = 32'h38842800;
      84886: inst = 32'h10a00001;
      84887: inst = 32'hca04b9b;
      84888: inst = 32'h13e00001;
      84889: inst = 32'hfe0d96a;
      84890: inst = 32'h5be00000;
      84891: inst = 32'h8c50000;
      84892: inst = 32'h24612800;
      84893: inst = 32'h10a00000;
      84894: inst = 32'hca00004;
      84895: inst = 32'h24822800;
      84896: inst = 32'h10a00000;
      84897: inst = 32'hca00004;
      84898: inst = 32'h38632800;
      84899: inst = 32'h38842800;
      84900: inst = 32'h10a00001;
      84901: inst = 32'hca04ba9;
      84902: inst = 32'h13e00001;
      84903: inst = 32'hfe0d96a;
      84904: inst = 32'h5be00000;
      84905: inst = 32'h8c50000;
      84906: inst = 32'h24612800;
      84907: inst = 32'h10a00000;
      84908: inst = 32'hca00005;
      84909: inst = 32'h24822800;
      84910: inst = 32'h10a00000;
      84911: inst = 32'hca00004;
      84912: inst = 32'h38632800;
      84913: inst = 32'h38842800;
      84914: inst = 32'h10a00001;
      84915: inst = 32'hca04bb7;
      84916: inst = 32'h13e00001;
      84917: inst = 32'hfe0d96a;
      84918: inst = 32'h5be00000;
      84919: inst = 32'h8c50000;
      84920: inst = 32'h24612800;
      84921: inst = 32'h10a00000;
      84922: inst = 32'hca00005;
      84923: inst = 32'h24822800;
      84924: inst = 32'h10a00000;
      84925: inst = 32'hca00004;
      84926: inst = 32'h38632800;
      84927: inst = 32'h38842800;
      84928: inst = 32'h10a00001;
      84929: inst = 32'hca04bc5;
      84930: inst = 32'h13e00001;
      84931: inst = 32'hfe0d96a;
      84932: inst = 32'h5be00000;
      84933: inst = 32'h8c50000;
      84934: inst = 32'h24612800;
      84935: inst = 32'h10a00000;
      84936: inst = 32'hca00005;
      84937: inst = 32'h24822800;
      84938: inst = 32'h10a00000;
      84939: inst = 32'hca00004;
      84940: inst = 32'h38632800;
      84941: inst = 32'h38842800;
      84942: inst = 32'h10a00001;
      84943: inst = 32'hca04bd3;
      84944: inst = 32'h13e00001;
      84945: inst = 32'hfe0d96a;
      84946: inst = 32'h5be00000;
      84947: inst = 32'h8c50000;
      84948: inst = 32'h24612800;
      84949: inst = 32'h10a00000;
      84950: inst = 32'hca00005;
      84951: inst = 32'h24822800;
      84952: inst = 32'h10a00000;
      84953: inst = 32'hca00004;
      84954: inst = 32'h38632800;
      84955: inst = 32'h38842800;
      84956: inst = 32'h10a00001;
      84957: inst = 32'hca04be1;
      84958: inst = 32'h13e00001;
      84959: inst = 32'hfe0d96a;
      84960: inst = 32'h5be00000;
      84961: inst = 32'h8c50000;
      84962: inst = 32'h24612800;
      84963: inst = 32'h10a00000;
      84964: inst = 32'hca00005;
      84965: inst = 32'h24822800;
      84966: inst = 32'h10a00000;
      84967: inst = 32'hca00004;
      84968: inst = 32'h38632800;
      84969: inst = 32'h38842800;
      84970: inst = 32'h10a00001;
      84971: inst = 32'hca04bef;
      84972: inst = 32'h13e00001;
      84973: inst = 32'hfe0d96a;
      84974: inst = 32'h5be00000;
      84975: inst = 32'h8c50000;
      84976: inst = 32'h24612800;
      84977: inst = 32'h10a00000;
      84978: inst = 32'hca00005;
      84979: inst = 32'h24822800;
      84980: inst = 32'h10a00000;
      84981: inst = 32'hca00004;
      84982: inst = 32'h38632800;
      84983: inst = 32'h38842800;
      84984: inst = 32'h10a00001;
      84985: inst = 32'hca04bfd;
      84986: inst = 32'h13e00001;
      84987: inst = 32'hfe0d96a;
      84988: inst = 32'h5be00000;
      84989: inst = 32'h8c50000;
      84990: inst = 32'h24612800;
      84991: inst = 32'h10a00000;
      84992: inst = 32'hca00005;
      84993: inst = 32'h24822800;
      84994: inst = 32'h10a00000;
      84995: inst = 32'hca00004;
      84996: inst = 32'h38632800;
      84997: inst = 32'h38842800;
      84998: inst = 32'h10a00001;
      84999: inst = 32'hca04c0b;
      85000: inst = 32'h13e00001;
      85001: inst = 32'hfe0d96a;
      85002: inst = 32'h5be00000;
      85003: inst = 32'h8c50000;
      85004: inst = 32'h24612800;
      85005: inst = 32'h10a00000;
      85006: inst = 32'hca00005;
      85007: inst = 32'h24822800;
      85008: inst = 32'h10a00000;
      85009: inst = 32'hca00004;
      85010: inst = 32'h38632800;
      85011: inst = 32'h38842800;
      85012: inst = 32'h10a00001;
      85013: inst = 32'hca04c19;
      85014: inst = 32'h13e00001;
      85015: inst = 32'hfe0d96a;
      85016: inst = 32'h5be00000;
      85017: inst = 32'h8c50000;
      85018: inst = 32'h24612800;
      85019: inst = 32'h10a00000;
      85020: inst = 32'hca00005;
      85021: inst = 32'h24822800;
      85022: inst = 32'h10a00000;
      85023: inst = 32'hca00004;
      85024: inst = 32'h38632800;
      85025: inst = 32'h38842800;
      85026: inst = 32'h10a00001;
      85027: inst = 32'hca04c27;
      85028: inst = 32'h13e00001;
      85029: inst = 32'hfe0d96a;
      85030: inst = 32'h5be00000;
      85031: inst = 32'h8c50000;
      85032: inst = 32'h24612800;
      85033: inst = 32'h10a00000;
      85034: inst = 32'hca00005;
      85035: inst = 32'h24822800;
      85036: inst = 32'h10a00000;
      85037: inst = 32'hca00004;
      85038: inst = 32'h38632800;
      85039: inst = 32'h38842800;
      85040: inst = 32'h10a00001;
      85041: inst = 32'hca04c35;
      85042: inst = 32'h13e00001;
      85043: inst = 32'hfe0d96a;
      85044: inst = 32'h5be00000;
      85045: inst = 32'h8c50000;
      85046: inst = 32'h24612800;
      85047: inst = 32'h10a00000;
      85048: inst = 32'hca00005;
      85049: inst = 32'h24822800;
      85050: inst = 32'h10a00000;
      85051: inst = 32'hca00004;
      85052: inst = 32'h38632800;
      85053: inst = 32'h38842800;
      85054: inst = 32'h10a00001;
      85055: inst = 32'hca04c43;
      85056: inst = 32'h13e00001;
      85057: inst = 32'hfe0d96a;
      85058: inst = 32'h5be00000;
      85059: inst = 32'h8c50000;
      85060: inst = 32'h24612800;
      85061: inst = 32'h10a00000;
      85062: inst = 32'hca00005;
      85063: inst = 32'h24822800;
      85064: inst = 32'h10a00000;
      85065: inst = 32'hca00004;
      85066: inst = 32'h38632800;
      85067: inst = 32'h38842800;
      85068: inst = 32'h10a00001;
      85069: inst = 32'hca04c51;
      85070: inst = 32'h13e00001;
      85071: inst = 32'hfe0d96a;
      85072: inst = 32'h5be00000;
      85073: inst = 32'h8c50000;
      85074: inst = 32'h24612800;
      85075: inst = 32'h10a00000;
      85076: inst = 32'hca00005;
      85077: inst = 32'h24822800;
      85078: inst = 32'h10a00000;
      85079: inst = 32'hca00004;
      85080: inst = 32'h38632800;
      85081: inst = 32'h38842800;
      85082: inst = 32'h10a00001;
      85083: inst = 32'hca04c5f;
      85084: inst = 32'h13e00001;
      85085: inst = 32'hfe0d96a;
      85086: inst = 32'h5be00000;
      85087: inst = 32'h8c50000;
      85088: inst = 32'h24612800;
      85089: inst = 32'h10a00000;
      85090: inst = 32'hca00005;
      85091: inst = 32'h24822800;
      85092: inst = 32'h10a00000;
      85093: inst = 32'hca00004;
      85094: inst = 32'h38632800;
      85095: inst = 32'h38842800;
      85096: inst = 32'h10a00001;
      85097: inst = 32'hca04c6d;
      85098: inst = 32'h13e00001;
      85099: inst = 32'hfe0d96a;
      85100: inst = 32'h5be00000;
      85101: inst = 32'h8c50000;
      85102: inst = 32'h24612800;
      85103: inst = 32'h10a00000;
      85104: inst = 32'hca00005;
      85105: inst = 32'h24822800;
      85106: inst = 32'h10a00000;
      85107: inst = 32'hca00004;
      85108: inst = 32'h38632800;
      85109: inst = 32'h38842800;
      85110: inst = 32'h10a00001;
      85111: inst = 32'hca04c7b;
      85112: inst = 32'h13e00001;
      85113: inst = 32'hfe0d96a;
      85114: inst = 32'h5be00000;
      85115: inst = 32'h8c50000;
      85116: inst = 32'h24612800;
      85117: inst = 32'h10a00000;
      85118: inst = 32'hca00005;
      85119: inst = 32'h24822800;
      85120: inst = 32'h10a00000;
      85121: inst = 32'hca00004;
      85122: inst = 32'h38632800;
      85123: inst = 32'h38842800;
      85124: inst = 32'h10a00001;
      85125: inst = 32'hca04c89;
      85126: inst = 32'h13e00001;
      85127: inst = 32'hfe0d96a;
      85128: inst = 32'h5be00000;
      85129: inst = 32'h8c50000;
      85130: inst = 32'h24612800;
      85131: inst = 32'h10a00000;
      85132: inst = 32'hca00005;
      85133: inst = 32'h24822800;
      85134: inst = 32'h10a00000;
      85135: inst = 32'hca00004;
      85136: inst = 32'h38632800;
      85137: inst = 32'h38842800;
      85138: inst = 32'h10a00001;
      85139: inst = 32'hca04c97;
      85140: inst = 32'h13e00001;
      85141: inst = 32'hfe0d96a;
      85142: inst = 32'h5be00000;
      85143: inst = 32'h8c50000;
      85144: inst = 32'h24612800;
      85145: inst = 32'h10a00000;
      85146: inst = 32'hca00005;
      85147: inst = 32'h24822800;
      85148: inst = 32'h10a00000;
      85149: inst = 32'hca00004;
      85150: inst = 32'h38632800;
      85151: inst = 32'h38842800;
      85152: inst = 32'h10a00001;
      85153: inst = 32'hca04ca5;
      85154: inst = 32'h13e00001;
      85155: inst = 32'hfe0d96a;
      85156: inst = 32'h5be00000;
      85157: inst = 32'h8c50000;
      85158: inst = 32'h24612800;
      85159: inst = 32'h10a00000;
      85160: inst = 32'hca00005;
      85161: inst = 32'h24822800;
      85162: inst = 32'h10a00000;
      85163: inst = 32'hca00004;
      85164: inst = 32'h38632800;
      85165: inst = 32'h38842800;
      85166: inst = 32'h10a00001;
      85167: inst = 32'hca04cb3;
      85168: inst = 32'h13e00001;
      85169: inst = 32'hfe0d96a;
      85170: inst = 32'h5be00000;
      85171: inst = 32'h8c50000;
      85172: inst = 32'h24612800;
      85173: inst = 32'h10a00000;
      85174: inst = 32'hca00005;
      85175: inst = 32'h24822800;
      85176: inst = 32'h10a00000;
      85177: inst = 32'hca00004;
      85178: inst = 32'h38632800;
      85179: inst = 32'h38842800;
      85180: inst = 32'h10a00001;
      85181: inst = 32'hca04cc1;
      85182: inst = 32'h13e00001;
      85183: inst = 32'hfe0d96a;
      85184: inst = 32'h5be00000;
      85185: inst = 32'h8c50000;
      85186: inst = 32'h24612800;
      85187: inst = 32'h10a00000;
      85188: inst = 32'hca00005;
      85189: inst = 32'h24822800;
      85190: inst = 32'h10a00000;
      85191: inst = 32'hca00004;
      85192: inst = 32'h38632800;
      85193: inst = 32'h38842800;
      85194: inst = 32'h10a00001;
      85195: inst = 32'hca04ccf;
      85196: inst = 32'h13e00001;
      85197: inst = 32'hfe0d96a;
      85198: inst = 32'h5be00000;
      85199: inst = 32'h8c50000;
      85200: inst = 32'h24612800;
      85201: inst = 32'h10a00000;
      85202: inst = 32'hca00005;
      85203: inst = 32'h24822800;
      85204: inst = 32'h10a00000;
      85205: inst = 32'hca00004;
      85206: inst = 32'h38632800;
      85207: inst = 32'h38842800;
      85208: inst = 32'h10a00001;
      85209: inst = 32'hca04cdd;
      85210: inst = 32'h13e00001;
      85211: inst = 32'hfe0d96a;
      85212: inst = 32'h5be00000;
      85213: inst = 32'h8c50000;
      85214: inst = 32'h24612800;
      85215: inst = 32'h10a00000;
      85216: inst = 32'hca00005;
      85217: inst = 32'h24822800;
      85218: inst = 32'h10a00000;
      85219: inst = 32'hca00004;
      85220: inst = 32'h38632800;
      85221: inst = 32'h38842800;
      85222: inst = 32'h10a00001;
      85223: inst = 32'hca04ceb;
      85224: inst = 32'h13e00001;
      85225: inst = 32'hfe0d96a;
      85226: inst = 32'h5be00000;
      85227: inst = 32'h8c50000;
      85228: inst = 32'h24612800;
      85229: inst = 32'h10a00000;
      85230: inst = 32'hca00005;
      85231: inst = 32'h24822800;
      85232: inst = 32'h10a00000;
      85233: inst = 32'hca00004;
      85234: inst = 32'h38632800;
      85235: inst = 32'h38842800;
      85236: inst = 32'h10a00001;
      85237: inst = 32'hca04cf9;
      85238: inst = 32'h13e00001;
      85239: inst = 32'hfe0d96a;
      85240: inst = 32'h5be00000;
      85241: inst = 32'h8c50000;
      85242: inst = 32'h24612800;
      85243: inst = 32'h10a00000;
      85244: inst = 32'hca00005;
      85245: inst = 32'h24822800;
      85246: inst = 32'h10a00000;
      85247: inst = 32'hca00004;
      85248: inst = 32'h38632800;
      85249: inst = 32'h38842800;
      85250: inst = 32'h10a00001;
      85251: inst = 32'hca04d07;
      85252: inst = 32'h13e00001;
      85253: inst = 32'hfe0d96a;
      85254: inst = 32'h5be00000;
      85255: inst = 32'h8c50000;
      85256: inst = 32'h24612800;
      85257: inst = 32'h10a00000;
      85258: inst = 32'hca00005;
      85259: inst = 32'h24822800;
      85260: inst = 32'h10a00000;
      85261: inst = 32'hca00004;
      85262: inst = 32'h38632800;
      85263: inst = 32'h38842800;
      85264: inst = 32'h10a00001;
      85265: inst = 32'hca04d15;
      85266: inst = 32'h13e00001;
      85267: inst = 32'hfe0d96a;
      85268: inst = 32'h5be00000;
      85269: inst = 32'h8c50000;
      85270: inst = 32'h24612800;
      85271: inst = 32'h10a00000;
      85272: inst = 32'hca00005;
      85273: inst = 32'h24822800;
      85274: inst = 32'h10a00000;
      85275: inst = 32'hca00004;
      85276: inst = 32'h38632800;
      85277: inst = 32'h38842800;
      85278: inst = 32'h10a00001;
      85279: inst = 32'hca04d23;
      85280: inst = 32'h13e00001;
      85281: inst = 32'hfe0d96a;
      85282: inst = 32'h5be00000;
      85283: inst = 32'h8c50000;
      85284: inst = 32'h24612800;
      85285: inst = 32'h10a00000;
      85286: inst = 32'hca00005;
      85287: inst = 32'h24822800;
      85288: inst = 32'h10a00000;
      85289: inst = 32'hca00004;
      85290: inst = 32'h38632800;
      85291: inst = 32'h38842800;
      85292: inst = 32'h10a00001;
      85293: inst = 32'hca04d31;
      85294: inst = 32'h13e00001;
      85295: inst = 32'hfe0d96a;
      85296: inst = 32'h5be00000;
      85297: inst = 32'h8c50000;
      85298: inst = 32'h24612800;
      85299: inst = 32'h10a00000;
      85300: inst = 32'hca00005;
      85301: inst = 32'h24822800;
      85302: inst = 32'h10a00000;
      85303: inst = 32'hca00004;
      85304: inst = 32'h38632800;
      85305: inst = 32'h38842800;
      85306: inst = 32'h10a00001;
      85307: inst = 32'hca04d3f;
      85308: inst = 32'h13e00001;
      85309: inst = 32'hfe0d96a;
      85310: inst = 32'h5be00000;
      85311: inst = 32'h8c50000;
      85312: inst = 32'h24612800;
      85313: inst = 32'h10a00000;
      85314: inst = 32'hca00005;
      85315: inst = 32'h24822800;
      85316: inst = 32'h10a00000;
      85317: inst = 32'hca00004;
      85318: inst = 32'h38632800;
      85319: inst = 32'h38842800;
      85320: inst = 32'h10a00001;
      85321: inst = 32'hca04d4d;
      85322: inst = 32'h13e00001;
      85323: inst = 32'hfe0d96a;
      85324: inst = 32'h5be00000;
      85325: inst = 32'h8c50000;
      85326: inst = 32'h24612800;
      85327: inst = 32'h10a00000;
      85328: inst = 32'hca00005;
      85329: inst = 32'h24822800;
      85330: inst = 32'h10a00000;
      85331: inst = 32'hca00004;
      85332: inst = 32'h38632800;
      85333: inst = 32'h38842800;
      85334: inst = 32'h10a00001;
      85335: inst = 32'hca04d5b;
      85336: inst = 32'h13e00001;
      85337: inst = 32'hfe0d96a;
      85338: inst = 32'h5be00000;
      85339: inst = 32'h8c50000;
      85340: inst = 32'h24612800;
      85341: inst = 32'h10a00000;
      85342: inst = 32'hca00005;
      85343: inst = 32'h24822800;
      85344: inst = 32'h10a00000;
      85345: inst = 32'hca00004;
      85346: inst = 32'h38632800;
      85347: inst = 32'h38842800;
      85348: inst = 32'h10a00001;
      85349: inst = 32'hca04d69;
      85350: inst = 32'h13e00001;
      85351: inst = 32'hfe0d96a;
      85352: inst = 32'h5be00000;
      85353: inst = 32'h8c50000;
      85354: inst = 32'h24612800;
      85355: inst = 32'h10a00000;
      85356: inst = 32'hca00005;
      85357: inst = 32'h24822800;
      85358: inst = 32'h10a00000;
      85359: inst = 32'hca00004;
      85360: inst = 32'h38632800;
      85361: inst = 32'h38842800;
      85362: inst = 32'h10a00001;
      85363: inst = 32'hca04d77;
      85364: inst = 32'h13e00001;
      85365: inst = 32'hfe0d96a;
      85366: inst = 32'h5be00000;
      85367: inst = 32'h8c50000;
      85368: inst = 32'h24612800;
      85369: inst = 32'h10a00000;
      85370: inst = 32'hca00005;
      85371: inst = 32'h24822800;
      85372: inst = 32'h10a00000;
      85373: inst = 32'hca00004;
      85374: inst = 32'h38632800;
      85375: inst = 32'h38842800;
      85376: inst = 32'h10a00001;
      85377: inst = 32'hca04d85;
      85378: inst = 32'h13e00001;
      85379: inst = 32'hfe0d96a;
      85380: inst = 32'h5be00000;
      85381: inst = 32'h8c50000;
      85382: inst = 32'h24612800;
      85383: inst = 32'h10a00000;
      85384: inst = 32'hca00005;
      85385: inst = 32'h24822800;
      85386: inst = 32'h10a00000;
      85387: inst = 32'hca00004;
      85388: inst = 32'h38632800;
      85389: inst = 32'h38842800;
      85390: inst = 32'h10a00001;
      85391: inst = 32'hca04d93;
      85392: inst = 32'h13e00001;
      85393: inst = 32'hfe0d96a;
      85394: inst = 32'h5be00000;
      85395: inst = 32'h8c50000;
      85396: inst = 32'h24612800;
      85397: inst = 32'h10a00000;
      85398: inst = 32'hca00005;
      85399: inst = 32'h24822800;
      85400: inst = 32'h10a00000;
      85401: inst = 32'hca00004;
      85402: inst = 32'h38632800;
      85403: inst = 32'h38842800;
      85404: inst = 32'h10a00001;
      85405: inst = 32'hca04da1;
      85406: inst = 32'h13e00001;
      85407: inst = 32'hfe0d96a;
      85408: inst = 32'h5be00000;
      85409: inst = 32'h8c50000;
      85410: inst = 32'h24612800;
      85411: inst = 32'h10a00000;
      85412: inst = 32'hca00005;
      85413: inst = 32'h24822800;
      85414: inst = 32'h10a00000;
      85415: inst = 32'hca00004;
      85416: inst = 32'h38632800;
      85417: inst = 32'h38842800;
      85418: inst = 32'h10a00001;
      85419: inst = 32'hca04daf;
      85420: inst = 32'h13e00001;
      85421: inst = 32'hfe0d96a;
      85422: inst = 32'h5be00000;
      85423: inst = 32'h8c50000;
      85424: inst = 32'h24612800;
      85425: inst = 32'h10a00000;
      85426: inst = 32'hca00005;
      85427: inst = 32'h24822800;
      85428: inst = 32'h10a00000;
      85429: inst = 32'hca00004;
      85430: inst = 32'h38632800;
      85431: inst = 32'h38842800;
      85432: inst = 32'h10a00001;
      85433: inst = 32'hca04dbd;
      85434: inst = 32'h13e00001;
      85435: inst = 32'hfe0d96a;
      85436: inst = 32'h5be00000;
      85437: inst = 32'h8c50000;
      85438: inst = 32'h24612800;
      85439: inst = 32'h10a00000;
      85440: inst = 32'hca00005;
      85441: inst = 32'h24822800;
      85442: inst = 32'h10a00000;
      85443: inst = 32'hca00004;
      85444: inst = 32'h38632800;
      85445: inst = 32'h38842800;
      85446: inst = 32'h10a00001;
      85447: inst = 32'hca04dcb;
      85448: inst = 32'h13e00001;
      85449: inst = 32'hfe0d96a;
      85450: inst = 32'h5be00000;
      85451: inst = 32'h8c50000;
      85452: inst = 32'h24612800;
      85453: inst = 32'h10a00000;
      85454: inst = 32'hca00005;
      85455: inst = 32'h24822800;
      85456: inst = 32'h10a00000;
      85457: inst = 32'hca00004;
      85458: inst = 32'h38632800;
      85459: inst = 32'h38842800;
      85460: inst = 32'h10a00001;
      85461: inst = 32'hca04dd9;
      85462: inst = 32'h13e00001;
      85463: inst = 32'hfe0d96a;
      85464: inst = 32'h5be00000;
      85465: inst = 32'h8c50000;
      85466: inst = 32'h24612800;
      85467: inst = 32'h10a00000;
      85468: inst = 32'hca00005;
      85469: inst = 32'h24822800;
      85470: inst = 32'h10a00000;
      85471: inst = 32'hca00004;
      85472: inst = 32'h38632800;
      85473: inst = 32'h38842800;
      85474: inst = 32'h10a00001;
      85475: inst = 32'hca04de7;
      85476: inst = 32'h13e00001;
      85477: inst = 32'hfe0d96a;
      85478: inst = 32'h5be00000;
      85479: inst = 32'h8c50000;
      85480: inst = 32'h24612800;
      85481: inst = 32'h10a00000;
      85482: inst = 32'hca00005;
      85483: inst = 32'h24822800;
      85484: inst = 32'h10a00000;
      85485: inst = 32'hca00004;
      85486: inst = 32'h38632800;
      85487: inst = 32'h38842800;
      85488: inst = 32'h10a00001;
      85489: inst = 32'hca04df5;
      85490: inst = 32'h13e00001;
      85491: inst = 32'hfe0d96a;
      85492: inst = 32'h5be00000;
      85493: inst = 32'h8c50000;
      85494: inst = 32'h24612800;
      85495: inst = 32'h10a00000;
      85496: inst = 32'hca00005;
      85497: inst = 32'h24822800;
      85498: inst = 32'h10a00000;
      85499: inst = 32'hca00004;
      85500: inst = 32'h38632800;
      85501: inst = 32'h38842800;
      85502: inst = 32'h10a00001;
      85503: inst = 32'hca04e03;
      85504: inst = 32'h13e00001;
      85505: inst = 32'hfe0d96a;
      85506: inst = 32'h5be00000;
      85507: inst = 32'h8c50000;
      85508: inst = 32'h24612800;
      85509: inst = 32'h10a00000;
      85510: inst = 32'hca00005;
      85511: inst = 32'h24822800;
      85512: inst = 32'h10a00000;
      85513: inst = 32'hca00004;
      85514: inst = 32'h38632800;
      85515: inst = 32'h38842800;
      85516: inst = 32'h10a00001;
      85517: inst = 32'hca04e11;
      85518: inst = 32'h13e00001;
      85519: inst = 32'hfe0d96a;
      85520: inst = 32'h5be00000;
      85521: inst = 32'h8c50000;
      85522: inst = 32'h24612800;
      85523: inst = 32'h10a00000;
      85524: inst = 32'hca00005;
      85525: inst = 32'h24822800;
      85526: inst = 32'h10a00000;
      85527: inst = 32'hca00004;
      85528: inst = 32'h38632800;
      85529: inst = 32'h38842800;
      85530: inst = 32'h10a00001;
      85531: inst = 32'hca04e1f;
      85532: inst = 32'h13e00001;
      85533: inst = 32'hfe0d96a;
      85534: inst = 32'h5be00000;
      85535: inst = 32'h8c50000;
      85536: inst = 32'h24612800;
      85537: inst = 32'h10a00000;
      85538: inst = 32'hca00005;
      85539: inst = 32'h24822800;
      85540: inst = 32'h10a00000;
      85541: inst = 32'hca00004;
      85542: inst = 32'h38632800;
      85543: inst = 32'h38842800;
      85544: inst = 32'h10a00001;
      85545: inst = 32'hca04e2d;
      85546: inst = 32'h13e00001;
      85547: inst = 32'hfe0d96a;
      85548: inst = 32'h5be00000;
      85549: inst = 32'h8c50000;
      85550: inst = 32'h24612800;
      85551: inst = 32'h10a00000;
      85552: inst = 32'hca00005;
      85553: inst = 32'h24822800;
      85554: inst = 32'h10a00000;
      85555: inst = 32'hca00004;
      85556: inst = 32'h38632800;
      85557: inst = 32'h38842800;
      85558: inst = 32'h10a00001;
      85559: inst = 32'hca04e3b;
      85560: inst = 32'h13e00001;
      85561: inst = 32'hfe0d96a;
      85562: inst = 32'h5be00000;
      85563: inst = 32'h8c50000;
      85564: inst = 32'h24612800;
      85565: inst = 32'h10a00000;
      85566: inst = 32'hca00005;
      85567: inst = 32'h24822800;
      85568: inst = 32'h10a00000;
      85569: inst = 32'hca00004;
      85570: inst = 32'h38632800;
      85571: inst = 32'h38842800;
      85572: inst = 32'h10a00001;
      85573: inst = 32'hca04e49;
      85574: inst = 32'h13e00001;
      85575: inst = 32'hfe0d96a;
      85576: inst = 32'h5be00000;
      85577: inst = 32'h8c50000;
      85578: inst = 32'h24612800;
      85579: inst = 32'h10a00000;
      85580: inst = 32'hca00005;
      85581: inst = 32'h24822800;
      85582: inst = 32'h10a00000;
      85583: inst = 32'hca00004;
      85584: inst = 32'h38632800;
      85585: inst = 32'h38842800;
      85586: inst = 32'h10a00001;
      85587: inst = 32'hca04e57;
      85588: inst = 32'h13e00001;
      85589: inst = 32'hfe0d96a;
      85590: inst = 32'h5be00000;
      85591: inst = 32'h8c50000;
      85592: inst = 32'h24612800;
      85593: inst = 32'h10a00000;
      85594: inst = 32'hca00005;
      85595: inst = 32'h24822800;
      85596: inst = 32'h10a00000;
      85597: inst = 32'hca00004;
      85598: inst = 32'h38632800;
      85599: inst = 32'h38842800;
      85600: inst = 32'h10a00001;
      85601: inst = 32'hca04e65;
      85602: inst = 32'h13e00001;
      85603: inst = 32'hfe0d96a;
      85604: inst = 32'h5be00000;
      85605: inst = 32'h8c50000;
      85606: inst = 32'h24612800;
      85607: inst = 32'h10a00000;
      85608: inst = 32'hca00005;
      85609: inst = 32'h24822800;
      85610: inst = 32'h10a00000;
      85611: inst = 32'hca00004;
      85612: inst = 32'h38632800;
      85613: inst = 32'h38842800;
      85614: inst = 32'h10a00001;
      85615: inst = 32'hca04e73;
      85616: inst = 32'h13e00001;
      85617: inst = 32'hfe0d96a;
      85618: inst = 32'h5be00000;
      85619: inst = 32'h8c50000;
      85620: inst = 32'h24612800;
      85621: inst = 32'h10a00000;
      85622: inst = 32'hca00005;
      85623: inst = 32'h24822800;
      85624: inst = 32'h10a00000;
      85625: inst = 32'hca00004;
      85626: inst = 32'h38632800;
      85627: inst = 32'h38842800;
      85628: inst = 32'h10a00001;
      85629: inst = 32'hca04e81;
      85630: inst = 32'h13e00001;
      85631: inst = 32'hfe0d96a;
      85632: inst = 32'h5be00000;
      85633: inst = 32'h8c50000;
      85634: inst = 32'h24612800;
      85635: inst = 32'h10a00000;
      85636: inst = 32'hca00005;
      85637: inst = 32'h24822800;
      85638: inst = 32'h10a00000;
      85639: inst = 32'hca00004;
      85640: inst = 32'h38632800;
      85641: inst = 32'h38842800;
      85642: inst = 32'h10a00001;
      85643: inst = 32'hca04e8f;
      85644: inst = 32'h13e00001;
      85645: inst = 32'hfe0d96a;
      85646: inst = 32'h5be00000;
      85647: inst = 32'h8c50000;
      85648: inst = 32'h24612800;
      85649: inst = 32'h10a00000;
      85650: inst = 32'hca00005;
      85651: inst = 32'h24822800;
      85652: inst = 32'h10a00000;
      85653: inst = 32'hca00004;
      85654: inst = 32'h38632800;
      85655: inst = 32'h38842800;
      85656: inst = 32'h10a00001;
      85657: inst = 32'hca04e9d;
      85658: inst = 32'h13e00001;
      85659: inst = 32'hfe0d96a;
      85660: inst = 32'h5be00000;
      85661: inst = 32'h8c50000;
      85662: inst = 32'h24612800;
      85663: inst = 32'h10a00000;
      85664: inst = 32'hca00005;
      85665: inst = 32'h24822800;
      85666: inst = 32'h10a00000;
      85667: inst = 32'hca00004;
      85668: inst = 32'h38632800;
      85669: inst = 32'h38842800;
      85670: inst = 32'h10a00001;
      85671: inst = 32'hca04eab;
      85672: inst = 32'h13e00001;
      85673: inst = 32'hfe0d96a;
      85674: inst = 32'h5be00000;
      85675: inst = 32'h8c50000;
      85676: inst = 32'h24612800;
      85677: inst = 32'h10a00000;
      85678: inst = 32'hca00005;
      85679: inst = 32'h24822800;
      85680: inst = 32'h10a00000;
      85681: inst = 32'hca00004;
      85682: inst = 32'h38632800;
      85683: inst = 32'h38842800;
      85684: inst = 32'h10a00001;
      85685: inst = 32'hca04eb9;
      85686: inst = 32'h13e00001;
      85687: inst = 32'hfe0d96a;
      85688: inst = 32'h5be00000;
      85689: inst = 32'h8c50000;
      85690: inst = 32'h24612800;
      85691: inst = 32'h10a00000;
      85692: inst = 32'hca00005;
      85693: inst = 32'h24822800;
      85694: inst = 32'h10a00000;
      85695: inst = 32'hca00004;
      85696: inst = 32'h38632800;
      85697: inst = 32'h38842800;
      85698: inst = 32'h10a00001;
      85699: inst = 32'hca04ec7;
      85700: inst = 32'h13e00001;
      85701: inst = 32'hfe0d96a;
      85702: inst = 32'h5be00000;
      85703: inst = 32'h8c50000;
      85704: inst = 32'h24612800;
      85705: inst = 32'h10a00000;
      85706: inst = 32'hca00005;
      85707: inst = 32'h24822800;
      85708: inst = 32'h10a00000;
      85709: inst = 32'hca00004;
      85710: inst = 32'h38632800;
      85711: inst = 32'h38842800;
      85712: inst = 32'h10a00001;
      85713: inst = 32'hca04ed5;
      85714: inst = 32'h13e00001;
      85715: inst = 32'hfe0d96a;
      85716: inst = 32'h5be00000;
      85717: inst = 32'h8c50000;
      85718: inst = 32'h24612800;
      85719: inst = 32'h10a00000;
      85720: inst = 32'hca00005;
      85721: inst = 32'h24822800;
      85722: inst = 32'h10a00000;
      85723: inst = 32'hca00004;
      85724: inst = 32'h38632800;
      85725: inst = 32'h38842800;
      85726: inst = 32'h10a00001;
      85727: inst = 32'hca04ee3;
      85728: inst = 32'h13e00001;
      85729: inst = 32'hfe0d96a;
      85730: inst = 32'h5be00000;
      85731: inst = 32'h8c50000;
      85732: inst = 32'h24612800;
      85733: inst = 32'h10a00000;
      85734: inst = 32'hca00005;
      85735: inst = 32'h24822800;
      85736: inst = 32'h10a00000;
      85737: inst = 32'hca00004;
      85738: inst = 32'h38632800;
      85739: inst = 32'h38842800;
      85740: inst = 32'h10a00001;
      85741: inst = 32'hca04ef1;
      85742: inst = 32'h13e00001;
      85743: inst = 32'hfe0d96a;
      85744: inst = 32'h5be00000;
      85745: inst = 32'h8c50000;
      85746: inst = 32'h24612800;
      85747: inst = 32'h10a00000;
      85748: inst = 32'hca00005;
      85749: inst = 32'h24822800;
      85750: inst = 32'h10a00000;
      85751: inst = 32'hca00004;
      85752: inst = 32'h38632800;
      85753: inst = 32'h38842800;
      85754: inst = 32'h10a00001;
      85755: inst = 32'hca04eff;
      85756: inst = 32'h13e00001;
      85757: inst = 32'hfe0d96a;
      85758: inst = 32'h5be00000;
      85759: inst = 32'h8c50000;
      85760: inst = 32'h24612800;
      85761: inst = 32'h10a00000;
      85762: inst = 32'hca00005;
      85763: inst = 32'h24822800;
      85764: inst = 32'h10a00000;
      85765: inst = 32'hca00004;
      85766: inst = 32'h38632800;
      85767: inst = 32'h38842800;
      85768: inst = 32'h10a00001;
      85769: inst = 32'hca04f0d;
      85770: inst = 32'h13e00001;
      85771: inst = 32'hfe0d96a;
      85772: inst = 32'h5be00000;
      85773: inst = 32'h8c50000;
      85774: inst = 32'h24612800;
      85775: inst = 32'h10a00000;
      85776: inst = 32'hca00005;
      85777: inst = 32'h24822800;
      85778: inst = 32'h10a00000;
      85779: inst = 32'hca00004;
      85780: inst = 32'h38632800;
      85781: inst = 32'h38842800;
      85782: inst = 32'h10a00001;
      85783: inst = 32'hca04f1b;
      85784: inst = 32'h13e00001;
      85785: inst = 32'hfe0d96a;
      85786: inst = 32'h5be00000;
      85787: inst = 32'h8c50000;
      85788: inst = 32'h24612800;
      85789: inst = 32'h10a00000;
      85790: inst = 32'hca00005;
      85791: inst = 32'h24822800;
      85792: inst = 32'h10a00000;
      85793: inst = 32'hca00004;
      85794: inst = 32'h38632800;
      85795: inst = 32'h38842800;
      85796: inst = 32'h10a00001;
      85797: inst = 32'hca04f29;
      85798: inst = 32'h13e00001;
      85799: inst = 32'hfe0d96a;
      85800: inst = 32'h5be00000;
      85801: inst = 32'h8c50000;
      85802: inst = 32'h24612800;
      85803: inst = 32'h10a00000;
      85804: inst = 32'hca00005;
      85805: inst = 32'h24822800;
      85806: inst = 32'h10a00000;
      85807: inst = 32'hca00004;
      85808: inst = 32'h38632800;
      85809: inst = 32'h38842800;
      85810: inst = 32'h10a00001;
      85811: inst = 32'hca04f37;
      85812: inst = 32'h13e00001;
      85813: inst = 32'hfe0d96a;
      85814: inst = 32'h5be00000;
      85815: inst = 32'h8c50000;
      85816: inst = 32'h24612800;
      85817: inst = 32'h10a00000;
      85818: inst = 32'hca00005;
      85819: inst = 32'h24822800;
      85820: inst = 32'h10a00000;
      85821: inst = 32'hca00004;
      85822: inst = 32'h38632800;
      85823: inst = 32'h38842800;
      85824: inst = 32'h10a00001;
      85825: inst = 32'hca04f45;
      85826: inst = 32'h13e00001;
      85827: inst = 32'hfe0d96a;
      85828: inst = 32'h5be00000;
      85829: inst = 32'h8c50000;
      85830: inst = 32'h24612800;
      85831: inst = 32'h10a00000;
      85832: inst = 32'hca00005;
      85833: inst = 32'h24822800;
      85834: inst = 32'h10a00000;
      85835: inst = 32'hca00004;
      85836: inst = 32'h38632800;
      85837: inst = 32'h38842800;
      85838: inst = 32'h10a00001;
      85839: inst = 32'hca04f53;
      85840: inst = 32'h13e00001;
      85841: inst = 32'hfe0d96a;
      85842: inst = 32'h5be00000;
      85843: inst = 32'h8c50000;
      85844: inst = 32'h24612800;
      85845: inst = 32'h10a00000;
      85846: inst = 32'hca00005;
      85847: inst = 32'h24822800;
      85848: inst = 32'h10a00000;
      85849: inst = 32'hca00004;
      85850: inst = 32'h38632800;
      85851: inst = 32'h38842800;
      85852: inst = 32'h10a00001;
      85853: inst = 32'hca04f61;
      85854: inst = 32'h13e00001;
      85855: inst = 32'hfe0d96a;
      85856: inst = 32'h5be00000;
      85857: inst = 32'h8c50000;
      85858: inst = 32'h24612800;
      85859: inst = 32'h10a00000;
      85860: inst = 32'hca00005;
      85861: inst = 32'h24822800;
      85862: inst = 32'h10a00000;
      85863: inst = 32'hca00004;
      85864: inst = 32'h38632800;
      85865: inst = 32'h38842800;
      85866: inst = 32'h10a00001;
      85867: inst = 32'hca04f6f;
      85868: inst = 32'h13e00001;
      85869: inst = 32'hfe0d96a;
      85870: inst = 32'h5be00000;
      85871: inst = 32'h8c50000;
      85872: inst = 32'h24612800;
      85873: inst = 32'h10a00000;
      85874: inst = 32'hca00005;
      85875: inst = 32'h24822800;
      85876: inst = 32'h10a00000;
      85877: inst = 32'hca00004;
      85878: inst = 32'h38632800;
      85879: inst = 32'h38842800;
      85880: inst = 32'h10a00001;
      85881: inst = 32'hca04f7d;
      85882: inst = 32'h13e00001;
      85883: inst = 32'hfe0d96a;
      85884: inst = 32'h5be00000;
      85885: inst = 32'h8c50000;
      85886: inst = 32'h24612800;
      85887: inst = 32'h10a00000;
      85888: inst = 32'hca00005;
      85889: inst = 32'h24822800;
      85890: inst = 32'h10a00000;
      85891: inst = 32'hca00004;
      85892: inst = 32'h38632800;
      85893: inst = 32'h38842800;
      85894: inst = 32'h10a00001;
      85895: inst = 32'hca04f8b;
      85896: inst = 32'h13e00001;
      85897: inst = 32'hfe0d96a;
      85898: inst = 32'h5be00000;
      85899: inst = 32'h8c50000;
      85900: inst = 32'h24612800;
      85901: inst = 32'h10a00000;
      85902: inst = 32'hca00005;
      85903: inst = 32'h24822800;
      85904: inst = 32'h10a00000;
      85905: inst = 32'hca00004;
      85906: inst = 32'h38632800;
      85907: inst = 32'h38842800;
      85908: inst = 32'h10a00001;
      85909: inst = 32'hca04f99;
      85910: inst = 32'h13e00001;
      85911: inst = 32'hfe0d96a;
      85912: inst = 32'h5be00000;
      85913: inst = 32'h8c50000;
      85914: inst = 32'h24612800;
      85915: inst = 32'h10a00000;
      85916: inst = 32'hca00005;
      85917: inst = 32'h24822800;
      85918: inst = 32'h10a00000;
      85919: inst = 32'hca00004;
      85920: inst = 32'h38632800;
      85921: inst = 32'h38842800;
      85922: inst = 32'h10a00001;
      85923: inst = 32'hca04fa7;
      85924: inst = 32'h13e00001;
      85925: inst = 32'hfe0d96a;
      85926: inst = 32'h5be00000;
      85927: inst = 32'h8c50000;
      85928: inst = 32'h24612800;
      85929: inst = 32'h10a00000;
      85930: inst = 32'hca00005;
      85931: inst = 32'h24822800;
      85932: inst = 32'h10a00000;
      85933: inst = 32'hca00004;
      85934: inst = 32'h38632800;
      85935: inst = 32'h38842800;
      85936: inst = 32'h10a00001;
      85937: inst = 32'hca04fb5;
      85938: inst = 32'h13e00001;
      85939: inst = 32'hfe0d96a;
      85940: inst = 32'h5be00000;
      85941: inst = 32'h8c50000;
      85942: inst = 32'h24612800;
      85943: inst = 32'h10a00000;
      85944: inst = 32'hca00005;
      85945: inst = 32'h24822800;
      85946: inst = 32'h10a00000;
      85947: inst = 32'hca00004;
      85948: inst = 32'h38632800;
      85949: inst = 32'h38842800;
      85950: inst = 32'h10a00001;
      85951: inst = 32'hca04fc3;
      85952: inst = 32'h13e00001;
      85953: inst = 32'hfe0d96a;
      85954: inst = 32'h5be00000;
      85955: inst = 32'h8c50000;
      85956: inst = 32'h24612800;
      85957: inst = 32'h10a00000;
      85958: inst = 32'hca00005;
      85959: inst = 32'h24822800;
      85960: inst = 32'h10a00000;
      85961: inst = 32'hca00004;
      85962: inst = 32'h38632800;
      85963: inst = 32'h38842800;
      85964: inst = 32'h10a00001;
      85965: inst = 32'hca04fd1;
      85966: inst = 32'h13e00001;
      85967: inst = 32'hfe0d96a;
      85968: inst = 32'h5be00000;
      85969: inst = 32'h8c50000;
      85970: inst = 32'h24612800;
      85971: inst = 32'h10a00000;
      85972: inst = 32'hca00005;
      85973: inst = 32'h24822800;
      85974: inst = 32'h10a00000;
      85975: inst = 32'hca00004;
      85976: inst = 32'h38632800;
      85977: inst = 32'h38842800;
      85978: inst = 32'h10a00001;
      85979: inst = 32'hca04fdf;
      85980: inst = 32'h13e00001;
      85981: inst = 32'hfe0d96a;
      85982: inst = 32'h5be00000;
      85983: inst = 32'h8c50000;
      85984: inst = 32'h24612800;
      85985: inst = 32'h10a00000;
      85986: inst = 32'hca00005;
      85987: inst = 32'h24822800;
      85988: inst = 32'h10a00000;
      85989: inst = 32'hca00004;
      85990: inst = 32'h38632800;
      85991: inst = 32'h38842800;
      85992: inst = 32'h10a00001;
      85993: inst = 32'hca04fed;
      85994: inst = 32'h13e00001;
      85995: inst = 32'hfe0d96a;
      85996: inst = 32'h5be00000;
      85997: inst = 32'h8c50000;
      85998: inst = 32'h24612800;
      85999: inst = 32'h10a00000;
      86000: inst = 32'hca00005;
      86001: inst = 32'h24822800;
      86002: inst = 32'h10a00000;
      86003: inst = 32'hca00004;
      86004: inst = 32'h38632800;
      86005: inst = 32'h38842800;
      86006: inst = 32'h10a00001;
      86007: inst = 32'hca04ffb;
      86008: inst = 32'h13e00001;
      86009: inst = 32'hfe0d96a;
      86010: inst = 32'h5be00000;
      86011: inst = 32'h8c50000;
      86012: inst = 32'h24612800;
      86013: inst = 32'h10a00000;
      86014: inst = 32'hca00005;
      86015: inst = 32'h24822800;
      86016: inst = 32'h10a00000;
      86017: inst = 32'hca00004;
      86018: inst = 32'h38632800;
      86019: inst = 32'h38842800;
      86020: inst = 32'h10a00001;
      86021: inst = 32'hca05009;
      86022: inst = 32'h13e00001;
      86023: inst = 32'hfe0d96a;
      86024: inst = 32'h5be00000;
      86025: inst = 32'h8c50000;
      86026: inst = 32'h24612800;
      86027: inst = 32'h10a00000;
      86028: inst = 32'hca00005;
      86029: inst = 32'h24822800;
      86030: inst = 32'h10a00000;
      86031: inst = 32'hca00004;
      86032: inst = 32'h38632800;
      86033: inst = 32'h38842800;
      86034: inst = 32'h10a00001;
      86035: inst = 32'hca05017;
      86036: inst = 32'h13e00001;
      86037: inst = 32'hfe0d96a;
      86038: inst = 32'h5be00000;
      86039: inst = 32'h8c50000;
      86040: inst = 32'h24612800;
      86041: inst = 32'h10a00000;
      86042: inst = 32'hca00005;
      86043: inst = 32'h24822800;
      86044: inst = 32'h10a00000;
      86045: inst = 32'hca00004;
      86046: inst = 32'h38632800;
      86047: inst = 32'h38842800;
      86048: inst = 32'h10a00001;
      86049: inst = 32'hca05025;
      86050: inst = 32'h13e00001;
      86051: inst = 32'hfe0d96a;
      86052: inst = 32'h5be00000;
      86053: inst = 32'h8c50000;
      86054: inst = 32'h24612800;
      86055: inst = 32'h10a00000;
      86056: inst = 32'hca00005;
      86057: inst = 32'h24822800;
      86058: inst = 32'h10a00000;
      86059: inst = 32'hca00004;
      86060: inst = 32'h38632800;
      86061: inst = 32'h38842800;
      86062: inst = 32'h10a00001;
      86063: inst = 32'hca05033;
      86064: inst = 32'h13e00001;
      86065: inst = 32'hfe0d96a;
      86066: inst = 32'h5be00000;
      86067: inst = 32'h8c50000;
      86068: inst = 32'h24612800;
      86069: inst = 32'h10a00000;
      86070: inst = 32'hca00005;
      86071: inst = 32'h24822800;
      86072: inst = 32'h10a00000;
      86073: inst = 32'hca00004;
      86074: inst = 32'h38632800;
      86075: inst = 32'h38842800;
      86076: inst = 32'h10a00001;
      86077: inst = 32'hca05041;
      86078: inst = 32'h13e00001;
      86079: inst = 32'hfe0d96a;
      86080: inst = 32'h5be00000;
      86081: inst = 32'h8c50000;
      86082: inst = 32'h24612800;
      86083: inst = 32'h10a00000;
      86084: inst = 32'hca00005;
      86085: inst = 32'h24822800;
      86086: inst = 32'h10a00000;
      86087: inst = 32'hca00004;
      86088: inst = 32'h38632800;
      86089: inst = 32'h38842800;
      86090: inst = 32'h10a00001;
      86091: inst = 32'hca0504f;
      86092: inst = 32'h13e00001;
      86093: inst = 32'hfe0d96a;
      86094: inst = 32'h5be00000;
      86095: inst = 32'h8c50000;
      86096: inst = 32'h24612800;
      86097: inst = 32'h10a00000;
      86098: inst = 32'hca00005;
      86099: inst = 32'h24822800;
      86100: inst = 32'h10a00000;
      86101: inst = 32'hca00004;
      86102: inst = 32'h38632800;
      86103: inst = 32'h38842800;
      86104: inst = 32'h10a00001;
      86105: inst = 32'hca0505d;
      86106: inst = 32'h13e00001;
      86107: inst = 32'hfe0d96a;
      86108: inst = 32'h5be00000;
      86109: inst = 32'h8c50000;
      86110: inst = 32'h24612800;
      86111: inst = 32'h10a00000;
      86112: inst = 32'hca00005;
      86113: inst = 32'h24822800;
      86114: inst = 32'h10a00000;
      86115: inst = 32'hca00004;
      86116: inst = 32'h38632800;
      86117: inst = 32'h38842800;
      86118: inst = 32'h10a00001;
      86119: inst = 32'hca0506b;
      86120: inst = 32'h13e00001;
      86121: inst = 32'hfe0d96a;
      86122: inst = 32'h5be00000;
      86123: inst = 32'h8c50000;
      86124: inst = 32'h24612800;
      86125: inst = 32'h10a00000;
      86126: inst = 32'hca00005;
      86127: inst = 32'h24822800;
      86128: inst = 32'h10a00000;
      86129: inst = 32'hca00004;
      86130: inst = 32'h38632800;
      86131: inst = 32'h38842800;
      86132: inst = 32'h10a00001;
      86133: inst = 32'hca05079;
      86134: inst = 32'h13e00001;
      86135: inst = 32'hfe0d96a;
      86136: inst = 32'h5be00000;
      86137: inst = 32'h8c50000;
      86138: inst = 32'h24612800;
      86139: inst = 32'h10a00000;
      86140: inst = 32'hca00005;
      86141: inst = 32'h24822800;
      86142: inst = 32'h10a00000;
      86143: inst = 32'hca00004;
      86144: inst = 32'h38632800;
      86145: inst = 32'h38842800;
      86146: inst = 32'h10a00001;
      86147: inst = 32'hca05087;
      86148: inst = 32'h13e00001;
      86149: inst = 32'hfe0d96a;
      86150: inst = 32'h5be00000;
      86151: inst = 32'h8c50000;
      86152: inst = 32'h24612800;
      86153: inst = 32'h10a00000;
      86154: inst = 32'hca00005;
      86155: inst = 32'h24822800;
      86156: inst = 32'h10a00000;
      86157: inst = 32'hca00004;
      86158: inst = 32'h38632800;
      86159: inst = 32'h38842800;
      86160: inst = 32'h10a00001;
      86161: inst = 32'hca05095;
      86162: inst = 32'h13e00001;
      86163: inst = 32'hfe0d96a;
      86164: inst = 32'h5be00000;
      86165: inst = 32'h8c50000;
      86166: inst = 32'h24612800;
      86167: inst = 32'h10a00000;
      86168: inst = 32'hca00005;
      86169: inst = 32'h24822800;
      86170: inst = 32'h10a00000;
      86171: inst = 32'hca00004;
      86172: inst = 32'h38632800;
      86173: inst = 32'h38842800;
      86174: inst = 32'h10a00001;
      86175: inst = 32'hca050a3;
      86176: inst = 32'h13e00001;
      86177: inst = 32'hfe0d96a;
      86178: inst = 32'h5be00000;
      86179: inst = 32'h8c50000;
      86180: inst = 32'h24612800;
      86181: inst = 32'h10a00000;
      86182: inst = 32'hca00005;
      86183: inst = 32'h24822800;
      86184: inst = 32'h10a00000;
      86185: inst = 32'hca00004;
      86186: inst = 32'h38632800;
      86187: inst = 32'h38842800;
      86188: inst = 32'h10a00001;
      86189: inst = 32'hca050b1;
      86190: inst = 32'h13e00001;
      86191: inst = 32'hfe0d96a;
      86192: inst = 32'h5be00000;
      86193: inst = 32'h8c50000;
      86194: inst = 32'h24612800;
      86195: inst = 32'h10a00000;
      86196: inst = 32'hca00005;
      86197: inst = 32'h24822800;
      86198: inst = 32'h10a00000;
      86199: inst = 32'hca00004;
      86200: inst = 32'h38632800;
      86201: inst = 32'h38842800;
      86202: inst = 32'h10a00001;
      86203: inst = 32'hca050bf;
      86204: inst = 32'h13e00001;
      86205: inst = 32'hfe0d96a;
      86206: inst = 32'h5be00000;
      86207: inst = 32'h8c50000;
      86208: inst = 32'h24612800;
      86209: inst = 32'h10a00000;
      86210: inst = 32'hca00005;
      86211: inst = 32'h24822800;
      86212: inst = 32'h10a00000;
      86213: inst = 32'hca00004;
      86214: inst = 32'h38632800;
      86215: inst = 32'h38842800;
      86216: inst = 32'h10a00001;
      86217: inst = 32'hca050cd;
      86218: inst = 32'h13e00001;
      86219: inst = 32'hfe0d96a;
      86220: inst = 32'h5be00000;
      86221: inst = 32'h8c50000;
      86222: inst = 32'h24612800;
      86223: inst = 32'h10a00000;
      86224: inst = 32'hca00005;
      86225: inst = 32'h24822800;
      86226: inst = 32'h10a00000;
      86227: inst = 32'hca00004;
      86228: inst = 32'h38632800;
      86229: inst = 32'h38842800;
      86230: inst = 32'h10a00001;
      86231: inst = 32'hca050db;
      86232: inst = 32'h13e00001;
      86233: inst = 32'hfe0d96a;
      86234: inst = 32'h5be00000;
      86235: inst = 32'h8c50000;
      86236: inst = 32'h24612800;
      86237: inst = 32'h10a00000;
      86238: inst = 32'hca00005;
      86239: inst = 32'h24822800;
      86240: inst = 32'h10a00000;
      86241: inst = 32'hca00004;
      86242: inst = 32'h38632800;
      86243: inst = 32'h38842800;
      86244: inst = 32'h10a00001;
      86245: inst = 32'hca050e9;
      86246: inst = 32'h13e00001;
      86247: inst = 32'hfe0d96a;
      86248: inst = 32'h5be00000;
      86249: inst = 32'h8c50000;
      86250: inst = 32'h24612800;
      86251: inst = 32'h10a00000;
      86252: inst = 32'hca00006;
      86253: inst = 32'h24822800;
      86254: inst = 32'h10a00000;
      86255: inst = 32'hca00004;
      86256: inst = 32'h38632800;
      86257: inst = 32'h38842800;
      86258: inst = 32'h10a00001;
      86259: inst = 32'hca050f7;
      86260: inst = 32'h13e00001;
      86261: inst = 32'hfe0d96a;
      86262: inst = 32'h5be00000;
      86263: inst = 32'h8c50000;
      86264: inst = 32'h24612800;
      86265: inst = 32'h10a00000;
      86266: inst = 32'hca00006;
      86267: inst = 32'h24822800;
      86268: inst = 32'h10a00000;
      86269: inst = 32'hca00004;
      86270: inst = 32'h38632800;
      86271: inst = 32'h38842800;
      86272: inst = 32'h10a00001;
      86273: inst = 32'hca05105;
      86274: inst = 32'h13e00001;
      86275: inst = 32'hfe0d96a;
      86276: inst = 32'h5be00000;
      86277: inst = 32'h8c50000;
      86278: inst = 32'h24612800;
      86279: inst = 32'h10a00000;
      86280: inst = 32'hca00006;
      86281: inst = 32'h24822800;
      86282: inst = 32'h10a00000;
      86283: inst = 32'hca00004;
      86284: inst = 32'h38632800;
      86285: inst = 32'h38842800;
      86286: inst = 32'h10a00001;
      86287: inst = 32'hca05113;
      86288: inst = 32'h13e00001;
      86289: inst = 32'hfe0d96a;
      86290: inst = 32'h5be00000;
      86291: inst = 32'h8c50000;
      86292: inst = 32'h24612800;
      86293: inst = 32'h10a00000;
      86294: inst = 32'hca00006;
      86295: inst = 32'h24822800;
      86296: inst = 32'h10a00000;
      86297: inst = 32'hca00004;
      86298: inst = 32'h38632800;
      86299: inst = 32'h38842800;
      86300: inst = 32'h10a00001;
      86301: inst = 32'hca05121;
      86302: inst = 32'h13e00001;
      86303: inst = 32'hfe0d96a;
      86304: inst = 32'h5be00000;
      86305: inst = 32'h8c50000;
      86306: inst = 32'h24612800;
      86307: inst = 32'h10a00000;
      86308: inst = 32'hca00006;
      86309: inst = 32'h24822800;
      86310: inst = 32'h10a00000;
      86311: inst = 32'hca00004;
      86312: inst = 32'h38632800;
      86313: inst = 32'h38842800;
      86314: inst = 32'h10a00001;
      86315: inst = 32'hca0512f;
      86316: inst = 32'h13e00001;
      86317: inst = 32'hfe0d96a;
      86318: inst = 32'h5be00000;
      86319: inst = 32'h8c50000;
      86320: inst = 32'h24612800;
      86321: inst = 32'h10a00000;
      86322: inst = 32'hca00006;
      86323: inst = 32'h24822800;
      86324: inst = 32'h10a00000;
      86325: inst = 32'hca00004;
      86326: inst = 32'h38632800;
      86327: inst = 32'h38842800;
      86328: inst = 32'h10a00001;
      86329: inst = 32'hca0513d;
      86330: inst = 32'h13e00001;
      86331: inst = 32'hfe0d96a;
      86332: inst = 32'h5be00000;
      86333: inst = 32'h8c50000;
      86334: inst = 32'h24612800;
      86335: inst = 32'h10a00000;
      86336: inst = 32'hca00006;
      86337: inst = 32'h24822800;
      86338: inst = 32'h10a00000;
      86339: inst = 32'hca00004;
      86340: inst = 32'h38632800;
      86341: inst = 32'h38842800;
      86342: inst = 32'h10a00001;
      86343: inst = 32'hca0514b;
      86344: inst = 32'h13e00001;
      86345: inst = 32'hfe0d96a;
      86346: inst = 32'h5be00000;
      86347: inst = 32'h8c50000;
      86348: inst = 32'h24612800;
      86349: inst = 32'h10a00000;
      86350: inst = 32'hca00006;
      86351: inst = 32'h24822800;
      86352: inst = 32'h10a00000;
      86353: inst = 32'hca00004;
      86354: inst = 32'h38632800;
      86355: inst = 32'h38842800;
      86356: inst = 32'h10a00001;
      86357: inst = 32'hca05159;
      86358: inst = 32'h13e00001;
      86359: inst = 32'hfe0d96a;
      86360: inst = 32'h5be00000;
      86361: inst = 32'h8c50000;
      86362: inst = 32'h24612800;
      86363: inst = 32'h10a00000;
      86364: inst = 32'hca00006;
      86365: inst = 32'h24822800;
      86366: inst = 32'h10a00000;
      86367: inst = 32'hca00004;
      86368: inst = 32'h38632800;
      86369: inst = 32'h38842800;
      86370: inst = 32'h10a00001;
      86371: inst = 32'hca05167;
      86372: inst = 32'h13e00001;
      86373: inst = 32'hfe0d96a;
      86374: inst = 32'h5be00000;
      86375: inst = 32'h8c50000;
      86376: inst = 32'h24612800;
      86377: inst = 32'h10a00000;
      86378: inst = 32'hca00006;
      86379: inst = 32'h24822800;
      86380: inst = 32'h10a00000;
      86381: inst = 32'hca00004;
      86382: inst = 32'h38632800;
      86383: inst = 32'h38842800;
      86384: inst = 32'h10a00001;
      86385: inst = 32'hca05175;
      86386: inst = 32'h13e00001;
      86387: inst = 32'hfe0d96a;
      86388: inst = 32'h5be00000;
      86389: inst = 32'h8c50000;
      86390: inst = 32'h24612800;
      86391: inst = 32'h10a00000;
      86392: inst = 32'hca00006;
      86393: inst = 32'h24822800;
      86394: inst = 32'h10a00000;
      86395: inst = 32'hca00004;
      86396: inst = 32'h38632800;
      86397: inst = 32'h38842800;
      86398: inst = 32'h10a00001;
      86399: inst = 32'hca05183;
      86400: inst = 32'h13e00001;
      86401: inst = 32'hfe0d96a;
      86402: inst = 32'h5be00000;
      86403: inst = 32'h8c50000;
      86404: inst = 32'h24612800;
      86405: inst = 32'h10a00000;
      86406: inst = 32'hca00006;
      86407: inst = 32'h24822800;
      86408: inst = 32'h10a00000;
      86409: inst = 32'hca00004;
      86410: inst = 32'h38632800;
      86411: inst = 32'h38842800;
      86412: inst = 32'h10a00001;
      86413: inst = 32'hca05191;
      86414: inst = 32'h13e00001;
      86415: inst = 32'hfe0d96a;
      86416: inst = 32'h5be00000;
      86417: inst = 32'h8c50000;
      86418: inst = 32'h24612800;
      86419: inst = 32'h10a00000;
      86420: inst = 32'hca00006;
      86421: inst = 32'h24822800;
      86422: inst = 32'h10a00000;
      86423: inst = 32'hca00004;
      86424: inst = 32'h38632800;
      86425: inst = 32'h38842800;
      86426: inst = 32'h10a00001;
      86427: inst = 32'hca0519f;
      86428: inst = 32'h13e00001;
      86429: inst = 32'hfe0d96a;
      86430: inst = 32'h5be00000;
      86431: inst = 32'h8c50000;
      86432: inst = 32'h24612800;
      86433: inst = 32'h10a00000;
      86434: inst = 32'hca00006;
      86435: inst = 32'h24822800;
      86436: inst = 32'h10a00000;
      86437: inst = 32'hca00004;
      86438: inst = 32'h38632800;
      86439: inst = 32'h38842800;
      86440: inst = 32'h10a00001;
      86441: inst = 32'hca051ad;
      86442: inst = 32'h13e00001;
      86443: inst = 32'hfe0d96a;
      86444: inst = 32'h5be00000;
      86445: inst = 32'h8c50000;
      86446: inst = 32'h24612800;
      86447: inst = 32'h10a00000;
      86448: inst = 32'hca00006;
      86449: inst = 32'h24822800;
      86450: inst = 32'h10a00000;
      86451: inst = 32'hca00004;
      86452: inst = 32'h38632800;
      86453: inst = 32'h38842800;
      86454: inst = 32'h10a00001;
      86455: inst = 32'hca051bb;
      86456: inst = 32'h13e00001;
      86457: inst = 32'hfe0d96a;
      86458: inst = 32'h5be00000;
      86459: inst = 32'h8c50000;
      86460: inst = 32'h24612800;
      86461: inst = 32'h10a00000;
      86462: inst = 32'hca00006;
      86463: inst = 32'h24822800;
      86464: inst = 32'h10a00000;
      86465: inst = 32'hca00004;
      86466: inst = 32'h38632800;
      86467: inst = 32'h38842800;
      86468: inst = 32'h10a00001;
      86469: inst = 32'hca051c9;
      86470: inst = 32'h13e00001;
      86471: inst = 32'hfe0d96a;
      86472: inst = 32'h5be00000;
      86473: inst = 32'h8c50000;
      86474: inst = 32'h24612800;
      86475: inst = 32'h10a00000;
      86476: inst = 32'hca00006;
      86477: inst = 32'h24822800;
      86478: inst = 32'h10a00000;
      86479: inst = 32'hca00004;
      86480: inst = 32'h38632800;
      86481: inst = 32'h38842800;
      86482: inst = 32'h10a00001;
      86483: inst = 32'hca051d7;
      86484: inst = 32'h13e00001;
      86485: inst = 32'hfe0d96a;
      86486: inst = 32'h5be00000;
      86487: inst = 32'h8c50000;
      86488: inst = 32'h24612800;
      86489: inst = 32'h10a00000;
      86490: inst = 32'hca00006;
      86491: inst = 32'h24822800;
      86492: inst = 32'h10a00000;
      86493: inst = 32'hca00004;
      86494: inst = 32'h38632800;
      86495: inst = 32'h38842800;
      86496: inst = 32'h10a00001;
      86497: inst = 32'hca051e5;
      86498: inst = 32'h13e00001;
      86499: inst = 32'hfe0d96a;
      86500: inst = 32'h5be00000;
      86501: inst = 32'h8c50000;
      86502: inst = 32'h24612800;
      86503: inst = 32'h10a00000;
      86504: inst = 32'hca00006;
      86505: inst = 32'h24822800;
      86506: inst = 32'h10a00000;
      86507: inst = 32'hca00004;
      86508: inst = 32'h38632800;
      86509: inst = 32'h38842800;
      86510: inst = 32'h10a00001;
      86511: inst = 32'hca051f3;
      86512: inst = 32'h13e00001;
      86513: inst = 32'hfe0d96a;
      86514: inst = 32'h5be00000;
      86515: inst = 32'h8c50000;
      86516: inst = 32'h24612800;
      86517: inst = 32'h10a00000;
      86518: inst = 32'hca00006;
      86519: inst = 32'h24822800;
      86520: inst = 32'h10a00000;
      86521: inst = 32'hca00004;
      86522: inst = 32'h38632800;
      86523: inst = 32'h38842800;
      86524: inst = 32'h10a00001;
      86525: inst = 32'hca05201;
      86526: inst = 32'h13e00001;
      86527: inst = 32'hfe0d96a;
      86528: inst = 32'h5be00000;
      86529: inst = 32'h8c50000;
      86530: inst = 32'h24612800;
      86531: inst = 32'h10a00000;
      86532: inst = 32'hca00006;
      86533: inst = 32'h24822800;
      86534: inst = 32'h10a00000;
      86535: inst = 32'hca00004;
      86536: inst = 32'h38632800;
      86537: inst = 32'h38842800;
      86538: inst = 32'h10a00001;
      86539: inst = 32'hca0520f;
      86540: inst = 32'h13e00001;
      86541: inst = 32'hfe0d96a;
      86542: inst = 32'h5be00000;
      86543: inst = 32'h8c50000;
      86544: inst = 32'h24612800;
      86545: inst = 32'h10a00000;
      86546: inst = 32'hca00006;
      86547: inst = 32'h24822800;
      86548: inst = 32'h10a00000;
      86549: inst = 32'hca00004;
      86550: inst = 32'h38632800;
      86551: inst = 32'h38842800;
      86552: inst = 32'h10a00001;
      86553: inst = 32'hca0521d;
      86554: inst = 32'h13e00001;
      86555: inst = 32'hfe0d96a;
      86556: inst = 32'h5be00000;
      86557: inst = 32'h8c50000;
      86558: inst = 32'h24612800;
      86559: inst = 32'h10a00000;
      86560: inst = 32'hca00006;
      86561: inst = 32'h24822800;
      86562: inst = 32'h10a00000;
      86563: inst = 32'hca00004;
      86564: inst = 32'h38632800;
      86565: inst = 32'h38842800;
      86566: inst = 32'h10a00001;
      86567: inst = 32'hca0522b;
      86568: inst = 32'h13e00001;
      86569: inst = 32'hfe0d96a;
      86570: inst = 32'h5be00000;
      86571: inst = 32'h8c50000;
      86572: inst = 32'h24612800;
      86573: inst = 32'h10a00000;
      86574: inst = 32'hca00006;
      86575: inst = 32'h24822800;
      86576: inst = 32'h10a00000;
      86577: inst = 32'hca00004;
      86578: inst = 32'h38632800;
      86579: inst = 32'h38842800;
      86580: inst = 32'h10a00001;
      86581: inst = 32'hca05239;
      86582: inst = 32'h13e00001;
      86583: inst = 32'hfe0d96a;
      86584: inst = 32'h5be00000;
      86585: inst = 32'h8c50000;
      86586: inst = 32'h24612800;
      86587: inst = 32'h10a00000;
      86588: inst = 32'hca00006;
      86589: inst = 32'h24822800;
      86590: inst = 32'h10a00000;
      86591: inst = 32'hca00004;
      86592: inst = 32'h38632800;
      86593: inst = 32'h38842800;
      86594: inst = 32'h10a00001;
      86595: inst = 32'hca05247;
      86596: inst = 32'h13e00001;
      86597: inst = 32'hfe0d96a;
      86598: inst = 32'h5be00000;
      86599: inst = 32'h8c50000;
      86600: inst = 32'h24612800;
      86601: inst = 32'h10a00000;
      86602: inst = 32'hca00006;
      86603: inst = 32'h24822800;
      86604: inst = 32'h10a00000;
      86605: inst = 32'hca00004;
      86606: inst = 32'h38632800;
      86607: inst = 32'h38842800;
      86608: inst = 32'h10a00001;
      86609: inst = 32'hca05255;
      86610: inst = 32'h13e00001;
      86611: inst = 32'hfe0d96a;
      86612: inst = 32'h5be00000;
      86613: inst = 32'h8c50000;
      86614: inst = 32'h24612800;
      86615: inst = 32'h10a00000;
      86616: inst = 32'hca00006;
      86617: inst = 32'h24822800;
      86618: inst = 32'h10a00000;
      86619: inst = 32'hca00004;
      86620: inst = 32'h38632800;
      86621: inst = 32'h38842800;
      86622: inst = 32'h10a00001;
      86623: inst = 32'hca05263;
      86624: inst = 32'h13e00001;
      86625: inst = 32'hfe0d96a;
      86626: inst = 32'h5be00000;
      86627: inst = 32'h8c50000;
      86628: inst = 32'h24612800;
      86629: inst = 32'h10a00000;
      86630: inst = 32'hca00006;
      86631: inst = 32'h24822800;
      86632: inst = 32'h10a00000;
      86633: inst = 32'hca00004;
      86634: inst = 32'h38632800;
      86635: inst = 32'h38842800;
      86636: inst = 32'h10a00001;
      86637: inst = 32'hca05271;
      86638: inst = 32'h13e00001;
      86639: inst = 32'hfe0d96a;
      86640: inst = 32'h5be00000;
      86641: inst = 32'h8c50000;
      86642: inst = 32'h24612800;
      86643: inst = 32'h10a00000;
      86644: inst = 32'hca00006;
      86645: inst = 32'h24822800;
      86646: inst = 32'h10a00000;
      86647: inst = 32'hca00004;
      86648: inst = 32'h38632800;
      86649: inst = 32'h38842800;
      86650: inst = 32'h10a00001;
      86651: inst = 32'hca0527f;
      86652: inst = 32'h13e00001;
      86653: inst = 32'hfe0d96a;
      86654: inst = 32'h5be00000;
      86655: inst = 32'h8c50000;
      86656: inst = 32'h24612800;
      86657: inst = 32'h10a00000;
      86658: inst = 32'hca00006;
      86659: inst = 32'h24822800;
      86660: inst = 32'h10a00000;
      86661: inst = 32'hca00004;
      86662: inst = 32'h38632800;
      86663: inst = 32'h38842800;
      86664: inst = 32'h10a00001;
      86665: inst = 32'hca0528d;
      86666: inst = 32'h13e00001;
      86667: inst = 32'hfe0d96a;
      86668: inst = 32'h5be00000;
      86669: inst = 32'h8c50000;
      86670: inst = 32'h24612800;
      86671: inst = 32'h10a00000;
      86672: inst = 32'hca00006;
      86673: inst = 32'h24822800;
      86674: inst = 32'h10a00000;
      86675: inst = 32'hca00004;
      86676: inst = 32'h38632800;
      86677: inst = 32'h38842800;
      86678: inst = 32'h10a00001;
      86679: inst = 32'hca0529b;
      86680: inst = 32'h13e00001;
      86681: inst = 32'hfe0d96a;
      86682: inst = 32'h5be00000;
      86683: inst = 32'h8c50000;
      86684: inst = 32'h24612800;
      86685: inst = 32'h10a00000;
      86686: inst = 32'hca00006;
      86687: inst = 32'h24822800;
      86688: inst = 32'h10a00000;
      86689: inst = 32'hca00004;
      86690: inst = 32'h38632800;
      86691: inst = 32'h38842800;
      86692: inst = 32'h10a00001;
      86693: inst = 32'hca052a9;
      86694: inst = 32'h13e00001;
      86695: inst = 32'hfe0d96a;
      86696: inst = 32'h5be00000;
      86697: inst = 32'h8c50000;
      86698: inst = 32'h24612800;
      86699: inst = 32'h10a00000;
      86700: inst = 32'hca00006;
      86701: inst = 32'h24822800;
      86702: inst = 32'h10a00000;
      86703: inst = 32'hca00004;
      86704: inst = 32'h38632800;
      86705: inst = 32'h38842800;
      86706: inst = 32'h10a00001;
      86707: inst = 32'hca052b7;
      86708: inst = 32'h13e00001;
      86709: inst = 32'hfe0d96a;
      86710: inst = 32'h5be00000;
      86711: inst = 32'h8c50000;
      86712: inst = 32'h24612800;
      86713: inst = 32'h10a00000;
      86714: inst = 32'hca00006;
      86715: inst = 32'h24822800;
      86716: inst = 32'h10a00000;
      86717: inst = 32'hca00004;
      86718: inst = 32'h38632800;
      86719: inst = 32'h38842800;
      86720: inst = 32'h10a00001;
      86721: inst = 32'hca052c5;
      86722: inst = 32'h13e00001;
      86723: inst = 32'hfe0d96a;
      86724: inst = 32'h5be00000;
      86725: inst = 32'h8c50000;
      86726: inst = 32'h24612800;
      86727: inst = 32'h10a00000;
      86728: inst = 32'hca00006;
      86729: inst = 32'h24822800;
      86730: inst = 32'h10a00000;
      86731: inst = 32'hca00004;
      86732: inst = 32'h38632800;
      86733: inst = 32'h38842800;
      86734: inst = 32'h10a00001;
      86735: inst = 32'hca052d3;
      86736: inst = 32'h13e00001;
      86737: inst = 32'hfe0d96a;
      86738: inst = 32'h5be00000;
      86739: inst = 32'h8c50000;
      86740: inst = 32'h24612800;
      86741: inst = 32'h10a00000;
      86742: inst = 32'hca00006;
      86743: inst = 32'h24822800;
      86744: inst = 32'h10a00000;
      86745: inst = 32'hca00004;
      86746: inst = 32'h38632800;
      86747: inst = 32'h38842800;
      86748: inst = 32'h10a00001;
      86749: inst = 32'hca052e1;
      86750: inst = 32'h13e00001;
      86751: inst = 32'hfe0d96a;
      86752: inst = 32'h5be00000;
      86753: inst = 32'h8c50000;
      86754: inst = 32'h24612800;
      86755: inst = 32'h10a00000;
      86756: inst = 32'hca00006;
      86757: inst = 32'h24822800;
      86758: inst = 32'h10a00000;
      86759: inst = 32'hca00004;
      86760: inst = 32'h38632800;
      86761: inst = 32'h38842800;
      86762: inst = 32'h10a00001;
      86763: inst = 32'hca052ef;
      86764: inst = 32'h13e00001;
      86765: inst = 32'hfe0d96a;
      86766: inst = 32'h5be00000;
      86767: inst = 32'h8c50000;
      86768: inst = 32'h24612800;
      86769: inst = 32'h10a00000;
      86770: inst = 32'hca00006;
      86771: inst = 32'h24822800;
      86772: inst = 32'h10a00000;
      86773: inst = 32'hca00004;
      86774: inst = 32'h38632800;
      86775: inst = 32'h38842800;
      86776: inst = 32'h10a00001;
      86777: inst = 32'hca052fd;
      86778: inst = 32'h13e00001;
      86779: inst = 32'hfe0d96a;
      86780: inst = 32'h5be00000;
      86781: inst = 32'h8c50000;
      86782: inst = 32'h24612800;
      86783: inst = 32'h10a00000;
      86784: inst = 32'hca00006;
      86785: inst = 32'h24822800;
      86786: inst = 32'h10a00000;
      86787: inst = 32'hca00004;
      86788: inst = 32'h38632800;
      86789: inst = 32'h38842800;
      86790: inst = 32'h10a00001;
      86791: inst = 32'hca0530b;
      86792: inst = 32'h13e00001;
      86793: inst = 32'hfe0d96a;
      86794: inst = 32'h5be00000;
      86795: inst = 32'h8c50000;
      86796: inst = 32'h24612800;
      86797: inst = 32'h10a00000;
      86798: inst = 32'hca00006;
      86799: inst = 32'h24822800;
      86800: inst = 32'h10a00000;
      86801: inst = 32'hca00004;
      86802: inst = 32'h38632800;
      86803: inst = 32'h38842800;
      86804: inst = 32'h10a00001;
      86805: inst = 32'hca05319;
      86806: inst = 32'h13e00001;
      86807: inst = 32'hfe0d96a;
      86808: inst = 32'h5be00000;
      86809: inst = 32'h8c50000;
      86810: inst = 32'h24612800;
      86811: inst = 32'h10a00000;
      86812: inst = 32'hca00006;
      86813: inst = 32'h24822800;
      86814: inst = 32'h10a00000;
      86815: inst = 32'hca00004;
      86816: inst = 32'h38632800;
      86817: inst = 32'h38842800;
      86818: inst = 32'h10a00001;
      86819: inst = 32'hca05327;
      86820: inst = 32'h13e00001;
      86821: inst = 32'hfe0d96a;
      86822: inst = 32'h5be00000;
      86823: inst = 32'h8c50000;
      86824: inst = 32'h24612800;
      86825: inst = 32'h10a00000;
      86826: inst = 32'hca00006;
      86827: inst = 32'h24822800;
      86828: inst = 32'h10a00000;
      86829: inst = 32'hca00004;
      86830: inst = 32'h38632800;
      86831: inst = 32'h38842800;
      86832: inst = 32'h10a00001;
      86833: inst = 32'hca05335;
      86834: inst = 32'h13e00001;
      86835: inst = 32'hfe0d96a;
      86836: inst = 32'h5be00000;
      86837: inst = 32'h8c50000;
      86838: inst = 32'h24612800;
      86839: inst = 32'h10a00000;
      86840: inst = 32'hca00006;
      86841: inst = 32'h24822800;
      86842: inst = 32'h10a00000;
      86843: inst = 32'hca00004;
      86844: inst = 32'h38632800;
      86845: inst = 32'h38842800;
      86846: inst = 32'h10a00001;
      86847: inst = 32'hca05343;
      86848: inst = 32'h13e00001;
      86849: inst = 32'hfe0d96a;
      86850: inst = 32'h5be00000;
      86851: inst = 32'h8c50000;
      86852: inst = 32'h24612800;
      86853: inst = 32'h10a00000;
      86854: inst = 32'hca00006;
      86855: inst = 32'h24822800;
      86856: inst = 32'h10a00000;
      86857: inst = 32'hca00004;
      86858: inst = 32'h38632800;
      86859: inst = 32'h38842800;
      86860: inst = 32'h10a00001;
      86861: inst = 32'hca05351;
      86862: inst = 32'h13e00001;
      86863: inst = 32'hfe0d96a;
      86864: inst = 32'h5be00000;
      86865: inst = 32'h8c50000;
      86866: inst = 32'h24612800;
      86867: inst = 32'h10a00000;
      86868: inst = 32'hca00006;
      86869: inst = 32'h24822800;
      86870: inst = 32'h10a00000;
      86871: inst = 32'hca00004;
      86872: inst = 32'h38632800;
      86873: inst = 32'h38842800;
      86874: inst = 32'h10a00001;
      86875: inst = 32'hca0535f;
      86876: inst = 32'h13e00001;
      86877: inst = 32'hfe0d96a;
      86878: inst = 32'h5be00000;
      86879: inst = 32'h8c50000;
      86880: inst = 32'h24612800;
      86881: inst = 32'h10a00000;
      86882: inst = 32'hca00006;
      86883: inst = 32'h24822800;
      86884: inst = 32'h10a00000;
      86885: inst = 32'hca00004;
      86886: inst = 32'h38632800;
      86887: inst = 32'h38842800;
      86888: inst = 32'h10a00001;
      86889: inst = 32'hca0536d;
      86890: inst = 32'h13e00001;
      86891: inst = 32'hfe0d96a;
      86892: inst = 32'h5be00000;
      86893: inst = 32'h8c50000;
      86894: inst = 32'h24612800;
      86895: inst = 32'h10a00000;
      86896: inst = 32'hca00006;
      86897: inst = 32'h24822800;
      86898: inst = 32'h10a00000;
      86899: inst = 32'hca00004;
      86900: inst = 32'h38632800;
      86901: inst = 32'h38842800;
      86902: inst = 32'h10a00001;
      86903: inst = 32'hca0537b;
      86904: inst = 32'h13e00001;
      86905: inst = 32'hfe0d96a;
      86906: inst = 32'h5be00000;
      86907: inst = 32'h8c50000;
      86908: inst = 32'h24612800;
      86909: inst = 32'h10a00000;
      86910: inst = 32'hca00006;
      86911: inst = 32'h24822800;
      86912: inst = 32'h10a00000;
      86913: inst = 32'hca00004;
      86914: inst = 32'h38632800;
      86915: inst = 32'h38842800;
      86916: inst = 32'h10a00001;
      86917: inst = 32'hca05389;
      86918: inst = 32'h13e00001;
      86919: inst = 32'hfe0d96a;
      86920: inst = 32'h5be00000;
      86921: inst = 32'h8c50000;
      86922: inst = 32'h24612800;
      86923: inst = 32'h10a00000;
      86924: inst = 32'hca00006;
      86925: inst = 32'h24822800;
      86926: inst = 32'h10a00000;
      86927: inst = 32'hca00004;
      86928: inst = 32'h38632800;
      86929: inst = 32'h38842800;
      86930: inst = 32'h10a00001;
      86931: inst = 32'hca05397;
      86932: inst = 32'h13e00001;
      86933: inst = 32'hfe0d96a;
      86934: inst = 32'h5be00000;
      86935: inst = 32'h8c50000;
      86936: inst = 32'h24612800;
      86937: inst = 32'h10a00000;
      86938: inst = 32'hca00006;
      86939: inst = 32'h24822800;
      86940: inst = 32'h10a00000;
      86941: inst = 32'hca00004;
      86942: inst = 32'h38632800;
      86943: inst = 32'h38842800;
      86944: inst = 32'h10a00001;
      86945: inst = 32'hca053a5;
      86946: inst = 32'h13e00001;
      86947: inst = 32'hfe0d96a;
      86948: inst = 32'h5be00000;
      86949: inst = 32'h8c50000;
      86950: inst = 32'h24612800;
      86951: inst = 32'h10a00000;
      86952: inst = 32'hca00006;
      86953: inst = 32'h24822800;
      86954: inst = 32'h10a00000;
      86955: inst = 32'hca00004;
      86956: inst = 32'h38632800;
      86957: inst = 32'h38842800;
      86958: inst = 32'h10a00001;
      86959: inst = 32'hca053b3;
      86960: inst = 32'h13e00001;
      86961: inst = 32'hfe0d96a;
      86962: inst = 32'h5be00000;
      86963: inst = 32'h8c50000;
      86964: inst = 32'h24612800;
      86965: inst = 32'h10a00000;
      86966: inst = 32'hca00006;
      86967: inst = 32'h24822800;
      86968: inst = 32'h10a00000;
      86969: inst = 32'hca00004;
      86970: inst = 32'h38632800;
      86971: inst = 32'h38842800;
      86972: inst = 32'h10a00001;
      86973: inst = 32'hca053c1;
      86974: inst = 32'h13e00001;
      86975: inst = 32'hfe0d96a;
      86976: inst = 32'h5be00000;
      86977: inst = 32'h8c50000;
      86978: inst = 32'h24612800;
      86979: inst = 32'h10a00000;
      86980: inst = 32'hca00006;
      86981: inst = 32'h24822800;
      86982: inst = 32'h10a00000;
      86983: inst = 32'hca00004;
      86984: inst = 32'h38632800;
      86985: inst = 32'h38842800;
      86986: inst = 32'h10a00001;
      86987: inst = 32'hca053cf;
      86988: inst = 32'h13e00001;
      86989: inst = 32'hfe0d96a;
      86990: inst = 32'h5be00000;
      86991: inst = 32'h8c50000;
      86992: inst = 32'h24612800;
      86993: inst = 32'h10a00000;
      86994: inst = 32'hca00006;
      86995: inst = 32'h24822800;
      86996: inst = 32'h10a00000;
      86997: inst = 32'hca00004;
      86998: inst = 32'h38632800;
      86999: inst = 32'h38842800;
      87000: inst = 32'h10a00001;
      87001: inst = 32'hca053dd;
      87002: inst = 32'h13e00001;
      87003: inst = 32'hfe0d96a;
      87004: inst = 32'h5be00000;
      87005: inst = 32'h8c50000;
      87006: inst = 32'h24612800;
      87007: inst = 32'h10a00000;
      87008: inst = 32'hca00006;
      87009: inst = 32'h24822800;
      87010: inst = 32'h10a00000;
      87011: inst = 32'hca00004;
      87012: inst = 32'h38632800;
      87013: inst = 32'h38842800;
      87014: inst = 32'h10a00001;
      87015: inst = 32'hca053eb;
      87016: inst = 32'h13e00001;
      87017: inst = 32'hfe0d96a;
      87018: inst = 32'h5be00000;
      87019: inst = 32'h8c50000;
      87020: inst = 32'h24612800;
      87021: inst = 32'h10a00000;
      87022: inst = 32'hca00006;
      87023: inst = 32'h24822800;
      87024: inst = 32'h10a00000;
      87025: inst = 32'hca00004;
      87026: inst = 32'h38632800;
      87027: inst = 32'h38842800;
      87028: inst = 32'h10a00001;
      87029: inst = 32'hca053f9;
      87030: inst = 32'h13e00001;
      87031: inst = 32'hfe0d96a;
      87032: inst = 32'h5be00000;
      87033: inst = 32'h8c50000;
      87034: inst = 32'h24612800;
      87035: inst = 32'h10a00000;
      87036: inst = 32'hca00006;
      87037: inst = 32'h24822800;
      87038: inst = 32'h10a00000;
      87039: inst = 32'hca00004;
      87040: inst = 32'h38632800;
      87041: inst = 32'h38842800;
      87042: inst = 32'h10a00001;
      87043: inst = 32'hca05407;
      87044: inst = 32'h13e00001;
      87045: inst = 32'hfe0d96a;
      87046: inst = 32'h5be00000;
      87047: inst = 32'h8c50000;
      87048: inst = 32'h24612800;
      87049: inst = 32'h10a00000;
      87050: inst = 32'hca00006;
      87051: inst = 32'h24822800;
      87052: inst = 32'h10a00000;
      87053: inst = 32'hca00004;
      87054: inst = 32'h38632800;
      87055: inst = 32'h38842800;
      87056: inst = 32'h10a00001;
      87057: inst = 32'hca05415;
      87058: inst = 32'h13e00001;
      87059: inst = 32'hfe0d96a;
      87060: inst = 32'h5be00000;
      87061: inst = 32'h8c50000;
      87062: inst = 32'h24612800;
      87063: inst = 32'h10a00000;
      87064: inst = 32'hca00006;
      87065: inst = 32'h24822800;
      87066: inst = 32'h10a00000;
      87067: inst = 32'hca00004;
      87068: inst = 32'h38632800;
      87069: inst = 32'h38842800;
      87070: inst = 32'h10a00001;
      87071: inst = 32'hca05423;
      87072: inst = 32'h13e00001;
      87073: inst = 32'hfe0d96a;
      87074: inst = 32'h5be00000;
      87075: inst = 32'h8c50000;
      87076: inst = 32'h24612800;
      87077: inst = 32'h10a00000;
      87078: inst = 32'hca00006;
      87079: inst = 32'h24822800;
      87080: inst = 32'h10a00000;
      87081: inst = 32'hca00004;
      87082: inst = 32'h38632800;
      87083: inst = 32'h38842800;
      87084: inst = 32'h10a00001;
      87085: inst = 32'hca05431;
      87086: inst = 32'h13e00001;
      87087: inst = 32'hfe0d96a;
      87088: inst = 32'h5be00000;
      87089: inst = 32'h8c50000;
      87090: inst = 32'h24612800;
      87091: inst = 32'h10a00000;
      87092: inst = 32'hca00006;
      87093: inst = 32'h24822800;
      87094: inst = 32'h10a00000;
      87095: inst = 32'hca00004;
      87096: inst = 32'h38632800;
      87097: inst = 32'h38842800;
      87098: inst = 32'h10a00001;
      87099: inst = 32'hca0543f;
      87100: inst = 32'h13e00001;
      87101: inst = 32'hfe0d96a;
      87102: inst = 32'h5be00000;
      87103: inst = 32'h8c50000;
      87104: inst = 32'h24612800;
      87105: inst = 32'h10a00000;
      87106: inst = 32'hca00006;
      87107: inst = 32'h24822800;
      87108: inst = 32'h10a00000;
      87109: inst = 32'hca00004;
      87110: inst = 32'h38632800;
      87111: inst = 32'h38842800;
      87112: inst = 32'h10a00001;
      87113: inst = 32'hca0544d;
      87114: inst = 32'h13e00001;
      87115: inst = 32'hfe0d96a;
      87116: inst = 32'h5be00000;
      87117: inst = 32'h8c50000;
      87118: inst = 32'h24612800;
      87119: inst = 32'h10a00000;
      87120: inst = 32'hca00006;
      87121: inst = 32'h24822800;
      87122: inst = 32'h10a00000;
      87123: inst = 32'hca00004;
      87124: inst = 32'h38632800;
      87125: inst = 32'h38842800;
      87126: inst = 32'h10a00001;
      87127: inst = 32'hca0545b;
      87128: inst = 32'h13e00001;
      87129: inst = 32'hfe0d96a;
      87130: inst = 32'h5be00000;
      87131: inst = 32'h8c50000;
      87132: inst = 32'h24612800;
      87133: inst = 32'h10a00000;
      87134: inst = 32'hca00006;
      87135: inst = 32'h24822800;
      87136: inst = 32'h10a00000;
      87137: inst = 32'hca00004;
      87138: inst = 32'h38632800;
      87139: inst = 32'h38842800;
      87140: inst = 32'h10a00001;
      87141: inst = 32'hca05469;
      87142: inst = 32'h13e00001;
      87143: inst = 32'hfe0d96a;
      87144: inst = 32'h5be00000;
      87145: inst = 32'h8c50000;
      87146: inst = 32'h24612800;
      87147: inst = 32'h10a00000;
      87148: inst = 32'hca00006;
      87149: inst = 32'h24822800;
      87150: inst = 32'h10a00000;
      87151: inst = 32'hca00004;
      87152: inst = 32'h38632800;
      87153: inst = 32'h38842800;
      87154: inst = 32'h10a00001;
      87155: inst = 32'hca05477;
      87156: inst = 32'h13e00001;
      87157: inst = 32'hfe0d96a;
      87158: inst = 32'h5be00000;
      87159: inst = 32'h8c50000;
      87160: inst = 32'h24612800;
      87161: inst = 32'h10a00000;
      87162: inst = 32'hca00006;
      87163: inst = 32'h24822800;
      87164: inst = 32'h10a00000;
      87165: inst = 32'hca00004;
      87166: inst = 32'h38632800;
      87167: inst = 32'h38842800;
      87168: inst = 32'h10a00001;
      87169: inst = 32'hca05485;
      87170: inst = 32'h13e00001;
      87171: inst = 32'hfe0d96a;
      87172: inst = 32'h5be00000;
      87173: inst = 32'h8c50000;
      87174: inst = 32'h24612800;
      87175: inst = 32'h10a00000;
      87176: inst = 32'hca00006;
      87177: inst = 32'h24822800;
      87178: inst = 32'h10a00000;
      87179: inst = 32'hca00004;
      87180: inst = 32'h38632800;
      87181: inst = 32'h38842800;
      87182: inst = 32'h10a00001;
      87183: inst = 32'hca05493;
      87184: inst = 32'h13e00001;
      87185: inst = 32'hfe0d96a;
      87186: inst = 32'h5be00000;
      87187: inst = 32'h8c50000;
      87188: inst = 32'h24612800;
      87189: inst = 32'h10a00000;
      87190: inst = 32'hca00006;
      87191: inst = 32'h24822800;
      87192: inst = 32'h10a00000;
      87193: inst = 32'hca00004;
      87194: inst = 32'h38632800;
      87195: inst = 32'h38842800;
      87196: inst = 32'h10a00001;
      87197: inst = 32'hca054a1;
      87198: inst = 32'h13e00001;
      87199: inst = 32'hfe0d96a;
      87200: inst = 32'h5be00000;
      87201: inst = 32'h8c50000;
      87202: inst = 32'h24612800;
      87203: inst = 32'h10a00000;
      87204: inst = 32'hca00006;
      87205: inst = 32'h24822800;
      87206: inst = 32'h10a00000;
      87207: inst = 32'hca00004;
      87208: inst = 32'h38632800;
      87209: inst = 32'h38842800;
      87210: inst = 32'h10a00001;
      87211: inst = 32'hca054af;
      87212: inst = 32'h13e00001;
      87213: inst = 32'hfe0d96a;
      87214: inst = 32'h5be00000;
      87215: inst = 32'h8c50000;
      87216: inst = 32'h24612800;
      87217: inst = 32'h10a00000;
      87218: inst = 32'hca00006;
      87219: inst = 32'h24822800;
      87220: inst = 32'h10a00000;
      87221: inst = 32'hca00004;
      87222: inst = 32'h38632800;
      87223: inst = 32'h38842800;
      87224: inst = 32'h10a00001;
      87225: inst = 32'hca054bd;
      87226: inst = 32'h13e00001;
      87227: inst = 32'hfe0d96a;
      87228: inst = 32'h5be00000;
      87229: inst = 32'h8c50000;
      87230: inst = 32'h24612800;
      87231: inst = 32'h10a00000;
      87232: inst = 32'hca00006;
      87233: inst = 32'h24822800;
      87234: inst = 32'h10a00000;
      87235: inst = 32'hca00004;
      87236: inst = 32'h38632800;
      87237: inst = 32'h38842800;
      87238: inst = 32'h10a00001;
      87239: inst = 32'hca054cb;
      87240: inst = 32'h13e00001;
      87241: inst = 32'hfe0d96a;
      87242: inst = 32'h5be00000;
      87243: inst = 32'h8c50000;
      87244: inst = 32'h24612800;
      87245: inst = 32'h10a00000;
      87246: inst = 32'hca00006;
      87247: inst = 32'h24822800;
      87248: inst = 32'h10a00000;
      87249: inst = 32'hca00004;
      87250: inst = 32'h38632800;
      87251: inst = 32'h38842800;
      87252: inst = 32'h10a00001;
      87253: inst = 32'hca054d9;
      87254: inst = 32'h13e00001;
      87255: inst = 32'hfe0d96a;
      87256: inst = 32'h5be00000;
      87257: inst = 32'h8c50000;
      87258: inst = 32'h24612800;
      87259: inst = 32'h10a00000;
      87260: inst = 32'hca00006;
      87261: inst = 32'h24822800;
      87262: inst = 32'h10a00000;
      87263: inst = 32'hca00004;
      87264: inst = 32'h38632800;
      87265: inst = 32'h38842800;
      87266: inst = 32'h10a00001;
      87267: inst = 32'hca054e7;
      87268: inst = 32'h13e00001;
      87269: inst = 32'hfe0d96a;
      87270: inst = 32'h5be00000;
      87271: inst = 32'h8c50000;
      87272: inst = 32'h24612800;
      87273: inst = 32'h10a00000;
      87274: inst = 32'hca00006;
      87275: inst = 32'h24822800;
      87276: inst = 32'h10a00000;
      87277: inst = 32'hca00004;
      87278: inst = 32'h38632800;
      87279: inst = 32'h38842800;
      87280: inst = 32'h10a00001;
      87281: inst = 32'hca054f5;
      87282: inst = 32'h13e00001;
      87283: inst = 32'hfe0d96a;
      87284: inst = 32'h5be00000;
      87285: inst = 32'h8c50000;
      87286: inst = 32'h24612800;
      87287: inst = 32'h10a00000;
      87288: inst = 32'hca00006;
      87289: inst = 32'h24822800;
      87290: inst = 32'h10a00000;
      87291: inst = 32'hca00004;
      87292: inst = 32'h38632800;
      87293: inst = 32'h38842800;
      87294: inst = 32'h10a00001;
      87295: inst = 32'hca05503;
      87296: inst = 32'h13e00001;
      87297: inst = 32'hfe0d96a;
      87298: inst = 32'h5be00000;
      87299: inst = 32'h8c50000;
      87300: inst = 32'h24612800;
      87301: inst = 32'h10a00000;
      87302: inst = 32'hca00006;
      87303: inst = 32'h24822800;
      87304: inst = 32'h10a00000;
      87305: inst = 32'hca00004;
      87306: inst = 32'h38632800;
      87307: inst = 32'h38842800;
      87308: inst = 32'h10a00001;
      87309: inst = 32'hca05511;
      87310: inst = 32'h13e00001;
      87311: inst = 32'hfe0d96a;
      87312: inst = 32'h5be00000;
      87313: inst = 32'h8c50000;
      87314: inst = 32'h24612800;
      87315: inst = 32'h10a00000;
      87316: inst = 32'hca00006;
      87317: inst = 32'h24822800;
      87318: inst = 32'h10a00000;
      87319: inst = 32'hca00004;
      87320: inst = 32'h38632800;
      87321: inst = 32'h38842800;
      87322: inst = 32'h10a00001;
      87323: inst = 32'hca0551f;
      87324: inst = 32'h13e00001;
      87325: inst = 32'hfe0d96a;
      87326: inst = 32'h5be00000;
      87327: inst = 32'h8c50000;
      87328: inst = 32'h24612800;
      87329: inst = 32'h10a00000;
      87330: inst = 32'hca00006;
      87331: inst = 32'h24822800;
      87332: inst = 32'h10a00000;
      87333: inst = 32'hca00004;
      87334: inst = 32'h38632800;
      87335: inst = 32'h38842800;
      87336: inst = 32'h10a00001;
      87337: inst = 32'hca0552d;
      87338: inst = 32'h13e00001;
      87339: inst = 32'hfe0d96a;
      87340: inst = 32'h5be00000;
      87341: inst = 32'h8c50000;
      87342: inst = 32'h24612800;
      87343: inst = 32'h10a00000;
      87344: inst = 32'hca00006;
      87345: inst = 32'h24822800;
      87346: inst = 32'h10a00000;
      87347: inst = 32'hca00004;
      87348: inst = 32'h38632800;
      87349: inst = 32'h38842800;
      87350: inst = 32'h10a00001;
      87351: inst = 32'hca0553b;
      87352: inst = 32'h13e00001;
      87353: inst = 32'hfe0d96a;
      87354: inst = 32'h5be00000;
      87355: inst = 32'h8c50000;
      87356: inst = 32'h24612800;
      87357: inst = 32'h10a00000;
      87358: inst = 32'hca00006;
      87359: inst = 32'h24822800;
      87360: inst = 32'h10a00000;
      87361: inst = 32'hca00004;
      87362: inst = 32'h38632800;
      87363: inst = 32'h38842800;
      87364: inst = 32'h10a00001;
      87365: inst = 32'hca05549;
      87366: inst = 32'h13e00001;
      87367: inst = 32'hfe0d96a;
      87368: inst = 32'h5be00000;
      87369: inst = 32'h8c50000;
      87370: inst = 32'h24612800;
      87371: inst = 32'h10a00000;
      87372: inst = 32'hca00006;
      87373: inst = 32'h24822800;
      87374: inst = 32'h10a00000;
      87375: inst = 32'hca00004;
      87376: inst = 32'h38632800;
      87377: inst = 32'h38842800;
      87378: inst = 32'h10a00001;
      87379: inst = 32'hca05557;
      87380: inst = 32'h13e00001;
      87381: inst = 32'hfe0d96a;
      87382: inst = 32'h5be00000;
      87383: inst = 32'h8c50000;
      87384: inst = 32'h24612800;
      87385: inst = 32'h10a00000;
      87386: inst = 32'hca00006;
      87387: inst = 32'h24822800;
      87388: inst = 32'h10a00000;
      87389: inst = 32'hca00004;
      87390: inst = 32'h38632800;
      87391: inst = 32'h38842800;
      87392: inst = 32'h10a00001;
      87393: inst = 32'hca05565;
      87394: inst = 32'h13e00001;
      87395: inst = 32'hfe0d96a;
      87396: inst = 32'h5be00000;
      87397: inst = 32'h8c50000;
      87398: inst = 32'h24612800;
      87399: inst = 32'h10a00000;
      87400: inst = 32'hca00006;
      87401: inst = 32'h24822800;
      87402: inst = 32'h10a00000;
      87403: inst = 32'hca00004;
      87404: inst = 32'h38632800;
      87405: inst = 32'h38842800;
      87406: inst = 32'h10a00001;
      87407: inst = 32'hca05573;
      87408: inst = 32'h13e00001;
      87409: inst = 32'hfe0d96a;
      87410: inst = 32'h5be00000;
      87411: inst = 32'h8c50000;
      87412: inst = 32'h24612800;
      87413: inst = 32'h10a00000;
      87414: inst = 32'hca00006;
      87415: inst = 32'h24822800;
      87416: inst = 32'h10a00000;
      87417: inst = 32'hca00004;
      87418: inst = 32'h38632800;
      87419: inst = 32'h38842800;
      87420: inst = 32'h10a00001;
      87421: inst = 32'hca05581;
      87422: inst = 32'h13e00001;
      87423: inst = 32'hfe0d96a;
      87424: inst = 32'h5be00000;
      87425: inst = 32'h8c50000;
      87426: inst = 32'h24612800;
      87427: inst = 32'h10a00000;
      87428: inst = 32'hca00006;
      87429: inst = 32'h24822800;
      87430: inst = 32'h10a00000;
      87431: inst = 32'hca00004;
      87432: inst = 32'h38632800;
      87433: inst = 32'h38842800;
      87434: inst = 32'h10a00001;
      87435: inst = 32'hca0558f;
      87436: inst = 32'h13e00001;
      87437: inst = 32'hfe0d96a;
      87438: inst = 32'h5be00000;
      87439: inst = 32'h8c50000;
      87440: inst = 32'h24612800;
      87441: inst = 32'h10a00000;
      87442: inst = 32'hca00006;
      87443: inst = 32'h24822800;
      87444: inst = 32'h10a00000;
      87445: inst = 32'hca00004;
      87446: inst = 32'h38632800;
      87447: inst = 32'h38842800;
      87448: inst = 32'h10a00001;
      87449: inst = 32'hca0559d;
      87450: inst = 32'h13e00001;
      87451: inst = 32'hfe0d96a;
      87452: inst = 32'h5be00000;
      87453: inst = 32'h8c50000;
      87454: inst = 32'h24612800;
      87455: inst = 32'h10a00000;
      87456: inst = 32'hca00006;
      87457: inst = 32'h24822800;
      87458: inst = 32'h10a00000;
      87459: inst = 32'hca00004;
      87460: inst = 32'h38632800;
      87461: inst = 32'h38842800;
      87462: inst = 32'h10a00001;
      87463: inst = 32'hca055ab;
      87464: inst = 32'h13e00001;
      87465: inst = 32'hfe0d96a;
      87466: inst = 32'h5be00000;
      87467: inst = 32'h8c50000;
      87468: inst = 32'h24612800;
      87469: inst = 32'h10a00000;
      87470: inst = 32'hca00006;
      87471: inst = 32'h24822800;
      87472: inst = 32'h10a00000;
      87473: inst = 32'hca00004;
      87474: inst = 32'h38632800;
      87475: inst = 32'h38842800;
      87476: inst = 32'h10a00001;
      87477: inst = 32'hca055b9;
      87478: inst = 32'h13e00001;
      87479: inst = 32'hfe0d96a;
      87480: inst = 32'h5be00000;
      87481: inst = 32'h8c50000;
      87482: inst = 32'h24612800;
      87483: inst = 32'h10a00000;
      87484: inst = 32'hca00006;
      87485: inst = 32'h24822800;
      87486: inst = 32'h10a00000;
      87487: inst = 32'hca00004;
      87488: inst = 32'h38632800;
      87489: inst = 32'h38842800;
      87490: inst = 32'h10a00001;
      87491: inst = 32'hca055c7;
      87492: inst = 32'h13e00001;
      87493: inst = 32'hfe0d96a;
      87494: inst = 32'h5be00000;
      87495: inst = 32'h8c50000;
      87496: inst = 32'h24612800;
      87497: inst = 32'h10a00000;
      87498: inst = 32'hca00006;
      87499: inst = 32'h24822800;
      87500: inst = 32'h10a00000;
      87501: inst = 32'hca00004;
      87502: inst = 32'h38632800;
      87503: inst = 32'h38842800;
      87504: inst = 32'h10a00001;
      87505: inst = 32'hca055d5;
      87506: inst = 32'h13e00001;
      87507: inst = 32'hfe0d96a;
      87508: inst = 32'h5be00000;
      87509: inst = 32'h8c50000;
      87510: inst = 32'h24612800;
      87511: inst = 32'h10a00000;
      87512: inst = 32'hca00006;
      87513: inst = 32'h24822800;
      87514: inst = 32'h10a00000;
      87515: inst = 32'hca00004;
      87516: inst = 32'h38632800;
      87517: inst = 32'h38842800;
      87518: inst = 32'h10a00001;
      87519: inst = 32'hca055e3;
      87520: inst = 32'h13e00001;
      87521: inst = 32'hfe0d96a;
      87522: inst = 32'h5be00000;
      87523: inst = 32'h8c50000;
      87524: inst = 32'h24612800;
      87525: inst = 32'h10a00000;
      87526: inst = 32'hca00006;
      87527: inst = 32'h24822800;
      87528: inst = 32'h10a00000;
      87529: inst = 32'hca00004;
      87530: inst = 32'h38632800;
      87531: inst = 32'h38842800;
      87532: inst = 32'h10a00001;
      87533: inst = 32'hca055f1;
      87534: inst = 32'h13e00001;
      87535: inst = 32'hfe0d96a;
      87536: inst = 32'h5be00000;
      87537: inst = 32'h8c50000;
      87538: inst = 32'h24612800;
      87539: inst = 32'h10a00000;
      87540: inst = 32'hca00006;
      87541: inst = 32'h24822800;
      87542: inst = 32'h10a00000;
      87543: inst = 32'hca00004;
      87544: inst = 32'h38632800;
      87545: inst = 32'h38842800;
      87546: inst = 32'h10a00001;
      87547: inst = 32'hca055ff;
      87548: inst = 32'h13e00001;
      87549: inst = 32'hfe0d96a;
      87550: inst = 32'h5be00000;
      87551: inst = 32'h8c50000;
      87552: inst = 32'h24612800;
      87553: inst = 32'h10a00000;
      87554: inst = 32'hca00006;
      87555: inst = 32'h24822800;
      87556: inst = 32'h10a00000;
      87557: inst = 32'hca00004;
      87558: inst = 32'h38632800;
      87559: inst = 32'h38842800;
      87560: inst = 32'h10a00001;
      87561: inst = 32'hca0560d;
      87562: inst = 32'h13e00001;
      87563: inst = 32'hfe0d96a;
      87564: inst = 32'h5be00000;
      87565: inst = 32'h8c50000;
      87566: inst = 32'h24612800;
      87567: inst = 32'h10a00000;
      87568: inst = 32'hca00006;
      87569: inst = 32'h24822800;
      87570: inst = 32'h10a00000;
      87571: inst = 32'hca00004;
      87572: inst = 32'h38632800;
      87573: inst = 32'h38842800;
      87574: inst = 32'h10a00001;
      87575: inst = 32'hca0561b;
      87576: inst = 32'h13e00001;
      87577: inst = 32'hfe0d96a;
      87578: inst = 32'h5be00000;
      87579: inst = 32'h8c50000;
      87580: inst = 32'h24612800;
      87581: inst = 32'h10a00000;
      87582: inst = 32'hca00006;
      87583: inst = 32'h24822800;
      87584: inst = 32'h10a00000;
      87585: inst = 32'hca00004;
      87586: inst = 32'h38632800;
      87587: inst = 32'h38842800;
      87588: inst = 32'h10a00001;
      87589: inst = 32'hca05629;
      87590: inst = 32'h13e00001;
      87591: inst = 32'hfe0d96a;
      87592: inst = 32'h5be00000;
      87593: inst = 32'h8c50000;
      87594: inst = 32'h24612800;
      87595: inst = 32'h10a00000;
      87596: inst = 32'hca00007;
      87597: inst = 32'h24822800;
      87598: inst = 32'h10a00000;
      87599: inst = 32'hca00004;
      87600: inst = 32'h38632800;
      87601: inst = 32'h38842800;
      87602: inst = 32'h10a00001;
      87603: inst = 32'hca05637;
      87604: inst = 32'h13e00001;
      87605: inst = 32'hfe0d96a;
      87606: inst = 32'h5be00000;
      87607: inst = 32'h8c50000;
      87608: inst = 32'h24612800;
      87609: inst = 32'h10a00000;
      87610: inst = 32'hca00007;
      87611: inst = 32'h24822800;
      87612: inst = 32'h10a00000;
      87613: inst = 32'hca00004;
      87614: inst = 32'h38632800;
      87615: inst = 32'h38842800;
      87616: inst = 32'h10a00001;
      87617: inst = 32'hca05645;
      87618: inst = 32'h13e00001;
      87619: inst = 32'hfe0d96a;
      87620: inst = 32'h5be00000;
      87621: inst = 32'h8c50000;
      87622: inst = 32'h24612800;
      87623: inst = 32'h10a00000;
      87624: inst = 32'hca00007;
      87625: inst = 32'h24822800;
      87626: inst = 32'h10a00000;
      87627: inst = 32'hca00004;
      87628: inst = 32'h38632800;
      87629: inst = 32'h38842800;
      87630: inst = 32'h10a00001;
      87631: inst = 32'hca05653;
      87632: inst = 32'h13e00001;
      87633: inst = 32'hfe0d96a;
      87634: inst = 32'h5be00000;
      87635: inst = 32'h8c50000;
      87636: inst = 32'h24612800;
      87637: inst = 32'h10a00000;
      87638: inst = 32'hca00007;
      87639: inst = 32'h24822800;
      87640: inst = 32'h10a00000;
      87641: inst = 32'hca00004;
      87642: inst = 32'h38632800;
      87643: inst = 32'h38842800;
      87644: inst = 32'h10a00001;
      87645: inst = 32'hca05661;
      87646: inst = 32'h13e00001;
      87647: inst = 32'hfe0d96a;
      87648: inst = 32'h5be00000;
      87649: inst = 32'h8c50000;
      87650: inst = 32'h24612800;
      87651: inst = 32'h10a00000;
      87652: inst = 32'hca00007;
      87653: inst = 32'h24822800;
      87654: inst = 32'h10a00000;
      87655: inst = 32'hca00004;
      87656: inst = 32'h38632800;
      87657: inst = 32'h38842800;
      87658: inst = 32'h10a00001;
      87659: inst = 32'hca0566f;
      87660: inst = 32'h13e00001;
      87661: inst = 32'hfe0d96a;
      87662: inst = 32'h5be00000;
      87663: inst = 32'h8c50000;
      87664: inst = 32'h24612800;
      87665: inst = 32'h10a00000;
      87666: inst = 32'hca00007;
      87667: inst = 32'h24822800;
      87668: inst = 32'h10a00000;
      87669: inst = 32'hca00004;
      87670: inst = 32'h38632800;
      87671: inst = 32'h38842800;
      87672: inst = 32'h10a00001;
      87673: inst = 32'hca0567d;
      87674: inst = 32'h13e00001;
      87675: inst = 32'hfe0d96a;
      87676: inst = 32'h5be00000;
      87677: inst = 32'h8c50000;
      87678: inst = 32'h24612800;
      87679: inst = 32'h10a00000;
      87680: inst = 32'hca00007;
      87681: inst = 32'h24822800;
      87682: inst = 32'h10a00000;
      87683: inst = 32'hca00004;
      87684: inst = 32'h38632800;
      87685: inst = 32'h38842800;
      87686: inst = 32'h10a00001;
      87687: inst = 32'hca0568b;
      87688: inst = 32'h13e00001;
      87689: inst = 32'hfe0d96a;
      87690: inst = 32'h5be00000;
      87691: inst = 32'h8c50000;
      87692: inst = 32'h24612800;
      87693: inst = 32'h10a00000;
      87694: inst = 32'hca00007;
      87695: inst = 32'h24822800;
      87696: inst = 32'h10a00000;
      87697: inst = 32'hca00004;
      87698: inst = 32'h38632800;
      87699: inst = 32'h38842800;
      87700: inst = 32'h10a00001;
      87701: inst = 32'hca05699;
      87702: inst = 32'h13e00001;
      87703: inst = 32'hfe0d96a;
      87704: inst = 32'h5be00000;
      87705: inst = 32'h8c50000;
      87706: inst = 32'h24612800;
      87707: inst = 32'h10a00000;
      87708: inst = 32'hca00007;
      87709: inst = 32'h24822800;
      87710: inst = 32'h10a00000;
      87711: inst = 32'hca00004;
      87712: inst = 32'h38632800;
      87713: inst = 32'h38842800;
      87714: inst = 32'h10a00001;
      87715: inst = 32'hca056a7;
      87716: inst = 32'h13e00001;
      87717: inst = 32'hfe0d96a;
      87718: inst = 32'h5be00000;
      87719: inst = 32'h8c50000;
      87720: inst = 32'h24612800;
      87721: inst = 32'h10a00000;
      87722: inst = 32'hca00007;
      87723: inst = 32'h24822800;
      87724: inst = 32'h10a00000;
      87725: inst = 32'hca00004;
      87726: inst = 32'h38632800;
      87727: inst = 32'h38842800;
      87728: inst = 32'h10a00001;
      87729: inst = 32'hca056b5;
      87730: inst = 32'h13e00001;
      87731: inst = 32'hfe0d96a;
      87732: inst = 32'h5be00000;
      87733: inst = 32'h8c50000;
      87734: inst = 32'h24612800;
      87735: inst = 32'h10a00000;
      87736: inst = 32'hca00007;
      87737: inst = 32'h24822800;
      87738: inst = 32'h10a00000;
      87739: inst = 32'hca00004;
      87740: inst = 32'h38632800;
      87741: inst = 32'h38842800;
      87742: inst = 32'h10a00001;
      87743: inst = 32'hca056c3;
      87744: inst = 32'h13e00001;
      87745: inst = 32'hfe0d96a;
      87746: inst = 32'h5be00000;
      87747: inst = 32'h8c50000;
      87748: inst = 32'h24612800;
      87749: inst = 32'h10a00000;
      87750: inst = 32'hca00007;
      87751: inst = 32'h24822800;
      87752: inst = 32'h10a00000;
      87753: inst = 32'hca00004;
      87754: inst = 32'h38632800;
      87755: inst = 32'h38842800;
      87756: inst = 32'h10a00001;
      87757: inst = 32'hca056d1;
      87758: inst = 32'h13e00001;
      87759: inst = 32'hfe0d96a;
      87760: inst = 32'h5be00000;
      87761: inst = 32'h8c50000;
      87762: inst = 32'h24612800;
      87763: inst = 32'h10a00000;
      87764: inst = 32'hca00007;
      87765: inst = 32'h24822800;
      87766: inst = 32'h10a00000;
      87767: inst = 32'hca00004;
      87768: inst = 32'h38632800;
      87769: inst = 32'h38842800;
      87770: inst = 32'h10a00001;
      87771: inst = 32'hca056df;
      87772: inst = 32'h13e00001;
      87773: inst = 32'hfe0d96a;
      87774: inst = 32'h5be00000;
      87775: inst = 32'h8c50000;
      87776: inst = 32'h24612800;
      87777: inst = 32'h10a00000;
      87778: inst = 32'hca00007;
      87779: inst = 32'h24822800;
      87780: inst = 32'h10a00000;
      87781: inst = 32'hca00004;
      87782: inst = 32'h38632800;
      87783: inst = 32'h38842800;
      87784: inst = 32'h10a00001;
      87785: inst = 32'hca056ed;
      87786: inst = 32'h13e00001;
      87787: inst = 32'hfe0d96a;
      87788: inst = 32'h5be00000;
      87789: inst = 32'h8c50000;
      87790: inst = 32'h24612800;
      87791: inst = 32'h10a00000;
      87792: inst = 32'hca00007;
      87793: inst = 32'h24822800;
      87794: inst = 32'h10a00000;
      87795: inst = 32'hca00004;
      87796: inst = 32'h38632800;
      87797: inst = 32'h38842800;
      87798: inst = 32'h10a00001;
      87799: inst = 32'hca056fb;
      87800: inst = 32'h13e00001;
      87801: inst = 32'hfe0d96a;
      87802: inst = 32'h5be00000;
      87803: inst = 32'h8c50000;
      87804: inst = 32'h24612800;
      87805: inst = 32'h10a00000;
      87806: inst = 32'hca00007;
      87807: inst = 32'h24822800;
      87808: inst = 32'h10a00000;
      87809: inst = 32'hca00004;
      87810: inst = 32'h38632800;
      87811: inst = 32'h38842800;
      87812: inst = 32'h10a00001;
      87813: inst = 32'hca05709;
      87814: inst = 32'h13e00001;
      87815: inst = 32'hfe0d96a;
      87816: inst = 32'h5be00000;
      87817: inst = 32'h8c50000;
      87818: inst = 32'h24612800;
      87819: inst = 32'h10a00000;
      87820: inst = 32'hca00007;
      87821: inst = 32'h24822800;
      87822: inst = 32'h10a00000;
      87823: inst = 32'hca00004;
      87824: inst = 32'h38632800;
      87825: inst = 32'h38842800;
      87826: inst = 32'h10a00001;
      87827: inst = 32'hca05717;
      87828: inst = 32'h13e00001;
      87829: inst = 32'hfe0d96a;
      87830: inst = 32'h5be00000;
      87831: inst = 32'h8c50000;
      87832: inst = 32'h24612800;
      87833: inst = 32'h10a00000;
      87834: inst = 32'hca00007;
      87835: inst = 32'h24822800;
      87836: inst = 32'h10a00000;
      87837: inst = 32'hca00004;
      87838: inst = 32'h38632800;
      87839: inst = 32'h38842800;
      87840: inst = 32'h10a00001;
      87841: inst = 32'hca05725;
      87842: inst = 32'h13e00001;
      87843: inst = 32'hfe0d96a;
      87844: inst = 32'h5be00000;
      87845: inst = 32'h8c50000;
      87846: inst = 32'h24612800;
      87847: inst = 32'h10a00000;
      87848: inst = 32'hca00007;
      87849: inst = 32'h24822800;
      87850: inst = 32'h10a00000;
      87851: inst = 32'hca00004;
      87852: inst = 32'h38632800;
      87853: inst = 32'h38842800;
      87854: inst = 32'h10a00001;
      87855: inst = 32'hca05733;
      87856: inst = 32'h13e00001;
      87857: inst = 32'hfe0d96a;
      87858: inst = 32'h5be00000;
      87859: inst = 32'h8c50000;
      87860: inst = 32'h24612800;
      87861: inst = 32'h10a00000;
      87862: inst = 32'hca00007;
      87863: inst = 32'h24822800;
      87864: inst = 32'h10a00000;
      87865: inst = 32'hca00004;
      87866: inst = 32'h38632800;
      87867: inst = 32'h38842800;
      87868: inst = 32'h10a00001;
      87869: inst = 32'hca05741;
      87870: inst = 32'h13e00001;
      87871: inst = 32'hfe0d96a;
      87872: inst = 32'h5be00000;
      87873: inst = 32'h8c50000;
      87874: inst = 32'h24612800;
      87875: inst = 32'h10a00000;
      87876: inst = 32'hca00007;
      87877: inst = 32'h24822800;
      87878: inst = 32'h10a00000;
      87879: inst = 32'hca00004;
      87880: inst = 32'h38632800;
      87881: inst = 32'h38842800;
      87882: inst = 32'h10a00001;
      87883: inst = 32'hca0574f;
      87884: inst = 32'h13e00001;
      87885: inst = 32'hfe0d96a;
      87886: inst = 32'h5be00000;
      87887: inst = 32'h8c50000;
      87888: inst = 32'h24612800;
      87889: inst = 32'h10a00000;
      87890: inst = 32'hca00007;
      87891: inst = 32'h24822800;
      87892: inst = 32'h10a00000;
      87893: inst = 32'hca00004;
      87894: inst = 32'h38632800;
      87895: inst = 32'h38842800;
      87896: inst = 32'h10a00001;
      87897: inst = 32'hca0575d;
      87898: inst = 32'h13e00001;
      87899: inst = 32'hfe0d96a;
      87900: inst = 32'h5be00000;
      87901: inst = 32'h8c50000;
      87902: inst = 32'h24612800;
      87903: inst = 32'h10a00000;
      87904: inst = 32'hca00007;
      87905: inst = 32'h24822800;
      87906: inst = 32'h10a00000;
      87907: inst = 32'hca00004;
      87908: inst = 32'h38632800;
      87909: inst = 32'h38842800;
      87910: inst = 32'h10a00001;
      87911: inst = 32'hca0576b;
      87912: inst = 32'h13e00001;
      87913: inst = 32'hfe0d96a;
      87914: inst = 32'h5be00000;
      87915: inst = 32'h8c50000;
      87916: inst = 32'h24612800;
      87917: inst = 32'h10a00000;
      87918: inst = 32'hca00007;
      87919: inst = 32'h24822800;
      87920: inst = 32'h10a00000;
      87921: inst = 32'hca00004;
      87922: inst = 32'h38632800;
      87923: inst = 32'h38842800;
      87924: inst = 32'h10a00001;
      87925: inst = 32'hca05779;
      87926: inst = 32'h13e00001;
      87927: inst = 32'hfe0d96a;
      87928: inst = 32'h5be00000;
      87929: inst = 32'h8c50000;
      87930: inst = 32'h24612800;
      87931: inst = 32'h10a00000;
      87932: inst = 32'hca00007;
      87933: inst = 32'h24822800;
      87934: inst = 32'h10a00000;
      87935: inst = 32'hca00004;
      87936: inst = 32'h38632800;
      87937: inst = 32'h38842800;
      87938: inst = 32'h10a00001;
      87939: inst = 32'hca05787;
      87940: inst = 32'h13e00001;
      87941: inst = 32'hfe0d96a;
      87942: inst = 32'h5be00000;
      87943: inst = 32'h8c50000;
      87944: inst = 32'h24612800;
      87945: inst = 32'h10a00000;
      87946: inst = 32'hca00007;
      87947: inst = 32'h24822800;
      87948: inst = 32'h10a00000;
      87949: inst = 32'hca00004;
      87950: inst = 32'h38632800;
      87951: inst = 32'h38842800;
      87952: inst = 32'h10a00001;
      87953: inst = 32'hca05795;
      87954: inst = 32'h13e00001;
      87955: inst = 32'hfe0d96a;
      87956: inst = 32'h5be00000;
      87957: inst = 32'h8c50000;
      87958: inst = 32'h24612800;
      87959: inst = 32'h10a00000;
      87960: inst = 32'hca00007;
      87961: inst = 32'h24822800;
      87962: inst = 32'h10a00000;
      87963: inst = 32'hca00004;
      87964: inst = 32'h38632800;
      87965: inst = 32'h38842800;
      87966: inst = 32'h10a00001;
      87967: inst = 32'hca057a3;
      87968: inst = 32'h13e00001;
      87969: inst = 32'hfe0d96a;
      87970: inst = 32'h5be00000;
      87971: inst = 32'h8c50000;
      87972: inst = 32'h24612800;
      87973: inst = 32'h10a00000;
      87974: inst = 32'hca00007;
      87975: inst = 32'h24822800;
      87976: inst = 32'h10a00000;
      87977: inst = 32'hca00004;
      87978: inst = 32'h38632800;
      87979: inst = 32'h38842800;
      87980: inst = 32'h10a00001;
      87981: inst = 32'hca057b1;
      87982: inst = 32'h13e00001;
      87983: inst = 32'hfe0d96a;
      87984: inst = 32'h5be00000;
      87985: inst = 32'h8c50000;
      87986: inst = 32'h24612800;
      87987: inst = 32'h10a00000;
      87988: inst = 32'hca00007;
      87989: inst = 32'h24822800;
      87990: inst = 32'h10a00000;
      87991: inst = 32'hca00004;
      87992: inst = 32'h38632800;
      87993: inst = 32'h38842800;
      87994: inst = 32'h10a00001;
      87995: inst = 32'hca057bf;
      87996: inst = 32'h13e00001;
      87997: inst = 32'hfe0d96a;
      87998: inst = 32'h5be00000;
      87999: inst = 32'h8c50000;
      88000: inst = 32'h24612800;
      88001: inst = 32'h10a00000;
      88002: inst = 32'hca00007;
      88003: inst = 32'h24822800;
      88004: inst = 32'h10a00000;
      88005: inst = 32'hca00004;
      88006: inst = 32'h38632800;
      88007: inst = 32'h38842800;
      88008: inst = 32'h10a00001;
      88009: inst = 32'hca057cd;
      88010: inst = 32'h13e00001;
      88011: inst = 32'hfe0d96a;
      88012: inst = 32'h5be00000;
      88013: inst = 32'h8c50000;
      88014: inst = 32'h24612800;
      88015: inst = 32'h10a00000;
      88016: inst = 32'hca00007;
      88017: inst = 32'h24822800;
      88018: inst = 32'h10a00000;
      88019: inst = 32'hca00004;
      88020: inst = 32'h38632800;
      88021: inst = 32'h38842800;
      88022: inst = 32'h10a00001;
      88023: inst = 32'hca057db;
      88024: inst = 32'h13e00001;
      88025: inst = 32'hfe0d96a;
      88026: inst = 32'h5be00000;
      88027: inst = 32'h8c50000;
      88028: inst = 32'h24612800;
      88029: inst = 32'h10a00000;
      88030: inst = 32'hca00007;
      88031: inst = 32'h24822800;
      88032: inst = 32'h10a00000;
      88033: inst = 32'hca00004;
      88034: inst = 32'h38632800;
      88035: inst = 32'h38842800;
      88036: inst = 32'h10a00001;
      88037: inst = 32'hca057e9;
      88038: inst = 32'h13e00001;
      88039: inst = 32'hfe0d96a;
      88040: inst = 32'h5be00000;
      88041: inst = 32'h8c50000;
      88042: inst = 32'h24612800;
      88043: inst = 32'h10a00000;
      88044: inst = 32'hca00007;
      88045: inst = 32'h24822800;
      88046: inst = 32'h10a00000;
      88047: inst = 32'hca00004;
      88048: inst = 32'h38632800;
      88049: inst = 32'h38842800;
      88050: inst = 32'h10a00001;
      88051: inst = 32'hca057f7;
      88052: inst = 32'h13e00001;
      88053: inst = 32'hfe0d96a;
      88054: inst = 32'h5be00000;
      88055: inst = 32'h8c50000;
      88056: inst = 32'h24612800;
      88057: inst = 32'h10a00000;
      88058: inst = 32'hca00007;
      88059: inst = 32'h24822800;
      88060: inst = 32'h10a00000;
      88061: inst = 32'hca00004;
      88062: inst = 32'h38632800;
      88063: inst = 32'h38842800;
      88064: inst = 32'h10a00001;
      88065: inst = 32'hca05805;
      88066: inst = 32'h13e00001;
      88067: inst = 32'hfe0d96a;
      88068: inst = 32'h5be00000;
      88069: inst = 32'h8c50000;
      88070: inst = 32'h24612800;
      88071: inst = 32'h10a00000;
      88072: inst = 32'hca00007;
      88073: inst = 32'h24822800;
      88074: inst = 32'h10a00000;
      88075: inst = 32'hca00004;
      88076: inst = 32'h38632800;
      88077: inst = 32'h38842800;
      88078: inst = 32'h10a00001;
      88079: inst = 32'hca05813;
      88080: inst = 32'h13e00001;
      88081: inst = 32'hfe0d96a;
      88082: inst = 32'h5be00000;
      88083: inst = 32'h8c50000;
      88084: inst = 32'h24612800;
      88085: inst = 32'h10a00000;
      88086: inst = 32'hca00007;
      88087: inst = 32'h24822800;
      88088: inst = 32'h10a00000;
      88089: inst = 32'hca00004;
      88090: inst = 32'h38632800;
      88091: inst = 32'h38842800;
      88092: inst = 32'h10a00001;
      88093: inst = 32'hca05821;
      88094: inst = 32'h13e00001;
      88095: inst = 32'hfe0d96a;
      88096: inst = 32'h5be00000;
      88097: inst = 32'h8c50000;
      88098: inst = 32'h24612800;
      88099: inst = 32'h10a00000;
      88100: inst = 32'hca00007;
      88101: inst = 32'h24822800;
      88102: inst = 32'h10a00000;
      88103: inst = 32'hca00004;
      88104: inst = 32'h38632800;
      88105: inst = 32'h38842800;
      88106: inst = 32'h10a00001;
      88107: inst = 32'hca0582f;
      88108: inst = 32'h13e00001;
      88109: inst = 32'hfe0d96a;
      88110: inst = 32'h5be00000;
      88111: inst = 32'h8c50000;
      88112: inst = 32'h24612800;
      88113: inst = 32'h10a00000;
      88114: inst = 32'hca00007;
      88115: inst = 32'h24822800;
      88116: inst = 32'h10a00000;
      88117: inst = 32'hca00004;
      88118: inst = 32'h38632800;
      88119: inst = 32'h38842800;
      88120: inst = 32'h10a00001;
      88121: inst = 32'hca0583d;
      88122: inst = 32'h13e00001;
      88123: inst = 32'hfe0d96a;
      88124: inst = 32'h5be00000;
      88125: inst = 32'h8c50000;
      88126: inst = 32'h24612800;
      88127: inst = 32'h10a00000;
      88128: inst = 32'hca00007;
      88129: inst = 32'h24822800;
      88130: inst = 32'h10a00000;
      88131: inst = 32'hca00004;
      88132: inst = 32'h38632800;
      88133: inst = 32'h38842800;
      88134: inst = 32'h10a00001;
      88135: inst = 32'hca0584b;
      88136: inst = 32'h13e00001;
      88137: inst = 32'hfe0d96a;
      88138: inst = 32'h5be00000;
      88139: inst = 32'h8c50000;
      88140: inst = 32'h24612800;
      88141: inst = 32'h10a00000;
      88142: inst = 32'hca00007;
      88143: inst = 32'h24822800;
      88144: inst = 32'h10a00000;
      88145: inst = 32'hca00004;
      88146: inst = 32'h38632800;
      88147: inst = 32'h38842800;
      88148: inst = 32'h10a00001;
      88149: inst = 32'hca05859;
      88150: inst = 32'h13e00001;
      88151: inst = 32'hfe0d96a;
      88152: inst = 32'h5be00000;
      88153: inst = 32'h8c50000;
      88154: inst = 32'h24612800;
      88155: inst = 32'h10a00000;
      88156: inst = 32'hca00007;
      88157: inst = 32'h24822800;
      88158: inst = 32'h10a00000;
      88159: inst = 32'hca00004;
      88160: inst = 32'h38632800;
      88161: inst = 32'h38842800;
      88162: inst = 32'h10a00001;
      88163: inst = 32'hca05867;
      88164: inst = 32'h13e00001;
      88165: inst = 32'hfe0d96a;
      88166: inst = 32'h5be00000;
      88167: inst = 32'h8c50000;
      88168: inst = 32'h24612800;
      88169: inst = 32'h10a00000;
      88170: inst = 32'hca00007;
      88171: inst = 32'h24822800;
      88172: inst = 32'h10a00000;
      88173: inst = 32'hca00004;
      88174: inst = 32'h38632800;
      88175: inst = 32'h38842800;
      88176: inst = 32'h10a00001;
      88177: inst = 32'hca05875;
      88178: inst = 32'h13e00001;
      88179: inst = 32'hfe0d96a;
      88180: inst = 32'h5be00000;
      88181: inst = 32'h8c50000;
      88182: inst = 32'h24612800;
      88183: inst = 32'h10a00000;
      88184: inst = 32'hca00007;
      88185: inst = 32'h24822800;
      88186: inst = 32'h10a00000;
      88187: inst = 32'hca00004;
      88188: inst = 32'h38632800;
      88189: inst = 32'h38842800;
      88190: inst = 32'h10a00001;
      88191: inst = 32'hca05883;
      88192: inst = 32'h13e00001;
      88193: inst = 32'hfe0d96a;
      88194: inst = 32'h5be00000;
      88195: inst = 32'h8c50000;
      88196: inst = 32'h24612800;
      88197: inst = 32'h10a00000;
      88198: inst = 32'hca00007;
      88199: inst = 32'h24822800;
      88200: inst = 32'h10a00000;
      88201: inst = 32'hca00004;
      88202: inst = 32'h38632800;
      88203: inst = 32'h38842800;
      88204: inst = 32'h10a00001;
      88205: inst = 32'hca05891;
      88206: inst = 32'h13e00001;
      88207: inst = 32'hfe0d96a;
      88208: inst = 32'h5be00000;
      88209: inst = 32'h8c50000;
      88210: inst = 32'h24612800;
      88211: inst = 32'h10a00000;
      88212: inst = 32'hca00007;
      88213: inst = 32'h24822800;
      88214: inst = 32'h10a00000;
      88215: inst = 32'hca00004;
      88216: inst = 32'h38632800;
      88217: inst = 32'h38842800;
      88218: inst = 32'h10a00001;
      88219: inst = 32'hca0589f;
      88220: inst = 32'h13e00001;
      88221: inst = 32'hfe0d96a;
      88222: inst = 32'h5be00000;
      88223: inst = 32'h8c50000;
      88224: inst = 32'h24612800;
      88225: inst = 32'h10a00000;
      88226: inst = 32'hca00007;
      88227: inst = 32'h24822800;
      88228: inst = 32'h10a00000;
      88229: inst = 32'hca00004;
      88230: inst = 32'h38632800;
      88231: inst = 32'h38842800;
      88232: inst = 32'h10a00001;
      88233: inst = 32'hca058ad;
      88234: inst = 32'h13e00001;
      88235: inst = 32'hfe0d96a;
      88236: inst = 32'h5be00000;
      88237: inst = 32'h8c50000;
      88238: inst = 32'h24612800;
      88239: inst = 32'h10a00000;
      88240: inst = 32'hca00007;
      88241: inst = 32'h24822800;
      88242: inst = 32'h10a00000;
      88243: inst = 32'hca00004;
      88244: inst = 32'h38632800;
      88245: inst = 32'h38842800;
      88246: inst = 32'h10a00001;
      88247: inst = 32'hca058bb;
      88248: inst = 32'h13e00001;
      88249: inst = 32'hfe0d96a;
      88250: inst = 32'h5be00000;
      88251: inst = 32'h8c50000;
      88252: inst = 32'h24612800;
      88253: inst = 32'h10a00000;
      88254: inst = 32'hca00007;
      88255: inst = 32'h24822800;
      88256: inst = 32'h10a00000;
      88257: inst = 32'hca00004;
      88258: inst = 32'h38632800;
      88259: inst = 32'h38842800;
      88260: inst = 32'h10a00001;
      88261: inst = 32'hca058c9;
      88262: inst = 32'h13e00001;
      88263: inst = 32'hfe0d96a;
      88264: inst = 32'h5be00000;
      88265: inst = 32'h8c50000;
      88266: inst = 32'h24612800;
      88267: inst = 32'h10a00000;
      88268: inst = 32'hca00007;
      88269: inst = 32'h24822800;
      88270: inst = 32'h10a00000;
      88271: inst = 32'hca00004;
      88272: inst = 32'h38632800;
      88273: inst = 32'h38842800;
      88274: inst = 32'h10a00001;
      88275: inst = 32'hca058d7;
      88276: inst = 32'h13e00001;
      88277: inst = 32'hfe0d96a;
      88278: inst = 32'h5be00000;
      88279: inst = 32'h8c50000;
      88280: inst = 32'h24612800;
      88281: inst = 32'h10a00000;
      88282: inst = 32'hca00007;
      88283: inst = 32'h24822800;
      88284: inst = 32'h10a00000;
      88285: inst = 32'hca00004;
      88286: inst = 32'h38632800;
      88287: inst = 32'h38842800;
      88288: inst = 32'h10a00001;
      88289: inst = 32'hca058e5;
      88290: inst = 32'h13e00001;
      88291: inst = 32'hfe0d96a;
      88292: inst = 32'h5be00000;
      88293: inst = 32'h8c50000;
      88294: inst = 32'h24612800;
      88295: inst = 32'h10a00000;
      88296: inst = 32'hca00007;
      88297: inst = 32'h24822800;
      88298: inst = 32'h10a00000;
      88299: inst = 32'hca00004;
      88300: inst = 32'h38632800;
      88301: inst = 32'h38842800;
      88302: inst = 32'h10a00001;
      88303: inst = 32'hca058f3;
      88304: inst = 32'h13e00001;
      88305: inst = 32'hfe0d96a;
      88306: inst = 32'h5be00000;
      88307: inst = 32'h8c50000;
      88308: inst = 32'h24612800;
      88309: inst = 32'h10a00000;
      88310: inst = 32'hca00007;
      88311: inst = 32'h24822800;
      88312: inst = 32'h10a00000;
      88313: inst = 32'hca00004;
      88314: inst = 32'h38632800;
      88315: inst = 32'h38842800;
      88316: inst = 32'h10a00001;
      88317: inst = 32'hca05901;
      88318: inst = 32'h13e00001;
      88319: inst = 32'hfe0d96a;
      88320: inst = 32'h5be00000;
      88321: inst = 32'h8c50000;
      88322: inst = 32'h24612800;
      88323: inst = 32'h10a00000;
      88324: inst = 32'hca00007;
      88325: inst = 32'h24822800;
      88326: inst = 32'h10a00000;
      88327: inst = 32'hca00004;
      88328: inst = 32'h38632800;
      88329: inst = 32'h38842800;
      88330: inst = 32'h10a00001;
      88331: inst = 32'hca0590f;
      88332: inst = 32'h13e00001;
      88333: inst = 32'hfe0d96a;
      88334: inst = 32'h5be00000;
      88335: inst = 32'h8c50000;
      88336: inst = 32'h24612800;
      88337: inst = 32'h10a00000;
      88338: inst = 32'hca00007;
      88339: inst = 32'h24822800;
      88340: inst = 32'h10a00000;
      88341: inst = 32'hca00004;
      88342: inst = 32'h38632800;
      88343: inst = 32'h38842800;
      88344: inst = 32'h10a00001;
      88345: inst = 32'hca0591d;
      88346: inst = 32'h13e00001;
      88347: inst = 32'hfe0d96a;
      88348: inst = 32'h5be00000;
      88349: inst = 32'h8c50000;
      88350: inst = 32'h24612800;
      88351: inst = 32'h10a00000;
      88352: inst = 32'hca00007;
      88353: inst = 32'h24822800;
      88354: inst = 32'h10a00000;
      88355: inst = 32'hca00004;
      88356: inst = 32'h38632800;
      88357: inst = 32'h38842800;
      88358: inst = 32'h10a00001;
      88359: inst = 32'hca0592b;
      88360: inst = 32'h13e00001;
      88361: inst = 32'hfe0d96a;
      88362: inst = 32'h5be00000;
      88363: inst = 32'h8c50000;
      88364: inst = 32'h24612800;
      88365: inst = 32'h10a00000;
      88366: inst = 32'hca00007;
      88367: inst = 32'h24822800;
      88368: inst = 32'h10a00000;
      88369: inst = 32'hca00004;
      88370: inst = 32'h38632800;
      88371: inst = 32'h38842800;
      88372: inst = 32'h10a00001;
      88373: inst = 32'hca05939;
      88374: inst = 32'h13e00001;
      88375: inst = 32'hfe0d96a;
      88376: inst = 32'h5be00000;
      88377: inst = 32'h8c50000;
      88378: inst = 32'h24612800;
      88379: inst = 32'h10a00000;
      88380: inst = 32'hca00007;
      88381: inst = 32'h24822800;
      88382: inst = 32'h10a00000;
      88383: inst = 32'hca00004;
      88384: inst = 32'h38632800;
      88385: inst = 32'h38842800;
      88386: inst = 32'h10a00001;
      88387: inst = 32'hca05947;
      88388: inst = 32'h13e00001;
      88389: inst = 32'hfe0d96a;
      88390: inst = 32'h5be00000;
      88391: inst = 32'h8c50000;
      88392: inst = 32'h24612800;
      88393: inst = 32'h10a00000;
      88394: inst = 32'hca00007;
      88395: inst = 32'h24822800;
      88396: inst = 32'h10a00000;
      88397: inst = 32'hca00004;
      88398: inst = 32'h38632800;
      88399: inst = 32'h38842800;
      88400: inst = 32'h10a00001;
      88401: inst = 32'hca05955;
      88402: inst = 32'h13e00001;
      88403: inst = 32'hfe0d96a;
      88404: inst = 32'h5be00000;
      88405: inst = 32'h8c50000;
      88406: inst = 32'h24612800;
      88407: inst = 32'h10a00000;
      88408: inst = 32'hca00007;
      88409: inst = 32'h24822800;
      88410: inst = 32'h10a00000;
      88411: inst = 32'hca00004;
      88412: inst = 32'h38632800;
      88413: inst = 32'h38842800;
      88414: inst = 32'h10a00001;
      88415: inst = 32'hca05963;
      88416: inst = 32'h13e00001;
      88417: inst = 32'hfe0d96a;
      88418: inst = 32'h5be00000;
      88419: inst = 32'h8c50000;
      88420: inst = 32'h24612800;
      88421: inst = 32'h10a00000;
      88422: inst = 32'hca00007;
      88423: inst = 32'h24822800;
      88424: inst = 32'h10a00000;
      88425: inst = 32'hca00004;
      88426: inst = 32'h38632800;
      88427: inst = 32'h38842800;
      88428: inst = 32'h10a00001;
      88429: inst = 32'hca05971;
      88430: inst = 32'h13e00001;
      88431: inst = 32'hfe0d96a;
      88432: inst = 32'h5be00000;
      88433: inst = 32'h8c50000;
      88434: inst = 32'h24612800;
      88435: inst = 32'h10a00000;
      88436: inst = 32'hca00007;
      88437: inst = 32'h24822800;
      88438: inst = 32'h10a00000;
      88439: inst = 32'hca00004;
      88440: inst = 32'h38632800;
      88441: inst = 32'h38842800;
      88442: inst = 32'h10a00001;
      88443: inst = 32'hca0597f;
      88444: inst = 32'h13e00001;
      88445: inst = 32'hfe0d96a;
      88446: inst = 32'h5be00000;
      88447: inst = 32'h8c50000;
      88448: inst = 32'h24612800;
      88449: inst = 32'h10a00000;
      88450: inst = 32'hca00007;
      88451: inst = 32'h24822800;
      88452: inst = 32'h10a00000;
      88453: inst = 32'hca00004;
      88454: inst = 32'h38632800;
      88455: inst = 32'h38842800;
      88456: inst = 32'h10a00001;
      88457: inst = 32'hca0598d;
      88458: inst = 32'h13e00001;
      88459: inst = 32'hfe0d96a;
      88460: inst = 32'h5be00000;
      88461: inst = 32'h8c50000;
      88462: inst = 32'h24612800;
      88463: inst = 32'h10a00000;
      88464: inst = 32'hca00007;
      88465: inst = 32'h24822800;
      88466: inst = 32'h10a00000;
      88467: inst = 32'hca00004;
      88468: inst = 32'h38632800;
      88469: inst = 32'h38842800;
      88470: inst = 32'h10a00001;
      88471: inst = 32'hca0599b;
      88472: inst = 32'h13e00001;
      88473: inst = 32'hfe0d96a;
      88474: inst = 32'h5be00000;
      88475: inst = 32'h8c50000;
      88476: inst = 32'h24612800;
      88477: inst = 32'h10a00000;
      88478: inst = 32'hca00007;
      88479: inst = 32'h24822800;
      88480: inst = 32'h10a00000;
      88481: inst = 32'hca00004;
      88482: inst = 32'h38632800;
      88483: inst = 32'h38842800;
      88484: inst = 32'h10a00001;
      88485: inst = 32'hca059a9;
      88486: inst = 32'h13e00001;
      88487: inst = 32'hfe0d96a;
      88488: inst = 32'h5be00000;
      88489: inst = 32'h8c50000;
      88490: inst = 32'h24612800;
      88491: inst = 32'h10a00000;
      88492: inst = 32'hca00007;
      88493: inst = 32'h24822800;
      88494: inst = 32'h10a00000;
      88495: inst = 32'hca00004;
      88496: inst = 32'h38632800;
      88497: inst = 32'h38842800;
      88498: inst = 32'h10a00001;
      88499: inst = 32'hca059b7;
      88500: inst = 32'h13e00001;
      88501: inst = 32'hfe0d96a;
      88502: inst = 32'h5be00000;
      88503: inst = 32'h8c50000;
      88504: inst = 32'h24612800;
      88505: inst = 32'h10a00000;
      88506: inst = 32'hca00007;
      88507: inst = 32'h24822800;
      88508: inst = 32'h10a00000;
      88509: inst = 32'hca00004;
      88510: inst = 32'h38632800;
      88511: inst = 32'h38842800;
      88512: inst = 32'h10a00001;
      88513: inst = 32'hca059c5;
      88514: inst = 32'h13e00001;
      88515: inst = 32'hfe0d96a;
      88516: inst = 32'h5be00000;
      88517: inst = 32'h8c50000;
      88518: inst = 32'h24612800;
      88519: inst = 32'h10a00000;
      88520: inst = 32'hca00007;
      88521: inst = 32'h24822800;
      88522: inst = 32'h10a00000;
      88523: inst = 32'hca00004;
      88524: inst = 32'h38632800;
      88525: inst = 32'h38842800;
      88526: inst = 32'h10a00001;
      88527: inst = 32'hca059d3;
      88528: inst = 32'h13e00001;
      88529: inst = 32'hfe0d96a;
      88530: inst = 32'h5be00000;
      88531: inst = 32'h8c50000;
      88532: inst = 32'h24612800;
      88533: inst = 32'h10a00000;
      88534: inst = 32'hca00007;
      88535: inst = 32'h24822800;
      88536: inst = 32'h10a00000;
      88537: inst = 32'hca00004;
      88538: inst = 32'h38632800;
      88539: inst = 32'h38842800;
      88540: inst = 32'h10a00001;
      88541: inst = 32'hca059e1;
      88542: inst = 32'h13e00001;
      88543: inst = 32'hfe0d96a;
      88544: inst = 32'h5be00000;
      88545: inst = 32'h8c50000;
      88546: inst = 32'h24612800;
      88547: inst = 32'h10a00000;
      88548: inst = 32'hca00007;
      88549: inst = 32'h24822800;
      88550: inst = 32'h10a00000;
      88551: inst = 32'hca00004;
      88552: inst = 32'h38632800;
      88553: inst = 32'h38842800;
      88554: inst = 32'h10a00001;
      88555: inst = 32'hca059ef;
      88556: inst = 32'h13e00001;
      88557: inst = 32'hfe0d96a;
      88558: inst = 32'h5be00000;
      88559: inst = 32'h8c50000;
      88560: inst = 32'h24612800;
      88561: inst = 32'h10a00000;
      88562: inst = 32'hca00007;
      88563: inst = 32'h24822800;
      88564: inst = 32'h10a00000;
      88565: inst = 32'hca00004;
      88566: inst = 32'h38632800;
      88567: inst = 32'h38842800;
      88568: inst = 32'h10a00001;
      88569: inst = 32'hca059fd;
      88570: inst = 32'h13e00001;
      88571: inst = 32'hfe0d96a;
      88572: inst = 32'h5be00000;
      88573: inst = 32'h8c50000;
      88574: inst = 32'h24612800;
      88575: inst = 32'h10a00000;
      88576: inst = 32'hca00007;
      88577: inst = 32'h24822800;
      88578: inst = 32'h10a00000;
      88579: inst = 32'hca00004;
      88580: inst = 32'h38632800;
      88581: inst = 32'h38842800;
      88582: inst = 32'h10a00001;
      88583: inst = 32'hca05a0b;
      88584: inst = 32'h13e00001;
      88585: inst = 32'hfe0d96a;
      88586: inst = 32'h5be00000;
      88587: inst = 32'h8c50000;
      88588: inst = 32'h24612800;
      88589: inst = 32'h10a00000;
      88590: inst = 32'hca00007;
      88591: inst = 32'h24822800;
      88592: inst = 32'h10a00000;
      88593: inst = 32'hca00004;
      88594: inst = 32'h38632800;
      88595: inst = 32'h38842800;
      88596: inst = 32'h10a00001;
      88597: inst = 32'hca05a19;
      88598: inst = 32'h13e00001;
      88599: inst = 32'hfe0d96a;
      88600: inst = 32'h5be00000;
      88601: inst = 32'h8c50000;
      88602: inst = 32'h24612800;
      88603: inst = 32'h10a00000;
      88604: inst = 32'hca00007;
      88605: inst = 32'h24822800;
      88606: inst = 32'h10a00000;
      88607: inst = 32'hca00004;
      88608: inst = 32'h38632800;
      88609: inst = 32'h38842800;
      88610: inst = 32'h10a00001;
      88611: inst = 32'hca05a27;
      88612: inst = 32'h13e00001;
      88613: inst = 32'hfe0d96a;
      88614: inst = 32'h5be00000;
      88615: inst = 32'h8c50000;
      88616: inst = 32'h24612800;
      88617: inst = 32'h10a00000;
      88618: inst = 32'hca00007;
      88619: inst = 32'h24822800;
      88620: inst = 32'h10a00000;
      88621: inst = 32'hca00004;
      88622: inst = 32'h38632800;
      88623: inst = 32'h38842800;
      88624: inst = 32'h10a00001;
      88625: inst = 32'hca05a35;
      88626: inst = 32'h13e00001;
      88627: inst = 32'hfe0d96a;
      88628: inst = 32'h5be00000;
      88629: inst = 32'h8c50000;
      88630: inst = 32'h24612800;
      88631: inst = 32'h10a00000;
      88632: inst = 32'hca00007;
      88633: inst = 32'h24822800;
      88634: inst = 32'h10a00000;
      88635: inst = 32'hca00004;
      88636: inst = 32'h38632800;
      88637: inst = 32'h38842800;
      88638: inst = 32'h10a00001;
      88639: inst = 32'hca05a43;
      88640: inst = 32'h13e00001;
      88641: inst = 32'hfe0d96a;
      88642: inst = 32'h5be00000;
      88643: inst = 32'h8c50000;
      88644: inst = 32'h24612800;
      88645: inst = 32'h10a00000;
      88646: inst = 32'hca00007;
      88647: inst = 32'h24822800;
      88648: inst = 32'h10a00000;
      88649: inst = 32'hca00004;
      88650: inst = 32'h38632800;
      88651: inst = 32'h38842800;
      88652: inst = 32'h10a00001;
      88653: inst = 32'hca05a51;
      88654: inst = 32'h13e00001;
      88655: inst = 32'hfe0d96a;
      88656: inst = 32'h5be00000;
      88657: inst = 32'h8c50000;
      88658: inst = 32'h24612800;
      88659: inst = 32'h10a00000;
      88660: inst = 32'hca00007;
      88661: inst = 32'h24822800;
      88662: inst = 32'h10a00000;
      88663: inst = 32'hca00004;
      88664: inst = 32'h38632800;
      88665: inst = 32'h38842800;
      88666: inst = 32'h10a00001;
      88667: inst = 32'hca05a5f;
      88668: inst = 32'h13e00001;
      88669: inst = 32'hfe0d96a;
      88670: inst = 32'h5be00000;
      88671: inst = 32'h8c50000;
      88672: inst = 32'h24612800;
      88673: inst = 32'h10a00000;
      88674: inst = 32'hca00007;
      88675: inst = 32'h24822800;
      88676: inst = 32'h10a00000;
      88677: inst = 32'hca00004;
      88678: inst = 32'h38632800;
      88679: inst = 32'h38842800;
      88680: inst = 32'h10a00001;
      88681: inst = 32'hca05a6d;
      88682: inst = 32'h13e00001;
      88683: inst = 32'hfe0d96a;
      88684: inst = 32'h5be00000;
      88685: inst = 32'h8c50000;
      88686: inst = 32'h24612800;
      88687: inst = 32'h10a00000;
      88688: inst = 32'hca00007;
      88689: inst = 32'h24822800;
      88690: inst = 32'h10a00000;
      88691: inst = 32'hca00004;
      88692: inst = 32'h38632800;
      88693: inst = 32'h38842800;
      88694: inst = 32'h10a00001;
      88695: inst = 32'hca05a7b;
      88696: inst = 32'h13e00001;
      88697: inst = 32'hfe0d96a;
      88698: inst = 32'h5be00000;
      88699: inst = 32'h8c50000;
      88700: inst = 32'h24612800;
      88701: inst = 32'h10a00000;
      88702: inst = 32'hca00007;
      88703: inst = 32'h24822800;
      88704: inst = 32'h10a00000;
      88705: inst = 32'hca00004;
      88706: inst = 32'h38632800;
      88707: inst = 32'h38842800;
      88708: inst = 32'h10a00001;
      88709: inst = 32'hca05a89;
      88710: inst = 32'h13e00001;
      88711: inst = 32'hfe0d96a;
      88712: inst = 32'h5be00000;
      88713: inst = 32'h8c50000;
      88714: inst = 32'h24612800;
      88715: inst = 32'h10a00000;
      88716: inst = 32'hca00007;
      88717: inst = 32'h24822800;
      88718: inst = 32'h10a00000;
      88719: inst = 32'hca00004;
      88720: inst = 32'h38632800;
      88721: inst = 32'h38842800;
      88722: inst = 32'h10a00001;
      88723: inst = 32'hca05a97;
      88724: inst = 32'h13e00001;
      88725: inst = 32'hfe0d96a;
      88726: inst = 32'h5be00000;
      88727: inst = 32'h8c50000;
      88728: inst = 32'h24612800;
      88729: inst = 32'h10a00000;
      88730: inst = 32'hca00007;
      88731: inst = 32'h24822800;
      88732: inst = 32'h10a00000;
      88733: inst = 32'hca00004;
      88734: inst = 32'h38632800;
      88735: inst = 32'h38842800;
      88736: inst = 32'h10a00001;
      88737: inst = 32'hca05aa5;
      88738: inst = 32'h13e00001;
      88739: inst = 32'hfe0d96a;
      88740: inst = 32'h5be00000;
      88741: inst = 32'h8c50000;
      88742: inst = 32'h24612800;
      88743: inst = 32'h10a00000;
      88744: inst = 32'hca00007;
      88745: inst = 32'h24822800;
      88746: inst = 32'h10a00000;
      88747: inst = 32'hca00004;
      88748: inst = 32'h38632800;
      88749: inst = 32'h38842800;
      88750: inst = 32'h10a00001;
      88751: inst = 32'hca05ab3;
      88752: inst = 32'h13e00001;
      88753: inst = 32'hfe0d96a;
      88754: inst = 32'h5be00000;
      88755: inst = 32'h8c50000;
      88756: inst = 32'h24612800;
      88757: inst = 32'h10a00000;
      88758: inst = 32'hca00007;
      88759: inst = 32'h24822800;
      88760: inst = 32'h10a00000;
      88761: inst = 32'hca00004;
      88762: inst = 32'h38632800;
      88763: inst = 32'h38842800;
      88764: inst = 32'h10a00001;
      88765: inst = 32'hca05ac1;
      88766: inst = 32'h13e00001;
      88767: inst = 32'hfe0d96a;
      88768: inst = 32'h5be00000;
      88769: inst = 32'h8c50000;
      88770: inst = 32'h24612800;
      88771: inst = 32'h10a00000;
      88772: inst = 32'hca00007;
      88773: inst = 32'h24822800;
      88774: inst = 32'h10a00000;
      88775: inst = 32'hca00004;
      88776: inst = 32'h38632800;
      88777: inst = 32'h38842800;
      88778: inst = 32'h10a00001;
      88779: inst = 32'hca05acf;
      88780: inst = 32'h13e00001;
      88781: inst = 32'hfe0d96a;
      88782: inst = 32'h5be00000;
      88783: inst = 32'h8c50000;
      88784: inst = 32'h24612800;
      88785: inst = 32'h10a00000;
      88786: inst = 32'hca00007;
      88787: inst = 32'h24822800;
      88788: inst = 32'h10a00000;
      88789: inst = 32'hca00004;
      88790: inst = 32'h38632800;
      88791: inst = 32'h38842800;
      88792: inst = 32'h10a00001;
      88793: inst = 32'hca05add;
      88794: inst = 32'h13e00001;
      88795: inst = 32'hfe0d96a;
      88796: inst = 32'h5be00000;
      88797: inst = 32'h8c50000;
      88798: inst = 32'h24612800;
      88799: inst = 32'h10a00000;
      88800: inst = 32'hca00007;
      88801: inst = 32'h24822800;
      88802: inst = 32'h10a00000;
      88803: inst = 32'hca00004;
      88804: inst = 32'h38632800;
      88805: inst = 32'h38842800;
      88806: inst = 32'h10a00001;
      88807: inst = 32'hca05aeb;
      88808: inst = 32'h13e00001;
      88809: inst = 32'hfe0d96a;
      88810: inst = 32'h5be00000;
      88811: inst = 32'h8c50000;
      88812: inst = 32'h24612800;
      88813: inst = 32'h10a00000;
      88814: inst = 32'hca00007;
      88815: inst = 32'h24822800;
      88816: inst = 32'h10a00000;
      88817: inst = 32'hca00004;
      88818: inst = 32'h38632800;
      88819: inst = 32'h38842800;
      88820: inst = 32'h10a00001;
      88821: inst = 32'hca05af9;
      88822: inst = 32'h13e00001;
      88823: inst = 32'hfe0d96a;
      88824: inst = 32'h5be00000;
      88825: inst = 32'h8c50000;
      88826: inst = 32'h24612800;
      88827: inst = 32'h10a00000;
      88828: inst = 32'hca00007;
      88829: inst = 32'h24822800;
      88830: inst = 32'h10a00000;
      88831: inst = 32'hca00004;
      88832: inst = 32'h38632800;
      88833: inst = 32'h38842800;
      88834: inst = 32'h10a00001;
      88835: inst = 32'hca05b07;
      88836: inst = 32'h13e00001;
      88837: inst = 32'hfe0d96a;
      88838: inst = 32'h5be00000;
      88839: inst = 32'h8c50000;
      88840: inst = 32'h24612800;
      88841: inst = 32'h10a00000;
      88842: inst = 32'hca00007;
      88843: inst = 32'h24822800;
      88844: inst = 32'h10a00000;
      88845: inst = 32'hca00004;
      88846: inst = 32'h38632800;
      88847: inst = 32'h38842800;
      88848: inst = 32'h10a00001;
      88849: inst = 32'hca05b15;
      88850: inst = 32'h13e00001;
      88851: inst = 32'hfe0d96a;
      88852: inst = 32'h5be00000;
      88853: inst = 32'h8c50000;
      88854: inst = 32'h24612800;
      88855: inst = 32'h10a00000;
      88856: inst = 32'hca00007;
      88857: inst = 32'h24822800;
      88858: inst = 32'h10a00000;
      88859: inst = 32'hca00004;
      88860: inst = 32'h38632800;
      88861: inst = 32'h38842800;
      88862: inst = 32'h10a00001;
      88863: inst = 32'hca05b23;
      88864: inst = 32'h13e00001;
      88865: inst = 32'hfe0d96a;
      88866: inst = 32'h5be00000;
      88867: inst = 32'h8c50000;
      88868: inst = 32'h24612800;
      88869: inst = 32'h10a00000;
      88870: inst = 32'hca00007;
      88871: inst = 32'h24822800;
      88872: inst = 32'h10a00000;
      88873: inst = 32'hca00004;
      88874: inst = 32'h38632800;
      88875: inst = 32'h38842800;
      88876: inst = 32'h10a00001;
      88877: inst = 32'hca05b31;
      88878: inst = 32'h13e00001;
      88879: inst = 32'hfe0d96a;
      88880: inst = 32'h5be00000;
      88881: inst = 32'h8c50000;
      88882: inst = 32'h24612800;
      88883: inst = 32'h10a00000;
      88884: inst = 32'hca00007;
      88885: inst = 32'h24822800;
      88886: inst = 32'h10a00000;
      88887: inst = 32'hca00004;
      88888: inst = 32'h38632800;
      88889: inst = 32'h38842800;
      88890: inst = 32'h10a00001;
      88891: inst = 32'hca05b3f;
      88892: inst = 32'h13e00001;
      88893: inst = 32'hfe0d96a;
      88894: inst = 32'h5be00000;
      88895: inst = 32'h8c50000;
      88896: inst = 32'h24612800;
      88897: inst = 32'h10a00000;
      88898: inst = 32'hca00007;
      88899: inst = 32'h24822800;
      88900: inst = 32'h10a00000;
      88901: inst = 32'hca00004;
      88902: inst = 32'h38632800;
      88903: inst = 32'h38842800;
      88904: inst = 32'h10a00001;
      88905: inst = 32'hca05b4d;
      88906: inst = 32'h13e00001;
      88907: inst = 32'hfe0d96a;
      88908: inst = 32'h5be00000;
      88909: inst = 32'h8c50000;
      88910: inst = 32'h24612800;
      88911: inst = 32'h10a00000;
      88912: inst = 32'hca00007;
      88913: inst = 32'h24822800;
      88914: inst = 32'h10a00000;
      88915: inst = 32'hca00004;
      88916: inst = 32'h38632800;
      88917: inst = 32'h38842800;
      88918: inst = 32'h10a00001;
      88919: inst = 32'hca05b5b;
      88920: inst = 32'h13e00001;
      88921: inst = 32'hfe0d96a;
      88922: inst = 32'h5be00000;
      88923: inst = 32'h8c50000;
      88924: inst = 32'h24612800;
      88925: inst = 32'h10a00000;
      88926: inst = 32'hca00007;
      88927: inst = 32'h24822800;
      88928: inst = 32'h10a00000;
      88929: inst = 32'hca00004;
      88930: inst = 32'h38632800;
      88931: inst = 32'h38842800;
      88932: inst = 32'h10a00001;
      88933: inst = 32'hca05b69;
      88934: inst = 32'h13e00001;
      88935: inst = 32'hfe0d96a;
      88936: inst = 32'h5be00000;
      88937: inst = 32'h8c50000;
      88938: inst = 32'h24612800;
      88939: inst = 32'h10a00000;
      88940: inst = 32'hca00008;
      88941: inst = 32'h24822800;
      88942: inst = 32'h10a00000;
      88943: inst = 32'hca00004;
      88944: inst = 32'h38632800;
      88945: inst = 32'h38842800;
      88946: inst = 32'h10a00001;
      88947: inst = 32'hca05b77;
      88948: inst = 32'h13e00001;
      88949: inst = 32'hfe0d96a;
      88950: inst = 32'h5be00000;
      88951: inst = 32'h8c50000;
      88952: inst = 32'h24612800;
      88953: inst = 32'h10a00000;
      88954: inst = 32'hca00008;
      88955: inst = 32'h24822800;
      88956: inst = 32'h10a00000;
      88957: inst = 32'hca00004;
      88958: inst = 32'h38632800;
      88959: inst = 32'h38842800;
      88960: inst = 32'h10a00001;
      88961: inst = 32'hca05b85;
      88962: inst = 32'h13e00001;
      88963: inst = 32'hfe0d96a;
      88964: inst = 32'h5be00000;
      88965: inst = 32'h8c50000;
      88966: inst = 32'h24612800;
      88967: inst = 32'h10a00000;
      88968: inst = 32'hca00008;
      88969: inst = 32'h24822800;
      88970: inst = 32'h10a00000;
      88971: inst = 32'hca00004;
      88972: inst = 32'h38632800;
      88973: inst = 32'h38842800;
      88974: inst = 32'h10a00001;
      88975: inst = 32'hca05b93;
      88976: inst = 32'h13e00001;
      88977: inst = 32'hfe0d96a;
      88978: inst = 32'h5be00000;
      88979: inst = 32'h8c50000;
      88980: inst = 32'h24612800;
      88981: inst = 32'h10a00000;
      88982: inst = 32'hca00008;
      88983: inst = 32'h24822800;
      88984: inst = 32'h10a00000;
      88985: inst = 32'hca00004;
      88986: inst = 32'h38632800;
      88987: inst = 32'h38842800;
      88988: inst = 32'h10a00001;
      88989: inst = 32'hca05ba1;
      88990: inst = 32'h13e00001;
      88991: inst = 32'hfe0d96a;
      88992: inst = 32'h5be00000;
      88993: inst = 32'h8c50000;
      88994: inst = 32'h24612800;
      88995: inst = 32'h10a00000;
      88996: inst = 32'hca00008;
      88997: inst = 32'h24822800;
      88998: inst = 32'h10a00000;
      88999: inst = 32'hca00004;
      89000: inst = 32'h38632800;
      89001: inst = 32'h38842800;
      89002: inst = 32'h10a00001;
      89003: inst = 32'hca05baf;
      89004: inst = 32'h13e00001;
      89005: inst = 32'hfe0d96a;
      89006: inst = 32'h5be00000;
      89007: inst = 32'h8c50000;
      89008: inst = 32'h24612800;
      89009: inst = 32'h10a00000;
      89010: inst = 32'hca00008;
      89011: inst = 32'h24822800;
      89012: inst = 32'h10a00000;
      89013: inst = 32'hca00004;
      89014: inst = 32'h38632800;
      89015: inst = 32'h38842800;
      89016: inst = 32'h10a00001;
      89017: inst = 32'hca05bbd;
      89018: inst = 32'h13e00001;
      89019: inst = 32'hfe0d96a;
      89020: inst = 32'h5be00000;
      89021: inst = 32'h8c50000;
      89022: inst = 32'h24612800;
      89023: inst = 32'h10a00000;
      89024: inst = 32'hca00008;
      89025: inst = 32'h24822800;
      89026: inst = 32'h10a00000;
      89027: inst = 32'hca00004;
      89028: inst = 32'h38632800;
      89029: inst = 32'h38842800;
      89030: inst = 32'h10a00001;
      89031: inst = 32'hca05bcb;
      89032: inst = 32'h13e00001;
      89033: inst = 32'hfe0d96a;
      89034: inst = 32'h5be00000;
      89035: inst = 32'h8c50000;
      89036: inst = 32'h24612800;
      89037: inst = 32'h10a00000;
      89038: inst = 32'hca00008;
      89039: inst = 32'h24822800;
      89040: inst = 32'h10a00000;
      89041: inst = 32'hca00004;
      89042: inst = 32'h38632800;
      89043: inst = 32'h38842800;
      89044: inst = 32'h10a00001;
      89045: inst = 32'hca05bd9;
      89046: inst = 32'h13e00001;
      89047: inst = 32'hfe0d96a;
      89048: inst = 32'h5be00000;
      89049: inst = 32'h8c50000;
      89050: inst = 32'h24612800;
      89051: inst = 32'h10a00000;
      89052: inst = 32'hca00008;
      89053: inst = 32'h24822800;
      89054: inst = 32'h10a00000;
      89055: inst = 32'hca00004;
      89056: inst = 32'h38632800;
      89057: inst = 32'h38842800;
      89058: inst = 32'h10a00001;
      89059: inst = 32'hca05be7;
      89060: inst = 32'h13e00001;
      89061: inst = 32'hfe0d96a;
      89062: inst = 32'h5be00000;
      89063: inst = 32'h8c50000;
      89064: inst = 32'h24612800;
      89065: inst = 32'h10a00000;
      89066: inst = 32'hca00008;
      89067: inst = 32'h24822800;
      89068: inst = 32'h10a00000;
      89069: inst = 32'hca00004;
      89070: inst = 32'h38632800;
      89071: inst = 32'h38842800;
      89072: inst = 32'h10a00001;
      89073: inst = 32'hca05bf5;
      89074: inst = 32'h13e00001;
      89075: inst = 32'hfe0d96a;
      89076: inst = 32'h5be00000;
      89077: inst = 32'h8c50000;
      89078: inst = 32'h24612800;
      89079: inst = 32'h10a00000;
      89080: inst = 32'hca00008;
      89081: inst = 32'h24822800;
      89082: inst = 32'h10a00000;
      89083: inst = 32'hca00004;
      89084: inst = 32'h38632800;
      89085: inst = 32'h38842800;
      89086: inst = 32'h10a00001;
      89087: inst = 32'hca05c03;
      89088: inst = 32'h13e00001;
      89089: inst = 32'hfe0d96a;
      89090: inst = 32'h5be00000;
      89091: inst = 32'h8c50000;
      89092: inst = 32'h24612800;
      89093: inst = 32'h10a00000;
      89094: inst = 32'hca00008;
      89095: inst = 32'h24822800;
      89096: inst = 32'h10a00000;
      89097: inst = 32'hca00004;
      89098: inst = 32'h38632800;
      89099: inst = 32'h38842800;
      89100: inst = 32'h10a00001;
      89101: inst = 32'hca05c11;
      89102: inst = 32'h13e00001;
      89103: inst = 32'hfe0d96a;
      89104: inst = 32'h5be00000;
      89105: inst = 32'h8c50000;
      89106: inst = 32'h24612800;
      89107: inst = 32'h10a00000;
      89108: inst = 32'hca00008;
      89109: inst = 32'h24822800;
      89110: inst = 32'h10a00000;
      89111: inst = 32'hca00004;
      89112: inst = 32'h38632800;
      89113: inst = 32'h38842800;
      89114: inst = 32'h10a00001;
      89115: inst = 32'hca05c1f;
      89116: inst = 32'h13e00001;
      89117: inst = 32'hfe0d96a;
      89118: inst = 32'h5be00000;
      89119: inst = 32'h8c50000;
      89120: inst = 32'h24612800;
      89121: inst = 32'h10a00000;
      89122: inst = 32'hca00008;
      89123: inst = 32'h24822800;
      89124: inst = 32'h10a00000;
      89125: inst = 32'hca00004;
      89126: inst = 32'h38632800;
      89127: inst = 32'h38842800;
      89128: inst = 32'h10a00001;
      89129: inst = 32'hca05c2d;
      89130: inst = 32'h13e00001;
      89131: inst = 32'hfe0d96a;
      89132: inst = 32'h5be00000;
      89133: inst = 32'h8c50000;
      89134: inst = 32'h24612800;
      89135: inst = 32'h10a00000;
      89136: inst = 32'hca00008;
      89137: inst = 32'h24822800;
      89138: inst = 32'h10a00000;
      89139: inst = 32'hca00004;
      89140: inst = 32'h38632800;
      89141: inst = 32'h38842800;
      89142: inst = 32'h10a00001;
      89143: inst = 32'hca05c3b;
      89144: inst = 32'h13e00001;
      89145: inst = 32'hfe0d96a;
      89146: inst = 32'h5be00000;
      89147: inst = 32'h8c50000;
      89148: inst = 32'h24612800;
      89149: inst = 32'h10a00000;
      89150: inst = 32'hca00008;
      89151: inst = 32'h24822800;
      89152: inst = 32'h10a00000;
      89153: inst = 32'hca00004;
      89154: inst = 32'h38632800;
      89155: inst = 32'h38842800;
      89156: inst = 32'h10a00001;
      89157: inst = 32'hca05c49;
      89158: inst = 32'h13e00001;
      89159: inst = 32'hfe0d96a;
      89160: inst = 32'h5be00000;
      89161: inst = 32'h8c50000;
      89162: inst = 32'h24612800;
      89163: inst = 32'h10a00000;
      89164: inst = 32'hca00008;
      89165: inst = 32'h24822800;
      89166: inst = 32'h10a00000;
      89167: inst = 32'hca00004;
      89168: inst = 32'h38632800;
      89169: inst = 32'h38842800;
      89170: inst = 32'h10a00001;
      89171: inst = 32'hca05c57;
      89172: inst = 32'h13e00001;
      89173: inst = 32'hfe0d96a;
      89174: inst = 32'h5be00000;
      89175: inst = 32'h8c50000;
      89176: inst = 32'h24612800;
      89177: inst = 32'h10a00000;
      89178: inst = 32'hca00008;
      89179: inst = 32'h24822800;
      89180: inst = 32'h10a00000;
      89181: inst = 32'hca00004;
      89182: inst = 32'h38632800;
      89183: inst = 32'h38842800;
      89184: inst = 32'h10a00001;
      89185: inst = 32'hca05c65;
      89186: inst = 32'h13e00001;
      89187: inst = 32'hfe0d96a;
      89188: inst = 32'h5be00000;
      89189: inst = 32'h8c50000;
      89190: inst = 32'h24612800;
      89191: inst = 32'h10a00000;
      89192: inst = 32'hca00008;
      89193: inst = 32'h24822800;
      89194: inst = 32'h10a00000;
      89195: inst = 32'hca00004;
      89196: inst = 32'h38632800;
      89197: inst = 32'h38842800;
      89198: inst = 32'h10a00001;
      89199: inst = 32'hca05c73;
      89200: inst = 32'h13e00001;
      89201: inst = 32'hfe0d96a;
      89202: inst = 32'h5be00000;
      89203: inst = 32'h8c50000;
      89204: inst = 32'h24612800;
      89205: inst = 32'h10a00000;
      89206: inst = 32'hca00008;
      89207: inst = 32'h24822800;
      89208: inst = 32'h10a00000;
      89209: inst = 32'hca00004;
      89210: inst = 32'h38632800;
      89211: inst = 32'h38842800;
      89212: inst = 32'h10a00001;
      89213: inst = 32'hca05c81;
      89214: inst = 32'h13e00001;
      89215: inst = 32'hfe0d96a;
      89216: inst = 32'h5be00000;
      89217: inst = 32'h8c50000;
      89218: inst = 32'h24612800;
      89219: inst = 32'h10a00000;
      89220: inst = 32'hca00008;
      89221: inst = 32'h24822800;
      89222: inst = 32'h10a00000;
      89223: inst = 32'hca00004;
      89224: inst = 32'h38632800;
      89225: inst = 32'h38842800;
      89226: inst = 32'h10a00001;
      89227: inst = 32'hca05c8f;
      89228: inst = 32'h13e00001;
      89229: inst = 32'hfe0d96a;
      89230: inst = 32'h5be00000;
      89231: inst = 32'h8c50000;
      89232: inst = 32'h24612800;
      89233: inst = 32'h10a00000;
      89234: inst = 32'hca00008;
      89235: inst = 32'h24822800;
      89236: inst = 32'h10a00000;
      89237: inst = 32'hca00004;
      89238: inst = 32'h38632800;
      89239: inst = 32'h38842800;
      89240: inst = 32'h10a00001;
      89241: inst = 32'hca05c9d;
      89242: inst = 32'h13e00001;
      89243: inst = 32'hfe0d96a;
      89244: inst = 32'h5be00000;
      89245: inst = 32'h8c50000;
      89246: inst = 32'h24612800;
      89247: inst = 32'h10a00000;
      89248: inst = 32'hca00008;
      89249: inst = 32'h24822800;
      89250: inst = 32'h10a00000;
      89251: inst = 32'hca00004;
      89252: inst = 32'h38632800;
      89253: inst = 32'h38842800;
      89254: inst = 32'h10a00001;
      89255: inst = 32'hca05cab;
      89256: inst = 32'h13e00001;
      89257: inst = 32'hfe0d96a;
      89258: inst = 32'h5be00000;
      89259: inst = 32'h8c50000;
      89260: inst = 32'h24612800;
      89261: inst = 32'h10a00000;
      89262: inst = 32'hca00008;
      89263: inst = 32'h24822800;
      89264: inst = 32'h10a00000;
      89265: inst = 32'hca00004;
      89266: inst = 32'h38632800;
      89267: inst = 32'h38842800;
      89268: inst = 32'h10a00001;
      89269: inst = 32'hca05cb9;
      89270: inst = 32'h13e00001;
      89271: inst = 32'hfe0d96a;
      89272: inst = 32'h5be00000;
      89273: inst = 32'h8c50000;
      89274: inst = 32'h24612800;
      89275: inst = 32'h10a00000;
      89276: inst = 32'hca00008;
      89277: inst = 32'h24822800;
      89278: inst = 32'h10a00000;
      89279: inst = 32'hca00004;
      89280: inst = 32'h38632800;
      89281: inst = 32'h38842800;
      89282: inst = 32'h10a00001;
      89283: inst = 32'hca05cc7;
      89284: inst = 32'h13e00001;
      89285: inst = 32'hfe0d96a;
      89286: inst = 32'h5be00000;
      89287: inst = 32'h8c50000;
      89288: inst = 32'h24612800;
      89289: inst = 32'h10a00000;
      89290: inst = 32'hca00008;
      89291: inst = 32'h24822800;
      89292: inst = 32'h10a00000;
      89293: inst = 32'hca00004;
      89294: inst = 32'h38632800;
      89295: inst = 32'h38842800;
      89296: inst = 32'h10a00001;
      89297: inst = 32'hca05cd5;
      89298: inst = 32'h13e00001;
      89299: inst = 32'hfe0d96a;
      89300: inst = 32'h5be00000;
      89301: inst = 32'h8c50000;
      89302: inst = 32'h24612800;
      89303: inst = 32'h10a00000;
      89304: inst = 32'hca00008;
      89305: inst = 32'h24822800;
      89306: inst = 32'h10a00000;
      89307: inst = 32'hca00004;
      89308: inst = 32'h38632800;
      89309: inst = 32'h38842800;
      89310: inst = 32'h10a00001;
      89311: inst = 32'hca05ce3;
      89312: inst = 32'h13e00001;
      89313: inst = 32'hfe0d96a;
      89314: inst = 32'h5be00000;
      89315: inst = 32'h8c50000;
      89316: inst = 32'h24612800;
      89317: inst = 32'h10a00000;
      89318: inst = 32'hca00008;
      89319: inst = 32'h24822800;
      89320: inst = 32'h10a00000;
      89321: inst = 32'hca00004;
      89322: inst = 32'h38632800;
      89323: inst = 32'h38842800;
      89324: inst = 32'h10a00001;
      89325: inst = 32'hca05cf1;
      89326: inst = 32'h13e00001;
      89327: inst = 32'hfe0d96a;
      89328: inst = 32'h5be00000;
      89329: inst = 32'h8c50000;
      89330: inst = 32'h24612800;
      89331: inst = 32'h10a00000;
      89332: inst = 32'hca00008;
      89333: inst = 32'h24822800;
      89334: inst = 32'h10a00000;
      89335: inst = 32'hca00004;
      89336: inst = 32'h38632800;
      89337: inst = 32'h38842800;
      89338: inst = 32'h10a00001;
      89339: inst = 32'hca05cff;
      89340: inst = 32'h13e00001;
      89341: inst = 32'hfe0d96a;
      89342: inst = 32'h5be00000;
      89343: inst = 32'h8c50000;
      89344: inst = 32'h24612800;
      89345: inst = 32'h10a00000;
      89346: inst = 32'hca00008;
      89347: inst = 32'h24822800;
      89348: inst = 32'h10a00000;
      89349: inst = 32'hca00004;
      89350: inst = 32'h38632800;
      89351: inst = 32'h38842800;
      89352: inst = 32'h10a00001;
      89353: inst = 32'hca05d0d;
      89354: inst = 32'h13e00001;
      89355: inst = 32'hfe0d96a;
      89356: inst = 32'h5be00000;
      89357: inst = 32'h8c50000;
      89358: inst = 32'h24612800;
      89359: inst = 32'h10a00000;
      89360: inst = 32'hca00008;
      89361: inst = 32'h24822800;
      89362: inst = 32'h10a00000;
      89363: inst = 32'hca00004;
      89364: inst = 32'h38632800;
      89365: inst = 32'h38842800;
      89366: inst = 32'h10a00001;
      89367: inst = 32'hca05d1b;
      89368: inst = 32'h13e00001;
      89369: inst = 32'hfe0d96a;
      89370: inst = 32'h5be00000;
      89371: inst = 32'h8c50000;
      89372: inst = 32'h24612800;
      89373: inst = 32'h10a00000;
      89374: inst = 32'hca00008;
      89375: inst = 32'h24822800;
      89376: inst = 32'h10a00000;
      89377: inst = 32'hca00004;
      89378: inst = 32'h38632800;
      89379: inst = 32'h38842800;
      89380: inst = 32'h10a00001;
      89381: inst = 32'hca05d29;
      89382: inst = 32'h13e00001;
      89383: inst = 32'hfe0d96a;
      89384: inst = 32'h5be00000;
      89385: inst = 32'h8c50000;
      89386: inst = 32'h24612800;
      89387: inst = 32'h10a00000;
      89388: inst = 32'hca00008;
      89389: inst = 32'h24822800;
      89390: inst = 32'h10a00000;
      89391: inst = 32'hca00004;
      89392: inst = 32'h38632800;
      89393: inst = 32'h38842800;
      89394: inst = 32'h10a00001;
      89395: inst = 32'hca05d37;
      89396: inst = 32'h13e00001;
      89397: inst = 32'hfe0d96a;
      89398: inst = 32'h5be00000;
      89399: inst = 32'h8c50000;
      89400: inst = 32'h24612800;
      89401: inst = 32'h10a00000;
      89402: inst = 32'hca00008;
      89403: inst = 32'h24822800;
      89404: inst = 32'h10a00000;
      89405: inst = 32'hca00004;
      89406: inst = 32'h38632800;
      89407: inst = 32'h38842800;
      89408: inst = 32'h10a00001;
      89409: inst = 32'hca05d45;
      89410: inst = 32'h13e00001;
      89411: inst = 32'hfe0d96a;
      89412: inst = 32'h5be00000;
      89413: inst = 32'h8c50000;
      89414: inst = 32'h24612800;
      89415: inst = 32'h10a00000;
      89416: inst = 32'hca00008;
      89417: inst = 32'h24822800;
      89418: inst = 32'h10a00000;
      89419: inst = 32'hca00004;
      89420: inst = 32'h38632800;
      89421: inst = 32'h38842800;
      89422: inst = 32'h10a00001;
      89423: inst = 32'hca05d53;
      89424: inst = 32'h13e00001;
      89425: inst = 32'hfe0d96a;
      89426: inst = 32'h5be00000;
      89427: inst = 32'h8c50000;
      89428: inst = 32'h24612800;
      89429: inst = 32'h10a00000;
      89430: inst = 32'hca00008;
      89431: inst = 32'h24822800;
      89432: inst = 32'h10a00000;
      89433: inst = 32'hca00004;
      89434: inst = 32'h38632800;
      89435: inst = 32'h38842800;
      89436: inst = 32'h10a00001;
      89437: inst = 32'hca05d61;
      89438: inst = 32'h13e00001;
      89439: inst = 32'hfe0d96a;
      89440: inst = 32'h5be00000;
      89441: inst = 32'h8c50000;
      89442: inst = 32'h24612800;
      89443: inst = 32'h10a00000;
      89444: inst = 32'hca00008;
      89445: inst = 32'h24822800;
      89446: inst = 32'h10a00000;
      89447: inst = 32'hca00004;
      89448: inst = 32'h38632800;
      89449: inst = 32'h38842800;
      89450: inst = 32'h10a00001;
      89451: inst = 32'hca05d6f;
      89452: inst = 32'h13e00001;
      89453: inst = 32'hfe0d96a;
      89454: inst = 32'h5be00000;
      89455: inst = 32'h8c50000;
      89456: inst = 32'h24612800;
      89457: inst = 32'h10a00000;
      89458: inst = 32'hca00008;
      89459: inst = 32'h24822800;
      89460: inst = 32'h10a00000;
      89461: inst = 32'hca00004;
      89462: inst = 32'h38632800;
      89463: inst = 32'h38842800;
      89464: inst = 32'h10a00001;
      89465: inst = 32'hca05d7d;
      89466: inst = 32'h13e00001;
      89467: inst = 32'hfe0d96a;
      89468: inst = 32'h5be00000;
      89469: inst = 32'h8c50000;
      89470: inst = 32'h24612800;
      89471: inst = 32'h10a00000;
      89472: inst = 32'hca00008;
      89473: inst = 32'h24822800;
      89474: inst = 32'h10a00000;
      89475: inst = 32'hca00004;
      89476: inst = 32'h38632800;
      89477: inst = 32'h38842800;
      89478: inst = 32'h10a00001;
      89479: inst = 32'hca05d8b;
      89480: inst = 32'h13e00001;
      89481: inst = 32'hfe0d96a;
      89482: inst = 32'h5be00000;
      89483: inst = 32'h8c50000;
      89484: inst = 32'h24612800;
      89485: inst = 32'h10a00000;
      89486: inst = 32'hca00008;
      89487: inst = 32'h24822800;
      89488: inst = 32'h10a00000;
      89489: inst = 32'hca00004;
      89490: inst = 32'h38632800;
      89491: inst = 32'h38842800;
      89492: inst = 32'h10a00001;
      89493: inst = 32'hca05d99;
      89494: inst = 32'h13e00001;
      89495: inst = 32'hfe0d96a;
      89496: inst = 32'h5be00000;
      89497: inst = 32'h8c50000;
      89498: inst = 32'h24612800;
      89499: inst = 32'h10a00000;
      89500: inst = 32'hca00008;
      89501: inst = 32'h24822800;
      89502: inst = 32'h10a00000;
      89503: inst = 32'hca00004;
      89504: inst = 32'h38632800;
      89505: inst = 32'h38842800;
      89506: inst = 32'h10a00001;
      89507: inst = 32'hca05da7;
      89508: inst = 32'h13e00001;
      89509: inst = 32'hfe0d96a;
      89510: inst = 32'h5be00000;
      89511: inst = 32'h8c50000;
      89512: inst = 32'h24612800;
      89513: inst = 32'h10a00000;
      89514: inst = 32'hca00008;
      89515: inst = 32'h24822800;
      89516: inst = 32'h10a00000;
      89517: inst = 32'hca00004;
      89518: inst = 32'h38632800;
      89519: inst = 32'h38842800;
      89520: inst = 32'h10a00001;
      89521: inst = 32'hca05db5;
      89522: inst = 32'h13e00001;
      89523: inst = 32'hfe0d96a;
      89524: inst = 32'h5be00000;
      89525: inst = 32'h8c50000;
      89526: inst = 32'h24612800;
      89527: inst = 32'h10a00000;
      89528: inst = 32'hca00008;
      89529: inst = 32'h24822800;
      89530: inst = 32'h10a00000;
      89531: inst = 32'hca00004;
      89532: inst = 32'h38632800;
      89533: inst = 32'h38842800;
      89534: inst = 32'h10a00001;
      89535: inst = 32'hca05dc3;
      89536: inst = 32'h13e00001;
      89537: inst = 32'hfe0d96a;
      89538: inst = 32'h5be00000;
      89539: inst = 32'h8c50000;
      89540: inst = 32'h24612800;
      89541: inst = 32'h10a00000;
      89542: inst = 32'hca00008;
      89543: inst = 32'h24822800;
      89544: inst = 32'h10a00000;
      89545: inst = 32'hca00004;
      89546: inst = 32'h38632800;
      89547: inst = 32'h38842800;
      89548: inst = 32'h10a00001;
      89549: inst = 32'hca05dd1;
      89550: inst = 32'h13e00001;
      89551: inst = 32'hfe0d96a;
      89552: inst = 32'h5be00000;
      89553: inst = 32'h8c50000;
      89554: inst = 32'h24612800;
      89555: inst = 32'h10a00000;
      89556: inst = 32'hca00008;
      89557: inst = 32'h24822800;
      89558: inst = 32'h10a00000;
      89559: inst = 32'hca00004;
      89560: inst = 32'h38632800;
      89561: inst = 32'h38842800;
      89562: inst = 32'h10a00001;
      89563: inst = 32'hca05ddf;
      89564: inst = 32'h13e00001;
      89565: inst = 32'hfe0d96a;
      89566: inst = 32'h5be00000;
      89567: inst = 32'h8c50000;
      89568: inst = 32'h24612800;
      89569: inst = 32'h10a00000;
      89570: inst = 32'hca00008;
      89571: inst = 32'h24822800;
      89572: inst = 32'h10a00000;
      89573: inst = 32'hca00004;
      89574: inst = 32'h38632800;
      89575: inst = 32'h38842800;
      89576: inst = 32'h10a00001;
      89577: inst = 32'hca05ded;
      89578: inst = 32'h13e00001;
      89579: inst = 32'hfe0d96a;
      89580: inst = 32'h5be00000;
      89581: inst = 32'h8c50000;
      89582: inst = 32'h24612800;
      89583: inst = 32'h10a00000;
      89584: inst = 32'hca00008;
      89585: inst = 32'h24822800;
      89586: inst = 32'h10a00000;
      89587: inst = 32'hca00004;
      89588: inst = 32'h38632800;
      89589: inst = 32'h38842800;
      89590: inst = 32'h10a00001;
      89591: inst = 32'hca05dfb;
      89592: inst = 32'h13e00001;
      89593: inst = 32'hfe0d96a;
      89594: inst = 32'h5be00000;
      89595: inst = 32'h8c50000;
      89596: inst = 32'h24612800;
      89597: inst = 32'h10a00000;
      89598: inst = 32'hca00008;
      89599: inst = 32'h24822800;
      89600: inst = 32'h10a00000;
      89601: inst = 32'hca00004;
      89602: inst = 32'h38632800;
      89603: inst = 32'h38842800;
      89604: inst = 32'h10a00001;
      89605: inst = 32'hca05e09;
      89606: inst = 32'h13e00001;
      89607: inst = 32'hfe0d96a;
      89608: inst = 32'h5be00000;
      89609: inst = 32'h8c50000;
      89610: inst = 32'h24612800;
      89611: inst = 32'h10a00000;
      89612: inst = 32'hca00008;
      89613: inst = 32'h24822800;
      89614: inst = 32'h10a00000;
      89615: inst = 32'hca00004;
      89616: inst = 32'h38632800;
      89617: inst = 32'h38842800;
      89618: inst = 32'h10a00001;
      89619: inst = 32'hca05e17;
      89620: inst = 32'h13e00001;
      89621: inst = 32'hfe0d96a;
      89622: inst = 32'h5be00000;
      89623: inst = 32'h8c50000;
      89624: inst = 32'h24612800;
      89625: inst = 32'h10a00000;
      89626: inst = 32'hca00008;
      89627: inst = 32'h24822800;
      89628: inst = 32'h10a00000;
      89629: inst = 32'hca00004;
      89630: inst = 32'h38632800;
      89631: inst = 32'h38842800;
      89632: inst = 32'h10a00001;
      89633: inst = 32'hca05e25;
      89634: inst = 32'h13e00001;
      89635: inst = 32'hfe0d96a;
      89636: inst = 32'h5be00000;
      89637: inst = 32'h8c50000;
      89638: inst = 32'h24612800;
      89639: inst = 32'h10a00000;
      89640: inst = 32'hca00008;
      89641: inst = 32'h24822800;
      89642: inst = 32'h10a00000;
      89643: inst = 32'hca00004;
      89644: inst = 32'h38632800;
      89645: inst = 32'h38842800;
      89646: inst = 32'h10a00001;
      89647: inst = 32'hca05e33;
      89648: inst = 32'h13e00001;
      89649: inst = 32'hfe0d96a;
      89650: inst = 32'h5be00000;
      89651: inst = 32'h8c50000;
      89652: inst = 32'h24612800;
      89653: inst = 32'h10a00000;
      89654: inst = 32'hca00008;
      89655: inst = 32'h24822800;
      89656: inst = 32'h10a00000;
      89657: inst = 32'hca00004;
      89658: inst = 32'h38632800;
      89659: inst = 32'h38842800;
      89660: inst = 32'h10a00001;
      89661: inst = 32'hca05e41;
      89662: inst = 32'h13e00001;
      89663: inst = 32'hfe0d96a;
      89664: inst = 32'h5be00000;
      89665: inst = 32'h8c50000;
      89666: inst = 32'h24612800;
      89667: inst = 32'h10a00000;
      89668: inst = 32'hca00008;
      89669: inst = 32'h24822800;
      89670: inst = 32'h10a00000;
      89671: inst = 32'hca00004;
      89672: inst = 32'h38632800;
      89673: inst = 32'h38842800;
      89674: inst = 32'h10a00001;
      89675: inst = 32'hca05e4f;
      89676: inst = 32'h13e00001;
      89677: inst = 32'hfe0d96a;
      89678: inst = 32'h5be00000;
      89679: inst = 32'h8c50000;
      89680: inst = 32'h24612800;
      89681: inst = 32'h10a00000;
      89682: inst = 32'hca00008;
      89683: inst = 32'h24822800;
      89684: inst = 32'h10a00000;
      89685: inst = 32'hca00004;
      89686: inst = 32'h38632800;
      89687: inst = 32'h38842800;
      89688: inst = 32'h10a00001;
      89689: inst = 32'hca05e5d;
      89690: inst = 32'h13e00001;
      89691: inst = 32'hfe0d96a;
      89692: inst = 32'h5be00000;
      89693: inst = 32'h8c50000;
      89694: inst = 32'h24612800;
      89695: inst = 32'h10a00000;
      89696: inst = 32'hca00008;
      89697: inst = 32'h24822800;
      89698: inst = 32'h10a00000;
      89699: inst = 32'hca00004;
      89700: inst = 32'h38632800;
      89701: inst = 32'h38842800;
      89702: inst = 32'h10a00001;
      89703: inst = 32'hca05e6b;
      89704: inst = 32'h13e00001;
      89705: inst = 32'hfe0d96a;
      89706: inst = 32'h5be00000;
      89707: inst = 32'h8c50000;
      89708: inst = 32'h24612800;
      89709: inst = 32'h10a00000;
      89710: inst = 32'hca00008;
      89711: inst = 32'h24822800;
      89712: inst = 32'h10a00000;
      89713: inst = 32'hca00004;
      89714: inst = 32'h38632800;
      89715: inst = 32'h38842800;
      89716: inst = 32'h10a00001;
      89717: inst = 32'hca05e79;
      89718: inst = 32'h13e00001;
      89719: inst = 32'hfe0d96a;
      89720: inst = 32'h5be00000;
      89721: inst = 32'h8c50000;
      89722: inst = 32'h24612800;
      89723: inst = 32'h10a00000;
      89724: inst = 32'hca00008;
      89725: inst = 32'h24822800;
      89726: inst = 32'h10a00000;
      89727: inst = 32'hca00004;
      89728: inst = 32'h38632800;
      89729: inst = 32'h38842800;
      89730: inst = 32'h10a00001;
      89731: inst = 32'hca05e87;
      89732: inst = 32'h13e00001;
      89733: inst = 32'hfe0d96a;
      89734: inst = 32'h5be00000;
      89735: inst = 32'h8c50000;
      89736: inst = 32'h24612800;
      89737: inst = 32'h10a00000;
      89738: inst = 32'hca00008;
      89739: inst = 32'h24822800;
      89740: inst = 32'h10a00000;
      89741: inst = 32'hca00004;
      89742: inst = 32'h38632800;
      89743: inst = 32'h38842800;
      89744: inst = 32'h10a00001;
      89745: inst = 32'hca05e95;
      89746: inst = 32'h13e00001;
      89747: inst = 32'hfe0d96a;
      89748: inst = 32'h5be00000;
      89749: inst = 32'h8c50000;
      89750: inst = 32'h24612800;
      89751: inst = 32'h10a00000;
      89752: inst = 32'hca00008;
      89753: inst = 32'h24822800;
      89754: inst = 32'h10a00000;
      89755: inst = 32'hca00004;
      89756: inst = 32'h38632800;
      89757: inst = 32'h38842800;
      89758: inst = 32'h10a00001;
      89759: inst = 32'hca05ea3;
      89760: inst = 32'h13e00001;
      89761: inst = 32'hfe0d96a;
      89762: inst = 32'h5be00000;
      89763: inst = 32'h8c50000;
      89764: inst = 32'h24612800;
      89765: inst = 32'h10a00000;
      89766: inst = 32'hca00008;
      89767: inst = 32'h24822800;
      89768: inst = 32'h10a00000;
      89769: inst = 32'hca00004;
      89770: inst = 32'h38632800;
      89771: inst = 32'h38842800;
      89772: inst = 32'h10a00001;
      89773: inst = 32'hca05eb1;
      89774: inst = 32'h13e00001;
      89775: inst = 32'hfe0d96a;
      89776: inst = 32'h5be00000;
      89777: inst = 32'h8c50000;
      89778: inst = 32'h24612800;
      89779: inst = 32'h10a00000;
      89780: inst = 32'hca00008;
      89781: inst = 32'h24822800;
      89782: inst = 32'h10a00000;
      89783: inst = 32'hca00004;
      89784: inst = 32'h38632800;
      89785: inst = 32'h38842800;
      89786: inst = 32'h10a00001;
      89787: inst = 32'hca05ebf;
      89788: inst = 32'h13e00001;
      89789: inst = 32'hfe0d96a;
      89790: inst = 32'h5be00000;
      89791: inst = 32'h8c50000;
      89792: inst = 32'h24612800;
      89793: inst = 32'h10a00000;
      89794: inst = 32'hca00008;
      89795: inst = 32'h24822800;
      89796: inst = 32'h10a00000;
      89797: inst = 32'hca00004;
      89798: inst = 32'h38632800;
      89799: inst = 32'h38842800;
      89800: inst = 32'h10a00001;
      89801: inst = 32'hca05ecd;
      89802: inst = 32'h13e00001;
      89803: inst = 32'hfe0d96a;
      89804: inst = 32'h5be00000;
      89805: inst = 32'h8c50000;
      89806: inst = 32'h24612800;
      89807: inst = 32'h10a00000;
      89808: inst = 32'hca00008;
      89809: inst = 32'h24822800;
      89810: inst = 32'h10a00000;
      89811: inst = 32'hca00004;
      89812: inst = 32'h38632800;
      89813: inst = 32'h38842800;
      89814: inst = 32'h10a00001;
      89815: inst = 32'hca05edb;
      89816: inst = 32'h13e00001;
      89817: inst = 32'hfe0d96a;
      89818: inst = 32'h5be00000;
      89819: inst = 32'h8c50000;
      89820: inst = 32'h24612800;
      89821: inst = 32'h10a00000;
      89822: inst = 32'hca00008;
      89823: inst = 32'h24822800;
      89824: inst = 32'h10a00000;
      89825: inst = 32'hca00004;
      89826: inst = 32'h38632800;
      89827: inst = 32'h38842800;
      89828: inst = 32'h10a00001;
      89829: inst = 32'hca05ee9;
      89830: inst = 32'h13e00001;
      89831: inst = 32'hfe0d96a;
      89832: inst = 32'h5be00000;
      89833: inst = 32'h8c50000;
      89834: inst = 32'h24612800;
      89835: inst = 32'h10a00000;
      89836: inst = 32'hca00008;
      89837: inst = 32'h24822800;
      89838: inst = 32'h10a00000;
      89839: inst = 32'hca00004;
      89840: inst = 32'h38632800;
      89841: inst = 32'h38842800;
      89842: inst = 32'h10a00001;
      89843: inst = 32'hca05ef7;
      89844: inst = 32'h13e00001;
      89845: inst = 32'hfe0d96a;
      89846: inst = 32'h5be00000;
      89847: inst = 32'h8c50000;
      89848: inst = 32'h24612800;
      89849: inst = 32'h10a00000;
      89850: inst = 32'hca00008;
      89851: inst = 32'h24822800;
      89852: inst = 32'h10a00000;
      89853: inst = 32'hca00004;
      89854: inst = 32'h38632800;
      89855: inst = 32'h38842800;
      89856: inst = 32'h10a00001;
      89857: inst = 32'hca05f05;
      89858: inst = 32'h13e00001;
      89859: inst = 32'hfe0d96a;
      89860: inst = 32'h5be00000;
      89861: inst = 32'h8c50000;
      89862: inst = 32'h24612800;
      89863: inst = 32'h10a00000;
      89864: inst = 32'hca00008;
      89865: inst = 32'h24822800;
      89866: inst = 32'h10a00000;
      89867: inst = 32'hca00004;
      89868: inst = 32'h38632800;
      89869: inst = 32'h38842800;
      89870: inst = 32'h10a00001;
      89871: inst = 32'hca05f13;
      89872: inst = 32'h13e00001;
      89873: inst = 32'hfe0d96a;
      89874: inst = 32'h5be00000;
      89875: inst = 32'h8c50000;
      89876: inst = 32'h24612800;
      89877: inst = 32'h10a00000;
      89878: inst = 32'hca00008;
      89879: inst = 32'h24822800;
      89880: inst = 32'h10a00000;
      89881: inst = 32'hca00004;
      89882: inst = 32'h38632800;
      89883: inst = 32'h38842800;
      89884: inst = 32'h10a00001;
      89885: inst = 32'hca05f21;
      89886: inst = 32'h13e00001;
      89887: inst = 32'hfe0d96a;
      89888: inst = 32'h5be00000;
      89889: inst = 32'h8c50000;
      89890: inst = 32'h24612800;
      89891: inst = 32'h10a00000;
      89892: inst = 32'hca00008;
      89893: inst = 32'h24822800;
      89894: inst = 32'h10a00000;
      89895: inst = 32'hca00004;
      89896: inst = 32'h38632800;
      89897: inst = 32'h38842800;
      89898: inst = 32'h10a00001;
      89899: inst = 32'hca05f2f;
      89900: inst = 32'h13e00001;
      89901: inst = 32'hfe0d96a;
      89902: inst = 32'h5be00000;
      89903: inst = 32'h8c50000;
      89904: inst = 32'h24612800;
      89905: inst = 32'h10a00000;
      89906: inst = 32'hca00008;
      89907: inst = 32'h24822800;
      89908: inst = 32'h10a00000;
      89909: inst = 32'hca00004;
      89910: inst = 32'h38632800;
      89911: inst = 32'h38842800;
      89912: inst = 32'h10a00001;
      89913: inst = 32'hca05f3d;
      89914: inst = 32'h13e00001;
      89915: inst = 32'hfe0d96a;
      89916: inst = 32'h5be00000;
      89917: inst = 32'h8c50000;
      89918: inst = 32'h24612800;
      89919: inst = 32'h10a00000;
      89920: inst = 32'hca00008;
      89921: inst = 32'h24822800;
      89922: inst = 32'h10a00000;
      89923: inst = 32'hca00004;
      89924: inst = 32'h38632800;
      89925: inst = 32'h38842800;
      89926: inst = 32'h10a00001;
      89927: inst = 32'hca05f4b;
      89928: inst = 32'h13e00001;
      89929: inst = 32'hfe0d96a;
      89930: inst = 32'h5be00000;
      89931: inst = 32'h8c50000;
      89932: inst = 32'h24612800;
      89933: inst = 32'h10a00000;
      89934: inst = 32'hca00008;
      89935: inst = 32'h24822800;
      89936: inst = 32'h10a00000;
      89937: inst = 32'hca00004;
      89938: inst = 32'h38632800;
      89939: inst = 32'h38842800;
      89940: inst = 32'h10a00001;
      89941: inst = 32'hca05f59;
      89942: inst = 32'h13e00001;
      89943: inst = 32'hfe0d96a;
      89944: inst = 32'h5be00000;
      89945: inst = 32'h8c50000;
      89946: inst = 32'h24612800;
      89947: inst = 32'h10a00000;
      89948: inst = 32'hca00008;
      89949: inst = 32'h24822800;
      89950: inst = 32'h10a00000;
      89951: inst = 32'hca00004;
      89952: inst = 32'h38632800;
      89953: inst = 32'h38842800;
      89954: inst = 32'h10a00001;
      89955: inst = 32'hca05f67;
      89956: inst = 32'h13e00001;
      89957: inst = 32'hfe0d96a;
      89958: inst = 32'h5be00000;
      89959: inst = 32'h8c50000;
      89960: inst = 32'h24612800;
      89961: inst = 32'h10a00000;
      89962: inst = 32'hca00008;
      89963: inst = 32'h24822800;
      89964: inst = 32'h10a00000;
      89965: inst = 32'hca00004;
      89966: inst = 32'h38632800;
      89967: inst = 32'h38842800;
      89968: inst = 32'h10a00001;
      89969: inst = 32'hca05f75;
      89970: inst = 32'h13e00001;
      89971: inst = 32'hfe0d96a;
      89972: inst = 32'h5be00000;
      89973: inst = 32'h8c50000;
      89974: inst = 32'h24612800;
      89975: inst = 32'h10a00000;
      89976: inst = 32'hca00008;
      89977: inst = 32'h24822800;
      89978: inst = 32'h10a00000;
      89979: inst = 32'hca00004;
      89980: inst = 32'h38632800;
      89981: inst = 32'h38842800;
      89982: inst = 32'h10a00001;
      89983: inst = 32'hca05f83;
      89984: inst = 32'h13e00001;
      89985: inst = 32'hfe0d96a;
      89986: inst = 32'h5be00000;
      89987: inst = 32'h8c50000;
      89988: inst = 32'h24612800;
      89989: inst = 32'h10a00000;
      89990: inst = 32'hca00008;
      89991: inst = 32'h24822800;
      89992: inst = 32'h10a00000;
      89993: inst = 32'hca00004;
      89994: inst = 32'h38632800;
      89995: inst = 32'h38842800;
      89996: inst = 32'h10a00001;
      89997: inst = 32'hca05f91;
      89998: inst = 32'h13e00001;
      89999: inst = 32'hfe0d96a;
      90000: inst = 32'h5be00000;
      90001: inst = 32'h8c50000;
      90002: inst = 32'h24612800;
      90003: inst = 32'h10a00000;
      90004: inst = 32'hca00008;
      90005: inst = 32'h24822800;
      90006: inst = 32'h10a00000;
      90007: inst = 32'hca00004;
      90008: inst = 32'h38632800;
      90009: inst = 32'h38842800;
      90010: inst = 32'h10a00001;
      90011: inst = 32'hca05f9f;
      90012: inst = 32'h13e00001;
      90013: inst = 32'hfe0d96a;
      90014: inst = 32'h5be00000;
      90015: inst = 32'h8c50000;
      90016: inst = 32'h24612800;
      90017: inst = 32'h10a00000;
      90018: inst = 32'hca00008;
      90019: inst = 32'h24822800;
      90020: inst = 32'h10a00000;
      90021: inst = 32'hca00004;
      90022: inst = 32'h38632800;
      90023: inst = 32'h38842800;
      90024: inst = 32'h10a00001;
      90025: inst = 32'hca05fad;
      90026: inst = 32'h13e00001;
      90027: inst = 32'hfe0d96a;
      90028: inst = 32'h5be00000;
      90029: inst = 32'h8c50000;
      90030: inst = 32'h24612800;
      90031: inst = 32'h10a00000;
      90032: inst = 32'hca00008;
      90033: inst = 32'h24822800;
      90034: inst = 32'h10a00000;
      90035: inst = 32'hca00004;
      90036: inst = 32'h38632800;
      90037: inst = 32'h38842800;
      90038: inst = 32'h10a00001;
      90039: inst = 32'hca05fbb;
      90040: inst = 32'h13e00001;
      90041: inst = 32'hfe0d96a;
      90042: inst = 32'h5be00000;
      90043: inst = 32'h8c50000;
      90044: inst = 32'h24612800;
      90045: inst = 32'h10a00000;
      90046: inst = 32'hca00008;
      90047: inst = 32'h24822800;
      90048: inst = 32'h10a00000;
      90049: inst = 32'hca00004;
      90050: inst = 32'h38632800;
      90051: inst = 32'h38842800;
      90052: inst = 32'h10a00001;
      90053: inst = 32'hca05fc9;
      90054: inst = 32'h13e00001;
      90055: inst = 32'hfe0d96a;
      90056: inst = 32'h5be00000;
      90057: inst = 32'h8c50000;
      90058: inst = 32'h24612800;
      90059: inst = 32'h10a00000;
      90060: inst = 32'hca00008;
      90061: inst = 32'h24822800;
      90062: inst = 32'h10a00000;
      90063: inst = 32'hca00004;
      90064: inst = 32'h38632800;
      90065: inst = 32'h38842800;
      90066: inst = 32'h10a00001;
      90067: inst = 32'hca05fd7;
      90068: inst = 32'h13e00001;
      90069: inst = 32'hfe0d96a;
      90070: inst = 32'h5be00000;
      90071: inst = 32'h8c50000;
      90072: inst = 32'h24612800;
      90073: inst = 32'h10a00000;
      90074: inst = 32'hca00008;
      90075: inst = 32'h24822800;
      90076: inst = 32'h10a00000;
      90077: inst = 32'hca00004;
      90078: inst = 32'h38632800;
      90079: inst = 32'h38842800;
      90080: inst = 32'h10a00001;
      90081: inst = 32'hca05fe5;
      90082: inst = 32'h13e00001;
      90083: inst = 32'hfe0d96a;
      90084: inst = 32'h5be00000;
      90085: inst = 32'h8c50000;
      90086: inst = 32'h24612800;
      90087: inst = 32'h10a00000;
      90088: inst = 32'hca00008;
      90089: inst = 32'h24822800;
      90090: inst = 32'h10a00000;
      90091: inst = 32'hca00004;
      90092: inst = 32'h38632800;
      90093: inst = 32'h38842800;
      90094: inst = 32'h10a00001;
      90095: inst = 32'hca05ff3;
      90096: inst = 32'h13e00001;
      90097: inst = 32'hfe0d96a;
      90098: inst = 32'h5be00000;
      90099: inst = 32'h8c50000;
      90100: inst = 32'h24612800;
      90101: inst = 32'h10a00000;
      90102: inst = 32'hca00008;
      90103: inst = 32'h24822800;
      90104: inst = 32'h10a00000;
      90105: inst = 32'hca00004;
      90106: inst = 32'h38632800;
      90107: inst = 32'h38842800;
      90108: inst = 32'h10a00001;
      90109: inst = 32'hca06001;
      90110: inst = 32'h13e00001;
      90111: inst = 32'hfe0d96a;
      90112: inst = 32'h5be00000;
      90113: inst = 32'h8c50000;
      90114: inst = 32'h24612800;
      90115: inst = 32'h10a00000;
      90116: inst = 32'hca00008;
      90117: inst = 32'h24822800;
      90118: inst = 32'h10a00000;
      90119: inst = 32'hca00004;
      90120: inst = 32'h38632800;
      90121: inst = 32'h38842800;
      90122: inst = 32'h10a00001;
      90123: inst = 32'hca0600f;
      90124: inst = 32'h13e00001;
      90125: inst = 32'hfe0d96a;
      90126: inst = 32'h5be00000;
      90127: inst = 32'h8c50000;
      90128: inst = 32'h24612800;
      90129: inst = 32'h10a00000;
      90130: inst = 32'hca00008;
      90131: inst = 32'h24822800;
      90132: inst = 32'h10a00000;
      90133: inst = 32'hca00004;
      90134: inst = 32'h38632800;
      90135: inst = 32'h38842800;
      90136: inst = 32'h10a00001;
      90137: inst = 32'hca0601d;
      90138: inst = 32'h13e00001;
      90139: inst = 32'hfe0d96a;
      90140: inst = 32'h5be00000;
      90141: inst = 32'h8c50000;
      90142: inst = 32'h24612800;
      90143: inst = 32'h10a00000;
      90144: inst = 32'hca00008;
      90145: inst = 32'h24822800;
      90146: inst = 32'h10a00000;
      90147: inst = 32'hca00004;
      90148: inst = 32'h38632800;
      90149: inst = 32'h38842800;
      90150: inst = 32'h10a00001;
      90151: inst = 32'hca0602b;
      90152: inst = 32'h13e00001;
      90153: inst = 32'hfe0d96a;
      90154: inst = 32'h5be00000;
      90155: inst = 32'h8c50000;
      90156: inst = 32'h24612800;
      90157: inst = 32'h10a00000;
      90158: inst = 32'hca00008;
      90159: inst = 32'h24822800;
      90160: inst = 32'h10a00000;
      90161: inst = 32'hca00004;
      90162: inst = 32'h38632800;
      90163: inst = 32'h38842800;
      90164: inst = 32'h10a00001;
      90165: inst = 32'hca06039;
      90166: inst = 32'h13e00001;
      90167: inst = 32'hfe0d96a;
      90168: inst = 32'h5be00000;
      90169: inst = 32'h8c50000;
      90170: inst = 32'h24612800;
      90171: inst = 32'h10a00000;
      90172: inst = 32'hca00008;
      90173: inst = 32'h24822800;
      90174: inst = 32'h10a00000;
      90175: inst = 32'hca00004;
      90176: inst = 32'h38632800;
      90177: inst = 32'h38842800;
      90178: inst = 32'h10a00001;
      90179: inst = 32'hca06047;
      90180: inst = 32'h13e00001;
      90181: inst = 32'hfe0d96a;
      90182: inst = 32'h5be00000;
      90183: inst = 32'h8c50000;
      90184: inst = 32'h24612800;
      90185: inst = 32'h10a00000;
      90186: inst = 32'hca00008;
      90187: inst = 32'h24822800;
      90188: inst = 32'h10a00000;
      90189: inst = 32'hca00004;
      90190: inst = 32'h38632800;
      90191: inst = 32'h38842800;
      90192: inst = 32'h10a00001;
      90193: inst = 32'hca06055;
      90194: inst = 32'h13e00001;
      90195: inst = 32'hfe0d96a;
      90196: inst = 32'h5be00000;
      90197: inst = 32'h8c50000;
      90198: inst = 32'h24612800;
      90199: inst = 32'h10a00000;
      90200: inst = 32'hca00008;
      90201: inst = 32'h24822800;
      90202: inst = 32'h10a00000;
      90203: inst = 32'hca00004;
      90204: inst = 32'h38632800;
      90205: inst = 32'h38842800;
      90206: inst = 32'h10a00001;
      90207: inst = 32'hca06063;
      90208: inst = 32'h13e00001;
      90209: inst = 32'hfe0d96a;
      90210: inst = 32'h5be00000;
      90211: inst = 32'h8c50000;
      90212: inst = 32'h24612800;
      90213: inst = 32'h10a00000;
      90214: inst = 32'hca00008;
      90215: inst = 32'h24822800;
      90216: inst = 32'h10a00000;
      90217: inst = 32'hca00004;
      90218: inst = 32'h38632800;
      90219: inst = 32'h38842800;
      90220: inst = 32'h10a00001;
      90221: inst = 32'hca06071;
      90222: inst = 32'h13e00001;
      90223: inst = 32'hfe0d96a;
      90224: inst = 32'h5be00000;
      90225: inst = 32'h8c50000;
      90226: inst = 32'h24612800;
      90227: inst = 32'h10a00000;
      90228: inst = 32'hca00008;
      90229: inst = 32'h24822800;
      90230: inst = 32'h10a00000;
      90231: inst = 32'hca00004;
      90232: inst = 32'h38632800;
      90233: inst = 32'h38842800;
      90234: inst = 32'h10a00001;
      90235: inst = 32'hca0607f;
      90236: inst = 32'h13e00001;
      90237: inst = 32'hfe0d96a;
      90238: inst = 32'h5be00000;
      90239: inst = 32'h8c50000;
      90240: inst = 32'h24612800;
      90241: inst = 32'h10a00000;
      90242: inst = 32'hca00008;
      90243: inst = 32'h24822800;
      90244: inst = 32'h10a00000;
      90245: inst = 32'hca00004;
      90246: inst = 32'h38632800;
      90247: inst = 32'h38842800;
      90248: inst = 32'h10a00001;
      90249: inst = 32'hca0608d;
      90250: inst = 32'h13e00001;
      90251: inst = 32'hfe0d96a;
      90252: inst = 32'h5be00000;
      90253: inst = 32'h8c50000;
      90254: inst = 32'h24612800;
      90255: inst = 32'h10a00000;
      90256: inst = 32'hca00008;
      90257: inst = 32'h24822800;
      90258: inst = 32'h10a00000;
      90259: inst = 32'hca00004;
      90260: inst = 32'h38632800;
      90261: inst = 32'h38842800;
      90262: inst = 32'h10a00001;
      90263: inst = 32'hca0609b;
      90264: inst = 32'h13e00001;
      90265: inst = 32'hfe0d96a;
      90266: inst = 32'h5be00000;
      90267: inst = 32'h8c50000;
      90268: inst = 32'h24612800;
      90269: inst = 32'h10a00000;
      90270: inst = 32'hca00008;
      90271: inst = 32'h24822800;
      90272: inst = 32'h10a00000;
      90273: inst = 32'hca00004;
      90274: inst = 32'h38632800;
      90275: inst = 32'h38842800;
      90276: inst = 32'h10a00001;
      90277: inst = 32'hca060a9;
      90278: inst = 32'h13e00001;
      90279: inst = 32'hfe0d96a;
      90280: inst = 32'h5be00000;
      90281: inst = 32'h8c50000;
      90282: inst = 32'h24612800;
      90283: inst = 32'h10a00000;
      90284: inst = 32'hca00009;
      90285: inst = 32'h24822800;
      90286: inst = 32'h10a00000;
      90287: inst = 32'hca00004;
      90288: inst = 32'h38632800;
      90289: inst = 32'h38842800;
      90290: inst = 32'h10a00001;
      90291: inst = 32'hca060b7;
      90292: inst = 32'h13e00001;
      90293: inst = 32'hfe0d96a;
      90294: inst = 32'h5be00000;
      90295: inst = 32'h8c50000;
      90296: inst = 32'h24612800;
      90297: inst = 32'h10a00000;
      90298: inst = 32'hca00009;
      90299: inst = 32'h24822800;
      90300: inst = 32'h10a00000;
      90301: inst = 32'hca00004;
      90302: inst = 32'h38632800;
      90303: inst = 32'h38842800;
      90304: inst = 32'h10a00001;
      90305: inst = 32'hca060c5;
      90306: inst = 32'h13e00001;
      90307: inst = 32'hfe0d96a;
      90308: inst = 32'h5be00000;
      90309: inst = 32'h8c50000;
      90310: inst = 32'h24612800;
      90311: inst = 32'h10a00000;
      90312: inst = 32'hca00009;
      90313: inst = 32'h24822800;
      90314: inst = 32'h10a00000;
      90315: inst = 32'hca00004;
      90316: inst = 32'h38632800;
      90317: inst = 32'h38842800;
      90318: inst = 32'h10a00001;
      90319: inst = 32'hca060d3;
      90320: inst = 32'h13e00001;
      90321: inst = 32'hfe0d96a;
      90322: inst = 32'h5be00000;
      90323: inst = 32'h8c50000;
      90324: inst = 32'h24612800;
      90325: inst = 32'h10a00000;
      90326: inst = 32'hca00009;
      90327: inst = 32'h24822800;
      90328: inst = 32'h10a00000;
      90329: inst = 32'hca00004;
      90330: inst = 32'h38632800;
      90331: inst = 32'h38842800;
      90332: inst = 32'h10a00001;
      90333: inst = 32'hca060e1;
      90334: inst = 32'h13e00001;
      90335: inst = 32'hfe0d96a;
      90336: inst = 32'h5be00000;
      90337: inst = 32'h8c50000;
      90338: inst = 32'h24612800;
      90339: inst = 32'h10a00000;
      90340: inst = 32'hca00009;
      90341: inst = 32'h24822800;
      90342: inst = 32'h10a00000;
      90343: inst = 32'hca00004;
      90344: inst = 32'h38632800;
      90345: inst = 32'h38842800;
      90346: inst = 32'h10a00001;
      90347: inst = 32'hca060ef;
      90348: inst = 32'h13e00001;
      90349: inst = 32'hfe0d96a;
      90350: inst = 32'h5be00000;
      90351: inst = 32'h8c50000;
      90352: inst = 32'h24612800;
      90353: inst = 32'h10a00000;
      90354: inst = 32'hca00009;
      90355: inst = 32'h24822800;
      90356: inst = 32'h10a00000;
      90357: inst = 32'hca00004;
      90358: inst = 32'h38632800;
      90359: inst = 32'h38842800;
      90360: inst = 32'h10a00001;
      90361: inst = 32'hca060fd;
      90362: inst = 32'h13e00001;
      90363: inst = 32'hfe0d96a;
      90364: inst = 32'h5be00000;
      90365: inst = 32'h8c50000;
      90366: inst = 32'h24612800;
      90367: inst = 32'h10a00000;
      90368: inst = 32'hca00009;
      90369: inst = 32'h24822800;
      90370: inst = 32'h10a00000;
      90371: inst = 32'hca00004;
      90372: inst = 32'h38632800;
      90373: inst = 32'h38842800;
      90374: inst = 32'h10a00001;
      90375: inst = 32'hca0610b;
      90376: inst = 32'h13e00001;
      90377: inst = 32'hfe0d96a;
      90378: inst = 32'h5be00000;
      90379: inst = 32'h8c50000;
      90380: inst = 32'h24612800;
      90381: inst = 32'h10a00000;
      90382: inst = 32'hca00009;
      90383: inst = 32'h24822800;
      90384: inst = 32'h10a00000;
      90385: inst = 32'hca00004;
      90386: inst = 32'h38632800;
      90387: inst = 32'h38842800;
      90388: inst = 32'h10a00001;
      90389: inst = 32'hca06119;
      90390: inst = 32'h13e00001;
      90391: inst = 32'hfe0d96a;
      90392: inst = 32'h5be00000;
      90393: inst = 32'h8c50000;
      90394: inst = 32'h24612800;
      90395: inst = 32'h10a00000;
      90396: inst = 32'hca00009;
      90397: inst = 32'h24822800;
      90398: inst = 32'h10a00000;
      90399: inst = 32'hca00004;
      90400: inst = 32'h38632800;
      90401: inst = 32'h38842800;
      90402: inst = 32'h10a00001;
      90403: inst = 32'hca06127;
      90404: inst = 32'h13e00001;
      90405: inst = 32'hfe0d96a;
      90406: inst = 32'h5be00000;
      90407: inst = 32'h8c50000;
      90408: inst = 32'h24612800;
      90409: inst = 32'h10a00000;
      90410: inst = 32'hca00009;
      90411: inst = 32'h24822800;
      90412: inst = 32'h10a00000;
      90413: inst = 32'hca00004;
      90414: inst = 32'h38632800;
      90415: inst = 32'h38842800;
      90416: inst = 32'h10a00001;
      90417: inst = 32'hca06135;
      90418: inst = 32'h13e00001;
      90419: inst = 32'hfe0d96a;
      90420: inst = 32'h5be00000;
      90421: inst = 32'h8c50000;
      90422: inst = 32'h24612800;
      90423: inst = 32'h10a00000;
      90424: inst = 32'hca00009;
      90425: inst = 32'h24822800;
      90426: inst = 32'h10a00000;
      90427: inst = 32'hca00004;
      90428: inst = 32'h38632800;
      90429: inst = 32'h38842800;
      90430: inst = 32'h10a00001;
      90431: inst = 32'hca06143;
      90432: inst = 32'h13e00001;
      90433: inst = 32'hfe0d96a;
      90434: inst = 32'h5be00000;
      90435: inst = 32'h8c50000;
      90436: inst = 32'h24612800;
      90437: inst = 32'h10a00000;
      90438: inst = 32'hca00009;
      90439: inst = 32'h24822800;
      90440: inst = 32'h10a00000;
      90441: inst = 32'hca00004;
      90442: inst = 32'h38632800;
      90443: inst = 32'h38842800;
      90444: inst = 32'h10a00001;
      90445: inst = 32'hca06151;
      90446: inst = 32'h13e00001;
      90447: inst = 32'hfe0d96a;
      90448: inst = 32'h5be00000;
      90449: inst = 32'h8c50000;
      90450: inst = 32'h24612800;
      90451: inst = 32'h10a00000;
      90452: inst = 32'hca00009;
      90453: inst = 32'h24822800;
      90454: inst = 32'h10a00000;
      90455: inst = 32'hca00004;
      90456: inst = 32'h38632800;
      90457: inst = 32'h38842800;
      90458: inst = 32'h10a00001;
      90459: inst = 32'hca0615f;
      90460: inst = 32'h13e00001;
      90461: inst = 32'hfe0d96a;
      90462: inst = 32'h5be00000;
      90463: inst = 32'h8c50000;
      90464: inst = 32'h24612800;
      90465: inst = 32'h10a00000;
      90466: inst = 32'hca00009;
      90467: inst = 32'h24822800;
      90468: inst = 32'h10a00000;
      90469: inst = 32'hca00004;
      90470: inst = 32'h38632800;
      90471: inst = 32'h38842800;
      90472: inst = 32'h10a00001;
      90473: inst = 32'hca0616d;
      90474: inst = 32'h13e00001;
      90475: inst = 32'hfe0d96a;
      90476: inst = 32'h5be00000;
      90477: inst = 32'h8c50000;
      90478: inst = 32'h24612800;
      90479: inst = 32'h10a00000;
      90480: inst = 32'hca00009;
      90481: inst = 32'h24822800;
      90482: inst = 32'h10a00000;
      90483: inst = 32'hca00004;
      90484: inst = 32'h38632800;
      90485: inst = 32'h38842800;
      90486: inst = 32'h10a00001;
      90487: inst = 32'hca0617b;
      90488: inst = 32'h13e00001;
      90489: inst = 32'hfe0d96a;
      90490: inst = 32'h5be00000;
      90491: inst = 32'h8c50000;
      90492: inst = 32'h24612800;
      90493: inst = 32'h10a00000;
      90494: inst = 32'hca00009;
      90495: inst = 32'h24822800;
      90496: inst = 32'h10a00000;
      90497: inst = 32'hca00004;
      90498: inst = 32'h38632800;
      90499: inst = 32'h38842800;
      90500: inst = 32'h10a00001;
      90501: inst = 32'hca06189;
      90502: inst = 32'h13e00001;
      90503: inst = 32'hfe0d96a;
      90504: inst = 32'h5be00000;
      90505: inst = 32'h8c50000;
      90506: inst = 32'h24612800;
      90507: inst = 32'h10a00000;
      90508: inst = 32'hca00009;
      90509: inst = 32'h24822800;
      90510: inst = 32'h10a00000;
      90511: inst = 32'hca00004;
      90512: inst = 32'h38632800;
      90513: inst = 32'h38842800;
      90514: inst = 32'h10a00001;
      90515: inst = 32'hca06197;
      90516: inst = 32'h13e00001;
      90517: inst = 32'hfe0d96a;
      90518: inst = 32'h5be00000;
      90519: inst = 32'h8c50000;
      90520: inst = 32'h24612800;
      90521: inst = 32'h10a00000;
      90522: inst = 32'hca00009;
      90523: inst = 32'h24822800;
      90524: inst = 32'h10a00000;
      90525: inst = 32'hca00004;
      90526: inst = 32'h38632800;
      90527: inst = 32'h38842800;
      90528: inst = 32'h10a00001;
      90529: inst = 32'hca061a5;
      90530: inst = 32'h13e00001;
      90531: inst = 32'hfe0d96a;
      90532: inst = 32'h5be00000;
      90533: inst = 32'h8c50000;
      90534: inst = 32'h24612800;
      90535: inst = 32'h10a00000;
      90536: inst = 32'hca00009;
      90537: inst = 32'h24822800;
      90538: inst = 32'h10a00000;
      90539: inst = 32'hca00004;
      90540: inst = 32'h38632800;
      90541: inst = 32'h38842800;
      90542: inst = 32'h10a00001;
      90543: inst = 32'hca061b3;
      90544: inst = 32'h13e00001;
      90545: inst = 32'hfe0d96a;
      90546: inst = 32'h5be00000;
      90547: inst = 32'h8c50000;
      90548: inst = 32'h24612800;
      90549: inst = 32'h10a00000;
      90550: inst = 32'hca00009;
      90551: inst = 32'h24822800;
      90552: inst = 32'h10a00000;
      90553: inst = 32'hca00004;
      90554: inst = 32'h38632800;
      90555: inst = 32'h38842800;
      90556: inst = 32'h10a00001;
      90557: inst = 32'hca061c1;
      90558: inst = 32'h13e00001;
      90559: inst = 32'hfe0d96a;
      90560: inst = 32'h5be00000;
      90561: inst = 32'h8c50000;
      90562: inst = 32'h24612800;
      90563: inst = 32'h10a00000;
      90564: inst = 32'hca00009;
      90565: inst = 32'h24822800;
      90566: inst = 32'h10a00000;
      90567: inst = 32'hca00004;
      90568: inst = 32'h38632800;
      90569: inst = 32'h38842800;
      90570: inst = 32'h10a00001;
      90571: inst = 32'hca061cf;
      90572: inst = 32'h13e00001;
      90573: inst = 32'hfe0d96a;
      90574: inst = 32'h5be00000;
      90575: inst = 32'h8c50000;
      90576: inst = 32'h24612800;
      90577: inst = 32'h10a00000;
      90578: inst = 32'hca00009;
      90579: inst = 32'h24822800;
      90580: inst = 32'h10a00000;
      90581: inst = 32'hca00004;
      90582: inst = 32'h38632800;
      90583: inst = 32'h38842800;
      90584: inst = 32'h10a00001;
      90585: inst = 32'hca061dd;
      90586: inst = 32'h13e00001;
      90587: inst = 32'hfe0d96a;
      90588: inst = 32'h5be00000;
      90589: inst = 32'h8c50000;
      90590: inst = 32'h24612800;
      90591: inst = 32'h10a00000;
      90592: inst = 32'hca00009;
      90593: inst = 32'h24822800;
      90594: inst = 32'h10a00000;
      90595: inst = 32'hca00004;
      90596: inst = 32'h38632800;
      90597: inst = 32'h38842800;
      90598: inst = 32'h10a00001;
      90599: inst = 32'hca061eb;
      90600: inst = 32'h13e00001;
      90601: inst = 32'hfe0d96a;
      90602: inst = 32'h5be00000;
      90603: inst = 32'h8c50000;
      90604: inst = 32'h24612800;
      90605: inst = 32'h10a00000;
      90606: inst = 32'hca00009;
      90607: inst = 32'h24822800;
      90608: inst = 32'h10a00000;
      90609: inst = 32'hca00004;
      90610: inst = 32'h38632800;
      90611: inst = 32'h38842800;
      90612: inst = 32'h10a00001;
      90613: inst = 32'hca061f9;
      90614: inst = 32'h13e00001;
      90615: inst = 32'hfe0d96a;
      90616: inst = 32'h5be00000;
      90617: inst = 32'h8c50000;
      90618: inst = 32'h24612800;
      90619: inst = 32'h10a00000;
      90620: inst = 32'hca00009;
      90621: inst = 32'h24822800;
      90622: inst = 32'h10a00000;
      90623: inst = 32'hca00004;
      90624: inst = 32'h38632800;
      90625: inst = 32'h38842800;
      90626: inst = 32'h10a00001;
      90627: inst = 32'hca06207;
      90628: inst = 32'h13e00001;
      90629: inst = 32'hfe0d96a;
      90630: inst = 32'h5be00000;
      90631: inst = 32'h8c50000;
      90632: inst = 32'h24612800;
      90633: inst = 32'h10a00000;
      90634: inst = 32'hca00009;
      90635: inst = 32'h24822800;
      90636: inst = 32'h10a00000;
      90637: inst = 32'hca00004;
      90638: inst = 32'h38632800;
      90639: inst = 32'h38842800;
      90640: inst = 32'h10a00001;
      90641: inst = 32'hca06215;
      90642: inst = 32'h13e00001;
      90643: inst = 32'hfe0d96a;
      90644: inst = 32'h5be00000;
      90645: inst = 32'h8c50000;
      90646: inst = 32'h24612800;
      90647: inst = 32'h10a00000;
      90648: inst = 32'hca00009;
      90649: inst = 32'h24822800;
      90650: inst = 32'h10a00000;
      90651: inst = 32'hca00004;
      90652: inst = 32'h38632800;
      90653: inst = 32'h38842800;
      90654: inst = 32'h10a00001;
      90655: inst = 32'hca06223;
      90656: inst = 32'h13e00001;
      90657: inst = 32'hfe0d96a;
      90658: inst = 32'h5be00000;
      90659: inst = 32'h8c50000;
      90660: inst = 32'h24612800;
      90661: inst = 32'h10a00000;
      90662: inst = 32'hca00009;
      90663: inst = 32'h24822800;
      90664: inst = 32'h10a00000;
      90665: inst = 32'hca00004;
      90666: inst = 32'h38632800;
      90667: inst = 32'h38842800;
      90668: inst = 32'h10a00001;
      90669: inst = 32'hca06231;
      90670: inst = 32'h13e00001;
      90671: inst = 32'hfe0d96a;
      90672: inst = 32'h5be00000;
      90673: inst = 32'h8c50000;
      90674: inst = 32'h24612800;
      90675: inst = 32'h10a00000;
      90676: inst = 32'hca00009;
      90677: inst = 32'h24822800;
      90678: inst = 32'h10a00000;
      90679: inst = 32'hca00004;
      90680: inst = 32'h38632800;
      90681: inst = 32'h38842800;
      90682: inst = 32'h10a00001;
      90683: inst = 32'hca0623f;
      90684: inst = 32'h13e00001;
      90685: inst = 32'hfe0d96a;
      90686: inst = 32'h5be00000;
      90687: inst = 32'h8c50000;
      90688: inst = 32'h24612800;
      90689: inst = 32'h10a00000;
      90690: inst = 32'hca00009;
      90691: inst = 32'h24822800;
      90692: inst = 32'h10a00000;
      90693: inst = 32'hca00004;
      90694: inst = 32'h38632800;
      90695: inst = 32'h38842800;
      90696: inst = 32'h10a00001;
      90697: inst = 32'hca0624d;
      90698: inst = 32'h13e00001;
      90699: inst = 32'hfe0d96a;
      90700: inst = 32'h5be00000;
      90701: inst = 32'h8c50000;
      90702: inst = 32'h24612800;
      90703: inst = 32'h10a00000;
      90704: inst = 32'hca00009;
      90705: inst = 32'h24822800;
      90706: inst = 32'h10a00000;
      90707: inst = 32'hca00004;
      90708: inst = 32'h38632800;
      90709: inst = 32'h38842800;
      90710: inst = 32'h10a00001;
      90711: inst = 32'hca0625b;
      90712: inst = 32'h13e00001;
      90713: inst = 32'hfe0d96a;
      90714: inst = 32'h5be00000;
      90715: inst = 32'h8c50000;
      90716: inst = 32'h24612800;
      90717: inst = 32'h10a00000;
      90718: inst = 32'hca00009;
      90719: inst = 32'h24822800;
      90720: inst = 32'h10a00000;
      90721: inst = 32'hca00004;
      90722: inst = 32'h38632800;
      90723: inst = 32'h38842800;
      90724: inst = 32'h10a00001;
      90725: inst = 32'hca06269;
      90726: inst = 32'h13e00001;
      90727: inst = 32'hfe0d96a;
      90728: inst = 32'h5be00000;
      90729: inst = 32'h8c50000;
      90730: inst = 32'h24612800;
      90731: inst = 32'h10a00000;
      90732: inst = 32'hca00009;
      90733: inst = 32'h24822800;
      90734: inst = 32'h10a00000;
      90735: inst = 32'hca00004;
      90736: inst = 32'h38632800;
      90737: inst = 32'h38842800;
      90738: inst = 32'h10a00001;
      90739: inst = 32'hca06277;
      90740: inst = 32'h13e00001;
      90741: inst = 32'hfe0d96a;
      90742: inst = 32'h5be00000;
      90743: inst = 32'h8c50000;
      90744: inst = 32'h24612800;
      90745: inst = 32'h10a00000;
      90746: inst = 32'hca00009;
      90747: inst = 32'h24822800;
      90748: inst = 32'h10a00000;
      90749: inst = 32'hca00004;
      90750: inst = 32'h38632800;
      90751: inst = 32'h38842800;
      90752: inst = 32'h10a00001;
      90753: inst = 32'hca06285;
      90754: inst = 32'h13e00001;
      90755: inst = 32'hfe0d96a;
      90756: inst = 32'h5be00000;
      90757: inst = 32'h8c50000;
      90758: inst = 32'h24612800;
      90759: inst = 32'h10a00000;
      90760: inst = 32'hca00009;
      90761: inst = 32'h24822800;
      90762: inst = 32'h10a00000;
      90763: inst = 32'hca00004;
      90764: inst = 32'h38632800;
      90765: inst = 32'h38842800;
      90766: inst = 32'h10a00001;
      90767: inst = 32'hca06293;
      90768: inst = 32'h13e00001;
      90769: inst = 32'hfe0d96a;
      90770: inst = 32'h5be00000;
      90771: inst = 32'h8c50000;
      90772: inst = 32'h24612800;
      90773: inst = 32'h10a00000;
      90774: inst = 32'hca00009;
      90775: inst = 32'h24822800;
      90776: inst = 32'h10a00000;
      90777: inst = 32'hca00004;
      90778: inst = 32'h38632800;
      90779: inst = 32'h38842800;
      90780: inst = 32'h10a00001;
      90781: inst = 32'hca062a1;
      90782: inst = 32'h13e00001;
      90783: inst = 32'hfe0d96a;
      90784: inst = 32'h5be00000;
      90785: inst = 32'h8c50000;
      90786: inst = 32'h24612800;
      90787: inst = 32'h10a00000;
      90788: inst = 32'hca00009;
      90789: inst = 32'h24822800;
      90790: inst = 32'h10a00000;
      90791: inst = 32'hca00004;
      90792: inst = 32'h38632800;
      90793: inst = 32'h38842800;
      90794: inst = 32'h10a00001;
      90795: inst = 32'hca062af;
      90796: inst = 32'h13e00001;
      90797: inst = 32'hfe0d96a;
      90798: inst = 32'h5be00000;
      90799: inst = 32'h8c50000;
      90800: inst = 32'h24612800;
      90801: inst = 32'h10a00000;
      90802: inst = 32'hca00009;
      90803: inst = 32'h24822800;
      90804: inst = 32'h10a00000;
      90805: inst = 32'hca00004;
      90806: inst = 32'h38632800;
      90807: inst = 32'h38842800;
      90808: inst = 32'h10a00001;
      90809: inst = 32'hca062bd;
      90810: inst = 32'h13e00001;
      90811: inst = 32'hfe0d96a;
      90812: inst = 32'h5be00000;
      90813: inst = 32'h8c50000;
      90814: inst = 32'h24612800;
      90815: inst = 32'h10a00000;
      90816: inst = 32'hca00009;
      90817: inst = 32'h24822800;
      90818: inst = 32'h10a00000;
      90819: inst = 32'hca00004;
      90820: inst = 32'h38632800;
      90821: inst = 32'h38842800;
      90822: inst = 32'h10a00001;
      90823: inst = 32'hca062cb;
      90824: inst = 32'h13e00001;
      90825: inst = 32'hfe0d96a;
      90826: inst = 32'h5be00000;
      90827: inst = 32'h8c50000;
      90828: inst = 32'h24612800;
      90829: inst = 32'h10a00000;
      90830: inst = 32'hca00009;
      90831: inst = 32'h24822800;
      90832: inst = 32'h10a00000;
      90833: inst = 32'hca00004;
      90834: inst = 32'h38632800;
      90835: inst = 32'h38842800;
      90836: inst = 32'h10a00001;
      90837: inst = 32'hca062d9;
      90838: inst = 32'h13e00001;
      90839: inst = 32'hfe0d96a;
      90840: inst = 32'h5be00000;
      90841: inst = 32'h8c50000;
      90842: inst = 32'h24612800;
      90843: inst = 32'h10a00000;
      90844: inst = 32'hca00009;
      90845: inst = 32'h24822800;
      90846: inst = 32'h10a00000;
      90847: inst = 32'hca00004;
      90848: inst = 32'h38632800;
      90849: inst = 32'h38842800;
      90850: inst = 32'h10a00001;
      90851: inst = 32'hca062e7;
      90852: inst = 32'h13e00001;
      90853: inst = 32'hfe0d96a;
      90854: inst = 32'h5be00000;
      90855: inst = 32'h8c50000;
      90856: inst = 32'h24612800;
      90857: inst = 32'h10a00000;
      90858: inst = 32'hca00009;
      90859: inst = 32'h24822800;
      90860: inst = 32'h10a00000;
      90861: inst = 32'hca00004;
      90862: inst = 32'h38632800;
      90863: inst = 32'h38842800;
      90864: inst = 32'h10a00001;
      90865: inst = 32'hca062f5;
      90866: inst = 32'h13e00001;
      90867: inst = 32'hfe0d96a;
      90868: inst = 32'h5be00000;
      90869: inst = 32'h8c50000;
      90870: inst = 32'h24612800;
      90871: inst = 32'h10a00000;
      90872: inst = 32'hca00009;
      90873: inst = 32'h24822800;
      90874: inst = 32'h10a00000;
      90875: inst = 32'hca00004;
      90876: inst = 32'h38632800;
      90877: inst = 32'h38842800;
      90878: inst = 32'h10a00001;
      90879: inst = 32'hca06303;
      90880: inst = 32'h13e00001;
      90881: inst = 32'hfe0d96a;
      90882: inst = 32'h5be00000;
      90883: inst = 32'h8c50000;
      90884: inst = 32'h24612800;
      90885: inst = 32'h10a00000;
      90886: inst = 32'hca00009;
      90887: inst = 32'h24822800;
      90888: inst = 32'h10a00000;
      90889: inst = 32'hca00004;
      90890: inst = 32'h38632800;
      90891: inst = 32'h38842800;
      90892: inst = 32'h10a00001;
      90893: inst = 32'hca06311;
      90894: inst = 32'h13e00001;
      90895: inst = 32'hfe0d96a;
      90896: inst = 32'h5be00000;
      90897: inst = 32'h8c50000;
      90898: inst = 32'h24612800;
      90899: inst = 32'h10a00000;
      90900: inst = 32'hca00009;
      90901: inst = 32'h24822800;
      90902: inst = 32'h10a00000;
      90903: inst = 32'hca00004;
      90904: inst = 32'h38632800;
      90905: inst = 32'h38842800;
      90906: inst = 32'h10a00001;
      90907: inst = 32'hca0631f;
      90908: inst = 32'h13e00001;
      90909: inst = 32'hfe0d96a;
      90910: inst = 32'h5be00000;
      90911: inst = 32'h8c50000;
      90912: inst = 32'h24612800;
      90913: inst = 32'h10a00000;
      90914: inst = 32'hca00009;
      90915: inst = 32'h24822800;
      90916: inst = 32'h10a00000;
      90917: inst = 32'hca00004;
      90918: inst = 32'h38632800;
      90919: inst = 32'h38842800;
      90920: inst = 32'h10a00001;
      90921: inst = 32'hca0632d;
      90922: inst = 32'h13e00001;
      90923: inst = 32'hfe0d96a;
      90924: inst = 32'h5be00000;
      90925: inst = 32'h8c50000;
      90926: inst = 32'h24612800;
      90927: inst = 32'h10a00000;
      90928: inst = 32'hca00009;
      90929: inst = 32'h24822800;
      90930: inst = 32'h10a00000;
      90931: inst = 32'hca00004;
      90932: inst = 32'h38632800;
      90933: inst = 32'h38842800;
      90934: inst = 32'h10a00001;
      90935: inst = 32'hca0633b;
      90936: inst = 32'h13e00001;
      90937: inst = 32'hfe0d96a;
      90938: inst = 32'h5be00000;
      90939: inst = 32'h8c50000;
      90940: inst = 32'h24612800;
      90941: inst = 32'h10a00000;
      90942: inst = 32'hca00009;
      90943: inst = 32'h24822800;
      90944: inst = 32'h10a00000;
      90945: inst = 32'hca00004;
      90946: inst = 32'h38632800;
      90947: inst = 32'h38842800;
      90948: inst = 32'h10a00001;
      90949: inst = 32'hca06349;
      90950: inst = 32'h13e00001;
      90951: inst = 32'hfe0d96a;
      90952: inst = 32'h5be00000;
      90953: inst = 32'h8c50000;
      90954: inst = 32'h24612800;
      90955: inst = 32'h10a00000;
      90956: inst = 32'hca00009;
      90957: inst = 32'h24822800;
      90958: inst = 32'h10a00000;
      90959: inst = 32'hca00004;
      90960: inst = 32'h38632800;
      90961: inst = 32'h38842800;
      90962: inst = 32'h10a00001;
      90963: inst = 32'hca06357;
      90964: inst = 32'h13e00001;
      90965: inst = 32'hfe0d96a;
      90966: inst = 32'h5be00000;
      90967: inst = 32'h8c50000;
      90968: inst = 32'h24612800;
      90969: inst = 32'h10a00000;
      90970: inst = 32'hca00009;
      90971: inst = 32'h24822800;
      90972: inst = 32'h10a00000;
      90973: inst = 32'hca00004;
      90974: inst = 32'h38632800;
      90975: inst = 32'h38842800;
      90976: inst = 32'h10a00001;
      90977: inst = 32'hca06365;
      90978: inst = 32'h13e00001;
      90979: inst = 32'hfe0d96a;
      90980: inst = 32'h5be00000;
      90981: inst = 32'h8c50000;
      90982: inst = 32'h24612800;
      90983: inst = 32'h10a00000;
      90984: inst = 32'hca00009;
      90985: inst = 32'h24822800;
      90986: inst = 32'h10a00000;
      90987: inst = 32'hca00004;
      90988: inst = 32'h38632800;
      90989: inst = 32'h38842800;
      90990: inst = 32'h10a00001;
      90991: inst = 32'hca06373;
      90992: inst = 32'h13e00001;
      90993: inst = 32'hfe0d96a;
      90994: inst = 32'h5be00000;
      90995: inst = 32'h8c50000;
      90996: inst = 32'h24612800;
      90997: inst = 32'h10a00000;
      90998: inst = 32'hca00009;
      90999: inst = 32'h24822800;
      91000: inst = 32'h10a00000;
      91001: inst = 32'hca00004;
      91002: inst = 32'h38632800;
      91003: inst = 32'h38842800;
      91004: inst = 32'h10a00001;
      91005: inst = 32'hca06381;
      91006: inst = 32'h13e00001;
      91007: inst = 32'hfe0d96a;
      91008: inst = 32'h5be00000;
      91009: inst = 32'h8c50000;
      91010: inst = 32'h24612800;
      91011: inst = 32'h10a00000;
      91012: inst = 32'hca00009;
      91013: inst = 32'h24822800;
      91014: inst = 32'h10a00000;
      91015: inst = 32'hca00004;
      91016: inst = 32'h38632800;
      91017: inst = 32'h38842800;
      91018: inst = 32'h10a00001;
      91019: inst = 32'hca0638f;
      91020: inst = 32'h13e00001;
      91021: inst = 32'hfe0d96a;
      91022: inst = 32'h5be00000;
      91023: inst = 32'h8c50000;
      91024: inst = 32'h24612800;
      91025: inst = 32'h10a00000;
      91026: inst = 32'hca00009;
      91027: inst = 32'h24822800;
      91028: inst = 32'h10a00000;
      91029: inst = 32'hca00004;
      91030: inst = 32'h38632800;
      91031: inst = 32'h38842800;
      91032: inst = 32'h10a00001;
      91033: inst = 32'hca0639d;
      91034: inst = 32'h13e00001;
      91035: inst = 32'hfe0d96a;
      91036: inst = 32'h5be00000;
      91037: inst = 32'h8c50000;
      91038: inst = 32'h24612800;
      91039: inst = 32'h10a00000;
      91040: inst = 32'hca00009;
      91041: inst = 32'h24822800;
      91042: inst = 32'h10a00000;
      91043: inst = 32'hca00004;
      91044: inst = 32'h38632800;
      91045: inst = 32'h38842800;
      91046: inst = 32'h10a00001;
      91047: inst = 32'hca063ab;
      91048: inst = 32'h13e00001;
      91049: inst = 32'hfe0d96a;
      91050: inst = 32'h5be00000;
      91051: inst = 32'h8c50000;
      91052: inst = 32'h24612800;
      91053: inst = 32'h10a00000;
      91054: inst = 32'hca00009;
      91055: inst = 32'h24822800;
      91056: inst = 32'h10a00000;
      91057: inst = 32'hca00004;
      91058: inst = 32'h38632800;
      91059: inst = 32'h38842800;
      91060: inst = 32'h10a00001;
      91061: inst = 32'hca063b9;
      91062: inst = 32'h13e00001;
      91063: inst = 32'hfe0d96a;
      91064: inst = 32'h5be00000;
      91065: inst = 32'h8c50000;
      91066: inst = 32'h24612800;
      91067: inst = 32'h10a00000;
      91068: inst = 32'hca00009;
      91069: inst = 32'h24822800;
      91070: inst = 32'h10a00000;
      91071: inst = 32'hca00004;
      91072: inst = 32'h38632800;
      91073: inst = 32'h38842800;
      91074: inst = 32'h10a00001;
      91075: inst = 32'hca063c7;
      91076: inst = 32'h13e00001;
      91077: inst = 32'hfe0d96a;
      91078: inst = 32'h5be00000;
      91079: inst = 32'h8c50000;
      91080: inst = 32'h24612800;
      91081: inst = 32'h10a00000;
      91082: inst = 32'hca00009;
      91083: inst = 32'h24822800;
      91084: inst = 32'h10a00000;
      91085: inst = 32'hca00004;
      91086: inst = 32'h38632800;
      91087: inst = 32'h38842800;
      91088: inst = 32'h10a00001;
      91089: inst = 32'hca063d5;
      91090: inst = 32'h13e00001;
      91091: inst = 32'hfe0d96a;
      91092: inst = 32'h5be00000;
      91093: inst = 32'h8c50000;
      91094: inst = 32'h24612800;
      91095: inst = 32'h10a00000;
      91096: inst = 32'hca00009;
      91097: inst = 32'h24822800;
      91098: inst = 32'h10a00000;
      91099: inst = 32'hca00004;
      91100: inst = 32'h38632800;
      91101: inst = 32'h38842800;
      91102: inst = 32'h10a00001;
      91103: inst = 32'hca063e3;
      91104: inst = 32'h13e00001;
      91105: inst = 32'hfe0d96a;
      91106: inst = 32'h5be00000;
      91107: inst = 32'h8c50000;
      91108: inst = 32'h24612800;
      91109: inst = 32'h10a00000;
      91110: inst = 32'hca00009;
      91111: inst = 32'h24822800;
      91112: inst = 32'h10a00000;
      91113: inst = 32'hca00004;
      91114: inst = 32'h38632800;
      91115: inst = 32'h38842800;
      91116: inst = 32'h10a00001;
      91117: inst = 32'hca063f1;
      91118: inst = 32'h13e00001;
      91119: inst = 32'hfe0d96a;
      91120: inst = 32'h5be00000;
      91121: inst = 32'h8c50000;
      91122: inst = 32'h24612800;
      91123: inst = 32'h10a00000;
      91124: inst = 32'hca00009;
      91125: inst = 32'h24822800;
      91126: inst = 32'h10a00000;
      91127: inst = 32'hca00004;
      91128: inst = 32'h38632800;
      91129: inst = 32'h38842800;
      91130: inst = 32'h10a00001;
      91131: inst = 32'hca063ff;
      91132: inst = 32'h13e00001;
      91133: inst = 32'hfe0d96a;
      91134: inst = 32'h5be00000;
      91135: inst = 32'h8c50000;
      91136: inst = 32'h24612800;
      91137: inst = 32'h10a00000;
      91138: inst = 32'hca00009;
      91139: inst = 32'h24822800;
      91140: inst = 32'h10a00000;
      91141: inst = 32'hca00004;
      91142: inst = 32'h38632800;
      91143: inst = 32'h38842800;
      91144: inst = 32'h10a00001;
      91145: inst = 32'hca0640d;
      91146: inst = 32'h13e00001;
      91147: inst = 32'hfe0d96a;
      91148: inst = 32'h5be00000;
      91149: inst = 32'h8c50000;
      91150: inst = 32'h24612800;
      91151: inst = 32'h10a00000;
      91152: inst = 32'hca00009;
      91153: inst = 32'h24822800;
      91154: inst = 32'h10a00000;
      91155: inst = 32'hca00004;
      91156: inst = 32'h38632800;
      91157: inst = 32'h38842800;
      91158: inst = 32'h10a00001;
      91159: inst = 32'hca0641b;
      91160: inst = 32'h13e00001;
      91161: inst = 32'hfe0d96a;
      91162: inst = 32'h5be00000;
      91163: inst = 32'h8c50000;
      91164: inst = 32'h24612800;
      91165: inst = 32'h10a00000;
      91166: inst = 32'hca00009;
      91167: inst = 32'h24822800;
      91168: inst = 32'h10a00000;
      91169: inst = 32'hca00004;
      91170: inst = 32'h38632800;
      91171: inst = 32'h38842800;
      91172: inst = 32'h10a00001;
      91173: inst = 32'hca06429;
      91174: inst = 32'h13e00001;
      91175: inst = 32'hfe0d96a;
      91176: inst = 32'h5be00000;
      91177: inst = 32'h8c50000;
      91178: inst = 32'h24612800;
      91179: inst = 32'h10a00000;
      91180: inst = 32'hca00009;
      91181: inst = 32'h24822800;
      91182: inst = 32'h10a00000;
      91183: inst = 32'hca00004;
      91184: inst = 32'h38632800;
      91185: inst = 32'h38842800;
      91186: inst = 32'h10a00001;
      91187: inst = 32'hca06437;
      91188: inst = 32'h13e00001;
      91189: inst = 32'hfe0d96a;
      91190: inst = 32'h5be00000;
      91191: inst = 32'h8c50000;
      91192: inst = 32'h24612800;
      91193: inst = 32'h10a00000;
      91194: inst = 32'hca00009;
      91195: inst = 32'h24822800;
      91196: inst = 32'h10a00000;
      91197: inst = 32'hca00004;
      91198: inst = 32'h38632800;
      91199: inst = 32'h38842800;
      91200: inst = 32'h10a00001;
      91201: inst = 32'hca06445;
      91202: inst = 32'h13e00001;
      91203: inst = 32'hfe0d96a;
      91204: inst = 32'h5be00000;
      91205: inst = 32'h8c50000;
      91206: inst = 32'h24612800;
      91207: inst = 32'h10a00000;
      91208: inst = 32'hca00009;
      91209: inst = 32'h24822800;
      91210: inst = 32'h10a00000;
      91211: inst = 32'hca00004;
      91212: inst = 32'h38632800;
      91213: inst = 32'h38842800;
      91214: inst = 32'h10a00001;
      91215: inst = 32'hca06453;
      91216: inst = 32'h13e00001;
      91217: inst = 32'hfe0d96a;
      91218: inst = 32'h5be00000;
      91219: inst = 32'h8c50000;
      91220: inst = 32'h24612800;
      91221: inst = 32'h10a00000;
      91222: inst = 32'hca00009;
      91223: inst = 32'h24822800;
      91224: inst = 32'h10a00000;
      91225: inst = 32'hca00004;
      91226: inst = 32'h38632800;
      91227: inst = 32'h38842800;
      91228: inst = 32'h10a00001;
      91229: inst = 32'hca06461;
      91230: inst = 32'h13e00001;
      91231: inst = 32'hfe0d96a;
      91232: inst = 32'h5be00000;
      91233: inst = 32'h8c50000;
      91234: inst = 32'h24612800;
      91235: inst = 32'h10a00000;
      91236: inst = 32'hca00009;
      91237: inst = 32'h24822800;
      91238: inst = 32'h10a00000;
      91239: inst = 32'hca00004;
      91240: inst = 32'h38632800;
      91241: inst = 32'h38842800;
      91242: inst = 32'h10a00001;
      91243: inst = 32'hca0646f;
      91244: inst = 32'h13e00001;
      91245: inst = 32'hfe0d96a;
      91246: inst = 32'h5be00000;
      91247: inst = 32'h8c50000;
      91248: inst = 32'h24612800;
      91249: inst = 32'h10a00000;
      91250: inst = 32'hca00009;
      91251: inst = 32'h24822800;
      91252: inst = 32'h10a00000;
      91253: inst = 32'hca00004;
      91254: inst = 32'h38632800;
      91255: inst = 32'h38842800;
      91256: inst = 32'h10a00001;
      91257: inst = 32'hca0647d;
      91258: inst = 32'h13e00001;
      91259: inst = 32'hfe0d96a;
      91260: inst = 32'h5be00000;
      91261: inst = 32'h8c50000;
      91262: inst = 32'h24612800;
      91263: inst = 32'h10a00000;
      91264: inst = 32'hca00009;
      91265: inst = 32'h24822800;
      91266: inst = 32'h10a00000;
      91267: inst = 32'hca00004;
      91268: inst = 32'h38632800;
      91269: inst = 32'h38842800;
      91270: inst = 32'h10a00001;
      91271: inst = 32'hca0648b;
      91272: inst = 32'h13e00001;
      91273: inst = 32'hfe0d96a;
      91274: inst = 32'h5be00000;
      91275: inst = 32'h8c50000;
      91276: inst = 32'h24612800;
      91277: inst = 32'h10a00000;
      91278: inst = 32'hca00009;
      91279: inst = 32'h24822800;
      91280: inst = 32'h10a00000;
      91281: inst = 32'hca00004;
      91282: inst = 32'h38632800;
      91283: inst = 32'h38842800;
      91284: inst = 32'h10a00001;
      91285: inst = 32'hca06499;
      91286: inst = 32'h13e00001;
      91287: inst = 32'hfe0d96a;
      91288: inst = 32'h5be00000;
      91289: inst = 32'h8c50000;
      91290: inst = 32'h24612800;
      91291: inst = 32'h10a00000;
      91292: inst = 32'hca00009;
      91293: inst = 32'h24822800;
      91294: inst = 32'h10a00000;
      91295: inst = 32'hca00004;
      91296: inst = 32'h38632800;
      91297: inst = 32'h38842800;
      91298: inst = 32'h10a00001;
      91299: inst = 32'hca064a7;
      91300: inst = 32'h13e00001;
      91301: inst = 32'hfe0d96a;
      91302: inst = 32'h5be00000;
      91303: inst = 32'h8c50000;
      91304: inst = 32'h24612800;
      91305: inst = 32'h10a00000;
      91306: inst = 32'hca00009;
      91307: inst = 32'h24822800;
      91308: inst = 32'h10a00000;
      91309: inst = 32'hca00004;
      91310: inst = 32'h38632800;
      91311: inst = 32'h38842800;
      91312: inst = 32'h10a00001;
      91313: inst = 32'hca064b5;
      91314: inst = 32'h13e00001;
      91315: inst = 32'hfe0d96a;
      91316: inst = 32'h5be00000;
      91317: inst = 32'h8c50000;
      91318: inst = 32'h24612800;
      91319: inst = 32'h10a00000;
      91320: inst = 32'hca00009;
      91321: inst = 32'h24822800;
      91322: inst = 32'h10a00000;
      91323: inst = 32'hca00004;
      91324: inst = 32'h38632800;
      91325: inst = 32'h38842800;
      91326: inst = 32'h10a00001;
      91327: inst = 32'hca064c3;
      91328: inst = 32'h13e00001;
      91329: inst = 32'hfe0d96a;
      91330: inst = 32'h5be00000;
      91331: inst = 32'h8c50000;
      91332: inst = 32'h24612800;
      91333: inst = 32'h10a00000;
      91334: inst = 32'hca00009;
      91335: inst = 32'h24822800;
      91336: inst = 32'h10a00000;
      91337: inst = 32'hca00004;
      91338: inst = 32'h38632800;
      91339: inst = 32'h38842800;
      91340: inst = 32'h10a00001;
      91341: inst = 32'hca064d1;
      91342: inst = 32'h13e00001;
      91343: inst = 32'hfe0d96a;
      91344: inst = 32'h5be00000;
      91345: inst = 32'h8c50000;
      91346: inst = 32'h24612800;
      91347: inst = 32'h10a00000;
      91348: inst = 32'hca00009;
      91349: inst = 32'h24822800;
      91350: inst = 32'h10a00000;
      91351: inst = 32'hca00004;
      91352: inst = 32'h38632800;
      91353: inst = 32'h38842800;
      91354: inst = 32'h10a00001;
      91355: inst = 32'hca064df;
      91356: inst = 32'h13e00001;
      91357: inst = 32'hfe0d96a;
      91358: inst = 32'h5be00000;
      91359: inst = 32'h8c50000;
      91360: inst = 32'h24612800;
      91361: inst = 32'h10a00000;
      91362: inst = 32'hca00009;
      91363: inst = 32'h24822800;
      91364: inst = 32'h10a00000;
      91365: inst = 32'hca00004;
      91366: inst = 32'h38632800;
      91367: inst = 32'h38842800;
      91368: inst = 32'h10a00001;
      91369: inst = 32'hca064ed;
      91370: inst = 32'h13e00001;
      91371: inst = 32'hfe0d96a;
      91372: inst = 32'h5be00000;
      91373: inst = 32'h8c50000;
      91374: inst = 32'h24612800;
      91375: inst = 32'h10a00000;
      91376: inst = 32'hca00009;
      91377: inst = 32'h24822800;
      91378: inst = 32'h10a00000;
      91379: inst = 32'hca00004;
      91380: inst = 32'h38632800;
      91381: inst = 32'h38842800;
      91382: inst = 32'h10a00001;
      91383: inst = 32'hca064fb;
      91384: inst = 32'h13e00001;
      91385: inst = 32'hfe0d96a;
      91386: inst = 32'h5be00000;
      91387: inst = 32'h8c50000;
      91388: inst = 32'h24612800;
      91389: inst = 32'h10a00000;
      91390: inst = 32'hca00009;
      91391: inst = 32'h24822800;
      91392: inst = 32'h10a00000;
      91393: inst = 32'hca00004;
      91394: inst = 32'h38632800;
      91395: inst = 32'h38842800;
      91396: inst = 32'h10a00001;
      91397: inst = 32'hca06509;
      91398: inst = 32'h13e00001;
      91399: inst = 32'hfe0d96a;
      91400: inst = 32'h5be00000;
      91401: inst = 32'h8c50000;
      91402: inst = 32'h24612800;
      91403: inst = 32'h10a00000;
      91404: inst = 32'hca00009;
      91405: inst = 32'h24822800;
      91406: inst = 32'h10a00000;
      91407: inst = 32'hca00004;
      91408: inst = 32'h38632800;
      91409: inst = 32'h38842800;
      91410: inst = 32'h10a00001;
      91411: inst = 32'hca06517;
      91412: inst = 32'h13e00001;
      91413: inst = 32'hfe0d96a;
      91414: inst = 32'h5be00000;
      91415: inst = 32'h8c50000;
      91416: inst = 32'h24612800;
      91417: inst = 32'h10a00000;
      91418: inst = 32'hca00009;
      91419: inst = 32'h24822800;
      91420: inst = 32'h10a00000;
      91421: inst = 32'hca00004;
      91422: inst = 32'h38632800;
      91423: inst = 32'h38842800;
      91424: inst = 32'h10a00001;
      91425: inst = 32'hca06525;
      91426: inst = 32'h13e00001;
      91427: inst = 32'hfe0d96a;
      91428: inst = 32'h5be00000;
      91429: inst = 32'h8c50000;
      91430: inst = 32'h24612800;
      91431: inst = 32'h10a00000;
      91432: inst = 32'hca00009;
      91433: inst = 32'h24822800;
      91434: inst = 32'h10a00000;
      91435: inst = 32'hca00004;
      91436: inst = 32'h38632800;
      91437: inst = 32'h38842800;
      91438: inst = 32'h10a00001;
      91439: inst = 32'hca06533;
      91440: inst = 32'h13e00001;
      91441: inst = 32'hfe0d96a;
      91442: inst = 32'h5be00000;
      91443: inst = 32'h8c50000;
      91444: inst = 32'h24612800;
      91445: inst = 32'h10a00000;
      91446: inst = 32'hca00009;
      91447: inst = 32'h24822800;
      91448: inst = 32'h10a00000;
      91449: inst = 32'hca00004;
      91450: inst = 32'h38632800;
      91451: inst = 32'h38842800;
      91452: inst = 32'h10a00001;
      91453: inst = 32'hca06541;
      91454: inst = 32'h13e00001;
      91455: inst = 32'hfe0d96a;
      91456: inst = 32'h5be00000;
      91457: inst = 32'h8c50000;
      91458: inst = 32'h24612800;
      91459: inst = 32'h10a00000;
      91460: inst = 32'hca00009;
      91461: inst = 32'h24822800;
      91462: inst = 32'h10a00000;
      91463: inst = 32'hca00004;
      91464: inst = 32'h38632800;
      91465: inst = 32'h38842800;
      91466: inst = 32'h10a00001;
      91467: inst = 32'hca0654f;
      91468: inst = 32'h13e00001;
      91469: inst = 32'hfe0d96a;
      91470: inst = 32'h5be00000;
      91471: inst = 32'h8c50000;
      91472: inst = 32'h24612800;
      91473: inst = 32'h10a00000;
      91474: inst = 32'hca00009;
      91475: inst = 32'h24822800;
      91476: inst = 32'h10a00000;
      91477: inst = 32'hca00004;
      91478: inst = 32'h38632800;
      91479: inst = 32'h38842800;
      91480: inst = 32'h10a00001;
      91481: inst = 32'hca0655d;
      91482: inst = 32'h13e00001;
      91483: inst = 32'hfe0d96a;
      91484: inst = 32'h5be00000;
      91485: inst = 32'h8c50000;
      91486: inst = 32'h24612800;
      91487: inst = 32'h10a00000;
      91488: inst = 32'hca00009;
      91489: inst = 32'h24822800;
      91490: inst = 32'h10a00000;
      91491: inst = 32'hca00004;
      91492: inst = 32'h38632800;
      91493: inst = 32'h38842800;
      91494: inst = 32'h10a00001;
      91495: inst = 32'hca0656b;
      91496: inst = 32'h13e00001;
      91497: inst = 32'hfe0d96a;
      91498: inst = 32'h5be00000;
      91499: inst = 32'h8c50000;
      91500: inst = 32'h24612800;
      91501: inst = 32'h10a00000;
      91502: inst = 32'hca00009;
      91503: inst = 32'h24822800;
      91504: inst = 32'h10a00000;
      91505: inst = 32'hca00004;
      91506: inst = 32'h38632800;
      91507: inst = 32'h38842800;
      91508: inst = 32'h10a00001;
      91509: inst = 32'hca06579;
      91510: inst = 32'h13e00001;
      91511: inst = 32'hfe0d96a;
      91512: inst = 32'h5be00000;
      91513: inst = 32'h8c50000;
      91514: inst = 32'h24612800;
      91515: inst = 32'h10a00000;
      91516: inst = 32'hca00009;
      91517: inst = 32'h24822800;
      91518: inst = 32'h10a00000;
      91519: inst = 32'hca00004;
      91520: inst = 32'h38632800;
      91521: inst = 32'h38842800;
      91522: inst = 32'h10a00001;
      91523: inst = 32'hca06587;
      91524: inst = 32'h13e00001;
      91525: inst = 32'hfe0d96a;
      91526: inst = 32'h5be00000;
      91527: inst = 32'h8c50000;
      91528: inst = 32'h24612800;
      91529: inst = 32'h10a00000;
      91530: inst = 32'hca00009;
      91531: inst = 32'h24822800;
      91532: inst = 32'h10a00000;
      91533: inst = 32'hca00004;
      91534: inst = 32'h38632800;
      91535: inst = 32'h38842800;
      91536: inst = 32'h10a00001;
      91537: inst = 32'hca06595;
      91538: inst = 32'h13e00001;
      91539: inst = 32'hfe0d96a;
      91540: inst = 32'h5be00000;
      91541: inst = 32'h8c50000;
      91542: inst = 32'h24612800;
      91543: inst = 32'h10a00000;
      91544: inst = 32'hca00009;
      91545: inst = 32'h24822800;
      91546: inst = 32'h10a00000;
      91547: inst = 32'hca00004;
      91548: inst = 32'h38632800;
      91549: inst = 32'h38842800;
      91550: inst = 32'h10a00001;
      91551: inst = 32'hca065a3;
      91552: inst = 32'h13e00001;
      91553: inst = 32'hfe0d96a;
      91554: inst = 32'h5be00000;
      91555: inst = 32'h8c50000;
      91556: inst = 32'h24612800;
      91557: inst = 32'h10a00000;
      91558: inst = 32'hca00009;
      91559: inst = 32'h24822800;
      91560: inst = 32'h10a00000;
      91561: inst = 32'hca00004;
      91562: inst = 32'h38632800;
      91563: inst = 32'h38842800;
      91564: inst = 32'h10a00001;
      91565: inst = 32'hca065b1;
      91566: inst = 32'h13e00001;
      91567: inst = 32'hfe0d96a;
      91568: inst = 32'h5be00000;
      91569: inst = 32'h8c50000;
      91570: inst = 32'h24612800;
      91571: inst = 32'h10a00000;
      91572: inst = 32'hca00009;
      91573: inst = 32'h24822800;
      91574: inst = 32'h10a00000;
      91575: inst = 32'hca00004;
      91576: inst = 32'h38632800;
      91577: inst = 32'h38842800;
      91578: inst = 32'h10a00001;
      91579: inst = 32'hca065bf;
      91580: inst = 32'h13e00001;
      91581: inst = 32'hfe0d96a;
      91582: inst = 32'h5be00000;
      91583: inst = 32'h8c50000;
      91584: inst = 32'h24612800;
      91585: inst = 32'h10a00000;
      91586: inst = 32'hca00009;
      91587: inst = 32'h24822800;
      91588: inst = 32'h10a00000;
      91589: inst = 32'hca00004;
      91590: inst = 32'h38632800;
      91591: inst = 32'h38842800;
      91592: inst = 32'h10a00001;
      91593: inst = 32'hca065cd;
      91594: inst = 32'h13e00001;
      91595: inst = 32'hfe0d96a;
      91596: inst = 32'h5be00000;
      91597: inst = 32'h8c50000;
      91598: inst = 32'h24612800;
      91599: inst = 32'h10a00000;
      91600: inst = 32'hca00009;
      91601: inst = 32'h24822800;
      91602: inst = 32'h10a00000;
      91603: inst = 32'hca00004;
      91604: inst = 32'h38632800;
      91605: inst = 32'h38842800;
      91606: inst = 32'h10a00001;
      91607: inst = 32'hca065db;
      91608: inst = 32'h13e00001;
      91609: inst = 32'hfe0d96a;
      91610: inst = 32'h5be00000;
      91611: inst = 32'h8c50000;
      91612: inst = 32'h24612800;
      91613: inst = 32'h10a00000;
      91614: inst = 32'hca00009;
      91615: inst = 32'h24822800;
      91616: inst = 32'h10a00000;
      91617: inst = 32'hca00004;
      91618: inst = 32'h38632800;
      91619: inst = 32'h38842800;
      91620: inst = 32'h10a00001;
      91621: inst = 32'hca065e9;
      91622: inst = 32'h13e00001;
      91623: inst = 32'hfe0d96a;
      91624: inst = 32'h5be00000;
      91625: inst = 32'h8c50000;
      91626: inst = 32'h24612800;
      91627: inst = 32'h10a00000;
      91628: inst = 32'hca0000a;
      91629: inst = 32'h24822800;
      91630: inst = 32'h10a00000;
      91631: inst = 32'hca00004;
      91632: inst = 32'h38632800;
      91633: inst = 32'h38842800;
      91634: inst = 32'h10a00001;
      91635: inst = 32'hca065f7;
      91636: inst = 32'h13e00001;
      91637: inst = 32'hfe0d96a;
      91638: inst = 32'h5be00000;
      91639: inst = 32'h8c50000;
      91640: inst = 32'h24612800;
      91641: inst = 32'h10a00000;
      91642: inst = 32'hca0000a;
      91643: inst = 32'h24822800;
      91644: inst = 32'h10a00000;
      91645: inst = 32'hca00004;
      91646: inst = 32'h38632800;
      91647: inst = 32'h38842800;
      91648: inst = 32'h10a00001;
      91649: inst = 32'hca06605;
      91650: inst = 32'h13e00001;
      91651: inst = 32'hfe0d96a;
      91652: inst = 32'h5be00000;
      91653: inst = 32'h8c50000;
      91654: inst = 32'h24612800;
      91655: inst = 32'h10a00000;
      91656: inst = 32'hca0000a;
      91657: inst = 32'h24822800;
      91658: inst = 32'h10a00000;
      91659: inst = 32'hca00004;
      91660: inst = 32'h38632800;
      91661: inst = 32'h38842800;
      91662: inst = 32'h10a00001;
      91663: inst = 32'hca06613;
      91664: inst = 32'h13e00001;
      91665: inst = 32'hfe0d96a;
      91666: inst = 32'h5be00000;
      91667: inst = 32'h8c50000;
      91668: inst = 32'h24612800;
      91669: inst = 32'h10a00000;
      91670: inst = 32'hca0000a;
      91671: inst = 32'h24822800;
      91672: inst = 32'h10a00000;
      91673: inst = 32'hca00004;
      91674: inst = 32'h38632800;
      91675: inst = 32'h38842800;
      91676: inst = 32'h10a00001;
      91677: inst = 32'hca06621;
      91678: inst = 32'h13e00001;
      91679: inst = 32'hfe0d96a;
      91680: inst = 32'h5be00000;
      91681: inst = 32'h8c50000;
      91682: inst = 32'h24612800;
      91683: inst = 32'h10a00000;
      91684: inst = 32'hca0000a;
      91685: inst = 32'h24822800;
      91686: inst = 32'h10a00000;
      91687: inst = 32'hca00004;
      91688: inst = 32'h38632800;
      91689: inst = 32'h38842800;
      91690: inst = 32'h10a00001;
      91691: inst = 32'hca0662f;
      91692: inst = 32'h13e00001;
      91693: inst = 32'hfe0d96a;
      91694: inst = 32'h5be00000;
      91695: inst = 32'h8c50000;
      91696: inst = 32'h24612800;
      91697: inst = 32'h10a00000;
      91698: inst = 32'hca0000a;
      91699: inst = 32'h24822800;
      91700: inst = 32'h10a00000;
      91701: inst = 32'hca00004;
      91702: inst = 32'h38632800;
      91703: inst = 32'h38842800;
      91704: inst = 32'h10a00001;
      91705: inst = 32'hca0663d;
      91706: inst = 32'h13e00001;
      91707: inst = 32'hfe0d96a;
      91708: inst = 32'h5be00000;
      91709: inst = 32'h8c50000;
      91710: inst = 32'h24612800;
      91711: inst = 32'h10a00000;
      91712: inst = 32'hca0000a;
      91713: inst = 32'h24822800;
      91714: inst = 32'h10a00000;
      91715: inst = 32'hca00004;
      91716: inst = 32'h38632800;
      91717: inst = 32'h38842800;
      91718: inst = 32'h10a00001;
      91719: inst = 32'hca0664b;
      91720: inst = 32'h13e00001;
      91721: inst = 32'hfe0d96a;
      91722: inst = 32'h5be00000;
      91723: inst = 32'h8c50000;
      91724: inst = 32'h24612800;
      91725: inst = 32'h10a00000;
      91726: inst = 32'hca0000a;
      91727: inst = 32'h24822800;
      91728: inst = 32'h10a00000;
      91729: inst = 32'hca00004;
      91730: inst = 32'h38632800;
      91731: inst = 32'h38842800;
      91732: inst = 32'h10a00001;
      91733: inst = 32'hca06659;
      91734: inst = 32'h13e00001;
      91735: inst = 32'hfe0d96a;
      91736: inst = 32'h5be00000;
      91737: inst = 32'h8c50000;
      91738: inst = 32'h24612800;
      91739: inst = 32'h10a00000;
      91740: inst = 32'hca0000a;
      91741: inst = 32'h24822800;
      91742: inst = 32'h10a00000;
      91743: inst = 32'hca00004;
      91744: inst = 32'h38632800;
      91745: inst = 32'h38842800;
      91746: inst = 32'h10a00001;
      91747: inst = 32'hca06667;
      91748: inst = 32'h13e00001;
      91749: inst = 32'hfe0d96a;
      91750: inst = 32'h5be00000;
      91751: inst = 32'h8c50000;
      91752: inst = 32'h24612800;
      91753: inst = 32'h10a00000;
      91754: inst = 32'hca0000a;
      91755: inst = 32'h24822800;
      91756: inst = 32'h10a00000;
      91757: inst = 32'hca00004;
      91758: inst = 32'h38632800;
      91759: inst = 32'h38842800;
      91760: inst = 32'h10a00001;
      91761: inst = 32'hca06675;
      91762: inst = 32'h13e00001;
      91763: inst = 32'hfe0d96a;
      91764: inst = 32'h5be00000;
      91765: inst = 32'h8c50000;
      91766: inst = 32'h24612800;
      91767: inst = 32'h10a00000;
      91768: inst = 32'hca0000a;
      91769: inst = 32'h24822800;
      91770: inst = 32'h10a00000;
      91771: inst = 32'hca00004;
      91772: inst = 32'h38632800;
      91773: inst = 32'h38842800;
      91774: inst = 32'h10a00001;
      91775: inst = 32'hca06683;
      91776: inst = 32'h13e00001;
      91777: inst = 32'hfe0d96a;
      91778: inst = 32'h5be00000;
      91779: inst = 32'h8c50000;
      91780: inst = 32'h24612800;
      91781: inst = 32'h10a00000;
      91782: inst = 32'hca0000a;
      91783: inst = 32'h24822800;
      91784: inst = 32'h10a00000;
      91785: inst = 32'hca00004;
      91786: inst = 32'h38632800;
      91787: inst = 32'h38842800;
      91788: inst = 32'h10a00001;
      91789: inst = 32'hca06691;
      91790: inst = 32'h13e00001;
      91791: inst = 32'hfe0d96a;
      91792: inst = 32'h5be00000;
      91793: inst = 32'h8c50000;
      91794: inst = 32'h24612800;
      91795: inst = 32'h10a00000;
      91796: inst = 32'hca0000a;
      91797: inst = 32'h24822800;
      91798: inst = 32'h10a00000;
      91799: inst = 32'hca00004;
      91800: inst = 32'h38632800;
      91801: inst = 32'h38842800;
      91802: inst = 32'h10a00001;
      91803: inst = 32'hca0669f;
      91804: inst = 32'h13e00001;
      91805: inst = 32'hfe0d96a;
      91806: inst = 32'h5be00000;
      91807: inst = 32'h8c50000;
      91808: inst = 32'h24612800;
      91809: inst = 32'h10a00000;
      91810: inst = 32'hca0000a;
      91811: inst = 32'h24822800;
      91812: inst = 32'h10a00000;
      91813: inst = 32'hca00004;
      91814: inst = 32'h38632800;
      91815: inst = 32'h38842800;
      91816: inst = 32'h10a00001;
      91817: inst = 32'hca066ad;
      91818: inst = 32'h13e00001;
      91819: inst = 32'hfe0d96a;
      91820: inst = 32'h5be00000;
      91821: inst = 32'h8c50000;
      91822: inst = 32'h24612800;
      91823: inst = 32'h10a00000;
      91824: inst = 32'hca0000a;
      91825: inst = 32'h24822800;
      91826: inst = 32'h10a00000;
      91827: inst = 32'hca00004;
      91828: inst = 32'h38632800;
      91829: inst = 32'h38842800;
      91830: inst = 32'h10a00001;
      91831: inst = 32'hca066bb;
      91832: inst = 32'h13e00001;
      91833: inst = 32'hfe0d96a;
      91834: inst = 32'h5be00000;
      91835: inst = 32'h8c50000;
      91836: inst = 32'h24612800;
      91837: inst = 32'h10a00000;
      91838: inst = 32'hca0000a;
      91839: inst = 32'h24822800;
      91840: inst = 32'h10a00000;
      91841: inst = 32'hca00004;
      91842: inst = 32'h38632800;
      91843: inst = 32'h38842800;
      91844: inst = 32'h10a00001;
      91845: inst = 32'hca066c9;
      91846: inst = 32'h13e00001;
      91847: inst = 32'hfe0d96a;
      91848: inst = 32'h5be00000;
      91849: inst = 32'h8c50000;
      91850: inst = 32'h24612800;
      91851: inst = 32'h10a00000;
      91852: inst = 32'hca0000a;
      91853: inst = 32'h24822800;
      91854: inst = 32'h10a00000;
      91855: inst = 32'hca00004;
      91856: inst = 32'h38632800;
      91857: inst = 32'h38842800;
      91858: inst = 32'h10a00001;
      91859: inst = 32'hca066d7;
      91860: inst = 32'h13e00001;
      91861: inst = 32'hfe0d96a;
      91862: inst = 32'h5be00000;
      91863: inst = 32'h8c50000;
      91864: inst = 32'h24612800;
      91865: inst = 32'h10a00000;
      91866: inst = 32'hca0000a;
      91867: inst = 32'h24822800;
      91868: inst = 32'h10a00000;
      91869: inst = 32'hca00004;
      91870: inst = 32'h38632800;
      91871: inst = 32'h38842800;
      91872: inst = 32'h10a00001;
      91873: inst = 32'hca066e5;
      91874: inst = 32'h13e00001;
      91875: inst = 32'hfe0d96a;
      91876: inst = 32'h5be00000;
      91877: inst = 32'h8c50000;
      91878: inst = 32'h24612800;
      91879: inst = 32'h10a00000;
      91880: inst = 32'hca0000a;
      91881: inst = 32'h24822800;
      91882: inst = 32'h10a00000;
      91883: inst = 32'hca00004;
      91884: inst = 32'h38632800;
      91885: inst = 32'h38842800;
      91886: inst = 32'h10a00001;
      91887: inst = 32'hca066f3;
      91888: inst = 32'h13e00001;
      91889: inst = 32'hfe0d96a;
      91890: inst = 32'h5be00000;
      91891: inst = 32'h8c50000;
      91892: inst = 32'h24612800;
      91893: inst = 32'h10a00000;
      91894: inst = 32'hca0000a;
      91895: inst = 32'h24822800;
      91896: inst = 32'h10a00000;
      91897: inst = 32'hca00004;
      91898: inst = 32'h38632800;
      91899: inst = 32'h38842800;
      91900: inst = 32'h10a00001;
      91901: inst = 32'hca06701;
      91902: inst = 32'h13e00001;
      91903: inst = 32'hfe0d96a;
      91904: inst = 32'h5be00000;
      91905: inst = 32'h8c50000;
      91906: inst = 32'h24612800;
      91907: inst = 32'h10a00000;
      91908: inst = 32'hca0000a;
      91909: inst = 32'h24822800;
      91910: inst = 32'h10a00000;
      91911: inst = 32'hca00004;
      91912: inst = 32'h38632800;
      91913: inst = 32'h38842800;
      91914: inst = 32'h10a00001;
      91915: inst = 32'hca0670f;
      91916: inst = 32'h13e00001;
      91917: inst = 32'hfe0d96a;
      91918: inst = 32'h5be00000;
      91919: inst = 32'h8c50000;
      91920: inst = 32'h24612800;
      91921: inst = 32'h10a00000;
      91922: inst = 32'hca0000a;
      91923: inst = 32'h24822800;
      91924: inst = 32'h10a00000;
      91925: inst = 32'hca00004;
      91926: inst = 32'h38632800;
      91927: inst = 32'h38842800;
      91928: inst = 32'h10a00001;
      91929: inst = 32'hca0671d;
      91930: inst = 32'h13e00001;
      91931: inst = 32'hfe0d96a;
      91932: inst = 32'h5be00000;
      91933: inst = 32'h8c50000;
      91934: inst = 32'h24612800;
      91935: inst = 32'h10a00000;
      91936: inst = 32'hca0000a;
      91937: inst = 32'h24822800;
      91938: inst = 32'h10a00000;
      91939: inst = 32'hca00004;
      91940: inst = 32'h38632800;
      91941: inst = 32'h38842800;
      91942: inst = 32'h10a00001;
      91943: inst = 32'hca0672b;
      91944: inst = 32'h13e00001;
      91945: inst = 32'hfe0d96a;
      91946: inst = 32'h5be00000;
      91947: inst = 32'h8c50000;
      91948: inst = 32'h24612800;
      91949: inst = 32'h10a00000;
      91950: inst = 32'hca0000a;
      91951: inst = 32'h24822800;
      91952: inst = 32'h10a00000;
      91953: inst = 32'hca00004;
      91954: inst = 32'h38632800;
      91955: inst = 32'h38842800;
      91956: inst = 32'h10a00001;
      91957: inst = 32'hca06739;
      91958: inst = 32'h13e00001;
      91959: inst = 32'hfe0d96a;
      91960: inst = 32'h5be00000;
      91961: inst = 32'h8c50000;
      91962: inst = 32'h24612800;
      91963: inst = 32'h10a00000;
      91964: inst = 32'hca0000a;
      91965: inst = 32'h24822800;
      91966: inst = 32'h10a00000;
      91967: inst = 32'hca00004;
      91968: inst = 32'h38632800;
      91969: inst = 32'h38842800;
      91970: inst = 32'h10a00001;
      91971: inst = 32'hca06747;
      91972: inst = 32'h13e00001;
      91973: inst = 32'hfe0d96a;
      91974: inst = 32'h5be00000;
      91975: inst = 32'h8c50000;
      91976: inst = 32'h24612800;
      91977: inst = 32'h10a00000;
      91978: inst = 32'hca0000a;
      91979: inst = 32'h24822800;
      91980: inst = 32'h10a00000;
      91981: inst = 32'hca00004;
      91982: inst = 32'h38632800;
      91983: inst = 32'h38842800;
      91984: inst = 32'h10a00001;
      91985: inst = 32'hca06755;
      91986: inst = 32'h13e00001;
      91987: inst = 32'hfe0d96a;
      91988: inst = 32'h5be00000;
      91989: inst = 32'h8c50000;
      91990: inst = 32'h24612800;
      91991: inst = 32'h10a00000;
      91992: inst = 32'hca0000a;
      91993: inst = 32'h24822800;
      91994: inst = 32'h10a00000;
      91995: inst = 32'hca00004;
      91996: inst = 32'h38632800;
      91997: inst = 32'h38842800;
      91998: inst = 32'h10a00001;
      91999: inst = 32'hca06763;
      92000: inst = 32'h13e00001;
      92001: inst = 32'hfe0d96a;
      92002: inst = 32'h5be00000;
      92003: inst = 32'h8c50000;
      92004: inst = 32'h24612800;
      92005: inst = 32'h10a00000;
      92006: inst = 32'hca0000a;
      92007: inst = 32'h24822800;
      92008: inst = 32'h10a00000;
      92009: inst = 32'hca00004;
      92010: inst = 32'h38632800;
      92011: inst = 32'h38842800;
      92012: inst = 32'h10a00001;
      92013: inst = 32'hca06771;
      92014: inst = 32'h13e00001;
      92015: inst = 32'hfe0d96a;
      92016: inst = 32'h5be00000;
      92017: inst = 32'h8c50000;
      92018: inst = 32'h24612800;
      92019: inst = 32'h10a00000;
      92020: inst = 32'hca0000a;
      92021: inst = 32'h24822800;
      92022: inst = 32'h10a00000;
      92023: inst = 32'hca00004;
      92024: inst = 32'h38632800;
      92025: inst = 32'h38842800;
      92026: inst = 32'h10a00001;
      92027: inst = 32'hca0677f;
      92028: inst = 32'h13e00001;
      92029: inst = 32'hfe0d96a;
      92030: inst = 32'h5be00000;
      92031: inst = 32'h8c50000;
      92032: inst = 32'h24612800;
      92033: inst = 32'h10a00000;
      92034: inst = 32'hca0000a;
      92035: inst = 32'h24822800;
      92036: inst = 32'h10a00000;
      92037: inst = 32'hca00004;
      92038: inst = 32'h38632800;
      92039: inst = 32'h38842800;
      92040: inst = 32'h10a00001;
      92041: inst = 32'hca0678d;
      92042: inst = 32'h13e00001;
      92043: inst = 32'hfe0d96a;
      92044: inst = 32'h5be00000;
      92045: inst = 32'h8c50000;
      92046: inst = 32'h24612800;
      92047: inst = 32'h10a00000;
      92048: inst = 32'hca0000a;
      92049: inst = 32'h24822800;
      92050: inst = 32'h10a00000;
      92051: inst = 32'hca00004;
      92052: inst = 32'h38632800;
      92053: inst = 32'h38842800;
      92054: inst = 32'h10a00001;
      92055: inst = 32'hca0679b;
      92056: inst = 32'h13e00001;
      92057: inst = 32'hfe0d96a;
      92058: inst = 32'h5be00000;
      92059: inst = 32'h8c50000;
      92060: inst = 32'h24612800;
      92061: inst = 32'h10a00000;
      92062: inst = 32'hca0000a;
      92063: inst = 32'h24822800;
      92064: inst = 32'h10a00000;
      92065: inst = 32'hca00004;
      92066: inst = 32'h38632800;
      92067: inst = 32'h38842800;
      92068: inst = 32'h10a00001;
      92069: inst = 32'hca067a9;
      92070: inst = 32'h13e00001;
      92071: inst = 32'hfe0d96a;
      92072: inst = 32'h5be00000;
      92073: inst = 32'h8c50000;
      92074: inst = 32'h24612800;
      92075: inst = 32'h10a00000;
      92076: inst = 32'hca0000a;
      92077: inst = 32'h24822800;
      92078: inst = 32'h10a00000;
      92079: inst = 32'hca00004;
      92080: inst = 32'h38632800;
      92081: inst = 32'h38842800;
      92082: inst = 32'h10a00001;
      92083: inst = 32'hca067b7;
      92084: inst = 32'h13e00001;
      92085: inst = 32'hfe0d96a;
      92086: inst = 32'h5be00000;
      92087: inst = 32'h8c50000;
      92088: inst = 32'h24612800;
      92089: inst = 32'h10a00000;
      92090: inst = 32'hca0000a;
      92091: inst = 32'h24822800;
      92092: inst = 32'h10a00000;
      92093: inst = 32'hca00004;
      92094: inst = 32'h38632800;
      92095: inst = 32'h38842800;
      92096: inst = 32'h10a00001;
      92097: inst = 32'hca067c5;
      92098: inst = 32'h13e00001;
      92099: inst = 32'hfe0d96a;
      92100: inst = 32'h5be00000;
      92101: inst = 32'h8c50000;
      92102: inst = 32'h24612800;
      92103: inst = 32'h10a00000;
      92104: inst = 32'hca0000a;
      92105: inst = 32'h24822800;
      92106: inst = 32'h10a00000;
      92107: inst = 32'hca00004;
      92108: inst = 32'h38632800;
      92109: inst = 32'h38842800;
      92110: inst = 32'h10a00001;
      92111: inst = 32'hca067d3;
      92112: inst = 32'h13e00001;
      92113: inst = 32'hfe0d96a;
      92114: inst = 32'h5be00000;
      92115: inst = 32'h8c50000;
      92116: inst = 32'h24612800;
      92117: inst = 32'h10a00000;
      92118: inst = 32'hca0000a;
      92119: inst = 32'h24822800;
      92120: inst = 32'h10a00000;
      92121: inst = 32'hca00004;
      92122: inst = 32'h38632800;
      92123: inst = 32'h38842800;
      92124: inst = 32'h10a00001;
      92125: inst = 32'hca067e1;
      92126: inst = 32'h13e00001;
      92127: inst = 32'hfe0d96a;
      92128: inst = 32'h5be00000;
      92129: inst = 32'h8c50000;
      92130: inst = 32'h24612800;
      92131: inst = 32'h10a00000;
      92132: inst = 32'hca0000a;
      92133: inst = 32'h24822800;
      92134: inst = 32'h10a00000;
      92135: inst = 32'hca00004;
      92136: inst = 32'h38632800;
      92137: inst = 32'h38842800;
      92138: inst = 32'h10a00001;
      92139: inst = 32'hca067ef;
      92140: inst = 32'h13e00001;
      92141: inst = 32'hfe0d96a;
      92142: inst = 32'h5be00000;
      92143: inst = 32'h8c50000;
      92144: inst = 32'h24612800;
      92145: inst = 32'h10a00000;
      92146: inst = 32'hca0000a;
      92147: inst = 32'h24822800;
      92148: inst = 32'h10a00000;
      92149: inst = 32'hca00004;
      92150: inst = 32'h38632800;
      92151: inst = 32'h38842800;
      92152: inst = 32'h10a00001;
      92153: inst = 32'hca067fd;
      92154: inst = 32'h13e00001;
      92155: inst = 32'hfe0d96a;
      92156: inst = 32'h5be00000;
      92157: inst = 32'h8c50000;
      92158: inst = 32'h24612800;
      92159: inst = 32'h10a00000;
      92160: inst = 32'hca0000a;
      92161: inst = 32'h24822800;
      92162: inst = 32'h10a00000;
      92163: inst = 32'hca00004;
      92164: inst = 32'h38632800;
      92165: inst = 32'h38842800;
      92166: inst = 32'h10a00001;
      92167: inst = 32'hca0680b;
      92168: inst = 32'h13e00001;
      92169: inst = 32'hfe0d96a;
      92170: inst = 32'h5be00000;
      92171: inst = 32'h8c50000;
      92172: inst = 32'h24612800;
      92173: inst = 32'h10a00000;
      92174: inst = 32'hca0000a;
      92175: inst = 32'h24822800;
      92176: inst = 32'h10a00000;
      92177: inst = 32'hca00004;
      92178: inst = 32'h38632800;
      92179: inst = 32'h38842800;
      92180: inst = 32'h10a00001;
      92181: inst = 32'hca06819;
      92182: inst = 32'h13e00001;
      92183: inst = 32'hfe0d96a;
      92184: inst = 32'h5be00000;
      92185: inst = 32'h8c50000;
      92186: inst = 32'h24612800;
      92187: inst = 32'h10a00000;
      92188: inst = 32'hca0000a;
      92189: inst = 32'h24822800;
      92190: inst = 32'h10a00000;
      92191: inst = 32'hca00004;
      92192: inst = 32'h38632800;
      92193: inst = 32'h38842800;
      92194: inst = 32'h10a00001;
      92195: inst = 32'hca06827;
      92196: inst = 32'h13e00001;
      92197: inst = 32'hfe0d96a;
      92198: inst = 32'h5be00000;
      92199: inst = 32'h8c50000;
      92200: inst = 32'h24612800;
      92201: inst = 32'h10a00000;
      92202: inst = 32'hca0000a;
      92203: inst = 32'h24822800;
      92204: inst = 32'h10a00000;
      92205: inst = 32'hca00004;
      92206: inst = 32'h38632800;
      92207: inst = 32'h38842800;
      92208: inst = 32'h10a00001;
      92209: inst = 32'hca06835;
      92210: inst = 32'h13e00001;
      92211: inst = 32'hfe0d96a;
      92212: inst = 32'h5be00000;
      92213: inst = 32'h8c50000;
      92214: inst = 32'h24612800;
      92215: inst = 32'h10a00000;
      92216: inst = 32'hca0000a;
      92217: inst = 32'h24822800;
      92218: inst = 32'h10a00000;
      92219: inst = 32'hca00004;
      92220: inst = 32'h38632800;
      92221: inst = 32'h38842800;
      92222: inst = 32'h10a00001;
      92223: inst = 32'hca06843;
      92224: inst = 32'h13e00001;
      92225: inst = 32'hfe0d96a;
      92226: inst = 32'h5be00000;
      92227: inst = 32'h8c50000;
      92228: inst = 32'h24612800;
      92229: inst = 32'h10a00000;
      92230: inst = 32'hca0000a;
      92231: inst = 32'h24822800;
      92232: inst = 32'h10a00000;
      92233: inst = 32'hca00004;
      92234: inst = 32'h38632800;
      92235: inst = 32'h38842800;
      92236: inst = 32'h10a00001;
      92237: inst = 32'hca06851;
      92238: inst = 32'h13e00001;
      92239: inst = 32'hfe0d96a;
      92240: inst = 32'h5be00000;
      92241: inst = 32'h8c50000;
      92242: inst = 32'h24612800;
      92243: inst = 32'h10a00000;
      92244: inst = 32'hca0000a;
      92245: inst = 32'h24822800;
      92246: inst = 32'h10a00000;
      92247: inst = 32'hca00004;
      92248: inst = 32'h38632800;
      92249: inst = 32'h38842800;
      92250: inst = 32'h10a00001;
      92251: inst = 32'hca0685f;
      92252: inst = 32'h13e00001;
      92253: inst = 32'hfe0d96a;
      92254: inst = 32'h5be00000;
      92255: inst = 32'h8c50000;
      92256: inst = 32'h24612800;
      92257: inst = 32'h10a00000;
      92258: inst = 32'hca0000a;
      92259: inst = 32'h24822800;
      92260: inst = 32'h10a00000;
      92261: inst = 32'hca00004;
      92262: inst = 32'h38632800;
      92263: inst = 32'h38842800;
      92264: inst = 32'h10a00001;
      92265: inst = 32'hca0686d;
      92266: inst = 32'h13e00001;
      92267: inst = 32'hfe0d96a;
      92268: inst = 32'h5be00000;
      92269: inst = 32'h8c50000;
      92270: inst = 32'h24612800;
      92271: inst = 32'h10a00000;
      92272: inst = 32'hca0000a;
      92273: inst = 32'h24822800;
      92274: inst = 32'h10a00000;
      92275: inst = 32'hca00004;
      92276: inst = 32'h38632800;
      92277: inst = 32'h38842800;
      92278: inst = 32'h10a00001;
      92279: inst = 32'hca0687b;
      92280: inst = 32'h13e00001;
      92281: inst = 32'hfe0d96a;
      92282: inst = 32'h5be00000;
      92283: inst = 32'h8c50000;
      92284: inst = 32'h24612800;
      92285: inst = 32'h10a00000;
      92286: inst = 32'hca0000a;
      92287: inst = 32'h24822800;
      92288: inst = 32'h10a00000;
      92289: inst = 32'hca00004;
      92290: inst = 32'h38632800;
      92291: inst = 32'h38842800;
      92292: inst = 32'h10a00001;
      92293: inst = 32'hca06889;
      92294: inst = 32'h13e00001;
      92295: inst = 32'hfe0d96a;
      92296: inst = 32'h5be00000;
      92297: inst = 32'h8c50000;
      92298: inst = 32'h24612800;
      92299: inst = 32'h10a00000;
      92300: inst = 32'hca0000a;
      92301: inst = 32'h24822800;
      92302: inst = 32'h10a00000;
      92303: inst = 32'hca00004;
      92304: inst = 32'h38632800;
      92305: inst = 32'h38842800;
      92306: inst = 32'h10a00001;
      92307: inst = 32'hca06897;
      92308: inst = 32'h13e00001;
      92309: inst = 32'hfe0d96a;
      92310: inst = 32'h5be00000;
      92311: inst = 32'h8c50000;
      92312: inst = 32'h24612800;
      92313: inst = 32'h10a00000;
      92314: inst = 32'hca0000a;
      92315: inst = 32'h24822800;
      92316: inst = 32'h10a00000;
      92317: inst = 32'hca00004;
      92318: inst = 32'h38632800;
      92319: inst = 32'h38842800;
      92320: inst = 32'h10a00001;
      92321: inst = 32'hca068a5;
      92322: inst = 32'h13e00001;
      92323: inst = 32'hfe0d96a;
      92324: inst = 32'h5be00000;
      92325: inst = 32'h8c50000;
      92326: inst = 32'h24612800;
      92327: inst = 32'h10a00000;
      92328: inst = 32'hca0000a;
      92329: inst = 32'h24822800;
      92330: inst = 32'h10a00000;
      92331: inst = 32'hca00004;
      92332: inst = 32'h38632800;
      92333: inst = 32'h38842800;
      92334: inst = 32'h10a00001;
      92335: inst = 32'hca068b3;
      92336: inst = 32'h13e00001;
      92337: inst = 32'hfe0d96a;
      92338: inst = 32'h5be00000;
      92339: inst = 32'h8c50000;
      92340: inst = 32'h24612800;
      92341: inst = 32'h10a00000;
      92342: inst = 32'hca0000a;
      92343: inst = 32'h24822800;
      92344: inst = 32'h10a00000;
      92345: inst = 32'hca00004;
      92346: inst = 32'h38632800;
      92347: inst = 32'h38842800;
      92348: inst = 32'h10a00001;
      92349: inst = 32'hca068c1;
      92350: inst = 32'h13e00001;
      92351: inst = 32'hfe0d96a;
      92352: inst = 32'h5be00000;
      92353: inst = 32'h8c50000;
      92354: inst = 32'h24612800;
      92355: inst = 32'h10a00000;
      92356: inst = 32'hca0000a;
      92357: inst = 32'h24822800;
      92358: inst = 32'h10a00000;
      92359: inst = 32'hca00004;
      92360: inst = 32'h38632800;
      92361: inst = 32'h38842800;
      92362: inst = 32'h10a00001;
      92363: inst = 32'hca068cf;
      92364: inst = 32'h13e00001;
      92365: inst = 32'hfe0d96a;
      92366: inst = 32'h5be00000;
      92367: inst = 32'h8c50000;
      92368: inst = 32'h24612800;
      92369: inst = 32'h10a00000;
      92370: inst = 32'hca0000a;
      92371: inst = 32'h24822800;
      92372: inst = 32'h10a00000;
      92373: inst = 32'hca00004;
      92374: inst = 32'h38632800;
      92375: inst = 32'h38842800;
      92376: inst = 32'h10a00001;
      92377: inst = 32'hca068dd;
      92378: inst = 32'h13e00001;
      92379: inst = 32'hfe0d96a;
      92380: inst = 32'h5be00000;
      92381: inst = 32'h8c50000;
      92382: inst = 32'h24612800;
      92383: inst = 32'h10a00000;
      92384: inst = 32'hca0000a;
      92385: inst = 32'h24822800;
      92386: inst = 32'h10a00000;
      92387: inst = 32'hca00004;
      92388: inst = 32'h38632800;
      92389: inst = 32'h38842800;
      92390: inst = 32'h10a00001;
      92391: inst = 32'hca068eb;
      92392: inst = 32'h13e00001;
      92393: inst = 32'hfe0d96a;
      92394: inst = 32'h5be00000;
      92395: inst = 32'h8c50000;
      92396: inst = 32'h24612800;
      92397: inst = 32'h10a00000;
      92398: inst = 32'hca0000a;
      92399: inst = 32'h24822800;
      92400: inst = 32'h10a00000;
      92401: inst = 32'hca00004;
      92402: inst = 32'h38632800;
      92403: inst = 32'h38842800;
      92404: inst = 32'h10a00001;
      92405: inst = 32'hca068f9;
      92406: inst = 32'h13e00001;
      92407: inst = 32'hfe0d96a;
      92408: inst = 32'h5be00000;
      92409: inst = 32'h8c50000;
      92410: inst = 32'h24612800;
      92411: inst = 32'h10a00000;
      92412: inst = 32'hca0000a;
      92413: inst = 32'h24822800;
      92414: inst = 32'h10a00000;
      92415: inst = 32'hca00004;
      92416: inst = 32'h38632800;
      92417: inst = 32'h38842800;
      92418: inst = 32'h10a00001;
      92419: inst = 32'hca06907;
      92420: inst = 32'h13e00001;
      92421: inst = 32'hfe0d96a;
      92422: inst = 32'h5be00000;
      92423: inst = 32'h8c50000;
      92424: inst = 32'h24612800;
      92425: inst = 32'h10a00000;
      92426: inst = 32'hca0000a;
      92427: inst = 32'h24822800;
      92428: inst = 32'h10a00000;
      92429: inst = 32'hca00004;
      92430: inst = 32'h38632800;
      92431: inst = 32'h38842800;
      92432: inst = 32'h10a00001;
      92433: inst = 32'hca06915;
      92434: inst = 32'h13e00001;
      92435: inst = 32'hfe0d96a;
      92436: inst = 32'h5be00000;
      92437: inst = 32'h8c50000;
      92438: inst = 32'h24612800;
      92439: inst = 32'h10a00000;
      92440: inst = 32'hca0000a;
      92441: inst = 32'h24822800;
      92442: inst = 32'h10a00000;
      92443: inst = 32'hca00004;
      92444: inst = 32'h38632800;
      92445: inst = 32'h38842800;
      92446: inst = 32'h10a00001;
      92447: inst = 32'hca06923;
      92448: inst = 32'h13e00001;
      92449: inst = 32'hfe0d96a;
      92450: inst = 32'h5be00000;
      92451: inst = 32'h8c50000;
      92452: inst = 32'h24612800;
      92453: inst = 32'h10a00000;
      92454: inst = 32'hca0000a;
      92455: inst = 32'h24822800;
      92456: inst = 32'h10a00000;
      92457: inst = 32'hca00004;
      92458: inst = 32'h38632800;
      92459: inst = 32'h38842800;
      92460: inst = 32'h10a00001;
      92461: inst = 32'hca06931;
      92462: inst = 32'h13e00001;
      92463: inst = 32'hfe0d96a;
      92464: inst = 32'h5be00000;
      92465: inst = 32'h8c50000;
      92466: inst = 32'h24612800;
      92467: inst = 32'h10a00000;
      92468: inst = 32'hca0000a;
      92469: inst = 32'h24822800;
      92470: inst = 32'h10a00000;
      92471: inst = 32'hca00004;
      92472: inst = 32'h38632800;
      92473: inst = 32'h38842800;
      92474: inst = 32'h10a00001;
      92475: inst = 32'hca0693f;
      92476: inst = 32'h13e00001;
      92477: inst = 32'hfe0d96a;
      92478: inst = 32'h5be00000;
      92479: inst = 32'h8c50000;
      92480: inst = 32'h24612800;
      92481: inst = 32'h10a00000;
      92482: inst = 32'hca0000a;
      92483: inst = 32'h24822800;
      92484: inst = 32'h10a00000;
      92485: inst = 32'hca00004;
      92486: inst = 32'h38632800;
      92487: inst = 32'h38842800;
      92488: inst = 32'h10a00001;
      92489: inst = 32'hca0694d;
      92490: inst = 32'h13e00001;
      92491: inst = 32'hfe0d96a;
      92492: inst = 32'h5be00000;
      92493: inst = 32'h8c50000;
      92494: inst = 32'h24612800;
      92495: inst = 32'h10a00000;
      92496: inst = 32'hca0000a;
      92497: inst = 32'h24822800;
      92498: inst = 32'h10a00000;
      92499: inst = 32'hca00004;
      92500: inst = 32'h38632800;
      92501: inst = 32'h38842800;
      92502: inst = 32'h10a00001;
      92503: inst = 32'hca0695b;
      92504: inst = 32'h13e00001;
      92505: inst = 32'hfe0d96a;
      92506: inst = 32'h5be00000;
      92507: inst = 32'h8c50000;
      92508: inst = 32'h24612800;
      92509: inst = 32'h10a00000;
      92510: inst = 32'hca0000a;
      92511: inst = 32'h24822800;
      92512: inst = 32'h10a00000;
      92513: inst = 32'hca00004;
      92514: inst = 32'h38632800;
      92515: inst = 32'h38842800;
      92516: inst = 32'h10a00001;
      92517: inst = 32'hca06969;
      92518: inst = 32'h13e00001;
      92519: inst = 32'hfe0d96a;
      92520: inst = 32'h5be00000;
      92521: inst = 32'h8c50000;
      92522: inst = 32'h24612800;
      92523: inst = 32'h10a00000;
      92524: inst = 32'hca0000a;
      92525: inst = 32'h24822800;
      92526: inst = 32'h10a00000;
      92527: inst = 32'hca00004;
      92528: inst = 32'h38632800;
      92529: inst = 32'h38842800;
      92530: inst = 32'h10a00001;
      92531: inst = 32'hca06977;
      92532: inst = 32'h13e00001;
      92533: inst = 32'hfe0d96a;
      92534: inst = 32'h5be00000;
      92535: inst = 32'h8c50000;
      92536: inst = 32'h24612800;
      92537: inst = 32'h10a00000;
      92538: inst = 32'hca0000a;
      92539: inst = 32'h24822800;
      92540: inst = 32'h10a00000;
      92541: inst = 32'hca00004;
      92542: inst = 32'h38632800;
      92543: inst = 32'h38842800;
      92544: inst = 32'h10a00001;
      92545: inst = 32'hca06985;
      92546: inst = 32'h13e00001;
      92547: inst = 32'hfe0d96a;
      92548: inst = 32'h5be00000;
      92549: inst = 32'h8c50000;
      92550: inst = 32'h24612800;
      92551: inst = 32'h10a00000;
      92552: inst = 32'hca0000a;
      92553: inst = 32'h24822800;
      92554: inst = 32'h10a00000;
      92555: inst = 32'hca00004;
      92556: inst = 32'h38632800;
      92557: inst = 32'h38842800;
      92558: inst = 32'h10a00001;
      92559: inst = 32'hca06993;
      92560: inst = 32'h13e00001;
      92561: inst = 32'hfe0d96a;
      92562: inst = 32'h5be00000;
      92563: inst = 32'h8c50000;
      92564: inst = 32'h24612800;
      92565: inst = 32'h10a00000;
      92566: inst = 32'hca0000a;
      92567: inst = 32'h24822800;
      92568: inst = 32'h10a00000;
      92569: inst = 32'hca00004;
      92570: inst = 32'h38632800;
      92571: inst = 32'h38842800;
      92572: inst = 32'h10a00001;
      92573: inst = 32'hca069a1;
      92574: inst = 32'h13e00001;
      92575: inst = 32'hfe0d96a;
      92576: inst = 32'h5be00000;
      92577: inst = 32'h8c50000;
      92578: inst = 32'h24612800;
      92579: inst = 32'h10a00000;
      92580: inst = 32'hca0000a;
      92581: inst = 32'h24822800;
      92582: inst = 32'h10a00000;
      92583: inst = 32'hca00004;
      92584: inst = 32'h38632800;
      92585: inst = 32'h38842800;
      92586: inst = 32'h10a00001;
      92587: inst = 32'hca069af;
      92588: inst = 32'h13e00001;
      92589: inst = 32'hfe0d96a;
      92590: inst = 32'h5be00000;
      92591: inst = 32'h8c50000;
      92592: inst = 32'h24612800;
      92593: inst = 32'h10a00000;
      92594: inst = 32'hca0000a;
      92595: inst = 32'h24822800;
      92596: inst = 32'h10a00000;
      92597: inst = 32'hca00004;
      92598: inst = 32'h38632800;
      92599: inst = 32'h38842800;
      92600: inst = 32'h10a00001;
      92601: inst = 32'hca069bd;
      92602: inst = 32'h13e00001;
      92603: inst = 32'hfe0d96a;
      92604: inst = 32'h5be00000;
      92605: inst = 32'h8c50000;
      92606: inst = 32'h24612800;
      92607: inst = 32'h10a00000;
      92608: inst = 32'hca0000a;
      92609: inst = 32'h24822800;
      92610: inst = 32'h10a00000;
      92611: inst = 32'hca00004;
      92612: inst = 32'h38632800;
      92613: inst = 32'h38842800;
      92614: inst = 32'h10a00001;
      92615: inst = 32'hca069cb;
      92616: inst = 32'h13e00001;
      92617: inst = 32'hfe0d96a;
      92618: inst = 32'h5be00000;
      92619: inst = 32'h8c50000;
      92620: inst = 32'h24612800;
      92621: inst = 32'h10a00000;
      92622: inst = 32'hca0000a;
      92623: inst = 32'h24822800;
      92624: inst = 32'h10a00000;
      92625: inst = 32'hca00004;
      92626: inst = 32'h38632800;
      92627: inst = 32'h38842800;
      92628: inst = 32'h10a00001;
      92629: inst = 32'hca069d9;
      92630: inst = 32'h13e00001;
      92631: inst = 32'hfe0d96a;
      92632: inst = 32'h5be00000;
      92633: inst = 32'h8c50000;
      92634: inst = 32'h24612800;
      92635: inst = 32'h10a00000;
      92636: inst = 32'hca0000a;
      92637: inst = 32'h24822800;
      92638: inst = 32'h10a00000;
      92639: inst = 32'hca00004;
      92640: inst = 32'h38632800;
      92641: inst = 32'h38842800;
      92642: inst = 32'h10a00001;
      92643: inst = 32'hca069e7;
      92644: inst = 32'h13e00001;
      92645: inst = 32'hfe0d96a;
      92646: inst = 32'h5be00000;
      92647: inst = 32'h8c50000;
      92648: inst = 32'h24612800;
      92649: inst = 32'h10a00000;
      92650: inst = 32'hca0000a;
      92651: inst = 32'h24822800;
      92652: inst = 32'h10a00000;
      92653: inst = 32'hca00004;
      92654: inst = 32'h38632800;
      92655: inst = 32'h38842800;
      92656: inst = 32'h10a00001;
      92657: inst = 32'hca069f5;
      92658: inst = 32'h13e00001;
      92659: inst = 32'hfe0d96a;
      92660: inst = 32'h5be00000;
      92661: inst = 32'h8c50000;
      92662: inst = 32'h24612800;
      92663: inst = 32'h10a00000;
      92664: inst = 32'hca0000a;
      92665: inst = 32'h24822800;
      92666: inst = 32'h10a00000;
      92667: inst = 32'hca00004;
      92668: inst = 32'h38632800;
      92669: inst = 32'h38842800;
      92670: inst = 32'h10a00001;
      92671: inst = 32'hca06a03;
      92672: inst = 32'h13e00001;
      92673: inst = 32'hfe0d96a;
      92674: inst = 32'h5be00000;
      92675: inst = 32'h8c50000;
      92676: inst = 32'h24612800;
      92677: inst = 32'h10a00000;
      92678: inst = 32'hca0000a;
      92679: inst = 32'h24822800;
      92680: inst = 32'h10a00000;
      92681: inst = 32'hca00004;
      92682: inst = 32'h38632800;
      92683: inst = 32'h38842800;
      92684: inst = 32'h10a00001;
      92685: inst = 32'hca06a11;
      92686: inst = 32'h13e00001;
      92687: inst = 32'hfe0d96a;
      92688: inst = 32'h5be00000;
      92689: inst = 32'h8c50000;
      92690: inst = 32'h24612800;
      92691: inst = 32'h10a00000;
      92692: inst = 32'hca0000a;
      92693: inst = 32'h24822800;
      92694: inst = 32'h10a00000;
      92695: inst = 32'hca00004;
      92696: inst = 32'h38632800;
      92697: inst = 32'h38842800;
      92698: inst = 32'h10a00001;
      92699: inst = 32'hca06a1f;
      92700: inst = 32'h13e00001;
      92701: inst = 32'hfe0d96a;
      92702: inst = 32'h5be00000;
      92703: inst = 32'h8c50000;
      92704: inst = 32'h24612800;
      92705: inst = 32'h10a00000;
      92706: inst = 32'hca0000a;
      92707: inst = 32'h24822800;
      92708: inst = 32'h10a00000;
      92709: inst = 32'hca00004;
      92710: inst = 32'h38632800;
      92711: inst = 32'h38842800;
      92712: inst = 32'h10a00001;
      92713: inst = 32'hca06a2d;
      92714: inst = 32'h13e00001;
      92715: inst = 32'hfe0d96a;
      92716: inst = 32'h5be00000;
      92717: inst = 32'h8c50000;
      92718: inst = 32'h24612800;
      92719: inst = 32'h10a00000;
      92720: inst = 32'hca0000a;
      92721: inst = 32'h24822800;
      92722: inst = 32'h10a00000;
      92723: inst = 32'hca00004;
      92724: inst = 32'h38632800;
      92725: inst = 32'h38842800;
      92726: inst = 32'h10a00001;
      92727: inst = 32'hca06a3b;
      92728: inst = 32'h13e00001;
      92729: inst = 32'hfe0d96a;
      92730: inst = 32'h5be00000;
      92731: inst = 32'h8c50000;
      92732: inst = 32'h24612800;
      92733: inst = 32'h10a00000;
      92734: inst = 32'hca0000a;
      92735: inst = 32'h24822800;
      92736: inst = 32'h10a00000;
      92737: inst = 32'hca00004;
      92738: inst = 32'h38632800;
      92739: inst = 32'h38842800;
      92740: inst = 32'h10a00001;
      92741: inst = 32'hca06a49;
      92742: inst = 32'h13e00001;
      92743: inst = 32'hfe0d96a;
      92744: inst = 32'h5be00000;
      92745: inst = 32'h8c50000;
      92746: inst = 32'h24612800;
      92747: inst = 32'h10a00000;
      92748: inst = 32'hca0000a;
      92749: inst = 32'h24822800;
      92750: inst = 32'h10a00000;
      92751: inst = 32'hca00004;
      92752: inst = 32'h38632800;
      92753: inst = 32'h38842800;
      92754: inst = 32'h10a00001;
      92755: inst = 32'hca06a57;
      92756: inst = 32'h13e00001;
      92757: inst = 32'hfe0d96a;
      92758: inst = 32'h5be00000;
      92759: inst = 32'h8c50000;
      92760: inst = 32'h24612800;
      92761: inst = 32'h10a00000;
      92762: inst = 32'hca0000a;
      92763: inst = 32'h24822800;
      92764: inst = 32'h10a00000;
      92765: inst = 32'hca00004;
      92766: inst = 32'h38632800;
      92767: inst = 32'h38842800;
      92768: inst = 32'h10a00001;
      92769: inst = 32'hca06a65;
      92770: inst = 32'h13e00001;
      92771: inst = 32'hfe0d96a;
      92772: inst = 32'h5be00000;
      92773: inst = 32'h8c50000;
      92774: inst = 32'h24612800;
      92775: inst = 32'h10a00000;
      92776: inst = 32'hca0000a;
      92777: inst = 32'h24822800;
      92778: inst = 32'h10a00000;
      92779: inst = 32'hca00004;
      92780: inst = 32'h38632800;
      92781: inst = 32'h38842800;
      92782: inst = 32'h10a00001;
      92783: inst = 32'hca06a73;
      92784: inst = 32'h13e00001;
      92785: inst = 32'hfe0d96a;
      92786: inst = 32'h5be00000;
      92787: inst = 32'h8c50000;
      92788: inst = 32'h24612800;
      92789: inst = 32'h10a00000;
      92790: inst = 32'hca0000a;
      92791: inst = 32'h24822800;
      92792: inst = 32'h10a00000;
      92793: inst = 32'hca00004;
      92794: inst = 32'h38632800;
      92795: inst = 32'h38842800;
      92796: inst = 32'h10a00001;
      92797: inst = 32'hca06a81;
      92798: inst = 32'h13e00001;
      92799: inst = 32'hfe0d96a;
      92800: inst = 32'h5be00000;
      92801: inst = 32'h8c50000;
      92802: inst = 32'h24612800;
      92803: inst = 32'h10a00000;
      92804: inst = 32'hca0000a;
      92805: inst = 32'h24822800;
      92806: inst = 32'h10a00000;
      92807: inst = 32'hca00004;
      92808: inst = 32'h38632800;
      92809: inst = 32'h38842800;
      92810: inst = 32'h10a00001;
      92811: inst = 32'hca06a8f;
      92812: inst = 32'h13e00001;
      92813: inst = 32'hfe0d96a;
      92814: inst = 32'h5be00000;
      92815: inst = 32'h8c50000;
      92816: inst = 32'h24612800;
      92817: inst = 32'h10a00000;
      92818: inst = 32'hca0000a;
      92819: inst = 32'h24822800;
      92820: inst = 32'h10a00000;
      92821: inst = 32'hca00004;
      92822: inst = 32'h38632800;
      92823: inst = 32'h38842800;
      92824: inst = 32'h10a00001;
      92825: inst = 32'hca06a9d;
      92826: inst = 32'h13e00001;
      92827: inst = 32'hfe0d96a;
      92828: inst = 32'h5be00000;
      92829: inst = 32'h8c50000;
      92830: inst = 32'h24612800;
      92831: inst = 32'h10a00000;
      92832: inst = 32'hca0000a;
      92833: inst = 32'h24822800;
      92834: inst = 32'h10a00000;
      92835: inst = 32'hca00004;
      92836: inst = 32'h38632800;
      92837: inst = 32'h38842800;
      92838: inst = 32'h10a00001;
      92839: inst = 32'hca06aab;
      92840: inst = 32'h13e00001;
      92841: inst = 32'hfe0d96a;
      92842: inst = 32'h5be00000;
      92843: inst = 32'h8c50000;
      92844: inst = 32'h24612800;
      92845: inst = 32'h10a00000;
      92846: inst = 32'hca0000a;
      92847: inst = 32'h24822800;
      92848: inst = 32'h10a00000;
      92849: inst = 32'hca00004;
      92850: inst = 32'h38632800;
      92851: inst = 32'h38842800;
      92852: inst = 32'h10a00001;
      92853: inst = 32'hca06ab9;
      92854: inst = 32'h13e00001;
      92855: inst = 32'hfe0d96a;
      92856: inst = 32'h5be00000;
      92857: inst = 32'h8c50000;
      92858: inst = 32'h24612800;
      92859: inst = 32'h10a00000;
      92860: inst = 32'hca0000a;
      92861: inst = 32'h24822800;
      92862: inst = 32'h10a00000;
      92863: inst = 32'hca00004;
      92864: inst = 32'h38632800;
      92865: inst = 32'h38842800;
      92866: inst = 32'h10a00001;
      92867: inst = 32'hca06ac7;
      92868: inst = 32'h13e00001;
      92869: inst = 32'hfe0d96a;
      92870: inst = 32'h5be00000;
      92871: inst = 32'h8c50000;
      92872: inst = 32'h24612800;
      92873: inst = 32'h10a00000;
      92874: inst = 32'hca0000a;
      92875: inst = 32'h24822800;
      92876: inst = 32'h10a00000;
      92877: inst = 32'hca00004;
      92878: inst = 32'h38632800;
      92879: inst = 32'h38842800;
      92880: inst = 32'h10a00001;
      92881: inst = 32'hca06ad5;
      92882: inst = 32'h13e00001;
      92883: inst = 32'hfe0d96a;
      92884: inst = 32'h5be00000;
      92885: inst = 32'h8c50000;
      92886: inst = 32'h24612800;
      92887: inst = 32'h10a00000;
      92888: inst = 32'hca0000a;
      92889: inst = 32'h24822800;
      92890: inst = 32'h10a00000;
      92891: inst = 32'hca00004;
      92892: inst = 32'h38632800;
      92893: inst = 32'h38842800;
      92894: inst = 32'h10a00001;
      92895: inst = 32'hca06ae3;
      92896: inst = 32'h13e00001;
      92897: inst = 32'hfe0d96a;
      92898: inst = 32'h5be00000;
      92899: inst = 32'h8c50000;
      92900: inst = 32'h24612800;
      92901: inst = 32'h10a00000;
      92902: inst = 32'hca0000a;
      92903: inst = 32'h24822800;
      92904: inst = 32'h10a00000;
      92905: inst = 32'hca00004;
      92906: inst = 32'h38632800;
      92907: inst = 32'h38842800;
      92908: inst = 32'h10a00001;
      92909: inst = 32'hca06af1;
      92910: inst = 32'h13e00001;
      92911: inst = 32'hfe0d96a;
      92912: inst = 32'h5be00000;
      92913: inst = 32'h8c50000;
      92914: inst = 32'h24612800;
      92915: inst = 32'h10a00000;
      92916: inst = 32'hca0000a;
      92917: inst = 32'h24822800;
      92918: inst = 32'h10a00000;
      92919: inst = 32'hca00004;
      92920: inst = 32'h38632800;
      92921: inst = 32'h38842800;
      92922: inst = 32'h10a00001;
      92923: inst = 32'hca06aff;
      92924: inst = 32'h13e00001;
      92925: inst = 32'hfe0d96a;
      92926: inst = 32'h5be00000;
      92927: inst = 32'h8c50000;
      92928: inst = 32'h24612800;
      92929: inst = 32'h10a00000;
      92930: inst = 32'hca0000a;
      92931: inst = 32'h24822800;
      92932: inst = 32'h10a00000;
      92933: inst = 32'hca00004;
      92934: inst = 32'h38632800;
      92935: inst = 32'h38842800;
      92936: inst = 32'h10a00001;
      92937: inst = 32'hca06b0d;
      92938: inst = 32'h13e00001;
      92939: inst = 32'hfe0d96a;
      92940: inst = 32'h5be00000;
      92941: inst = 32'h8c50000;
      92942: inst = 32'h24612800;
      92943: inst = 32'h10a00000;
      92944: inst = 32'hca0000a;
      92945: inst = 32'h24822800;
      92946: inst = 32'h10a00000;
      92947: inst = 32'hca00004;
      92948: inst = 32'h38632800;
      92949: inst = 32'h38842800;
      92950: inst = 32'h10a00001;
      92951: inst = 32'hca06b1b;
      92952: inst = 32'h13e00001;
      92953: inst = 32'hfe0d96a;
      92954: inst = 32'h5be00000;
      92955: inst = 32'h8c50000;
      92956: inst = 32'h24612800;
      92957: inst = 32'h10a00000;
      92958: inst = 32'hca0000a;
      92959: inst = 32'h24822800;
      92960: inst = 32'h10a00000;
      92961: inst = 32'hca00004;
      92962: inst = 32'h38632800;
      92963: inst = 32'h38842800;
      92964: inst = 32'h10a00001;
      92965: inst = 32'hca06b29;
      92966: inst = 32'h13e00001;
      92967: inst = 32'hfe0d96a;
      92968: inst = 32'h5be00000;
      92969: inst = 32'h8c50000;
      92970: inst = 32'h24612800;
      92971: inst = 32'h10a00000;
      92972: inst = 32'hca0000b;
      92973: inst = 32'h24822800;
      92974: inst = 32'h10a00000;
      92975: inst = 32'hca00004;
      92976: inst = 32'h38632800;
      92977: inst = 32'h38842800;
      92978: inst = 32'h10a00001;
      92979: inst = 32'hca06b37;
      92980: inst = 32'h13e00001;
      92981: inst = 32'hfe0d96a;
      92982: inst = 32'h5be00000;
      92983: inst = 32'h8c50000;
      92984: inst = 32'h24612800;
      92985: inst = 32'h10a00000;
      92986: inst = 32'hca0000b;
      92987: inst = 32'h24822800;
      92988: inst = 32'h10a00000;
      92989: inst = 32'hca00004;
      92990: inst = 32'h38632800;
      92991: inst = 32'h38842800;
      92992: inst = 32'h10a00001;
      92993: inst = 32'hca06b45;
      92994: inst = 32'h13e00001;
      92995: inst = 32'hfe0d96a;
      92996: inst = 32'h5be00000;
      92997: inst = 32'h8c50000;
      92998: inst = 32'h24612800;
      92999: inst = 32'h10a00000;
      93000: inst = 32'hca0000b;
      93001: inst = 32'h24822800;
      93002: inst = 32'h10a00000;
      93003: inst = 32'hca00004;
      93004: inst = 32'h38632800;
      93005: inst = 32'h38842800;
      93006: inst = 32'h10a00001;
      93007: inst = 32'hca06b53;
      93008: inst = 32'h13e00001;
      93009: inst = 32'hfe0d96a;
      93010: inst = 32'h5be00000;
      93011: inst = 32'h8c50000;
      93012: inst = 32'h24612800;
      93013: inst = 32'h10a00000;
      93014: inst = 32'hca0000b;
      93015: inst = 32'h24822800;
      93016: inst = 32'h10a00000;
      93017: inst = 32'hca00004;
      93018: inst = 32'h38632800;
      93019: inst = 32'h38842800;
      93020: inst = 32'h10a00001;
      93021: inst = 32'hca06b61;
      93022: inst = 32'h13e00001;
      93023: inst = 32'hfe0d96a;
      93024: inst = 32'h5be00000;
      93025: inst = 32'h8c50000;
      93026: inst = 32'h24612800;
      93027: inst = 32'h10a00000;
      93028: inst = 32'hca0000b;
      93029: inst = 32'h24822800;
      93030: inst = 32'h10a00000;
      93031: inst = 32'hca00004;
      93032: inst = 32'h38632800;
      93033: inst = 32'h38842800;
      93034: inst = 32'h10a00001;
      93035: inst = 32'hca06b6f;
      93036: inst = 32'h13e00001;
      93037: inst = 32'hfe0d96a;
      93038: inst = 32'h5be00000;
      93039: inst = 32'h8c50000;
      93040: inst = 32'h24612800;
      93041: inst = 32'h10a00000;
      93042: inst = 32'hca0000b;
      93043: inst = 32'h24822800;
      93044: inst = 32'h10a00000;
      93045: inst = 32'hca00004;
      93046: inst = 32'h38632800;
      93047: inst = 32'h38842800;
      93048: inst = 32'h10a00001;
      93049: inst = 32'hca06b7d;
      93050: inst = 32'h13e00001;
      93051: inst = 32'hfe0d96a;
      93052: inst = 32'h5be00000;
      93053: inst = 32'h8c50000;
      93054: inst = 32'h24612800;
      93055: inst = 32'h10a00000;
      93056: inst = 32'hca0000b;
      93057: inst = 32'h24822800;
      93058: inst = 32'h10a00000;
      93059: inst = 32'hca00004;
      93060: inst = 32'h38632800;
      93061: inst = 32'h38842800;
      93062: inst = 32'h10a00001;
      93063: inst = 32'hca06b8b;
      93064: inst = 32'h13e00001;
      93065: inst = 32'hfe0d96a;
      93066: inst = 32'h5be00000;
      93067: inst = 32'h8c50000;
      93068: inst = 32'h24612800;
      93069: inst = 32'h10a00000;
      93070: inst = 32'hca0000b;
      93071: inst = 32'h24822800;
      93072: inst = 32'h10a00000;
      93073: inst = 32'hca00004;
      93074: inst = 32'h38632800;
      93075: inst = 32'h38842800;
      93076: inst = 32'h10a00001;
      93077: inst = 32'hca06b99;
      93078: inst = 32'h13e00001;
      93079: inst = 32'hfe0d96a;
      93080: inst = 32'h5be00000;
      93081: inst = 32'h8c50000;
      93082: inst = 32'h24612800;
      93083: inst = 32'h10a00000;
      93084: inst = 32'hca0000b;
      93085: inst = 32'h24822800;
      93086: inst = 32'h10a00000;
      93087: inst = 32'hca00004;
      93088: inst = 32'h38632800;
      93089: inst = 32'h38842800;
      93090: inst = 32'h10a00001;
      93091: inst = 32'hca06ba7;
      93092: inst = 32'h13e00001;
      93093: inst = 32'hfe0d96a;
      93094: inst = 32'h5be00000;
      93095: inst = 32'h8c50000;
      93096: inst = 32'h24612800;
      93097: inst = 32'h10a00000;
      93098: inst = 32'hca0000b;
      93099: inst = 32'h24822800;
      93100: inst = 32'h10a00000;
      93101: inst = 32'hca00004;
      93102: inst = 32'h38632800;
      93103: inst = 32'h38842800;
      93104: inst = 32'h10a00001;
      93105: inst = 32'hca06bb5;
      93106: inst = 32'h13e00001;
      93107: inst = 32'hfe0d96a;
      93108: inst = 32'h5be00000;
      93109: inst = 32'h8c50000;
      93110: inst = 32'h24612800;
      93111: inst = 32'h10a00000;
      93112: inst = 32'hca0000b;
      93113: inst = 32'h24822800;
      93114: inst = 32'h10a00000;
      93115: inst = 32'hca00004;
      93116: inst = 32'h38632800;
      93117: inst = 32'h38842800;
      93118: inst = 32'h10a00001;
      93119: inst = 32'hca06bc3;
      93120: inst = 32'h13e00001;
      93121: inst = 32'hfe0d96a;
      93122: inst = 32'h5be00000;
      93123: inst = 32'h8c50000;
      93124: inst = 32'h24612800;
      93125: inst = 32'h10a00000;
      93126: inst = 32'hca0000b;
      93127: inst = 32'h24822800;
      93128: inst = 32'h10a00000;
      93129: inst = 32'hca00004;
      93130: inst = 32'h38632800;
      93131: inst = 32'h38842800;
      93132: inst = 32'h10a00001;
      93133: inst = 32'hca06bd1;
      93134: inst = 32'h13e00001;
      93135: inst = 32'hfe0d96a;
      93136: inst = 32'h5be00000;
      93137: inst = 32'h8c50000;
      93138: inst = 32'h24612800;
      93139: inst = 32'h10a00000;
      93140: inst = 32'hca0000b;
      93141: inst = 32'h24822800;
      93142: inst = 32'h10a00000;
      93143: inst = 32'hca00004;
      93144: inst = 32'h38632800;
      93145: inst = 32'h38842800;
      93146: inst = 32'h10a00001;
      93147: inst = 32'hca06bdf;
      93148: inst = 32'h13e00001;
      93149: inst = 32'hfe0d96a;
      93150: inst = 32'h5be00000;
      93151: inst = 32'h8c50000;
      93152: inst = 32'h24612800;
      93153: inst = 32'h10a00000;
      93154: inst = 32'hca0000b;
      93155: inst = 32'h24822800;
      93156: inst = 32'h10a00000;
      93157: inst = 32'hca00004;
      93158: inst = 32'h38632800;
      93159: inst = 32'h38842800;
      93160: inst = 32'h10a00001;
      93161: inst = 32'hca06bed;
      93162: inst = 32'h13e00001;
      93163: inst = 32'hfe0d96a;
      93164: inst = 32'h5be00000;
      93165: inst = 32'h8c50000;
      93166: inst = 32'h24612800;
      93167: inst = 32'h10a00000;
      93168: inst = 32'hca0000b;
      93169: inst = 32'h24822800;
      93170: inst = 32'h10a00000;
      93171: inst = 32'hca00004;
      93172: inst = 32'h38632800;
      93173: inst = 32'h38842800;
      93174: inst = 32'h10a00001;
      93175: inst = 32'hca06bfb;
      93176: inst = 32'h13e00001;
      93177: inst = 32'hfe0d96a;
      93178: inst = 32'h5be00000;
      93179: inst = 32'h8c50000;
      93180: inst = 32'h24612800;
      93181: inst = 32'h10a00000;
      93182: inst = 32'hca0000b;
      93183: inst = 32'h24822800;
      93184: inst = 32'h10a00000;
      93185: inst = 32'hca00004;
      93186: inst = 32'h38632800;
      93187: inst = 32'h38842800;
      93188: inst = 32'h10a00001;
      93189: inst = 32'hca06c09;
      93190: inst = 32'h13e00001;
      93191: inst = 32'hfe0d96a;
      93192: inst = 32'h5be00000;
      93193: inst = 32'h8c50000;
      93194: inst = 32'h24612800;
      93195: inst = 32'h10a00000;
      93196: inst = 32'hca0000b;
      93197: inst = 32'h24822800;
      93198: inst = 32'h10a00000;
      93199: inst = 32'hca00004;
      93200: inst = 32'h38632800;
      93201: inst = 32'h38842800;
      93202: inst = 32'h10a00001;
      93203: inst = 32'hca06c17;
      93204: inst = 32'h13e00001;
      93205: inst = 32'hfe0d96a;
      93206: inst = 32'h5be00000;
      93207: inst = 32'h8c50000;
      93208: inst = 32'h24612800;
      93209: inst = 32'h10a00000;
      93210: inst = 32'hca0000b;
      93211: inst = 32'h24822800;
      93212: inst = 32'h10a00000;
      93213: inst = 32'hca00004;
      93214: inst = 32'h38632800;
      93215: inst = 32'h38842800;
      93216: inst = 32'h10a00001;
      93217: inst = 32'hca06c25;
      93218: inst = 32'h13e00001;
      93219: inst = 32'hfe0d96a;
      93220: inst = 32'h5be00000;
      93221: inst = 32'h8c50000;
      93222: inst = 32'h24612800;
      93223: inst = 32'h10a00000;
      93224: inst = 32'hca0000b;
      93225: inst = 32'h24822800;
      93226: inst = 32'h10a00000;
      93227: inst = 32'hca00004;
      93228: inst = 32'h38632800;
      93229: inst = 32'h38842800;
      93230: inst = 32'h10a00001;
      93231: inst = 32'hca06c33;
      93232: inst = 32'h13e00001;
      93233: inst = 32'hfe0d96a;
      93234: inst = 32'h5be00000;
      93235: inst = 32'h8c50000;
      93236: inst = 32'h24612800;
      93237: inst = 32'h10a00000;
      93238: inst = 32'hca0000b;
      93239: inst = 32'h24822800;
      93240: inst = 32'h10a00000;
      93241: inst = 32'hca00004;
      93242: inst = 32'h38632800;
      93243: inst = 32'h38842800;
      93244: inst = 32'h10a00001;
      93245: inst = 32'hca06c41;
      93246: inst = 32'h13e00001;
      93247: inst = 32'hfe0d96a;
      93248: inst = 32'h5be00000;
      93249: inst = 32'h8c50000;
      93250: inst = 32'h24612800;
      93251: inst = 32'h10a00000;
      93252: inst = 32'hca0000b;
      93253: inst = 32'h24822800;
      93254: inst = 32'h10a00000;
      93255: inst = 32'hca00004;
      93256: inst = 32'h38632800;
      93257: inst = 32'h38842800;
      93258: inst = 32'h10a00001;
      93259: inst = 32'hca06c4f;
      93260: inst = 32'h13e00001;
      93261: inst = 32'hfe0d96a;
      93262: inst = 32'h5be00000;
      93263: inst = 32'h8c50000;
      93264: inst = 32'h24612800;
      93265: inst = 32'h10a00000;
      93266: inst = 32'hca0000b;
      93267: inst = 32'h24822800;
      93268: inst = 32'h10a00000;
      93269: inst = 32'hca00004;
      93270: inst = 32'h38632800;
      93271: inst = 32'h38842800;
      93272: inst = 32'h10a00001;
      93273: inst = 32'hca06c5d;
      93274: inst = 32'h13e00001;
      93275: inst = 32'hfe0d96a;
      93276: inst = 32'h5be00000;
      93277: inst = 32'h8c50000;
      93278: inst = 32'h24612800;
      93279: inst = 32'h10a00000;
      93280: inst = 32'hca0000b;
      93281: inst = 32'h24822800;
      93282: inst = 32'h10a00000;
      93283: inst = 32'hca00004;
      93284: inst = 32'h38632800;
      93285: inst = 32'h38842800;
      93286: inst = 32'h10a00001;
      93287: inst = 32'hca06c6b;
      93288: inst = 32'h13e00001;
      93289: inst = 32'hfe0d96a;
      93290: inst = 32'h5be00000;
      93291: inst = 32'h8c50000;
      93292: inst = 32'h24612800;
      93293: inst = 32'h10a00000;
      93294: inst = 32'hca0000b;
      93295: inst = 32'h24822800;
      93296: inst = 32'h10a00000;
      93297: inst = 32'hca00004;
      93298: inst = 32'h38632800;
      93299: inst = 32'h38842800;
      93300: inst = 32'h10a00001;
      93301: inst = 32'hca06c79;
      93302: inst = 32'h13e00001;
      93303: inst = 32'hfe0d96a;
      93304: inst = 32'h5be00000;
      93305: inst = 32'h8c50000;
      93306: inst = 32'h24612800;
      93307: inst = 32'h10a00000;
      93308: inst = 32'hca0000b;
      93309: inst = 32'h24822800;
      93310: inst = 32'h10a00000;
      93311: inst = 32'hca00004;
      93312: inst = 32'h38632800;
      93313: inst = 32'h38842800;
      93314: inst = 32'h10a00001;
      93315: inst = 32'hca06c87;
      93316: inst = 32'h13e00001;
      93317: inst = 32'hfe0d96a;
      93318: inst = 32'h5be00000;
      93319: inst = 32'h8c50000;
      93320: inst = 32'h24612800;
      93321: inst = 32'h10a00000;
      93322: inst = 32'hca0000b;
      93323: inst = 32'h24822800;
      93324: inst = 32'h10a00000;
      93325: inst = 32'hca00004;
      93326: inst = 32'h38632800;
      93327: inst = 32'h38842800;
      93328: inst = 32'h10a00001;
      93329: inst = 32'hca06c95;
      93330: inst = 32'h13e00001;
      93331: inst = 32'hfe0d96a;
      93332: inst = 32'h5be00000;
      93333: inst = 32'h8c50000;
      93334: inst = 32'h24612800;
      93335: inst = 32'h10a00000;
      93336: inst = 32'hca0000b;
      93337: inst = 32'h24822800;
      93338: inst = 32'h10a00000;
      93339: inst = 32'hca00004;
      93340: inst = 32'h38632800;
      93341: inst = 32'h38842800;
      93342: inst = 32'h10a00001;
      93343: inst = 32'hca06ca3;
      93344: inst = 32'h13e00001;
      93345: inst = 32'hfe0d96a;
      93346: inst = 32'h5be00000;
      93347: inst = 32'h8c50000;
      93348: inst = 32'h24612800;
      93349: inst = 32'h10a00000;
      93350: inst = 32'hca0000b;
      93351: inst = 32'h24822800;
      93352: inst = 32'h10a00000;
      93353: inst = 32'hca00004;
      93354: inst = 32'h38632800;
      93355: inst = 32'h38842800;
      93356: inst = 32'h10a00001;
      93357: inst = 32'hca06cb1;
      93358: inst = 32'h13e00001;
      93359: inst = 32'hfe0d96a;
      93360: inst = 32'h5be00000;
      93361: inst = 32'h8c50000;
      93362: inst = 32'h24612800;
      93363: inst = 32'h10a00000;
      93364: inst = 32'hca0000b;
      93365: inst = 32'h24822800;
      93366: inst = 32'h10a00000;
      93367: inst = 32'hca00004;
      93368: inst = 32'h38632800;
      93369: inst = 32'h38842800;
      93370: inst = 32'h10a00001;
      93371: inst = 32'hca06cbf;
      93372: inst = 32'h13e00001;
      93373: inst = 32'hfe0d96a;
      93374: inst = 32'h5be00000;
      93375: inst = 32'h8c50000;
      93376: inst = 32'h24612800;
      93377: inst = 32'h10a00000;
      93378: inst = 32'hca0000b;
      93379: inst = 32'h24822800;
      93380: inst = 32'h10a00000;
      93381: inst = 32'hca00004;
      93382: inst = 32'h38632800;
      93383: inst = 32'h38842800;
      93384: inst = 32'h10a00001;
      93385: inst = 32'hca06ccd;
      93386: inst = 32'h13e00001;
      93387: inst = 32'hfe0d96a;
      93388: inst = 32'h5be00000;
      93389: inst = 32'h8c50000;
      93390: inst = 32'h24612800;
      93391: inst = 32'h10a00000;
      93392: inst = 32'hca0000b;
      93393: inst = 32'h24822800;
      93394: inst = 32'h10a00000;
      93395: inst = 32'hca00004;
      93396: inst = 32'h38632800;
      93397: inst = 32'h38842800;
      93398: inst = 32'h10a00001;
      93399: inst = 32'hca06cdb;
      93400: inst = 32'h13e00001;
      93401: inst = 32'hfe0d96a;
      93402: inst = 32'h5be00000;
      93403: inst = 32'h8c50000;
      93404: inst = 32'h24612800;
      93405: inst = 32'h10a00000;
      93406: inst = 32'hca0000b;
      93407: inst = 32'h24822800;
      93408: inst = 32'h10a00000;
      93409: inst = 32'hca00004;
      93410: inst = 32'h38632800;
      93411: inst = 32'h38842800;
      93412: inst = 32'h10a00001;
      93413: inst = 32'hca06ce9;
      93414: inst = 32'h13e00001;
      93415: inst = 32'hfe0d96a;
      93416: inst = 32'h5be00000;
      93417: inst = 32'h8c50000;
      93418: inst = 32'h24612800;
      93419: inst = 32'h10a00000;
      93420: inst = 32'hca0000b;
      93421: inst = 32'h24822800;
      93422: inst = 32'h10a00000;
      93423: inst = 32'hca00004;
      93424: inst = 32'h38632800;
      93425: inst = 32'h38842800;
      93426: inst = 32'h10a00001;
      93427: inst = 32'hca06cf7;
      93428: inst = 32'h13e00001;
      93429: inst = 32'hfe0d96a;
      93430: inst = 32'h5be00000;
      93431: inst = 32'h8c50000;
      93432: inst = 32'h24612800;
      93433: inst = 32'h10a00000;
      93434: inst = 32'hca0000b;
      93435: inst = 32'h24822800;
      93436: inst = 32'h10a00000;
      93437: inst = 32'hca00004;
      93438: inst = 32'h38632800;
      93439: inst = 32'h38842800;
      93440: inst = 32'h10a00001;
      93441: inst = 32'hca06d05;
      93442: inst = 32'h13e00001;
      93443: inst = 32'hfe0d96a;
      93444: inst = 32'h5be00000;
      93445: inst = 32'h8c50000;
      93446: inst = 32'h24612800;
      93447: inst = 32'h10a00000;
      93448: inst = 32'hca0000b;
      93449: inst = 32'h24822800;
      93450: inst = 32'h10a00000;
      93451: inst = 32'hca00004;
      93452: inst = 32'h38632800;
      93453: inst = 32'h38842800;
      93454: inst = 32'h10a00001;
      93455: inst = 32'hca06d13;
      93456: inst = 32'h13e00001;
      93457: inst = 32'hfe0d96a;
      93458: inst = 32'h5be00000;
      93459: inst = 32'h8c50000;
      93460: inst = 32'h24612800;
      93461: inst = 32'h10a00000;
      93462: inst = 32'hca0000b;
      93463: inst = 32'h24822800;
      93464: inst = 32'h10a00000;
      93465: inst = 32'hca00004;
      93466: inst = 32'h38632800;
      93467: inst = 32'h38842800;
      93468: inst = 32'h10a00001;
      93469: inst = 32'hca06d21;
      93470: inst = 32'h13e00001;
      93471: inst = 32'hfe0d96a;
      93472: inst = 32'h5be00000;
      93473: inst = 32'h8c50000;
      93474: inst = 32'h24612800;
      93475: inst = 32'h10a00000;
      93476: inst = 32'hca0000b;
      93477: inst = 32'h24822800;
      93478: inst = 32'h10a00000;
      93479: inst = 32'hca00004;
      93480: inst = 32'h38632800;
      93481: inst = 32'h38842800;
      93482: inst = 32'h10a00001;
      93483: inst = 32'hca06d2f;
      93484: inst = 32'h13e00001;
      93485: inst = 32'hfe0d96a;
      93486: inst = 32'h5be00000;
      93487: inst = 32'h8c50000;
      93488: inst = 32'h24612800;
      93489: inst = 32'h10a00000;
      93490: inst = 32'hca0000b;
      93491: inst = 32'h24822800;
      93492: inst = 32'h10a00000;
      93493: inst = 32'hca00004;
      93494: inst = 32'h38632800;
      93495: inst = 32'h38842800;
      93496: inst = 32'h10a00001;
      93497: inst = 32'hca06d3d;
      93498: inst = 32'h13e00001;
      93499: inst = 32'hfe0d96a;
      93500: inst = 32'h5be00000;
      93501: inst = 32'h8c50000;
      93502: inst = 32'h24612800;
      93503: inst = 32'h10a00000;
      93504: inst = 32'hca0000b;
      93505: inst = 32'h24822800;
      93506: inst = 32'h10a00000;
      93507: inst = 32'hca00004;
      93508: inst = 32'h38632800;
      93509: inst = 32'h38842800;
      93510: inst = 32'h10a00001;
      93511: inst = 32'hca06d4b;
      93512: inst = 32'h13e00001;
      93513: inst = 32'hfe0d96a;
      93514: inst = 32'h5be00000;
      93515: inst = 32'h8c50000;
      93516: inst = 32'h24612800;
      93517: inst = 32'h10a00000;
      93518: inst = 32'hca0000b;
      93519: inst = 32'h24822800;
      93520: inst = 32'h10a00000;
      93521: inst = 32'hca00004;
      93522: inst = 32'h38632800;
      93523: inst = 32'h38842800;
      93524: inst = 32'h10a00001;
      93525: inst = 32'hca06d59;
      93526: inst = 32'h13e00001;
      93527: inst = 32'hfe0d96a;
      93528: inst = 32'h5be00000;
      93529: inst = 32'h8c50000;
      93530: inst = 32'h24612800;
      93531: inst = 32'h10a00000;
      93532: inst = 32'hca0000b;
      93533: inst = 32'h24822800;
      93534: inst = 32'h10a00000;
      93535: inst = 32'hca00004;
      93536: inst = 32'h38632800;
      93537: inst = 32'h38842800;
      93538: inst = 32'h10a00001;
      93539: inst = 32'hca06d67;
      93540: inst = 32'h13e00001;
      93541: inst = 32'hfe0d96a;
      93542: inst = 32'h5be00000;
      93543: inst = 32'h8c50000;
      93544: inst = 32'h24612800;
      93545: inst = 32'h10a00000;
      93546: inst = 32'hca0000b;
      93547: inst = 32'h24822800;
      93548: inst = 32'h10a00000;
      93549: inst = 32'hca00004;
      93550: inst = 32'h38632800;
      93551: inst = 32'h38842800;
      93552: inst = 32'h10a00001;
      93553: inst = 32'hca06d75;
      93554: inst = 32'h13e00001;
      93555: inst = 32'hfe0d96a;
      93556: inst = 32'h5be00000;
      93557: inst = 32'h8c50000;
      93558: inst = 32'h24612800;
      93559: inst = 32'h10a00000;
      93560: inst = 32'hca0000b;
      93561: inst = 32'h24822800;
      93562: inst = 32'h10a00000;
      93563: inst = 32'hca00004;
      93564: inst = 32'h38632800;
      93565: inst = 32'h38842800;
      93566: inst = 32'h10a00001;
      93567: inst = 32'hca06d83;
      93568: inst = 32'h13e00001;
      93569: inst = 32'hfe0d96a;
      93570: inst = 32'h5be00000;
      93571: inst = 32'h8c50000;
      93572: inst = 32'h24612800;
      93573: inst = 32'h10a00000;
      93574: inst = 32'hca0000b;
      93575: inst = 32'h24822800;
      93576: inst = 32'h10a00000;
      93577: inst = 32'hca00004;
      93578: inst = 32'h38632800;
      93579: inst = 32'h38842800;
      93580: inst = 32'h10a00001;
      93581: inst = 32'hca06d91;
      93582: inst = 32'h13e00001;
      93583: inst = 32'hfe0d96a;
      93584: inst = 32'h5be00000;
      93585: inst = 32'h8c50000;
      93586: inst = 32'h24612800;
      93587: inst = 32'h10a00000;
      93588: inst = 32'hca0000b;
      93589: inst = 32'h24822800;
      93590: inst = 32'h10a00000;
      93591: inst = 32'hca00004;
      93592: inst = 32'h38632800;
      93593: inst = 32'h38842800;
      93594: inst = 32'h10a00001;
      93595: inst = 32'hca06d9f;
      93596: inst = 32'h13e00001;
      93597: inst = 32'hfe0d96a;
      93598: inst = 32'h5be00000;
      93599: inst = 32'h8c50000;
      93600: inst = 32'h24612800;
      93601: inst = 32'h10a00000;
      93602: inst = 32'hca0000b;
      93603: inst = 32'h24822800;
      93604: inst = 32'h10a00000;
      93605: inst = 32'hca00004;
      93606: inst = 32'h38632800;
      93607: inst = 32'h38842800;
      93608: inst = 32'h10a00001;
      93609: inst = 32'hca06dad;
      93610: inst = 32'h13e00001;
      93611: inst = 32'hfe0d96a;
      93612: inst = 32'h5be00000;
      93613: inst = 32'h8c50000;
      93614: inst = 32'h24612800;
      93615: inst = 32'h10a00000;
      93616: inst = 32'hca0000b;
      93617: inst = 32'h24822800;
      93618: inst = 32'h10a00000;
      93619: inst = 32'hca00004;
      93620: inst = 32'h38632800;
      93621: inst = 32'h38842800;
      93622: inst = 32'h10a00001;
      93623: inst = 32'hca06dbb;
      93624: inst = 32'h13e00001;
      93625: inst = 32'hfe0d96a;
      93626: inst = 32'h5be00000;
      93627: inst = 32'h8c50000;
      93628: inst = 32'h24612800;
      93629: inst = 32'h10a00000;
      93630: inst = 32'hca0000b;
      93631: inst = 32'h24822800;
      93632: inst = 32'h10a00000;
      93633: inst = 32'hca00004;
      93634: inst = 32'h38632800;
      93635: inst = 32'h38842800;
      93636: inst = 32'h10a00001;
      93637: inst = 32'hca06dc9;
      93638: inst = 32'h13e00001;
      93639: inst = 32'hfe0d96a;
      93640: inst = 32'h5be00000;
      93641: inst = 32'h8c50000;
      93642: inst = 32'h24612800;
      93643: inst = 32'h10a00000;
      93644: inst = 32'hca0000b;
      93645: inst = 32'h24822800;
      93646: inst = 32'h10a00000;
      93647: inst = 32'hca00004;
      93648: inst = 32'h38632800;
      93649: inst = 32'h38842800;
      93650: inst = 32'h10a00001;
      93651: inst = 32'hca06dd7;
      93652: inst = 32'h13e00001;
      93653: inst = 32'hfe0d96a;
      93654: inst = 32'h5be00000;
      93655: inst = 32'h8c50000;
      93656: inst = 32'h24612800;
      93657: inst = 32'h10a00000;
      93658: inst = 32'hca0000b;
      93659: inst = 32'h24822800;
      93660: inst = 32'h10a00000;
      93661: inst = 32'hca00004;
      93662: inst = 32'h38632800;
      93663: inst = 32'h38842800;
      93664: inst = 32'h10a00001;
      93665: inst = 32'hca06de5;
      93666: inst = 32'h13e00001;
      93667: inst = 32'hfe0d96a;
      93668: inst = 32'h5be00000;
      93669: inst = 32'h8c50000;
      93670: inst = 32'h24612800;
      93671: inst = 32'h10a00000;
      93672: inst = 32'hca0000b;
      93673: inst = 32'h24822800;
      93674: inst = 32'h10a00000;
      93675: inst = 32'hca00004;
      93676: inst = 32'h38632800;
      93677: inst = 32'h38842800;
      93678: inst = 32'h10a00001;
      93679: inst = 32'hca06df3;
      93680: inst = 32'h13e00001;
      93681: inst = 32'hfe0d96a;
      93682: inst = 32'h5be00000;
      93683: inst = 32'h8c50000;
      93684: inst = 32'h24612800;
      93685: inst = 32'h10a00000;
      93686: inst = 32'hca0000b;
      93687: inst = 32'h24822800;
      93688: inst = 32'h10a00000;
      93689: inst = 32'hca00004;
      93690: inst = 32'h38632800;
      93691: inst = 32'h38842800;
      93692: inst = 32'h10a00001;
      93693: inst = 32'hca06e01;
      93694: inst = 32'h13e00001;
      93695: inst = 32'hfe0d96a;
      93696: inst = 32'h5be00000;
      93697: inst = 32'h8c50000;
      93698: inst = 32'h24612800;
      93699: inst = 32'h10a00000;
      93700: inst = 32'hca0000b;
      93701: inst = 32'h24822800;
      93702: inst = 32'h10a00000;
      93703: inst = 32'hca00004;
      93704: inst = 32'h38632800;
      93705: inst = 32'h38842800;
      93706: inst = 32'h10a00001;
      93707: inst = 32'hca06e0f;
      93708: inst = 32'h13e00001;
      93709: inst = 32'hfe0d96a;
      93710: inst = 32'h5be00000;
      93711: inst = 32'h8c50000;
      93712: inst = 32'h24612800;
      93713: inst = 32'h10a00000;
      93714: inst = 32'hca0000b;
      93715: inst = 32'h24822800;
      93716: inst = 32'h10a00000;
      93717: inst = 32'hca00004;
      93718: inst = 32'h38632800;
      93719: inst = 32'h38842800;
      93720: inst = 32'h10a00001;
      93721: inst = 32'hca06e1d;
      93722: inst = 32'h13e00001;
      93723: inst = 32'hfe0d96a;
      93724: inst = 32'h5be00000;
      93725: inst = 32'h8c50000;
      93726: inst = 32'h24612800;
      93727: inst = 32'h10a00000;
      93728: inst = 32'hca0000b;
      93729: inst = 32'h24822800;
      93730: inst = 32'h10a00000;
      93731: inst = 32'hca00004;
      93732: inst = 32'h38632800;
      93733: inst = 32'h38842800;
      93734: inst = 32'h10a00001;
      93735: inst = 32'hca06e2b;
      93736: inst = 32'h13e00001;
      93737: inst = 32'hfe0d96a;
      93738: inst = 32'h5be00000;
      93739: inst = 32'h8c50000;
      93740: inst = 32'h24612800;
      93741: inst = 32'h10a00000;
      93742: inst = 32'hca0000b;
      93743: inst = 32'h24822800;
      93744: inst = 32'h10a00000;
      93745: inst = 32'hca00004;
      93746: inst = 32'h38632800;
      93747: inst = 32'h38842800;
      93748: inst = 32'h10a00001;
      93749: inst = 32'hca06e39;
      93750: inst = 32'h13e00001;
      93751: inst = 32'hfe0d96a;
      93752: inst = 32'h5be00000;
      93753: inst = 32'h8c50000;
      93754: inst = 32'h24612800;
      93755: inst = 32'h10a00000;
      93756: inst = 32'hca0000b;
      93757: inst = 32'h24822800;
      93758: inst = 32'h10a00000;
      93759: inst = 32'hca00004;
      93760: inst = 32'h38632800;
      93761: inst = 32'h38842800;
      93762: inst = 32'h10a00001;
      93763: inst = 32'hca06e47;
      93764: inst = 32'h13e00001;
      93765: inst = 32'hfe0d96a;
      93766: inst = 32'h5be00000;
      93767: inst = 32'h8c50000;
      93768: inst = 32'h24612800;
      93769: inst = 32'h10a00000;
      93770: inst = 32'hca0000b;
      93771: inst = 32'h24822800;
      93772: inst = 32'h10a00000;
      93773: inst = 32'hca00004;
      93774: inst = 32'h38632800;
      93775: inst = 32'h38842800;
      93776: inst = 32'h10a00001;
      93777: inst = 32'hca06e55;
      93778: inst = 32'h13e00001;
      93779: inst = 32'hfe0d96a;
      93780: inst = 32'h5be00000;
      93781: inst = 32'h8c50000;
      93782: inst = 32'h24612800;
      93783: inst = 32'h10a00000;
      93784: inst = 32'hca0000b;
      93785: inst = 32'h24822800;
      93786: inst = 32'h10a00000;
      93787: inst = 32'hca00004;
      93788: inst = 32'h38632800;
      93789: inst = 32'h38842800;
      93790: inst = 32'h10a00001;
      93791: inst = 32'hca06e63;
      93792: inst = 32'h13e00001;
      93793: inst = 32'hfe0d96a;
      93794: inst = 32'h5be00000;
      93795: inst = 32'h8c50000;
      93796: inst = 32'h24612800;
      93797: inst = 32'h10a00000;
      93798: inst = 32'hca0000b;
      93799: inst = 32'h24822800;
      93800: inst = 32'h10a00000;
      93801: inst = 32'hca00004;
      93802: inst = 32'h38632800;
      93803: inst = 32'h38842800;
      93804: inst = 32'h10a00001;
      93805: inst = 32'hca06e71;
      93806: inst = 32'h13e00001;
      93807: inst = 32'hfe0d96a;
      93808: inst = 32'h5be00000;
      93809: inst = 32'h8c50000;
      93810: inst = 32'h24612800;
      93811: inst = 32'h10a00000;
      93812: inst = 32'hca0000b;
      93813: inst = 32'h24822800;
      93814: inst = 32'h10a00000;
      93815: inst = 32'hca00004;
      93816: inst = 32'h38632800;
      93817: inst = 32'h38842800;
      93818: inst = 32'h10a00001;
      93819: inst = 32'hca06e7f;
      93820: inst = 32'h13e00001;
      93821: inst = 32'hfe0d96a;
      93822: inst = 32'h5be00000;
      93823: inst = 32'h8c50000;
      93824: inst = 32'h24612800;
      93825: inst = 32'h10a00000;
      93826: inst = 32'hca0000b;
      93827: inst = 32'h24822800;
      93828: inst = 32'h10a00000;
      93829: inst = 32'hca00004;
      93830: inst = 32'h38632800;
      93831: inst = 32'h38842800;
      93832: inst = 32'h10a00001;
      93833: inst = 32'hca06e8d;
      93834: inst = 32'h13e00001;
      93835: inst = 32'hfe0d96a;
      93836: inst = 32'h5be00000;
      93837: inst = 32'h8c50000;
      93838: inst = 32'h24612800;
      93839: inst = 32'h10a00000;
      93840: inst = 32'hca0000b;
      93841: inst = 32'h24822800;
      93842: inst = 32'h10a00000;
      93843: inst = 32'hca00004;
      93844: inst = 32'h38632800;
      93845: inst = 32'h38842800;
      93846: inst = 32'h10a00001;
      93847: inst = 32'hca06e9b;
      93848: inst = 32'h13e00001;
      93849: inst = 32'hfe0d96a;
      93850: inst = 32'h5be00000;
      93851: inst = 32'h8c50000;
      93852: inst = 32'h24612800;
      93853: inst = 32'h10a00000;
      93854: inst = 32'hca0000b;
      93855: inst = 32'h24822800;
      93856: inst = 32'h10a00000;
      93857: inst = 32'hca00004;
      93858: inst = 32'h38632800;
      93859: inst = 32'h38842800;
      93860: inst = 32'h10a00001;
      93861: inst = 32'hca06ea9;
      93862: inst = 32'h13e00001;
      93863: inst = 32'hfe0d96a;
      93864: inst = 32'h5be00000;
      93865: inst = 32'h8c50000;
      93866: inst = 32'h24612800;
      93867: inst = 32'h10a00000;
      93868: inst = 32'hca0000b;
      93869: inst = 32'h24822800;
      93870: inst = 32'h10a00000;
      93871: inst = 32'hca00004;
      93872: inst = 32'h38632800;
      93873: inst = 32'h38842800;
      93874: inst = 32'h10a00001;
      93875: inst = 32'hca06eb7;
      93876: inst = 32'h13e00001;
      93877: inst = 32'hfe0d96a;
      93878: inst = 32'h5be00000;
      93879: inst = 32'h8c50000;
      93880: inst = 32'h24612800;
      93881: inst = 32'h10a00000;
      93882: inst = 32'hca0000b;
      93883: inst = 32'h24822800;
      93884: inst = 32'h10a00000;
      93885: inst = 32'hca00004;
      93886: inst = 32'h38632800;
      93887: inst = 32'h38842800;
      93888: inst = 32'h10a00001;
      93889: inst = 32'hca06ec5;
      93890: inst = 32'h13e00001;
      93891: inst = 32'hfe0d96a;
      93892: inst = 32'h5be00000;
      93893: inst = 32'h8c50000;
      93894: inst = 32'h24612800;
      93895: inst = 32'h10a00000;
      93896: inst = 32'hca0000b;
      93897: inst = 32'h24822800;
      93898: inst = 32'h10a00000;
      93899: inst = 32'hca00004;
      93900: inst = 32'h38632800;
      93901: inst = 32'h38842800;
      93902: inst = 32'h10a00001;
      93903: inst = 32'hca06ed3;
      93904: inst = 32'h13e00001;
      93905: inst = 32'hfe0d96a;
      93906: inst = 32'h5be00000;
      93907: inst = 32'h8c50000;
      93908: inst = 32'h24612800;
      93909: inst = 32'h10a00000;
      93910: inst = 32'hca0000b;
      93911: inst = 32'h24822800;
      93912: inst = 32'h10a00000;
      93913: inst = 32'hca00004;
      93914: inst = 32'h38632800;
      93915: inst = 32'h38842800;
      93916: inst = 32'h10a00001;
      93917: inst = 32'hca06ee1;
      93918: inst = 32'h13e00001;
      93919: inst = 32'hfe0d96a;
      93920: inst = 32'h5be00000;
      93921: inst = 32'h8c50000;
      93922: inst = 32'h24612800;
      93923: inst = 32'h10a00000;
      93924: inst = 32'hca0000b;
      93925: inst = 32'h24822800;
      93926: inst = 32'h10a00000;
      93927: inst = 32'hca00004;
      93928: inst = 32'h38632800;
      93929: inst = 32'h38842800;
      93930: inst = 32'h10a00001;
      93931: inst = 32'hca06eef;
      93932: inst = 32'h13e00001;
      93933: inst = 32'hfe0d96a;
      93934: inst = 32'h5be00000;
      93935: inst = 32'h8c50000;
      93936: inst = 32'h24612800;
      93937: inst = 32'h10a00000;
      93938: inst = 32'hca0000b;
      93939: inst = 32'h24822800;
      93940: inst = 32'h10a00000;
      93941: inst = 32'hca00004;
      93942: inst = 32'h38632800;
      93943: inst = 32'h38842800;
      93944: inst = 32'h10a00001;
      93945: inst = 32'hca06efd;
      93946: inst = 32'h13e00001;
      93947: inst = 32'hfe0d96a;
      93948: inst = 32'h5be00000;
      93949: inst = 32'h8c50000;
      93950: inst = 32'h24612800;
      93951: inst = 32'h10a00000;
      93952: inst = 32'hca0000b;
      93953: inst = 32'h24822800;
      93954: inst = 32'h10a00000;
      93955: inst = 32'hca00004;
      93956: inst = 32'h38632800;
      93957: inst = 32'h38842800;
      93958: inst = 32'h10a00001;
      93959: inst = 32'hca06f0b;
      93960: inst = 32'h13e00001;
      93961: inst = 32'hfe0d96a;
      93962: inst = 32'h5be00000;
      93963: inst = 32'h8c50000;
      93964: inst = 32'h24612800;
      93965: inst = 32'h10a00000;
      93966: inst = 32'hca0000b;
      93967: inst = 32'h24822800;
      93968: inst = 32'h10a00000;
      93969: inst = 32'hca00004;
      93970: inst = 32'h38632800;
      93971: inst = 32'h38842800;
      93972: inst = 32'h10a00001;
      93973: inst = 32'hca06f19;
      93974: inst = 32'h13e00001;
      93975: inst = 32'hfe0d96a;
      93976: inst = 32'h5be00000;
      93977: inst = 32'h8c50000;
      93978: inst = 32'h24612800;
      93979: inst = 32'h10a00000;
      93980: inst = 32'hca0000b;
      93981: inst = 32'h24822800;
      93982: inst = 32'h10a00000;
      93983: inst = 32'hca00004;
      93984: inst = 32'h38632800;
      93985: inst = 32'h38842800;
      93986: inst = 32'h10a00001;
      93987: inst = 32'hca06f27;
      93988: inst = 32'h13e00001;
      93989: inst = 32'hfe0d96a;
      93990: inst = 32'h5be00000;
      93991: inst = 32'h8c50000;
      93992: inst = 32'h24612800;
      93993: inst = 32'h10a00000;
      93994: inst = 32'hca0000b;
      93995: inst = 32'h24822800;
      93996: inst = 32'h10a00000;
      93997: inst = 32'hca00004;
      93998: inst = 32'h38632800;
      93999: inst = 32'h38842800;
      94000: inst = 32'h10a00001;
      94001: inst = 32'hca06f35;
      94002: inst = 32'h13e00001;
      94003: inst = 32'hfe0d96a;
      94004: inst = 32'h5be00000;
      94005: inst = 32'h8c50000;
      94006: inst = 32'h24612800;
      94007: inst = 32'h10a00000;
      94008: inst = 32'hca0000b;
      94009: inst = 32'h24822800;
      94010: inst = 32'h10a00000;
      94011: inst = 32'hca00004;
      94012: inst = 32'h38632800;
      94013: inst = 32'h38842800;
      94014: inst = 32'h10a00001;
      94015: inst = 32'hca06f43;
      94016: inst = 32'h13e00001;
      94017: inst = 32'hfe0d96a;
      94018: inst = 32'h5be00000;
      94019: inst = 32'h8c50000;
      94020: inst = 32'h24612800;
      94021: inst = 32'h10a00000;
      94022: inst = 32'hca0000b;
      94023: inst = 32'h24822800;
      94024: inst = 32'h10a00000;
      94025: inst = 32'hca00004;
      94026: inst = 32'h38632800;
      94027: inst = 32'h38842800;
      94028: inst = 32'h10a00001;
      94029: inst = 32'hca06f51;
      94030: inst = 32'h13e00001;
      94031: inst = 32'hfe0d96a;
      94032: inst = 32'h5be00000;
      94033: inst = 32'h8c50000;
      94034: inst = 32'h24612800;
      94035: inst = 32'h10a00000;
      94036: inst = 32'hca0000b;
      94037: inst = 32'h24822800;
      94038: inst = 32'h10a00000;
      94039: inst = 32'hca00004;
      94040: inst = 32'h38632800;
      94041: inst = 32'h38842800;
      94042: inst = 32'h10a00001;
      94043: inst = 32'hca06f5f;
      94044: inst = 32'h13e00001;
      94045: inst = 32'hfe0d96a;
      94046: inst = 32'h5be00000;
      94047: inst = 32'h8c50000;
      94048: inst = 32'h24612800;
      94049: inst = 32'h10a00000;
      94050: inst = 32'hca0000b;
      94051: inst = 32'h24822800;
      94052: inst = 32'h10a00000;
      94053: inst = 32'hca00004;
      94054: inst = 32'h38632800;
      94055: inst = 32'h38842800;
      94056: inst = 32'h10a00001;
      94057: inst = 32'hca06f6d;
      94058: inst = 32'h13e00001;
      94059: inst = 32'hfe0d96a;
      94060: inst = 32'h5be00000;
      94061: inst = 32'h8c50000;
      94062: inst = 32'h24612800;
      94063: inst = 32'h10a00000;
      94064: inst = 32'hca0000b;
      94065: inst = 32'h24822800;
      94066: inst = 32'h10a00000;
      94067: inst = 32'hca00004;
      94068: inst = 32'h38632800;
      94069: inst = 32'h38842800;
      94070: inst = 32'h10a00001;
      94071: inst = 32'hca06f7b;
      94072: inst = 32'h13e00001;
      94073: inst = 32'hfe0d96a;
      94074: inst = 32'h5be00000;
      94075: inst = 32'h8c50000;
      94076: inst = 32'h24612800;
      94077: inst = 32'h10a00000;
      94078: inst = 32'hca0000b;
      94079: inst = 32'h24822800;
      94080: inst = 32'h10a00000;
      94081: inst = 32'hca00004;
      94082: inst = 32'h38632800;
      94083: inst = 32'h38842800;
      94084: inst = 32'h10a00001;
      94085: inst = 32'hca06f89;
      94086: inst = 32'h13e00001;
      94087: inst = 32'hfe0d96a;
      94088: inst = 32'h5be00000;
      94089: inst = 32'h8c50000;
      94090: inst = 32'h24612800;
      94091: inst = 32'h10a00000;
      94092: inst = 32'hca0000b;
      94093: inst = 32'h24822800;
      94094: inst = 32'h10a00000;
      94095: inst = 32'hca00004;
      94096: inst = 32'h38632800;
      94097: inst = 32'h38842800;
      94098: inst = 32'h10a00001;
      94099: inst = 32'hca06f97;
      94100: inst = 32'h13e00001;
      94101: inst = 32'hfe0d96a;
      94102: inst = 32'h5be00000;
      94103: inst = 32'h8c50000;
      94104: inst = 32'h24612800;
      94105: inst = 32'h10a00000;
      94106: inst = 32'hca0000b;
      94107: inst = 32'h24822800;
      94108: inst = 32'h10a00000;
      94109: inst = 32'hca00004;
      94110: inst = 32'h38632800;
      94111: inst = 32'h38842800;
      94112: inst = 32'h10a00001;
      94113: inst = 32'hca06fa5;
      94114: inst = 32'h13e00001;
      94115: inst = 32'hfe0d96a;
      94116: inst = 32'h5be00000;
      94117: inst = 32'h8c50000;
      94118: inst = 32'h24612800;
      94119: inst = 32'h10a00000;
      94120: inst = 32'hca0000b;
      94121: inst = 32'h24822800;
      94122: inst = 32'h10a00000;
      94123: inst = 32'hca00004;
      94124: inst = 32'h38632800;
      94125: inst = 32'h38842800;
      94126: inst = 32'h10a00001;
      94127: inst = 32'hca06fb3;
      94128: inst = 32'h13e00001;
      94129: inst = 32'hfe0d96a;
      94130: inst = 32'h5be00000;
      94131: inst = 32'h8c50000;
      94132: inst = 32'h24612800;
      94133: inst = 32'h10a00000;
      94134: inst = 32'hca0000b;
      94135: inst = 32'h24822800;
      94136: inst = 32'h10a00000;
      94137: inst = 32'hca00004;
      94138: inst = 32'h38632800;
      94139: inst = 32'h38842800;
      94140: inst = 32'h10a00001;
      94141: inst = 32'hca06fc1;
      94142: inst = 32'h13e00001;
      94143: inst = 32'hfe0d96a;
      94144: inst = 32'h5be00000;
      94145: inst = 32'h8c50000;
      94146: inst = 32'h24612800;
      94147: inst = 32'h10a00000;
      94148: inst = 32'hca0000b;
      94149: inst = 32'h24822800;
      94150: inst = 32'h10a00000;
      94151: inst = 32'hca00004;
      94152: inst = 32'h38632800;
      94153: inst = 32'h38842800;
      94154: inst = 32'h10a00001;
      94155: inst = 32'hca06fcf;
      94156: inst = 32'h13e00001;
      94157: inst = 32'hfe0d96a;
      94158: inst = 32'h5be00000;
      94159: inst = 32'h8c50000;
      94160: inst = 32'h24612800;
      94161: inst = 32'h10a00000;
      94162: inst = 32'hca0000b;
      94163: inst = 32'h24822800;
      94164: inst = 32'h10a00000;
      94165: inst = 32'hca00004;
      94166: inst = 32'h38632800;
      94167: inst = 32'h38842800;
      94168: inst = 32'h10a00001;
      94169: inst = 32'hca06fdd;
      94170: inst = 32'h13e00001;
      94171: inst = 32'hfe0d96a;
      94172: inst = 32'h5be00000;
      94173: inst = 32'h8c50000;
      94174: inst = 32'h24612800;
      94175: inst = 32'h10a00000;
      94176: inst = 32'hca0000b;
      94177: inst = 32'h24822800;
      94178: inst = 32'h10a00000;
      94179: inst = 32'hca00004;
      94180: inst = 32'h38632800;
      94181: inst = 32'h38842800;
      94182: inst = 32'h10a00001;
      94183: inst = 32'hca06feb;
      94184: inst = 32'h13e00001;
      94185: inst = 32'hfe0d96a;
      94186: inst = 32'h5be00000;
      94187: inst = 32'h8c50000;
      94188: inst = 32'h24612800;
      94189: inst = 32'h10a00000;
      94190: inst = 32'hca0000b;
      94191: inst = 32'h24822800;
      94192: inst = 32'h10a00000;
      94193: inst = 32'hca00004;
      94194: inst = 32'h38632800;
      94195: inst = 32'h38842800;
      94196: inst = 32'h10a00001;
      94197: inst = 32'hca06ff9;
      94198: inst = 32'h13e00001;
      94199: inst = 32'hfe0d96a;
      94200: inst = 32'h5be00000;
      94201: inst = 32'h8c50000;
      94202: inst = 32'h24612800;
      94203: inst = 32'h10a00000;
      94204: inst = 32'hca0000b;
      94205: inst = 32'h24822800;
      94206: inst = 32'h10a00000;
      94207: inst = 32'hca00004;
      94208: inst = 32'h38632800;
      94209: inst = 32'h38842800;
      94210: inst = 32'h10a00001;
      94211: inst = 32'hca07007;
      94212: inst = 32'h13e00001;
      94213: inst = 32'hfe0d96a;
      94214: inst = 32'h5be00000;
      94215: inst = 32'h8c50000;
      94216: inst = 32'h24612800;
      94217: inst = 32'h10a00000;
      94218: inst = 32'hca0000b;
      94219: inst = 32'h24822800;
      94220: inst = 32'h10a00000;
      94221: inst = 32'hca00004;
      94222: inst = 32'h38632800;
      94223: inst = 32'h38842800;
      94224: inst = 32'h10a00001;
      94225: inst = 32'hca07015;
      94226: inst = 32'h13e00001;
      94227: inst = 32'hfe0d96a;
      94228: inst = 32'h5be00000;
      94229: inst = 32'h8c50000;
      94230: inst = 32'h24612800;
      94231: inst = 32'h10a00000;
      94232: inst = 32'hca0000b;
      94233: inst = 32'h24822800;
      94234: inst = 32'h10a00000;
      94235: inst = 32'hca00004;
      94236: inst = 32'h38632800;
      94237: inst = 32'h38842800;
      94238: inst = 32'h10a00001;
      94239: inst = 32'hca07023;
      94240: inst = 32'h13e00001;
      94241: inst = 32'hfe0d96a;
      94242: inst = 32'h5be00000;
      94243: inst = 32'h8c50000;
      94244: inst = 32'h24612800;
      94245: inst = 32'h10a00000;
      94246: inst = 32'hca0000b;
      94247: inst = 32'h24822800;
      94248: inst = 32'h10a00000;
      94249: inst = 32'hca00004;
      94250: inst = 32'h38632800;
      94251: inst = 32'h38842800;
      94252: inst = 32'h10a00001;
      94253: inst = 32'hca07031;
      94254: inst = 32'h13e00001;
      94255: inst = 32'hfe0d96a;
      94256: inst = 32'h5be00000;
      94257: inst = 32'h8c50000;
      94258: inst = 32'h24612800;
      94259: inst = 32'h10a00000;
      94260: inst = 32'hca0000b;
      94261: inst = 32'h24822800;
      94262: inst = 32'h10a00000;
      94263: inst = 32'hca00004;
      94264: inst = 32'h38632800;
      94265: inst = 32'h38842800;
      94266: inst = 32'h10a00001;
      94267: inst = 32'hca0703f;
      94268: inst = 32'h13e00001;
      94269: inst = 32'hfe0d96a;
      94270: inst = 32'h5be00000;
      94271: inst = 32'h8c50000;
      94272: inst = 32'h24612800;
      94273: inst = 32'h10a00000;
      94274: inst = 32'hca0000b;
      94275: inst = 32'h24822800;
      94276: inst = 32'h10a00000;
      94277: inst = 32'hca00004;
      94278: inst = 32'h38632800;
      94279: inst = 32'h38842800;
      94280: inst = 32'h10a00001;
      94281: inst = 32'hca0704d;
      94282: inst = 32'h13e00001;
      94283: inst = 32'hfe0d96a;
      94284: inst = 32'h5be00000;
      94285: inst = 32'h8c50000;
      94286: inst = 32'h24612800;
      94287: inst = 32'h10a00000;
      94288: inst = 32'hca0000b;
      94289: inst = 32'h24822800;
      94290: inst = 32'h10a00000;
      94291: inst = 32'hca00004;
      94292: inst = 32'h38632800;
      94293: inst = 32'h38842800;
      94294: inst = 32'h10a00001;
      94295: inst = 32'hca0705b;
      94296: inst = 32'h13e00001;
      94297: inst = 32'hfe0d96a;
      94298: inst = 32'h5be00000;
      94299: inst = 32'h8c50000;
      94300: inst = 32'h24612800;
      94301: inst = 32'h10a00000;
      94302: inst = 32'hca0000b;
      94303: inst = 32'h24822800;
      94304: inst = 32'h10a00000;
      94305: inst = 32'hca00004;
      94306: inst = 32'h38632800;
      94307: inst = 32'h38842800;
      94308: inst = 32'h10a00001;
      94309: inst = 32'hca07069;
      94310: inst = 32'h13e00001;
      94311: inst = 32'hfe0d96a;
      94312: inst = 32'h5be00000;
      94313: inst = 32'h8c50000;
      94314: inst = 32'h24612800;
      94315: inst = 32'h10a00000;
      94316: inst = 32'hca0000c;
      94317: inst = 32'h24822800;
      94318: inst = 32'h10a00000;
      94319: inst = 32'hca00004;
      94320: inst = 32'h38632800;
      94321: inst = 32'h38842800;
      94322: inst = 32'h10a00001;
      94323: inst = 32'hca07077;
      94324: inst = 32'h13e00001;
      94325: inst = 32'hfe0d96a;
      94326: inst = 32'h5be00000;
      94327: inst = 32'h8c50000;
      94328: inst = 32'h24612800;
      94329: inst = 32'h10a00000;
      94330: inst = 32'hca0000c;
      94331: inst = 32'h24822800;
      94332: inst = 32'h10a00000;
      94333: inst = 32'hca00004;
      94334: inst = 32'h38632800;
      94335: inst = 32'h38842800;
      94336: inst = 32'h10a00001;
      94337: inst = 32'hca07085;
      94338: inst = 32'h13e00001;
      94339: inst = 32'hfe0d96a;
      94340: inst = 32'h5be00000;
      94341: inst = 32'h8c50000;
      94342: inst = 32'h24612800;
      94343: inst = 32'h10a00000;
      94344: inst = 32'hca0000c;
      94345: inst = 32'h24822800;
      94346: inst = 32'h10a00000;
      94347: inst = 32'hca00004;
      94348: inst = 32'h38632800;
      94349: inst = 32'h38842800;
      94350: inst = 32'h10a00001;
      94351: inst = 32'hca07093;
      94352: inst = 32'h13e00001;
      94353: inst = 32'hfe0d96a;
      94354: inst = 32'h5be00000;
      94355: inst = 32'h8c50000;
      94356: inst = 32'h24612800;
      94357: inst = 32'h10a00000;
      94358: inst = 32'hca0000c;
      94359: inst = 32'h24822800;
      94360: inst = 32'h10a00000;
      94361: inst = 32'hca00004;
      94362: inst = 32'h38632800;
      94363: inst = 32'h38842800;
      94364: inst = 32'h10a00001;
      94365: inst = 32'hca070a1;
      94366: inst = 32'h13e00001;
      94367: inst = 32'hfe0d96a;
      94368: inst = 32'h5be00000;
      94369: inst = 32'h8c50000;
      94370: inst = 32'h24612800;
      94371: inst = 32'h10a00000;
      94372: inst = 32'hca0000c;
      94373: inst = 32'h24822800;
      94374: inst = 32'h10a00000;
      94375: inst = 32'hca00004;
      94376: inst = 32'h38632800;
      94377: inst = 32'h38842800;
      94378: inst = 32'h10a00001;
      94379: inst = 32'hca070af;
      94380: inst = 32'h13e00001;
      94381: inst = 32'hfe0d96a;
      94382: inst = 32'h5be00000;
      94383: inst = 32'h8c50000;
      94384: inst = 32'h24612800;
      94385: inst = 32'h10a00000;
      94386: inst = 32'hca0000c;
      94387: inst = 32'h24822800;
      94388: inst = 32'h10a00000;
      94389: inst = 32'hca00004;
      94390: inst = 32'h38632800;
      94391: inst = 32'h38842800;
      94392: inst = 32'h10a00001;
      94393: inst = 32'hca070bd;
      94394: inst = 32'h13e00001;
      94395: inst = 32'hfe0d96a;
      94396: inst = 32'h5be00000;
      94397: inst = 32'h8c50000;
      94398: inst = 32'h24612800;
      94399: inst = 32'h10a00000;
      94400: inst = 32'hca0000c;
      94401: inst = 32'h24822800;
      94402: inst = 32'h10a00000;
      94403: inst = 32'hca00004;
      94404: inst = 32'h38632800;
      94405: inst = 32'h38842800;
      94406: inst = 32'h10a00001;
      94407: inst = 32'hca070cb;
      94408: inst = 32'h13e00001;
      94409: inst = 32'hfe0d96a;
      94410: inst = 32'h5be00000;
      94411: inst = 32'h8c50000;
      94412: inst = 32'h24612800;
      94413: inst = 32'h10a00000;
      94414: inst = 32'hca0000c;
      94415: inst = 32'h24822800;
      94416: inst = 32'h10a00000;
      94417: inst = 32'hca00004;
      94418: inst = 32'h38632800;
      94419: inst = 32'h38842800;
      94420: inst = 32'h10a00001;
      94421: inst = 32'hca070d9;
      94422: inst = 32'h13e00001;
      94423: inst = 32'hfe0d96a;
      94424: inst = 32'h5be00000;
      94425: inst = 32'h8c50000;
      94426: inst = 32'h24612800;
      94427: inst = 32'h10a00000;
      94428: inst = 32'hca0000c;
      94429: inst = 32'h24822800;
      94430: inst = 32'h10a00000;
      94431: inst = 32'hca00004;
      94432: inst = 32'h38632800;
      94433: inst = 32'h38842800;
      94434: inst = 32'h10a00001;
      94435: inst = 32'hca070e7;
      94436: inst = 32'h13e00001;
      94437: inst = 32'hfe0d96a;
      94438: inst = 32'h5be00000;
      94439: inst = 32'h8c50000;
      94440: inst = 32'h24612800;
      94441: inst = 32'h10a00000;
      94442: inst = 32'hca0000c;
      94443: inst = 32'h24822800;
      94444: inst = 32'h10a00000;
      94445: inst = 32'hca00004;
      94446: inst = 32'h38632800;
      94447: inst = 32'h38842800;
      94448: inst = 32'h10a00001;
      94449: inst = 32'hca070f5;
      94450: inst = 32'h13e00001;
      94451: inst = 32'hfe0d96a;
      94452: inst = 32'h5be00000;
      94453: inst = 32'h8c50000;
      94454: inst = 32'h24612800;
      94455: inst = 32'h10a00000;
      94456: inst = 32'hca0000c;
      94457: inst = 32'h24822800;
      94458: inst = 32'h10a00000;
      94459: inst = 32'hca00004;
      94460: inst = 32'h38632800;
      94461: inst = 32'h38842800;
      94462: inst = 32'h10a00001;
      94463: inst = 32'hca07103;
      94464: inst = 32'h13e00001;
      94465: inst = 32'hfe0d96a;
      94466: inst = 32'h5be00000;
      94467: inst = 32'h8c50000;
      94468: inst = 32'h24612800;
      94469: inst = 32'h10a00000;
      94470: inst = 32'hca0000c;
      94471: inst = 32'h24822800;
      94472: inst = 32'h10a00000;
      94473: inst = 32'hca00004;
      94474: inst = 32'h38632800;
      94475: inst = 32'h38842800;
      94476: inst = 32'h10a00001;
      94477: inst = 32'hca07111;
      94478: inst = 32'h13e00001;
      94479: inst = 32'hfe0d96a;
      94480: inst = 32'h5be00000;
      94481: inst = 32'h8c50000;
      94482: inst = 32'h24612800;
      94483: inst = 32'h10a00000;
      94484: inst = 32'hca0000c;
      94485: inst = 32'h24822800;
      94486: inst = 32'h10a00000;
      94487: inst = 32'hca00004;
      94488: inst = 32'h38632800;
      94489: inst = 32'h38842800;
      94490: inst = 32'h10a00001;
      94491: inst = 32'hca0711f;
      94492: inst = 32'h13e00001;
      94493: inst = 32'hfe0d96a;
      94494: inst = 32'h5be00000;
      94495: inst = 32'h8c50000;
      94496: inst = 32'h24612800;
      94497: inst = 32'h10a00000;
      94498: inst = 32'hca0000c;
      94499: inst = 32'h24822800;
      94500: inst = 32'h10a00000;
      94501: inst = 32'hca00004;
      94502: inst = 32'h38632800;
      94503: inst = 32'h38842800;
      94504: inst = 32'h10a00001;
      94505: inst = 32'hca0712d;
      94506: inst = 32'h13e00001;
      94507: inst = 32'hfe0d96a;
      94508: inst = 32'h5be00000;
      94509: inst = 32'h8c50000;
      94510: inst = 32'h24612800;
      94511: inst = 32'h10a00000;
      94512: inst = 32'hca0000c;
      94513: inst = 32'h24822800;
      94514: inst = 32'h10a00000;
      94515: inst = 32'hca00004;
      94516: inst = 32'h38632800;
      94517: inst = 32'h38842800;
      94518: inst = 32'h10a00001;
      94519: inst = 32'hca0713b;
      94520: inst = 32'h13e00001;
      94521: inst = 32'hfe0d96a;
      94522: inst = 32'h5be00000;
      94523: inst = 32'h8c50000;
      94524: inst = 32'h24612800;
      94525: inst = 32'h10a00000;
      94526: inst = 32'hca0000c;
      94527: inst = 32'h24822800;
      94528: inst = 32'h10a00000;
      94529: inst = 32'hca00004;
      94530: inst = 32'h38632800;
      94531: inst = 32'h38842800;
      94532: inst = 32'h10a00001;
      94533: inst = 32'hca07149;
      94534: inst = 32'h13e00001;
      94535: inst = 32'hfe0d96a;
      94536: inst = 32'h5be00000;
      94537: inst = 32'h8c50000;
      94538: inst = 32'h24612800;
      94539: inst = 32'h10a00000;
      94540: inst = 32'hca0000c;
      94541: inst = 32'h24822800;
      94542: inst = 32'h10a00000;
      94543: inst = 32'hca00004;
      94544: inst = 32'h38632800;
      94545: inst = 32'h38842800;
      94546: inst = 32'h10a00001;
      94547: inst = 32'hca07157;
      94548: inst = 32'h13e00001;
      94549: inst = 32'hfe0d96a;
      94550: inst = 32'h5be00000;
      94551: inst = 32'h8c50000;
      94552: inst = 32'h24612800;
      94553: inst = 32'h10a00000;
      94554: inst = 32'hca0000c;
      94555: inst = 32'h24822800;
      94556: inst = 32'h10a00000;
      94557: inst = 32'hca00004;
      94558: inst = 32'h38632800;
      94559: inst = 32'h38842800;
      94560: inst = 32'h10a00001;
      94561: inst = 32'hca07165;
      94562: inst = 32'h13e00001;
      94563: inst = 32'hfe0d96a;
      94564: inst = 32'h5be00000;
      94565: inst = 32'h8c50000;
      94566: inst = 32'h24612800;
      94567: inst = 32'h10a00000;
      94568: inst = 32'hca0000c;
      94569: inst = 32'h24822800;
      94570: inst = 32'h10a00000;
      94571: inst = 32'hca00004;
      94572: inst = 32'h38632800;
      94573: inst = 32'h38842800;
      94574: inst = 32'h10a00001;
      94575: inst = 32'hca07173;
      94576: inst = 32'h13e00001;
      94577: inst = 32'hfe0d96a;
      94578: inst = 32'h5be00000;
      94579: inst = 32'h8c50000;
      94580: inst = 32'h24612800;
      94581: inst = 32'h10a00000;
      94582: inst = 32'hca0000c;
      94583: inst = 32'h24822800;
      94584: inst = 32'h10a00000;
      94585: inst = 32'hca00004;
      94586: inst = 32'h38632800;
      94587: inst = 32'h38842800;
      94588: inst = 32'h10a00001;
      94589: inst = 32'hca07181;
      94590: inst = 32'h13e00001;
      94591: inst = 32'hfe0d96a;
      94592: inst = 32'h5be00000;
      94593: inst = 32'h8c50000;
      94594: inst = 32'h24612800;
      94595: inst = 32'h10a00000;
      94596: inst = 32'hca0000c;
      94597: inst = 32'h24822800;
      94598: inst = 32'h10a00000;
      94599: inst = 32'hca00004;
      94600: inst = 32'h38632800;
      94601: inst = 32'h38842800;
      94602: inst = 32'h10a00001;
      94603: inst = 32'hca0718f;
      94604: inst = 32'h13e00001;
      94605: inst = 32'hfe0d96a;
      94606: inst = 32'h5be00000;
      94607: inst = 32'h8c50000;
      94608: inst = 32'h24612800;
      94609: inst = 32'h10a00000;
      94610: inst = 32'hca0000c;
      94611: inst = 32'h24822800;
      94612: inst = 32'h10a00000;
      94613: inst = 32'hca00004;
      94614: inst = 32'h38632800;
      94615: inst = 32'h38842800;
      94616: inst = 32'h10a00001;
      94617: inst = 32'hca0719d;
      94618: inst = 32'h13e00001;
      94619: inst = 32'hfe0d96a;
      94620: inst = 32'h5be00000;
      94621: inst = 32'h8c50000;
      94622: inst = 32'h24612800;
      94623: inst = 32'h10a00000;
      94624: inst = 32'hca0000c;
      94625: inst = 32'h24822800;
      94626: inst = 32'h10a00000;
      94627: inst = 32'hca00004;
      94628: inst = 32'h38632800;
      94629: inst = 32'h38842800;
      94630: inst = 32'h10a00001;
      94631: inst = 32'hca071ab;
      94632: inst = 32'h13e00001;
      94633: inst = 32'hfe0d96a;
      94634: inst = 32'h5be00000;
      94635: inst = 32'h8c50000;
      94636: inst = 32'h24612800;
      94637: inst = 32'h10a00000;
      94638: inst = 32'hca0000c;
      94639: inst = 32'h24822800;
      94640: inst = 32'h10a00000;
      94641: inst = 32'hca00004;
      94642: inst = 32'h38632800;
      94643: inst = 32'h38842800;
      94644: inst = 32'h10a00001;
      94645: inst = 32'hca071b9;
      94646: inst = 32'h13e00001;
      94647: inst = 32'hfe0d96a;
      94648: inst = 32'h5be00000;
      94649: inst = 32'h8c50000;
      94650: inst = 32'h24612800;
      94651: inst = 32'h10a00000;
      94652: inst = 32'hca0000c;
      94653: inst = 32'h24822800;
      94654: inst = 32'h10a00000;
      94655: inst = 32'hca00004;
      94656: inst = 32'h38632800;
      94657: inst = 32'h38842800;
      94658: inst = 32'h10a00001;
      94659: inst = 32'hca071c7;
      94660: inst = 32'h13e00001;
      94661: inst = 32'hfe0d96a;
      94662: inst = 32'h5be00000;
      94663: inst = 32'h8c50000;
      94664: inst = 32'h24612800;
      94665: inst = 32'h10a00000;
      94666: inst = 32'hca0000c;
      94667: inst = 32'h24822800;
      94668: inst = 32'h10a00000;
      94669: inst = 32'hca00004;
      94670: inst = 32'h38632800;
      94671: inst = 32'h38842800;
      94672: inst = 32'h10a00001;
      94673: inst = 32'hca071d5;
      94674: inst = 32'h13e00001;
      94675: inst = 32'hfe0d96a;
      94676: inst = 32'h5be00000;
      94677: inst = 32'h8c50000;
      94678: inst = 32'h24612800;
      94679: inst = 32'h10a00000;
      94680: inst = 32'hca0000c;
      94681: inst = 32'h24822800;
      94682: inst = 32'h10a00000;
      94683: inst = 32'hca00004;
      94684: inst = 32'h38632800;
      94685: inst = 32'h38842800;
      94686: inst = 32'h10a00001;
      94687: inst = 32'hca071e3;
      94688: inst = 32'h13e00001;
      94689: inst = 32'hfe0d96a;
      94690: inst = 32'h5be00000;
      94691: inst = 32'h8c50000;
      94692: inst = 32'h24612800;
      94693: inst = 32'h10a00000;
      94694: inst = 32'hca0000c;
      94695: inst = 32'h24822800;
      94696: inst = 32'h10a00000;
      94697: inst = 32'hca00004;
      94698: inst = 32'h38632800;
      94699: inst = 32'h38842800;
      94700: inst = 32'h10a00001;
      94701: inst = 32'hca071f1;
      94702: inst = 32'h13e00001;
      94703: inst = 32'hfe0d96a;
      94704: inst = 32'h5be00000;
      94705: inst = 32'h8c50000;
      94706: inst = 32'h24612800;
      94707: inst = 32'h10a00000;
      94708: inst = 32'hca0000c;
      94709: inst = 32'h24822800;
      94710: inst = 32'h10a00000;
      94711: inst = 32'hca00004;
      94712: inst = 32'h38632800;
      94713: inst = 32'h38842800;
      94714: inst = 32'h10a00001;
      94715: inst = 32'hca071ff;
      94716: inst = 32'h13e00001;
      94717: inst = 32'hfe0d96a;
      94718: inst = 32'h5be00000;
      94719: inst = 32'h8c50000;
      94720: inst = 32'h24612800;
      94721: inst = 32'h10a00000;
      94722: inst = 32'hca0000c;
      94723: inst = 32'h24822800;
      94724: inst = 32'h10a00000;
      94725: inst = 32'hca00004;
      94726: inst = 32'h38632800;
      94727: inst = 32'h38842800;
      94728: inst = 32'h10a00001;
      94729: inst = 32'hca0720d;
      94730: inst = 32'h13e00001;
      94731: inst = 32'hfe0d96a;
      94732: inst = 32'h5be00000;
      94733: inst = 32'h8c50000;
      94734: inst = 32'h24612800;
      94735: inst = 32'h10a00000;
      94736: inst = 32'hca0000c;
      94737: inst = 32'h24822800;
      94738: inst = 32'h10a00000;
      94739: inst = 32'hca00004;
      94740: inst = 32'h38632800;
      94741: inst = 32'h38842800;
      94742: inst = 32'h10a00001;
      94743: inst = 32'hca0721b;
      94744: inst = 32'h13e00001;
      94745: inst = 32'hfe0d96a;
      94746: inst = 32'h5be00000;
      94747: inst = 32'h8c50000;
      94748: inst = 32'h24612800;
      94749: inst = 32'h10a00000;
      94750: inst = 32'hca0000c;
      94751: inst = 32'h24822800;
      94752: inst = 32'h10a00000;
      94753: inst = 32'hca00004;
      94754: inst = 32'h38632800;
      94755: inst = 32'h38842800;
      94756: inst = 32'h10a00001;
      94757: inst = 32'hca07229;
      94758: inst = 32'h13e00001;
      94759: inst = 32'hfe0d96a;
      94760: inst = 32'h5be00000;
      94761: inst = 32'h8c50000;
      94762: inst = 32'h24612800;
      94763: inst = 32'h10a00000;
      94764: inst = 32'hca0000c;
      94765: inst = 32'h24822800;
      94766: inst = 32'h10a00000;
      94767: inst = 32'hca00004;
      94768: inst = 32'h38632800;
      94769: inst = 32'h38842800;
      94770: inst = 32'h10a00001;
      94771: inst = 32'hca07237;
      94772: inst = 32'h13e00001;
      94773: inst = 32'hfe0d96a;
      94774: inst = 32'h5be00000;
      94775: inst = 32'h8c50000;
      94776: inst = 32'h24612800;
      94777: inst = 32'h10a00000;
      94778: inst = 32'hca0000c;
      94779: inst = 32'h24822800;
      94780: inst = 32'h10a00000;
      94781: inst = 32'hca00004;
      94782: inst = 32'h38632800;
      94783: inst = 32'h38842800;
      94784: inst = 32'h10a00001;
      94785: inst = 32'hca07245;
      94786: inst = 32'h13e00001;
      94787: inst = 32'hfe0d96a;
      94788: inst = 32'h5be00000;
      94789: inst = 32'h8c50000;
      94790: inst = 32'h24612800;
      94791: inst = 32'h10a00000;
      94792: inst = 32'hca0000c;
      94793: inst = 32'h24822800;
      94794: inst = 32'h10a00000;
      94795: inst = 32'hca00004;
      94796: inst = 32'h38632800;
      94797: inst = 32'h38842800;
      94798: inst = 32'h10a00001;
      94799: inst = 32'hca07253;
      94800: inst = 32'h13e00001;
      94801: inst = 32'hfe0d96a;
      94802: inst = 32'h5be00000;
      94803: inst = 32'h8c50000;
      94804: inst = 32'h24612800;
      94805: inst = 32'h10a00000;
      94806: inst = 32'hca0000c;
      94807: inst = 32'h24822800;
      94808: inst = 32'h10a00000;
      94809: inst = 32'hca00004;
      94810: inst = 32'h38632800;
      94811: inst = 32'h38842800;
      94812: inst = 32'h10a00001;
      94813: inst = 32'hca07261;
      94814: inst = 32'h13e00001;
      94815: inst = 32'hfe0d96a;
      94816: inst = 32'h5be00000;
      94817: inst = 32'h8c50000;
      94818: inst = 32'h24612800;
      94819: inst = 32'h10a00000;
      94820: inst = 32'hca0000c;
      94821: inst = 32'h24822800;
      94822: inst = 32'h10a00000;
      94823: inst = 32'hca00004;
      94824: inst = 32'h38632800;
      94825: inst = 32'h38842800;
      94826: inst = 32'h10a00001;
      94827: inst = 32'hca0726f;
      94828: inst = 32'h13e00001;
      94829: inst = 32'hfe0d96a;
      94830: inst = 32'h5be00000;
      94831: inst = 32'h8c50000;
      94832: inst = 32'h24612800;
      94833: inst = 32'h10a00000;
      94834: inst = 32'hca0000c;
      94835: inst = 32'h24822800;
      94836: inst = 32'h10a00000;
      94837: inst = 32'hca00004;
      94838: inst = 32'h38632800;
      94839: inst = 32'h38842800;
      94840: inst = 32'h10a00001;
      94841: inst = 32'hca0727d;
      94842: inst = 32'h13e00001;
      94843: inst = 32'hfe0d96a;
      94844: inst = 32'h5be00000;
      94845: inst = 32'h8c50000;
      94846: inst = 32'h24612800;
      94847: inst = 32'h10a00000;
      94848: inst = 32'hca0000c;
      94849: inst = 32'h24822800;
      94850: inst = 32'h10a00000;
      94851: inst = 32'hca00004;
      94852: inst = 32'h38632800;
      94853: inst = 32'h38842800;
      94854: inst = 32'h10a00001;
      94855: inst = 32'hca0728b;
      94856: inst = 32'h13e00001;
      94857: inst = 32'hfe0d96a;
      94858: inst = 32'h5be00000;
      94859: inst = 32'h8c50000;
      94860: inst = 32'h24612800;
      94861: inst = 32'h10a00000;
      94862: inst = 32'hca0000c;
      94863: inst = 32'h24822800;
      94864: inst = 32'h10a00000;
      94865: inst = 32'hca00004;
      94866: inst = 32'h38632800;
      94867: inst = 32'h38842800;
      94868: inst = 32'h10a00001;
      94869: inst = 32'hca07299;
      94870: inst = 32'h13e00001;
      94871: inst = 32'hfe0d96a;
      94872: inst = 32'h5be00000;
      94873: inst = 32'h8c50000;
      94874: inst = 32'h24612800;
      94875: inst = 32'h10a00000;
      94876: inst = 32'hca0000c;
      94877: inst = 32'h24822800;
      94878: inst = 32'h10a00000;
      94879: inst = 32'hca00004;
      94880: inst = 32'h38632800;
      94881: inst = 32'h38842800;
      94882: inst = 32'h10a00001;
      94883: inst = 32'hca072a7;
      94884: inst = 32'h13e00001;
      94885: inst = 32'hfe0d96a;
      94886: inst = 32'h5be00000;
      94887: inst = 32'h8c50000;
      94888: inst = 32'h24612800;
      94889: inst = 32'h10a00000;
      94890: inst = 32'hca0000c;
      94891: inst = 32'h24822800;
      94892: inst = 32'h10a00000;
      94893: inst = 32'hca00004;
      94894: inst = 32'h38632800;
      94895: inst = 32'h38842800;
      94896: inst = 32'h10a00001;
      94897: inst = 32'hca072b5;
      94898: inst = 32'h13e00001;
      94899: inst = 32'hfe0d96a;
      94900: inst = 32'h5be00000;
      94901: inst = 32'h8c50000;
      94902: inst = 32'h24612800;
      94903: inst = 32'h10a00000;
      94904: inst = 32'hca0000c;
      94905: inst = 32'h24822800;
      94906: inst = 32'h10a00000;
      94907: inst = 32'hca00004;
      94908: inst = 32'h38632800;
      94909: inst = 32'h38842800;
      94910: inst = 32'h10a00001;
      94911: inst = 32'hca072c3;
      94912: inst = 32'h13e00001;
      94913: inst = 32'hfe0d96a;
      94914: inst = 32'h5be00000;
      94915: inst = 32'h8c50000;
      94916: inst = 32'h24612800;
      94917: inst = 32'h10a00000;
      94918: inst = 32'hca0000c;
      94919: inst = 32'h24822800;
      94920: inst = 32'h10a00000;
      94921: inst = 32'hca00004;
      94922: inst = 32'h38632800;
      94923: inst = 32'h38842800;
      94924: inst = 32'h10a00001;
      94925: inst = 32'hca072d1;
      94926: inst = 32'h13e00001;
      94927: inst = 32'hfe0d96a;
      94928: inst = 32'h5be00000;
      94929: inst = 32'h8c50000;
      94930: inst = 32'h24612800;
      94931: inst = 32'h10a00000;
      94932: inst = 32'hca0000c;
      94933: inst = 32'h24822800;
      94934: inst = 32'h10a00000;
      94935: inst = 32'hca00004;
      94936: inst = 32'h38632800;
      94937: inst = 32'h38842800;
      94938: inst = 32'h10a00001;
      94939: inst = 32'hca072df;
      94940: inst = 32'h13e00001;
      94941: inst = 32'hfe0d96a;
      94942: inst = 32'h5be00000;
      94943: inst = 32'h8c50000;
      94944: inst = 32'h24612800;
      94945: inst = 32'h10a00000;
      94946: inst = 32'hca0000c;
      94947: inst = 32'h24822800;
      94948: inst = 32'h10a00000;
      94949: inst = 32'hca00004;
      94950: inst = 32'h38632800;
      94951: inst = 32'h38842800;
      94952: inst = 32'h10a00001;
      94953: inst = 32'hca072ed;
      94954: inst = 32'h13e00001;
      94955: inst = 32'hfe0d96a;
      94956: inst = 32'h5be00000;
      94957: inst = 32'h8c50000;
      94958: inst = 32'h24612800;
      94959: inst = 32'h10a00000;
      94960: inst = 32'hca0000c;
      94961: inst = 32'h24822800;
      94962: inst = 32'h10a00000;
      94963: inst = 32'hca00004;
      94964: inst = 32'h38632800;
      94965: inst = 32'h38842800;
      94966: inst = 32'h10a00001;
      94967: inst = 32'hca072fb;
      94968: inst = 32'h13e00001;
      94969: inst = 32'hfe0d96a;
      94970: inst = 32'h5be00000;
      94971: inst = 32'h8c50000;
      94972: inst = 32'h24612800;
      94973: inst = 32'h10a00000;
      94974: inst = 32'hca0000c;
      94975: inst = 32'h24822800;
      94976: inst = 32'h10a00000;
      94977: inst = 32'hca00004;
      94978: inst = 32'h38632800;
      94979: inst = 32'h38842800;
      94980: inst = 32'h10a00001;
      94981: inst = 32'hca07309;
      94982: inst = 32'h13e00001;
      94983: inst = 32'hfe0d96a;
      94984: inst = 32'h5be00000;
      94985: inst = 32'h8c50000;
      94986: inst = 32'h24612800;
      94987: inst = 32'h10a00000;
      94988: inst = 32'hca0000c;
      94989: inst = 32'h24822800;
      94990: inst = 32'h10a00000;
      94991: inst = 32'hca00004;
      94992: inst = 32'h38632800;
      94993: inst = 32'h38842800;
      94994: inst = 32'h10a00001;
      94995: inst = 32'hca07317;
      94996: inst = 32'h13e00001;
      94997: inst = 32'hfe0d96a;
      94998: inst = 32'h5be00000;
      94999: inst = 32'h8c50000;
      95000: inst = 32'h24612800;
      95001: inst = 32'h10a00000;
      95002: inst = 32'hca0000c;
      95003: inst = 32'h24822800;
      95004: inst = 32'h10a00000;
      95005: inst = 32'hca00004;
      95006: inst = 32'h38632800;
      95007: inst = 32'h38842800;
      95008: inst = 32'h10a00001;
      95009: inst = 32'hca07325;
      95010: inst = 32'h13e00001;
      95011: inst = 32'hfe0d96a;
      95012: inst = 32'h5be00000;
      95013: inst = 32'h8c50000;
      95014: inst = 32'h24612800;
      95015: inst = 32'h10a00000;
      95016: inst = 32'hca0000c;
      95017: inst = 32'h24822800;
      95018: inst = 32'h10a00000;
      95019: inst = 32'hca00004;
      95020: inst = 32'h38632800;
      95021: inst = 32'h38842800;
      95022: inst = 32'h10a00001;
      95023: inst = 32'hca07333;
      95024: inst = 32'h13e00001;
      95025: inst = 32'hfe0d96a;
      95026: inst = 32'h5be00000;
      95027: inst = 32'h8c50000;
      95028: inst = 32'h24612800;
      95029: inst = 32'h10a00000;
      95030: inst = 32'hca0000c;
      95031: inst = 32'h24822800;
      95032: inst = 32'h10a00000;
      95033: inst = 32'hca00004;
      95034: inst = 32'h38632800;
      95035: inst = 32'h38842800;
      95036: inst = 32'h10a00001;
      95037: inst = 32'hca07341;
      95038: inst = 32'h13e00001;
      95039: inst = 32'hfe0d96a;
      95040: inst = 32'h5be00000;
      95041: inst = 32'h8c50000;
      95042: inst = 32'h24612800;
      95043: inst = 32'h10a00000;
      95044: inst = 32'hca0000c;
      95045: inst = 32'h24822800;
      95046: inst = 32'h10a00000;
      95047: inst = 32'hca00004;
      95048: inst = 32'h38632800;
      95049: inst = 32'h38842800;
      95050: inst = 32'h10a00001;
      95051: inst = 32'hca0734f;
      95052: inst = 32'h13e00001;
      95053: inst = 32'hfe0d96a;
      95054: inst = 32'h5be00000;
      95055: inst = 32'h8c50000;
      95056: inst = 32'h24612800;
      95057: inst = 32'h10a00000;
      95058: inst = 32'hca0000c;
      95059: inst = 32'h24822800;
      95060: inst = 32'h10a00000;
      95061: inst = 32'hca00004;
      95062: inst = 32'h38632800;
      95063: inst = 32'h38842800;
      95064: inst = 32'h10a00001;
      95065: inst = 32'hca0735d;
      95066: inst = 32'h13e00001;
      95067: inst = 32'hfe0d96a;
      95068: inst = 32'h5be00000;
      95069: inst = 32'h8c50000;
      95070: inst = 32'h24612800;
      95071: inst = 32'h10a00000;
      95072: inst = 32'hca0000c;
      95073: inst = 32'h24822800;
      95074: inst = 32'h10a00000;
      95075: inst = 32'hca00004;
      95076: inst = 32'h38632800;
      95077: inst = 32'h38842800;
      95078: inst = 32'h10a00001;
      95079: inst = 32'hca0736b;
      95080: inst = 32'h13e00001;
      95081: inst = 32'hfe0d96a;
      95082: inst = 32'h5be00000;
      95083: inst = 32'h8c50000;
      95084: inst = 32'h24612800;
      95085: inst = 32'h10a00000;
      95086: inst = 32'hca0000c;
      95087: inst = 32'h24822800;
      95088: inst = 32'h10a00000;
      95089: inst = 32'hca00004;
      95090: inst = 32'h38632800;
      95091: inst = 32'h38842800;
      95092: inst = 32'h10a00001;
      95093: inst = 32'hca07379;
      95094: inst = 32'h13e00001;
      95095: inst = 32'hfe0d96a;
      95096: inst = 32'h5be00000;
      95097: inst = 32'h8c50000;
      95098: inst = 32'h24612800;
      95099: inst = 32'h10a00000;
      95100: inst = 32'hca0000c;
      95101: inst = 32'h24822800;
      95102: inst = 32'h10a00000;
      95103: inst = 32'hca00004;
      95104: inst = 32'h38632800;
      95105: inst = 32'h38842800;
      95106: inst = 32'h10a00001;
      95107: inst = 32'hca07387;
      95108: inst = 32'h13e00001;
      95109: inst = 32'hfe0d96a;
      95110: inst = 32'h5be00000;
      95111: inst = 32'h8c50000;
      95112: inst = 32'h24612800;
      95113: inst = 32'h10a00000;
      95114: inst = 32'hca0000c;
      95115: inst = 32'h24822800;
      95116: inst = 32'h10a00000;
      95117: inst = 32'hca00004;
      95118: inst = 32'h38632800;
      95119: inst = 32'h38842800;
      95120: inst = 32'h10a00001;
      95121: inst = 32'hca07395;
      95122: inst = 32'h13e00001;
      95123: inst = 32'hfe0d96a;
      95124: inst = 32'h5be00000;
      95125: inst = 32'h8c50000;
      95126: inst = 32'h24612800;
      95127: inst = 32'h10a00000;
      95128: inst = 32'hca0000c;
      95129: inst = 32'h24822800;
      95130: inst = 32'h10a00000;
      95131: inst = 32'hca00004;
      95132: inst = 32'h38632800;
      95133: inst = 32'h38842800;
      95134: inst = 32'h10a00001;
      95135: inst = 32'hca073a3;
      95136: inst = 32'h13e00001;
      95137: inst = 32'hfe0d96a;
      95138: inst = 32'h5be00000;
      95139: inst = 32'h8c50000;
      95140: inst = 32'h24612800;
      95141: inst = 32'h10a00000;
      95142: inst = 32'hca0000c;
      95143: inst = 32'h24822800;
      95144: inst = 32'h10a00000;
      95145: inst = 32'hca00004;
      95146: inst = 32'h38632800;
      95147: inst = 32'h38842800;
      95148: inst = 32'h10a00001;
      95149: inst = 32'hca073b1;
      95150: inst = 32'h13e00001;
      95151: inst = 32'hfe0d96a;
      95152: inst = 32'h5be00000;
      95153: inst = 32'h8c50000;
      95154: inst = 32'h24612800;
      95155: inst = 32'h10a00000;
      95156: inst = 32'hca0000c;
      95157: inst = 32'h24822800;
      95158: inst = 32'h10a00000;
      95159: inst = 32'hca00004;
      95160: inst = 32'h38632800;
      95161: inst = 32'h38842800;
      95162: inst = 32'h10a00001;
      95163: inst = 32'hca073bf;
      95164: inst = 32'h13e00001;
      95165: inst = 32'hfe0d96a;
      95166: inst = 32'h5be00000;
      95167: inst = 32'h8c50000;
      95168: inst = 32'h24612800;
      95169: inst = 32'h10a00000;
      95170: inst = 32'hca0000c;
      95171: inst = 32'h24822800;
      95172: inst = 32'h10a00000;
      95173: inst = 32'hca00004;
      95174: inst = 32'h38632800;
      95175: inst = 32'h38842800;
      95176: inst = 32'h10a00001;
      95177: inst = 32'hca073cd;
      95178: inst = 32'h13e00001;
      95179: inst = 32'hfe0d96a;
      95180: inst = 32'h5be00000;
      95181: inst = 32'h8c50000;
      95182: inst = 32'h24612800;
      95183: inst = 32'h10a00000;
      95184: inst = 32'hca0000c;
      95185: inst = 32'h24822800;
      95186: inst = 32'h10a00000;
      95187: inst = 32'hca00004;
      95188: inst = 32'h38632800;
      95189: inst = 32'h38842800;
      95190: inst = 32'h10a00001;
      95191: inst = 32'hca073db;
      95192: inst = 32'h13e00001;
      95193: inst = 32'hfe0d96a;
      95194: inst = 32'h5be00000;
      95195: inst = 32'h8c50000;
      95196: inst = 32'h24612800;
      95197: inst = 32'h10a00000;
      95198: inst = 32'hca0000c;
      95199: inst = 32'h24822800;
      95200: inst = 32'h10a00000;
      95201: inst = 32'hca00004;
      95202: inst = 32'h38632800;
      95203: inst = 32'h38842800;
      95204: inst = 32'h10a00001;
      95205: inst = 32'hca073e9;
      95206: inst = 32'h13e00001;
      95207: inst = 32'hfe0d96a;
      95208: inst = 32'h5be00000;
      95209: inst = 32'h8c50000;
      95210: inst = 32'h24612800;
      95211: inst = 32'h10a00000;
      95212: inst = 32'hca0000c;
      95213: inst = 32'h24822800;
      95214: inst = 32'h10a00000;
      95215: inst = 32'hca00004;
      95216: inst = 32'h38632800;
      95217: inst = 32'h38842800;
      95218: inst = 32'h10a00001;
      95219: inst = 32'hca073f7;
      95220: inst = 32'h13e00001;
      95221: inst = 32'hfe0d96a;
      95222: inst = 32'h5be00000;
      95223: inst = 32'h8c50000;
      95224: inst = 32'h24612800;
      95225: inst = 32'h10a00000;
      95226: inst = 32'hca0000c;
      95227: inst = 32'h24822800;
      95228: inst = 32'h10a00000;
      95229: inst = 32'hca00004;
      95230: inst = 32'h38632800;
      95231: inst = 32'h38842800;
      95232: inst = 32'h10a00001;
      95233: inst = 32'hca07405;
      95234: inst = 32'h13e00001;
      95235: inst = 32'hfe0d96a;
      95236: inst = 32'h5be00000;
      95237: inst = 32'h8c50000;
      95238: inst = 32'h24612800;
      95239: inst = 32'h10a00000;
      95240: inst = 32'hca0000c;
      95241: inst = 32'h24822800;
      95242: inst = 32'h10a00000;
      95243: inst = 32'hca00004;
      95244: inst = 32'h38632800;
      95245: inst = 32'h38842800;
      95246: inst = 32'h10a00001;
      95247: inst = 32'hca07413;
      95248: inst = 32'h13e00001;
      95249: inst = 32'hfe0d96a;
      95250: inst = 32'h5be00000;
      95251: inst = 32'h8c50000;
      95252: inst = 32'h24612800;
      95253: inst = 32'h10a00000;
      95254: inst = 32'hca0000c;
      95255: inst = 32'h24822800;
      95256: inst = 32'h10a00000;
      95257: inst = 32'hca00004;
      95258: inst = 32'h38632800;
      95259: inst = 32'h38842800;
      95260: inst = 32'h10a00001;
      95261: inst = 32'hca07421;
      95262: inst = 32'h13e00001;
      95263: inst = 32'hfe0d96a;
      95264: inst = 32'h5be00000;
      95265: inst = 32'h8c50000;
      95266: inst = 32'h24612800;
      95267: inst = 32'h10a00000;
      95268: inst = 32'hca0000c;
      95269: inst = 32'h24822800;
      95270: inst = 32'h10a00000;
      95271: inst = 32'hca00004;
      95272: inst = 32'h38632800;
      95273: inst = 32'h38842800;
      95274: inst = 32'h10a00001;
      95275: inst = 32'hca0742f;
      95276: inst = 32'h13e00001;
      95277: inst = 32'hfe0d96a;
      95278: inst = 32'h5be00000;
      95279: inst = 32'h8c50000;
      95280: inst = 32'h24612800;
      95281: inst = 32'h10a00000;
      95282: inst = 32'hca0000c;
      95283: inst = 32'h24822800;
      95284: inst = 32'h10a00000;
      95285: inst = 32'hca00004;
      95286: inst = 32'h38632800;
      95287: inst = 32'h38842800;
      95288: inst = 32'h10a00001;
      95289: inst = 32'hca0743d;
      95290: inst = 32'h13e00001;
      95291: inst = 32'hfe0d96a;
      95292: inst = 32'h5be00000;
      95293: inst = 32'h8c50000;
      95294: inst = 32'h24612800;
      95295: inst = 32'h10a00000;
      95296: inst = 32'hca0000c;
      95297: inst = 32'h24822800;
      95298: inst = 32'h10a00000;
      95299: inst = 32'hca00004;
      95300: inst = 32'h38632800;
      95301: inst = 32'h38842800;
      95302: inst = 32'h10a00001;
      95303: inst = 32'hca0744b;
      95304: inst = 32'h13e00001;
      95305: inst = 32'hfe0d96a;
      95306: inst = 32'h5be00000;
      95307: inst = 32'h8c50000;
      95308: inst = 32'h24612800;
      95309: inst = 32'h10a00000;
      95310: inst = 32'hca0000c;
      95311: inst = 32'h24822800;
      95312: inst = 32'h10a00000;
      95313: inst = 32'hca00004;
      95314: inst = 32'h38632800;
      95315: inst = 32'h38842800;
      95316: inst = 32'h10a00001;
      95317: inst = 32'hca07459;
      95318: inst = 32'h13e00001;
      95319: inst = 32'hfe0d96a;
      95320: inst = 32'h5be00000;
      95321: inst = 32'h8c50000;
      95322: inst = 32'h24612800;
      95323: inst = 32'h10a00000;
      95324: inst = 32'hca0000c;
      95325: inst = 32'h24822800;
      95326: inst = 32'h10a00000;
      95327: inst = 32'hca00004;
      95328: inst = 32'h38632800;
      95329: inst = 32'h38842800;
      95330: inst = 32'h10a00001;
      95331: inst = 32'hca07467;
      95332: inst = 32'h13e00001;
      95333: inst = 32'hfe0d96a;
      95334: inst = 32'h5be00000;
      95335: inst = 32'h8c50000;
      95336: inst = 32'h24612800;
      95337: inst = 32'h10a00000;
      95338: inst = 32'hca0000c;
      95339: inst = 32'h24822800;
      95340: inst = 32'h10a00000;
      95341: inst = 32'hca00004;
      95342: inst = 32'h38632800;
      95343: inst = 32'h38842800;
      95344: inst = 32'h10a00001;
      95345: inst = 32'hca07475;
      95346: inst = 32'h13e00001;
      95347: inst = 32'hfe0d96a;
      95348: inst = 32'h5be00000;
      95349: inst = 32'h8c50000;
      95350: inst = 32'h24612800;
      95351: inst = 32'h10a00000;
      95352: inst = 32'hca0000c;
      95353: inst = 32'h24822800;
      95354: inst = 32'h10a00000;
      95355: inst = 32'hca00004;
      95356: inst = 32'h38632800;
      95357: inst = 32'h38842800;
      95358: inst = 32'h10a00001;
      95359: inst = 32'hca07483;
      95360: inst = 32'h13e00001;
      95361: inst = 32'hfe0d96a;
      95362: inst = 32'h5be00000;
      95363: inst = 32'h8c50000;
      95364: inst = 32'h24612800;
      95365: inst = 32'h10a00000;
      95366: inst = 32'hca0000c;
      95367: inst = 32'h24822800;
      95368: inst = 32'h10a00000;
      95369: inst = 32'hca00004;
      95370: inst = 32'h38632800;
      95371: inst = 32'h38842800;
      95372: inst = 32'h10a00001;
      95373: inst = 32'hca07491;
      95374: inst = 32'h13e00001;
      95375: inst = 32'hfe0d96a;
      95376: inst = 32'h5be00000;
      95377: inst = 32'h8c50000;
      95378: inst = 32'h24612800;
      95379: inst = 32'h10a00000;
      95380: inst = 32'hca0000c;
      95381: inst = 32'h24822800;
      95382: inst = 32'h10a00000;
      95383: inst = 32'hca00004;
      95384: inst = 32'h38632800;
      95385: inst = 32'h38842800;
      95386: inst = 32'h10a00001;
      95387: inst = 32'hca0749f;
      95388: inst = 32'h13e00001;
      95389: inst = 32'hfe0d96a;
      95390: inst = 32'h5be00000;
      95391: inst = 32'h8c50000;
      95392: inst = 32'h24612800;
      95393: inst = 32'h10a00000;
      95394: inst = 32'hca0000c;
      95395: inst = 32'h24822800;
      95396: inst = 32'h10a00000;
      95397: inst = 32'hca00004;
      95398: inst = 32'h38632800;
      95399: inst = 32'h38842800;
      95400: inst = 32'h10a00001;
      95401: inst = 32'hca074ad;
      95402: inst = 32'h13e00001;
      95403: inst = 32'hfe0d96a;
      95404: inst = 32'h5be00000;
      95405: inst = 32'h8c50000;
      95406: inst = 32'h24612800;
      95407: inst = 32'h10a00000;
      95408: inst = 32'hca0000c;
      95409: inst = 32'h24822800;
      95410: inst = 32'h10a00000;
      95411: inst = 32'hca00004;
      95412: inst = 32'h38632800;
      95413: inst = 32'h38842800;
      95414: inst = 32'h10a00001;
      95415: inst = 32'hca074bb;
      95416: inst = 32'h13e00001;
      95417: inst = 32'hfe0d96a;
      95418: inst = 32'h5be00000;
      95419: inst = 32'h8c50000;
      95420: inst = 32'h24612800;
      95421: inst = 32'h10a00000;
      95422: inst = 32'hca0000c;
      95423: inst = 32'h24822800;
      95424: inst = 32'h10a00000;
      95425: inst = 32'hca00004;
      95426: inst = 32'h38632800;
      95427: inst = 32'h38842800;
      95428: inst = 32'h10a00001;
      95429: inst = 32'hca074c9;
      95430: inst = 32'h13e00001;
      95431: inst = 32'hfe0d96a;
      95432: inst = 32'h5be00000;
      95433: inst = 32'h8c50000;
      95434: inst = 32'h24612800;
      95435: inst = 32'h10a00000;
      95436: inst = 32'hca0000c;
      95437: inst = 32'h24822800;
      95438: inst = 32'h10a00000;
      95439: inst = 32'hca00004;
      95440: inst = 32'h38632800;
      95441: inst = 32'h38842800;
      95442: inst = 32'h10a00001;
      95443: inst = 32'hca074d7;
      95444: inst = 32'h13e00001;
      95445: inst = 32'hfe0d96a;
      95446: inst = 32'h5be00000;
      95447: inst = 32'h8c50000;
      95448: inst = 32'h24612800;
      95449: inst = 32'h10a00000;
      95450: inst = 32'hca0000c;
      95451: inst = 32'h24822800;
      95452: inst = 32'h10a00000;
      95453: inst = 32'hca00004;
      95454: inst = 32'h38632800;
      95455: inst = 32'h38842800;
      95456: inst = 32'h10a00001;
      95457: inst = 32'hca074e5;
      95458: inst = 32'h13e00001;
      95459: inst = 32'hfe0d96a;
      95460: inst = 32'h5be00000;
      95461: inst = 32'h8c50000;
      95462: inst = 32'h24612800;
      95463: inst = 32'h10a00000;
      95464: inst = 32'hca0000c;
      95465: inst = 32'h24822800;
      95466: inst = 32'h10a00000;
      95467: inst = 32'hca00004;
      95468: inst = 32'h38632800;
      95469: inst = 32'h38842800;
      95470: inst = 32'h10a00001;
      95471: inst = 32'hca074f3;
      95472: inst = 32'h13e00001;
      95473: inst = 32'hfe0d96a;
      95474: inst = 32'h5be00000;
      95475: inst = 32'h8c50000;
      95476: inst = 32'h24612800;
      95477: inst = 32'h10a00000;
      95478: inst = 32'hca0000c;
      95479: inst = 32'h24822800;
      95480: inst = 32'h10a00000;
      95481: inst = 32'hca00004;
      95482: inst = 32'h38632800;
      95483: inst = 32'h38842800;
      95484: inst = 32'h10a00001;
      95485: inst = 32'hca07501;
      95486: inst = 32'h13e00001;
      95487: inst = 32'hfe0d96a;
      95488: inst = 32'h5be00000;
      95489: inst = 32'h8c50000;
      95490: inst = 32'h24612800;
      95491: inst = 32'h10a00000;
      95492: inst = 32'hca0000c;
      95493: inst = 32'h24822800;
      95494: inst = 32'h10a00000;
      95495: inst = 32'hca00004;
      95496: inst = 32'h38632800;
      95497: inst = 32'h38842800;
      95498: inst = 32'h10a00001;
      95499: inst = 32'hca0750f;
      95500: inst = 32'h13e00001;
      95501: inst = 32'hfe0d96a;
      95502: inst = 32'h5be00000;
      95503: inst = 32'h8c50000;
      95504: inst = 32'h24612800;
      95505: inst = 32'h10a00000;
      95506: inst = 32'hca0000c;
      95507: inst = 32'h24822800;
      95508: inst = 32'h10a00000;
      95509: inst = 32'hca00004;
      95510: inst = 32'h38632800;
      95511: inst = 32'h38842800;
      95512: inst = 32'h10a00001;
      95513: inst = 32'hca0751d;
      95514: inst = 32'h13e00001;
      95515: inst = 32'hfe0d96a;
      95516: inst = 32'h5be00000;
      95517: inst = 32'h8c50000;
      95518: inst = 32'h24612800;
      95519: inst = 32'h10a00000;
      95520: inst = 32'hca0000c;
      95521: inst = 32'h24822800;
      95522: inst = 32'h10a00000;
      95523: inst = 32'hca00004;
      95524: inst = 32'h38632800;
      95525: inst = 32'h38842800;
      95526: inst = 32'h10a00001;
      95527: inst = 32'hca0752b;
      95528: inst = 32'h13e00001;
      95529: inst = 32'hfe0d96a;
      95530: inst = 32'h5be00000;
      95531: inst = 32'h8c50000;
      95532: inst = 32'h24612800;
      95533: inst = 32'h10a00000;
      95534: inst = 32'hca0000c;
      95535: inst = 32'h24822800;
      95536: inst = 32'h10a00000;
      95537: inst = 32'hca00004;
      95538: inst = 32'h38632800;
      95539: inst = 32'h38842800;
      95540: inst = 32'h10a00001;
      95541: inst = 32'hca07539;
      95542: inst = 32'h13e00001;
      95543: inst = 32'hfe0d96a;
      95544: inst = 32'h5be00000;
      95545: inst = 32'h8c50000;
      95546: inst = 32'h24612800;
      95547: inst = 32'h10a00000;
      95548: inst = 32'hca0000c;
      95549: inst = 32'h24822800;
      95550: inst = 32'h10a00000;
      95551: inst = 32'hca00004;
      95552: inst = 32'h38632800;
      95553: inst = 32'h38842800;
      95554: inst = 32'h10a00001;
      95555: inst = 32'hca07547;
      95556: inst = 32'h13e00001;
      95557: inst = 32'hfe0d96a;
      95558: inst = 32'h5be00000;
      95559: inst = 32'h8c50000;
      95560: inst = 32'h24612800;
      95561: inst = 32'h10a00000;
      95562: inst = 32'hca0000c;
      95563: inst = 32'h24822800;
      95564: inst = 32'h10a00000;
      95565: inst = 32'hca00004;
      95566: inst = 32'h38632800;
      95567: inst = 32'h38842800;
      95568: inst = 32'h10a00001;
      95569: inst = 32'hca07555;
      95570: inst = 32'h13e00001;
      95571: inst = 32'hfe0d96a;
      95572: inst = 32'h5be00000;
      95573: inst = 32'h8c50000;
      95574: inst = 32'h24612800;
      95575: inst = 32'h10a00000;
      95576: inst = 32'hca0000c;
      95577: inst = 32'h24822800;
      95578: inst = 32'h10a00000;
      95579: inst = 32'hca00004;
      95580: inst = 32'h38632800;
      95581: inst = 32'h38842800;
      95582: inst = 32'h10a00001;
      95583: inst = 32'hca07563;
      95584: inst = 32'h13e00001;
      95585: inst = 32'hfe0d96a;
      95586: inst = 32'h5be00000;
      95587: inst = 32'h8c50000;
      95588: inst = 32'h24612800;
      95589: inst = 32'h10a00000;
      95590: inst = 32'hca0000c;
      95591: inst = 32'h24822800;
      95592: inst = 32'h10a00000;
      95593: inst = 32'hca00004;
      95594: inst = 32'h38632800;
      95595: inst = 32'h38842800;
      95596: inst = 32'h10a00001;
      95597: inst = 32'hca07571;
      95598: inst = 32'h13e00001;
      95599: inst = 32'hfe0d96a;
      95600: inst = 32'h5be00000;
      95601: inst = 32'h8c50000;
      95602: inst = 32'h24612800;
      95603: inst = 32'h10a00000;
      95604: inst = 32'hca0000c;
      95605: inst = 32'h24822800;
      95606: inst = 32'h10a00000;
      95607: inst = 32'hca00004;
      95608: inst = 32'h38632800;
      95609: inst = 32'h38842800;
      95610: inst = 32'h10a00001;
      95611: inst = 32'hca0757f;
      95612: inst = 32'h13e00001;
      95613: inst = 32'hfe0d96a;
      95614: inst = 32'h5be00000;
      95615: inst = 32'h8c50000;
      95616: inst = 32'h24612800;
      95617: inst = 32'h10a00000;
      95618: inst = 32'hca0000c;
      95619: inst = 32'h24822800;
      95620: inst = 32'h10a00000;
      95621: inst = 32'hca00004;
      95622: inst = 32'h38632800;
      95623: inst = 32'h38842800;
      95624: inst = 32'h10a00001;
      95625: inst = 32'hca0758d;
      95626: inst = 32'h13e00001;
      95627: inst = 32'hfe0d96a;
      95628: inst = 32'h5be00000;
      95629: inst = 32'h8c50000;
      95630: inst = 32'h24612800;
      95631: inst = 32'h10a00000;
      95632: inst = 32'hca0000c;
      95633: inst = 32'h24822800;
      95634: inst = 32'h10a00000;
      95635: inst = 32'hca00004;
      95636: inst = 32'h38632800;
      95637: inst = 32'h38842800;
      95638: inst = 32'h10a00001;
      95639: inst = 32'hca0759b;
      95640: inst = 32'h13e00001;
      95641: inst = 32'hfe0d96a;
      95642: inst = 32'h5be00000;
      95643: inst = 32'h8c50000;
      95644: inst = 32'h24612800;
      95645: inst = 32'h10a00000;
      95646: inst = 32'hca0000c;
      95647: inst = 32'h24822800;
      95648: inst = 32'h10a00000;
      95649: inst = 32'hca00004;
      95650: inst = 32'h38632800;
      95651: inst = 32'h38842800;
      95652: inst = 32'h10a00001;
      95653: inst = 32'hca075a9;
      95654: inst = 32'h13e00001;
      95655: inst = 32'hfe0d96a;
      95656: inst = 32'h5be00000;
      95657: inst = 32'h8c50000;
      95658: inst = 32'h24612800;
      95659: inst = 32'h10a00000;
      95660: inst = 32'hca0000d;
      95661: inst = 32'h24822800;
      95662: inst = 32'h10a00000;
      95663: inst = 32'hca00004;
      95664: inst = 32'h38632800;
      95665: inst = 32'h38842800;
      95666: inst = 32'h10a00001;
      95667: inst = 32'hca075b7;
      95668: inst = 32'h13e00001;
      95669: inst = 32'hfe0d96a;
      95670: inst = 32'h5be00000;
      95671: inst = 32'h8c50000;
      95672: inst = 32'h24612800;
      95673: inst = 32'h10a00000;
      95674: inst = 32'hca0000d;
      95675: inst = 32'h24822800;
      95676: inst = 32'h10a00000;
      95677: inst = 32'hca00004;
      95678: inst = 32'h38632800;
      95679: inst = 32'h38842800;
      95680: inst = 32'h10a00001;
      95681: inst = 32'hca075c5;
      95682: inst = 32'h13e00001;
      95683: inst = 32'hfe0d96a;
      95684: inst = 32'h5be00000;
      95685: inst = 32'h8c50000;
      95686: inst = 32'h24612800;
      95687: inst = 32'h10a00000;
      95688: inst = 32'hca0000d;
      95689: inst = 32'h24822800;
      95690: inst = 32'h10a00000;
      95691: inst = 32'hca00004;
      95692: inst = 32'h38632800;
      95693: inst = 32'h38842800;
      95694: inst = 32'h10a00001;
      95695: inst = 32'hca075d3;
      95696: inst = 32'h13e00001;
      95697: inst = 32'hfe0d96a;
      95698: inst = 32'h5be00000;
      95699: inst = 32'h8c50000;
      95700: inst = 32'h24612800;
      95701: inst = 32'h10a00000;
      95702: inst = 32'hca0000d;
      95703: inst = 32'h24822800;
      95704: inst = 32'h10a00000;
      95705: inst = 32'hca00004;
      95706: inst = 32'h38632800;
      95707: inst = 32'h38842800;
      95708: inst = 32'h10a00001;
      95709: inst = 32'hca075e1;
      95710: inst = 32'h13e00001;
      95711: inst = 32'hfe0d96a;
      95712: inst = 32'h5be00000;
      95713: inst = 32'h8c50000;
      95714: inst = 32'h24612800;
      95715: inst = 32'h10a00000;
      95716: inst = 32'hca0000d;
      95717: inst = 32'h24822800;
      95718: inst = 32'h10a00000;
      95719: inst = 32'hca00004;
      95720: inst = 32'h38632800;
      95721: inst = 32'h38842800;
      95722: inst = 32'h10a00001;
      95723: inst = 32'hca075ef;
      95724: inst = 32'h13e00001;
      95725: inst = 32'hfe0d96a;
      95726: inst = 32'h5be00000;
      95727: inst = 32'h8c50000;
      95728: inst = 32'h24612800;
      95729: inst = 32'h10a00000;
      95730: inst = 32'hca0000d;
      95731: inst = 32'h24822800;
      95732: inst = 32'h10a00000;
      95733: inst = 32'hca00004;
      95734: inst = 32'h38632800;
      95735: inst = 32'h38842800;
      95736: inst = 32'h10a00001;
      95737: inst = 32'hca075fd;
      95738: inst = 32'h13e00001;
      95739: inst = 32'hfe0d96a;
      95740: inst = 32'h5be00000;
      95741: inst = 32'h8c50000;
      95742: inst = 32'h24612800;
      95743: inst = 32'h10a00000;
      95744: inst = 32'hca0000d;
      95745: inst = 32'h24822800;
      95746: inst = 32'h10a00000;
      95747: inst = 32'hca00004;
      95748: inst = 32'h38632800;
      95749: inst = 32'h38842800;
      95750: inst = 32'h10a00001;
      95751: inst = 32'hca0760b;
      95752: inst = 32'h13e00001;
      95753: inst = 32'hfe0d96a;
      95754: inst = 32'h5be00000;
      95755: inst = 32'h8c50000;
      95756: inst = 32'h24612800;
      95757: inst = 32'h10a00000;
      95758: inst = 32'hca0000d;
      95759: inst = 32'h24822800;
      95760: inst = 32'h10a00000;
      95761: inst = 32'hca00004;
      95762: inst = 32'h38632800;
      95763: inst = 32'h38842800;
      95764: inst = 32'h10a00001;
      95765: inst = 32'hca07619;
      95766: inst = 32'h13e00001;
      95767: inst = 32'hfe0d96a;
      95768: inst = 32'h5be00000;
      95769: inst = 32'h8c50000;
      95770: inst = 32'h24612800;
      95771: inst = 32'h10a00000;
      95772: inst = 32'hca0000d;
      95773: inst = 32'h24822800;
      95774: inst = 32'h10a00000;
      95775: inst = 32'hca00004;
      95776: inst = 32'h38632800;
      95777: inst = 32'h38842800;
      95778: inst = 32'h10a00001;
      95779: inst = 32'hca07627;
      95780: inst = 32'h13e00001;
      95781: inst = 32'hfe0d96a;
      95782: inst = 32'h5be00000;
      95783: inst = 32'h8c50000;
      95784: inst = 32'h24612800;
      95785: inst = 32'h10a00000;
      95786: inst = 32'hca0000d;
      95787: inst = 32'h24822800;
      95788: inst = 32'h10a00000;
      95789: inst = 32'hca00004;
      95790: inst = 32'h38632800;
      95791: inst = 32'h38842800;
      95792: inst = 32'h10a00001;
      95793: inst = 32'hca07635;
      95794: inst = 32'h13e00001;
      95795: inst = 32'hfe0d96a;
      95796: inst = 32'h5be00000;
      95797: inst = 32'h8c50000;
      95798: inst = 32'h24612800;
      95799: inst = 32'h10a00000;
      95800: inst = 32'hca0000d;
      95801: inst = 32'h24822800;
      95802: inst = 32'h10a00000;
      95803: inst = 32'hca00004;
      95804: inst = 32'h38632800;
      95805: inst = 32'h38842800;
      95806: inst = 32'h10a00001;
      95807: inst = 32'hca07643;
      95808: inst = 32'h13e00001;
      95809: inst = 32'hfe0d96a;
      95810: inst = 32'h5be00000;
      95811: inst = 32'h8c50000;
      95812: inst = 32'h24612800;
      95813: inst = 32'h10a00000;
      95814: inst = 32'hca0000d;
      95815: inst = 32'h24822800;
      95816: inst = 32'h10a00000;
      95817: inst = 32'hca00004;
      95818: inst = 32'h38632800;
      95819: inst = 32'h38842800;
      95820: inst = 32'h10a00001;
      95821: inst = 32'hca07651;
      95822: inst = 32'h13e00001;
      95823: inst = 32'hfe0d96a;
      95824: inst = 32'h5be00000;
      95825: inst = 32'h8c50000;
      95826: inst = 32'h24612800;
      95827: inst = 32'h10a00000;
      95828: inst = 32'hca0000d;
      95829: inst = 32'h24822800;
      95830: inst = 32'h10a00000;
      95831: inst = 32'hca00004;
      95832: inst = 32'h38632800;
      95833: inst = 32'h38842800;
      95834: inst = 32'h10a00001;
      95835: inst = 32'hca0765f;
      95836: inst = 32'h13e00001;
      95837: inst = 32'hfe0d96a;
      95838: inst = 32'h5be00000;
      95839: inst = 32'h8c50000;
      95840: inst = 32'h24612800;
      95841: inst = 32'h10a00000;
      95842: inst = 32'hca0000d;
      95843: inst = 32'h24822800;
      95844: inst = 32'h10a00000;
      95845: inst = 32'hca00004;
      95846: inst = 32'h38632800;
      95847: inst = 32'h38842800;
      95848: inst = 32'h10a00001;
      95849: inst = 32'hca0766d;
      95850: inst = 32'h13e00001;
      95851: inst = 32'hfe0d96a;
      95852: inst = 32'h5be00000;
      95853: inst = 32'h8c50000;
      95854: inst = 32'h24612800;
      95855: inst = 32'h10a00000;
      95856: inst = 32'hca0000d;
      95857: inst = 32'h24822800;
      95858: inst = 32'h10a00000;
      95859: inst = 32'hca00004;
      95860: inst = 32'h38632800;
      95861: inst = 32'h38842800;
      95862: inst = 32'h10a00001;
      95863: inst = 32'hca0767b;
      95864: inst = 32'h13e00001;
      95865: inst = 32'hfe0d96a;
      95866: inst = 32'h5be00000;
      95867: inst = 32'h8c50000;
      95868: inst = 32'h24612800;
      95869: inst = 32'h10a00000;
      95870: inst = 32'hca0000d;
      95871: inst = 32'h24822800;
      95872: inst = 32'h10a00000;
      95873: inst = 32'hca00004;
      95874: inst = 32'h38632800;
      95875: inst = 32'h38842800;
      95876: inst = 32'h10a00001;
      95877: inst = 32'hca07689;
      95878: inst = 32'h13e00001;
      95879: inst = 32'hfe0d96a;
      95880: inst = 32'h5be00000;
      95881: inst = 32'h8c50000;
      95882: inst = 32'h24612800;
      95883: inst = 32'h10a00000;
      95884: inst = 32'hca0000d;
      95885: inst = 32'h24822800;
      95886: inst = 32'h10a00000;
      95887: inst = 32'hca00004;
      95888: inst = 32'h38632800;
      95889: inst = 32'h38842800;
      95890: inst = 32'h10a00001;
      95891: inst = 32'hca07697;
      95892: inst = 32'h13e00001;
      95893: inst = 32'hfe0d96a;
      95894: inst = 32'h5be00000;
      95895: inst = 32'h8c50000;
      95896: inst = 32'h24612800;
      95897: inst = 32'h10a00000;
      95898: inst = 32'hca0000d;
      95899: inst = 32'h24822800;
      95900: inst = 32'h10a00000;
      95901: inst = 32'hca00004;
      95902: inst = 32'h38632800;
      95903: inst = 32'h38842800;
      95904: inst = 32'h10a00001;
      95905: inst = 32'hca076a5;
      95906: inst = 32'h13e00001;
      95907: inst = 32'hfe0d96a;
      95908: inst = 32'h5be00000;
      95909: inst = 32'h8c50000;
      95910: inst = 32'h24612800;
      95911: inst = 32'h10a00000;
      95912: inst = 32'hca0000d;
      95913: inst = 32'h24822800;
      95914: inst = 32'h10a00000;
      95915: inst = 32'hca00004;
      95916: inst = 32'h38632800;
      95917: inst = 32'h38842800;
      95918: inst = 32'h10a00001;
      95919: inst = 32'hca076b3;
      95920: inst = 32'h13e00001;
      95921: inst = 32'hfe0d96a;
      95922: inst = 32'h5be00000;
      95923: inst = 32'h8c50000;
      95924: inst = 32'h24612800;
      95925: inst = 32'h10a00000;
      95926: inst = 32'hca0000d;
      95927: inst = 32'h24822800;
      95928: inst = 32'h10a00000;
      95929: inst = 32'hca00004;
      95930: inst = 32'h38632800;
      95931: inst = 32'h38842800;
      95932: inst = 32'h10a00001;
      95933: inst = 32'hca076c1;
      95934: inst = 32'h13e00001;
      95935: inst = 32'hfe0d96a;
      95936: inst = 32'h5be00000;
      95937: inst = 32'h8c50000;
      95938: inst = 32'h24612800;
      95939: inst = 32'h10a00000;
      95940: inst = 32'hca0000d;
      95941: inst = 32'h24822800;
      95942: inst = 32'h10a00000;
      95943: inst = 32'hca00004;
      95944: inst = 32'h38632800;
      95945: inst = 32'h38842800;
      95946: inst = 32'h10a00001;
      95947: inst = 32'hca076cf;
      95948: inst = 32'h13e00001;
      95949: inst = 32'hfe0d96a;
      95950: inst = 32'h5be00000;
      95951: inst = 32'h8c50000;
      95952: inst = 32'h24612800;
      95953: inst = 32'h10a00000;
      95954: inst = 32'hca0000d;
      95955: inst = 32'h24822800;
      95956: inst = 32'h10a00000;
      95957: inst = 32'hca00004;
      95958: inst = 32'h38632800;
      95959: inst = 32'h38842800;
      95960: inst = 32'h10a00001;
      95961: inst = 32'hca076dd;
      95962: inst = 32'h13e00001;
      95963: inst = 32'hfe0d96a;
      95964: inst = 32'h5be00000;
      95965: inst = 32'h8c50000;
      95966: inst = 32'h24612800;
      95967: inst = 32'h10a00000;
      95968: inst = 32'hca0000d;
      95969: inst = 32'h24822800;
      95970: inst = 32'h10a00000;
      95971: inst = 32'hca00004;
      95972: inst = 32'h38632800;
      95973: inst = 32'h38842800;
      95974: inst = 32'h10a00001;
      95975: inst = 32'hca076eb;
      95976: inst = 32'h13e00001;
      95977: inst = 32'hfe0d96a;
      95978: inst = 32'h5be00000;
      95979: inst = 32'h8c50000;
      95980: inst = 32'h24612800;
      95981: inst = 32'h10a00000;
      95982: inst = 32'hca0000d;
      95983: inst = 32'h24822800;
      95984: inst = 32'h10a00000;
      95985: inst = 32'hca00004;
      95986: inst = 32'h38632800;
      95987: inst = 32'h38842800;
      95988: inst = 32'h10a00001;
      95989: inst = 32'hca076f9;
      95990: inst = 32'h13e00001;
      95991: inst = 32'hfe0d96a;
      95992: inst = 32'h5be00000;
      95993: inst = 32'h8c50000;
      95994: inst = 32'h24612800;
      95995: inst = 32'h10a00000;
      95996: inst = 32'hca0000d;
      95997: inst = 32'h24822800;
      95998: inst = 32'h10a00000;
      95999: inst = 32'hca00004;
      96000: inst = 32'h38632800;
      96001: inst = 32'h38842800;
      96002: inst = 32'h10a00001;
      96003: inst = 32'hca07707;
      96004: inst = 32'h13e00001;
      96005: inst = 32'hfe0d96a;
      96006: inst = 32'h5be00000;
      96007: inst = 32'h8c50000;
      96008: inst = 32'h24612800;
      96009: inst = 32'h10a00000;
      96010: inst = 32'hca0000d;
      96011: inst = 32'h24822800;
      96012: inst = 32'h10a00000;
      96013: inst = 32'hca00004;
      96014: inst = 32'h38632800;
      96015: inst = 32'h38842800;
      96016: inst = 32'h10a00001;
      96017: inst = 32'hca07715;
      96018: inst = 32'h13e00001;
      96019: inst = 32'hfe0d96a;
      96020: inst = 32'h5be00000;
      96021: inst = 32'h8c50000;
      96022: inst = 32'h24612800;
      96023: inst = 32'h10a00000;
      96024: inst = 32'hca0000d;
      96025: inst = 32'h24822800;
      96026: inst = 32'h10a00000;
      96027: inst = 32'hca00004;
      96028: inst = 32'h38632800;
      96029: inst = 32'h38842800;
      96030: inst = 32'h10a00001;
      96031: inst = 32'hca07723;
      96032: inst = 32'h13e00001;
      96033: inst = 32'hfe0d96a;
      96034: inst = 32'h5be00000;
      96035: inst = 32'h8c50000;
      96036: inst = 32'h24612800;
      96037: inst = 32'h10a00000;
      96038: inst = 32'hca0000d;
      96039: inst = 32'h24822800;
      96040: inst = 32'h10a00000;
      96041: inst = 32'hca00004;
      96042: inst = 32'h38632800;
      96043: inst = 32'h38842800;
      96044: inst = 32'h10a00001;
      96045: inst = 32'hca07731;
      96046: inst = 32'h13e00001;
      96047: inst = 32'hfe0d96a;
      96048: inst = 32'h5be00000;
      96049: inst = 32'h8c50000;
      96050: inst = 32'h24612800;
      96051: inst = 32'h10a00000;
      96052: inst = 32'hca0000d;
      96053: inst = 32'h24822800;
      96054: inst = 32'h10a00000;
      96055: inst = 32'hca00004;
      96056: inst = 32'h38632800;
      96057: inst = 32'h38842800;
      96058: inst = 32'h10a00001;
      96059: inst = 32'hca0773f;
      96060: inst = 32'h13e00001;
      96061: inst = 32'hfe0d96a;
      96062: inst = 32'h5be00000;
      96063: inst = 32'h8c50000;
      96064: inst = 32'h24612800;
      96065: inst = 32'h10a00000;
      96066: inst = 32'hca0000d;
      96067: inst = 32'h24822800;
      96068: inst = 32'h10a00000;
      96069: inst = 32'hca00004;
      96070: inst = 32'h38632800;
      96071: inst = 32'h38842800;
      96072: inst = 32'h10a00001;
      96073: inst = 32'hca0774d;
      96074: inst = 32'h13e00001;
      96075: inst = 32'hfe0d96a;
      96076: inst = 32'h5be00000;
      96077: inst = 32'h8c50000;
      96078: inst = 32'h24612800;
      96079: inst = 32'h10a00000;
      96080: inst = 32'hca0000d;
      96081: inst = 32'h24822800;
      96082: inst = 32'h10a00000;
      96083: inst = 32'hca00004;
      96084: inst = 32'h38632800;
      96085: inst = 32'h38842800;
      96086: inst = 32'h10a00001;
      96087: inst = 32'hca0775b;
      96088: inst = 32'h13e00001;
      96089: inst = 32'hfe0d96a;
      96090: inst = 32'h5be00000;
      96091: inst = 32'h8c50000;
      96092: inst = 32'h24612800;
      96093: inst = 32'h10a00000;
      96094: inst = 32'hca0000d;
      96095: inst = 32'h24822800;
      96096: inst = 32'h10a00000;
      96097: inst = 32'hca00004;
      96098: inst = 32'h38632800;
      96099: inst = 32'h38842800;
      96100: inst = 32'h10a00001;
      96101: inst = 32'hca07769;
      96102: inst = 32'h13e00001;
      96103: inst = 32'hfe0d96a;
      96104: inst = 32'h5be00000;
      96105: inst = 32'h8c50000;
      96106: inst = 32'h24612800;
      96107: inst = 32'h10a00000;
      96108: inst = 32'hca0000d;
      96109: inst = 32'h24822800;
      96110: inst = 32'h10a00000;
      96111: inst = 32'hca00004;
      96112: inst = 32'h38632800;
      96113: inst = 32'h38842800;
      96114: inst = 32'h10a00001;
      96115: inst = 32'hca07777;
      96116: inst = 32'h13e00001;
      96117: inst = 32'hfe0d96a;
      96118: inst = 32'h5be00000;
      96119: inst = 32'h8c50000;
      96120: inst = 32'h24612800;
      96121: inst = 32'h10a00000;
      96122: inst = 32'hca0000d;
      96123: inst = 32'h24822800;
      96124: inst = 32'h10a00000;
      96125: inst = 32'hca00004;
      96126: inst = 32'h38632800;
      96127: inst = 32'h38842800;
      96128: inst = 32'h10a00001;
      96129: inst = 32'hca07785;
      96130: inst = 32'h13e00001;
      96131: inst = 32'hfe0d96a;
      96132: inst = 32'h5be00000;
      96133: inst = 32'h8c50000;
      96134: inst = 32'h24612800;
      96135: inst = 32'h10a00000;
      96136: inst = 32'hca0000d;
      96137: inst = 32'h24822800;
      96138: inst = 32'h10a00000;
      96139: inst = 32'hca00004;
      96140: inst = 32'h38632800;
      96141: inst = 32'h38842800;
      96142: inst = 32'h10a00001;
      96143: inst = 32'hca07793;
      96144: inst = 32'h13e00001;
      96145: inst = 32'hfe0d96a;
      96146: inst = 32'h5be00000;
      96147: inst = 32'h8c50000;
      96148: inst = 32'h24612800;
      96149: inst = 32'h10a00000;
      96150: inst = 32'hca0000d;
      96151: inst = 32'h24822800;
      96152: inst = 32'h10a00000;
      96153: inst = 32'hca00004;
      96154: inst = 32'h38632800;
      96155: inst = 32'h38842800;
      96156: inst = 32'h10a00001;
      96157: inst = 32'hca077a1;
      96158: inst = 32'h13e00001;
      96159: inst = 32'hfe0d96a;
      96160: inst = 32'h5be00000;
      96161: inst = 32'h8c50000;
      96162: inst = 32'h24612800;
      96163: inst = 32'h10a00000;
      96164: inst = 32'hca0000d;
      96165: inst = 32'h24822800;
      96166: inst = 32'h10a00000;
      96167: inst = 32'hca00004;
      96168: inst = 32'h38632800;
      96169: inst = 32'h38842800;
      96170: inst = 32'h10a00001;
      96171: inst = 32'hca077af;
      96172: inst = 32'h13e00001;
      96173: inst = 32'hfe0d96a;
      96174: inst = 32'h5be00000;
      96175: inst = 32'h8c50000;
      96176: inst = 32'h24612800;
      96177: inst = 32'h10a00000;
      96178: inst = 32'hca0000d;
      96179: inst = 32'h24822800;
      96180: inst = 32'h10a00000;
      96181: inst = 32'hca00004;
      96182: inst = 32'h38632800;
      96183: inst = 32'h38842800;
      96184: inst = 32'h10a00001;
      96185: inst = 32'hca077bd;
      96186: inst = 32'h13e00001;
      96187: inst = 32'hfe0d96a;
      96188: inst = 32'h5be00000;
      96189: inst = 32'h8c50000;
      96190: inst = 32'h24612800;
      96191: inst = 32'h10a00000;
      96192: inst = 32'hca0000d;
      96193: inst = 32'h24822800;
      96194: inst = 32'h10a00000;
      96195: inst = 32'hca00004;
      96196: inst = 32'h38632800;
      96197: inst = 32'h38842800;
      96198: inst = 32'h10a00001;
      96199: inst = 32'hca077cb;
      96200: inst = 32'h13e00001;
      96201: inst = 32'hfe0d96a;
      96202: inst = 32'h5be00000;
      96203: inst = 32'h8c50000;
      96204: inst = 32'h24612800;
      96205: inst = 32'h10a00000;
      96206: inst = 32'hca0000d;
      96207: inst = 32'h24822800;
      96208: inst = 32'h10a00000;
      96209: inst = 32'hca00004;
      96210: inst = 32'h38632800;
      96211: inst = 32'h38842800;
      96212: inst = 32'h10a00001;
      96213: inst = 32'hca077d9;
      96214: inst = 32'h13e00001;
      96215: inst = 32'hfe0d96a;
      96216: inst = 32'h5be00000;
      96217: inst = 32'h8c50000;
      96218: inst = 32'h24612800;
      96219: inst = 32'h10a00000;
      96220: inst = 32'hca0000d;
      96221: inst = 32'h24822800;
      96222: inst = 32'h10a00000;
      96223: inst = 32'hca00004;
      96224: inst = 32'h38632800;
      96225: inst = 32'h38842800;
      96226: inst = 32'h10a00001;
      96227: inst = 32'hca077e7;
      96228: inst = 32'h13e00001;
      96229: inst = 32'hfe0d96a;
      96230: inst = 32'h5be00000;
      96231: inst = 32'h8c50000;
      96232: inst = 32'h24612800;
      96233: inst = 32'h10a00000;
      96234: inst = 32'hca0000d;
      96235: inst = 32'h24822800;
      96236: inst = 32'h10a00000;
      96237: inst = 32'hca00004;
      96238: inst = 32'h38632800;
      96239: inst = 32'h38842800;
      96240: inst = 32'h10a00001;
      96241: inst = 32'hca077f5;
      96242: inst = 32'h13e00001;
      96243: inst = 32'hfe0d96a;
      96244: inst = 32'h5be00000;
      96245: inst = 32'h8c50000;
      96246: inst = 32'h24612800;
      96247: inst = 32'h10a00000;
      96248: inst = 32'hca0000d;
      96249: inst = 32'h24822800;
      96250: inst = 32'h10a00000;
      96251: inst = 32'hca00004;
      96252: inst = 32'h38632800;
      96253: inst = 32'h38842800;
      96254: inst = 32'h10a00001;
      96255: inst = 32'hca07803;
      96256: inst = 32'h13e00001;
      96257: inst = 32'hfe0d96a;
      96258: inst = 32'h5be00000;
      96259: inst = 32'h8c50000;
      96260: inst = 32'h24612800;
      96261: inst = 32'h10a00000;
      96262: inst = 32'hca0000d;
      96263: inst = 32'h24822800;
      96264: inst = 32'h10a00000;
      96265: inst = 32'hca00004;
      96266: inst = 32'h38632800;
      96267: inst = 32'h38842800;
      96268: inst = 32'h10a00001;
      96269: inst = 32'hca07811;
      96270: inst = 32'h13e00001;
      96271: inst = 32'hfe0d96a;
      96272: inst = 32'h5be00000;
      96273: inst = 32'h8c50000;
      96274: inst = 32'h24612800;
      96275: inst = 32'h10a00000;
      96276: inst = 32'hca0000d;
      96277: inst = 32'h24822800;
      96278: inst = 32'h10a00000;
      96279: inst = 32'hca00004;
      96280: inst = 32'h38632800;
      96281: inst = 32'h38842800;
      96282: inst = 32'h10a00001;
      96283: inst = 32'hca0781f;
      96284: inst = 32'h13e00001;
      96285: inst = 32'hfe0d96a;
      96286: inst = 32'h5be00000;
      96287: inst = 32'h8c50000;
      96288: inst = 32'h24612800;
      96289: inst = 32'h10a00000;
      96290: inst = 32'hca0000d;
      96291: inst = 32'h24822800;
      96292: inst = 32'h10a00000;
      96293: inst = 32'hca00004;
      96294: inst = 32'h38632800;
      96295: inst = 32'h38842800;
      96296: inst = 32'h10a00001;
      96297: inst = 32'hca0782d;
      96298: inst = 32'h13e00001;
      96299: inst = 32'hfe0d96a;
      96300: inst = 32'h5be00000;
      96301: inst = 32'h8c50000;
      96302: inst = 32'h24612800;
      96303: inst = 32'h10a00000;
      96304: inst = 32'hca0000d;
      96305: inst = 32'h24822800;
      96306: inst = 32'h10a00000;
      96307: inst = 32'hca00004;
      96308: inst = 32'h38632800;
      96309: inst = 32'h38842800;
      96310: inst = 32'h10a00001;
      96311: inst = 32'hca0783b;
      96312: inst = 32'h13e00001;
      96313: inst = 32'hfe0d96a;
      96314: inst = 32'h5be00000;
      96315: inst = 32'h8c50000;
      96316: inst = 32'h24612800;
      96317: inst = 32'h10a00000;
      96318: inst = 32'hca0000d;
      96319: inst = 32'h24822800;
      96320: inst = 32'h10a00000;
      96321: inst = 32'hca00004;
      96322: inst = 32'h38632800;
      96323: inst = 32'h38842800;
      96324: inst = 32'h10a00001;
      96325: inst = 32'hca07849;
      96326: inst = 32'h13e00001;
      96327: inst = 32'hfe0d96a;
      96328: inst = 32'h5be00000;
      96329: inst = 32'h8c50000;
      96330: inst = 32'h24612800;
      96331: inst = 32'h10a00000;
      96332: inst = 32'hca0000d;
      96333: inst = 32'h24822800;
      96334: inst = 32'h10a00000;
      96335: inst = 32'hca00004;
      96336: inst = 32'h38632800;
      96337: inst = 32'h38842800;
      96338: inst = 32'h10a00001;
      96339: inst = 32'hca07857;
      96340: inst = 32'h13e00001;
      96341: inst = 32'hfe0d96a;
      96342: inst = 32'h5be00000;
      96343: inst = 32'h8c50000;
      96344: inst = 32'h24612800;
      96345: inst = 32'h10a00000;
      96346: inst = 32'hca0000d;
      96347: inst = 32'h24822800;
      96348: inst = 32'h10a00000;
      96349: inst = 32'hca00004;
      96350: inst = 32'h38632800;
      96351: inst = 32'h38842800;
      96352: inst = 32'h10a00001;
      96353: inst = 32'hca07865;
      96354: inst = 32'h13e00001;
      96355: inst = 32'hfe0d96a;
      96356: inst = 32'h5be00000;
      96357: inst = 32'h8c50000;
      96358: inst = 32'h24612800;
      96359: inst = 32'h10a00000;
      96360: inst = 32'hca0000d;
      96361: inst = 32'h24822800;
      96362: inst = 32'h10a00000;
      96363: inst = 32'hca00004;
      96364: inst = 32'h38632800;
      96365: inst = 32'h38842800;
      96366: inst = 32'h10a00001;
      96367: inst = 32'hca07873;
      96368: inst = 32'h13e00001;
      96369: inst = 32'hfe0d96a;
      96370: inst = 32'h5be00000;
      96371: inst = 32'h8c50000;
      96372: inst = 32'h24612800;
      96373: inst = 32'h10a00000;
      96374: inst = 32'hca0000d;
      96375: inst = 32'h24822800;
      96376: inst = 32'h10a00000;
      96377: inst = 32'hca00004;
      96378: inst = 32'h38632800;
      96379: inst = 32'h38842800;
      96380: inst = 32'h10a00001;
      96381: inst = 32'hca07881;
      96382: inst = 32'h13e00001;
      96383: inst = 32'hfe0d96a;
      96384: inst = 32'h5be00000;
      96385: inst = 32'h8c50000;
      96386: inst = 32'h24612800;
      96387: inst = 32'h10a00000;
      96388: inst = 32'hca0000d;
      96389: inst = 32'h24822800;
      96390: inst = 32'h10a00000;
      96391: inst = 32'hca00004;
      96392: inst = 32'h38632800;
      96393: inst = 32'h38842800;
      96394: inst = 32'h10a00001;
      96395: inst = 32'hca0788f;
      96396: inst = 32'h13e00001;
      96397: inst = 32'hfe0d96a;
      96398: inst = 32'h5be00000;
      96399: inst = 32'h8c50000;
      96400: inst = 32'h24612800;
      96401: inst = 32'h10a00000;
      96402: inst = 32'hca0000d;
      96403: inst = 32'h24822800;
      96404: inst = 32'h10a00000;
      96405: inst = 32'hca00004;
      96406: inst = 32'h38632800;
      96407: inst = 32'h38842800;
      96408: inst = 32'h10a00001;
      96409: inst = 32'hca0789d;
      96410: inst = 32'h13e00001;
      96411: inst = 32'hfe0d96a;
      96412: inst = 32'h5be00000;
      96413: inst = 32'h8c50000;
      96414: inst = 32'h24612800;
      96415: inst = 32'h10a00000;
      96416: inst = 32'hca0000d;
      96417: inst = 32'h24822800;
      96418: inst = 32'h10a00000;
      96419: inst = 32'hca00004;
      96420: inst = 32'h38632800;
      96421: inst = 32'h38842800;
      96422: inst = 32'h10a00001;
      96423: inst = 32'hca078ab;
      96424: inst = 32'h13e00001;
      96425: inst = 32'hfe0d96a;
      96426: inst = 32'h5be00000;
      96427: inst = 32'h8c50000;
      96428: inst = 32'h24612800;
      96429: inst = 32'h10a00000;
      96430: inst = 32'hca0000d;
      96431: inst = 32'h24822800;
      96432: inst = 32'h10a00000;
      96433: inst = 32'hca00004;
      96434: inst = 32'h38632800;
      96435: inst = 32'h38842800;
      96436: inst = 32'h10a00001;
      96437: inst = 32'hca078b9;
      96438: inst = 32'h13e00001;
      96439: inst = 32'hfe0d96a;
      96440: inst = 32'h5be00000;
      96441: inst = 32'h8c50000;
      96442: inst = 32'h24612800;
      96443: inst = 32'h10a00000;
      96444: inst = 32'hca0000d;
      96445: inst = 32'h24822800;
      96446: inst = 32'h10a00000;
      96447: inst = 32'hca00004;
      96448: inst = 32'h38632800;
      96449: inst = 32'h38842800;
      96450: inst = 32'h10a00001;
      96451: inst = 32'hca078c7;
      96452: inst = 32'h13e00001;
      96453: inst = 32'hfe0d96a;
      96454: inst = 32'h5be00000;
      96455: inst = 32'h8c50000;
      96456: inst = 32'h24612800;
      96457: inst = 32'h10a00000;
      96458: inst = 32'hca0000d;
      96459: inst = 32'h24822800;
      96460: inst = 32'h10a00000;
      96461: inst = 32'hca00004;
      96462: inst = 32'h38632800;
      96463: inst = 32'h38842800;
      96464: inst = 32'h10a00001;
      96465: inst = 32'hca078d5;
      96466: inst = 32'h13e00001;
      96467: inst = 32'hfe0d96a;
      96468: inst = 32'h5be00000;
      96469: inst = 32'h8c50000;
      96470: inst = 32'h24612800;
      96471: inst = 32'h10a00000;
      96472: inst = 32'hca0000d;
      96473: inst = 32'h24822800;
      96474: inst = 32'h10a00000;
      96475: inst = 32'hca00004;
      96476: inst = 32'h38632800;
      96477: inst = 32'h38842800;
      96478: inst = 32'h10a00001;
      96479: inst = 32'hca078e3;
      96480: inst = 32'h13e00001;
      96481: inst = 32'hfe0d96a;
      96482: inst = 32'h5be00000;
      96483: inst = 32'h8c50000;
      96484: inst = 32'h24612800;
      96485: inst = 32'h10a00000;
      96486: inst = 32'hca0000d;
      96487: inst = 32'h24822800;
      96488: inst = 32'h10a00000;
      96489: inst = 32'hca00004;
      96490: inst = 32'h38632800;
      96491: inst = 32'h38842800;
      96492: inst = 32'h10a00001;
      96493: inst = 32'hca078f1;
      96494: inst = 32'h13e00001;
      96495: inst = 32'hfe0d96a;
      96496: inst = 32'h5be00000;
      96497: inst = 32'h8c50000;
      96498: inst = 32'h24612800;
      96499: inst = 32'h10a00000;
      96500: inst = 32'hca0000d;
      96501: inst = 32'h24822800;
      96502: inst = 32'h10a00000;
      96503: inst = 32'hca00004;
      96504: inst = 32'h38632800;
      96505: inst = 32'h38842800;
      96506: inst = 32'h10a00001;
      96507: inst = 32'hca078ff;
      96508: inst = 32'h13e00001;
      96509: inst = 32'hfe0d96a;
      96510: inst = 32'h5be00000;
      96511: inst = 32'h8c50000;
      96512: inst = 32'h24612800;
      96513: inst = 32'h10a00000;
      96514: inst = 32'hca0000d;
      96515: inst = 32'h24822800;
      96516: inst = 32'h10a00000;
      96517: inst = 32'hca00004;
      96518: inst = 32'h38632800;
      96519: inst = 32'h38842800;
      96520: inst = 32'h10a00001;
      96521: inst = 32'hca0790d;
      96522: inst = 32'h13e00001;
      96523: inst = 32'hfe0d96a;
      96524: inst = 32'h5be00000;
      96525: inst = 32'h8c50000;
      96526: inst = 32'h24612800;
      96527: inst = 32'h10a00000;
      96528: inst = 32'hca0000d;
      96529: inst = 32'h24822800;
      96530: inst = 32'h10a00000;
      96531: inst = 32'hca00004;
      96532: inst = 32'h38632800;
      96533: inst = 32'h38842800;
      96534: inst = 32'h10a00001;
      96535: inst = 32'hca0791b;
      96536: inst = 32'h13e00001;
      96537: inst = 32'hfe0d96a;
      96538: inst = 32'h5be00000;
      96539: inst = 32'h8c50000;
      96540: inst = 32'h24612800;
      96541: inst = 32'h10a00000;
      96542: inst = 32'hca0000d;
      96543: inst = 32'h24822800;
      96544: inst = 32'h10a00000;
      96545: inst = 32'hca00004;
      96546: inst = 32'h38632800;
      96547: inst = 32'h38842800;
      96548: inst = 32'h10a00001;
      96549: inst = 32'hca07929;
      96550: inst = 32'h13e00001;
      96551: inst = 32'hfe0d96a;
      96552: inst = 32'h5be00000;
      96553: inst = 32'h8c50000;
      96554: inst = 32'h24612800;
      96555: inst = 32'h10a00000;
      96556: inst = 32'hca0000d;
      96557: inst = 32'h24822800;
      96558: inst = 32'h10a00000;
      96559: inst = 32'hca00004;
      96560: inst = 32'h38632800;
      96561: inst = 32'h38842800;
      96562: inst = 32'h10a00001;
      96563: inst = 32'hca07937;
      96564: inst = 32'h13e00001;
      96565: inst = 32'hfe0d96a;
      96566: inst = 32'h5be00000;
      96567: inst = 32'h8c50000;
      96568: inst = 32'h24612800;
      96569: inst = 32'h10a00000;
      96570: inst = 32'hca0000d;
      96571: inst = 32'h24822800;
      96572: inst = 32'h10a00000;
      96573: inst = 32'hca00004;
      96574: inst = 32'h38632800;
      96575: inst = 32'h38842800;
      96576: inst = 32'h10a00001;
      96577: inst = 32'hca07945;
      96578: inst = 32'h13e00001;
      96579: inst = 32'hfe0d96a;
      96580: inst = 32'h5be00000;
      96581: inst = 32'h8c50000;
      96582: inst = 32'h24612800;
      96583: inst = 32'h10a00000;
      96584: inst = 32'hca0000d;
      96585: inst = 32'h24822800;
      96586: inst = 32'h10a00000;
      96587: inst = 32'hca00004;
      96588: inst = 32'h38632800;
      96589: inst = 32'h38842800;
      96590: inst = 32'h10a00001;
      96591: inst = 32'hca07953;
      96592: inst = 32'h13e00001;
      96593: inst = 32'hfe0d96a;
      96594: inst = 32'h5be00000;
      96595: inst = 32'h8c50000;
      96596: inst = 32'h24612800;
      96597: inst = 32'h10a00000;
      96598: inst = 32'hca0000d;
      96599: inst = 32'h24822800;
      96600: inst = 32'h10a00000;
      96601: inst = 32'hca00004;
      96602: inst = 32'h38632800;
      96603: inst = 32'h38842800;
      96604: inst = 32'h10a00001;
      96605: inst = 32'hca07961;
      96606: inst = 32'h13e00001;
      96607: inst = 32'hfe0d96a;
      96608: inst = 32'h5be00000;
      96609: inst = 32'h8c50000;
      96610: inst = 32'h24612800;
      96611: inst = 32'h10a00000;
      96612: inst = 32'hca0000d;
      96613: inst = 32'h24822800;
      96614: inst = 32'h10a00000;
      96615: inst = 32'hca00004;
      96616: inst = 32'h38632800;
      96617: inst = 32'h38842800;
      96618: inst = 32'h10a00001;
      96619: inst = 32'hca0796f;
      96620: inst = 32'h13e00001;
      96621: inst = 32'hfe0d96a;
      96622: inst = 32'h5be00000;
      96623: inst = 32'h8c50000;
      96624: inst = 32'h24612800;
      96625: inst = 32'h10a00000;
      96626: inst = 32'hca0000d;
      96627: inst = 32'h24822800;
      96628: inst = 32'h10a00000;
      96629: inst = 32'hca00004;
      96630: inst = 32'h38632800;
      96631: inst = 32'h38842800;
      96632: inst = 32'h10a00001;
      96633: inst = 32'hca0797d;
      96634: inst = 32'h13e00001;
      96635: inst = 32'hfe0d96a;
      96636: inst = 32'h5be00000;
      96637: inst = 32'h8c50000;
      96638: inst = 32'h24612800;
      96639: inst = 32'h10a00000;
      96640: inst = 32'hca0000d;
      96641: inst = 32'h24822800;
      96642: inst = 32'h10a00000;
      96643: inst = 32'hca00004;
      96644: inst = 32'h38632800;
      96645: inst = 32'h38842800;
      96646: inst = 32'h10a00001;
      96647: inst = 32'hca0798b;
      96648: inst = 32'h13e00001;
      96649: inst = 32'hfe0d96a;
      96650: inst = 32'h5be00000;
      96651: inst = 32'h8c50000;
      96652: inst = 32'h24612800;
      96653: inst = 32'h10a00000;
      96654: inst = 32'hca0000d;
      96655: inst = 32'h24822800;
      96656: inst = 32'h10a00000;
      96657: inst = 32'hca00004;
      96658: inst = 32'h38632800;
      96659: inst = 32'h38842800;
      96660: inst = 32'h10a00001;
      96661: inst = 32'hca07999;
      96662: inst = 32'h13e00001;
      96663: inst = 32'hfe0d96a;
      96664: inst = 32'h5be00000;
      96665: inst = 32'h8c50000;
      96666: inst = 32'h24612800;
      96667: inst = 32'h10a00000;
      96668: inst = 32'hca0000d;
      96669: inst = 32'h24822800;
      96670: inst = 32'h10a00000;
      96671: inst = 32'hca00004;
      96672: inst = 32'h38632800;
      96673: inst = 32'h38842800;
      96674: inst = 32'h10a00001;
      96675: inst = 32'hca079a7;
      96676: inst = 32'h13e00001;
      96677: inst = 32'hfe0d96a;
      96678: inst = 32'h5be00000;
      96679: inst = 32'h8c50000;
      96680: inst = 32'h24612800;
      96681: inst = 32'h10a00000;
      96682: inst = 32'hca0000d;
      96683: inst = 32'h24822800;
      96684: inst = 32'h10a00000;
      96685: inst = 32'hca00004;
      96686: inst = 32'h38632800;
      96687: inst = 32'h38842800;
      96688: inst = 32'h10a00001;
      96689: inst = 32'hca079b5;
      96690: inst = 32'h13e00001;
      96691: inst = 32'hfe0d96a;
      96692: inst = 32'h5be00000;
      96693: inst = 32'h8c50000;
      96694: inst = 32'h24612800;
      96695: inst = 32'h10a00000;
      96696: inst = 32'hca0000d;
      96697: inst = 32'h24822800;
      96698: inst = 32'h10a00000;
      96699: inst = 32'hca00004;
      96700: inst = 32'h38632800;
      96701: inst = 32'h38842800;
      96702: inst = 32'h10a00001;
      96703: inst = 32'hca079c3;
      96704: inst = 32'h13e00001;
      96705: inst = 32'hfe0d96a;
      96706: inst = 32'h5be00000;
      96707: inst = 32'h8c50000;
      96708: inst = 32'h24612800;
      96709: inst = 32'h10a00000;
      96710: inst = 32'hca0000d;
      96711: inst = 32'h24822800;
      96712: inst = 32'h10a00000;
      96713: inst = 32'hca00004;
      96714: inst = 32'h38632800;
      96715: inst = 32'h38842800;
      96716: inst = 32'h10a00001;
      96717: inst = 32'hca079d1;
      96718: inst = 32'h13e00001;
      96719: inst = 32'hfe0d96a;
      96720: inst = 32'h5be00000;
      96721: inst = 32'h8c50000;
      96722: inst = 32'h24612800;
      96723: inst = 32'h10a00000;
      96724: inst = 32'hca0000d;
      96725: inst = 32'h24822800;
      96726: inst = 32'h10a00000;
      96727: inst = 32'hca00004;
      96728: inst = 32'h38632800;
      96729: inst = 32'h38842800;
      96730: inst = 32'h10a00001;
      96731: inst = 32'hca079df;
      96732: inst = 32'h13e00001;
      96733: inst = 32'hfe0d96a;
      96734: inst = 32'h5be00000;
      96735: inst = 32'h8c50000;
      96736: inst = 32'h24612800;
      96737: inst = 32'h10a00000;
      96738: inst = 32'hca0000d;
      96739: inst = 32'h24822800;
      96740: inst = 32'h10a00000;
      96741: inst = 32'hca00004;
      96742: inst = 32'h38632800;
      96743: inst = 32'h38842800;
      96744: inst = 32'h10a00001;
      96745: inst = 32'hca079ed;
      96746: inst = 32'h13e00001;
      96747: inst = 32'hfe0d96a;
      96748: inst = 32'h5be00000;
      96749: inst = 32'h8c50000;
      96750: inst = 32'h24612800;
      96751: inst = 32'h10a00000;
      96752: inst = 32'hca0000d;
      96753: inst = 32'h24822800;
      96754: inst = 32'h10a00000;
      96755: inst = 32'hca00004;
      96756: inst = 32'h38632800;
      96757: inst = 32'h38842800;
      96758: inst = 32'h10a00001;
      96759: inst = 32'hca079fb;
      96760: inst = 32'h13e00001;
      96761: inst = 32'hfe0d96a;
      96762: inst = 32'h5be00000;
      96763: inst = 32'h8c50000;
      96764: inst = 32'h24612800;
      96765: inst = 32'h10a00000;
      96766: inst = 32'hca0000d;
      96767: inst = 32'h24822800;
      96768: inst = 32'h10a00000;
      96769: inst = 32'hca00004;
      96770: inst = 32'h38632800;
      96771: inst = 32'h38842800;
      96772: inst = 32'h10a00001;
      96773: inst = 32'hca07a09;
      96774: inst = 32'h13e00001;
      96775: inst = 32'hfe0d96a;
      96776: inst = 32'h5be00000;
      96777: inst = 32'h8c50000;
      96778: inst = 32'h24612800;
      96779: inst = 32'h10a00000;
      96780: inst = 32'hca0000d;
      96781: inst = 32'h24822800;
      96782: inst = 32'h10a00000;
      96783: inst = 32'hca00004;
      96784: inst = 32'h38632800;
      96785: inst = 32'h38842800;
      96786: inst = 32'h10a00001;
      96787: inst = 32'hca07a17;
      96788: inst = 32'h13e00001;
      96789: inst = 32'hfe0d96a;
      96790: inst = 32'h5be00000;
      96791: inst = 32'h8c50000;
      96792: inst = 32'h24612800;
      96793: inst = 32'h10a00000;
      96794: inst = 32'hca0000d;
      96795: inst = 32'h24822800;
      96796: inst = 32'h10a00000;
      96797: inst = 32'hca00004;
      96798: inst = 32'h38632800;
      96799: inst = 32'h38842800;
      96800: inst = 32'h10a00001;
      96801: inst = 32'hca07a25;
      96802: inst = 32'h13e00001;
      96803: inst = 32'hfe0d96a;
      96804: inst = 32'h5be00000;
      96805: inst = 32'h8c50000;
      96806: inst = 32'h24612800;
      96807: inst = 32'h10a00000;
      96808: inst = 32'hca0000d;
      96809: inst = 32'h24822800;
      96810: inst = 32'h10a00000;
      96811: inst = 32'hca00004;
      96812: inst = 32'h38632800;
      96813: inst = 32'h38842800;
      96814: inst = 32'h10a00001;
      96815: inst = 32'hca07a33;
      96816: inst = 32'h13e00001;
      96817: inst = 32'hfe0d96a;
      96818: inst = 32'h5be00000;
      96819: inst = 32'h8c50000;
      96820: inst = 32'h24612800;
      96821: inst = 32'h10a00000;
      96822: inst = 32'hca0000d;
      96823: inst = 32'h24822800;
      96824: inst = 32'h10a00000;
      96825: inst = 32'hca00004;
      96826: inst = 32'h38632800;
      96827: inst = 32'h38842800;
      96828: inst = 32'h10a00001;
      96829: inst = 32'hca07a41;
      96830: inst = 32'h13e00001;
      96831: inst = 32'hfe0d96a;
      96832: inst = 32'h5be00000;
      96833: inst = 32'h8c50000;
      96834: inst = 32'h24612800;
      96835: inst = 32'h10a00000;
      96836: inst = 32'hca0000d;
      96837: inst = 32'h24822800;
      96838: inst = 32'h10a00000;
      96839: inst = 32'hca00004;
      96840: inst = 32'h38632800;
      96841: inst = 32'h38842800;
      96842: inst = 32'h10a00001;
      96843: inst = 32'hca07a4f;
      96844: inst = 32'h13e00001;
      96845: inst = 32'hfe0d96a;
      96846: inst = 32'h5be00000;
      96847: inst = 32'h8c50000;
      96848: inst = 32'h24612800;
      96849: inst = 32'h10a00000;
      96850: inst = 32'hca0000d;
      96851: inst = 32'h24822800;
      96852: inst = 32'h10a00000;
      96853: inst = 32'hca00004;
      96854: inst = 32'h38632800;
      96855: inst = 32'h38842800;
      96856: inst = 32'h10a00001;
      96857: inst = 32'hca07a5d;
      96858: inst = 32'h13e00001;
      96859: inst = 32'hfe0d96a;
      96860: inst = 32'h5be00000;
      96861: inst = 32'h8c50000;
      96862: inst = 32'h24612800;
      96863: inst = 32'h10a00000;
      96864: inst = 32'hca0000d;
      96865: inst = 32'h24822800;
      96866: inst = 32'h10a00000;
      96867: inst = 32'hca00004;
      96868: inst = 32'h38632800;
      96869: inst = 32'h38842800;
      96870: inst = 32'h10a00001;
      96871: inst = 32'hca07a6b;
      96872: inst = 32'h13e00001;
      96873: inst = 32'hfe0d96a;
      96874: inst = 32'h5be00000;
      96875: inst = 32'h8c50000;
      96876: inst = 32'h24612800;
      96877: inst = 32'h10a00000;
      96878: inst = 32'hca0000d;
      96879: inst = 32'h24822800;
      96880: inst = 32'h10a00000;
      96881: inst = 32'hca00004;
      96882: inst = 32'h38632800;
      96883: inst = 32'h38842800;
      96884: inst = 32'h10a00001;
      96885: inst = 32'hca07a79;
      96886: inst = 32'h13e00001;
      96887: inst = 32'hfe0d96a;
      96888: inst = 32'h5be00000;
      96889: inst = 32'h8c50000;
      96890: inst = 32'h24612800;
      96891: inst = 32'h10a00000;
      96892: inst = 32'hca0000d;
      96893: inst = 32'h24822800;
      96894: inst = 32'h10a00000;
      96895: inst = 32'hca00004;
      96896: inst = 32'h38632800;
      96897: inst = 32'h38842800;
      96898: inst = 32'h10a00001;
      96899: inst = 32'hca07a87;
      96900: inst = 32'h13e00001;
      96901: inst = 32'hfe0d96a;
      96902: inst = 32'h5be00000;
      96903: inst = 32'h8c50000;
      96904: inst = 32'h24612800;
      96905: inst = 32'h10a00000;
      96906: inst = 32'hca0000d;
      96907: inst = 32'h24822800;
      96908: inst = 32'h10a00000;
      96909: inst = 32'hca00004;
      96910: inst = 32'h38632800;
      96911: inst = 32'h38842800;
      96912: inst = 32'h10a00001;
      96913: inst = 32'hca07a95;
      96914: inst = 32'h13e00001;
      96915: inst = 32'hfe0d96a;
      96916: inst = 32'h5be00000;
      96917: inst = 32'h8c50000;
      96918: inst = 32'h24612800;
      96919: inst = 32'h10a00000;
      96920: inst = 32'hca0000d;
      96921: inst = 32'h24822800;
      96922: inst = 32'h10a00000;
      96923: inst = 32'hca00004;
      96924: inst = 32'h38632800;
      96925: inst = 32'h38842800;
      96926: inst = 32'h10a00001;
      96927: inst = 32'hca07aa3;
      96928: inst = 32'h13e00001;
      96929: inst = 32'hfe0d96a;
      96930: inst = 32'h5be00000;
      96931: inst = 32'h8c50000;
      96932: inst = 32'h24612800;
      96933: inst = 32'h10a00000;
      96934: inst = 32'hca0000d;
      96935: inst = 32'h24822800;
      96936: inst = 32'h10a00000;
      96937: inst = 32'hca00004;
      96938: inst = 32'h38632800;
      96939: inst = 32'h38842800;
      96940: inst = 32'h10a00001;
      96941: inst = 32'hca07ab1;
      96942: inst = 32'h13e00001;
      96943: inst = 32'hfe0d96a;
      96944: inst = 32'h5be00000;
      96945: inst = 32'h8c50000;
      96946: inst = 32'h24612800;
      96947: inst = 32'h10a00000;
      96948: inst = 32'hca0000d;
      96949: inst = 32'h24822800;
      96950: inst = 32'h10a00000;
      96951: inst = 32'hca00004;
      96952: inst = 32'h38632800;
      96953: inst = 32'h38842800;
      96954: inst = 32'h10a00001;
      96955: inst = 32'hca07abf;
      96956: inst = 32'h13e00001;
      96957: inst = 32'hfe0d96a;
      96958: inst = 32'h5be00000;
      96959: inst = 32'h8c50000;
      96960: inst = 32'h24612800;
      96961: inst = 32'h10a00000;
      96962: inst = 32'hca0000d;
      96963: inst = 32'h24822800;
      96964: inst = 32'h10a00000;
      96965: inst = 32'hca00004;
      96966: inst = 32'h38632800;
      96967: inst = 32'h38842800;
      96968: inst = 32'h10a00001;
      96969: inst = 32'hca07acd;
      96970: inst = 32'h13e00001;
      96971: inst = 32'hfe0d96a;
      96972: inst = 32'h5be00000;
      96973: inst = 32'h8c50000;
      96974: inst = 32'h24612800;
      96975: inst = 32'h10a00000;
      96976: inst = 32'hca0000d;
      96977: inst = 32'h24822800;
      96978: inst = 32'h10a00000;
      96979: inst = 32'hca00004;
      96980: inst = 32'h38632800;
      96981: inst = 32'h38842800;
      96982: inst = 32'h10a00001;
      96983: inst = 32'hca07adb;
      96984: inst = 32'h13e00001;
      96985: inst = 32'hfe0d96a;
      96986: inst = 32'h5be00000;
      96987: inst = 32'h8c50000;
      96988: inst = 32'h24612800;
      96989: inst = 32'h10a00000;
      96990: inst = 32'hca0000d;
      96991: inst = 32'h24822800;
      96992: inst = 32'h10a00000;
      96993: inst = 32'hca00004;
      96994: inst = 32'h38632800;
      96995: inst = 32'h38842800;
      96996: inst = 32'h10a00001;
      96997: inst = 32'hca07ae9;
      96998: inst = 32'h13e00001;
      96999: inst = 32'hfe0d96a;
      97000: inst = 32'h5be00000;
      97001: inst = 32'h8c50000;
      97002: inst = 32'h24612800;
      97003: inst = 32'h10a00000;
      97004: inst = 32'hca0000e;
      97005: inst = 32'h24822800;
      97006: inst = 32'h10a00000;
      97007: inst = 32'hca00004;
      97008: inst = 32'h38632800;
      97009: inst = 32'h38842800;
      97010: inst = 32'h10a00001;
      97011: inst = 32'hca07af7;
      97012: inst = 32'h13e00001;
      97013: inst = 32'hfe0d96a;
      97014: inst = 32'h5be00000;
      97015: inst = 32'h8c50000;
      97016: inst = 32'h24612800;
      97017: inst = 32'h10a00000;
      97018: inst = 32'hca0000e;
      97019: inst = 32'h24822800;
      97020: inst = 32'h10a00000;
      97021: inst = 32'hca00004;
      97022: inst = 32'h38632800;
      97023: inst = 32'h38842800;
      97024: inst = 32'h10a00001;
      97025: inst = 32'hca07b05;
      97026: inst = 32'h13e00001;
      97027: inst = 32'hfe0d96a;
      97028: inst = 32'h5be00000;
      97029: inst = 32'h8c50000;
      97030: inst = 32'h24612800;
      97031: inst = 32'h10a00000;
      97032: inst = 32'hca0000e;
      97033: inst = 32'h24822800;
      97034: inst = 32'h10a00000;
      97035: inst = 32'hca00004;
      97036: inst = 32'h38632800;
      97037: inst = 32'h38842800;
      97038: inst = 32'h10a00001;
      97039: inst = 32'hca07b13;
      97040: inst = 32'h13e00001;
      97041: inst = 32'hfe0d96a;
      97042: inst = 32'h5be00000;
      97043: inst = 32'h8c50000;
      97044: inst = 32'h24612800;
      97045: inst = 32'h10a00000;
      97046: inst = 32'hca0000e;
      97047: inst = 32'h24822800;
      97048: inst = 32'h10a00000;
      97049: inst = 32'hca00004;
      97050: inst = 32'h38632800;
      97051: inst = 32'h38842800;
      97052: inst = 32'h10a00001;
      97053: inst = 32'hca07b21;
      97054: inst = 32'h13e00001;
      97055: inst = 32'hfe0d96a;
      97056: inst = 32'h5be00000;
      97057: inst = 32'h8c50000;
      97058: inst = 32'h24612800;
      97059: inst = 32'h10a00000;
      97060: inst = 32'hca0000e;
      97061: inst = 32'h24822800;
      97062: inst = 32'h10a00000;
      97063: inst = 32'hca00004;
      97064: inst = 32'h38632800;
      97065: inst = 32'h38842800;
      97066: inst = 32'h10a00001;
      97067: inst = 32'hca07b2f;
      97068: inst = 32'h13e00001;
      97069: inst = 32'hfe0d96a;
      97070: inst = 32'h5be00000;
      97071: inst = 32'h8c50000;
      97072: inst = 32'h24612800;
      97073: inst = 32'h10a00000;
      97074: inst = 32'hca0000e;
      97075: inst = 32'h24822800;
      97076: inst = 32'h10a00000;
      97077: inst = 32'hca00004;
      97078: inst = 32'h38632800;
      97079: inst = 32'h38842800;
      97080: inst = 32'h10a00001;
      97081: inst = 32'hca07b3d;
      97082: inst = 32'h13e00001;
      97083: inst = 32'hfe0d96a;
      97084: inst = 32'h5be00000;
      97085: inst = 32'h8c50000;
      97086: inst = 32'h24612800;
      97087: inst = 32'h10a00000;
      97088: inst = 32'hca0000e;
      97089: inst = 32'h24822800;
      97090: inst = 32'h10a00000;
      97091: inst = 32'hca00004;
      97092: inst = 32'h38632800;
      97093: inst = 32'h38842800;
      97094: inst = 32'h10a00001;
      97095: inst = 32'hca07b4b;
      97096: inst = 32'h13e00001;
      97097: inst = 32'hfe0d96a;
      97098: inst = 32'h5be00000;
      97099: inst = 32'h8c50000;
      97100: inst = 32'h24612800;
      97101: inst = 32'h10a00000;
      97102: inst = 32'hca0000e;
      97103: inst = 32'h24822800;
      97104: inst = 32'h10a00000;
      97105: inst = 32'hca00004;
      97106: inst = 32'h38632800;
      97107: inst = 32'h38842800;
      97108: inst = 32'h10a00001;
      97109: inst = 32'hca07b59;
      97110: inst = 32'h13e00001;
      97111: inst = 32'hfe0d96a;
      97112: inst = 32'h5be00000;
      97113: inst = 32'h8c50000;
      97114: inst = 32'h24612800;
      97115: inst = 32'h10a00000;
      97116: inst = 32'hca0000e;
      97117: inst = 32'h24822800;
      97118: inst = 32'h10a00000;
      97119: inst = 32'hca00004;
      97120: inst = 32'h38632800;
      97121: inst = 32'h38842800;
      97122: inst = 32'h10a00001;
      97123: inst = 32'hca07b67;
      97124: inst = 32'h13e00001;
      97125: inst = 32'hfe0d96a;
      97126: inst = 32'h5be00000;
      97127: inst = 32'h8c50000;
      97128: inst = 32'h24612800;
      97129: inst = 32'h10a00000;
      97130: inst = 32'hca0000e;
      97131: inst = 32'h24822800;
      97132: inst = 32'h10a00000;
      97133: inst = 32'hca00004;
      97134: inst = 32'h38632800;
      97135: inst = 32'h38842800;
      97136: inst = 32'h10a00001;
      97137: inst = 32'hca07b75;
      97138: inst = 32'h13e00001;
      97139: inst = 32'hfe0d96a;
      97140: inst = 32'h5be00000;
      97141: inst = 32'h8c50000;
      97142: inst = 32'h24612800;
      97143: inst = 32'h10a00000;
      97144: inst = 32'hca0000e;
      97145: inst = 32'h24822800;
      97146: inst = 32'h10a00000;
      97147: inst = 32'hca00004;
      97148: inst = 32'h38632800;
      97149: inst = 32'h38842800;
      97150: inst = 32'h10a00001;
      97151: inst = 32'hca07b83;
      97152: inst = 32'h13e00001;
      97153: inst = 32'hfe0d96a;
      97154: inst = 32'h5be00000;
      97155: inst = 32'h8c50000;
      97156: inst = 32'h24612800;
      97157: inst = 32'h10a00000;
      97158: inst = 32'hca0000e;
      97159: inst = 32'h24822800;
      97160: inst = 32'h10a00000;
      97161: inst = 32'hca00004;
      97162: inst = 32'h38632800;
      97163: inst = 32'h38842800;
      97164: inst = 32'h10a00001;
      97165: inst = 32'hca07b91;
      97166: inst = 32'h13e00001;
      97167: inst = 32'hfe0d96a;
      97168: inst = 32'h5be00000;
      97169: inst = 32'h8c50000;
      97170: inst = 32'h24612800;
      97171: inst = 32'h10a00000;
      97172: inst = 32'hca0000e;
      97173: inst = 32'h24822800;
      97174: inst = 32'h10a00000;
      97175: inst = 32'hca00004;
      97176: inst = 32'h38632800;
      97177: inst = 32'h38842800;
      97178: inst = 32'h10a00001;
      97179: inst = 32'hca07b9f;
      97180: inst = 32'h13e00001;
      97181: inst = 32'hfe0d96a;
      97182: inst = 32'h5be00000;
      97183: inst = 32'h8c50000;
      97184: inst = 32'h24612800;
      97185: inst = 32'h10a00000;
      97186: inst = 32'hca0000e;
      97187: inst = 32'h24822800;
      97188: inst = 32'h10a00000;
      97189: inst = 32'hca00004;
      97190: inst = 32'h38632800;
      97191: inst = 32'h38842800;
      97192: inst = 32'h10a00001;
      97193: inst = 32'hca07bad;
      97194: inst = 32'h13e00001;
      97195: inst = 32'hfe0d96a;
      97196: inst = 32'h5be00000;
      97197: inst = 32'h8c50000;
      97198: inst = 32'h24612800;
      97199: inst = 32'h10a00000;
      97200: inst = 32'hca0000e;
      97201: inst = 32'h24822800;
      97202: inst = 32'h10a00000;
      97203: inst = 32'hca00004;
      97204: inst = 32'h38632800;
      97205: inst = 32'h38842800;
      97206: inst = 32'h10a00001;
      97207: inst = 32'hca07bbb;
      97208: inst = 32'h13e00001;
      97209: inst = 32'hfe0d96a;
      97210: inst = 32'h5be00000;
      97211: inst = 32'h8c50000;
      97212: inst = 32'h24612800;
      97213: inst = 32'h10a00000;
      97214: inst = 32'hca0000e;
      97215: inst = 32'h24822800;
      97216: inst = 32'h10a00000;
      97217: inst = 32'hca00004;
      97218: inst = 32'h38632800;
      97219: inst = 32'h38842800;
      97220: inst = 32'h10a00001;
      97221: inst = 32'hca07bc9;
      97222: inst = 32'h13e00001;
      97223: inst = 32'hfe0d96a;
      97224: inst = 32'h5be00000;
      97225: inst = 32'h8c50000;
      97226: inst = 32'h24612800;
      97227: inst = 32'h10a00000;
      97228: inst = 32'hca0000e;
      97229: inst = 32'h24822800;
      97230: inst = 32'h10a00000;
      97231: inst = 32'hca00004;
      97232: inst = 32'h38632800;
      97233: inst = 32'h38842800;
      97234: inst = 32'h10a00001;
      97235: inst = 32'hca07bd7;
      97236: inst = 32'h13e00001;
      97237: inst = 32'hfe0d96a;
      97238: inst = 32'h5be00000;
      97239: inst = 32'h8c50000;
      97240: inst = 32'h24612800;
      97241: inst = 32'h10a00000;
      97242: inst = 32'hca0000e;
      97243: inst = 32'h24822800;
      97244: inst = 32'h10a00000;
      97245: inst = 32'hca00004;
      97246: inst = 32'h38632800;
      97247: inst = 32'h38842800;
      97248: inst = 32'h10a00001;
      97249: inst = 32'hca07be5;
      97250: inst = 32'h13e00001;
      97251: inst = 32'hfe0d96a;
      97252: inst = 32'h5be00000;
      97253: inst = 32'h8c50000;
      97254: inst = 32'h24612800;
      97255: inst = 32'h10a00000;
      97256: inst = 32'hca0000e;
      97257: inst = 32'h24822800;
      97258: inst = 32'h10a00000;
      97259: inst = 32'hca00004;
      97260: inst = 32'h38632800;
      97261: inst = 32'h38842800;
      97262: inst = 32'h10a00001;
      97263: inst = 32'hca07bf3;
      97264: inst = 32'h13e00001;
      97265: inst = 32'hfe0d96a;
      97266: inst = 32'h5be00000;
      97267: inst = 32'h8c50000;
      97268: inst = 32'h24612800;
      97269: inst = 32'h10a00000;
      97270: inst = 32'hca0000e;
      97271: inst = 32'h24822800;
      97272: inst = 32'h10a00000;
      97273: inst = 32'hca00004;
      97274: inst = 32'h38632800;
      97275: inst = 32'h38842800;
      97276: inst = 32'h10a00001;
      97277: inst = 32'hca07c01;
      97278: inst = 32'h13e00001;
      97279: inst = 32'hfe0d96a;
      97280: inst = 32'h5be00000;
      97281: inst = 32'h8c50000;
      97282: inst = 32'h24612800;
      97283: inst = 32'h10a00000;
      97284: inst = 32'hca0000e;
      97285: inst = 32'h24822800;
      97286: inst = 32'h10a00000;
      97287: inst = 32'hca00004;
      97288: inst = 32'h38632800;
      97289: inst = 32'h38842800;
      97290: inst = 32'h10a00001;
      97291: inst = 32'hca07c0f;
      97292: inst = 32'h13e00001;
      97293: inst = 32'hfe0d96a;
      97294: inst = 32'h5be00000;
      97295: inst = 32'h8c50000;
      97296: inst = 32'h24612800;
      97297: inst = 32'h10a00000;
      97298: inst = 32'hca0000e;
      97299: inst = 32'h24822800;
      97300: inst = 32'h10a00000;
      97301: inst = 32'hca00004;
      97302: inst = 32'h38632800;
      97303: inst = 32'h38842800;
      97304: inst = 32'h10a00001;
      97305: inst = 32'hca07c1d;
      97306: inst = 32'h13e00001;
      97307: inst = 32'hfe0d96a;
      97308: inst = 32'h5be00000;
      97309: inst = 32'h8c50000;
      97310: inst = 32'h24612800;
      97311: inst = 32'h10a00000;
      97312: inst = 32'hca0000e;
      97313: inst = 32'h24822800;
      97314: inst = 32'h10a00000;
      97315: inst = 32'hca00004;
      97316: inst = 32'h38632800;
      97317: inst = 32'h38842800;
      97318: inst = 32'h10a00001;
      97319: inst = 32'hca07c2b;
      97320: inst = 32'h13e00001;
      97321: inst = 32'hfe0d96a;
      97322: inst = 32'h5be00000;
      97323: inst = 32'h8c50000;
      97324: inst = 32'h24612800;
      97325: inst = 32'h10a00000;
      97326: inst = 32'hca0000e;
      97327: inst = 32'h24822800;
      97328: inst = 32'h10a00000;
      97329: inst = 32'hca00004;
      97330: inst = 32'h38632800;
      97331: inst = 32'h38842800;
      97332: inst = 32'h10a00001;
      97333: inst = 32'hca07c39;
      97334: inst = 32'h13e00001;
      97335: inst = 32'hfe0d96a;
      97336: inst = 32'h5be00000;
      97337: inst = 32'h8c50000;
      97338: inst = 32'h24612800;
      97339: inst = 32'h10a00000;
      97340: inst = 32'hca0000e;
      97341: inst = 32'h24822800;
      97342: inst = 32'h10a00000;
      97343: inst = 32'hca00004;
      97344: inst = 32'h38632800;
      97345: inst = 32'h38842800;
      97346: inst = 32'h10a00001;
      97347: inst = 32'hca07c47;
      97348: inst = 32'h13e00001;
      97349: inst = 32'hfe0d96a;
      97350: inst = 32'h5be00000;
      97351: inst = 32'h8c50000;
      97352: inst = 32'h24612800;
      97353: inst = 32'h10a00000;
      97354: inst = 32'hca0000e;
      97355: inst = 32'h24822800;
      97356: inst = 32'h10a00000;
      97357: inst = 32'hca00004;
      97358: inst = 32'h38632800;
      97359: inst = 32'h38842800;
      97360: inst = 32'h10a00001;
      97361: inst = 32'hca07c55;
      97362: inst = 32'h13e00001;
      97363: inst = 32'hfe0d96a;
      97364: inst = 32'h5be00000;
      97365: inst = 32'h8c50000;
      97366: inst = 32'h24612800;
      97367: inst = 32'h10a00000;
      97368: inst = 32'hca0000e;
      97369: inst = 32'h24822800;
      97370: inst = 32'h10a00000;
      97371: inst = 32'hca00004;
      97372: inst = 32'h38632800;
      97373: inst = 32'h38842800;
      97374: inst = 32'h10a00001;
      97375: inst = 32'hca07c63;
      97376: inst = 32'h13e00001;
      97377: inst = 32'hfe0d96a;
      97378: inst = 32'h5be00000;
      97379: inst = 32'h8c50000;
      97380: inst = 32'h24612800;
      97381: inst = 32'h10a00000;
      97382: inst = 32'hca0000e;
      97383: inst = 32'h24822800;
      97384: inst = 32'h10a00000;
      97385: inst = 32'hca00004;
      97386: inst = 32'h38632800;
      97387: inst = 32'h38842800;
      97388: inst = 32'h10a00001;
      97389: inst = 32'hca07c71;
      97390: inst = 32'h13e00001;
      97391: inst = 32'hfe0d96a;
      97392: inst = 32'h5be00000;
      97393: inst = 32'h8c50000;
      97394: inst = 32'h24612800;
      97395: inst = 32'h10a00000;
      97396: inst = 32'hca0000e;
      97397: inst = 32'h24822800;
      97398: inst = 32'h10a00000;
      97399: inst = 32'hca00004;
      97400: inst = 32'h38632800;
      97401: inst = 32'h38842800;
      97402: inst = 32'h10a00001;
      97403: inst = 32'hca07c7f;
      97404: inst = 32'h13e00001;
      97405: inst = 32'hfe0d96a;
      97406: inst = 32'h5be00000;
      97407: inst = 32'h8c50000;
      97408: inst = 32'h24612800;
      97409: inst = 32'h10a00000;
      97410: inst = 32'hca0000e;
      97411: inst = 32'h24822800;
      97412: inst = 32'h10a00000;
      97413: inst = 32'hca00004;
      97414: inst = 32'h38632800;
      97415: inst = 32'h38842800;
      97416: inst = 32'h10a00001;
      97417: inst = 32'hca07c8d;
      97418: inst = 32'h13e00001;
      97419: inst = 32'hfe0d96a;
      97420: inst = 32'h5be00000;
      97421: inst = 32'h8c50000;
      97422: inst = 32'h24612800;
      97423: inst = 32'h10a00000;
      97424: inst = 32'hca0000e;
      97425: inst = 32'h24822800;
      97426: inst = 32'h10a00000;
      97427: inst = 32'hca00004;
      97428: inst = 32'h38632800;
      97429: inst = 32'h38842800;
      97430: inst = 32'h10a00001;
      97431: inst = 32'hca07c9b;
      97432: inst = 32'h13e00001;
      97433: inst = 32'hfe0d96a;
      97434: inst = 32'h5be00000;
      97435: inst = 32'h8c50000;
      97436: inst = 32'h24612800;
      97437: inst = 32'h10a00000;
      97438: inst = 32'hca0000e;
      97439: inst = 32'h24822800;
      97440: inst = 32'h10a00000;
      97441: inst = 32'hca00004;
      97442: inst = 32'h38632800;
      97443: inst = 32'h38842800;
      97444: inst = 32'h10a00001;
      97445: inst = 32'hca07ca9;
      97446: inst = 32'h13e00001;
      97447: inst = 32'hfe0d96a;
      97448: inst = 32'h5be00000;
      97449: inst = 32'h8c50000;
      97450: inst = 32'h24612800;
      97451: inst = 32'h10a00000;
      97452: inst = 32'hca0000e;
      97453: inst = 32'h24822800;
      97454: inst = 32'h10a00000;
      97455: inst = 32'hca00004;
      97456: inst = 32'h38632800;
      97457: inst = 32'h38842800;
      97458: inst = 32'h10a00001;
      97459: inst = 32'hca07cb7;
      97460: inst = 32'h13e00001;
      97461: inst = 32'hfe0d96a;
      97462: inst = 32'h5be00000;
      97463: inst = 32'h8c50000;
      97464: inst = 32'h24612800;
      97465: inst = 32'h10a00000;
      97466: inst = 32'hca0000e;
      97467: inst = 32'h24822800;
      97468: inst = 32'h10a00000;
      97469: inst = 32'hca00004;
      97470: inst = 32'h38632800;
      97471: inst = 32'h38842800;
      97472: inst = 32'h10a00001;
      97473: inst = 32'hca07cc5;
      97474: inst = 32'h13e00001;
      97475: inst = 32'hfe0d96a;
      97476: inst = 32'h5be00000;
      97477: inst = 32'h8c50000;
      97478: inst = 32'h24612800;
      97479: inst = 32'h10a00000;
      97480: inst = 32'hca0000e;
      97481: inst = 32'h24822800;
      97482: inst = 32'h10a00000;
      97483: inst = 32'hca00004;
      97484: inst = 32'h38632800;
      97485: inst = 32'h38842800;
      97486: inst = 32'h10a00001;
      97487: inst = 32'hca07cd3;
      97488: inst = 32'h13e00001;
      97489: inst = 32'hfe0d96a;
      97490: inst = 32'h5be00000;
      97491: inst = 32'h8c50000;
      97492: inst = 32'h24612800;
      97493: inst = 32'h10a00000;
      97494: inst = 32'hca0000e;
      97495: inst = 32'h24822800;
      97496: inst = 32'h10a00000;
      97497: inst = 32'hca00004;
      97498: inst = 32'h38632800;
      97499: inst = 32'h38842800;
      97500: inst = 32'h10a00001;
      97501: inst = 32'hca07ce1;
      97502: inst = 32'h13e00001;
      97503: inst = 32'hfe0d96a;
      97504: inst = 32'h5be00000;
      97505: inst = 32'h8c50000;
      97506: inst = 32'h24612800;
      97507: inst = 32'h10a00000;
      97508: inst = 32'hca0000e;
      97509: inst = 32'h24822800;
      97510: inst = 32'h10a00000;
      97511: inst = 32'hca00004;
      97512: inst = 32'h38632800;
      97513: inst = 32'h38842800;
      97514: inst = 32'h10a00001;
      97515: inst = 32'hca07cef;
      97516: inst = 32'h13e00001;
      97517: inst = 32'hfe0d96a;
      97518: inst = 32'h5be00000;
      97519: inst = 32'h8c50000;
      97520: inst = 32'h24612800;
      97521: inst = 32'h10a00000;
      97522: inst = 32'hca0000e;
      97523: inst = 32'h24822800;
      97524: inst = 32'h10a00000;
      97525: inst = 32'hca00004;
      97526: inst = 32'h38632800;
      97527: inst = 32'h38842800;
      97528: inst = 32'h10a00001;
      97529: inst = 32'hca07cfd;
      97530: inst = 32'h13e00001;
      97531: inst = 32'hfe0d96a;
      97532: inst = 32'h5be00000;
      97533: inst = 32'h8c50000;
      97534: inst = 32'h24612800;
      97535: inst = 32'h10a00000;
      97536: inst = 32'hca0000e;
      97537: inst = 32'h24822800;
      97538: inst = 32'h10a00000;
      97539: inst = 32'hca00004;
      97540: inst = 32'h38632800;
      97541: inst = 32'h38842800;
      97542: inst = 32'h10a00001;
      97543: inst = 32'hca07d0b;
      97544: inst = 32'h13e00001;
      97545: inst = 32'hfe0d96a;
      97546: inst = 32'h5be00000;
      97547: inst = 32'h8c50000;
      97548: inst = 32'h24612800;
      97549: inst = 32'h10a00000;
      97550: inst = 32'hca0000e;
      97551: inst = 32'h24822800;
      97552: inst = 32'h10a00000;
      97553: inst = 32'hca00004;
      97554: inst = 32'h38632800;
      97555: inst = 32'h38842800;
      97556: inst = 32'h10a00001;
      97557: inst = 32'hca07d19;
      97558: inst = 32'h13e00001;
      97559: inst = 32'hfe0d96a;
      97560: inst = 32'h5be00000;
      97561: inst = 32'h8c50000;
      97562: inst = 32'h24612800;
      97563: inst = 32'h10a00000;
      97564: inst = 32'hca0000e;
      97565: inst = 32'h24822800;
      97566: inst = 32'h10a00000;
      97567: inst = 32'hca00004;
      97568: inst = 32'h38632800;
      97569: inst = 32'h38842800;
      97570: inst = 32'h10a00001;
      97571: inst = 32'hca07d27;
      97572: inst = 32'h13e00001;
      97573: inst = 32'hfe0d96a;
      97574: inst = 32'h5be00000;
      97575: inst = 32'h8c50000;
      97576: inst = 32'h24612800;
      97577: inst = 32'h10a00000;
      97578: inst = 32'hca0000e;
      97579: inst = 32'h24822800;
      97580: inst = 32'h10a00000;
      97581: inst = 32'hca00004;
      97582: inst = 32'h38632800;
      97583: inst = 32'h38842800;
      97584: inst = 32'h10a00001;
      97585: inst = 32'hca07d35;
      97586: inst = 32'h13e00001;
      97587: inst = 32'hfe0d96a;
      97588: inst = 32'h5be00000;
      97589: inst = 32'h8c50000;
      97590: inst = 32'h24612800;
      97591: inst = 32'h10a00000;
      97592: inst = 32'hca0000e;
      97593: inst = 32'h24822800;
      97594: inst = 32'h10a00000;
      97595: inst = 32'hca00004;
      97596: inst = 32'h38632800;
      97597: inst = 32'h38842800;
      97598: inst = 32'h10a00001;
      97599: inst = 32'hca07d43;
      97600: inst = 32'h13e00001;
      97601: inst = 32'hfe0d96a;
      97602: inst = 32'h5be00000;
      97603: inst = 32'h8c50000;
      97604: inst = 32'h24612800;
      97605: inst = 32'h10a00000;
      97606: inst = 32'hca0000e;
      97607: inst = 32'h24822800;
      97608: inst = 32'h10a00000;
      97609: inst = 32'hca00004;
      97610: inst = 32'h38632800;
      97611: inst = 32'h38842800;
      97612: inst = 32'h10a00001;
      97613: inst = 32'hca07d51;
      97614: inst = 32'h13e00001;
      97615: inst = 32'hfe0d96a;
      97616: inst = 32'h5be00000;
      97617: inst = 32'h8c50000;
      97618: inst = 32'h24612800;
      97619: inst = 32'h10a00000;
      97620: inst = 32'hca0000e;
      97621: inst = 32'h24822800;
      97622: inst = 32'h10a00000;
      97623: inst = 32'hca00004;
      97624: inst = 32'h38632800;
      97625: inst = 32'h38842800;
      97626: inst = 32'h10a00001;
      97627: inst = 32'hca07d5f;
      97628: inst = 32'h13e00001;
      97629: inst = 32'hfe0d96a;
      97630: inst = 32'h5be00000;
      97631: inst = 32'h8c50000;
      97632: inst = 32'h24612800;
      97633: inst = 32'h10a00000;
      97634: inst = 32'hca0000e;
      97635: inst = 32'h24822800;
      97636: inst = 32'h10a00000;
      97637: inst = 32'hca00004;
      97638: inst = 32'h38632800;
      97639: inst = 32'h38842800;
      97640: inst = 32'h10a00001;
      97641: inst = 32'hca07d6d;
      97642: inst = 32'h13e00001;
      97643: inst = 32'hfe0d96a;
      97644: inst = 32'h5be00000;
      97645: inst = 32'h8c50000;
      97646: inst = 32'h24612800;
      97647: inst = 32'h10a00000;
      97648: inst = 32'hca0000e;
      97649: inst = 32'h24822800;
      97650: inst = 32'h10a00000;
      97651: inst = 32'hca00004;
      97652: inst = 32'h38632800;
      97653: inst = 32'h38842800;
      97654: inst = 32'h10a00001;
      97655: inst = 32'hca07d7b;
      97656: inst = 32'h13e00001;
      97657: inst = 32'hfe0d96a;
      97658: inst = 32'h5be00000;
      97659: inst = 32'h8c50000;
      97660: inst = 32'h24612800;
      97661: inst = 32'h10a00000;
      97662: inst = 32'hca0000e;
      97663: inst = 32'h24822800;
      97664: inst = 32'h10a00000;
      97665: inst = 32'hca00004;
      97666: inst = 32'h38632800;
      97667: inst = 32'h38842800;
      97668: inst = 32'h10a00001;
      97669: inst = 32'hca07d89;
      97670: inst = 32'h13e00001;
      97671: inst = 32'hfe0d96a;
      97672: inst = 32'h5be00000;
      97673: inst = 32'h8c50000;
      97674: inst = 32'h24612800;
      97675: inst = 32'h10a00000;
      97676: inst = 32'hca0000e;
      97677: inst = 32'h24822800;
      97678: inst = 32'h10a00000;
      97679: inst = 32'hca00004;
      97680: inst = 32'h38632800;
      97681: inst = 32'h38842800;
      97682: inst = 32'h10a00001;
      97683: inst = 32'hca07d97;
      97684: inst = 32'h13e00001;
      97685: inst = 32'hfe0d96a;
      97686: inst = 32'h5be00000;
      97687: inst = 32'h8c50000;
      97688: inst = 32'h24612800;
      97689: inst = 32'h10a00000;
      97690: inst = 32'hca0000e;
      97691: inst = 32'h24822800;
      97692: inst = 32'h10a00000;
      97693: inst = 32'hca00004;
      97694: inst = 32'h38632800;
      97695: inst = 32'h38842800;
      97696: inst = 32'h10a00001;
      97697: inst = 32'hca07da5;
      97698: inst = 32'h13e00001;
      97699: inst = 32'hfe0d96a;
      97700: inst = 32'h5be00000;
      97701: inst = 32'h8c50000;
      97702: inst = 32'h24612800;
      97703: inst = 32'h10a00000;
      97704: inst = 32'hca0000e;
      97705: inst = 32'h24822800;
      97706: inst = 32'h10a00000;
      97707: inst = 32'hca00004;
      97708: inst = 32'h38632800;
      97709: inst = 32'h38842800;
      97710: inst = 32'h10a00001;
      97711: inst = 32'hca07db3;
      97712: inst = 32'h13e00001;
      97713: inst = 32'hfe0d96a;
      97714: inst = 32'h5be00000;
      97715: inst = 32'h8c50000;
      97716: inst = 32'h24612800;
      97717: inst = 32'h10a00000;
      97718: inst = 32'hca0000e;
      97719: inst = 32'h24822800;
      97720: inst = 32'h10a00000;
      97721: inst = 32'hca00004;
      97722: inst = 32'h38632800;
      97723: inst = 32'h38842800;
      97724: inst = 32'h10a00001;
      97725: inst = 32'hca07dc1;
      97726: inst = 32'h13e00001;
      97727: inst = 32'hfe0d96a;
      97728: inst = 32'h5be00000;
      97729: inst = 32'h8c50000;
      97730: inst = 32'h24612800;
      97731: inst = 32'h10a00000;
      97732: inst = 32'hca0000e;
      97733: inst = 32'h24822800;
      97734: inst = 32'h10a00000;
      97735: inst = 32'hca00004;
      97736: inst = 32'h38632800;
      97737: inst = 32'h38842800;
      97738: inst = 32'h10a00001;
      97739: inst = 32'hca07dcf;
      97740: inst = 32'h13e00001;
      97741: inst = 32'hfe0d96a;
      97742: inst = 32'h5be00000;
      97743: inst = 32'h8c50000;
      97744: inst = 32'h24612800;
      97745: inst = 32'h10a00000;
      97746: inst = 32'hca0000e;
      97747: inst = 32'h24822800;
      97748: inst = 32'h10a00000;
      97749: inst = 32'hca00004;
      97750: inst = 32'h38632800;
      97751: inst = 32'h38842800;
      97752: inst = 32'h10a00001;
      97753: inst = 32'hca07ddd;
      97754: inst = 32'h13e00001;
      97755: inst = 32'hfe0d96a;
      97756: inst = 32'h5be00000;
      97757: inst = 32'h8c50000;
      97758: inst = 32'h24612800;
      97759: inst = 32'h10a00000;
      97760: inst = 32'hca0000e;
      97761: inst = 32'h24822800;
      97762: inst = 32'h10a00000;
      97763: inst = 32'hca00004;
      97764: inst = 32'h38632800;
      97765: inst = 32'h38842800;
      97766: inst = 32'h10a00001;
      97767: inst = 32'hca07deb;
      97768: inst = 32'h13e00001;
      97769: inst = 32'hfe0d96a;
      97770: inst = 32'h5be00000;
      97771: inst = 32'h8c50000;
      97772: inst = 32'h24612800;
      97773: inst = 32'h10a00000;
      97774: inst = 32'hca0000e;
      97775: inst = 32'h24822800;
      97776: inst = 32'h10a00000;
      97777: inst = 32'hca00004;
      97778: inst = 32'h38632800;
      97779: inst = 32'h38842800;
      97780: inst = 32'h10a00001;
      97781: inst = 32'hca07df9;
      97782: inst = 32'h13e00001;
      97783: inst = 32'hfe0d96a;
      97784: inst = 32'h5be00000;
      97785: inst = 32'h8c50000;
      97786: inst = 32'h24612800;
      97787: inst = 32'h10a00000;
      97788: inst = 32'hca0000e;
      97789: inst = 32'h24822800;
      97790: inst = 32'h10a00000;
      97791: inst = 32'hca00004;
      97792: inst = 32'h38632800;
      97793: inst = 32'h38842800;
      97794: inst = 32'h10a00001;
      97795: inst = 32'hca07e07;
      97796: inst = 32'h13e00001;
      97797: inst = 32'hfe0d96a;
      97798: inst = 32'h5be00000;
      97799: inst = 32'h8c50000;
      97800: inst = 32'h24612800;
      97801: inst = 32'h10a00000;
      97802: inst = 32'hca0000e;
      97803: inst = 32'h24822800;
      97804: inst = 32'h10a00000;
      97805: inst = 32'hca00004;
      97806: inst = 32'h38632800;
      97807: inst = 32'h38842800;
      97808: inst = 32'h10a00001;
      97809: inst = 32'hca07e15;
      97810: inst = 32'h13e00001;
      97811: inst = 32'hfe0d96a;
      97812: inst = 32'h5be00000;
      97813: inst = 32'h8c50000;
      97814: inst = 32'h24612800;
      97815: inst = 32'h10a00000;
      97816: inst = 32'hca0000e;
      97817: inst = 32'h24822800;
      97818: inst = 32'h10a00000;
      97819: inst = 32'hca00004;
      97820: inst = 32'h38632800;
      97821: inst = 32'h38842800;
      97822: inst = 32'h10a00001;
      97823: inst = 32'hca07e23;
      97824: inst = 32'h13e00001;
      97825: inst = 32'hfe0d96a;
      97826: inst = 32'h5be00000;
      97827: inst = 32'h8c50000;
      97828: inst = 32'h24612800;
      97829: inst = 32'h10a00000;
      97830: inst = 32'hca0000e;
      97831: inst = 32'h24822800;
      97832: inst = 32'h10a00000;
      97833: inst = 32'hca00004;
      97834: inst = 32'h38632800;
      97835: inst = 32'h38842800;
      97836: inst = 32'h10a00001;
      97837: inst = 32'hca07e31;
      97838: inst = 32'h13e00001;
      97839: inst = 32'hfe0d96a;
      97840: inst = 32'h5be00000;
      97841: inst = 32'h8c50000;
      97842: inst = 32'h24612800;
      97843: inst = 32'h10a00000;
      97844: inst = 32'hca0000e;
      97845: inst = 32'h24822800;
      97846: inst = 32'h10a00000;
      97847: inst = 32'hca00004;
      97848: inst = 32'h38632800;
      97849: inst = 32'h38842800;
      97850: inst = 32'h10a00001;
      97851: inst = 32'hca07e3f;
      97852: inst = 32'h13e00001;
      97853: inst = 32'hfe0d96a;
      97854: inst = 32'h5be00000;
      97855: inst = 32'h8c50000;
      97856: inst = 32'h24612800;
      97857: inst = 32'h10a00000;
      97858: inst = 32'hca0000e;
      97859: inst = 32'h24822800;
      97860: inst = 32'h10a00000;
      97861: inst = 32'hca00004;
      97862: inst = 32'h38632800;
      97863: inst = 32'h38842800;
      97864: inst = 32'h10a00001;
      97865: inst = 32'hca07e4d;
      97866: inst = 32'h13e00001;
      97867: inst = 32'hfe0d96a;
      97868: inst = 32'h5be00000;
      97869: inst = 32'h8c50000;
      97870: inst = 32'h24612800;
      97871: inst = 32'h10a00000;
      97872: inst = 32'hca0000e;
      97873: inst = 32'h24822800;
      97874: inst = 32'h10a00000;
      97875: inst = 32'hca00004;
      97876: inst = 32'h38632800;
      97877: inst = 32'h38842800;
      97878: inst = 32'h10a00001;
      97879: inst = 32'hca07e5b;
      97880: inst = 32'h13e00001;
      97881: inst = 32'hfe0d96a;
      97882: inst = 32'h5be00000;
      97883: inst = 32'h8c50000;
      97884: inst = 32'h24612800;
      97885: inst = 32'h10a00000;
      97886: inst = 32'hca0000e;
      97887: inst = 32'h24822800;
      97888: inst = 32'h10a00000;
      97889: inst = 32'hca00004;
      97890: inst = 32'h38632800;
      97891: inst = 32'h38842800;
      97892: inst = 32'h10a00001;
      97893: inst = 32'hca07e69;
      97894: inst = 32'h13e00001;
      97895: inst = 32'hfe0d96a;
      97896: inst = 32'h5be00000;
      97897: inst = 32'h8c50000;
      97898: inst = 32'h24612800;
      97899: inst = 32'h10a00000;
      97900: inst = 32'hca0000e;
      97901: inst = 32'h24822800;
      97902: inst = 32'h10a00000;
      97903: inst = 32'hca00004;
      97904: inst = 32'h38632800;
      97905: inst = 32'h38842800;
      97906: inst = 32'h10a00001;
      97907: inst = 32'hca07e77;
      97908: inst = 32'h13e00001;
      97909: inst = 32'hfe0d96a;
      97910: inst = 32'h5be00000;
      97911: inst = 32'h8c50000;
      97912: inst = 32'h24612800;
      97913: inst = 32'h10a00000;
      97914: inst = 32'hca0000e;
      97915: inst = 32'h24822800;
      97916: inst = 32'h10a00000;
      97917: inst = 32'hca00004;
      97918: inst = 32'h38632800;
      97919: inst = 32'h38842800;
      97920: inst = 32'h10a00001;
      97921: inst = 32'hca07e85;
      97922: inst = 32'h13e00001;
      97923: inst = 32'hfe0d96a;
      97924: inst = 32'h5be00000;
      97925: inst = 32'h8c50000;
      97926: inst = 32'h24612800;
      97927: inst = 32'h10a00000;
      97928: inst = 32'hca0000e;
      97929: inst = 32'h24822800;
      97930: inst = 32'h10a00000;
      97931: inst = 32'hca00004;
      97932: inst = 32'h38632800;
      97933: inst = 32'h38842800;
      97934: inst = 32'h10a00001;
      97935: inst = 32'hca07e93;
      97936: inst = 32'h13e00001;
      97937: inst = 32'hfe0d96a;
      97938: inst = 32'h5be00000;
      97939: inst = 32'h8c50000;
      97940: inst = 32'h24612800;
      97941: inst = 32'h10a00000;
      97942: inst = 32'hca0000e;
      97943: inst = 32'h24822800;
      97944: inst = 32'h10a00000;
      97945: inst = 32'hca00004;
      97946: inst = 32'h38632800;
      97947: inst = 32'h38842800;
      97948: inst = 32'h10a00001;
      97949: inst = 32'hca07ea1;
      97950: inst = 32'h13e00001;
      97951: inst = 32'hfe0d96a;
      97952: inst = 32'h5be00000;
      97953: inst = 32'h8c50000;
      97954: inst = 32'h24612800;
      97955: inst = 32'h10a00000;
      97956: inst = 32'hca0000e;
      97957: inst = 32'h24822800;
      97958: inst = 32'h10a00000;
      97959: inst = 32'hca00004;
      97960: inst = 32'h38632800;
      97961: inst = 32'h38842800;
      97962: inst = 32'h10a00001;
      97963: inst = 32'hca07eaf;
      97964: inst = 32'h13e00001;
      97965: inst = 32'hfe0d96a;
      97966: inst = 32'h5be00000;
      97967: inst = 32'h8c50000;
      97968: inst = 32'h24612800;
      97969: inst = 32'h10a00000;
      97970: inst = 32'hca0000e;
      97971: inst = 32'h24822800;
      97972: inst = 32'h10a00000;
      97973: inst = 32'hca00004;
      97974: inst = 32'h38632800;
      97975: inst = 32'h38842800;
      97976: inst = 32'h10a00001;
      97977: inst = 32'hca07ebd;
      97978: inst = 32'h13e00001;
      97979: inst = 32'hfe0d96a;
      97980: inst = 32'h5be00000;
      97981: inst = 32'h8c50000;
      97982: inst = 32'h24612800;
      97983: inst = 32'h10a00000;
      97984: inst = 32'hca0000e;
      97985: inst = 32'h24822800;
      97986: inst = 32'h10a00000;
      97987: inst = 32'hca00004;
      97988: inst = 32'h38632800;
      97989: inst = 32'h38842800;
      97990: inst = 32'h10a00001;
      97991: inst = 32'hca07ecb;
      97992: inst = 32'h13e00001;
      97993: inst = 32'hfe0d96a;
      97994: inst = 32'h5be00000;
      97995: inst = 32'h8c50000;
      97996: inst = 32'h24612800;
      97997: inst = 32'h10a00000;
      97998: inst = 32'hca0000e;
      97999: inst = 32'h24822800;
      98000: inst = 32'h10a00000;
      98001: inst = 32'hca00004;
      98002: inst = 32'h38632800;
      98003: inst = 32'h38842800;
      98004: inst = 32'h10a00001;
      98005: inst = 32'hca07ed9;
      98006: inst = 32'h13e00001;
      98007: inst = 32'hfe0d96a;
      98008: inst = 32'h5be00000;
      98009: inst = 32'h8c50000;
      98010: inst = 32'h24612800;
      98011: inst = 32'h10a00000;
      98012: inst = 32'hca0000e;
      98013: inst = 32'h24822800;
      98014: inst = 32'h10a00000;
      98015: inst = 32'hca00004;
      98016: inst = 32'h38632800;
      98017: inst = 32'h38842800;
      98018: inst = 32'h10a00001;
      98019: inst = 32'hca07ee7;
      98020: inst = 32'h13e00001;
      98021: inst = 32'hfe0d96a;
      98022: inst = 32'h5be00000;
      98023: inst = 32'h8c50000;
      98024: inst = 32'h24612800;
      98025: inst = 32'h10a00000;
      98026: inst = 32'hca0000e;
      98027: inst = 32'h24822800;
      98028: inst = 32'h10a00000;
      98029: inst = 32'hca00004;
      98030: inst = 32'h38632800;
      98031: inst = 32'h38842800;
      98032: inst = 32'h10a00001;
      98033: inst = 32'hca07ef5;
      98034: inst = 32'h13e00001;
      98035: inst = 32'hfe0d96a;
      98036: inst = 32'h5be00000;
      98037: inst = 32'h8c50000;
      98038: inst = 32'h24612800;
      98039: inst = 32'h10a00000;
      98040: inst = 32'hca0000e;
      98041: inst = 32'h24822800;
      98042: inst = 32'h10a00000;
      98043: inst = 32'hca00004;
      98044: inst = 32'h38632800;
      98045: inst = 32'h38842800;
      98046: inst = 32'h10a00001;
      98047: inst = 32'hca07f03;
      98048: inst = 32'h13e00001;
      98049: inst = 32'hfe0d96a;
      98050: inst = 32'h5be00000;
      98051: inst = 32'h8c50000;
      98052: inst = 32'h24612800;
      98053: inst = 32'h10a00000;
      98054: inst = 32'hca0000e;
      98055: inst = 32'h24822800;
      98056: inst = 32'h10a00000;
      98057: inst = 32'hca00004;
      98058: inst = 32'h38632800;
      98059: inst = 32'h38842800;
      98060: inst = 32'h10a00001;
      98061: inst = 32'hca07f11;
      98062: inst = 32'h13e00001;
      98063: inst = 32'hfe0d96a;
      98064: inst = 32'h5be00000;
      98065: inst = 32'h8c50000;
      98066: inst = 32'h24612800;
      98067: inst = 32'h10a00000;
      98068: inst = 32'hca0000e;
      98069: inst = 32'h24822800;
      98070: inst = 32'h10a00000;
      98071: inst = 32'hca00004;
      98072: inst = 32'h38632800;
      98073: inst = 32'h38842800;
      98074: inst = 32'h10a00001;
      98075: inst = 32'hca07f1f;
      98076: inst = 32'h13e00001;
      98077: inst = 32'hfe0d96a;
      98078: inst = 32'h5be00000;
      98079: inst = 32'h8c50000;
      98080: inst = 32'h24612800;
      98081: inst = 32'h10a00000;
      98082: inst = 32'hca0000e;
      98083: inst = 32'h24822800;
      98084: inst = 32'h10a00000;
      98085: inst = 32'hca00004;
      98086: inst = 32'h38632800;
      98087: inst = 32'h38842800;
      98088: inst = 32'h10a00001;
      98089: inst = 32'hca07f2d;
      98090: inst = 32'h13e00001;
      98091: inst = 32'hfe0d96a;
      98092: inst = 32'h5be00000;
      98093: inst = 32'h8c50000;
      98094: inst = 32'h24612800;
      98095: inst = 32'h10a00000;
      98096: inst = 32'hca0000e;
      98097: inst = 32'h24822800;
      98098: inst = 32'h10a00000;
      98099: inst = 32'hca00004;
      98100: inst = 32'h38632800;
      98101: inst = 32'h38842800;
      98102: inst = 32'h10a00001;
      98103: inst = 32'hca07f3b;
      98104: inst = 32'h13e00001;
      98105: inst = 32'hfe0d96a;
      98106: inst = 32'h5be00000;
      98107: inst = 32'h8c50000;
      98108: inst = 32'h24612800;
      98109: inst = 32'h10a00000;
      98110: inst = 32'hca0000e;
      98111: inst = 32'h24822800;
      98112: inst = 32'h10a00000;
      98113: inst = 32'hca00004;
      98114: inst = 32'h38632800;
      98115: inst = 32'h38842800;
      98116: inst = 32'h10a00001;
      98117: inst = 32'hca07f49;
      98118: inst = 32'h13e00001;
      98119: inst = 32'hfe0d96a;
      98120: inst = 32'h5be00000;
      98121: inst = 32'h8c50000;
      98122: inst = 32'h24612800;
      98123: inst = 32'h10a00000;
      98124: inst = 32'hca0000e;
      98125: inst = 32'h24822800;
      98126: inst = 32'h10a00000;
      98127: inst = 32'hca00004;
      98128: inst = 32'h38632800;
      98129: inst = 32'h38842800;
      98130: inst = 32'h10a00001;
      98131: inst = 32'hca07f57;
      98132: inst = 32'h13e00001;
      98133: inst = 32'hfe0d96a;
      98134: inst = 32'h5be00000;
      98135: inst = 32'h8c50000;
      98136: inst = 32'h24612800;
      98137: inst = 32'h10a00000;
      98138: inst = 32'hca0000e;
      98139: inst = 32'h24822800;
      98140: inst = 32'h10a00000;
      98141: inst = 32'hca00004;
      98142: inst = 32'h38632800;
      98143: inst = 32'h38842800;
      98144: inst = 32'h10a00001;
      98145: inst = 32'hca07f65;
      98146: inst = 32'h13e00001;
      98147: inst = 32'hfe0d96a;
      98148: inst = 32'h5be00000;
      98149: inst = 32'h8c50000;
      98150: inst = 32'h24612800;
      98151: inst = 32'h10a00000;
      98152: inst = 32'hca0000e;
      98153: inst = 32'h24822800;
      98154: inst = 32'h10a00000;
      98155: inst = 32'hca00004;
      98156: inst = 32'h38632800;
      98157: inst = 32'h38842800;
      98158: inst = 32'h10a00001;
      98159: inst = 32'hca07f73;
      98160: inst = 32'h13e00001;
      98161: inst = 32'hfe0d96a;
      98162: inst = 32'h5be00000;
      98163: inst = 32'h8c50000;
      98164: inst = 32'h24612800;
      98165: inst = 32'h10a00000;
      98166: inst = 32'hca0000e;
      98167: inst = 32'h24822800;
      98168: inst = 32'h10a00000;
      98169: inst = 32'hca00004;
      98170: inst = 32'h38632800;
      98171: inst = 32'h38842800;
      98172: inst = 32'h10a00001;
      98173: inst = 32'hca07f81;
      98174: inst = 32'h13e00001;
      98175: inst = 32'hfe0d96a;
      98176: inst = 32'h5be00000;
      98177: inst = 32'h8c50000;
      98178: inst = 32'h24612800;
      98179: inst = 32'h10a00000;
      98180: inst = 32'hca0000e;
      98181: inst = 32'h24822800;
      98182: inst = 32'h10a00000;
      98183: inst = 32'hca00004;
      98184: inst = 32'h38632800;
      98185: inst = 32'h38842800;
      98186: inst = 32'h10a00001;
      98187: inst = 32'hca07f8f;
      98188: inst = 32'h13e00001;
      98189: inst = 32'hfe0d96a;
      98190: inst = 32'h5be00000;
      98191: inst = 32'h8c50000;
      98192: inst = 32'h24612800;
      98193: inst = 32'h10a00000;
      98194: inst = 32'hca0000e;
      98195: inst = 32'h24822800;
      98196: inst = 32'h10a00000;
      98197: inst = 32'hca00004;
      98198: inst = 32'h38632800;
      98199: inst = 32'h38842800;
      98200: inst = 32'h10a00001;
      98201: inst = 32'hca07f9d;
      98202: inst = 32'h13e00001;
      98203: inst = 32'hfe0d96a;
      98204: inst = 32'h5be00000;
      98205: inst = 32'h8c50000;
      98206: inst = 32'h24612800;
      98207: inst = 32'h10a00000;
      98208: inst = 32'hca0000e;
      98209: inst = 32'h24822800;
      98210: inst = 32'h10a00000;
      98211: inst = 32'hca00004;
      98212: inst = 32'h38632800;
      98213: inst = 32'h38842800;
      98214: inst = 32'h10a00001;
      98215: inst = 32'hca07fab;
      98216: inst = 32'h13e00001;
      98217: inst = 32'hfe0d96a;
      98218: inst = 32'h5be00000;
      98219: inst = 32'h8c50000;
      98220: inst = 32'h24612800;
      98221: inst = 32'h10a00000;
      98222: inst = 32'hca0000e;
      98223: inst = 32'h24822800;
      98224: inst = 32'h10a00000;
      98225: inst = 32'hca00004;
      98226: inst = 32'h38632800;
      98227: inst = 32'h38842800;
      98228: inst = 32'h10a00001;
      98229: inst = 32'hca07fb9;
      98230: inst = 32'h13e00001;
      98231: inst = 32'hfe0d96a;
      98232: inst = 32'h5be00000;
      98233: inst = 32'h8c50000;
      98234: inst = 32'h24612800;
      98235: inst = 32'h10a00000;
      98236: inst = 32'hca0000e;
      98237: inst = 32'h24822800;
      98238: inst = 32'h10a00000;
      98239: inst = 32'hca00004;
      98240: inst = 32'h38632800;
      98241: inst = 32'h38842800;
      98242: inst = 32'h10a00001;
      98243: inst = 32'hca07fc7;
      98244: inst = 32'h13e00001;
      98245: inst = 32'hfe0d96a;
      98246: inst = 32'h5be00000;
      98247: inst = 32'h8c50000;
      98248: inst = 32'h24612800;
      98249: inst = 32'h10a00000;
      98250: inst = 32'hca0000e;
      98251: inst = 32'h24822800;
      98252: inst = 32'h10a00000;
      98253: inst = 32'hca00004;
      98254: inst = 32'h38632800;
      98255: inst = 32'h38842800;
      98256: inst = 32'h10a00001;
      98257: inst = 32'hca07fd5;
      98258: inst = 32'h13e00001;
      98259: inst = 32'hfe0d96a;
      98260: inst = 32'h5be00000;
      98261: inst = 32'h8c50000;
      98262: inst = 32'h24612800;
      98263: inst = 32'h10a00000;
      98264: inst = 32'hca0000e;
      98265: inst = 32'h24822800;
      98266: inst = 32'h10a00000;
      98267: inst = 32'hca00004;
      98268: inst = 32'h38632800;
      98269: inst = 32'h38842800;
      98270: inst = 32'h10a00001;
      98271: inst = 32'hca07fe3;
      98272: inst = 32'h13e00001;
      98273: inst = 32'hfe0d96a;
      98274: inst = 32'h5be00000;
      98275: inst = 32'h8c50000;
      98276: inst = 32'h24612800;
      98277: inst = 32'h10a00000;
      98278: inst = 32'hca0000e;
      98279: inst = 32'h24822800;
      98280: inst = 32'h10a00000;
      98281: inst = 32'hca00004;
      98282: inst = 32'h38632800;
      98283: inst = 32'h38842800;
      98284: inst = 32'h10a00001;
      98285: inst = 32'hca07ff1;
      98286: inst = 32'h13e00001;
      98287: inst = 32'hfe0d96a;
      98288: inst = 32'h5be00000;
      98289: inst = 32'h8c50000;
      98290: inst = 32'h24612800;
      98291: inst = 32'h10a00000;
      98292: inst = 32'hca0000e;
      98293: inst = 32'h24822800;
      98294: inst = 32'h10a00000;
      98295: inst = 32'hca00004;
      98296: inst = 32'h38632800;
      98297: inst = 32'h38842800;
      98298: inst = 32'h10a00001;
      98299: inst = 32'hca07fff;
      98300: inst = 32'h13e00001;
      98301: inst = 32'hfe0d96a;
      98302: inst = 32'h5be00000;
      98303: inst = 32'h8c50000;
      98304: inst = 32'h24612800;
      98305: inst = 32'h10a00000;
      98306: inst = 32'hca0000e;
      98307: inst = 32'h24822800;
      98308: inst = 32'h10a00000;
      98309: inst = 32'hca00004;
      98310: inst = 32'h38632800;
      98311: inst = 32'h38842800;
      98312: inst = 32'h10a00001;
      98313: inst = 32'hca0800d;
      98314: inst = 32'h13e00001;
      98315: inst = 32'hfe0d96a;
      98316: inst = 32'h5be00000;
      98317: inst = 32'h8c50000;
      98318: inst = 32'h24612800;
      98319: inst = 32'h10a00000;
      98320: inst = 32'hca0000e;
      98321: inst = 32'h24822800;
      98322: inst = 32'h10a00000;
      98323: inst = 32'hca00004;
      98324: inst = 32'h38632800;
      98325: inst = 32'h38842800;
      98326: inst = 32'h10a00001;
      98327: inst = 32'hca0801b;
      98328: inst = 32'h13e00001;
      98329: inst = 32'hfe0d96a;
      98330: inst = 32'h5be00000;
      98331: inst = 32'h8c50000;
      98332: inst = 32'h24612800;
      98333: inst = 32'h10a00000;
      98334: inst = 32'hca0000e;
      98335: inst = 32'h24822800;
      98336: inst = 32'h10a00000;
      98337: inst = 32'hca00004;
      98338: inst = 32'h38632800;
      98339: inst = 32'h38842800;
      98340: inst = 32'h10a00001;
      98341: inst = 32'hca08029;
      98342: inst = 32'h13e00001;
      98343: inst = 32'hfe0d96a;
      98344: inst = 32'h5be00000;
      98345: inst = 32'h8c50000;
      98346: inst = 32'h24612800;
      98347: inst = 32'h10a00000;
      98348: inst = 32'hca0000f;
      98349: inst = 32'h24822800;
      98350: inst = 32'h10a00000;
      98351: inst = 32'hca00004;
      98352: inst = 32'h38632800;
      98353: inst = 32'h38842800;
      98354: inst = 32'h10a00001;
      98355: inst = 32'hca08037;
      98356: inst = 32'h13e00001;
      98357: inst = 32'hfe0d96a;
      98358: inst = 32'h5be00000;
      98359: inst = 32'h8c50000;
      98360: inst = 32'h24612800;
      98361: inst = 32'h10a00000;
      98362: inst = 32'hca0000f;
      98363: inst = 32'h24822800;
      98364: inst = 32'h10a00000;
      98365: inst = 32'hca00004;
      98366: inst = 32'h38632800;
      98367: inst = 32'h38842800;
      98368: inst = 32'h10a00001;
      98369: inst = 32'hca08045;
      98370: inst = 32'h13e00001;
      98371: inst = 32'hfe0d96a;
      98372: inst = 32'h5be00000;
      98373: inst = 32'h8c50000;
      98374: inst = 32'h24612800;
      98375: inst = 32'h10a00000;
      98376: inst = 32'hca0000f;
      98377: inst = 32'h24822800;
      98378: inst = 32'h10a00000;
      98379: inst = 32'hca00004;
      98380: inst = 32'h38632800;
      98381: inst = 32'h38842800;
      98382: inst = 32'h10a00001;
      98383: inst = 32'hca08053;
      98384: inst = 32'h13e00001;
      98385: inst = 32'hfe0d96a;
      98386: inst = 32'h5be00000;
      98387: inst = 32'h8c50000;
      98388: inst = 32'h24612800;
      98389: inst = 32'h10a00000;
      98390: inst = 32'hca0000f;
      98391: inst = 32'h24822800;
      98392: inst = 32'h10a00000;
      98393: inst = 32'hca00004;
      98394: inst = 32'h38632800;
      98395: inst = 32'h38842800;
      98396: inst = 32'h10a00001;
      98397: inst = 32'hca08061;
      98398: inst = 32'h13e00001;
      98399: inst = 32'hfe0d96a;
      98400: inst = 32'h5be00000;
      98401: inst = 32'h8c50000;
      98402: inst = 32'h24612800;
      98403: inst = 32'h10a00000;
      98404: inst = 32'hca0000f;
      98405: inst = 32'h24822800;
      98406: inst = 32'h10a00000;
      98407: inst = 32'hca00004;
      98408: inst = 32'h38632800;
      98409: inst = 32'h38842800;
      98410: inst = 32'h10a00001;
      98411: inst = 32'hca0806f;
      98412: inst = 32'h13e00001;
      98413: inst = 32'hfe0d96a;
      98414: inst = 32'h5be00000;
      98415: inst = 32'h8c50000;
      98416: inst = 32'h24612800;
      98417: inst = 32'h10a00000;
      98418: inst = 32'hca0000f;
      98419: inst = 32'h24822800;
      98420: inst = 32'h10a00000;
      98421: inst = 32'hca00004;
      98422: inst = 32'h38632800;
      98423: inst = 32'h38842800;
      98424: inst = 32'h10a00001;
      98425: inst = 32'hca0807d;
      98426: inst = 32'h13e00001;
      98427: inst = 32'hfe0d96a;
      98428: inst = 32'h5be00000;
      98429: inst = 32'h8c50000;
      98430: inst = 32'h24612800;
      98431: inst = 32'h10a00000;
      98432: inst = 32'hca0000f;
      98433: inst = 32'h24822800;
      98434: inst = 32'h10a00000;
      98435: inst = 32'hca00004;
      98436: inst = 32'h38632800;
      98437: inst = 32'h38842800;
      98438: inst = 32'h10a00001;
      98439: inst = 32'hca0808b;
      98440: inst = 32'h13e00001;
      98441: inst = 32'hfe0d96a;
      98442: inst = 32'h5be00000;
      98443: inst = 32'h8c50000;
      98444: inst = 32'h24612800;
      98445: inst = 32'h10a00000;
      98446: inst = 32'hca0000f;
      98447: inst = 32'h24822800;
      98448: inst = 32'h10a00000;
      98449: inst = 32'hca00004;
      98450: inst = 32'h38632800;
      98451: inst = 32'h38842800;
      98452: inst = 32'h10a00001;
      98453: inst = 32'hca08099;
      98454: inst = 32'h13e00001;
      98455: inst = 32'hfe0d96a;
      98456: inst = 32'h5be00000;
      98457: inst = 32'h8c50000;
      98458: inst = 32'h24612800;
      98459: inst = 32'h10a00000;
      98460: inst = 32'hca0000f;
      98461: inst = 32'h24822800;
      98462: inst = 32'h10a00000;
      98463: inst = 32'hca00004;
      98464: inst = 32'h38632800;
      98465: inst = 32'h38842800;
      98466: inst = 32'h10a00001;
      98467: inst = 32'hca080a7;
      98468: inst = 32'h13e00001;
      98469: inst = 32'hfe0d96a;
      98470: inst = 32'h5be00000;
      98471: inst = 32'h8c50000;
      98472: inst = 32'h24612800;
      98473: inst = 32'h10a00000;
      98474: inst = 32'hca0000f;
      98475: inst = 32'h24822800;
      98476: inst = 32'h10a00000;
      98477: inst = 32'hca00004;
      98478: inst = 32'h38632800;
      98479: inst = 32'h38842800;
      98480: inst = 32'h10a00001;
      98481: inst = 32'hca080b5;
      98482: inst = 32'h13e00001;
      98483: inst = 32'hfe0d96a;
      98484: inst = 32'h5be00000;
      98485: inst = 32'h8c50000;
      98486: inst = 32'h24612800;
      98487: inst = 32'h10a00000;
      98488: inst = 32'hca0000f;
      98489: inst = 32'h24822800;
      98490: inst = 32'h10a00000;
      98491: inst = 32'hca00004;
      98492: inst = 32'h38632800;
      98493: inst = 32'h38842800;
      98494: inst = 32'h10a00001;
      98495: inst = 32'hca080c3;
      98496: inst = 32'h13e00001;
      98497: inst = 32'hfe0d96a;
      98498: inst = 32'h5be00000;
      98499: inst = 32'h8c50000;
      98500: inst = 32'h24612800;
      98501: inst = 32'h10a00000;
      98502: inst = 32'hca0000f;
      98503: inst = 32'h24822800;
      98504: inst = 32'h10a00000;
      98505: inst = 32'hca00004;
      98506: inst = 32'h38632800;
      98507: inst = 32'h38842800;
      98508: inst = 32'h10a00001;
      98509: inst = 32'hca080d1;
      98510: inst = 32'h13e00001;
      98511: inst = 32'hfe0d96a;
      98512: inst = 32'h5be00000;
      98513: inst = 32'h8c50000;
      98514: inst = 32'h24612800;
      98515: inst = 32'h10a00000;
      98516: inst = 32'hca0000f;
      98517: inst = 32'h24822800;
      98518: inst = 32'h10a00000;
      98519: inst = 32'hca00004;
      98520: inst = 32'h38632800;
      98521: inst = 32'h38842800;
      98522: inst = 32'h10a00001;
      98523: inst = 32'hca080df;
      98524: inst = 32'h13e00001;
      98525: inst = 32'hfe0d96a;
      98526: inst = 32'h5be00000;
      98527: inst = 32'h8c50000;
      98528: inst = 32'h24612800;
      98529: inst = 32'h10a00000;
      98530: inst = 32'hca0000f;
      98531: inst = 32'h24822800;
      98532: inst = 32'h10a00000;
      98533: inst = 32'hca00004;
      98534: inst = 32'h38632800;
      98535: inst = 32'h38842800;
      98536: inst = 32'h10a00001;
      98537: inst = 32'hca080ed;
      98538: inst = 32'h13e00001;
      98539: inst = 32'hfe0d96a;
      98540: inst = 32'h5be00000;
      98541: inst = 32'h8c50000;
      98542: inst = 32'h24612800;
      98543: inst = 32'h10a00000;
      98544: inst = 32'hca0000f;
      98545: inst = 32'h24822800;
      98546: inst = 32'h10a00000;
      98547: inst = 32'hca00004;
      98548: inst = 32'h38632800;
      98549: inst = 32'h38842800;
      98550: inst = 32'h10a00001;
      98551: inst = 32'hca080fb;
      98552: inst = 32'h13e00001;
      98553: inst = 32'hfe0d96a;
      98554: inst = 32'h5be00000;
      98555: inst = 32'h8c50000;
      98556: inst = 32'h24612800;
      98557: inst = 32'h10a00000;
      98558: inst = 32'hca0000f;
      98559: inst = 32'h24822800;
      98560: inst = 32'h10a00000;
      98561: inst = 32'hca00004;
      98562: inst = 32'h38632800;
      98563: inst = 32'h38842800;
      98564: inst = 32'h10a00001;
      98565: inst = 32'hca08109;
      98566: inst = 32'h13e00001;
      98567: inst = 32'hfe0d96a;
      98568: inst = 32'h5be00000;
      98569: inst = 32'h8c50000;
      98570: inst = 32'h24612800;
      98571: inst = 32'h10a00000;
      98572: inst = 32'hca0000f;
      98573: inst = 32'h24822800;
      98574: inst = 32'h10a00000;
      98575: inst = 32'hca00004;
      98576: inst = 32'h38632800;
      98577: inst = 32'h38842800;
      98578: inst = 32'h10a00001;
      98579: inst = 32'hca08117;
      98580: inst = 32'h13e00001;
      98581: inst = 32'hfe0d96a;
      98582: inst = 32'h5be00000;
      98583: inst = 32'h8c50000;
      98584: inst = 32'h24612800;
      98585: inst = 32'h10a00000;
      98586: inst = 32'hca0000f;
      98587: inst = 32'h24822800;
      98588: inst = 32'h10a00000;
      98589: inst = 32'hca00004;
      98590: inst = 32'h38632800;
      98591: inst = 32'h38842800;
      98592: inst = 32'h10a00001;
      98593: inst = 32'hca08125;
      98594: inst = 32'h13e00001;
      98595: inst = 32'hfe0d96a;
      98596: inst = 32'h5be00000;
      98597: inst = 32'h8c50000;
      98598: inst = 32'h24612800;
      98599: inst = 32'h10a00000;
      98600: inst = 32'hca0000f;
      98601: inst = 32'h24822800;
      98602: inst = 32'h10a00000;
      98603: inst = 32'hca00004;
      98604: inst = 32'h38632800;
      98605: inst = 32'h38842800;
      98606: inst = 32'h10a00001;
      98607: inst = 32'hca08133;
      98608: inst = 32'h13e00001;
      98609: inst = 32'hfe0d96a;
      98610: inst = 32'h5be00000;
      98611: inst = 32'h8c50000;
      98612: inst = 32'h24612800;
      98613: inst = 32'h10a00000;
      98614: inst = 32'hca0000f;
      98615: inst = 32'h24822800;
      98616: inst = 32'h10a00000;
      98617: inst = 32'hca00004;
      98618: inst = 32'h38632800;
      98619: inst = 32'h38842800;
      98620: inst = 32'h10a00001;
      98621: inst = 32'hca08141;
      98622: inst = 32'h13e00001;
      98623: inst = 32'hfe0d96a;
      98624: inst = 32'h5be00000;
      98625: inst = 32'h8c50000;
      98626: inst = 32'h24612800;
      98627: inst = 32'h10a00000;
      98628: inst = 32'hca0000f;
      98629: inst = 32'h24822800;
      98630: inst = 32'h10a00000;
      98631: inst = 32'hca00004;
      98632: inst = 32'h38632800;
      98633: inst = 32'h38842800;
      98634: inst = 32'h10a00001;
      98635: inst = 32'hca0814f;
      98636: inst = 32'h13e00001;
      98637: inst = 32'hfe0d96a;
      98638: inst = 32'h5be00000;
      98639: inst = 32'h8c50000;
      98640: inst = 32'h24612800;
      98641: inst = 32'h10a00000;
      98642: inst = 32'hca0000f;
      98643: inst = 32'h24822800;
      98644: inst = 32'h10a00000;
      98645: inst = 32'hca00004;
      98646: inst = 32'h38632800;
      98647: inst = 32'h38842800;
      98648: inst = 32'h10a00001;
      98649: inst = 32'hca0815d;
      98650: inst = 32'h13e00001;
      98651: inst = 32'hfe0d96a;
      98652: inst = 32'h5be00000;
      98653: inst = 32'h8c50000;
      98654: inst = 32'h24612800;
      98655: inst = 32'h10a00000;
      98656: inst = 32'hca0000f;
      98657: inst = 32'h24822800;
      98658: inst = 32'h10a00000;
      98659: inst = 32'hca00004;
      98660: inst = 32'h38632800;
      98661: inst = 32'h38842800;
      98662: inst = 32'h10a00001;
      98663: inst = 32'hca0816b;
      98664: inst = 32'h13e00001;
      98665: inst = 32'hfe0d96a;
      98666: inst = 32'h5be00000;
      98667: inst = 32'h8c50000;
      98668: inst = 32'h24612800;
      98669: inst = 32'h10a00000;
      98670: inst = 32'hca0000f;
      98671: inst = 32'h24822800;
      98672: inst = 32'h10a00000;
      98673: inst = 32'hca00004;
      98674: inst = 32'h38632800;
      98675: inst = 32'h38842800;
      98676: inst = 32'h10a00001;
      98677: inst = 32'hca08179;
      98678: inst = 32'h13e00001;
      98679: inst = 32'hfe0d96a;
      98680: inst = 32'h5be00000;
      98681: inst = 32'h8c50000;
      98682: inst = 32'h24612800;
      98683: inst = 32'h10a00000;
      98684: inst = 32'hca0000f;
      98685: inst = 32'h24822800;
      98686: inst = 32'h10a00000;
      98687: inst = 32'hca00004;
      98688: inst = 32'h38632800;
      98689: inst = 32'h38842800;
      98690: inst = 32'h10a00001;
      98691: inst = 32'hca08187;
      98692: inst = 32'h13e00001;
      98693: inst = 32'hfe0d96a;
      98694: inst = 32'h5be00000;
      98695: inst = 32'h8c50000;
      98696: inst = 32'h24612800;
      98697: inst = 32'h10a00000;
      98698: inst = 32'hca0000f;
      98699: inst = 32'h24822800;
      98700: inst = 32'h10a00000;
      98701: inst = 32'hca00004;
      98702: inst = 32'h38632800;
      98703: inst = 32'h38842800;
      98704: inst = 32'h10a00001;
      98705: inst = 32'hca08195;
      98706: inst = 32'h13e00001;
      98707: inst = 32'hfe0d96a;
      98708: inst = 32'h5be00000;
      98709: inst = 32'h8c50000;
      98710: inst = 32'h24612800;
      98711: inst = 32'h10a00000;
      98712: inst = 32'hca0000f;
      98713: inst = 32'h24822800;
      98714: inst = 32'h10a00000;
      98715: inst = 32'hca00004;
      98716: inst = 32'h38632800;
      98717: inst = 32'h38842800;
      98718: inst = 32'h10a00001;
      98719: inst = 32'hca081a3;
      98720: inst = 32'h13e00001;
      98721: inst = 32'hfe0d96a;
      98722: inst = 32'h5be00000;
      98723: inst = 32'h8c50000;
      98724: inst = 32'h24612800;
      98725: inst = 32'h10a00000;
      98726: inst = 32'hca0000f;
      98727: inst = 32'h24822800;
      98728: inst = 32'h10a00000;
      98729: inst = 32'hca00004;
      98730: inst = 32'h38632800;
      98731: inst = 32'h38842800;
      98732: inst = 32'h10a00001;
      98733: inst = 32'hca081b1;
      98734: inst = 32'h13e00001;
      98735: inst = 32'hfe0d96a;
      98736: inst = 32'h5be00000;
      98737: inst = 32'h8c50000;
      98738: inst = 32'h24612800;
      98739: inst = 32'h10a00000;
      98740: inst = 32'hca0000f;
      98741: inst = 32'h24822800;
      98742: inst = 32'h10a00000;
      98743: inst = 32'hca00004;
      98744: inst = 32'h38632800;
      98745: inst = 32'h38842800;
      98746: inst = 32'h10a00001;
      98747: inst = 32'hca081bf;
      98748: inst = 32'h13e00001;
      98749: inst = 32'hfe0d96a;
      98750: inst = 32'h5be00000;
      98751: inst = 32'h8c50000;
      98752: inst = 32'h24612800;
      98753: inst = 32'h10a00000;
      98754: inst = 32'hca0000f;
      98755: inst = 32'h24822800;
      98756: inst = 32'h10a00000;
      98757: inst = 32'hca00004;
      98758: inst = 32'h38632800;
      98759: inst = 32'h38842800;
      98760: inst = 32'h10a00001;
      98761: inst = 32'hca081cd;
      98762: inst = 32'h13e00001;
      98763: inst = 32'hfe0d96a;
      98764: inst = 32'h5be00000;
      98765: inst = 32'h8c50000;
      98766: inst = 32'h24612800;
      98767: inst = 32'h10a00000;
      98768: inst = 32'hca0000f;
      98769: inst = 32'h24822800;
      98770: inst = 32'h10a00000;
      98771: inst = 32'hca00004;
      98772: inst = 32'h38632800;
      98773: inst = 32'h38842800;
      98774: inst = 32'h10a00001;
      98775: inst = 32'hca081db;
      98776: inst = 32'h13e00001;
      98777: inst = 32'hfe0d96a;
      98778: inst = 32'h5be00000;
      98779: inst = 32'h8c50000;
      98780: inst = 32'h24612800;
      98781: inst = 32'h10a00000;
      98782: inst = 32'hca0000f;
      98783: inst = 32'h24822800;
      98784: inst = 32'h10a00000;
      98785: inst = 32'hca00004;
      98786: inst = 32'h38632800;
      98787: inst = 32'h38842800;
      98788: inst = 32'h10a00001;
      98789: inst = 32'hca081e9;
      98790: inst = 32'h13e00001;
      98791: inst = 32'hfe0d96a;
      98792: inst = 32'h5be00000;
      98793: inst = 32'h8c50000;
      98794: inst = 32'h24612800;
      98795: inst = 32'h10a00000;
      98796: inst = 32'hca0000f;
      98797: inst = 32'h24822800;
      98798: inst = 32'h10a00000;
      98799: inst = 32'hca00004;
      98800: inst = 32'h38632800;
      98801: inst = 32'h38842800;
      98802: inst = 32'h10a00001;
      98803: inst = 32'hca081f7;
      98804: inst = 32'h13e00001;
      98805: inst = 32'hfe0d96a;
      98806: inst = 32'h5be00000;
      98807: inst = 32'h8c50000;
      98808: inst = 32'h24612800;
      98809: inst = 32'h10a00000;
      98810: inst = 32'hca0000f;
      98811: inst = 32'h24822800;
      98812: inst = 32'h10a00000;
      98813: inst = 32'hca00004;
      98814: inst = 32'h38632800;
      98815: inst = 32'h38842800;
      98816: inst = 32'h10a00001;
      98817: inst = 32'hca08205;
      98818: inst = 32'h13e00001;
      98819: inst = 32'hfe0d96a;
      98820: inst = 32'h5be00000;
      98821: inst = 32'h8c50000;
      98822: inst = 32'h24612800;
      98823: inst = 32'h10a00000;
      98824: inst = 32'hca0000f;
      98825: inst = 32'h24822800;
      98826: inst = 32'h10a00000;
      98827: inst = 32'hca00004;
      98828: inst = 32'h38632800;
      98829: inst = 32'h38842800;
      98830: inst = 32'h10a00001;
      98831: inst = 32'hca08213;
      98832: inst = 32'h13e00001;
      98833: inst = 32'hfe0d96a;
      98834: inst = 32'h5be00000;
      98835: inst = 32'h8c50000;
      98836: inst = 32'h24612800;
      98837: inst = 32'h10a00000;
      98838: inst = 32'hca0000f;
      98839: inst = 32'h24822800;
      98840: inst = 32'h10a00000;
      98841: inst = 32'hca00004;
      98842: inst = 32'h38632800;
      98843: inst = 32'h38842800;
      98844: inst = 32'h10a00001;
      98845: inst = 32'hca08221;
      98846: inst = 32'h13e00001;
      98847: inst = 32'hfe0d96a;
      98848: inst = 32'h5be00000;
      98849: inst = 32'h8c50000;
      98850: inst = 32'h24612800;
      98851: inst = 32'h10a00000;
      98852: inst = 32'hca0000f;
      98853: inst = 32'h24822800;
      98854: inst = 32'h10a00000;
      98855: inst = 32'hca00004;
      98856: inst = 32'h38632800;
      98857: inst = 32'h38842800;
      98858: inst = 32'h10a00001;
      98859: inst = 32'hca0822f;
      98860: inst = 32'h13e00001;
      98861: inst = 32'hfe0d96a;
      98862: inst = 32'h5be00000;
      98863: inst = 32'h8c50000;
      98864: inst = 32'h24612800;
      98865: inst = 32'h10a00000;
      98866: inst = 32'hca0000f;
      98867: inst = 32'h24822800;
      98868: inst = 32'h10a00000;
      98869: inst = 32'hca00004;
      98870: inst = 32'h38632800;
      98871: inst = 32'h38842800;
      98872: inst = 32'h10a00001;
      98873: inst = 32'hca0823d;
      98874: inst = 32'h13e00001;
      98875: inst = 32'hfe0d96a;
      98876: inst = 32'h5be00000;
      98877: inst = 32'h8c50000;
      98878: inst = 32'h24612800;
      98879: inst = 32'h10a00000;
      98880: inst = 32'hca0000f;
      98881: inst = 32'h24822800;
      98882: inst = 32'h10a00000;
      98883: inst = 32'hca00004;
      98884: inst = 32'h38632800;
      98885: inst = 32'h38842800;
      98886: inst = 32'h10a00001;
      98887: inst = 32'hca0824b;
      98888: inst = 32'h13e00001;
      98889: inst = 32'hfe0d96a;
      98890: inst = 32'h5be00000;
      98891: inst = 32'h8c50000;
      98892: inst = 32'h24612800;
      98893: inst = 32'h10a00000;
      98894: inst = 32'hca0000f;
      98895: inst = 32'h24822800;
      98896: inst = 32'h10a00000;
      98897: inst = 32'hca00004;
      98898: inst = 32'h38632800;
      98899: inst = 32'h38842800;
      98900: inst = 32'h10a00001;
      98901: inst = 32'hca08259;
      98902: inst = 32'h13e00001;
      98903: inst = 32'hfe0d96a;
      98904: inst = 32'h5be00000;
      98905: inst = 32'h8c50000;
      98906: inst = 32'h24612800;
      98907: inst = 32'h10a00000;
      98908: inst = 32'hca0000f;
      98909: inst = 32'h24822800;
      98910: inst = 32'h10a00000;
      98911: inst = 32'hca00004;
      98912: inst = 32'h38632800;
      98913: inst = 32'h38842800;
      98914: inst = 32'h10a00001;
      98915: inst = 32'hca08267;
      98916: inst = 32'h13e00001;
      98917: inst = 32'hfe0d96a;
      98918: inst = 32'h5be00000;
      98919: inst = 32'h8c50000;
      98920: inst = 32'h24612800;
      98921: inst = 32'h10a00000;
      98922: inst = 32'hca0000f;
      98923: inst = 32'h24822800;
      98924: inst = 32'h10a00000;
      98925: inst = 32'hca00004;
      98926: inst = 32'h38632800;
      98927: inst = 32'h38842800;
      98928: inst = 32'h10a00001;
      98929: inst = 32'hca08275;
      98930: inst = 32'h13e00001;
      98931: inst = 32'hfe0d96a;
      98932: inst = 32'h5be00000;
      98933: inst = 32'h8c50000;
      98934: inst = 32'h24612800;
      98935: inst = 32'h10a00000;
      98936: inst = 32'hca0000f;
      98937: inst = 32'h24822800;
      98938: inst = 32'h10a00000;
      98939: inst = 32'hca00004;
      98940: inst = 32'h38632800;
      98941: inst = 32'h38842800;
      98942: inst = 32'h10a00001;
      98943: inst = 32'hca08283;
      98944: inst = 32'h13e00001;
      98945: inst = 32'hfe0d96a;
      98946: inst = 32'h5be00000;
      98947: inst = 32'h8c50000;
      98948: inst = 32'h24612800;
      98949: inst = 32'h10a00000;
      98950: inst = 32'hca0000f;
      98951: inst = 32'h24822800;
      98952: inst = 32'h10a00000;
      98953: inst = 32'hca00004;
      98954: inst = 32'h38632800;
      98955: inst = 32'h38842800;
      98956: inst = 32'h10a00001;
      98957: inst = 32'hca08291;
      98958: inst = 32'h13e00001;
      98959: inst = 32'hfe0d96a;
      98960: inst = 32'h5be00000;
      98961: inst = 32'h8c50000;
      98962: inst = 32'h24612800;
      98963: inst = 32'h10a00000;
      98964: inst = 32'hca0000f;
      98965: inst = 32'h24822800;
      98966: inst = 32'h10a00000;
      98967: inst = 32'hca00004;
      98968: inst = 32'h38632800;
      98969: inst = 32'h38842800;
      98970: inst = 32'h10a00001;
      98971: inst = 32'hca0829f;
      98972: inst = 32'h13e00001;
      98973: inst = 32'hfe0d96a;
      98974: inst = 32'h5be00000;
      98975: inst = 32'h8c50000;
      98976: inst = 32'h24612800;
      98977: inst = 32'h10a00000;
      98978: inst = 32'hca0000f;
      98979: inst = 32'h24822800;
      98980: inst = 32'h10a00000;
      98981: inst = 32'hca00004;
      98982: inst = 32'h38632800;
      98983: inst = 32'h38842800;
      98984: inst = 32'h10a00001;
      98985: inst = 32'hca082ad;
      98986: inst = 32'h13e00001;
      98987: inst = 32'hfe0d96a;
      98988: inst = 32'h5be00000;
      98989: inst = 32'h8c50000;
      98990: inst = 32'h24612800;
      98991: inst = 32'h10a00000;
      98992: inst = 32'hca0000f;
      98993: inst = 32'h24822800;
      98994: inst = 32'h10a00000;
      98995: inst = 32'hca00004;
      98996: inst = 32'h38632800;
      98997: inst = 32'h38842800;
      98998: inst = 32'h10a00001;
      98999: inst = 32'hca082bb;
      99000: inst = 32'h13e00001;
      99001: inst = 32'hfe0d96a;
      99002: inst = 32'h5be00000;
      99003: inst = 32'h8c50000;
      99004: inst = 32'h24612800;
      99005: inst = 32'h10a00000;
      99006: inst = 32'hca0000f;
      99007: inst = 32'h24822800;
      99008: inst = 32'h10a00000;
      99009: inst = 32'hca00004;
      99010: inst = 32'h38632800;
      99011: inst = 32'h38842800;
      99012: inst = 32'h10a00001;
      99013: inst = 32'hca082c9;
      99014: inst = 32'h13e00001;
      99015: inst = 32'hfe0d96a;
      99016: inst = 32'h5be00000;
      99017: inst = 32'h8c50000;
      99018: inst = 32'h24612800;
      99019: inst = 32'h10a00000;
      99020: inst = 32'hca0000f;
      99021: inst = 32'h24822800;
      99022: inst = 32'h10a00000;
      99023: inst = 32'hca00004;
      99024: inst = 32'h38632800;
      99025: inst = 32'h38842800;
      99026: inst = 32'h10a00001;
      99027: inst = 32'hca082d7;
      99028: inst = 32'h13e00001;
      99029: inst = 32'hfe0d96a;
      99030: inst = 32'h5be00000;
      99031: inst = 32'h8c50000;
      99032: inst = 32'h24612800;
      99033: inst = 32'h10a00000;
      99034: inst = 32'hca0000f;
      99035: inst = 32'h24822800;
      99036: inst = 32'h10a00000;
      99037: inst = 32'hca00004;
      99038: inst = 32'h38632800;
      99039: inst = 32'h38842800;
      99040: inst = 32'h10a00001;
      99041: inst = 32'hca082e5;
      99042: inst = 32'h13e00001;
      99043: inst = 32'hfe0d96a;
      99044: inst = 32'h5be00000;
      99045: inst = 32'h8c50000;
      99046: inst = 32'h24612800;
      99047: inst = 32'h10a00000;
      99048: inst = 32'hca0000f;
      99049: inst = 32'h24822800;
      99050: inst = 32'h10a00000;
      99051: inst = 32'hca00004;
      99052: inst = 32'h38632800;
      99053: inst = 32'h38842800;
      99054: inst = 32'h10a00001;
      99055: inst = 32'hca082f3;
      99056: inst = 32'h13e00001;
      99057: inst = 32'hfe0d96a;
      99058: inst = 32'h5be00000;
      99059: inst = 32'h8c50000;
      99060: inst = 32'h24612800;
      99061: inst = 32'h10a00000;
      99062: inst = 32'hca0000f;
      99063: inst = 32'h24822800;
      99064: inst = 32'h10a00000;
      99065: inst = 32'hca00004;
      99066: inst = 32'h38632800;
      99067: inst = 32'h38842800;
      99068: inst = 32'h10a00001;
      99069: inst = 32'hca08301;
      99070: inst = 32'h13e00001;
      99071: inst = 32'hfe0d96a;
      99072: inst = 32'h5be00000;
      99073: inst = 32'h8c50000;
      99074: inst = 32'h24612800;
      99075: inst = 32'h10a00000;
      99076: inst = 32'hca0000f;
      99077: inst = 32'h24822800;
      99078: inst = 32'h10a00000;
      99079: inst = 32'hca00004;
      99080: inst = 32'h38632800;
      99081: inst = 32'h38842800;
      99082: inst = 32'h10a00001;
      99083: inst = 32'hca0830f;
      99084: inst = 32'h13e00001;
      99085: inst = 32'hfe0d96a;
      99086: inst = 32'h5be00000;
      99087: inst = 32'h8c50000;
      99088: inst = 32'h24612800;
      99089: inst = 32'h10a00000;
      99090: inst = 32'hca0000f;
      99091: inst = 32'h24822800;
      99092: inst = 32'h10a00000;
      99093: inst = 32'hca00004;
      99094: inst = 32'h38632800;
      99095: inst = 32'h38842800;
      99096: inst = 32'h10a00001;
      99097: inst = 32'hca0831d;
      99098: inst = 32'h13e00001;
      99099: inst = 32'hfe0d96a;
      99100: inst = 32'h5be00000;
      99101: inst = 32'h8c50000;
      99102: inst = 32'h24612800;
      99103: inst = 32'h10a00000;
      99104: inst = 32'hca0000f;
      99105: inst = 32'h24822800;
      99106: inst = 32'h10a00000;
      99107: inst = 32'hca00004;
      99108: inst = 32'h38632800;
      99109: inst = 32'h38842800;
      99110: inst = 32'h10a00001;
      99111: inst = 32'hca0832b;
      99112: inst = 32'h13e00001;
      99113: inst = 32'hfe0d96a;
      99114: inst = 32'h5be00000;
      99115: inst = 32'h8c50000;
      99116: inst = 32'h24612800;
      99117: inst = 32'h10a00000;
      99118: inst = 32'hca0000f;
      99119: inst = 32'h24822800;
      99120: inst = 32'h10a00000;
      99121: inst = 32'hca00004;
      99122: inst = 32'h38632800;
      99123: inst = 32'h38842800;
      99124: inst = 32'h10a00001;
      99125: inst = 32'hca08339;
      99126: inst = 32'h13e00001;
      99127: inst = 32'hfe0d96a;
      99128: inst = 32'h5be00000;
      99129: inst = 32'h8c50000;
      99130: inst = 32'h24612800;
      99131: inst = 32'h10a00000;
      99132: inst = 32'hca0000f;
      99133: inst = 32'h24822800;
      99134: inst = 32'h10a00000;
      99135: inst = 32'hca00004;
      99136: inst = 32'h38632800;
      99137: inst = 32'h38842800;
      99138: inst = 32'h10a00001;
      99139: inst = 32'hca08347;
      99140: inst = 32'h13e00001;
      99141: inst = 32'hfe0d96a;
      99142: inst = 32'h5be00000;
      99143: inst = 32'h8c50000;
      99144: inst = 32'h24612800;
      99145: inst = 32'h10a00000;
      99146: inst = 32'hca0000f;
      99147: inst = 32'h24822800;
      99148: inst = 32'h10a00000;
      99149: inst = 32'hca00004;
      99150: inst = 32'h38632800;
      99151: inst = 32'h38842800;
      99152: inst = 32'h10a00001;
      99153: inst = 32'hca08355;
      99154: inst = 32'h13e00001;
      99155: inst = 32'hfe0d96a;
      99156: inst = 32'h5be00000;
      99157: inst = 32'h8c50000;
      99158: inst = 32'h24612800;
      99159: inst = 32'h10a00000;
      99160: inst = 32'hca0000f;
      99161: inst = 32'h24822800;
      99162: inst = 32'h10a00000;
      99163: inst = 32'hca00004;
      99164: inst = 32'h38632800;
      99165: inst = 32'h38842800;
      99166: inst = 32'h10a00001;
      99167: inst = 32'hca08363;
      99168: inst = 32'h13e00001;
      99169: inst = 32'hfe0d96a;
      99170: inst = 32'h5be00000;
      99171: inst = 32'h8c50000;
      99172: inst = 32'h24612800;
      99173: inst = 32'h10a00000;
      99174: inst = 32'hca0000f;
      99175: inst = 32'h24822800;
      99176: inst = 32'h10a00000;
      99177: inst = 32'hca00004;
      99178: inst = 32'h38632800;
      99179: inst = 32'h38842800;
      99180: inst = 32'h10a00001;
      99181: inst = 32'hca08371;
      99182: inst = 32'h13e00001;
      99183: inst = 32'hfe0d96a;
      99184: inst = 32'h5be00000;
      99185: inst = 32'h8c50000;
      99186: inst = 32'h24612800;
      99187: inst = 32'h10a00000;
      99188: inst = 32'hca0000f;
      99189: inst = 32'h24822800;
      99190: inst = 32'h10a00000;
      99191: inst = 32'hca00004;
      99192: inst = 32'h38632800;
      99193: inst = 32'h38842800;
      99194: inst = 32'h10a00001;
      99195: inst = 32'hca0837f;
      99196: inst = 32'h13e00001;
      99197: inst = 32'hfe0d96a;
      99198: inst = 32'h5be00000;
      99199: inst = 32'h8c50000;
      99200: inst = 32'h24612800;
      99201: inst = 32'h10a00000;
      99202: inst = 32'hca0000f;
      99203: inst = 32'h24822800;
      99204: inst = 32'h10a00000;
      99205: inst = 32'hca00004;
      99206: inst = 32'h38632800;
      99207: inst = 32'h38842800;
      99208: inst = 32'h10a00001;
      99209: inst = 32'hca0838d;
      99210: inst = 32'h13e00001;
      99211: inst = 32'hfe0d96a;
      99212: inst = 32'h5be00000;
      99213: inst = 32'h8c50000;
      99214: inst = 32'h24612800;
      99215: inst = 32'h10a00000;
      99216: inst = 32'hca0000f;
      99217: inst = 32'h24822800;
      99218: inst = 32'h10a00000;
      99219: inst = 32'hca00004;
      99220: inst = 32'h38632800;
      99221: inst = 32'h38842800;
      99222: inst = 32'h10a00001;
      99223: inst = 32'hca0839b;
      99224: inst = 32'h13e00001;
      99225: inst = 32'hfe0d96a;
      99226: inst = 32'h5be00000;
      99227: inst = 32'h8c50000;
      99228: inst = 32'h24612800;
      99229: inst = 32'h10a00000;
      99230: inst = 32'hca0000f;
      99231: inst = 32'h24822800;
      99232: inst = 32'h10a00000;
      99233: inst = 32'hca00004;
      99234: inst = 32'h38632800;
      99235: inst = 32'h38842800;
      99236: inst = 32'h10a00001;
      99237: inst = 32'hca083a9;
      99238: inst = 32'h13e00001;
      99239: inst = 32'hfe0d96a;
      99240: inst = 32'h5be00000;
      99241: inst = 32'h8c50000;
      99242: inst = 32'h24612800;
      99243: inst = 32'h10a00000;
      99244: inst = 32'hca0000f;
      99245: inst = 32'h24822800;
      99246: inst = 32'h10a00000;
      99247: inst = 32'hca00004;
      99248: inst = 32'h38632800;
      99249: inst = 32'h38842800;
      99250: inst = 32'h10a00001;
      99251: inst = 32'hca083b7;
      99252: inst = 32'h13e00001;
      99253: inst = 32'hfe0d96a;
      99254: inst = 32'h5be00000;
      99255: inst = 32'h8c50000;
      99256: inst = 32'h24612800;
      99257: inst = 32'h10a00000;
      99258: inst = 32'hca0000f;
      99259: inst = 32'h24822800;
      99260: inst = 32'h10a00000;
      99261: inst = 32'hca00004;
      99262: inst = 32'h38632800;
      99263: inst = 32'h38842800;
      99264: inst = 32'h10a00001;
      99265: inst = 32'hca083c5;
      99266: inst = 32'h13e00001;
      99267: inst = 32'hfe0d96a;
      99268: inst = 32'h5be00000;
      99269: inst = 32'h8c50000;
      99270: inst = 32'h24612800;
      99271: inst = 32'h10a00000;
      99272: inst = 32'hca0000f;
      99273: inst = 32'h24822800;
      99274: inst = 32'h10a00000;
      99275: inst = 32'hca00004;
      99276: inst = 32'h38632800;
      99277: inst = 32'h38842800;
      99278: inst = 32'h10a00001;
      99279: inst = 32'hca083d3;
      99280: inst = 32'h13e00001;
      99281: inst = 32'hfe0d96a;
      99282: inst = 32'h5be00000;
      99283: inst = 32'h8c50000;
      99284: inst = 32'h24612800;
      99285: inst = 32'h10a00000;
      99286: inst = 32'hca0000f;
      99287: inst = 32'h24822800;
      99288: inst = 32'h10a00000;
      99289: inst = 32'hca00004;
      99290: inst = 32'h38632800;
      99291: inst = 32'h38842800;
      99292: inst = 32'h10a00001;
      99293: inst = 32'hca083e1;
      99294: inst = 32'h13e00001;
      99295: inst = 32'hfe0d96a;
      99296: inst = 32'h5be00000;
      99297: inst = 32'h8c50000;
      99298: inst = 32'h24612800;
      99299: inst = 32'h10a00000;
      99300: inst = 32'hca0000f;
      99301: inst = 32'h24822800;
      99302: inst = 32'h10a00000;
      99303: inst = 32'hca00004;
      99304: inst = 32'h38632800;
      99305: inst = 32'h38842800;
      99306: inst = 32'h10a00001;
      99307: inst = 32'hca083ef;
      99308: inst = 32'h13e00001;
      99309: inst = 32'hfe0d96a;
      99310: inst = 32'h5be00000;
      99311: inst = 32'h8c50000;
      99312: inst = 32'h24612800;
      99313: inst = 32'h10a00000;
      99314: inst = 32'hca0000f;
      99315: inst = 32'h24822800;
      99316: inst = 32'h10a00000;
      99317: inst = 32'hca00004;
      99318: inst = 32'h38632800;
      99319: inst = 32'h38842800;
      99320: inst = 32'h10a00001;
      99321: inst = 32'hca083fd;
      99322: inst = 32'h13e00001;
      99323: inst = 32'hfe0d96a;
      99324: inst = 32'h5be00000;
      99325: inst = 32'h8c50000;
      99326: inst = 32'h24612800;
      99327: inst = 32'h10a00000;
      99328: inst = 32'hca0000f;
      99329: inst = 32'h24822800;
      99330: inst = 32'h10a00000;
      99331: inst = 32'hca00004;
      99332: inst = 32'h38632800;
      99333: inst = 32'h38842800;
      99334: inst = 32'h10a00001;
      99335: inst = 32'hca0840b;
      99336: inst = 32'h13e00001;
      99337: inst = 32'hfe0d96a;
      99338: inst = 32'h5be00000;
      99339: inst = 32'h8c50000;
      99340: inst = 32'h24612800;
      99341: inst = 32'h10a00000;
      99342: inst = 32'hca0000f;
      99343: inst = 32'h24822800;
      99344: inst = 32'h10a00000;
      99345: inst = 32'hca00004;
      99346: inst = 32'h38632800;
      99347: inst = 32'h38842800;
      99348: inst = 32'h10a00001;
      99349: inst = 32'hca08419;
      99350: inst = 32'h13e00001;
      99351: inst = 32'hfe0d96a;
      99352: inst = 32'h5be00000;
      99353: inst = 32'h8c50000;
      99354: inst = 32'h24612800;
      99355: inst = 32'h10a00000;
      99356: inst = 32'hca0000f;
      99357: inst = 32'h24822800;
      99358: inst = 32'h10a00000;
      99359: inst = 32'hca00004;
      99360: inst = 32'h38632800;
      99361: inst = 32'h38842800;
      99362: inst = 32'h10a00001;
      99363: inst = 32'hca08427;
      99364: inst = 32'h13e00001;
      99365: inst = 32'hfe0d96a;
      99366: inst = 32'h5be00000;
      99367: inst = 32'h8c50000;
      99368: inst = 32'h24612800;
      99369: inst = 32'h10a00000;
      99370: inst = 32'hca0000f;
      99371: inst = 32'h24822800;
      99372: inst = 32'h10a00000;
      99373: inst = 32'hca00004;
      99374: inst = 32'h38632800;
      99375: inst = 32'h38842800;
      99376: inst = 32'h10a00001;
      99377: inst = 32'hca08435;
      99378: inst = 32'h13e00001;
      99379: inst = 32'hfe0d96a;
      99380: inst = 32'h5be00000;
      99381: inst = 32'h8c50000;
      99382: inst = 32'h24612800;
      99383: inst = 32'h10a00000;
      99384: inst = 32'hca0000f;
      99385: inst = 32'h24822800;
      99386: inst = 32'h10a00000;
      99387: inst = 32'hca00004;
      99388: inst = 32'h38632800;
      99389: inst = 32'h38842800;
      99390: inst = 32'h10a00001;
      99391: inst = 32'hca08443;
      99392: inst = 32'h13e00001;
      99393: inst = 32'hfe0d96a;
      99394: inst = 32'h5be00000;
      99395: inst = 32'h8c50000;
      99396: inst = 32'h24612800;
      99397: inst = 32'h10a00000;
      99398: inst = 32'hca0000f;
      99399: inst = 32'h24822800;
      99400: inst = 32'h10a00000;
      99401: inst = 32'hca00004;
      99402: inst = 32'h38632800;
      99403: inst = 32'h38842800;
      99404: inst = 32'h10a00001;
      99405: inst = 32'hca08451;
      99406: inst = 32'h13e00001;
      99407: inst = 32'hfe0d96a;
      99408: inst = 32'h5be00000;
      99409: inst = 32'h8c50000;
      99410: inst = 32'h24612800;
      99411: inst = 32'h10a00000;
      99412: inst = 32'hca0000f;
      99413: inst = 32'h24822800;
      99414: inst = 32'h10a00000;
      99415: inst = 32'hca00004;
      99416: inst = 32'h38632800;
      99417: inst = 32'h38842800;
      99418: inst = 32'h10a00001;
      99419: inst = 32'hca0845f;
      99420: inst = 32'h13e00001;
      99421: inst = 32'hfe0d96a;
      99422: inst = 32'h5be00000;
      99423: inst = 32'h8c50000;
      99424: inst = 32'h24612800;
      99425: inst = 32'h10a00000;
      99426: inst = 32'hca0000f;
      99427: inst = 32'h24822800;
      99428: inst = 32'h10a00000;
      99429: inst = 32'hca00004;
      99430: inst = 32'h38632800;
      99431: inst = 32'h38842800;
      99432: inst = 32'h10a00001;
      99433: inst = 32'hca0846d;
      99434: inst = 32'h13e00001;
      99435: inst = 32'hfe0d96a;
      99436: inst = 32'h5be00000;
      99437: inst = 32'h8c50000;
      99438: inst = 32'h24612800;
      99439: inst = 32'h10a00000;
      99440: inst = 32'hca0000f;
      99441: inst = 32'h24822800;
      99442: inst = 32'h10a00000;
      99443: inst = 32'hca00004;
      99444: inst = 32'h38632800;
      99445: inst = 32'h38842800;
      99446: inst = 32'h10a00001;
      99447: inst = 32'hca0847b;
      99448: inst = 32'h13e00001;
      99449: inst = 32'hfe0d96a;
      99450: inst = 32'h5be00000;
      99451: inst = 32'h8c50000;
      99452: inst = 32'h24612800;
      99453: inst = 32'h10a00000;
      99454: inst = 32'hca0000f;
      99455: inst = 32'h24822800;
      99456: inst = 32'h10a00000;
      99457: inst = 32'hca00004;
      99458: inst = 32'h38632800;
      99459: inst = 32'h38842800;
      99460: inst = 32'h10a00001;
      99461: inst = 32'hca08489;
      99462: inst = 32'h13e00001;
      99463: inst = 32'hfe0d96a;
      99464: inst = 32'h5be00000;
      99465: inst = 32'h8c50000;
      99466: inst = 32'h24612800;
      99467: inst = 32'h10a00000;
      99468: inst = 32'hca0000f;
      99469: inst = 32'h24822800;
      99470: inst = 32'h10a00000;
      99471: inst = 32'hca00004;
      99472: inst = 32'h38632800;
      99473: inst = 32'h38842800;
      99474: inst = 32'h10a00001;
      99475: inst = 32'hca08497;
      99476: inst = 32'h13e00001;
      99477: inst = 32'hfe0d96a;
      99478: inst = 32'h5be00000;
      99479: inst = 32'h8c50000;
      99480: inst = 32'h24612800;
      99481: inst = 32'h10a00000;
      99482: inst = 32'hca0000f;
      99483: inst = 32'h24822800;
      99484: inst = 32'h10a00000;
      99485: inst = 32'hca00004;
      99486: inst = 32'h38632800;
      99487: inst = 32'h38842800;
      99488: inst = 32'h10a00001;
      99489: inst = 32'hca084a5;
      99490: inst = 32'h13e00001;
      99491: inst = 32'hfe0d96a;
      99492: inst = 32'h5be00000;
      99493: inst = 32'h8c50000;
      99494: inst = 32'h24612800;
      99495: inst = 32'h10a00000;
      99496: inst = 32'hca0000f;
      99497: inst = 32'h24822800;
      99498: inst = 32'h10a00000;
      99499: inst = 32'hca00004;
      99500: inst = 32'h38632800;
      99501: inst = 32'h38842800;
      99502: inst = 32'h10a00001;
      99503: inst = 32'hca084b3;
      99504: inst = 32'h13e00001;
      99505: inst = 32'hfe0d96a;
      99506: inst = 32'h5be00000;
      99507: inst = 32'h8c50000;
      99508: inst = 32'h24612800;
      99509: inst = 32'h10a00000;
      99510: inst = 32'hca0000f;
      99511: inst = 32'h24822800;
      99512: inst = 32'h10a00000;
      99513: inst = 32'hca00004;
      99514: inst = 32'h38632800;
      99515: inst = 32'h38842800;
      99516: inst = 32'h10a00001;
      99517: inst = 32'hca084c1;
      99518: inst = 32'h13e00001;
      99519: inst = 32'hfe0d96a;
      99520: inst = 32'h5be00000;
      99521: inst = 32'h8c50000;
      99522: inst = 32'h24612800;
      99523: inst = 32'h10a00000;
      99524: inst = 32'hca0000f;
      99525: inst = 32'h24822800;
      99526: inst = 32'h10a00000;
      99527: inst = 32'hca00004;
      99528: inst = 32'h38632800;
      99529: inst = 32'h38842800;
      99530: inst = 32'h10a00001;
      99531: inst = 32'hca084cf;
      99532: inst = 32'h13e00001;
      99533: inst = 32'hfe0d96a;
      99534: inst = 32'h5be00000;
      99535: inst = 32'h8c50000;
      99536: inst = 32'h24612800;
      99537: inst = 32'h10a00000;
      99538: inst = 32'hca0000f;
      99539: inst = 32'h24822800;
      99540: inst = 32'h10a00000;
      99541: inst = 32'hca00004;
      99542: inst = 32'h38632800;
      99543: inst = 32'h38842800;
      99544: inst = 32'h10a00001;
      99545: inst = 32'hca084dd;
      99546: inst = 32'h13e00001;
      99547: inst = 32'hfe0d96a;
      99548: inst = 32'h5be00000;
      99549: inst = 32'h8c50000;
      99550: inst = 32'h24612800;
      99551: inst = 32'h10a00000;
      99552: inst = 32'hca0000f;
      99553: inst = 32'h24822800;
      99554: inst = 32'h10a00000;
      99555: inst = 32'hca00004;
      99556: inst = 32'h38632800;
      99557: inst = 32'h38842800;
      99558: inst = 32'h10a00001;
      99559: inst = 32'hca084eb;
      99560: inst = 32'h13e00001;
      99561: inst = 32'hfe0d96a;
      99562: inst = 32'h5be00000;
      99563: inst = 32'h8c50000;
      99564: inst = 32'h24612800;
      99565: inst = 32'h10a00000;
      99566: inst = 32'hca0000f;
      99567: inst = 32'h24822800;
      99568: inst = 32'h10a00000;
      99569: inst = 32'hca00004;
      99570: inst = 32'h38632800;
      99571: inst = 32'h38842800;
      99572: inst = 32'h10a00001;
      99573: inst = 32'hca084f9;
      99574: inst = 32'h13e00001;
      99575: inst = 32'hfe0d96a;
      99576: inst = 32'h5be00000;
      99577: inst = 32'h8c50000;
      99578: inst = 32'h24612800;
      99579: inst = 32'h10a00000;
      99580: inst = 32'hca0000f;
      99581: inst = 32'h24822800;
      99582: inst = 32'h10a00000;
      99583: inst = 32'hca00004;
      99584: inst = 32'h38632800;
      99585: inst = 32'h38842800;
      99586: inst = 32'h10a00001;
      99587: inst = 32'hca08507;
      99588: inst = 32'h13e00001;
      99589: inst = 32'hfe0d96a;
      99590: inst = 32'h5be00000;
      99591: inst = 32'h8c50000;
      99592: inst = 32'h24612800;
      99593: inst = 32'h10a00000;
      99594: inst = 32'hca0000f;
      99595: inst = 32'h24822800;
      99596: inst = 32'h10a00000;
      99597: inst = 32'hca00004;
      99598: inst = 32'h38632800;
      99599: inst = 32'h38842800;
      99600: inst = 32'h10a00001;
      99601: inst = 32'hca08515;
      99602: inst = 32'h13e00001;
      99603: inst = 32'hfe0d96a;
      99604: inst = 32'h5be00000;
      99605: inst = 32'h8c50000;
      99606: inst = 32'h24612800;
      99607: inst = 32'h10a00000;
      99608: inst = 32'hca0000f;
      99609: inst = 32'h24822800;
      99610: inst = 32'h10a00000;
      99611: inst = 32'hca00004;
      99612: inst = 32'h38632800;
      99613: inst = 32'h38842800;
      99614: inst = 32'h10a00001;
      99615: inst = 32'hca08523;
      99616: inst = 32'h13e00001;
      99617: inst = 32'hfe0d96a;
      99618: inst = 32'h5be00000;
      99619: inst = 32'h8c50000;
      99620: inst = 32'h24612800;
      99621: inst = 32'h10a00000;
      99622: inst = 32'hca0000f;
      99623: inst = 32'h24822800;
      99624: inst = 32'h10a00000;
      99625: inst = 32'hca00004;
      99626: inst = 32'h38632800;
      99627: inst = 32'h38842800;
      99628: inst = 32'h10a00001;
      99629: inst = 32'hca08531;
      99630: inst = 32'h13e00001;
      99631: inst = 32'hfe0d96a;
      99632: inst = 32'h5be00000;
      99633: inst = 32'h8c50000;
      99634: inst = 32'h24612800;
      99635: inst = 32'h10a00000;
      99636: inst = 32'hca0000f;
      99637: inst = 32'h24822800;
      99638: inst = 32'h10a00000;
      99639: inst = 32'hca00004;
      99640: inst = 32'h38632800;
      99641: inst = 32'h38842800;
      99642: inst = 32'h10a00001;
      99643: inst = 32'hca0853f;
      99644: inst = 32'h13e00001;
      99645: inst = 32'hfe0d96a;
      99646: inst = 32'h5be00000;
      99647: inst = 32'h8c50000;
      99648: inst = 32'h24612800;
      99649: inst = 32'h10a00000;
      99650: inst = 32'hca0000f;
      99651: inst = 32'h24822800;
      99652: inst = 32'h10a00000;
      99653: inst = 32'hca00004;
      99654: inst = 32'h38632800;
      99655: inst = 32'h38842800;
      99656: inst = 32'h10a00001;
      99657: inst = 32'hca0854d;
      99658: inst = 32'h13e00001;
      99659: inst = 32'hfe0d96a;
      99660: inst = 32'h5be00000;
      99661: inst = 32'h8c50000;
      99662: inst = 32'h24612800;
      99663: inst = 32'h10a00000;
      99664: inst = 32'hca0000f;
      99665: inst = 32'h24822800;
      99666: inst = 32'h10a00000;
      99667: inst = 32'hca00004;
      99668: inst = 32'h38632800;
      99669: inst = 32'h38842800;
      99670: inst = 32'h10a00001;
      99671: inst = 32'hca0855b;
      99672: inst = 32'h13e00001;
      99673: inst = 32'hfe0d96a;
      99674: inst = 32'h5be00000;
      99675: inst = 32'h8c50000;
      99676: inst = 32'h24612800;
      99677: inst = 32'h10a00000;
      99678: inst = 32'hca0000f;
      99679: inst = 32'h24822800;
      99680: inst = 32'h10a00000;
      99681: inst = 32'hca00004;
      99682: inst = 32'h38632800;
      99683: inst = 32'h38842800;
      99684: inst = 32'h10a00001;
      99685: inst = 32'hca08569;
      99686: inst = 32'h13e00001;
      99687: inst = 32'hfe0d96a;
      99688: inst = 32'h5be00000;
      99689: inst = 32'h8c50000;
      99690: inst = 32'h24612800;
      99691: inst = 32'h10a00000;
      99692: inst = 32'hca00010;
      99693: inst = 32'h24822800;
      99694: inst = 32'h10a00000;
      99695: inst = 32'hca00004;
      99696: inst = 32'h38632800;
      99697: inst = 32'h38842800;
      99698: inst = 32'h10a00001;
      99699: inst = 32'hca08577;
      99700: inst = 32'h13e00001;
      99701: inst = 32'hfe0d96a;
      99702: inst = 32'h5be00000;
      99703: inst = 32'h8c50000;
      99704: inst = 32'h24612800;
      99705: inst = 32'h10a00000;
      99706: inst = 32'hca00010;
      99707: inst = 32'h24822800;
      99708: inst = 32'h10a00000;
      99709: inst = 32'hca00004;
      99710: inst = 32'h38632800;
      99711: inst = 32'h38842800;
      99712: inst = 32'h10a00001;
      99713: inst = 32'hca08585;
      99714: inst = 32'h13e00001;
      99715: inst = 32'hfe0d96a;
      99716: inst = 32'h5be00000;
      99717: inst = 32'h8c50000;
      99718: inst = 32'h24612800;
      99719: inst = 32'h10a00000;
      99720: inst = 32'hca00010;
      99721: inst = 32'h24822800;
      99722: inst = 32'h10a00000;
      99723: inst = 32'hca00004;
      99724: inst = 32'h38632800;
      99725: inst = 32'h38842800;
      99726: inst = 32'h10a00001;
      99727: inst = 32'hca08593;
      99728: inst = 32'h13e00001;
      99729: inst = 32'hfe0d96a;
      99730: inst = 32'h5be00000;
      99731: inst = 32'h8c50000;
      99732: inst = 32'h24612800;
      99733: inst = 32'h10a00000;
      99734: inst = 32'hca00010;
      99735: inst = 32'h24822800;
      99736: inst = 32'h10a00000;
      99737: inst = 32'hca00004;
      99738: inst = 32'h38632800;
      99739: inst = 32'h38842800;
      99740: inst = 32'h10a00001;
      99741: inst = 32'hca085a1;
      99742: inst = 32'h13e00001;
      99743: inst = 32'hfe0d96a;
      99744: inst = 32'h5be00000;
      99745: inst = 32'h8c50000;
      99746: inst = 32'h24612800;
      99747: inst = 32'h10a00000;
      99748: inst = 32'hca00010;
      99749: inst = 32'h24822800;
      99750: inst = 32'h10a00000;
      99751: inst = 32'hca00004;
      99752: inst = 32'h38632800;
      99753: inst = 32'h38842800;
      99754: inst = 32'h10a00001;
      99755: inst = 32'hca085af;
      99756: inst = 32'h13e00001;
      99757: inst = 32'hfe0d96a;
      99758: inst = 32'h5be00000;
      99759: inst = 32'h8c50000;
      99760: inst = 32'h24612800;
      99761: inst = 32'h10a00000;
      99762: inst = 32'hca00010;
      99763: inst = 32'h24822800;
      99764: inst = 32'h10a00000;
      99765: inst = 32'hca00004;
      99766: inst = 32'h38632800;
      99767: inst = 32'h38842800;
      99768: inst = 32'h10a00001;
      99769: inst = 32'hca085bd;
      99770: inst = 32'h13e00001;
      99771: inst = 32'hfe0d96a;
      99772: inst = 32'h5be00000;
      99773: inst = 32'h8c50000;
      99774: inst = 32'h24612800;
      99775: inst = 32'h10a00000;
      99776: inst = 32'hca00010;
      99777: inst = 32'h24822800;
      99778: inst = 32'h10a00000;
      99779: inst = 32'hca00004;
      99780: inst = 32'h38632800;
      99781: inst = 32'h38842800;
      99782: inst = 32'h10a00001;
      99783: inst = 32'hca085cb;
      99784: inst = 32'h13e00001;
      99785: inst = 32'hfe0d96a;
      99786: inst = 32'h5be00000;
      99787: inst = 32'h8c50000;
      99788: inst = 32'h24612800;
      99789: inst = 32'h10a00000;
      99790: inst = 32'hca00010;
      99791: inst = 32'h24822800;
      99792: inst = 32'h10a00000;
      99793: inst = 32'hca00004;
      99794: inst = 32'h38632800;
      99795: inst = 32'h38842800;
      99796: inst = 32'h10a00001;
      99797: inst = 32'hca085d9;
      99798: inst = 32'h13e00001;
      99799: inst = 32'hfe0d96a;
      99800: inst = 32'h5be00000;
      99801: inst = 32'h8c50000;
      99802: inst = 32'h24612800;
      99803: inst = 32'h10a00000;
      99804: inst = 32'hca00010;
      99805: inst = 32'h24822800;
      99806: inst = 32'h10a00000;
      99807: inst = 32'hca00004;
      99808: inst = 32'h38632800;
      99809: inst = 32'h38842800;
      99810: inst = 32'h10a00001;
      99811: inst = 32'hca085e7;
      99812: inst = 32'h13e00001;
      99813: inst = 32'hfe0d96a;
      99814: inst = 32'h5be00000;
      99815: inst = 32'h8c50000;
      99816: inst = 32'h24612800;
      99817: inst = 32'h10a00000;
      99818: inst = 32'hca00010;
      99819: inst = 32'h24822800;
      99820: inst = 32'h10a00000;
      99821: inst = 32'hca00004;
      99822: inst = 32'h38632800;
      99823: inst = 32'h38842800;
      99824: inst = 32'h10a00001;
      99825: inst = 32'hca085f5;
      99826: inst = 32'h13e00001;
      99827: inst = 32'hfe0d96a;
      99828: inst = 32'h5be00000;
      99829: inst = 32'h8c50000;
      99830: inst = 32'h24612800;
      99831: inst = 32'h10a00000;
      99832: inst = 32'hca00010;
      99833: inst = 32'h24822800;
      99834: inst = 32'h10a00000;
      99835: inst = 32'hca00004;
      99836: inst = 32'h38632800;
      99837: inst = 32'h38842800;
      99838: inst = 32'h10a00001;
      99839: inst = 32'hca08603;
      99840: inst = 32'h13e00001;
      99841: inst = 32'hfe0d96a;
      99842: inst = 32'h5be00000;
      99843: inst = 32'h8c50000;
      99844: inst = 32'h24612800;
      99845: inst = 32'h10a00000;
      99846: inst = 32'hca00010;
      99847: inst = 32'h24822800;
      99848: inst = 32'h10a00000;
      99849: inst = 32'hca00004;
      99850: inst = 32'h38632800;
      99851: inst = 32'h38842800;
      99852: inst = 32'h10a00001;
      99853: inst = 32'hca08611;
      99854: inst = 32'h13e00001;
      99855: inst = 32'hfe0d96a;
      99856: inst = 32'h5be00000;
      99857: inst = 32'h8c50000;
      99858: inst = 32'h24612800;
      99859: inst = 32'h10a00000;
      99860: inst = 32'hca00010;
      99861: inst = 32'h24822800;
      99862: inst = 32'h10a00000;
      99863: inst = 32'hca00004;
      99864: inst = 32'h38632800;
      99865: inst = 32'h38842800;
      99866: inst = 32'h10a00001;
      99867: inst = 32'hca0861f;
      99868: inst = 32'h13e00001;
      99869: inst = 32'hfe0d96a;
      99870: inst = 32'h5be00000;
      99871: inst = 32'h8c50000;
      99872: inst = 32'h24612800;
      99873: inst = 32'h10a00000;
      99874: inst = 32'hca00010;
      99875: inst = 32'h24822800;
      99876: inst = 32'h10a00000;
      99877: inst = 32'hca00004;
      99878: inst = 32'h38632800;
      99879: inst = 32'h38842800;
      99880: inst = 32'h10a00001;
      99881: inst = 32'hca0862d;
      99882: inst = 32'h13e00001;
      99883: inst = 32'hfe0d96a;
      99884: inst = 32'h5be00000;
      99885: inst = 32'h8c50000;
      99886: inst = 32'h24612800;
      99887: inst = 32'h10a00000;
      99888: inst = 32'hca00010;
      99889: inst = 32'h24822800;
      99890: inst = 32'h10a00000;
      99891: inst = 32'hca00004;
      99892: inst = 32'h38632800;
      99893: inst = 32'h38842800;
      99894: inst = 32'h10a00001;
      99895: inst = 32'hca0863b;
      99896: inst = 32'h13e00001;
      99897: inst = 32'hfe0d96a;
      99898: inst = 32'h5be00000;
      99899: inst = 32'h8c50000;
      99900: inst = 32'h24612800;
      99901: inst = 32'h10a00000;
      99902: inst = 32'hca00010;
      99903: inst = 32'h24822800;
      99904: inst = 32'h10a00000;
      99905: inst = 32'hca00004;
      99906: inst = 32'h38632800;
      99907: inst = 32'h38842800;
      99908: inst = 32'h10a00001;
      99909: inst = 32'hca08649;
      99910: inst = 32'h13e00001;
      99911: inst = 32'hfe0d96a;
      99912: inst = 32'h5be00000;
      99913: inst = 32'h8c50000;
      99914: inst = 32'h24612800;
      99915: inst = 32'h10a00000;
      99916: inst = 32'hca00010;
      99917: inst = 32'h24822800;
      99918: inst = 32'h10a00000;
      99919: inst = 32'hca00004;
      99920: inst = 32'h38632800;
      99921: inst = 32'h38842800;
      99922: inst = 32'h10a00001;
      99923: inst = 32'hca08657;
      99924: inst = 32'h13e00001;
      99925: inst = 32'hfe0d96a;
      99926: inst = 32'h5be00000;
      99927: inst = 32'h8c50000;
      99928: inst = 32'h24612800;
      99929: inst = 32'h10a00000;
      99930: inst = 32'hca00010;
      99931: inst = 32'h24822800;
      99932: inst = 32'h10a00000;
      99933: inst = 32'hca00004;
      99934: inst = 32'h38632800;
      99935: inst = 32'h38842800;
      99936: inst = 32'h10a00001;
      99937: inst = 32'hca08665;
      99938: inst = 32'h13e00001;
      99939: inst = 32'hfe0d96a;
      99940: inst = 32'h5be00000;
      99941: inst = 32'h8c50000;
      99942: inst = 32'h24612800;
      99943: inst = 32'h10a00000;
      99944: inst = 32'hca00010;
      99945: inst = 32'h24822800;
      99946: inst = 32'h10a00000;
      99947: inst = 32'hca00004;
      99948: inst = 32'h38632800;
      99949: inst = 32'h38842800;
      99950: inst = 32'h10a00001;
      99951: inst = 32'hca08673;
      99952: inst = 32'h13e00001;
      99953: inst = 32'hfe0d96a;
      99954: inst = 32'h5be00000;
      99955: inst = 32'h8c50000;
      99956: inst = 32'h24612800;
      99957: inst = 32'h10a00000;
      99958: inst = 32'hca00010;
      99959: inst = 32'h24822800;
      99960: inst = 32'h10a00000;
      99961: inst = 32'hca00004;
      99962: inst = 32'h38632800;
      99963: inst = 32'h38842800;
      99964: inst = 32'h10a00001;
      99965: inst = 32'hca08681;
      99966: inst = 32'h13e00001;
      99967: inst = 32'hfe0d96a;
      99968: inst = 32'h5be00000;
      99969: inst = 32'h8c50000;
      99970: inst = 32'h24612800;
      99971: inst = 32'h10a00000;
      99972: inst = 32'hca00010;
      99973: inst = 32'h24822800;
      99974: inst = 32'h10a00000;
      99975: inst = 32'hca00004;
      99976: inst = 32'h38632800;
      99977: inst = 32'h38842800;
      99978: inst = 32'h10a00001;
      99979: inst = 32'hca0868f;
      99980: inst = 32'h13e00001;
      99981: inst = 32'hfe0d96a;
      99982: inst = 32'h5be00000;
      99983: inst = 32'h8c50000;
      99984: inst = 32'h24612800;
      99985: inst = 32'h10a00000;
      99986: inst = 32'hca00010;
      99987: inst = 32'h24822800;
      99988: inst = 32'h10a00000;
      99989: inst = 32'hca00004;
      99990: inst = 32'h38632800;
      99991: inst = 32'h38842800;
      99992: inst = 32'h10a00001;
      99993: inst = 32'hca0869d;
      99994: inst = 32'h13e00001;
      99995: inst = 32'hfe0d96a;
      99996: inst = 32'h5be00000;
      99997: inst = 32'h8c50000;
      99998: inst = 32'h24612800;
      99999: inst = 32'h10a00000;
      100000: inst = 32'hca00010;
      100001: inst = 32'h24822800;
      100002: inst = 32'h10a00000;
      100003: inst = 32'hca00004;
      100004: inst = 32'h38632800;
      100005: inst = 32'h38842800;
      100006: inst = 32'h10a00001;
      100007: inst = 32'hca086ab;
      100008: inst = 32'h13e00001;
      100009: inst = 32'hfe0d96a;
      100010: inst = 32'h5be00000;
      100011: inst = 32'h8c50000;
      100012: inst = 32'h24612800;
      100013: inst = 32'h10a00000;
      100014: inst = 32'hca00010;
      100015: inst = 32'h24822800;
      100016: inst = 32'h10a00000;
      100017: inst = 32'hca00004;
      100018: inst = 32'h38632800;
      100019: inst = 32'h38842800;
      100020: inst = 32'h10a00001;
      100021: inst = 32'hca086b9;
      100022: inst = 32'h13e00001;
      100023: inst = 32'hfe0d96a;
      100024: inst = 32'h5be00000;
      100025: inst = 32'h8c50000;
      100026: inst = 32'h24612800;
      100027: inst = 32'h10a00000;
      100028: inst = 32'hca00010;
      100029: inst = 32'h24822800;
      100030: inst = 32'h10a00000;
      100031: inst = 32'hca00004;
      100032: inst = 32'h38632800;
      100033: inst = 32'h38842800;
      100034: inst = 32'h10a00001;
      100035: inst = 32'hca086c7;
      100036: inst = 32'h13e00001;
      100037: inst = 32'hfe0d96a;
      100038: inst = 32'h5be00000;
      100039: inst = 32'h8c50000;
      100040: inst = 32'h24612800;
      100041: inst = 32'h10a00000;
      100042: inst = 32'hca00010;
      100043: inst = 32'h24822800;
      100044: inst = 32'h10a00000;
      100045: inst = 32'hca00004;
      100046: inst = 32'h38632800;
      100047: inst = 32'h38842800;
      100048: inst = 32'h10a00001;
      100049: inst = 32'hca086d5;
      100050: inst = 32'h13e00001;
      100051: inst = 32'hfe0d96a;
      100052: inst = 32'h5be00000;
      100053: inst = 32'h8c50000;
      100054: inst = 32'h24612800;
      100055: inst = 32'h10a00000;
      100056: inst = 32'hca00010;
      100057: inst = 32'h24822800;
      100058: inst = 32'h10a00000;
      100059: inst = 32'hca00004;
      100060: inst = 32'h38632800;
      100061: inst = 32'h38842800;
      100062: inst = 32'h10a00001;
      100063: inst = 32'hca086e3;
      100064: inst = 32'h13e00001;
      100065: inst = 32'hfe0d96a;
      100066: inst = 32'h5be00000;
      100067: inst = 32'h8c50000;
      100068: inst = 32'h24612800;
      100069: inst = 32'h10a00000;
      100070: inst = 32'hca00010;
      100071: inst = 32'h24822800;
      100072: inst = 32'h10a00000;
      100073: inst = 32'hca00004;
      100074: inst = 32'h38632800;
      100075: inst = 32'h38842800;
      100076: inst = 32'h10a00001;
      100077: inst = 32'hca086f1;
      100078: inst = 32'h13e00001;
      100079: inst = 32'hfe0d96a;
      100080: inst = 32'h5be00000;
      100081: inst = 32'h8c50000;
      100082: inst = 32'h24612800;
      100083: inst = 32'h10a00000;
      100084: inst = 32'hca00010;
      100085: inst = 32'h24822800;
      100086: inst = 32'h10a00000;
      100087: inst = 32'hca00004;
      100088: inst = 32'h38632800;
      100089: inst = 32'h38842800;
      100090: inst = 32'h10a00001;
      100091: inst = 32'hca086ff;
      100092: inst = 32'h13e00001;
      100093: inst = 32'hfe0d96a;
      100094: inst = 32'h5be00000;
      100095: inst = 32'h8c50000;
      100096: inst = 32'h24612800;
      100097: inst = 32'h10a00000;
      100098: inst = 32'hca00010;
      100099: inst = 32'h24822800;
      100100: inst = 32'h10a00000;
      100101: inst = 32'hca00004;
      100102: inst = 32'h38632800;
      100103: inst = 32'h38842800;
      100104: inst = 32'h10a00001;
      100105: inst = 32'hca0870d;
      100106: inst = 32'h13e00001;
      100107: inst = 32'hfe0d96a;
      100108: inst = 32'h5be00000;
      100109: inst = 32'h8c50000;
      100110: inst = 32'h24612800;
      100111: inst = 32'h10a00000;
      100112: inst = 32'hca00010;
      100113: inst = 32'h24822800;
      100114: inst = 32'h10a00000;
      100115: inst = 32'hca00004;
      100116: inst = 32'h38632800;
      100117: inst = 32'h38842800;
      100118: inst = 32'h10a00001;
      100119: inst = 32'hca0871b;
      100120: inst = 32'h13e00001;
      100121: inst = 32'hfe0d96a;
      100122: inst = 32'h5be00000;
      100123: inst = 32'h8c50000;
      100124: inst = 32'h24612800;
      100125: inst = 32'h10a00000;
      100126: inst = 32'hca00010;
      100127: inst = 32'h24822800;
      100128: inst = 32'h10a00000;
      100129: inst = 32'hca00004;
      100130: inst = 32'h38632800;
      100131: inst = 32'h38842800;
      100132: inst = 32'h10a00001;
      100133: inst = 32'hca08729;
      100134: inst = 32'h13e00001;
      100135: inst = 32'hfe0d96a;
      100136: inst = 32'h5be00000;
      100137: inst = 32'h8c50000;
      100138: inst = 32'h24612800;
      100139: inst = 32'h10a00000;
      100140: inst = 32'hca00010;
      100141: inst = 32'h24822800;
      100142: inst = 32'h10a00000;
      100143: inst = 32'hca00004;
      100144: inst = 32'h38632800;
      100145: inst = 32'h38842800;
      100146: inst = 32'h10a00001;
      100147: inst = 32'hca08737;
      100148: inst = 32'h13e00001;
      100149: inst = 32'hfe0d96a;
      100150: inst = 32'h5be00000;
      100151: inst = 32'h8c50000;
      100152: inst = 32'h24612800;
      100153: inst = 32'h10a00000;
      100154: inst = 32'hca00010;
      100155: inst = 32'h24822800;
      100156: inst = 32'h10a00000;
      100157: inst = 32'hca00004;
      100158: inst = 32'h38632800;
      100159: inst = 32'h38842800;
      100160: inst = 32'h10a00001;
      100161: inst = 32'hca08745;
      100162: inst = 32'h13e00001;
      100163: inst = 32'hfe0d96a;
      100164: inst = 32'h5be00000;
      100165: inst = 32'h8c50000;
      100166: inst = 32'h24612800;
      100167: inst = 32'h10a00000;
      100168: inst = 32'hca00010;
      100169: inst = 32'h24822800;
      100170: inst = 32'h10a00000;
      100171: inst = 32'hca00004;
      100172: inst = 32'h38632800;
      100173: inst = 32'h38842800;
      100174: inst = 32'h10a00001;
      100175: inst = 32'hca08753;
      100176: inst = 32'h13e00001;
      100177: inst = 32'hfe0d96a;
      100178: inst = 32'h5be00000;
      100179: inst = 32'h8c50000;
      100180: inst = 32'h24612800;
      100181: inst = 32'h10a00000;
      100182: inst = 32'hca00010;
      100183: inst = 32'h24822800;
      100184: inst = 32'h10a00000;
      100185: inst = 32'hca00004;
      100186: inst = 32'h38632800;
      100187: inst = 32'h38842800;
      100188: inst = 32'h10a00001;
      100189: inst = 32'hca08761;
      100190: inst = 32'h13e00001;
      100191: inst = 32'hfe0d96a;
      100192: inst = 32'h5be00000;
      100193: inst = 32'h8c50000;
      100194: inst = 32'h24612800;
      100195: inst = 32'h10a00000;
      100196: inst = 32'hca00010;
      100197: inst = 32'h24822800;
      100198: inst = 32'h10a00000;
      100199: inst = 32'hca00004;
      100200: inst = 32'h38632800;
      100201: inst = 32'h38842800;
      100202: inst = 32'h10a00001;
      100203: inst = 32'hca0876f;
      100204: inst = 32'h13e00001;
      100205: inst = 32'hfe0d96a;
      100206: inst = 32'h5be00000;
      100207: inst = 32'h8c50000;
      100208: inst = 32'h24612800;
      100209: inst = 32'h10a00000;
      100210: inst = 32'hca00010;
      100211: inst = 32'h24822800;
      100212: inst = 32'h10a00000;
      100213: inst = 32'hca00004;
      100214: inst = 32'h38632800;
      100215: inst = 32'h38842800;
      100216: inst = 32'h10a00001;
      100217: inst = 32'hca0877d;
      100218: inst = 32'h13e00001;
      100219: inst = 32'hfe0d96a;
      100220: inst = 32'h5be00000;
      100221: inst = 32'h8c50000;
      100222: inst = 32'h24612800;
      100223: inst = 32'h10a00000;
      100224: inst = 32'hca00010;
      100225: inst = 32'h24822800;
      100226: inst = 32'h10a00000;
      100227: inst = 32'hca00004;
      100228: inst = 32'h38632800;
      100229: inst = 32'h38842800;
      100230: inst = 32'h10a00001;
      100231: inst = 32'hca0878b;
      100232: inst = 32'h13e00001;
      100233: inst = 32'hfe0d96a;
      100234: inst = 32'h5be00000;
      100235: inst = 32'h8c50000;
      100236: inst = 32'h24612800;
      100237: inst = 32'h10a00000;
      100238: inst = 32'hca00010;
      100239: inst = 32'h24822800;
      100240: inst = 32'h10a00000;
      100241: inst = 32'hca00004;
      100242: inst = 32'h38632800;
      100243: inst = 32'h38842800;
      100244: inst = 32'h10a00001;
      100245: inst = 32'hca08799;
      100246: inst = 32'h13e00001;
      100247: inst = 32'hfe0d96a;
      100248: inst = 32'h5be00000;
      100249: inst = 32'h8c50000;
      100250: inst = 32'h24612800;
      100251: inst = 32'h10a00000;
      100252: inst = 32'hca00010;
      100253: inst = 32'h24822800;
      100254: inst = 32'h10a00000;
      100255: inst = 32'hca00004;
      100256: inst = 32'h38632800;
      100257: inst = 32'h38842800;
      100258: inst = 32'h10a00001;
      100259: inst = 32'hca087a7;
      100260: inst = 32'h13e00001;
      100261: inst = 32'hfe0d96a;
      100262: inst = 32'h5be00000;
      100263: inst = 32'h8c50000;
      100264: inst = 32'h24612800;
      100265: inst = 32'h10a00000;
      100266: inst = 32'hca00010;
      100267: inst = 32'h24822800;
      100268: inst = 32'h10a00000;
      100269: inst = 32'hca00004;
      100270: inst = 32'h38632800;
      100271: inst = 32'h38842800;
      100272: inst = 32'h10a00001;
      100273: inst = 32'hca087b5;
      100274: inst = 32'h13e00001;
      100275: inst = 32'hfe0d96a;
      100276: inst = 32'h5be00000;
      100277: inst = 32'h8c50000;
      100278: inst = 32'h24612800;
      100279: inst = 32'h10a00000;
      100280: inst = 32'hca00010;
      100281: inst = 32'h24822800;
      100282: inst = 32'h10a00000;
      100283: inst = 32'hca00004;
      100284: inst = 32'h38632800;
      100285: inst = 32'h38842800;
      100286: inst = 32'h10a00001;
      100287: inst = 32'hca087c3;
      100288: inst = 32'h13e00001;
      100289: inst = 32'hfe0d96a;
      100290: inst = 32'h5be00000;
      100291: inst = 32'h8c50000;
      100292: inst = 32'h24612800;
      100293: inst = 32'h10a00000;
      100294: inst = 32'hca00010;
      100295: inst = 32'h24822800;
      100296: inst = 32'h10a00000;
      100297: inst = 32'hca00004;
      100298: inst = 32'h38632800;
      100299: inst = 32'h38842800;
      100300: inst = 32'h10a00001;
      100301: inst = 32'hca087d1;
      100302: inst = 32'h13e00001;
      100303: inst = 32'hfe0d96a;
      100304: inst = 32'h5be00000;
      100305: inst = 32'h8c50000;
      100306: inst = 32'h24612800;
      100307: inst = 32'h10a00000;
      100308: inst = 32'hca00010;
      100309: inst = 32'h24822800;
      100310: inst = 32'h10a00000;
      100311: inst = 32'hca00004;
      100312: inst = 32'h38632800;
      100313: inst = 32'h38842800;
      100314: inst = 32'h10a00001;
      100315: inst = 32'hca087df;
      100316: inst = 32'h13e00001;
      100317: inst = 32'hfe0d96a;
      100318: inst = 32'h5be00000;
      100319: inst = 32'h8c50000;
      100320: inst = 32'h24612800;
      100321: inst = 32'h10a00000;
      100322: inst = 32'hca00010;
      100323: inst = 32'h24822800;
      100324: inst = 32'h10a00000;
      100325: inst = 32'hca00004;
      100326: inst = 32'h38632800;
      100327: inst = 32'h38842800;
      100328: inst = 32'h10a00001;
      100329: inst = 32'hca087ed;
      100330: inst = 32'h13e00001;
      100331: inst = 32'hfe0d96a;
      100332: inst = 32'h5be00000;
      100333: inst = 32'h8c50000;
      100334: inst = 32'h24612800;
      100335: inst = 32'h10a00000;
      100336: inst = 32'hca00010;
      100337: inst = 32'h24822800;
      100338: inst = 32'h10a00000;
      100339: inst = 32'hca00004;
      100340: inst = 32'h38632800;
      100341: inst = 32'h38842800;
      100342: inst = 32'h10a00001;
      100343: inst = 32'hca087fb;
      100344: inst = 32'h13e00001;
      100345: inst = 32'hfe0d96a;
      100346: inst = 32'h5be00000;
      100347: inst = 32'h8c50000;
      100348: inst = 32'h24612800;
      100349: inst = 32'h10a00000;
      100350: inst = 32'hca00010;
      100351: inst = 32'h24822800;
      100352: inst = 32'h10a00000;
      100353: inst = 32'hca00004;
      100354: inst = 32'h38632800;
      100355: inst = 32'h38842800;
      100356: inst = 32'h10a00001;
      100357: inst = 32'hca08809;
      100358: inst = 32'h13e00001;
      100359: inst = 32'hfe0d96a;
      100360: inst = 32'h5be00000;
      100361: inst = 32'h8c50000;
      100362: inst = 32'h24612800;
      100363: inst = 32'h10a00000;
      100364: inst = 32'hca00010;
      100365: inst = 32'h24822800;
      100366: inst = 32'h10a00000;
      100367: inst = 32'hca00004;
      100368: inst = 32'h38632800;
      100369: inst = 32'h38842800;
      100370: inst = 32'h10a00001;
      100371: inst = 32'hca08817;
      100372: inst = 32'h13e00001;
      100373: inst = 32'hfe0d96a;
      100374: inst = 32'h5be00000;
      100375: inst = 32'h8c50000;
      100376: inst = 32'h24612800;
      100377: inst = 32'h10a00000;
      100378: inst = 32'hca00010;
      100379: inst = 32'h24822800;
      100380: inst = 32'h10a00000;
      100381: inst = 32'hca00004;
      100382: inst = 32'h38632800;
      100383: inst = 32'h38842800;
      100384: inst = 32'h10a00001;
      100385: inst = 32'hca08825;
      100386: inst = 32'h13e00001;
      100387: inst = 32'hfe0d96a;
      100388: inst = 32'h5be00000;
      100389: inst = 32'h8c50000;
      100390: inst = 32'h24612800;
      100391: inst = 32'h10a00000;
      100392: inst = 32'hca00010;
      100393: inst = 32'h24822800;
      100394: inst = 32'h10a00000;
      100395: inst = 32'hca00004;
      100396: inst = 32'h38632800;
      100397: inst = 32'h38842800;
      100398: inst = 32'h10a00001;
      100399: inst = 32'hca08833;
      100400: inst = 32'h13e00001;
      100401: inst = 32'hfe0d96a;
      100402: inst = 32'h5be00000;
      100403: inst = 32'h8c50000;
      100404: inst = 32'h24612800;
      100405: inst = 32'h10a00000;
      100406: inst = 32'hca00010;
      100407: inst = 32'h24822800;
      100408: inst = 32'h10a00000;
      100409: inst = 32'hca00004;
      100410: inst = 32'h38632800;
      100411: inst = 32'h38842800;
      100412: inst = 32'h10a00001;
      100413: inst = 32'hca08841;
      100414: inst = 32'h13e00001;
      100415: inst = 32'hfe0d96a;
      100416: inst = 32'h5be00000;
      100417: inst = 32'h8c50000;
      100418: inst = 32'h24612800;
      100419: inst = 32'h10a00000;
      100420: inst = 32'hca00010;
      100421: inst = 32'h24822800;
      100422: inst = 32'h10a00000;
      100423: inst = 32'hca00004;
      100424: inst = 32'h38632800;
      100425: inst = 32'h38842800;
      100426: inst = 32'h10a00001;
      100427: inst = 32'hca0884f;
      100428: inst = 32'h13e00001;
      100429: inst = 32'hfe0d96a;
      100430: inst = 32'h5be00000;
      100431: inst = 32'h8c50000;
      100432: inst = 32'h24612800;
      100433: inst = 32'h10a00000;
      100434: inst = 32'hca00010;
      100435: inst = 32'h24822800;
      100436: inst = 32'h10a00000;
      100437: inst = 32'hca00004;
      100438: inst = 32'h38632800;
      100439: inst = 32'h38842800;
      100440: inst = 32'h10a00001;
      100441: inst = 32'hca0885d;
      100442: inst = 32'h13e00001;
      100443: inst = 32'hfe0d96a;
      100444: inst = 32'h5be00000;
      100445: inst = 32'h8c50000;
      100446: inst = 32'h24612800;
      100447: inst = 32'h10a00000;
      100448: inst = 32'hca00010;
      100449: inst = 32'h24822800;
      100450: inst = 32'h10a00000;
      100451: inst = 32'hca00004;
      100452: inst = 32'h38632800;
      100453: inst = 32'h38842800;
      100454: inst = 32'h10a00001;
      100455: inst = 32'hca0886b;
      100456: inst = 32'h13e00001;
      100457: inst = 32'hfe0d96a;
      100458: inst = 32'h5be00000;
      100459: inst = 32'h8c50000;
      100460: inst = 32'h24612800;
      100461: inst = 32'h10a00000;
      100462: inst = 32'hca00010;
      100463: inst = 32'h24822800;
      100464: inst = 32'h10a00000;
      100465: inst = 32'hca00004;
      100466: inst = 32'h38632800;
      100467: inst = 32'h38842800;
      100468: inst = 32'h10a00001;
      100469: inst = 32'hca08879;
      100470: inst = 32'h13e00001;
      100471: inst = 32'hfe0d96a;
      100472: inst = 32'h5be00000;
      100473: inst = 32'h8c50000;
      100474: inst = 32'h24612800;
      100475: inst = 32'h10a00000;
      100476: inst = 32'hca00010;
      100477: inst = 32'h24822800;
      100478: inst = 32'h10a00000;
      100479: inst = 32'hca00004;
      100480: inst = 32'h38632800;
      100481: inst = 32'h38842800;
      100482: inst = 32'h10a00001;
      100483: inst = 32'hca08887;
      100484: inst = 32'h13e00001;
      100485: inst = 32'hfe0d96a;
      100486: inst = 32'h5be00000;
      100487: inst = 32'h8c50000;
      100488: inst = 32'h24612800;
      100489: inst = 32'h10a00000;
      100490: inst = 32'hca00010;
      100491: inst = 32'h24822800;
      100492: inst = 32'h10a00000;
      100493: inst = 32'hca00004;
      100494: inst = 32'h38632800;
      100495: inst = 32'h38842800;
      100496: inst = 32'h10a00001;
      100497: inst = 32'hca08895;
      100498: inst = 32'h13e00001;
      100499: inst = 32'hfe0d96a;
      100500: inst = 32'h5be00000;
      100501: inst = 32'h8c50000;
      100502: inst = 32'h24612800;
      100503: inst = 32'h10a00000;
      100504: inst = 32'hca00010;
      100505: inst = 32'h24822800;
      100506: inst = 32'h10a00000;
      100507: inst = 32'hca00004;
      100508: inst = 32'h38632800;
      100509: inst = 32'h38842800;
      100510: inst = 32'h10a00001;
      100511: inst = 32'hca088a3;
      100512: inst = 32'h13e00001;
      100513: inst = 32'hfe0d96a;
      100514: inst = 32'h5be00000;
      100515: inst = 32'h8c50000;
      100516: inst = 32'h24612800;
      100517: inst = 32'h10a00000;
      100518: inst = 32'hca00010;
      100519: inst = 32'h24822800;
      100520: inst = 32'h10a00000;
      100521: inst = 32'hca00004;
      100522: inst = 32'h38632800;
      100523: inst = 32'h38842800;
      100524: inst = 32'h10a00001;
      100525: inst = 32'hca088b1;
      100526: inst = 32'h13e00001;
      100527: inst = 32'hfe0d96a;
      100528: inst = 32'h5be00000;
      100529: inst = 32'h8c50000;
      100530: inst = 32'h24612800;
      100531: inst = 32'h10a00000;
      100532: inst = 32'hca00010;
      100533: inst = 32'h24822800;
      100534: inst = 32'h10a00000;
      100535: inst = 32'hca00004;
      100536: inst = 32'h38632800;
      100537: inst = 32'h38842800;
      100538: inst = 32'h10a00001;
      100539: inst = 32'hca088bf;
      100540: inst = 32'h13e00001;
      100541: inst = 32'hfe0d96a;
      100542: inst = 32'h5be00000;
      100543: inst = 32'h8c50000;
      100544: inst = 32'h24612800;
      100545: inst = 32'h10a00000;
      100546: inst = 32'hca00010;
      100547: inst = 32'h24822800;
      100548: inst = 32'h10a00000;
      100549: inst = 32'hca00004;
      100550: inst = 32'h38632800;
      100551: inst = 32'h38842800;
      100552: inst = 32'h10a00001;
      100553: inst = 32'hca088cd;
      100554: inst = 32'h13e00001;
      100555: inst = 32'hfe0d96a;
      100556: inst = 32'h5be00000;
      100557: inst = 32'h8c50000;
      100558: inst = 32'h24612800;
      100559: inst = 32'h10a00000;
      100560: inst = 32'hca00010;
      100561: inst = 32'h24822800;
      100562: inst = 32'h10a00000;
      100563: inst = 32'hca00004;
      100564: inst = 32'h38632800;
      100565: inst = 32'h38842800;
      100566: inst = 32'h10a00001;
      100567: inst = 32'hca088db;
      100568: inst = 32'h13e00001;
      100569: inst = 32'hfe0d96a;
      100570: inst = 32'h5be00000;
      100571: inst = 32'h8c50000;
      100572: inst = 32'h24612800;
      100573: inst = 32'h10a00000;
      100574: inst = 32'hca00010;
      100575: inst = 32'h24822800;
      100576: inst = 32'h10a00000;
      100577: inst = 32'hca00004;
      100578: inst = 32'h38632800;
      100579: inst = 32'h38842800;
      100580: inst = 32'h10a00001;
      100581: inst = 32'hca088e9;
      100582: inst = 32'h13e00001;
      100583: inst = 32'hfe0d96a;
      100584: inst = 32'h5be00000;
      100585: inst = 32'h8c50000;
      100586: inst = 32'h24612800;
      100587: inst = 32'h10a00000;
      100588: inst = 32'hca00010;
      100589: inst = 32'h24822800;
      100590: inst = 32'h10a00000;
      100591: inst = 32'hca00004;
      100592: inst = 32'h38632800;
      100593: inst = 32'h38842800;
      100594: inst = 32'h10a00001;
      100595: inst = 32'hca088f7;
      100596: inst = 32'h13e00001;
      100597: inst = 32'hfe0d96a;
      100598: inst = 32'h5be00000;
      100599: inst = 32'h8c50000;
      100600: inst = 32'h24612800;
      100601: inst = 32'h10a00000;
      100602: inst = 32'hca00010;
      100603: inst = 32'h24822800;
      100604: inst = 32'h10a00000;
      100605: inst = 32'hca00004;
      100606: inst = 32'h38632800;
      100607: inst = 32'h38842800;
      100608: inst = 32'h10a00001;
      100609: inst = 32'hca08905;
      100610: inst = 32'h13e00001;
      100611: inst = 32'hfe0d96a;
      100612: inst = 32'h5be00000;
      100613: inst = 32'h8c50000;
      100614: inst = 32'h24612800;
      100615: inst = 32'h10a00000;
      100616: inst = 32'hca00010;
      100617: inst = 32'h24822800;
      100618: inst = 32'h10a00000;
      100619: inst = 32'hca00004;
      100620: inst = 32'h38632800;
      100621: inst = 32'h38842800;
      100622: inst = 32'h10a00001;
      100623: inst = 32'hca08913;
      100624: inst = 32'h13e00001;
      100625: inst = 32'hfe0d96a;
      100626: inst = 32'h5be00000;
      100627: inst = 32'h8c50000;
      100628: inst = 32'h24612800;
      100629: inst = 32'h10a00000;
      100630: inst = 32'hca00010;
      100631: inst = 32'h24822800;
      100632: inst = 32'h10a00000;
      100633: inst = 32'hca00004;
      100634: inst = 32'h38632800;
      100635: inst = 32'h38842800;
      100636: inst = 32'h10a00001;
      100637: inst = 32'hca08921;
      100638: inst = 32'h13e00001;
      100639: inst = 32'hfe0d96a;
      100640: inst = 32'h5be00000;
      100641: inst = 32'h8c50000;
      100642: inst = 32'h24612800;
      100643: inst = 32'h10a00000;
      100644: inst = 32'hca00010;
      100645: inst = 32'h24822800;
      100646: inst = 32'h10a00000;
      100647: inst = 32'hca00004;
      100648: inst = 32'h38632800;
      100649: inst = 32'h38842800;
      100650: inst = 32'h10a00001;
      100651: inst = 32'hca0892f;
      100652: inst = 32'h13e00001;
      100653: inst = 32'hfe0d96a;
      100654: inst = 32'h5be00000;
      100655: inst = 32'h8c50000;
      100656: inst = 32'h24612800;
      100657: inst = 32'h10a00000;
      100658: inst = 32'hca00010;
      100659: inst = 32'h24822800;
      100660: inst = 32'h10a00000;
      100661: inst = 32'hca00004;
      100662: inst = 32'h38632800;
      100663: inst = 32'h38842800;
      100664: inst = 32'h10a00001;
      100665: inst = 32'hca0893d;
      100666: inst = 32'h13e00001;
      100667: inst = 32'hfe0d96a;
      100668: inst = 32'h5be00000;
      100669: inst = 32'h8c50000;
      100670: inst = 32'h24612800;
      100671: inst = 32'h10a00000;
      100672: inst = 32'hca00010;
      100673: inst = 32'h24822800;
      100674: inst = 32'h10a00000;
      100675: inst = 32'hca00004;
      100676: inst = 32'h38632800;
      100677: inst = 32'h38842800;
      100678: inst = 32'h10a00001;
      100679: inst = 32'hca0894b;
      100680: inst = 32'h13e00001;
      100681: inst = 32'hfe0d96a;
      100682: inst = 32'h5be00000;
      100683: inst = 32'h8c50000;
      100684: inst = 32'h24612800;
      100685: inst = 32'h10a00000;
      100686: inst = 32'hca00010;
      100687: inst = 32'h24822800;
      100688: inst = 32'h10a00000;
      100689: inst = 32'hca00004;
      100690: inst = 32'h38632800;
      100691: inst = 32'h38842800;
      100692: inst = 32'h10a00001;
      100693: inst = 32'hca08959;
      100694: inst = 32'h13e00001;
      100695: inst = 32'hfe0d96a;
      100696: inst = 32'h5be00000;
      100697: inst = 32'h8c50000;
      100698: inst = 32'h24612800;
      100699: inst = 32'h10a00000;
      100700: inst = 32'hca00010;
      100701: inst = 32'h24822800;
      100702: inst = 32'h10a00000;
      100703: inst = 32'hca00004;
      100704: inst = 32'h38632800;
      100705: inst = 32'h38842800;
      100706: inst = 32'h10a00001;
      100707: inst = 32'hca08967;
      100708: inst = 32'h13e00001;
      100709: inst = 32'hfe0d96a;
      100710: inst = 32'h5be00000;
      100711: inst = 32'h8c50000;
      100712: inst = 32'h24612800;
      100713: inst = 32'h10a00000;
      100714: inst = 32'hca00010;
      100715: inst = 32'h24822800;
      100716: inst = 32'h10a00000;
      100717: inst = 32'hca00004;
      100718: inst = 32'h38632800;
      100719: inst = 32'h38842800;
      100720: inst = 32'h10a00001;
      100721: inst = 32'hca08975;
      100722: inst = 32'h13e00001;
      100723: inst = 32'hfe0d96a;
      100724: inst = 32'h5be00000;
      100725: inst = 32'h8c50000;
      100726: inst = 32'h24612800;
      100727: inst = 32'h10a00000;
      100728: inst = 32'hca00010;
      100729: inst = 32'h24822800;
      100730: inst = 32'h10a00000;
      100731: inst = 32'hca00004;
      100732: inst = 32'h38632800;
      100733: inst = 32'h38842800;
      100734: inst = 32'h10a00001;
      100735: inst = 32'hca08983;
      100736: inst = 32'h13e00001;
      100737: inst = 32'hfe0d96a;
      100738: inst = 32'h5be00000;
      100739: inst = 32'h8c50000;
      100740: inst = 32'h24612800;
      100741: inst = 32'h10a00000;
      100742: inst = 32'hca00010;
      100743: inst = 32'h24822800;
      100744: inst = 32'h10a00000;
      100745: inst = 32'hca00004;
      100746: inst = 32'h38632800;
      100747: inst = 32'h38842800;
      100748: inst = 32'h10a00001;
      100749: inst = 32'hca08991;
      100750: inst = 32'h13e00001;
      100751: inst = 32'hfe0d96a;
      100752: inst = 32'h5be00000;
      100753: inst = 32'h8c50000;
      100754: inst = 32'h24612800;
      100755: inst = 32'h10a00000;
      100756: inst = 32'hca00010;
      100757: inst = 32'h24822800;
      100758: inst = 32'h10a00000;
      100759: inst = 32'hca00004;
      100760: inst = 32'h38632800;
      100761: inst = 32'h38842800;
      100762: inst = 32'h10a00001;
      100763: inst = 32'hca0899f;
      100764: inst = 32'h13e00001;
      100765: inst = 32'hfe0d96a;
      100766: inst = 32'h5be00000;
      100767: inst = 32'h8c50000;
      100768: inst = 32'h24612800;
      100769: inst = 32'h10a00000;
      100770: inst = 32'hca00010;
      100771: inst = 32'h24822800;
      100772: inst = 32'h10a00000;
      100773: inst = 32'hca00004;
      100774: inst = 32'h38632800;
      100775: inst = 32'h38842800;
      100776: inst = 32'h10a00001;
      100777: inst = 32'hca089ad;
      100778: inst = 32'h13e00001;
      100779: inst = 32'hfe0d96a;
      100780: inst = 32'h5be00000;
      100781: inst = 32'h8c50000;
      100782: inst = 32'h24612800;
      100783: inst = 32'h10a00000;
      100784: inst = 32'hca00010;
      100785: inst = 32'h24822800;
      100786: inst = 32'h10a00000;
      100787: inst = 32'hca00004;
      100788: inst = 32'h38632800;
      100789: inst = 32'h38842800;
      100790: inst = 32'h10a00001;
      100791: inst = 32'hca089bb;
      100792: inst = 32'h13e00001;
      100793: inst = 32'hfe0d96a;
      100794: inst = 32'h5be00000;
      100795: inst = 32'h8c50000;
      100796: inst = 32'h24612800;
      100797: inst = 32'h10a00000;
      100798: inst = 32'hca00010;
      100799: inst = 32'h24822800;
      100800: inst = 32'h10a00000;
      100801: inst = 32'hca00004;
      100802: inst = 32'h38632800;
      100803: inst = 32'h38842800;
      100804: inst = 32'h10a00001;
      100805: inst = 32'hca089c9;
      100806: inst = 32'h13e00001;
      100807: inst = 32'hfe0d96a;
      100808: inst = 32'h5be00000;
      100809: inst = 32'h8c50000;
      100810: inst = 32'h24612800;
      100811: inst = 32'h10a00000;
      100812: inst = 32'hca00010;
      100813: inst = 32'h24822800;
      100814: inst = 32'h10a00000;
      100815: inst = 32'hca00004;
      100816: inst = 32'h38632800;
      100817: inst = 32'h38842800;
      100818: inst = 32'h10a00001;
      100819: inst = 32'hca089d7;
      100820: inst = 32'h13e00001;
      100821: inst = 32'hfe0d96a;
      100822: inst = 32'h5be00000;
      100823: inst = 32'h8c50000;
      100824: inst = 32'h24612800;
      100825: inst = 32'h10a00000;
      100826: inst = 32'hca00010;
      100827: inst = 32'h24822800;
      100828: inst = 32'h10a00000;
      100829: inst = 32'hca00004;
      100830: inst = 32'h38632800;
      100831: inst = 32'h38842800;
      100832: inst = 32'h10a00001;
      100833: inst = 32'hca089e5;
      100834: inst = 32'h13e00001;
      100835: inst = 32'hfe0d96a;
      100836: inst = 32'h5be00000;
      100837: inst = 32'h8c50000;
      100838: inst = 32'h24612800;
      100839: inst = 32'h10a00000;
      100840: inst = 32'hca00010;
      100841: inst = 32'h24822800;
      100842: inst = 32'h10a00000;
      100843: inst = 32'hca00004;
      100844: inst = 32'h38632800;
      100845: inst = 32'h38842800;
      100846: inst = 32'h10a00001;
      100847: inst = 32'hca089f3;
      100848: inst = 32'h13e00001;
      100849: inst = 32'hfe0d96a;
      100850: inst = 32'h5be00000;
      100851: inst = 32'h8c50000;
      100852: inst = 32'h24612800;
      100853: inst = 32'h10a00000;
      100854: inst = 32'hca00010;
      100855: inst = 32'h24822800;
      100856: inst = 32'h10a00000;
      100857: inst = 32'hca00004;
      100858: inst = 32'h38632800;
      100859: inst = 32'h38842800;
      100860: inst = 32'h10a00001;
      100861: inst = 32'hca08a01;
      100862: inst = 32'h13e00001;
      100863: inst = 32'hfe0d96a;
      100864: inst = 32'h5be00000;
      100865: inst = 32'h8c50000;
      100866: inst = 32'h24612800;
      100867: inst = 32'h10a00000;
      100868: inst = 32'hca00010;
      100869: inst = 32'h24822800;
      100870: inst = 32'h10a00000;
      100871: inst = 32'hca00004;
      100872: inst = 32'h38632800;
      100873: inst = 32'h38842800;
      100874: inst = 32'h10a00001;
      100875: inst = 32'hca08a0f;
      100876: inst = 32'h13e00001;
      100877: inst = 32'hfe0d96a;
      100878: inst = 32'h5be00000;
      100879: inst = 32'h8c50000;
      100880: inst = 32'h24612800;
      100881: inst = 32'h10a00000;
      100882: inst = 32'hca00010;
      100883: inst = 32'h24822800;
      100884: inst = 32'h10a00000;
      100885: inst = 32'hca00004;
      100886: inst = 32'h38632800;
      100887: inst = 32'h38842800;
      100888: inst = 32'h10a00001;
      100889: inst = 32'hca08a1d;
      100890: inst = 32'h13e00001;
      100891: inst = 32'hfe0d96a;
      100892: inst = 32'h5be00000;
      100893: inst = 32'h8c50000;
      100894: inst = 32'h24612800;
      100895: inst = 32'h10a00000;
      100896: inst = 32'hca00010;
      100897: inst = 32'h24822800;
      100898: inst = 32'h10a00000;
      100899: inst = 32'hca00004;
      100900: inst = 32'h38632800;
      100901: inst = 32'h38842800;
      100902: inst = 32'h10a00001;
      100903: inst = 32'hca08a2b;
      100904: inst = 32'h13e00001;
      100905: inst = 32'hfe0d96a;
      100906: inst = 32'h5be00000;
      100907: inst = 32'h8c50000;
      100908: inst = 32'h24612800;
      100909: inst = 32'h10a00000;
      100910: inst = 32'hca00010;
      100911: inst = 32'h24822800;
      100912: inst = 32'h10a00000;
      100913: inst = 32'hca00004;
      100914: inst = 32'h38632800;
      100915: inst = 32'h38842800;
      100916: inst = 32'h10a00001;
      100917: inst = 32'hca08a39;
      100918: inst = 32'h13e00001;
      100919: inst = 32'hfe0d96a;
      100920: inst = 32'h5be00000;
      100921: inst = 32'h8c50000;
      100922: inst = 32'h24612800;
      100923: inst = 32'h10a00000;
      100924: inst = 32'hca00010;
      100925: inst = 32'h24822800;
      100926: inst = 32'h10a00000;
      100927: inst = 32'hca00004;
      100928: inst = 32'h38632800;
      100929: inst = 32'h38842800;
      100930: inst = 32'h10a00001;
      100931: inst = 32'hca08a47;
      100932: inst = 32'h13e00001;
      100933: inst = 32'hfe0d96a;
      100934: inst = 32'h5be00000;
      100935: inst = 32'h8c50000;
      100936: inst = 32'h24612800;
      100937: inst = 32'h10a00000;
      100938: inst = 32'hca00010;
      100939: inst = 32'h24822800;
      100940: inst = 32'h10a00000;
      100941: inst = 32'hca00004;
      100942: inst = 32'h38632800;
      100943: inst = 32'h38842800;
      100944: inst = 32'h10a00001;
      100945: inst = 32'hca08a55;
      100946: inst = 32'h13e00001;
      100947: inst = 32'hfe0d96a;
      100948: inst = 32'h5be00000;
      100949: inst = 32'h8c50000;
      100950: inst = 32'h24612800;
      100951: inst = 32'h10a00000;
      100952: inst = 32'hca00010;
      100953: inst = 32'h24822800;
      100954: inst = 32'h10a00000;
      100955: inst = 32'hca00004;
      100956: inst = 32'h38632800;
      100957: inst = 32'h38842800;
      100958: inst = 32'h10a00001;
      100959: inst = 32'hca08a63;
      100960: inst = 32'h13e00001;
      100961: inst = 32'hfe0d96a;
      100962: inst = 32'h5be00000;
      100963: inst = 32'h8c50000;
      100964: inst = 32'h24612800;
      100965: inst = 32'h10a00000;
      100966: inst = 32'hca00010;
      100967: inst = 32'h24822800;
      100968: inst = 32'h10a00000;
      100969: inst = 32'hca00004;
      100970: inst = 32'h38632800;
      100971: inst = 32'h38842800;
      100972: inst = 32'h10a00001;
      100973: inst = 32'hca08a71;
      100974: inst = 32'h13e00001;
      100975: inst = 32'hfe0d96a;
      100976: inst = 32'h5be00000;
      100977: inst = 32'h8c50000;
      100978: inst = 32'h24612800;
      100979: inst = 32'h10a00000;
      100980: inst = 32'hca00010;
      100981: inst = 32'h24822800;
      100982: inst = 32'h10a00000;
      100983: inst = 32'hca00004;
      100984: inst = 32'h38632800;
      100985: inst = 32'h38842800;
      100986: inst = 32'h10a00001;
      100987: inst = 32'hca08a7f;
      100988: inst = 32'h13e00001;
      100989: inst = 32'hfe0d96a;
      100990: inst = 32'h5be00000;
      100991: inst = 32'h8c50000;
      100992: inst = 32'h24612800;
      100993: inst = 32'h10a00000;
      100994: inst = 32'hca00010;
      100995: inst = 32'h24822800;
      100996: inst = 32'h10a00000;
      100997: inst = 32'hca00004;
      100998: inst = 32'h38632800;
      100999: inst = 32'h38842800;
      101000: inst = 32'h10a00001;
      101001: inst = 32'hca08a8d;
      101002: inst = 32'h13e00001;
      101003: inst = 32'hfe0d96a;
      101004: inst = 32'h5be00000;
      101005: inst = 32'h8c50000;
      101006: inst = 32'h24612800;
      101007: inst = 32'h10a00000;
      101008: inst = 32'hca00010;
      101009: inst = 32'h24822800;
      101010: inst = 32'h10a00000;
      101011: inst = 32'hca00004;
      101012: inst = 32'h38632800;
      101013: inst = 32'h38842800;
      101014: inst = 32'h10a00001;
      101015: inst = 32'hca08a9b;
      101016: inst = 32'h13e00001;
      101017: inst = 32'hfe0d96a;
      101018: inst = 32'h5be00000;
      101019: inst = 32'h8c50000;
      101020: inst = 32'h24612800;
      101021: inst = 32'h10a00000;
      101022: inst = 32'hca00010;
      101023: inst = 32'h24822800;
      101024: inst = 32'h10a00000;
      101025: inst = 32'hca00004;
      101026: inst = 32'h38632800;
      101027: inst = 32'h38842800;
      101028: inst = 32'h10a00001;
      101029: inst = 32'hca08aa9;
      101030: inst = 32'h13e00001;
      101031: inst = 32'hfe0d96a;
      101032: inst = 32'h5be00000;
      101033: inst = 32'h8c50000;
      101034: inst = 32'h24612800;
      101035: inst = 32'h10a00000;
      101036: inst = 32'hca00011;
      101037: inst = 32'h24822800;
      101038: inst = 32'h10a00000;
      101039: inst = 32'hca00004;
      101040: inst = 32'h38632800;
      101041: inst = 32'h38842800;
      101042: inst = 32'h10a00001;
      101043: inst = 32'hca08ab7;
      101044: inst = 32'h13e00001;
      101045: inst = 32'hfe0d96a;
      101046: inst = 32'h5be00000;
      101047: inst = 32'h8c50000;
      101048: inst = 32'h24612800;
      101049: inst = 32'h10a00000;
      101050: inst = 32'hca00011;
      101051: inst = 32'h24822800;
      101052: inst = 32'h10a00000;
      101053: inst = 32'hca00004;
      101054: inst = 32'h38632800;
      101055: inst = 32'h38842800;
      101056: inst = 32'h10a00001;
      101057: inst = 32'hca08ac5;
      101058: inst = 32'h13e00001;
      101059: inst = 32'hfe0d96a;
      101060: inst = 32'h5be00000;
      101061: inst = 32'h8c50000;
      101062: inst = 32'h24612800;
      101063: inst = 32'h10a00000;
      101064: inst = 32'hca00011;
      101065: inst = 32'h24822800;
      101066: inst = 32'h10a00000;
      101067: inst = 32'hca00004;
      101068: inst = 32'h38632800;
      101069: inst = 32'h38842800;
      101070: inst = 32'h10a00001;
      101071: inst = 32'hca08ad3;
      101072: inst = 32'h13e00001;
      101073: inst = 32'hfe0d96a;
      101074: inst = 32'h5be00000;
      101075: inst = 32'h8c50000;
      101076: inst = 32'h24612800;
      101077: inst = 32'h10a00000;
      101078: inst = 32'hca00011;
      101079: inst = 32'h24822800;
      101080: inst = 32'h10a00000;
      101081: inst = 32'hca00004;
      101082: inst = 32'h38632800;
      101083: inst = 32'h38842800;
      101084: inst = 32'h10a00001;
      101085: inst = 32'hca08ae1;
      101086: inst = 32'h13e00001;
      101087: inst = 32'hfe0d96a;
      101088: inst = 32'h5be00000;
      101089: inst = 32'h8c50000;
      101090: inst = 32'h24612800;
      101091: inst = 32'h10a00000;
      101092: inst = 32'hca00011;
      101093: inst = 32'h24822800;
      101094: inst = 32'h10a00000;
      101095: inst = 32'hca00004;
      101096: inst = 32'h38632800;
      101097: inst = 32'h38842800;
      101098: inst = 32'h10a00001;
      101099: inst = 32'hca08aef;
      101100: inst = 32'h13e00001;
      101101: inst = 32'hfe0d96a;
      101102: inst = 32'h5be00000;
      101103: inst = 32'h8c50000;
      101104: inst = 32'h24612800;
      101105: inst = 32'h10a00000;
      101106: inst = 32'hca00011;
      101107: inst = 32'h24822800;
      101108: inst = 32'h10a00000;
      101109: inst = 32'hca00004;
      101110: inst = 32'h38632800;
      101111: inst = 32'h38842800;
      101112: inst = 32'h10a00001;
      101113: inst = 32'hca08afd;
      101114: inst = 32'h13e00001;
      101115: inst = 32'hfe0d96a;
      101116: inst = 32'h5be00000;
      101117: inst = 32'h8c50000;
      101118: inst = 32'h24612800;
      101119: inst = 32'h10a00000;
      101120: inst = 32'hca00011;
      101121: inst = 32'h24822800;
      101122: inst = 32'h10a00000;
      101123: inst = 32'hca00004;
      101124: inst = 32'h38632800;
      101125: inst = 32'h38842800;
      101126: inst = 32'h10a00001;
      101127: inst = 32'hca08b0b;
      101128: inst = 32'h13e00001;
      101129: inst = 32'hfe0d96a;
      101130: inst = 32'h5be00000;
      101131: inst = 32'h8c50000;
      101132: inst = 32'h24612800;
      101133: inst = 32'h10a00000;
      101134: inst = 32'hca00011;
      101135: inst = 32'h24822800;
      101136: inst = 32'h10a00000;
      101137: inst = 32'hca00004;
      101138: inst = 32'h38632800;
      101139: inst = 32'h38842800;
      101140: inst = 32'h10a00001;
      101141: inst = 32'hca08b19;
      101142: inst = 32'h13e00001;
      101143: inst = 32'hfe0d96a;
      101144: inst = 32'h5be00000;
      101145: inst = 32'h8c50000;
      101146: inst = 32'h24612800;
      101147: inst = 32'h10a00000;
      101148: inst = 32'hca00011;
      101149: inst = 32'h24822800;
      101150: inst = 32'h10a00000;
      101151: inst = 32'hca00004;
      101152: inst = 32'h38632800;
      101153: inst = 32'h38842800;
      101154: inst = 32'h10a00001;
      101155: inst = 32'hca08b27;
      101156: inst = 32'h13e00001;
      101157: inst = 32'hfe0d96a;
      101158: inst = 32'h5be00000;
      101159: inst = 32'h8c50000;
      101160: inst = 32'h24612800;
      101161: inst = 32'h10a00000;
      101162: inst = 32'hca00011;
      101163: inst = 32'h24822800;
      101164: inst = 32'h10a00000;
      101165: inst = 32'hca00004;
      101166: inst = 32'h38632800;
      101167: inst = 32'h38842800;
      101168: inst = 32'h10a00001;
      101169: inst = 32'hca08b35;
      101170: inst = 32'h13e00001;
      101171: inst = 32'hfe0d96a;
      101172: inst = 32'h5be00000;
      101173: inst = 32'h8c50000;
      101174: inst = 32'h24612800;
      101175: inst = 32'h10a00000;
      101176: inst = 32'hca00011;
      101177: inst = 32'h24822800;
      101178: inst = 32'h10a00000;
      101179: inst = 32'hca00004;
      101180: inst = 32'h38632800;
      101181: inst = 32'h38842800;
      101182: inst = 32'h10a00001;
      101183: inst = 32'hca08b43;
      101184: inst = 32'h13e00001;
      101185: inst = 32'hfe0d96a;
      101186: inst = 32'h5be00000;
      101187: inst = 32'h8c50000;
      101188: inst = 32'h24612800;
      101189: inst = 32'h10a00000;
      101190: inst = 32'hca00011;
      101191: inst = 32'h24822800;
      101192: inst = 32'h10a00000;
      101193: inst = 32'hca00004;
      101194: inst = 32'h38632800;
      101195: inst = 32'h38842800;
      101196: inst = 32'h10a00001;
      101197: inst = 32'hca08b51;
      101198: inst = 32'h13e00001;
      101199: inst = 32'hfe0d96a;
      101200: inst = 32'h5be00000;
      101201: inst = 32'h8c50000;
      101202: inst = 32'h24612800;
      101203: inst = 32'h10a00000;
      101204: inst = 32'hca00011;
      101205: inst = 32'h24822800;
      101206: inst = 32'h10a00000;
      101207: inst = 32'hca00004;
      101208: inst = 32'h38632800;
      101209: inst = 32'h38842800;
      101210: inst = 32'h10a00001;
      101211: inst = 32'hca08b5f;
      101212: inst = 32'h13e00001;
      101213: inst = 32'hfe0d96a;
      101214: inst = 32'h5be00000;
      101215: inst = 32'h8c50000;
      101216: inst = 32'h24612800;
      101217: inst = 32'h10a00000;
      101218: inst = 32'hca00011;
      101219: inst = 32'h24822800;
      101220: inst = 32'h10a00000;
      101221: inst = 32'hca00004;
      101222: inst = 32'h38632800;
      101223: inst = 32'h38842800;
      101224: inst = 32'h10a00001;
      101225: inst = 32'hca08b6d;
      101226: inst = 32'h13e00001;
      101227: inst = 32'hfe0d96a;
      101228: inst = 32'h5be00000;
      101229: inst = 32'h8c50000;
      101230: inst = 32'h24612800;
      101231: inst = 32'h10a00000;
      101232: inst = 32'hca00011;
      101233: inst = 32'h24822800;
      101234: inst = 32'h10a00000;
      101235: inst = 32'hca00004;
      101236: inst = 32'h38632800;
      101237: inst = 32'h38842800;
      101238: inst = 32'h10a00001;
      101239: inst = 32'hca08b7b;
      101240: inst = 32'h13e00001;
      101241: inst = 32'hfe0d96a;
      101242: inst = 32'h5be00000;
      101243: inst = 32'h8c50000;
      101244: inst = 32'h24612800;
      101245: inst = 32'h10a00000;
      101246: inst = 32'hca00011;
      101247: inst = 32'h24822800;
      101248: inst = 32'h10a00000;
      101249: inst = 32'hca00004;
      101250: inst = 32'h38632800;
      101251: inst = 32'h38842800;
      101252: inst = 32'h10a00001;
      101253: inst = 32'hca08b89;
      101254: inst = 32'h13e00001;
      101255: inst = 32'hfe0d96a;
      101256: inst = 32'h5be00000;
      101257: inst = 32'h8c50000;
      101258: inst = 32'h24612800;
      101259: inst = 32'h10a00000;
      101260: inst = 32'hca00011;
      101261: inst = 32'h24822800;
      101262: inst = 32'h10a00000;
      101263: inst = 32'hca00004;
      101264: inst = 32'h38632800;
      101265: inst = 32'h38842800;
      101266: inst = 32'h10a00001;
      101267: inst = 32'hca08b97;
      101268: inst = 32'h13e00001;
      101269: inst = 32'hfe0d96a;
      101270: inst = 32'h5be00000;
      101271: inst = 32'h8c50000;
      101272: inst = 32'h24612800;
      101273: inst = 32'h10a00000;
      101274: inst = 32'hca00011;
      101275: inst = 32'h24822800;
      101276: inst = 32'h10a00000;
      101277: inst = 32'hca00004;
      101278: inst = 32'h38632800;
      101279: inst = 32'h38842800;
      101280: inst = 32'h10a00001;
      101281: inst = 32'hca08ba5;
      101282: inst = 32'h13e00001;
      101283: inst = 32'hfe0d96a;
      101284: inst = 32'h5be00000;
      101285: inst = 32'h8c50000;
      101286: inst = 32'h24612800;
      101287: inst = 32'h10a00000;
      101288: inst = 32'hca00011;
      101289: inst = 32'h24822800;
      101290: inst = 32'h10a00000;
      101291: inst = 32'hca00004;
      101292: inst = 32'h38632800;
      101293: inst = 32'h38842800;
      101294: inst = 32'h10a00001;
      101295: inst = 32'hca08bb3;
      101296: inst = 32'h13e00001;
      101297: inst = 32'hfe0d96a;
      101298: inst = 32'h5be00000;
      101299: inst = 32'h8c50000;
      101300: inst = 32'h24612800;
      101301: inst = 32'h10a00000;
      101302: inst = 32'hca00011;
      101303: inst = 32'h24822800;
      101304: inst = 32'h10a00000;
      101305: inst = 32'hca00004;
      101306: inst = 32'h38632800;
      101307: inst = 32'h38842800;
      101308: inst = 32'h10a00001;
      101309: inst = 32'hca08bc1;
      101310: inst = 32'h13e00001;
      101311: inst = 32'hfe0d96a;
      101312: inst = 32'h5be00000;
      101313: inst = 32'h8c50000;
      101314: inst = 32'h24612800;
      101315: inst = 32'h10a00000;
      101316: inst = 32'hca00011;
      101317: inst = 32'h24822800;
      101318: inst = 32'h10a00000;
      101319: inst = 32'hca00004;
      101320: inst = 32'h38632800;
      101321: inst = 32'h38842800;
      101322: inst = 32'h10a00001;
      101323: inst = 32'hca08bcf;
      101324: inst = 32'h13e00001;
      101325: inst = 32'hfe0d96a;
      101326: inst = 32'h5be00000;
      101327: inst = 32'h8c50000;
      101328: inst = 32'h24612800;
      101329: inst = 32'h10a00000;
      101330: inst = 32'hca00011;
      101331: inst = 32'h24822800;
      101332: inst = 32'h10a00000;
      101333: inst = 32'hca00004;
      101334: inst = 32'h38632800;
      101335: inst = 32'h38842800;
      101336: inst = 32'h10a00001;
      101337: inst = 32'hca08bdd;
      101338: inst = 32'h13e00001;
      101339: inst = 32'hfe0d96a;
      101340: inst = 32'h5be00000;
      101341: inst = 32'h8c50000;
      101342: inst = 32'h24612800;
      101343: inst = 32'h10a00000;
      101344: inst = 32'hca00011;
      101345: inst = 32'h24822800;
      101346: inst = 32'h10a00000;
      101347: inst = 32'hca00004;
      101348: inst = 32'h38632800;
      101349: inst = 32'h38842800;
      101350: inst = 32'h10a00001;
      101351: inst = 32'hca08beb;
      101352: inst = 32'h13e00001;
      101353: inst = 32'hfe0d96a;
      101354: inst = 32'h5be00000;
      101355: inst = 32'h8c50000;
      101356: inst = 32'h24612800;
      101357: inst = 32'h10a00000;
      101358: inst = 32'hca00011;
      101359: inst = 32'h24822800;
      101360: inst = 32'h10a00000;
      101361: inst = 32'hca00004;
      101362: inst = 32'h38632800;
      101363: inst = 32'h38842800;
      101364: inst = 32'h10a00001;
      101365: inst = 32'hca08bf9;
      101366: inst = 32'h13e00001;
      101367: inst = 32'hfe0d96a;
      101368: inst = 32'h5be00000;
      101369: inst = 32'h8c50000;
      101370: inst = 32'h24612800;
      101371: inst = 32'h10a00000;
      101372: inst = 32'hca00011;
      101373: inst = 32'h24822800;
      101374: inst = 32'h10a00000;
      101375: inst = 32'hca00004;
      101376: inst = 32'h38632800;
      101377: inst = 32'h38842800;
      101378: inst = 32'h10a00001;
      101379: inst = 32'hca08c07;
      101380: inst = 32'h13e00001;
      101381: inst = 32'hfe0d96a;
      101382: inst = 32'h5be00000;
      101383: inst = 32'h8c50000;
      101384: inst = 32'h24612800;
      101385: inst = 32'h10a00000;
      101386: inst = 32'hca00011;
      101387: inst = 32'h24822800;
      101388: inst = 32'h10a00000;
      101389: inst = 32'hca00004;
      101390: inst = 32'h38632800;
      101391: inst = 32'h38842800;
      101392: inst = 32'h10a00001;
      101393: inst = 32'hca08c15;
      101394: inst = 32'h13e00001;
      101395: inst = 32'hfe0d96a;
      101396: inst = 32'h5be00000;
      101397: inst = 32'h8c50000;
      101398: inst = 32'h24612800;
      101399: inst = 32'h10a00000;
      101400: inst = 32'hca00011;
      101401: inst = 32'h24822800;
      101402: inst = 32'h10a00000;
      101403: inst = 32'hca00004;
      101404: inst = 32'h38632800;
      101405: inst = 32'h38842800;
      101406: inst = 32'h10a00001;
      101407: inst = 32'hca08c23;
      101408: inst = 32'h13e00001;
      101409: inst = 32'hfe0d96a;
      101410: inst = 32'h5be00000;
      101411: inst = 32'h8c50000;
      101412: inst = 32'h24612800;
      101413: inst = 32'h10a00000;
      101414: inst = 32'hca00011;
      101415: inst = 32'h24822800;
      101416: inst = 32'h10a00000;
      101417: inst = 32'hca00004;
      101418: inst = 32'h38632800;
      101419: inst = 32'h38842800;
      101420: inst = 32'h10a00001;
      101421: inst = 32'hca08c31;
      101422: inst = 32'h13e00001;
      101423: inst = 32'hfe0d96a;
      101424: inst = 32'h5be00000;
      101425: inst = 32'h8c50000;
      101426: inst = 32'h24612800;
      101427: inst = 32'h10a00000;
      101428: inst = 32'hca00011;
      101429: inst = 32'h24822800;
      101430: inst = 32'h10a00000;
      101431: inst = 32'hca00004;
      101432: inst = 32'h38632800;
      101433: inst = 32'h38842800;
      101434: inst = 32'h10a00001;
      101435: inst = 32'hca08c3f;
      101436: inst = 32'h13e00001;
      101437: inst = 32'hfe0d96a;
      101438: inst = 32'h5be00000;
      101439: inst = 32'h8c50000;
      101440: inst = 32'h24612800;
      101441: inst = 32'h10a00000;
      101442: inst = 32'hca00011;
      101443: inst = 32'h24822800;
      101444: inst = 32'h10a00000;
      101445: inst = 32'hca00004;
      101446: inst = 32'h38632800;
      101447: inst = 32'h38842800;
      101448: inst = 32'h10a00001;
      101449: inst = 32'hca08c4d;
      101450: inst = 32'h13e00001;
      101451: inst = 32'hfe0d96a;
      101452: inst = 32'h5be00000;
      101453: inst = 32'h8c50000;
      101454: inst = 32'h24612800;
      101455: inst = 32'h10a00000;
      101456: inst = 32'hca00011;
      101457: inst = 32'h24822800;
      101458: inst = 32'h10a00000;
      101459: inst = 32'hca00004;
      101460: inst = 32'h38632800;
      101461: inst = 32'h38842800;
      101462: inst = 32'h10a00001;
      101463: inst = 32'hca08c5b;
      101464: inst = 32'h13e00001;
      101465: inst = 32'hfe0d96a;
      101466: inst = 32'h5be00000;
      101467: inst = 32'h8c50000;
      101468: inst = 32'h24612800;
      101469: inst = 32'h10a00000;
      101470: inst = 32'hca00011;
      101471: inst = 32'h24822800;
      101472: inst = 32'h10a00000;
      101473: inst = 32'hca00004;
      101474: inst = 32'h38632800;
      101475: inst = 32'h38842800;
      101476: inst = 32'h10a00001;
      101477: inst = 32'hca08c69;
      101478: inst = 32'h13e00001;
      101479: inst = 32'hfe0d96a;
      101480: inst = 32'h5be00000;
      101481: inst = 32'h8c50000;
      101482: inst = 32'h24612800;
      101483: inst = 32'h10a00000;
      101484: inst = 32'hca00011;
      101485: inst = 32'h24822800;
      101486: inst = 32'h10a00000;
      101487: inst = 32'hca00004;
      101488: inst = 32'h38632800;
      101489: inst = 32'h38842800;
      101490: inst = 32'h10a00001;
      101491: inst = 32'hca08c77;
      101492: inst = 32'h13e00001;
      101493: inst = 32'hfe0d96a;
      101494: inst = 32'h5be00000;
      101495: inst = 32'h8c50000;
      101496: inst = 32'h24612800;
      101497: inst = 32'h10a00000;
      101498: inst = 32'hca00011;
      101499: inst = 32'h24822800;
      101500: inst = 32'h10a00000;
      101501: inst = 32'hca00004;
      101502: inst = 32'h38632800;
      101503: inst = 32'h38842800;
      101504: inst = 32'h10a00001;
      101505: inst = 32'hca08c85;
      101506: inst = 32'h13e00001;
      101507: inst = 32'hfe0d96a;
      101508: inst = 32'h5be00000;
      101509: inst = 32'h8c50000;
      101510: inst = 32'h24612800;
      101511: inst = 32'h10a00000;
      101512: inst = 32'hca00011;
      101513: inst = 32'h24822800;
      101514: inst = 32'h10a00000;
      101515: inst = 32'hca00004;
      101516: inst = 32'h38632800;
      101517: inst = 32'h38842800;
      101518: inst = 32'h10a00001;
      101519: inst = 32'hca08c93;
      101520: inst = 32'h13e00001;
      101521: inst = 32'hfe0d96a;
      101522: inst = 32'h5be00000;
      101523: inst = 32'h8c50000;
      101524: inst = 32'h24612800;
      101525: inst = 32'h10a00000;
      101526: inst = 32'hca00011;
      101527: inst = 32'h24822800;
      101528: inst = 32'h10a00000;
      101529: inst = 32'hca00004;
      101530: inst = 32'h38632800;
      101531: inst = 32'h38842800;
      101532: inst = 32'h10a00001;
      101533: inst = 32'hca08ca1;
      101534: inst = 32'h13e00001;
      101535: inst = 32'hfe0d96a;
      101536: inst = 32'h5be00000;
      101537: inst = 32'h8c50000;
      101538: inst = 32'h24612800;
      101539: inst = 32'h10a00000;
      101540: inst = 32'hca00011;
      101541: inst = 32'h24822800;
      101542: inst = 32'h10a00000;
      101543: inst = 32'hca00004;
      101544: inst = 32'h38632800;
      101545: inst = 32'h38842800;
      101546: inst = 32'h10a00001;
      101547: inst = 32'hca08caf;
      101548: inst = 32'h13e00001;
      101549: inst = 32'hfe0d96a;
      101550: inst = 32'h5be00000;
      101551: inst = 32'h8c50000;
      101552: inst = 32'h24612800;
      101553: inst = 32'h10a00000;
      101554: inst = 32'hca00011;
      101555: inst = 32'h24822800;
      101556: inst = 32'h10a00000;
      101557: inst = 32'hca00004;
      101558: inst = 32'h38632800;
      101559: inst = 32'h38842800;
      101560: inst = 32'h10a00001;
      101561: inst = 32'hca08cbd;
      101562: inst = 32'h13e00001;
      101563: inst = 32'hfe0d96a;
      101564: inst = 32'h5be00000;
      101565: inst = 32'h8c50000;
      101566: inst = 32'h24612800;
      101567: inst = 32'h10a00000;
      101568: inst = 32'hca00011;
      101569: inst = 32'h24822800;
      101570: inst = 32'h10a00000;
      101571: inst = 32'hca00004;
      101572: inst = 32'h38632800;
      101573: inst = 32'h38842800;
      101574: inst = 32'h10a00001;
      101575: inst = 32'hca08ccb;
      101576: inst = 32'h13e00001;
      101577: inst = 32'hfe0d96a;
      101578: inst = 32'h5be00000;
      101579: inst = 32'h8c50000;
      101580: inst = 32'h24612800;
      101581: inst = 32'h10a00000;
      101582: inst = 32'hca00011;
      101583: inst = 32'h24822800;
      101584: inst = 32'h10a00000;
      101585: inst = 32'hca00004;
      101586: inst = 32'h38632800;
      101587: inst = 32'h38842800;
      101588: inst = 32'h10a00001;
      101589: inst = 32'hca08cd9;
      101590: inst = 32'h13e00001;
      101591: inst = 32'hfe0d96a;
      101592: inst = 32'h5be00000;
      101593: inst = 32'h8c50000;
      101594: inst = 32'h24612800;
      101595: inst = 32'h10a00000;
      101596: inst = 32'hca00011;
      101597: inst = 32'h24822800;
      101598: inst = 32'h10a00000;
      101599: inst = 32'hca00004;
      101600: inst = 32'h38632800;
      101601: inst = 32'h38842800;
      101602: inst = 32'h10a00001;
      101603: inst = 32'hca08ce7;
      101604: inst = 32'h13e00001;
      101605: inst = 32'hfe0d96a;
      101606: inst = 32'h5be00000;
      101607: inst = 32'h8c50000;
      101608: inst = 32'h24612800;
      101609: inst = 32'h10a00000;
      101610: inst = 32'hca00011;
      101611: inst = 32'h24822800;
      101612: inst = 32'h10a00000;
      101613: inst = 32'hca00004;
      101614: inst = 32'h38632800;
      101615: inst = 32'h38842800;
      101616: inst = 32'h10a00001;
      101617: inst = 32'hca08cf5;
      101618: inst = 32'h13e00001;
      101619: inst = 32'hfe0d96a;
      101620: inst = 32'h5be00000;
      101621: inst = 32'h8c50000;
      101622: inst = 32'h24612800;
      101623: inst = 32'h10a00000;
      101624: inst = 32'hca00011;
      101625: inst = 32'h24822800;
      101626: inst = 32'h10a00000;
      101627: inst = 32'hca00004;
      101628: inst = 32'h38632800;
      101629: inst = 32'h38842800;
      101630: inst = 32'h10a00001;
      101631: inst = 32'hca08d03;
      101632: inst = 32'h13e00001;
      101633: inst = 32'hfe0d96a;
      101634: inst = 32'h5be00000;
      101635: inst = 32'h8c50000;
      101636: inst = 32'h24612800;
      101637: inst = 32'h10a00000;
      101638: inst = 32'hca00011;
      101639: inst = 32'h24822800;
      101640: inst = 32'h10a00000;
      101641: inst = 32'hca00004;
      101642: inst = 32'h38632800;
      101643: inst = 32'h38842800;
      101644: inst = 32'h10a00001;
      101645: inst = 32'hca08d11;
      101646: inst = 32'h13e00001;
      101647: inst = 32'hfe0d96a;
      101648: inst = 32'h5be00000;
      101649: inst = 32'h8c50000;
      101650: inst = 32'h24612800;
      101651: inst = 32'h10a00000;
      101652: inst = 32'hca00011;
      101653: inst = 32'h24822800;
      101654: inst = 32'h10a00000;
      101655: inst = 32'hca00004;
      101656: inst = 32'h38632800;
      101657: inst = 32'h38842800;
      101658: inst = 32'h10a00001;
      101659: inst = 32'hca08d1f;
      101660: inst = 32'h13e00001;
      101661: inst = 32'hfe0d96a;
      101662: inst = 32'h5be00000;
      101663: inst = 32'h8c50000;
      101664: inst = 32'h24612800;
      101665: inst = 32'h10a00000;
      101666: inst = 32'hca00011;
      101667: inst = 32'h24822800;
      101668: inst = 32'h10a00000;
      101669: inst = 32'hca00004;
      101670: inst = 32'h38632800;
      101671: inst = 32'h38842800;
      101672: inst = 32'h10a00001;
      101673: inst = 32'hca08d2d;
      101674: inst = 32'h13e00001;
      101675: inst = 32'hfe0d96a;
      101676: inst = 32'h5be00000;
      101677: inst = 32'h8c50000;
      101678: inst = 32'h24612800;
      101679: inst = 32'h10a00000;
      101680: inst = 32'hca00011;
      101681: inst = 32'h24822800;
      101682: inst = 32'h10a00000;
      101683: inst = 32'hca00004;
      101684: inst = 32'h38632800;
      101685: inst = 32'h38842800;
      101686: inst = 32'h10a00001;
      101687: inst = 32'hca08d3b;
      101688: inst = 32'h13e00001;
      101689: inst = 32'hfe0d96a;
      101690: inst = 32'h5be00000;
      101691: inst = 32'h8c50000;
      101692: inst = 32'h24612800;
      101693: inst = 32'h10a00000;
      101694: inst = 32'hca00011;
      101695: inst = 32'h24822800;
      101696: inst = 32'h10a00000;
      101697: inst = 32'hca00004;
      101698: inst = 32'h38632800;
      101699: inst = 32'h38842800;
      101700: inst = 32'h10a00001;
      101701: inst = 32'hca08d49;
      101702: inst = 32'h13e00001;
      101703: inst = 32'hfe0d96a;
      101704: inst = 32'h5be00000;
      101705: inst = 32'h8c50000;
      101706: inst = 32'h24612800;
      101707: inst = 32'h10a00000;
      101708: inst = 32'hca00011;
      101709: inst = 32'h24822800;
      101710: inst = 32'h10a00000;
      101711: inst = 32'hca00004;
      101712: inst = 32'h38632800;
      101713: inst = 32'h38842800;
      101714: inst = 32'h10a00001;
      101715: inst = 32'hca08d57;
      101716: inst = 32'h13e00001;
      101717: inst = 32'hfe0d96a;
      101718: inst = 32'h5be00000;
      101719: inst = 32'h8c50000;
      101720: inst = 32'h24612800;
      101721: inst = 32'h10a00000;
      101722: inst = 32'hca00011;
      101723: inst = 32'h24822800;
      101724: inst = 32'h10a00000;
      101725: inst = 32'hca00004;
      101726: inst = 32'h38632800;
      101727: inst = 32'h38842800;
      101728: inst = 32'h10a00001;
      101729: inst = 32'hca08d65;
      101730: inst = 32'h13e00001;
      101731: inst = 32'hfe0d96a;
      101732: inst = 32'h5be00000;
      101733: inst = 32'h8c50000;
      101734: inst = 32'h24612800;
      101735: inst = 32'h10a00000;
      101736: inst = 32'hca00011;
      101737: inst = 32'h24822800;
      101738: inst = 32'h10a00000;
      101739: inst = 32'hca00004;
      101740: inst = 32'h38632800;
      101741: inst = 32'h38842800;
      101742: inst = 32'h10a00001;
      101743: inst = 32'hca08d73;
      101744: inst = 32'h13e00001;
      101745: inst = 32'hfe0d96a;
      101746: inst = 32'h5be00000;
      101747: inst = 32'h8c50000;
      101748: inst = 32'h24612800;
      101749: inst = 32'h10a00000;
      101750: inst = 32'hca00011;
      101751: inst = 32'h24822800;
      101752: inst = 32'h10a00000;
      101753: inst = 32'hca00004;
      101754: inst = 32'h38632800;
      101755: inst = 32'h38842800;
      101756: inst = 32'h10a00001;
      101757: inst = 32'hca08d81;
      101758: inst = 32'h13e00001;
      101759: inst = 32'hfe0d96a;
      101760: inst = 32'h5be00000;
      101761: inst = 32'h8c50000;
      101762: inst = 32'h24612800;
      101763: inst = 32'h10a00000;
      101764: inst = 32'hca00011;
      101765: inst = 32'h24822800;
      101766: inst = 32'h10a00000;
      101767: inst = 32'hca00004;
      101768: inst = 32'h38632800;
      101769: inst = 32'h38842800;
      101770: inst = 32'h10a00001;
      101771: inst = 32'hca08d8f;
      101772: inst = 32'h13e00001;
      101773: inst = 32'hfe0d96a;
      101774: inst = 32'h5be00000;
      101775: inst = 32'h8c50000;
      101776: inst = 32'h24612800;
      101777: inst = 32'h10a00000;
      101778: inst = 32'hca00011;
      101779: inst = 32'h24822800;
      101780: inst = 32'h10a00000;
      101781: inst = 32'hca00004;
      101782: inst = 32'h38632800;
      101783: inst = 32'h38842800;
      101784: inst = 32'h10a00001;
      101785: inst = 32'hca08d9d;
      101786: inst = 32'h13e00001;
      101787: inst = 32'hfe0d96a;
      101788: inst = 32'h5be00000;
      101789: inst = 32'h8c50000;
      101790: inst = 32'h24612800;
      101791: inst = 32'h10a00000;
      101792: inst = 32'hca00011;
      101793: inst = 32'h24822800;
      101794: inst = 32'h10a00000;
      101795: inst = 32'hca00004;
      101796: inst = 32'h38632800;
      101797: inst = 32'h38842800;
      101798: inst = 32'h10a00001;
      101799: inst = 32'hca08dab;
      101800: inst = 32'h13e00001;
      101801: inst = 32'hfe0d96a;
      101802: inst = 32'h5be00000;
      101803: inst = 32'h8c50000;
      101804: inst = 32'h24612800;
      101805: inst = 32'h10a00000;
      101806: inst = 32'hca00011;
      101807: inst = 32'h24822800;
      101808: inst = 32'h10a00000;
      101809: inst = 32'hca00004;
      101810: inst = 32'h38632800;
      101811: inst = 32'h38842800;
      101812: inst = 32'h10a00001;
      101813: inst = 32'hca08db9;
      101814: inst = 32'h13e00001;
      101815: inst = 32'hfe0d96a;
      101816: inst = 32'h5be00000;
      101817: inst = 32'h8c50000;
      101818: inst = 32'h24612800;
      101819: inst = 32'h10a00000;
      101820: inst = 32'hca00011;
      101821: inst = 32'h24822800;
      101822: inst = 32'h10a00000;
      101823: inst = 32'hca00004;
      101824: inst = 32'h38632800;
      101825: inst = 32'h38842800;
      101826: inst = 32'h10a00001;
      101827: inst = 32'hca08dc7;
      101828: inst = 32'h13e00001;
      101829: inst = 32'hfe0d96a;
      101830: inst = 32'h5be00000;
      101831: inst = 32'h8c50000;
      101832: inst = 32'h24612800;
      101833: inst = 32'h10a00000;
      101834: inst = 32'hca00011;
      101835: inst = 32'h24822800;
      101836: inst = 32'h10a00000;
      101837: inst = 32'hca00004;
      101838: inst = 32'h38632800;
      101839: inst = 32'h38842800;
      101840: inst = 32'h10a00001;
      101841: inst = 32'hca08dd5;
      101842: inst = 32'h13e00001;
      101843: inst = 32'hfe0d96a;
      101844: inst = 32'h5be00000;
      101845: inst = 32'h8c50000;
      101846: inst = 32'h24612800;
      101847: inst = 32'h10a00000;
      101848: inst = 32'hca00011;
      101849: inst = 32'h24822800;
      101850: inst = 32'h10a00000;
      101851: inst = 32'hca00004;
      101852: inst = 32'h38632800;
      101853: inst = 32'h38842800;
      101854: inst = 32'h10a00001;
      101855: inst = 32'hca08de3;
      101856: inst = 32'h13e00001;
      101857: inst = 32'hfe0d96a;
      101858: inst = 32'h5be00000;
      101859: inst = 32'h8c50000;
      101860: inst = 32'h24612800;
      101861: inst = 32'h10a00000;
      101862: inst = 32'hca00011;
      101863: inst = 32'h24822800;
      101864: inst = 32'h10a00000;
      101865: inst = 32'hca00004;
      101866: inst = 32'h38632800;
      101867: inst = 32'h38842800;
      101868: inst = 32'h10a00001;
      101869: inst = 32'hca08df1;
      101870: inst = 32'h13e00001;
      101871: inst = 32'hfe0d96a;
      101872: inst = 32'h5be00000;
      101873: inst = 32'h8c50000;
      101874: inst = 32'h24612800;
      101875: inst = 32'h10a00000;
      101876: inst = 32'hca00011;
      101877: inst = 32'h24822800;
      101878: inst = 32'h10a00000;
      101879: inst = 32'hca00004;
      101880: inst = 32'h38632800;
      101881: inst = 32'h38842800;
      101882: inst = 32'h10a00001;
      101883: inst = 32'hca08dff;
      101884: inst = 32'h13e00001;
      101885: inst = 32'hfe0d96a;
      101886: inst = 32'h5be00000;
      101887: inst = 32'h8c50000;
      101888: inst = 32'h24612800;
      101889: inst = 32'h10a00000;
      101890: inst = 32'hca00011;
      101891: inst = 32'h24822800;
      101892: inst = 32'h10a00000;
      101893: inst = 32'hca00004;
      101894: inst = 32'h38632800;
      101895: inst = 32'h38842800;
      101896: inst = 32'h10a00001;
      101897: inst = 32'hca08e0d;
      101898: inst = 32'h13e00001;
      101899: inst = 32'hfe0d96a;
      101900: inst = 32'h5be00000;
      101901: inst = 32'h8c50000;
      101902: inst = 32'h24612800;
      101903: inst = 32'h10a00000;
      101904: inst = 32'hca00011;
      101905: inst = 32'h24822800;
      101906: inst = 32'h10a00000;
      101907: inst = 32'hca00004;
      101908: inst = 32'h38632800;
      101909: inst = 32'h38842800;
      101910: inst = 32'h10a00001;
      101911: inst = 32'hca08e1b;
      101912: inst = 32'h13e00001;
      101913: inst = 32'hfe0d96a;
      101914: inst = 32'h5be00000;
      101915: inst = 32'h8c50000;
      101916: inst = 32'h24612800;
      101917: inst = 32'h10a00000;
      101918: inst = 32'hca00011;
      101919: inst = 32'h24822800;
      101920: inst = 32'h10a00000;
      101921: inst = 32'hca00004;
      101922: inst = 32'h38632800;
      101923: inst = 32'h38842800;
      101924: inst = 32'h10a00001;
      101925: inst = 32'hca08e29;
      101926: inst = 32'h13e00001;
      101927: inst = 32'hfe0d96a;
      101928: inst = 32'h5be00000;
      101929: inst = 32'h8c50000;
      101930: inst = 32'h24612800;
      101931: inst = 32'h10a00000;
      101932: inst = 32'hca00011;
      101933: inst = 32'h24822800;
      101934: inst = 32'h10a00000;
      101935: inst = 32'hca00004;
      101936: inst = 32'h38632800;
      101937: inst = 32'h38842800;
      101938: inst = 32'h10a00001;
      101939: inst = 32'hca08e37;
      101940: inst = 32'h13e00001;
      101941: inst = 32'hfe0d96a;
      101942: inst = 32'h5be00000;
      101943: inst = 32'h8c50000;
      101944: inst = 32'h24612800;
      101945: inst = 32'h10a00000;
      101946: inst = 32'hca00011;
      101947: inst = 32'h24822800;
      101948: inst = 32'h10a00000;
      101949: inst = 32'hca00004;
      101950: inst = 32'h38632800;
      101951: inst = 32'h38842800;
      101952: inst = 32'h10a00001;
      101953: inst = 32'hca08e45;
      101954: inst = 32'h13e00001;
      101955: inst = 32'hfe0d96a;
      101956: inst = 32'h5be00000;
      101957: inst = 32'h8c50000;
      101958: inst = 32'h24612800;
      101959: inst = 32'h10a00000;
      101960: inst = 32'hca00011;
      101961: inst = 32'h24822800;
      101962: inst = 32'h10a00000;
      101963: inst = 32'hca00004;
      101964: inst = 32'h38632800;
      101965: inst = 32'h38842800;
      101966: inst = 32'h10a00001;
      101967: inst = 32'hca08e53;
      101968: inst = 32'h13e00001;
      101969: inst = 32'hfe0d96a;
      101970: inst = 32'h5be00000;
      101971: inst = 32'h8c50000;
      101972: inst = 32'h24612800;
      101973: inst = 32'h10a00000;
      101974: inst = 32'hca00011;
      101975: inst = 32'h24822800;
      101976: inst = 32'h10a00000;
      101977: inst = 32'hca00004;
      101978: inst = 32'h38632800;
      101979: inst = 32'h38842800;
      101980: inst = 32'h10a00001;
      101981: inst = 32'hca08e61;
      101982: inst = 32'h13e00001;
      101983: inst = 32'hfe0d96a;
      101984: inst = 32'h5be00000;
      101985: inst = 32'h8c50000;
      101986: inst = 32'h24612800;
      101987: inst = 32'h10a00000;
      101988: inst = 32'hca00011;
      101989: inst = 32'h24822800;
      101990: inst = 32'h10a00000;
      101991: inst = 32'hca00004;
      101992: inst = 32'h38632800;
      101993: inst = 32'h38842800;
      101994: inst = 32'h10a00001;
      101995: inst = 32'hca08e6f;
      101996: inst = 32'h13e00001;
      101997: inst = 32'hfe0d96a;
      101998: inst = 32'h5be00000;
      101999: inst = 32'h8c50000;
      102000: inst = 32'h24612800;
      102001: inst = 32'h10a00000;
      102002: inst = 32'hca00011;
      102003: inst = 32'h24822800;
      102004: inst = 32'h10a00000;
      102005: inst = 32'hca00004;
      102006: inst = 32'h38632800;
      102007: inst = 32'h38842800;
      102008: inst = 32'h10a00001;
      102009: inst = 32'hca08e7d;
      102010: inst = 32'h13e00001;
      102011: inst = 32'hfe0d96a;
      102012: inst = 32'h5be00000;
      102013: inst = 32'h8c50000;
      102014: inst = 32'h24612800;
      102015: inst = 32'h10a00000;
      102016: inst = 32'hca00011;
      102017: inst = 32'h24822800;
      102018: inst = 32'h10a00000;
      102019: inst = 32'hca00004;
      102020: inst = 32'h38632800;
      102021: inst = 32'h38842800;
      102022: inst = 32'h10a00001;
      102023: inst = 32'hca08e8b;
      102024: inst = 32'h13e00001;
      102025: inst = 32'hfe0d96a;
      102026: inst = 32'h5be00000;
      102027: inst = 32'h8c50000;
      102028: inst = 32'h24612800;
      102029: inst = 32'h10a00000;
      102030: inst = 32'hca00011;
      102031: inst = 32'h24822800;
      102032: inst = 32'h10a00000;
      102033: inst = 32'hca00004;
      102034: inst = 32'h38632800;
      102035: inst = 32'h38842800;
      102036: inst = 32'h10a00001;
      102037: inst = 32'hca08e99;
      102038: inst = 32'h13e00001;
      102039: inst = 32'hfe0d96a;
      102040: inst = 32'h5be00000;
      102041: inst = 32'h8c50000;
      102042: inst = 32'h24612800;
      102043: inst = 32'h10a00000;
      102044: inst = 32'hca00011;
      102045: inst = 32'h24822800;
      102046: inst = 32'h10a00000;
      102047: inst = 32'hca00004;
      102048: inst = 32'h38632800;
      102049: inst = 32'h38842800;
      102050: inst = 32'h10a00001;
      102051: inst = 32'hca08ea7;
      102052: inst = 32'h13e00001;
      102053: inst = 32'hfe0d96a;
      102054: inst = 32'h5be00000;
      102055: inst = 32'h8c50000;
      102056: inst = 32'h24612800;
      102057: inst = 32'h10a00000;
      102058: inst = 32'hca00011;
      102059: inst = 32'h24822800;
      102060: inst = 32'h10a00000;
      102061: inst = 32'hca00004;
      102062: inst = 32'h38632800;
      102063: inst = 32'h38842800;
      102064: inst = 32'h10a00001;
      102065: inst = 32'hca08eb5;
      102066: inst = 32'h13e00001;
      102067: inst = 32'hfe0d96a;
      102068: inst = 32'h5be00000;
      102069: inst = 32'h8c50000;
      102070: inst = 32'h24612800;
      102071: inst = 32'h10a00000;
      102072: inst = 32'hca00011;
      102073: inst = 32'h24822800;
      102074: inst = 32'h10a00000;
      102075: inst = 32'hca00004;
      102076: inst = 32'h38632800;
      102077: inst = 32'h38842800;
      102078: inst = 32'h10a00001;
      102079: inst = 32'hca08ec3;
      102080: inst = 32'h13e00001;
      102081: inst = 32'hfe0d96a;
      102082: inst = 32'h5be00000;
      102083: inst = 32'h8c50000;
      102084: inst = 32'h24612800;
      102085: inst = 32'h10a00000;
      102086: inst = 32'hca00011;
      102087: inst = 32'h24822800;
      102088: inst = 32'h10a00000;
      102089: inst = 32'hca00004;
      102090: inst = 32'h38632800;
      102091: inst = 32'h38842800;
      102092: inst = 32'h10a00001;
      102093: inst = 32'hca08ed1;
      102094: inst = 32'h13e00001;
      102095: inst = 32'hfe0d96a;
      102096: inst = 32'h5be00000;
      102097: inst = 32'h8c50000;
      102098: inst = 32'h24612800;
      102099: inst = 32'h10a00000;
      102100: inst = 32'hca00011;
      102101: inst = 32'h24822800;
      102102: inst = 32'h10a00000;
      102103: inst = 32'hca00004;
      102104: inst = 32'h38632800;
      102105: inst = 32'h38842800;
      102106: inst = 32'h10a00001;
      102107: inst = 32'hca08edf;
      102108: inst = 32'h13e00001;
      102109: inst = 32'hfe0d96a;
      102110: inst = 32'h5be00000;
      102111: inst = 32'h8c50000;
      102112: inst = 32'h24612800;
      102113: inst = 32'h10a00000;
      102114: inst = 32'hca00011;
      102115: inst = 32'h24822800;
      102116: inst = 32'h10a00000;
      102117: inst = 32'hca00004;
      102118: inst = 32'h38632800;
      102119: inst = 32'h38842800;
      102120: inst = 32'h10a00001;
      102121: inst = 32'hca08eed;
      102122: inst = 32'h13e00001;
      102123: inst = 32'hfe0d96a;
      102124: inst = 32'h5be00000;
      102125: inst = 32'h8c50000;
      102126: inst = 32'h24612800;
      102127: inst = 32'h10a00000;
      102128: inst = 32'hca00011;
      102129: inst = 32'h24822800;
      102130: inst = 32'h10a00000;
      102131: inst = 32'hca00004;
      102132: inst = 32'h38632800;
      102133: inst = 32'h38842800;
      102134: inst = 32'h10a00001;
      102135: inst = 32'hca08efb;
      102136: inst = 32'h13e00001;
      102137: inst = 32'hfe0d96a;
      102138: inst = 32'h5be00000;
      102139: inst = 32'h8c50000;
      102140: inst = 32'h24612800;
      102141: inst = 32'h10a00000;
      102142: inst = 32'hca00011;
      102143: inst = 32'h24822800;
      102144: inst = 32'h10a00000;
      102145: inst = 32'hca00004;
      102146: inst = 32'h38632800;
      102147: inst = 32'h38842800;
      102148: inst = 32'h10a00001;
      102149: inst = 32'hca08f09;
      102150: inst = 32'h13e00001;
      102151: inst = 32'hfe0d96a;
      102152: inst = 32'h5be00000;
      102153: inst = 32'h8c50000;
      102154: inst = 32'h24612800;
      102155: inst = 32'h10a00000;
      102156: inst = 32'hca00011;
      102157: inst = 32'h24822800;
      102158: inst = 32'h10a00000;
      102159: inst = 32'hca00004;
      102160: inst = 32'h38632800;
      102161: inst = 32'h38842800;
      102162: inst = 32'h10a00001;
      102163: inst = 32'hca08f17;
      102164: inst = 32'h13e00001;
      102165: inst = 32'hfe0d96a;
      102166: inst = 32'h5be00000;
      102167: inst = 32'h8c50000;
      102168: inst = 32'h24612800;
      102169: inst = 32'h10a00000;
      102170: inst = 32'hca00011;
      102171: inst = 32'h24822800;
      102172: inst = 32'h10a00000;
      102173: inst = 32'hca00004;
      102174: inst = 32'h38632800;
      102175: inst = 32'h38842800;
      102176: inst = 32'h10a00001;
      102177: inst = 32'hca08f25;
      102178: inst = 32'h13e00001;
      102179: inst = 32'hfe0d96a;
      102180: inst = 32'h5be00000;
      102181: inst = 32'h8c50000;
      102182: inst = 32'h24612800;
      102183: inst = 32'h10a00000;
      102184: inst = 32'hca00011;
      102185: inst = 32'h24822800;
      102186: inst = 32'h10a00000;
      102187: inst = 32'hca00004;
      102188: inst = 32'h38632800;
      102189: inst = 32'h38842800;
      102190: inst = 32'h10a00001;
      102191: inst = 32'hca08f33;
      102192: inst = 32'h13e00001;
      102193: inst = 32'hfe0d96a;
      102194: inst = 32'h5be00000;
      102195: inst = 32'h8c50000;
      102196: inst = 32'h24612800;
      102197: inst = 32'h10a00000;
      102198: inst = 32'hca00011;
      102199: inst = 32'h24822800;
      102200: inst = 32'h10a00000;
      102201: inst = 32'hca00004;
      102202: inst = 32'h38632800;
      102203: inst = 32'h38842800;
      102204: inst = 32'h10a00001;
      102205: inst = 32'hca08f41;
      102206: inst = 32'h13e00001;
      102207: inst = 32'hfe0d96a;
      102208: inst = 32'h5be00000;
      102209: inst = 32'h8c50000;
      102210: inst = 32'h24612800;
      102211: inst = 32'h10a00000;
      102212: inst = 32'hca00011;
      102213: inst = 32'h24822800;
      102214: inst = 32'h10a00000;
      102215: inst = 32'hca00004;
      102216: inst = 32'h38632800;
      102217: inst = 32'h38842800;
      102218: inst = 32'h10a00001;
      102219: inst = 32'hca08f4f;
      102220: inst = 32'h13e00001;
      102221: inst = 32'hfe0d96a;
      102222: inst = 32'h5be00000;
      102223: inst = 32'h8c50000;
      102224: inst = 32'h24612800;
      102225: inst = 32'h10a00000;
      102226: inst = 32'hca00011;
      102227: inst = 32'h24822800;
      102228: inst = 32'h10a00000;
      102229: inst = 32'hca00004;
      102230: inst = 32'h38632800;
      102231: inst = 32'h38842800;
      102232: inst = 32'h10a00001;
      102233: inst = 32'hca08f5d;
      102234: inst = 32'h13e00001;
      102235: inst = 32'hfe0d96a;
      102236: inst = 32'h5be00000;
      102237: inst = 32'h8c50000;
      102238: inst = 32'h24612800;
      102239: inst = 32'h10a00000;
      102240: inst = 32'hca00011;
      102241: inst = 32'h24822800;
      102242: inst = 32'h10a00000;
      102243: inst = 32'hca00004;
      102244: inst = 32'h38632800;
      102245: inst = 32'h38842800;
      102246: inst = 32'h10a00001;
      102247: inst = 32'hca08f6b;
      102248: inst = 32'h13e00001;
      102249: inst = 32'hfe0d96a;
      102250: inst = 32'h5be00000;
      102251: inst = 32'h8c50000;
      102252: inst = 32'h24612800;
      102253: inst = 32'h10a00000;
      102254: inst = 32'hca00011;
      102255: inst = 32'h24822800;
      102256: inst = 32'h10a00000;
      102257: inst = 32'hca00004;
      102258: inst = 32'h38632800;
      102259: inst = 32'h38842800;
      102260: inst = 32'h10a00001;
      102261: inst = 32'hca08f79;
      102262: inst = 32'h13e00001;
      102263: inst = 32'hfe0d96a;
      102264: inst = 32'h5be00000;
      102265: inst = 32'h8c50000;
      102266: inst = 32'h24612800;
      102267: inst = 32'h10a00000;
      102268: inst = 32'hca00011;
      102269: inst = 32'h24822800;
      102270: inst = 32'h10a00000;
      102271: inst = 32'hca00004;
      102272: inst = 32'h38632800;
      102273: inst = 32'h38842800;
      102274: inst = 32'h10a00001;
      102275: inst = 32'hca08f87;
      102276: inst = 32'h13e00001;
      102277: inst = 32'hfe0d96a;
      102278: inst = 32'h5be00000;
      102279: inst = 32'h8c50000;
      102280: inst = 32'h24612800;
      102281: inst = 32'h10a00000;
      102282: inst = 32'hca00011;
      102283: inst = 32'h24822800;
      102284: inst = 32'h10a00000;
      102285: inst = 32'hca00004;
      102286: inst = 32'h38632800;
      102287: inst = 32'h38842800;
      102288: inst = 32'h10a00001;
      102289: inst = 32'hca08f95;
      102290: inst = 32'h13e00001;
      102291: inst = 32'hfe0d96a;
      102292: inst = 32'h5be00000;
      102293: inst = 32'h8c50000;
      102294: inst = 32'h24612800;
      102295: inst = 32'h10a00000;
      102296: inst = 32'hca00011;
      102297: inst = 32'h24822800;
      102298: inst = 32'h10a00000;
      102299: inst = 32'hca00004;
      102300: inst = 32'h38632800;
      102301: inst = 32'h38842800;
      102302: inst = 32'h10a00001;
      102303: inst = 32'hca08fa3;
      102304: inst = 32'h13e00001;
      102305: inst = 32'hfe0d96a;
      102306: inst = 32'h5be00000;
      102307: inst = 32'h8c50000;
      102308: inst = 32'h24612800;
      102309: inst = 32'h10a00000;
      102310: inst = 32'hca00011;
      102311: inst = 32'h24822800;
      102312: inst = 32'h10a00000;
      102313: inst = 32'hca00004;
      102314: inst = 32'h38632800;
      102315: inst = 32'h38842800;
      102316: inst = 32'h10a00001;
      102317: inst = 32'hca08fb1;
      102318: inst = 32'h13e00001;
      102319: inst = 32'hfe0d96a;
      102320: inst = 32'h5be00000;
      102321: inst = 32'h8c50000;
      102322: inst = 32'h24612800;
      102323: inst = 32'h10a00000;
      102324: inst = 32'hca00011;
      102325: inst = 32'h24822800;
      102326: inst = 32'h10a00000;
      102327: inst = 32'hca00004;
      102328: inst = 32'h38632800;
      102329: inst = 32'h38842800;
      102330: inst = 32'h10a00001;
      102331: inst = 32'hca08fbf;
      102332: inst = 32'h13e00001;
      102333: inst = 32'hfe0d96a;
      102334: inst = 32'h5be00000;
      102335: inst = 32'h8c50000;
      102336: inst = 32'h24612800;
      102337: inst = 32'h10a00000;
      102338: inst = 32'hca00011;
      102339: inst = 32'h24822800;
      102340: inst = 32'h10a00000;
      102341: inst = 32'hca00004;
      102342: inst = 32'h38632800;
      102343: inst = 32'h38842800;
      102344: inst = 32'h10a00001;
      102345: inst = 32'hca08fcd;
      102346: inst = 32'h13e00001;
      102347: inst = 32'hfe0d96a;
      102348: inst = 32'h5be00000;
      102349: inst = 32'h8c50000;
      102350: inst = 32'h24612800;
      102351: inst = 32'h10a00000;
      102352: inst = 32'hca00011;
      102353: inst = 32'h24822800;
      102354: inst = 32'h10a00000;
      102355: inst = 32'hca00004;
      102356: inst = 32'h38632800;
      102357: inst = 32'h38842800;
      102358: inst = 32'h10a00001;
      102359: inst = 32'hca08fdb;
      102360: inst = 32'h13e00001;
      102361: inst = 32'hfe0d96a;
      102362: inst = 32'h5be00000;
      102363: inst = 32'h8c50000;
      102364: inst = 32'h24612800;
      102365: inst = 32'h10a00000;
      102366: inst = 32'hca00011;
      102367: inst = 32'h24822800;
      102368: inst = 32'h10a00000;
      102369: inst = 32'hca00004;
      102370: inst = 32'h38632800;
      102371: inst = 32'h38842800;
      102372: inst = 32'h10a00001;
      102373: inst = 32'hca08fe9;
      102374: inst = 32'h13e00001;
      102375: inst = 32'hfe0d96a;
      102376: inst = 32'h5be00000;
      102377: inst = 32'h8c50000;
      102378: inst = 32'h24612800;
      102379: inst = 32'h10a00000;
      102380: inst = 32'hca00012;
      102381: inst = 32'h24822800;
      102382: inst = 32'h10a00000;
      102383: inst = 32'hca00004;
      102384: inst = 32'h38632800;
      102385: inst = 32'h38842800;
      102386: inst = 32'h10a00001;
      102387: inst = 32'hca08ff7;
      102388: inst = 32'h13e00001;
      102389: inst = 32'hfe0d96a;
      102390: inst = 32'h5be00000;
      102391: inst = 32'h8c50000;
      102392: inst = 32'h24612800;
      102393: inst = 32'h10a00000;
      102394: inst = 32'hca00012;
      102395: inst = 32'h24822800;
      102396: inst = 32'h10a00000;
      102397: inst = 32'hca00004;
      102398: inst = 32'h38632800;
      102399: inst = 32'h38842800;
      102400: inst = 32'h10a00001;
      102401: inst = 32'hca09005;
      102402: inst = 32'h13e00001;
      102403: inst = 32'hfe0d96a;
      102404: inst = 32'h5be00000;
      102405: inst = 32'h8c50000;
      102406: inst = 32'h24612800;
      102407: inst = 32'h10a00000;
      102408: inst = 32'hca00012;
      102409: inst = 32'h24822800;
      102410: inst = 32'h10a00000;
      102411: inst = 32'hca00004;
      102412: inst = 32'h38632800;
      102413: inst = 32'h38842800;
      102414: inst = 32'h10a00001;
      102415: inst = 32'hca09013;
      102416: inst = 32'h13e00001;
      102417: inst = 32'hfe0d96a;
      102418: inst = 32'h5be00000;
      102419: inst = 32'h8c50000;
      102420: inst = 32'h24612800;
      102421: inst = 32'h10a00000;
      102422: inst = 32'hca00012;
      102423: inst = 32'h24822800;
      102424: inst = 32'h10a00000;
      102425: inst = 32'hca00004;
      102426: inst = 32'h38632800;
      102427: inst = 32'h38842800;
      102428: inst = 32'h10a00001;
      102429: inst = 32'hca09021;
      102430: inst = 32'h13e00001;
      102431: inst = 32'hfe0d96a;
      102432: inst = 32'h5be00000;
      102433: inst = 32'h8c50000;
      102434: inst = 32'h24612800;
      102435: inst = 32'h10a00000;
      102436: inst = 32'hca00012;
      102437: inst = 32'h24822800;
      102438: inst = 32'h10a00000;
      102439: inst = 32'hca00004;
      102440: inst = 32'h38632800;
      102441: inst = 32'h38842800;
      102442: inst = 32'h10a00001;
      102443: inst = 32'hca0902f;
      102444: inst = 32'h13e00001;
      102445: inst = 32'hfe0d96a;
      102446: inst = 32'h5be00000;
      102447: inst = 32'h8c50000;
      102448: inst = 32'h24612800;
      102449: inst = 32'h10a00000;
      102450: inst = 32'hca00012;
      102451: inst = 32'h24822800;
      102452: inst = 32'h10a00000;
      102453: inst = 32'hca00004;
      102454: inst = 32'h38632800;
      102455: inst = 32'h38842800;
      102456: inst = 32'h10a00001;
      102457: inst = 32'hca0903d;
      102458: inst = 32'h13e00001;
      102459: inst = 32'hfe0d96a;
      102460: inst = 32'h5be00000;
      102461: inst = 32'h8c50000;
      102462: inst = 32'h24612800;
      102463: inst = 32'h10a00000;
      102464: inst = 32'hca00012;
      102465: inst = 32'h24822800;
      102466: inst = 32'h10a00000;
      102467: inst = 32'hca00004;
      102468: inst = 32'h38632800;
      102469: inst = 32'h38842800;
      102470: inst = 32'h10a00001;
      102471: inst = 32'hca0904b;
      102472: inst = 32'h13e00001;
      102473: inst = 32'hfe0d96a;
      102474: inst = 32'h5be00000;
      102475: inst = 32'h8c50000;
      102476: inst = 32'h24612800;
      102477: inst = 32'h10a00000;
      102478: inst = 32'hca00012;
      102479: inst = 32'h24822800;
      102480: inst = 32'h10a00000;
      102481: inst = 32'hca00004;
      102482: inst = 32'h38632800;
      102483: inst = 32'h38842800;
      102484: inst = 32'h10a00001;
      102485: inst = 32'hca09059;
      102486: inst = 32'h13e00001;
      102487: inst = 32'hfe0d96a;
      102488: inst = 32'h5be00000;
      102489: inst = 32'h8c50000;
      102490: inst = 32'h24612800;
      102491: inst = 32'h10a00000;
      102492: inst = 32'hca00012;
      102493: inst = 32'h24822800;
      102494: inst = 32'h10a00000;
      102495: inst = 32'hca00004;
      102496: inst = 32'h38632800;
      102497: inst = 32'h38842800;
      102498: inst = 32'h10a00001;
      102499: inst = 32'hca09067;
      102500: inst = 32'h13e00001;
      102501: inst = 32'hfe0d96a;
      102502: inst = 32'h5be00000;
      102503: inst = 32'h8c50000;
      102504: inst = 32'h24612800;
      102505: inst = 32'h10a00000;
      102506: inst = 32'hca00012;
      102507: inst = 32'h24822800;
      102508: inst = 32'h10a00000;
      102509: inst = 32'hca00004;
      102510: inst = 32'h38632800;
      102511: inst = 32'h38842800;
      102512: inst = 32'h10a00001;
      102513: inst = 32'hca09075;
      102514: inst = 32'h13e00001;
      102515: inst = 32'hfe0d96a;
      102516: inst = 32'h5be00000;
      102517: inst = 32'h8c50000;
      102518: inst = 32'h24612800;
      102519: inst = 32'h10a00000;
      102520: inst = 32'hca00012;
      102521: inst = 32'h24822800;
      102522: inst = 32'h10a00000;
      102523: inst = 32'hca00004;
      102524: inst = 32'h38632800;
      102525: inst = 32'h38842800;
      102526: inst = 32'h10a00001;
      102527: inst = 32'hca09083;
      102528: inst = 32'h13e00001;
      102529: inst = 32'hfe0d96a;
      102530: inst = 32'h5be00000;
      102531: inst = 32'h8c50000;
      102532: inst = 32'h24612800;
      102533: inst = 32'h10a00000;
      102534: inst = 32'hca00012;
      102535: inst = 32'h24822800;
      102536: inst = 32'h10a00000;
      102537: inst = 32'hca00004;
      102538: inst = 32'h38632800;
      102539: inst = 32'h38842800;
      102540: inst = 32'h10a00001;
      102541: inst = 32'hca09091;
      102542: inst = 32'h13e00001;
      102543: inst = 32'hfe0d96a;
      102544: inst = 32'h5be00000;
      102545: inst = 32'h8c50000;
      102546: inst = 32'h24612800;
      102547: inst = 32'h10a00000;
      102548: inst = 32'hca00012;
      102549: inst = 32'h24822800;
      102550: inst = 32'h10a00000;
      102551: inst = 32'hca00004;
      102552: inst = 32'h38632800;
      102553: inst = 32'h38842800;
      102554: inst = 32'h10a00001;
      102555: inst = 32'hca0909f;
      102556: inst = 32'h13e00001;
      102557: inst = 32'hfe0d96a;
      102558: inst = 32'h5be00000;
      102559: inst = 32'h8c50000;
      102560: inst = 32'h24612800;
      102561: inst = 32'h10a00000;
      102562: inst = 32'hca00012;
      102563: inst = 32'h24822800;
      102564: inst = 32'h10a00000;
      102565: inst = 32'hca00004;
      102566: inst = 32'h38632800;
      102567: inst = 32'h38842800;
      102568: inst = 32'h10a00001;
      102569: inst = 32'hca090ad;
      102570: inst = 32'h13e00001;
      102571: inst = 32'hfe0d96a;
      102572: inst = 32'h5be00000;
      102573: inst = 32'h8c50000;
      102574: inst = 32'h24612800;
      102575: inst = 32'h10a00000;
      102576: inst = 32'hca00012;
      102577: inst = 32'h24822800;
      102578: inst = 32'h10a00000;
      102579: inst = 32'hca00004;
      102580: inst = 32'h38632800;
      102581: inst = 32'h38842800;
      102582: inst = 32'h10a00001;
      102583: inst = 32'hca090bb;
      102584: inst = 32'h13e00001;
      102585: inst = 32'hfe0d96a;
      102586: inst = 32'h5be00000;
      102587: inst = 32'h8c50000;
      102588: inst = 32'h24612800;
      102589: inst = 32'h10a00000;
      102590: inst = 32'hca00012;
      102591: inst = 32'h24822800;
      102592: inst = 32'h10a00000;
      102593: inst = 32'hca00004;
      102594: inst = 32'h38632800;
      102595: inst = 32'h38842800;
      102596: inst = 32'h10a00001;
      102597: inst = 32'hca090c9;
      102598: inst = 32'h13e00001;
      102599: inst = 32'hfe0d96a;
      102600: inst = 32'h5be00000;
      102601: inst = 32'h8c50000;
      102602: inst = 32'h24612800;
      102603: inst = 32'h10a00000;
      102604: inst = 32'hca00012;
      102605: inst = 32'h24822800;
      102606: inst = 32'h10a00000;
      102607: inst = 32'hca00004;
      102608: inst = 32'h38632800;
      102609: inst = 32'h38842800;
      102610: inst = 32'h10a00001;
      102611: inst = 32'hca090d7;
      102612: inst = 32'h13e00001;
      102613: inst = 32'hfe0d96a;
      102614: inst = 32'h5be00000;
      102615: inst = 32'h8c50000;
      102616: inst = 32'h24612800;
      102617: inst = 32'h10a00000;
      102618: inst = 32'hca00012;
      102619: inst = 32'h24822800;
      102620: inst = 32'h10a00000;
      102621: inst = 32'hca00004;
      102622: inst = 32'h38632800;
      102623: inst = 32'h38842800;
      102624: inst = 32'h10a00001;
      102625: inst = 32'hca090e5;
      102626: inst = 32'h13e00001;
      102627: inst = 32'hfe0d96a;
      102628: inst = 32'h5be00000;
      102629: inst = 32'h8c50000;
      102630: inst = 32'h24612800;
      102631: inst = 32'h10a00000;
      102632: inst = 32'hca00012;
      102633: inst = 32'h24822800;
      102634: inst = 32'h10a00000;
      102635: inst = 32'hca00004;
      102636: inst = 32'h38632800;
      102637: inst = 32'h38842800;
      102638: inst = 32'h10a00001;
      102639: inst = 32'hca090f3;
      102640: inst = 32'h13e00001;
      102641: inst = 32'hfe0d96a;
      102642: inst = 32'h5be00000;
      102643: inst = 32'h8c50000;
      102644: inst = 32'h24612800;
      102645: inst = 32'h10a00000;
      102646: inst = 32'hca00012;
      102647: inst = 32'h24822800;
      102648: inst = 32'h10a00000;
      102649: inst = 32'hca00004;
      102650: inst = 32'h38632800;
      102651: inst = 32'h38842800;
      102652: inst = 32'h10a00001;
      102653: inst = 32'hca09101;
      102654: inst = 32'h13e00001;
      102655: inst = 32'hfe0d96a;
      102656: inst = 32'h5be00000;
      102657: inst = 32'h8c50000;
      102658: inst = 32'h24612800;
      102659: inst = 32'h10a00000;
      102660: inst = 32'hca00012;
      102661: inst = 32'h24822800;
      102662: inst = 32'h10a00000;
      102663: inst = 32'hca00004;
      102664: inst = 32'h38632800;
      102665: inst = 32'h38842800;
      102666: inst = 32'h10a00001;
      102667: inst = 32'hca0910f;
      102668: inst = 32'h13e00001;
      102669: inst = 32'hfe0d96a;
      102670: inst = 32'h5be00000;
      102671: inst = 32'h8c50000;
      102672: inst = 32'h24612800;
      102673: inst = 32'h10a00000;
      102674: inst = 32'hca00012;
      102675: inst = 32'h24822800;
      102676: inst = 32'h10a00000;
      102677: inst = 32'hca00004;
      102678: inst = 32'h38632800;
      102679: inst = 32'h38842800;
      102680: inst = 32'h10a00001;
      102681: inst = 32'hca0911d;
      102682: inst = 32'h13e00001;
      102683: inst = 32'hfe0d96a;
      102684: inst = 32'h5be00000;
      102685: inst = 32'h8c50000;
      102686: inst = 32'h24612800;
      102687: inst = 32'h10a00000;
      102688: inst = 32'hca00012;
      102689: inst = 32'h24822800;
      102690: inst = 32'h10a00000;
      102691: inst = 32'hca00004;
      102692: inst = 32'h38632800;
      102693: inst = 32'h38842800;
      102694: inst = 32'h10a00001;
      102695: inst = 32'hca0912b;
      102696: inst = 32'h13e00001;
      102697: inst = 32'hfe0d96a;
      102698: inst = 32'h5be00000;
      102699: inst = 32'h8c50000;
      102700: inst = 32'h24612800;
      102701: inst = 32'h10a00000;
      102702: inst = 32'hca00012;
      102703: inst = 32'h24822800;
      102704: inst = 32'h10a00000;
      102705: inst = 32'hca00004;
      102706: inst = 32'h38632800;
      102707: inst = 32'h38842800;
      102708: inst = 32'h10a00001;
      102709: inst = 32'hca09139;
      102710: inst = 32'h13e00001;
      102711: inst = 32'hfe0d96a;
      102712: inst = 32'h5be00000;
      102713: inst = 32'h8c50000;
      102714: inst = 32'h24612800;
      102715: inst = 32'h10a00000;
      102716: inst = 32'hca00012;
      102717: inst = 32'h24822800;
      102718: inst = 32'h10a00000;
      102719: inst = 32'hca00004;
      102720: inst = 32'h38632800;
      102721: inst = 32'h38842800;
      102722: inst = 32'h10a00001;
      102723: inst = 32'hca09147;
      102724: inst = 32'h13e00001;
      102725: inst = 32'hfe0d96a;
      102726: inst = 32'h5be00000;
      102727: inst = 32'h8c50000;
      102728: inst = 32'h24612800;
      102729: inst = 32'h10a00000;
      102730: inst = 32'hca00012;
      102731: inst = 32'h24822800;
      102732: inst = 32'h10a00000;
      102733: inst = 32'hca00004;
      102734: inst = 32'h38632800;
      102735: inst = 32'h38842800;
      102736: inst = 32'h10a00001;
      102737: inst = 32'hca09155;
      102738: inst = 32'h13e00001;
      102739: inst = 32'hfe0d96a;
      102740: inst = 32'h5be00000;
      102741: inst = 32'h8c50000;
      102742: inst = 32'h24612800;
      102743: inst = 32'h10a00000;
      102744: inst = 32'hca00012;
      102745: inst = 32'h24822800;
      102746: inst = 32'h10a00000;
      102747: inst = 32'hca00004;
      102748: inst = 32'h38632800;
      102749: inst = 32'h38842800;
      102750: inst = 32'h10a00001;
      102751: inst = 32'hca09163;
      102752: inst = 32'h13e00001;
      102753: inst = 32'hfe0d96a;
      102754: inst = 32'h5be00000;
      102755: inst = 32'h8c50000;
      102756: inst = 32'h24612800;
      102757: inst = 32'h10a00000;
      102758: inst = 32'hca00012;
      102759: inst = 32'h24822800;
      102760: inst = 32'h10a00000;
      102761: inst = 32'hca00004;
      102762: inst = 32'h38632800;
      102763: inst = 32'h38842800;
      102764: inst = 32'h10a00001;
      102765: inst = 32'hca09171;
      102766: inst = 32'h13e00001;
      102767: inst = 32'hfe0d96a;
      102768: inst = 32'h5be00000;
      102769: inst = 32'h8c50000;
      102770: inst = 32'h24612800;
      102771: inst = 32'h10a00000;
      102772: inst = 32'hca00012;
      102773: inst = 32'h24822800;
      102774: inst = 32'h10a00000;
      102775: inst = 32'hca00004;
      102776: inst = 32'h38632800;
      102777: inst = 32'h38842800;
      102778: inst = 32'h10a00001;
      102779: inst = 32'hca0917f;
      102780: inst = 32'h13e00001;
      102781: inst = 32'hfe0d96a;
      102782: inst = 32'h5be00000;
      102783: inst = 32'h8c50000;
      102784: inst = 32'h24612800;
      102785: inst = 32'h10a00000;
      102786: inst = 32'hca00012;
      102787: inst = 32'h24822800;
      102788: inst = 32'h10a00000;
      102789: inst = 32'hca00004;
      102790: inst = 32'h38632800;
      102791: inst = 32'h38842800;
      102792: inst = 32'h10a00001;
      102793: inst = 32'hca0918d;
      102794: inst = 32'h13e00001;
      102795: inst = 32'hfe0d96a;
      102796: inst = 32'h5be00000;
      102797: inst = 32'h8c50000;
      102798: inst = 32'h24612800;
      102799: inst = 32'h10a00000;
      102800: inst = 32'hca00012;
      102801: inst = 32'h24822800;
      102802: inst = 32'h10a00000;
      102803: inst = 32'hca00004;
      102804: inst = 32'h38632800;
      102805: inst = 32'h38842800;
      102806: inst = 32'h10a00001;
      102807: inst = 32'hca0919b;
      102808: inst = 32'h13e00001;
      102809: inst = 32'hfe0d96a;
      102810: inst = 32'h5be00000;
      102811: inst = 32'h8c50000;
      102812: inst = 32'h24612800;
      102813: inst = 32'h10a00000;
      102814: inst = 32'hca00012;
      102815: inst = 32'h24822800;
      102816: inst = 32'h10a00000;
      102817: inst = 32'hca00004;
      102818: inst = 32'h38632800;
      102819: inst = 32'h38842800;
      102820: inst = 32'h10a00001;
      102821: inst = 32'hca091a9;
      102822: inst = 32'h13e00001;
      102823: inst = 32'hfe0d96a;
      102824: inst = 32'h5be00000;
      102825: inst = 32'h8c50000;
      102826: inst = 32'h24612800;
      102827: inst = 32'h10a00000;
      102828: inst = 32'hca00012;
      102829: inst = 32'h24822800;
      102830: inst = 32'h10a00000;
      102831: inst = 32'hca00004;
      102832: inst = 32'h38632800;
      102833: inst = 32'h38842800;
      102834: inst = 32'h10a00001;
      102835: inst = 32'hca091b7;
      102836: inst = 32'h13e00001;
      102837: inst = 32'hfe0d96a;
      102838: inst = 32'h5be00000;
      102839: inst = 32'h8c50000;
      102840: inst = 32'h24612800;
      102841: inst = 32'h10a00000;
      102842: inst = 32'hca00012;
      102843: inst = 32'h24822800;
      102844: inst = 32'h10a00000;
      102845: inst = 32'hca00004;
      102846: inst = 32'h38632800;
      102847: inst = 32'h38842800;
      102848: inst = 32'h10a00001;
      102849: inst = 32'hca091c5;
      102850: inst = 32'h13e00001;
      102851: inst = 32'hfe0d96a;
      102852: inst = 32'h5be00000;
      102853: inst = 32'h8c50000;
      102854: inst = 32'h24612800;
      102855: inst = 32'h10a00000;
      102856: inst = 32'hca00012;
      102857: inst = 32'h24822800;
      102858: inst = 32'h10a00000;
      102859: inst = 32'hca00004;
      102860: inst = 32'h38632800;
      102861: inst = 32'h38842800;
      102862: inst = 32'h10a00001;
      102863: inst = 32'hca091d3;
      102864: inst = 32'h13e00001;
      102865: inst = 32'hfe0d96a;
      102866: inst = 32'h5be00000;
      102867: inst = 32'h8c50000;
      102868: inst = 32'h24612800;
      102869: inst = 32'h10a00000;
      102870: inst = 32'hca00012;
      102871: inst = 32'h24822800;
      102872: inst = 32'h10a00000;
      102873: inst = 32'hca00004;
      102874: inst = 32'h38632800;
      102875: inst = 32'h38842800;
      102876: inst = 32'h10a00001;
      102877: inst = 32'hca091e1;
      102878: inst = 32'h13e00001;
      102879: inst = 32'hfe0d96a;
      102880: inst = 32'h5be00000;
      102881: inst = 32'h8c50000;
      102882: inst = 32'h24612800;
      102883: inst = 32'h10a00000;
      102884: inst = 32'hca00012;
      102885: inst = 32'h24822800;
      102886: inst = 32'h10a00000;
      102887: inst = 32'hca00004;
      102888: inst = 32'h38632800;
      102889: inst = 32'h38842800;
      102890: inst = 32'h10a00001;
      102891: inst = 32'hca091ef;
      102892: inst = 32'h13e00001;
      102893: inst = 32'hfe0d96a;
      102894: inst = 32'h5be00000;
      102895: inst = 32'h8c50000;
      102896: inst = 32'h24612800;
      102897: inst = 32'h10a00000;
      102898: inst = 32'hca00012;
      102899: inst = 32'h24822800;
      102900: inst = 32'h10a00000;
      102901: inst = 32'hca00004;
      102902: inst = 32'h38632800;
      102903: inst = 32'h38842800;
      102904: inst = 32'h10a00001;
      102905: inst = 32'hca091fd;
      102906: inst = 32'h13e00001;
      102907: inst = 32'hfe0d96a;
      102908: inst = 32'h5be00000;
      102909: inst = 32'h8c50000;
      102910: inst = 32'h24612800;
      102911: inst = 32'h10a00000;
      102912: inst = 32'hca00012;
      102913: inst = 32'h24822800;
      102914: inst = 32'h10a00000;
      102915: inst = 32'hca00004;
      102916: inst = 32'h38632800;
      102917: inst = 32'h38842800;
      102918: inst = 32'h10a00001;
      102919: inst = 32'hca0920b;
      102920: inst = 32'h13e00001;
      102921: inst = 32'hfe0d96a;
      102922: inst = 32'h5be00000;
      102923: inst = 32'h8c50000;
      102924: inst = 32'h24612800;
      102925: inst = 32'h10a00000;
      102926: inst = 32'hca00012;
      102927: inst = 32'h24822800;
      102928: inst = 32'h10a00000;
      102929: inst = 32'hca00004;
      102930: inst = 32'h38632800;
      102931: inst = 32'h38842800;
      102932: inst = 32'h10a00001;
      102933: inst = 32'hca09219;
      102934: inst = 32'h13e00001;
      102935: inst = 32'hfe0d96a;
      102936: inst = 32'h5be00000;
      102937: inst = 32'h8c50000;
      102938: inst = 32'h24612800;
      102939: inst = 32'h10a00000;
      102940: inst = 32'hca00012;
      102941: inst = 32'h24822800;
      102942: inst = 32'h10a00000;
      102943: inst = 32'hca00004;
      102944: inst = 32'h38632800;
      102945: inst = 32'h38842800;
      102946: inst = 32'h10a00001;
      102947: inst = 32'hca09227;
      102948: inst = 32'h13e00001;
      102949: inst = 32'hfe0d96a;
      102950: inst = 32'h5be00000;
      102951: inst = 32'h8c50000;
      102952: inst = 32'h24612800;
      102953: inst = 32'h10a00000;
      102954: inst = 32'hca00012;
      102955: inst = 32'h24822800;
      102956: inst = 32'h10a00000;
      102957: inst = 32'hca00004;
      102958: inst = 32'h38632800;
      102959: inst = 32'h38842800;
      102960: inst = 32'h10a00001;
      102961: inst = 32'hca09235;
      102962: inst = 32'h13e00001;
      102963: inst = 32'hfe0d96a;
      102964: inst = 32'h5be00000;
      102965: inst = 32'h8c50000;
      102966: inst = 32'h24612800;
      102967: inst = 32'h10a00000;
      102968: inst = 32'hca00012;
      102969: inst = 32'h24822800;
      102970: inst = 32'h10a00000;
      102971: inst = 32'hca00004;
      102972: inst = 32'h38632800;
      102973: inst = 32'h38842800;
      102974: inst = 32'h10a00001;
      102975: inst = 32'hca09243;
      102976: inst = 32'h13e00001;
      102977: inst = 32'hfe0d96a;
      102978: inst = 32'h5be00000;
      102979: inst = 32'h8c50000;
      102980: inst = 32'h24612800;
      102981: inst = 32'h10a00000;
      102982: inst = 32'hca00012;
      102983: inst = 32'h24822800;
      102984: inst = 32'h10a00000;
      102985: inst = 32'hca00004;
      102986: inst = 32'h38632800;
      102987: inst = 32'h38842800;
      102988: inst = 32'h10a00001;
      102989: inst = 32'hca09251;
      102990: inst = 32'h13e00001;
      102991: inst = 32'hfe0d96a;
      102992: inst = 32'h5be00000;
      102993: inst = 32'h8c50000;
      102994: inst = 32'h24612800;
      102995: inst = 32'h10a00000;
      102996: inst = 32'hca00012;
      102997: inst = 32'h24822800;
      102998: inst = 32'h10a00000;
      102999: inst = 32'hca00004;
      103000: inst = 32'h38632800;
      103001: inst = 32'h38842800;
      103002: inst = 32'h10a00001;
      103003: inst = 32'hca0925f;
      103004: inst = 32'h13e00001;
      103005: inst = 32'hfe0d96a;
      103006: inst = 32'h5be00000;
      103007: inst = 32'h8c50000;
      103008: inst = 32'h24612800;
      103009: inst = 32'h10a00000;
      103010: inst = 32'hca00012;
      103011: inst = 32'h24822800;
      103012: inst = 32'h10a00000;
      103013: inst = 32'hca00004;
      103014: inst = 32'h38632800;
      103015: inst = 32'h38842800;
      103016: inst = 32'h10a00001;
      103017: inst = 32'hca0926d;
      103018: inst = 32'h13e00001;
      103019: inst = 32'hfe0d96a;
      103020: inst = 32'h5be00000;
      103021: inst = 32'h8c50000;
      103022: inst = 32'h24612800;
      103023: inst = 32'h10a00000;
      103024: inst = 32'hca00012;
      103025: inst = 32'h24822800;
      103026: inst = 32'h10a00000;
      103027: inst = 32'hca00004;
      103028: inst = 32'h38632800;
      103029: inst = 32'h38842800;
      103030: inst = 32'h10a00001;
      103031: inst = 32'hca0927b;
      103032: inst = 32'h13e00001;
      103033: inst = 32'hfe0d96a;
      103034: inst = 32'h5be00000;
      103035: inst = 32'h8c50000;
      103036: inst = 32'h24612800;
      103037: inst = 32'h10a00000;
      103038: inst = 32'hca00012;
      103039: inst = 32'h24822800;
      103040: inst = 32'h10a00000;
      103041: inst = 32'hca00004;
      103042: inst = 32'h38632800;
      103043: inst = 32'h38842800;
      103044: inst = 32'h10a00001;
      103045: inst = 32'hca09289;
      103046: inst = 32'h13e00001;
      103047: inst = 32'hfe0d96a;
      103048: inst = 32'h5be00000;
      103049: inst = 32'h8c50000;
      103050: inst = 32'h24612800;
      103051: inst = 32'h10a00000;
      103052: inst = 32'hca00012;
      103053: inst = 32'h24822800;
      103054: inst = 32'h10a00000;
      103055: inst = 32'hca00004;
      103056: inst = 32'h38632800;
      103057: inst = 32'h38842800;
      103058: inst = 32'h10a00001;
      103059: inst = 32'hca09297;
      103060: inst = 32'h13e00001;
      103061: inst = 32'hfe0d96a;
      103062: inst = 32'h5be00000;
      103063: inst = 32'h8c50000;
      103064: inst = 32'h24612800;
      103065: inst = 32'h10a00000;
      103066: inst = 32'hca00012;
      103067: inst = 32'h24822800;
      103068: inst = 32'h10a00000;
      103069: inst = 32'hca00004;
      103070: inst = 32'h38632800;
      103071: inst = 32'h38842800;
      103072: inst = 32'h10a00001;
      103073: inst = 32'hca092a5;
      103074: inst = 32'h13e00001;
      103075: inst = 32'hfe0d96a;
      103076: inst = 32'h5be00000;
      103077: inst = 32'h8c50000;
      103078: inst = 32'h24612800;
      103079: inst = 32'h10a00000;
      103080: inst = 32'hca00012;
      103081: inst = 32'h24822800;
      103082: inst = 32'h10a00000;
      103083: inst = 32'hca00004;
      103084: inst = 32'h38632800;
      103085: inst = 32'h38842800;
      103086: inst = 32'h10a00001;
      103087: inst = 32'hca092b3;
      103088: inst = 32'h13e00001;
      103089: inst = 32'hfe0d96a;
      103090: inst = 32'h5be00000;
      103091: inst = 32'h8c50000;
      103092: inst = 32'h24612800;
      103093: inst = 32'h10a00000;
      103094: inst = 32'hca00012;
      103095: inst = 32'h24822800;
      103096: inst = 32'h10a00000;
      103097: inst = 32'hca00004;
      103098: inst = 32'h38632800;
      103099: inst = 32'h38842800;
      103100: inst = 32'h10a00001;
      103101: inst = 32'hca092c1;
      103102: inst = 32'h13e00001;
      103103: inst = 32'hfe0d96a;
      103104: inst = 32'h5be00000;
      103105: inst = 32'h8c50000;
      103106: inst = 32'h24612800;
      103107: inst = 32'h10a00000;
      103108: inst = 32'hca00012;
      103109: inst = 32'h24822800;
      103110: inst = 32'h10a00000;
      103111: inst = 32'hca00004;
      103112: inst = 32'h38632800;
      103113: inst = 32'h38842800;
      103114: inst = 32'h10a00001;
      103115: inst = 32'hca092cf;
      103116: inst = 32'h13e00001;
      103117: inst = 32'hfe0d96a;
      103118: inst = 32'h5be00000;
      103119: inst = 32'h8c50000;
      103120: inst = 32'h24612800;
      103121: inst = 32'h10a00000;
      103122: inst = 32'hca00012;
      103123: inst = 32'h24822800;
      103124: inst = 32'h10a00000;
      103125: inst = 32'hca00004;
      103126: inst = 32'h38632800;
      103127: inst = 32'h38842800;
      103128: inst = 32'h10a00001;
      103129: inst = 32'hca092dd;
      103130: inst = 32'h13e00001;
      103131: inst = 32'hfe0d96a;
      103132: inst = 32'h5be00000;
      103133: inst = 32'h8c50000;
      103134: inst = 32'h24612800;
      103135: inst = 32'h10a00000;
      103136: inst = 32'hca00012;
      103137: inst = 32'h24822800;
      103138: inst = 32'h10a00000;
      103139: inst = 32'hca00004;
      103140: inst = 32'h38632800;
      103141: inst = 32'h38842800;
      103142: inst = 32'h10a00001;
      103143: inst = 32'hca092eb;
      103144: inst = 32'h13e00001;
      103145: inst = 32'hfe0d96a;
      103146: inst = 32'h5be00000;
      103147: inst = 32'h8c50000;
      103148: inst = 32'h24612800;
      103149: inst = 32'h10a00000;
      103150: inst = 32'hca00012;
      103151: inst = 32'h24822800;
      103152: inst = 32'h10a00000;
      103153: inst = 32'hca00004;
      103154: inst = 32'h38632800;
      103155: inst = 32'h38842800;
      103156: inst = 32'h10a00001;
      103157: inst = 32'hca092f9;
      103158: inst = 32'h13e00001;
      103159: inst = 32'hfe0d96a;
      103160: inst = 32'h5be00000;
      103161: inst = 32'h8c50000;
      103162: inst = 32'h24612800;
      103163: inst = 32'h10a00000;
      103164: inst = 32'hca00012;
      103165: inst = 32'h24822800;
      103166: inst = 32'h10a00000;
      103167: inst = 32'hca00004;
      103168: inst = 32'h38632800;
      103169: inst = 32'h38842800;
      103170: inst = 32'h10a00001;
      103171: inst = 32'hca09307;
      103172: inst = 32'h13e00001;
      103173: inst = 32'hfe0d96a;
      103174: inst = 32'h5be00000;
      103175: inst = 32'h8c50000;
      103176: inst = 32'h24612800;
      103177: inst = 32'h10a00000;
      103178: inst = 32'hca00012;
      103179: inst = 32'h24822800;
      103180: inst = 32'h10a00000;
      103181: inst = 32'hca00004;
      103182: inst = 32'h38632800;
      103183: inst = 32'h38842800;
      103184: inst = 32'h10a00001;
      103185: inst = 32'hca09315;
      103186: inst = 32'h13e00001;
      103187: inst = 32'hfe0d96a;
      103188: inst = 32'h5be00000;
      103189: inst = 32'h8c50000;
      103190: inst = 32'h24612800;
      103191: inst = 32'h10a00000;
      103192: inst = 32'hca00012;
      103193: inst = 32'h24822800;
      103194: inst = 32'h10a00000;
      103195: inst = 32'hca00004;
      103196: inst = 32'h38632800;
      103197: inst = 32'h38842800;
      103198: inst = 32'h10a00001;
      103199: inst = 32'hca09323;
      103200: inst = 32'h13e00001;
      103201: inst = 32'hfe0d96a;
      103202: inst = 32'h5be00000;
      103203: inst = 32'h8c50000;
      103204: inst = 32'h24612800;
      103205: inst = 32'h10a00000;
      103206: inst = 32'hca00012;
      103207: inst = 32'h24822800;
      103208: inst = 32'h10a00000;
      103209: inst = 32'hca00004;
      103210: inst = 32'h38632800;
      103211: inst = 32'h38842800;
      103212: inst = 32'h10a00001;
      103213: inst = 32'hca09331;
      103214: inst = 32'h13e00001;
      103215: inst = 32'hfe0d96a;
      103216: inst = 32'h5be00000;
      103217: inst = 32'h8c50000;
      103218: inst = 32'h24612800;
      103219: inst = 32'h10a00000;
      103220: inst = 32'hca00012;
      103221: inst = 32'h24822800;
      103222: inst = 32'h10a00000;
      103223: inst = 32'hca00004;
      103224: inst = 32'h38632800;
      103225: inst = 32'h38842800;
      103226: inst = 32'h10a00001;
      103227: inst = 32'hca0933f;
      103228: inst = 32'h13e00001;
      103229: inst = 32'hfe0d96a;
      103230: inst = 32'h5be00000;
      103231: inst = 32'h8c50000;
      103232: inst = 32'h24612800;
      103233: inst = 32'h10a00000;
      103234: inst = 32'hca00012;
      103235: inst = 32'h24822800;
      103236: inst = 32'h10a00000;
      103237: inst = 32'hca00004;
      103238: inst = 32'h38632800;
      103239: inst = 32'h38842800;
      103240: inst = 32'h10a00001;
      103241: inst = 32'hca0934d;
      103242: inst = 32'h13e00001;
      103243: inst = 32'hfe0d96a;
      103244: inst = 32'h5be00000;
      103245: inst = 32'h8c50000;
      103246: inst = 32'h24612800;
      103247: inst = 32'h10a00000;
      103248: inst = 32'hca00012;
      103249: inst = 32'h24822800;
      103250: inst = 32'h10a00000;
      103251: inst = 32'hca00004;
      103252: inst = 32'h38632800;
      103253: inst = 32'h38842800;
      103254: inst = 32'h10a00001;
      103255: inst = 32'hca0935b;
      103256: inst = 32'h13e00001;
      103257: inst = 32'hfe0d96a;
      103258: inst = 32'h5be00000;
      103259: inst = 32'h8c50000;
      103260: inst = 32'h24612800;
      103261: inst = 32'h10a00000;
      103262: inst = 32'hca00012;
      103263: inst = 32'h24822800;
      103264: inst = 32'h10a00000;
      103265: inst = 32'hca00004;
      103266: inst = 32'h38632800;
      103267: inst = 32'h38842800;
      103268: inst = 32'h10a00001;
      103269: inst = 32'hca09369;
      103270: inst = 32'h13e00001;
      103271: inst = 32'hfe0d96a;
      103272: inst = 32'h5be00000;
      103273: inst = 32'h8c50000;
      103274: inst = 32'h24612800;
      103275: inst = 32'h10a00000;
      103276: inst = 32'hca00012;
      103277: inst = 32'h24822800;
      103278: inst = 32'h10a00000;
      103279: inst = 32'hca00004;
      103280: inst = 32'h38632800;
      103281: inst = 32'h38842800;
      103282: inst = 32'h10a00001;
      103283: inst = 32'hca09377;
      103284: inst = 32'h13e00001;
      103285: inst = 32'hfe0d96a;
      103286: inst = 32'h5be00000;
      103287: inst = 32'h8c50000;
      103288: inst = 32'h24612800;
      103289: inst = 32'h10a00000;
      103290: inst = 32'hca00012;
      103291: inst = 32'h24822800;
      103292: inst = 32'h10a00000;
      103293: inst = 32'hca00004;
      103294: inst = 32'h38632800;
      103295: inst = 32'h38842800;
      103296: inst = 32'h10a00001;
      103297: inst = 32'hca09385;
      103298: inst = 32'h13e00001;
      103299: inst = 32'hfe0d96a;
      103300: inst = 32'h5be00000;
      103301: inst = 32'h8c50000;
      103302: inst = 32'h24612800;
      103303: inst = 32'h10a00000;
      103304: inst = 32'hca00012;
      103305: inst = 32'h24822800;
      103306: inst = 32'h10a00000;
      103307: inst = 32'hca00004;
      103308: inst = 32'h38632800;
      103309: inst = 32'h38842800;
      103310: inst = 32'h10a00001;
      103311: inst = 32'hca09393;
      103312: inst = 32'h13e00001;
      103313: inst = 32'hfe0d96a;
      103314: inst = 32'h5be00000;
      103315: inst = 32'h8c50000;
      103316: inst = 32'h24612800;
      103317: inst = 32'h10a00000;
      103318: inst = 32'hca00012;
      103319: inst = 32'h24822800;
      103320: inst = 32'h10a00000;
      103321: inst = 32'hca00004;
      103322: inst = 32'h38632800;
      103323: inst = 32'h38842800;
      103324: inst = 32'h10a00001;
      103325: inst = 32'hca093a1;
      103326: inst = 32'h13e00001;
      103327: inst = 32'hfe0d96a;
      103328: inst = 32'h5be00000;
      103329: inst = 32'h8c50000;
      103330: inst = 32'h24612800;
      103331: inst = 32'h10a00000;
      103332: inst = 32'hca00012;
      103333: inst = 32'h24822800;
      103334: inst = 32'h10a00000;
      103335: inst = 32'hca00004;
      103336: inst = 32'h38632800;
      103337: inst = 32'h38842800;
      103338: inst = 32'h10a00001;
      103339: inst = 32'hca093af;
      103340: inst = 32'h13e00001;
      103341: inst = 32'hfe0d96a;
      103342: inst = 32'h5be00000;
      103343: inst = 32'h8c50000;
      103344: inst = 32'h24612800;
      103345: inst = 32'h10a00000;
      103346: inst = 32'hca00012;
      103347: inst = 32'h24822800;
      103348: inst = 32'h10a00000;
      103349: inst = 32'hca00004;
      103350: inst = 32'h38632800;
      103351: inst = 32'h38842800;
      103352: inst = 32'h10a00001;
      103353: inst = 32'hca093bd;
      103354: inst = 32'h13e00001;
      103355: inst = 32'hfe0d96a;
      103356: inst = 32'h5be00000;
      103357: inst = 32'h8c50000;
      103358: inst = 32'h24612800;
      103359: inst = 32'h10a00000;
      103360: inst = 32'hca00012;
      103361: inst = 32'h24822800;
      103362: inst = 32'h10a00000;
      103363: inst = 32'hca00004;
      103364: inst = 32'h38632800;
      103365: inst = 32'h38842800;
      103366: inst = 32'h10a00001;
      103367: inst = 32'hca093cb;
      103368: inst = 32'h13e00001;
      103369: inst = 32'hfe0d96a;
      103370: inst = 32'h5be00000;
      103371: inst = 32'h8c50000;
      103372: inst = 32'h24612800;
      103373: inst = 32'h10a00000;
      103374: inst = 32'hca00012;
      103375: inst = 32'h24822800;
      103376: inst = 32'h10a00000;
      103377: inst = 32'hca00004;
      103378: inst = 32'h38632800;
      103379: inst = 32'h38842800;
      103380: inst = 32'h10a00001;
      103381: inst = 32'hca093d9;
      103382: inst = 32'h13e00001;
      103383: inst = 32'hfe0d96a;
      103384: inst = 32'h5be00000;
      103385: inst = 32'h8c50000;
      103386: inst = 32'h24612800;
      103387: inst = 32'h10a00000;
      103388: inst = 32'hca00012;
      103389: inst = 32'h24822800;
      103390: inst = 32'h10a00000;
      103391: inst = 32'hca00004;
      103392: inst = 32'h38632800;
      103393: inst = 32'h38842800;
      103394: inst = 32'h10a00001;
      103395: inst = 32'hca093e7;
      103396: inst = 32'h13e00001;
      103397: inst = 32'hfe0d96a;
      103398: inst = 32'h5be00000;
      103399: inst = 32'h8c50000;
      103400: inst = 32'h24612800;
      103401: inst = 32'h10a00000;
      103402: inst = 32'hca00012;
      103403: inst = 32'h24822800;
      103404: inst = 32'h10a00000;
      103405: inst = 32'hca00004;
      103406: inst = 32'h38632800;
      103407: inst = 32'h38842800;
      103408: inst = 32'h10a00001;
      103409: inst = 32'hca093f5;
      103410: inst = 32'h13e00001;
      103411: inst = 32'hfe0d96a;
      103412: inst = 32'h5be00000;
      103413: inst = 32'h8c50000;
      103414: inst = 32'h24612800;
      103415: inst = 32'h10a00000;
      103416: inst = 32'hca00012;
      103417: inst = 32'h24822800;
      103418: inst = 32'h10a00000;
      103419: inst = 32'hca00004;
      103420: inst = 32'h38632800;
      103421: inst = 32'h38842800;
      103422: inst = 32'h10a00001;
      103423: inst = 32'hca09403;
      103424: inst = 32'h13e00001;
      103425: inst = 32'hfe0d96a;
      103426: inst = 32'h5be00000;
      103427: inst = 32'h8c50000;
      103428: inst = 32'h24612800;
      103429: inst = 32'h10a00000;
      103430: inst = 32'hca00012;
      103431: inst = 32'h24822800;
      103432: inst = 32'h10a00000;
      103433: inst = 32'hca00004;
      103434: inst = 32'h38632800;
      103435: inst = 32'h38842800;
      103436: inst = 32'h10a00001;
      103437: inst = 32'hca09411;
      103438: inst = 32'h13e00001;
      103439: inst = 32'hfe0d96a;
      103440: inst = 32'h5be00000;
      103441: inst = 32'h8c50000;
      103442: inst = 32'h24612800;
      103443: inst = 32'h10a00000;
      103444: inst = 32'hca00012;
      103445: inst = 32'h24822800;
      103446: inst = 32'h10a00000;
      103447: inst = 32'hca00004;
      103448: inst = 32'h38632800;
      103449: inst = 32'h38842800;
      103450: inst = 32'h10a00001;
      103451: inst = 32'hca0941f;
      103452: inst = 32'h13e00001;
      103453: inst = 32'hfe0d96a;
      103454: inst = 32'h5be00000;
      103455: inst = 32'h8c50000;
      103456: inst = 32'h24612800;
      103457: inst = 32'h10a00000;
      103458: inst = 32'hca00012;
      103459: inst = 32'h24822800;
      103460: inst = 32'h10a00000;
      103461: inst = 32'hca00004;
      103462: inst = 32'h38632800;
      103463: inst = 32'h38842800;
      103464: inst = 32'h10a00001;
      103465: inst = 32'hca0942d;
      103466: inst = 32'h13e00001;
      103467: inst = 32'hfe0d96a;
      103468: inst = 32'h5be00000;
      103469: inst = 32'h8c50000;
      103470: inst = 32'h24612800;
      103471: inst = 32'h10a00000;
      103472: inst = 32'hca00012;
      103473: inst = 32'h24822800;
      103474: inst = 32'h10a00000;
      103475: inst = 32'hca00004;
      103476: inst = 32'h38632800;
      103477: inst = 32'h38842800;
      103478: inst = 32'h10a00001;
      103479: inst = 32'hca0943b;
      103480: inst = 32'h13e00001;
      103481: inst = 32'hfe0d96a;
      103482: inst = 32'h5be00000;
      103483: inst = 32'h8c50000;
      103484: inst = 32'h24612800;
      103485: inst = 32'h10a00000;
      103486: inst = 32'hca00012;
      103487: inst = 32'h24822800;
      103488: inst = 32'h10a00000;
      103489: inst = 32'hca00004;
      103490: inst = 32'h38632800;
      103491: inst = 32'h38842800;
      103492: inst = 32'h10a00001;
      103493: inst = 32'hca09449;
      103494: inst = 32'h13e00001;
      103495: inst = 32'hfe0d96a;
      103496: inst = 32'h5be00000;
      103497: inst = 32'h8c50000;
      103498: inst = 32'h24612800;
      103499: inst = 32'h10a00000;
      103500: inst = 32'hca00012;
      103501: inst = 32'h24822800;
      103502: inst = 32'h10a00000;
      103503: inst = 32'hca00004;
      103504: inst = 32'h38632800;
      103505: inst = 32'h38842800;
      103506: inst = 32'h10a00001;
      103507: inst = 32'hca09457;
      103508: inst = 32'h13e00001;
      103509: inst = 32'hfe0d96a;
      103510: inst = 32'h5be00000;
      103511: inst = 32'h8c50000;
      103512: inst = 32'h24612800;
      103513: inst = 32'h10a00000;
      103514: inst = 32'hca00012;
      103515: inst = 32'h24822800;
      103516: inst = 32'h10a00000;
      103517: inst = 32'hca00004;
      103518: inst = 32'h38632800;
      103519: inst = 32'h38842800;
      103520: inst = 32'h10a00001;
      103521: inst = 32'hca09465;
      103522: inst = 32'h13e00001;
      103523: inst = 32'hfe0d96a;
      103524: inst = 32'h5be00000;
      103525: inst = 32'h8c50000;
      103526: inst = 32'h24612800;
      103527: inst = 32'h10a00000;
      103528: inst = 32'hca00012;
      103529: inst = 32'h24822800;
      103530: inst = 32'h10a00000;
      103531: inst = 32'hca00004;
      103532: inst = 32'h38632800;
      103533: inst = 32'h38842800;
      103534: inst = 32'h10a00001;
      103535: inst = 32'hca09473;
      103536: inst = 32'h13e00001;
      103537: inst = 32'hfe0d96a;
      103538: inst = 32'h5be00000;
      103539: inst = 32'h8c50000;
      103540: inst = 32'h24612800;
      103541: inst = 32'h10a00000;
      103542: inst = 32'hca00012;
      103543: inst = 32'h24822800;
      103544: inst = 32'h10a00000;
      103545: inst = 32'hca00004;
      103546: inst = 32'h38632800;
      103547: inst = 32'h38842800;
      103548: inst = 32'h10a00001;
      103549: inst = 32'hca09481;
      103550: inst = 32'h13e00001;
      103551: inst = 32'hfe0d96a;
      103552: inst = 32'h5be00000;
      103553: inst = 32'h8c50000;
      103554: inst = 32'h24612800;
      103555: inst = 32'h10a00000;
      103556: inst = 32'hca00012;
      103557: inst = 32'h24822800;
      103558: inst = 32'h10a00000;
      103559: inst = 32'hca00004;
      103560: inst = 32'h38632800;
      103561: inst = 32'h38842800;
      103562: inst = 32'h10a00001;
      103563: inst = 32'hca0948f;
      103564: inst = 32'h13e00001;
      103565: inst = 32'hfe0d96a;
      103566: inst = 32'h5be00000;
      103567: inst = 32'h8c50000;
      103568: inst = 32'h24612800;
      103569: inst = 32'h10a00000;
      103570: inst = 32'hca00012;
      103571: inst = 32'h24822800;
      103572: inst = 32'h10a00000;
      103573: inst = 32'hca00004;
      103574: inst = 32'h38632800;
      103575: inst = 32'h38842800;
      103576: inst = 32'h10a00001;
      103577: inst = 32'hca0949d;
      103578: inst = 32'h13e00001;
      103579: inst = 32'hfe0d96a;
      103580: inst = 32'h5be00000;
      103581: inst = 32'h8c50000;
      103582: inst = 32'h24612800;
      103583: inst = 32'h10a00000;
      103584: inst = 32'hca00012;
      103585: inst = 32'h24822800;
      103586: inst = 32'h10a00000;
      103587: inst = 32'hca00004;
      103588: inst = 32'h38632800;
      103589: inst = 32'h38842800;
      103590: inst = 32'h10a00001;
      103591: inst = 32'hca094ab;
      103592: inst = 32'h13e00001;
      103593: inst = 32'hfe0d96a;
      103594: inst = 32'h5be00000;
      103595: inst = 32'h8c50000;
      103596: inst = 32'h24612800;
      103597: inst = 32'h10a00000;
      103598: inst = 32'hca00012;
      103599: inst = 32'h24822800;
      103600: inst = 32'h10a00000;
      103601: inst = 32'hca00004;
      103602: inst = 32'h38632800;
      103603: inst = 32'h38842800;
      103604: inst = 32'h10a00001;
      103605: inst = 32'hca094b9;
      103606: inst = 32'h13e00001;
      103607: inst = 32'hfe0d96a;
      103608: inst = 32'h5be00000;
      103609: inst = 32'h8c50000;
      103610: inst = 32'h24612800;
      103611: inst = 32'h10a00000;
      103612: inst = 32'hca00012;
      103613: inst = 32'h24822800;
      103614: inst = 32'h10a00000;
      103615: inst = 32'hca00004;
      103616: inst = 32'h38632800;
      103617: inst = 32'h38842800;
      103618: inst = 32'h10a00001;
      103619: inst = 32'hca094c7;
      103620: inst = 32'h13e00001;
      103621: inst = 32'hfe0d96a;
      103622: inst = 32'h5be00000;
      103623: inst = 32'h8c50000;
      103624: inst = 32'h24612800;
      103625: inst = 32'h10a00000;
      103626: inst = 32'hca00012;
      103627: inst = 32'h24822800;
      103628: inst = 32'h10a00000;
      103629: inst = 32'hca00004;
      103630: inst = 32'h38632800;
      103631: inst = 32'h38842800;
      103632: inst = 32'h10a00001;
      103633: inst = 32'hca094d5;
      103634: inst = 32'h13e00001;
      103635: inst = 32'hfe0d96a;
      103636: inst = 32'h5be00000;
      103637: inst = 32'h8c50000;
      103638: inst = 32'h24612800;
      103639: inst = 32'h10a00000;
      103640: inst = 32'hca00012;
      103641: inst = 32'h24822800;
      103642: inst = 32'h10a00000;
      103643: inst = 32'hca00004;
      103644: inst = 32'h38632800;
      103645: inst = 32'h38842800;
      103646: inst = 32'h10a00001;
      103647: inst = 32'hca094e3;
      103648: inst = 32'h13e00001;
      103649: inst = 32'hfe0d96a;
      103650: inst = 32'h5be00000;
      103651: inst = 32'h8c50000;
      103652: inst = 32'h24612800;
      103653: inst = 32'h10a00000;
      103654: inst = 32'hca00012;
      103655: inst = 32'h24822800;
      103656: inst = 32'h10a00000;
      103657: inst = 32'hca00004;
      103658: inst = 32'h38632800;
      103659: inst = 32'h38842800;
      103660: inst = 32'h10a00001;
      103661: inst = 32'hca094f1;
      103662: inst = 32'h13e00001;
      103663: inst = 32'hfe0d96a;
      103664: inst = 32'h5be00000;
      103665: inst = 32'h8c50000;
      103666: inst = 32'h24612800;
      103667: inst = 32'h10a00000;
      103668: inst = 32'hca00012;
      103669: inst = 32'h24822800;
      103670: inst = 32'h10a00000;
      103671: inst = 32'hca00004;
      103672: inst = 32'h38632800;
      103673: inst = 32'h38842800;
      103674: inst = 32'h10a00001;
      103675: inst = 32'hca094ff;
      103676: inst = 32'h13e00001;
      103677: inst = 32'hfe0d96a;
      103678: inst = 32'h5be00000;
      103679: inst = 32'h8c50000;
      103680: inst = 32'h24612800;
      103681: inst = 32'h10a00000;
      103682: inst = 32'hca00012;
      103683: inst = 32'h24822800;
      103684: inst = 32'h10a00000;
      103685: inst = 32'hca00004;
      103686: inst = 32'h38632800;
      103687: inst = 32'h38842800;
      103688: inst = 32'h10a00001;
      103689: inst = 32'hca0950d;
      103690: inst = 32'h13e00001;
      103691: inst = 32'hfe0d96a;
      103692: inst = 32'h5be00000;
      103693: inst = 32'h8c50000;
      103694: inst = 32'h24612800;
      103695: inst = 32'h10a00000;
      103696: inst = 32'hca00012;
      103697: inst = 32'h24822800;
      103698: inst = 32'h10a00000;
      103699: inst = 32'hca00004;
      103700: inst = 32'h38632800;
      103701: inst = 32'h38842800;
      103702: inst = 32'h10a00001;
      103703: inst = 32'hca0951b;
      103704: inst = 32'h13e00001;
      103705: inst = 32'hfe0d96a;
      103706: inst = 32'h5be00000;
      103707: inst = 32'h8c50000;
      103708: inst = 32'h24612800;
      103709: inst = 32'h10a00000;
      103710: inst = 32'hca00012;
      103711: inst = 32'h24822800;
      103712: inst = 32'h10a00000;
      103713: inst = 32'hca00004;
      103714: inst = 32'h38632800;
      103715: inst = 32'h38842800;
      103716: inst = 32'h10a00001;
      103717: inst = 32'hca09529;
      103718: inst = 32'h13e00001;
      103719: inst = 32'hfe0d96a;
      103720: inst = 32'h5be00000;
      103721: inst = 32'h8c50000;
      103722: inst = 32'h24612800;
      103723: inst = 32'h10a00000;
      103724: inst = 32'hca00013;
      103725: inst = 32'h24822800;
      103726: inst = 32'h10a00000;
      103727: inst = 32'hca00004;
      103728: inst = 32'h38632800;
      103729: inst = 32'h38842800;
      103730: inst = 32'h10a00001;
      103731: inst = 32'hca09537;
      103732: inst = 32'h13e00001;
      103733: inst = 32'hfe0d96a;
      103734: inst = 32'h5be00000;
      103735: inst = 32'h8c50000;
      103736: inst = 32'h24612800;
      103737: inst = 32'h10a00000;
      103738: inst = 32'hca00013;
      103739: inst = 32'h24822800;
      103740: inst = 32'h10a00000;
      103741: inst = 32'hca00004;
      103742: inst = 32'h38632800;
      103743: inst = 32'h38842800;
      103744: inst = 32'h10a00001;
      103745: inst = 32'hca09545;
      103746: inst = 32'h13e00001;
      103747: inst = 32'hfe0d96a;
      103748: inst = 32'h5be00000;
      103749: inst = 32'h8c50000;
      103750: inst = 32'h24612800;
      103751: inst = 32'h10a00000;
      103752: inst = 32'hca00013;
      103753: inst = 32'h24822800;
      103754: inst = 32'h10a00000;
      103755: inst = 32'hca00004;
      103756: inst = 32'h38632800;
      103757: inst = 32'h38842800;
      103758: inst = 32'h10a00001;
      103759: inst = 32'hca09553;
      103760: inst = 32'h13e00001;
      103761: inst = 32'hfe0d96a;
      103762: inst = 32'h5be00000;
      103763: inst = 32'h8c50000;
      103764: inst = 32'h24612800;
      103765: inst = 32'h10a00000;
      103766: inst = 32'hca00013;
      103767: inst = 32'h24822800;
      103768: inst = 32'h10a00000;
      103769: inst = 32'hca00004;
      103770: inst = 32'h38632800;
      103771: inst = 32'h38842800;
      103772: inst = 32'h10a00001;
      103773: inst = 32'hca09561;
      103774: inst = 32'h13e00001;
      103775: inst = 32'hfe0d96a;
      103776: inst = 32'h5be00000;
      103777: inst = 32'h8c50000;
      103778: inst = 32'h24612800;
      103779: inst = 32'h10a00000;
      103780: inst = 32'hca00013;
      103781: inst = 32'h24822800;
      103782: inst = 32'h10a00000;
      103783: inst = 32'hca00004;
      103784: inst = 32'h38632800;
      103785: inst = 32'h38842800;
      103786: inst = 32'h10a00001;
      103787: inst = 32'hca0956f;
      103788: inst = 32'h13e00001;
      103789: inst = 32'hfe0d96a;
      103790: inst = 32'h5be00000;
      103791: inst = 32'h8c50000;
      103792: inst = 32'h24612800;
      103793: inst = 32'h10a00000;
      103794: inst = 32'hca00013;
      103795: inst = 32'h24822800;
      103796: inst = 32'h10a00000;
      103797: inst = 32'hca00004;
      103798: inst = 32'h38632800;
      103799: inst = 32'h38842800;
      103800: inst = 32'h10a00001;
      103801: inst = 32'hca0957d;
      103802: inst = 32'h13e00001;
      103803: inst = 32'hfe0d96a;
      103804: inst = 32'h5be00000;
      103805: inst = 32'h8c50000;
      103806: inst = 32'h24612800;
      103807: inst = 32'h10a00000;
      103808: inst = 32'hca00013;
      103809: inst = 32'h24822800;
      103810: inst = 32'h10a00000;
      103811: inst = 32'hca00004;
      103812: inst = 32'h38632800;
      103813: inst = 32'h38842800;
      103814: inst = 32'h10a00001;
      103815: inst = 32'hca0958b;
      103816: inst = 32'h13e00001;
      103817: inst = 32'hfe0d96a;
      103818: inst = 32'h5be00000;
      103819: inst = 32'h8c50000;
      103820: inst = 32'h24612800;
      103821: inst = 32'h10a00000;
      103822: inst = 32'hca00013;
      103823: inst = 32'h24822800;
      103824: inst = 32'h10a00000;
      103825: inst = 32'hca00004;
      103826: inst = 32'h38632800;
      103827: inst = 32'h38842800;
      103828: inst = 32'h10a00001;
      103829: inst = 32'hca09599;
      103830: inst = 32'h13e00001;
      103831: inst = 32'hfe0d96a;
      103832: inst = 32'h5be00000;
      103833: inst = 32'h8c50000;
      103834: inst = 32'h24612800;
      103835: inst = 32'h10a00000;
      103836: inst = 32'hca00013;
      103837: inst = 32'h24822800;
      103838: inst = 32'h10a00000;
      103839: inst = 32'hca00004;
      103840: inst = 32'h38632800;
      103841: inst = 32'h38842800;
      103842: inst = 32'h10a00001;
      103843: inst = 32'hca095a7;
      103844: inst = 32'h13e00001;
      103845: inst = 32'hfe0d96a;
      103846: inst = 32'h5be00000;
      103847: inst = 32'h8c50000;
      103848: inst = 32'h24612800;
      103849: inst = 32'h10a00000;
      103850: inst = 32'hca00013;
      103851: inst = 32'h24822800;
      103852: inst = 32'h10a00000;
      103853: inst = 32'hca00004;
      103854: inst = 32'h38632800;
      103855: inst = 32'h38842800;
      103856: inst = 32'h10a00001;
      103857: inst = 32'hca095b5;
      103858: inst = 32'h13e00001;
      103859: inst = 32'hfe0d96a;
      103860: inst = 32'h5be00000;
      103861: inst = 32'h8c50000;
      103862: inst = 32'h24612800;
      103863: inst = 32'h10a00000;
      103864: inst = 32'hca00013;
      103865: inst = 32'h24822800;
      103866: inst = 32'h10a00000;
      103867: inst = 32'hca00004;
      103868: inst = 32'h38632800;
      103869: inst = 32'h38842800;
      103870: inst = 32'h10a00001;
      103871: inst = 32'hca095c3;
      103872: inst = 32'h13e00001;
      103873: inst = 32'hfe0d96a;
      103874: inst = 32'h5be00000;
      103875: inst = 32'h8c50000;
      103876: inst = 32'h24612800;
      103877: inst = 32'h10a00000;
      103878: inst = 32'hca00013;
      103879: inst = 32'h24822800;
      103880: inst = 32'h10a00000;
      103881: inst = 32'hca00004;
      103882: inst = 32'h38632800;
      103883: inst = 32'h38842800;
      103884: inst = 32'h10a00001;
      103885: inst = 32'hca095d1;
      103886: inst = 32'h13e00001;
      103887: inst = 32'hfe0d96a;
      103888: inst = 32'h5be00000;
      103889: inst = 32'h8c50000;
      103890: inst = 32'h24612800;
      103891: inst = 32'h10a00000;
      103892: inst = 32'hca00013;
      103893: inst = 32'h24822800;
      103894: inst = 32'h10a00000;
      103895: inst = 32'hca00004;
      103896: inst = 32'h38632800;
      103897: inst = 32'h38842800;
      103898: inst = 32'h10a00001;
      103899: inst = 32'hca095df;
      103900: inst = 32'h13e00001;
      103901: inst = 32'hfe0d96a;
      103902: inst = 32'h5be00000;
      103903: inst = 32'h8c50000;
      103904: inst = 32'h24612800;
      103905: inst = 32'h10a00000;
      103906: inst = 32'hca00013;
      103907: inst = 32'h24822800;
      103908: inst = 32'h10a00000;
      103909: inst = 32'hca00004;
      103910: inst = 32'h38632800;
      103911: inst = 32'h38842800;
      103912: inst = 32'h10a00001;
      103913: inst = 32'hca095ed;
      103914: inst = 32'h13e00001;
      103915: inst = 32'hfe0d96a;
      103916: inst = 32'h5be00000;
      103917: inst = 32'h8c50000;
      103918: inst = 32'h24612800;
      103919: inst = 32'h10a00000;
      103920: inst = 32'hca00013;
      103921: inst = 32'h24822800;
      103922: inst = 32'h10a00000;
      103923: inst = 32'hca00004;
      103924: inst = 32'h38632800;
      103925: inst = 32'h38842800;
      103926: inst = 32'h10a00001;
      103927: inst = 32'hca095fb;
      103928: inst = 32'h13e00001;
      103929: inst = 32'hfe0d96a;
      103930: inst = 32'h5be00000;
      103931: inst = 32'h8c50000;
      103932: inst = 32'h24612800;
      103933: inst = 32'h10a00000;
      103934: inst = 32'hca00013;
      103935: inst = 32'h24822800;
      103936: inst = 32'h10a00000;
      103937: inst = 32'hca00004;
      103938: inst = 32'h38632800;
      103939: inst = 32'h38842800;
      103940: inst = 32'h10a00001;
      103941: inst = 32'hca09609;
      103942: inst = 32'h13e00001;
      103943: inst = 32'hfe0d96a;
      103944: inst = 32'h5be00000;
      103945: inst = 32'h8c50000;
      103946: inst = 32'h24612800;
      103947: inst = 32'h10a00000;
      103948: inst = 32'hca00013;
      103949: inst = 32'h24822800;
      103950: inst = 32'h10a00000;
      103951: inst = 32'hca00004;
      103952: inst = 32'h38632800;
      103953: inst = 32'h38842800;
      103954: inst = 32'h10a00001;
      103955: inst = 32'hca09617;
      103956: inst = 32'h13e00001;
      103957: inst = 32'hfe0d96a;
      103958: inst = 32'h5be00000;
      103959: inst = 32'h8c50000;
      103960: inst = 32'h24612800;
      103961: inst = 32'h10a00000;
      103962: inst = 32'hca00013;
      103963: inst = 32'h24822800;
      103964: inst = 32'h10a00000;
      103965: inst = 32'hca00004;
      103966: inst = 32'h38632800;
      103967: inst = 32'h38842800;
      103968: inst = 32'h10a00001;
      103969: inst = 32'hca09625;
      103970: inst = 32'h13e00001;
      103971: inst = 32'hfe0d96a;
      103972: inst = 32'h5be00000;
      103973: inst = 32'h8c50000;
      103974: inst = 32'h24612800;
      103975: inst = 32'h10a00000;
      103976: inst = 32'hca00013;
      103977: inst = 32'h24822800;
      103978: inst = 32'h10a00000;
      103979: inst = 32'hca00004;
      103980: inst = 32'h38632800;
      103981: inst = 32'h38842800;
      103982: inst = 32'h10a00001;
      103983: inst = 32'hca09633;
      103984: inst = 32'h13e00001;
      103985: inst = 32'hfe0d96a;
      103986: inst = 32'h5be00000;
      103987: inst = 32'h8c50000;
      103988: inst = 32'h24612800;
      103989: inst = 32'h10a00000;
      103990: inst = 32'hca00013;
      103991: inst = 32'h24822800;
      103992: inst = 32'h10a00000;
      103993: inst = 32'hca00004;
      103994: inst = 32'h38632800;
      103995: inst = 32'h38842800;
      103996: inst = 32'h10a00001;
      103997: inst = 32'hca09641;
      103998: inst = 32'h13e00001;
      103999: inst = 32'hfe0d96a;
      104000: inst = 32'h5be00000;
      104001: inst = 32'h8c50000;
      104002: inst = 32'h24612800;
      104003: inst = 32'h10a00000;
      104004: inst = 32'hca00013;
      104005: inst = 32'h24822800;
      104006: inst = 32'h10a00000;
      104007: inst = 32'hca00004;
      104008: inst = 32'h38632800;
      104009: inst = 32'h38842800;
      104010: inst = 32'h10a00001;
      104011: inst = 32'hca0964f;
      104012: inst = 32'h13e00001;
      104013: inst = 32'hfe0d96a;
      104014: inst = 32'h5be00000;
      104015: inst = 32'h8c50000;
      104016: inst = 32'h24612800;
      104017: inst = 32'h10a00000;
      104018: inst = 32'hca00013;
      104019: inst = 32'h24822800;
      104020: inst = 32'h10a00000;
      104021: inst = 32'hca00004;
      104022: inst = 32'h38632800;
      104023: inst = 32'h38842800;
      104024: inst = 32'h10a00001;
      104025: inst = 32'hca0965d;
      104026: inst = 32'h13e00001;
      104027: inst = 32'hfe0d96a;
      104028: inst = 32'h5be00000;
      104029: inst = 32'h8c50000;
      104030: inst = 32'h24612800;
      104031: inst = 32'h10a00000;
      104032: inst = 32'hca00013;
      104033: inst = 32'h24822800;
      104034: inst = 32'h10a00000;
      104035: inst = 32'hca00004;
      104036: inst = 32'h38632800;
      104037: inst = 32'h38842800;
      104038: inst = 32'h10a00001;
      104039: inst = 32'hca0966b;
      104040: inst = 32'h13e00001;
      104041: inst = 32'hfe0d96a;
      104042: inst = 32'h5be00000;
      104043: inst = 32'h8c50000;
      104044: inst = 32'h24612800;
      104045: inst = 32'h10a00000;
      104046: inst = 32'hca00013;
      104047: inst = 32'h24822800;
      104048: inst = 32'h10a00000;
      104049: inst = 32'hca00004;
      104050: inst = 32'h38632800;
      104051: inst = 32'h38842800;
      104052: inst = 32'h10a00001;
      104053: inst = 32'hca09679;
      104054: inst = 32'h13e00001;
      104055: inst = 32'hfe0d96a;
      104056: inst = 32'h5be00000;
      104057: inst = 32'h8c50000;
      104058: inst = 32'h24612800;
      104059: inst = 32'h10a00000;
      104060: inst = 32'hca00013;
      104061: inst = 32'h24822800;
      104062: inst = 32'h10a00000;
      104063: inst = 32'hca00004;
      104064: inst = 32'h38632800;
      104065: inst = 32'h38842800;
      104066: inst = 32'h10a00001;
      104067: inst = 32'hca09687;
      104068: inst = 32'h13e00001;
      104069: inst = 32'hfe0d96a;
      104070: inst = 32'h5be00000;
      104071: inst = 32'h8c50000;
      104072: inst = 32'h24612800;
      104073: inst = 32'h10a00000;
      104074: inst = 32'hca00013;
      104075: inst = 32'h24822800;
      104076: inst = 32'h10a00000;
      104077: inst = 32'hca00004;
      104078: inst = 32'h38632800;
      104079: inst = 32'h38842800;
      104080: inst = 32'h10a00001;
      104081: inst = 32'hca09695;
      104082: inst = 32'h13e00001;
      104083: inst = 32'hfe0d96a;
      104084: inst = 32'h5be00000;
      104085: inst = 32'h8c50000;
      104086: inst = 32'h24612800;
      104087: inst = 32'h10a00000;
      104088: inst = 32'hca00013;
      104089: inst = 32'h24822800;
      104090: inst = 32'h10a00000;
      104091: inst = 32'hca00004;
      104092: inst = 32'h38632800;
      104093: inst = 32'h38842800;
      104094: inst = 32'h10a00001;
      104095: inst = 32'hca096a3;
      104096: inst = 32'h13e00001;
      104097: inst = 32'hfe0d96a;
      104098: inst = 32'h5be00000;
      104099: inst = 32'h8c50000;
      104100: inst = 32'h24612800;
      104101: inst = 32'h10a00000;
      104102: inst = 32'hca00013;
      104103: inst = 32'h24822800;
      104104: inst = 32'h10a00000;
      104105: inst = 32'hca00004;
      104106: inst = 32'h38632800;
      104107: inst = 32'h38842800;
      104108: inst = 32'h10a00001;
      104109: inst = 32'hca096b1;
      104110: inst = 32'h13e00001;
      104111: inst = 32'hfe0d96a;
      104112: inst = 32'h5be00000;
      104113: inst = 32'h8c50000;
      104114: inst = 32'h24612800;
      104115: inst = 32'h10a00000;
      104116: inst = 32'hca00013;
      104117: inst = 32'h24822800;
      104118: inst = 32'h10a00000;
      104119: inst = 32'hca00004;
      104120: inst = 32'h38632800;
      104121: inst = 32'h38842800;
      104122: inst = 32'h10a00001;
      104123: inst = 32'hca096bf;
      104124: inst = 32'h13e00001;
      104125: inst = 32'hfe0d96a;
      104126: inst = 32'h5be00000;
      104127: inst = 32'h8c50000;
      104128: inst = 32'h24612800;
      104129: inst = 32'h10a00000;
      104130: inst = 32'hca00013;
      104131: inst = 32'h24822800;
      104132: inst = 32'h10a00000;
      104133: inst = 32'hca00004;
      104134: inst = 32'h38632800;
      104135: inst = 32'h38842800;
      104136: inst = 32'h10a00001;
      104137: inst = 32'hca096cd;
      104138: inst = 32'h13e00001;
      104139: inst = 32'hfe0d96a;
      104140: inst = 32'h5be00000;
      104141: inst = 32'h8c50000;
      104142: inst = 32'h24612800;
      104143: inst = 32'h10a00000;
      104144: inst = 32'hca00013;
      104145: inst = 32'h24822800;
      104146: inst = 32'h10a00000;
      104147: inst = 32'hca00004;
      104148: inst = 32'h38632800;
      104149: inst = 32'h38842800;
      104150: inst = 32'h10a00001;
      104151: inst = 32'hca096db;
      104152: inst = 32'h13e00001;
      104153: inst = 32'hfe0d96a;
      104154: inst = 32'h5be00000;
      104155: inst = 32'h8c50000;
      104156: inst = 32'h24612800;
      104157: inst = 32'h10a00000;
      104158: inst = 32'hca00013;
      104159: inst = 32'h24822800;
      104160: inst = 32'h10a00000;
      104161: inst = 32'hca00004;
      104162: inst = 32'h38632800;
      104163: inst = 32'h38842800;
      104164: inst = 32'h10a00001;
      104165: inst = 32'hca096e9;
      104166: inst = 32'h13e00001;
      104167: inst = 32'hfe0d96a;
      104168: inst = 32'h5be00000;
      104169: inst = 32'h8c50000;
      104170: inst = 32'h24612800;
      104171: inst = 32'h10a00000;
      104172: inst = 32'hca00013;
      104173: inst = 32'h24822800;
      104174: inst = 32'h10a00000;
      104175: inst = 32'hca00004;
      104176: inst = 32'h38632800;
      104177: inst = 32'h38842800;
      104178: inst = 32'h10a00001;
      104179: inst = 32'hca096f7;
      104180: inst = 32'h13e00001;
      104181: inst = 32'hfe0d96a;
      104182: inst = 32'h5be00000;
      104183: inst = 32'h8c50000;
      104184: inst = 32'h24612800;
      104185: inst = 32'h10a00000;
      104186: inst = 32'hca00013;
      104187: inst = 32'h24822800;
      104188: inst = 32'h10a00000;
      104189: inst = 32'hca00004;
      104190: inst = 32'h38632800;
      104191: inst = 32'h38842800;
      104192: inst = 32'h10a00001;
      104193: inst = 32'hca09705;
      104194: inst = 32'h13e00001;
      104195: inst = 32'hfe0d96a;
      104196: inst = 32'h5be00000;
      104197: inst = 32'h8c50000;
      104198: inst = 32'h24612800;
      104199: inst = 32'h10a00000;
      104200: inst = 32'hca00013;
      104201: inst = 32'h24822800;
      104202: inst = 32'h10a00000;
      104203: inst = 32'hca00004;
      104204: inst = 32'h38632800;
      104205: inst = 32'h38842800;
      104206: inst = 32'h10a00001;
      104207: inst = 32'hca09713;
      104208: inst = 32'h13e00001;
      104209: inst = 32'hfe0d96a;
      104210: inst = 32'h5be00000;
      104211: inst = 32'h8c50000;
      104212: inst = 32'h24612800;
      104213: inst = 32'h10a00000;
      104214: inst = 32'hca00013;
      104215: inst = 32'h24822800;
      104216: inst = 32'h10a00000;
      104217: inst = 32'hca00004;
      104218: inst = 32'h38632800;
      104219: inst = 32'h38842800;
      104220: inst = 32'h10a00001;
      104221: inst = 32'hca09721;
      104222: inst = 32'h13e00001;
      104223: inst = 32'hfe0d96a;
      104224: inst = 32'h5be00000;
      104225: inst = 32'h8c50000;
      104226: inst = 32'h24612800;
      104227: inst = 32'h10a00000;
      104228: inst = 32'hca00013;
      104229: inst = 32'h24822800;
      104230: inst = 32'h10a00000;
      104231: inst = 32'hca00004;
      104232: inst = 32'h38632800;
      104233: inst = 32'h38842800;
      104234: inst = 32'h10a00001;
      104235: inst = 32'hca0972f;
      104236: inst = 32'h13e00001;
      104237: inst = 32'hfe0d96a;
      104238: inst = 32'h5be00000;
      104239: inst = 32'h8c50000;
      104240: inst = 32'h24612800;
      104241: inst = 32'h10a00000;
      104242: inst = 32'hca00013;
      104243: inst = 32'h24822800;
      104244: inst = 32'h10a00000;
      104245: inst = 32'hca00004;
      104246: inst = 32'h38632800;
      104247: inst = 32'h38842800;
      104248: inst = 32'h10a00001;
      104249: inst = 32'hca0973d;
      104250: inst = 32'h13e00001;
      104251: inst = 32'hfe0d96a;
      104252: inst = 32'h5be00000;
      104253: inst = 32'h8c50000;
      104254: inst = 32'h24612800;
      104255: inst = 32'h10a00000;
      104256: inst = 32'hca00013;
      104257: inst = 32'h24822800;
      104258: inst = 32'h10a00000;
      104259: inst = 32'hca00004;
      104260: inst = 32'h38632800;
      104261: inst = 32'h38842800;
      104262: inst = 32'h10a00001;
      104263: inst = 32'hca0974b;
      104264: inst = 32'h13e00001;
      104265: inst = 32'hfe0d96a;
      104266: inst = 32'h5be00000;
      104267: inst = 32'h8c50000;
      104268: inst = 32'h24612800;
      104269: inst = 32'h10a00000;
      104270: inst = 32'hca00013;
      104271: inst = 32'h24822800;
      104272: inst = 32'h10a00000;
      104273: inst = 32'hca00004;
      104274: inst = 32'h38632800;
      104275: inst = 32'h38842800;
      104276: inst = 32'h10a00001;
      104277: inst = 32'hca09759;
      104278: inst = 32'h13e00001;
      104279: inst = 32'hfe0d96a;
      104280: inst = 32'h5be00000;
      104281: inst = 32'h8c50000;
      104282: inst = 32'h24612800;
      104283: inst = 32'h10a00000;
      104284: inst = 32'hca00013;
      104285: inst = 32'h24822800;
      104286: inst = 32'h10a00000;
      104287: inst = 32'hca00004;
      104288: inst = 32'h38632800;
      104289: inst = 32'h38842800;
      104290: inst = 32'h10a00001;
      104291: inst = 32'hca09767;
      104292: inst = 32'h13e00001;
      104293: inst = 32'hfe0d96a;
      104294: inst = 32'h5be00000;
      104295: inst = 32'h8c50000;
      104296: inst = 32'h24612800;
      104297: inst = 32'h10a00000;
      104298: inst = 32'hca00013;
      104299: inst = 32'h24822800;
      104300: inst = 32'h10a00000;
      104301: inst = 32'hca00004;
      104302: inst = 32'h38632800;
      104303: inst = 32'h38842800;
      104304: inst = 32'h10a00001;
      104305: inst = 32'hca09775;
      104306: inst = 32'h13e00001;
      104307: inst = 32'hfe0d96a;
      104308: inst = 32'h5be00000;
      104309: inst = 32'h8c50000;
      104310: inst = 32'h24612800;
      104311: inst = 32'h10a00000;
      104312: inst = 32'hca00013;
      104313: inst = 32'h24822800;
      104314: inst = 32'h10a00000;
      104315: inst = 32'hca00004;
      104316: inst = 32'h38632800;
      104317: inst = 32'h38842800;
      104318: inst = 32'h10a00001;
      104319: inst = 32'hca09783;
      104320: inst = 32'h13e00001;
      104321: inst = 32'hfe0d96a;
      104322: inst = 32'h5be00000;
      104323: inst = 32'h8c50000;
      104324: inst = 32'h24612800;
      104325: inst = 32'h10a00000;
      104326: inst = 32'hca00013;
      104327: inst = 32'h24822800;
      104328: inst = 32'h10a00000;
      104329: inst = 32'hca00004;
      104330: inst = 32'h38632800;
      104331: inst = 32'h38842800;
      104332: inst = 32'h10a00001;
      104333: inst = 32'hca09791;
      104334: inst = 32'h13e00001;
      104335: inst = 32'hfe0d96a;
      104336: inst = 32'h5be00000;
      104337: inst = 32'h8c50000;
      104338: inst = 32'h24612800;
      104339: inst = 32'h10a00000;
      104340: inst = 32'hca00013;
      104341: inst = 32'h24822800;
      104342: inst = 32'h10a00000;
      104343: inst = 32'hca00004;
      104344: inst = 32'h38632800;
      104345: inst = 32'h38842800;
      104346: inst = 32'h10a00001;
      104347: inst = 32'hca0979f;
      104348: inst = 32'h13e00001;
      104349: inst = 32'hfe0d96a;
      104350: inst = 32'h5be00000;
      104351: inst = 32'h8c50000;
      104352: inst = 32'h24612800;
      104353: inst = 32'h10a00000;
      104354: inst = 32'hca00013;
      104355: inst = 32'h24822800;
      104356: inst = 32'h10a00000;
      104357: inst = 32'hca00004;
      104358: inst = 32'h38632800;
      104359: inst = 32'h38842800;
      104360: inst = 32'h10a00001;
      104361: inst = 32'hca097ad;
      104362: inst = 32'h13e00001;
      104363: inst = 32'hfe0d96a;
      104364: inst = 32'h5be00000;
      104365: inst = 32'h8c50000;
      104366: inst = 32'h24612800;
      104367: inst = 32'h10a00000;
      104368: inst = 32'hca00013;
      104369: inst = 32'h24822800;
      104370: inst = 32'h10a00000;
      104371: inst = 32'hca00004;
      104372: inst = 32'h38632800;
      104373: inst = 32'h38842800;
      104374: inst = 32'h10a00001;
      104375: inst = 32'hca097bb;
      104376: inst = 32'h13e00001;
      104377: inst = 32'hfe0d96a;
      104378: inst = 32'h5be00000;
      104379: inst = 32'h8c50000;
      104380: inst = 32'h24612800;
      104381: inst = 32'h10a00000;
      104382: inst = 32'hca00013;
      104383: inst = 32'h24822800;
      104384: inst = 32'h10a00000;
      104385: inst = 32'hca00004;
      104386: inst = 32'h38632800;
      104387: inst = 32'h38842800;
      104388: inst = 32'h10a00001;
      104389: inst = 32'hca097c9;
      104390: inst = 32'h13e00001;
      104391: inst = 32'hfe0d96a;
      104392: inst = 32'h5be00000;
      104393: inst = 32'h8c50000;
      104394: inst = 32'h24612800;
      104395: inst = 32'h10a00000;
      104396: inst = 32'hca00013;
      104397: inst = 32'h24822800;
      104398: inst = 32'h10a00000;
      104399: inst = 32'hca00004;
      104400: inst = 32'h38632800;
      104401: inst = 32'h38842800;
      104402: inst = 32'h10a00001;
      104403: inst = 32'hca097d7;
      104404: inst = 32'h13e00001;
      104405: inst = 32'hfe0d96a;
      104406: inst = 32'h5be00000;
      104407: inst = 32'h8c50000;
      104408: inst = 32'h24612800;
      104409: inst = 32'h10a00000;
      104410: inst = 32'hca00013;
      104411: inst = 32'h24822800;
      104412: inst = 32'h10a00000;
      104413: inst = 32'hca00004;
      104414: inst = 32'h38632800;
      104415: inst = 32'h38842800;
      104416: inst = 32'h10a00001;
      104417: inst = 32'hca097e5;
      104418: inst = 32'h13e00001;
      104419: inst = 32'hfe0d96a;
      104420: inst = 32'h5be00000;
      104421: inst = 32'h8c50000;
      104422: inst = 32'h24612800;
      104423: inst = 32'h10a00000;
      104424: inst = 32'hca00013;
      104425: inst = 32'h24822800;
      104426: inst = 32'h10a00000;
      104427: inst = 32'hca00004;
      104428: inst = 32'h38632800;
      104429: inst = 32'h38842800;
      104430: inst = 32'h10a00001;
      104431: inst = 32'hca097f3;
      104432: inst = 32'h13e00001;
      104433: inst = 32'hfe0d96a;
      104434: inst = 32'h5be00000;
      104435: inst = 32'h8c50000;
      104436: inst = 32'h24612800;
      104437: inst = 32'h10a00000;
      104438: inst = 32'hca00013;
      104439: inst = 32'h24822800;
      104440: inst = 32'h10a00000;
      104441: inst = 32'hca00004;
      104442: inst = 32'h38632800;
      104443: inst = 32'h38842800;
      104444: inst = 32'h10a00001;
      104445: inst = 32'hca09801;
      104446: inst = 32'h13e00001;
      104447: inst = 32'hfe0d96a;
      104448: inst = 32'h5be00000;
      104449: inst = 32'h8c50000;
      104450: inst = 32'h24612800;
      104451: inst = 32'h10a00000;
      104452: inst = 32'hca00013;
      104453: inst = 32'h24822800;
      104454: inst = 32'h10a00000;
      104455: inst = 32'hca00004;
      104456: inst = 32'h38632800;
      104457: inst = 32'h38842800;
      104458: inst = 32'h10a00001;
      104459: inst = 32'hca0980f;
      104460: inst = 32'h13e00001;
      104461: inst = 32'hfe0d96a;
      104462: inst = 32'h5be00000;
      104463: inst = 32'h8c50000;
      104464: inst = 32'h24612800;
      104465: inst = 32'h10a00000;
      104466: inst = 32'hca00013;
      104467: inst = 32'h24822800;
      104468: inst = 32'h10a00000;
      104469: inst = 32'hca00004;
      104470: inst = 32'h38632800;
      104471: inst = 32'h38842800;
      104472: inst = 32'h10a00001;
      104473: inst = 32'hca0981d;
      104474: inst = 32'h13e00001;
      104475: inst = 32'hfe0d96a;
      104476: inst = 32'h5be00000;
      104477: inst = 32'h8c50000;
      104478: inst = 32'h24612800;
      104479: inst = 32'h10a00000;
      104480: inst = 32'hca00013;
      104481: inst = 32'h24822800;
      104482: inst = 32'h10a00000;
      104483: inst = 32'hca00004;
      104484: inst = 32'h38632800;
      104485: inst = 32'h38842800;
      104486: inst = 32'h10a00001;
      104487: inst = 32'hca0982b;
      104488: inst = 32'h13e00001;
      104489: inst = 32'hfe0d96a;
      104490: inst = 32'h5be00000;
      104491: inst = 32'h8c50000;
      104492: inst = 32'h24612800;
      104493: inst = 32'h10a00000;
      104494: inst = 32'hca00013;
      104495: inst = 32'h24822800;
      104496: inst = 32'h10a00000;
      104497: inst = 32'hca00004;
      104498: inst = 32'h38632800;
      104499: inst = 32'h38842800;
      104500: inst = 32'h10a00001;
      104501: inst = 32'hca09839;
      104502: inst = 32'h13e00001;
      104503: inst = 32'hfe0d96a;
      104504: inst = 32'h5be00000;
      104505: inst = 32'h8c50000;
      104506: inst = 32'h24612800;
      104507: inst = 32'h10a00000;
      104508: inst = 32'hca00013;
      104509: inst = 32'h24822800;
      104510: inst = 32'h10a00000;
      104511: inst = 32'hca00004;
      104512: inst = 32'h38632800;
      104513: inst = 32'h38842800;
      104514: inst = 32'h10a00001;
      104515: inst = 32'hca09847;
      104516: inst = 32'h13e00001;
      104517: inst = 32'hfe0d96a;
      104518: inst = 32'h5be00000;
      104519: inst = 32'h8c50000;
      104520: inst = 32'h24612800;
      104521: inst = 32'h10a00000;
      104522: inst = 32'hca00013;
      104523: inst = 32'h24822800;
      104524: inst = 32'h10a00000;
      104525: inst = 32'hca00004;
      104526: inst = 32'h38632800;
      104527: inst = 32'h38842800;
      104528: inst = 32'h10a00001;
      104529: inst = 32'hca09855;
      104530: inst = 32'h13e00001;
      104531: inst = 32'hfe0d96a;
      104532: inst = 32'h5be00000;
      104533: inst = 32'h8c50000;
      104534: inst = 32'h24612800;
      104535: inst = 32'h10a00000;
      104536: inst = 32'hca00013;
      104537: inst = 32'h24822800;
      104538: inst = 32'h10a00000;
      104539: inst = 32'hca00004;
      104540: inst = 32'h38632800;
      104541: inst = 32'h38842800;
      104542: inst = 32'h10a00001;
      104543: inst = 32'hca09863;
      104544: inst = 32'h13e00001;
      104545: inst = 32'hfe0d96a;
      104546: inst = 32'h5be00000;
      104547: inst = 32'h8c50000;
      104548: inst = 32'h24612800;
      104549: inst = 32'h10a00000;
      104550: inst = 32'hca00013;
      104551: inst = 32'h24822800;
      104552: inst = 32'h10a00000;
      104553: inst = 32'hca00004;
      104554: inst = 32'h38632800;
      104555: inst = 32'h38842800;
      104556: inst = 32'h10a00001;
      104557: inst = 32'hca09871;
      104558: inst = 32'h13e00001;
      104559: inst = 32'hfe0d96a;
      104560: inst = 32'h5be00000;
      104561: inst = 32'h8c50000;
      104562: inst = 32'h24612800;
      104563: inst = 32'h10a00000;
      104564: inst = 32'hca00013;
      104565: inst = 32'h24822800;
      104566: inst = 32'h10a00000;
      104567: inst = 32'hca00004;
      104568: inst = 32'h38632800;
      104569: inst = 32'h38842800;
      104570: inst = 32'h10a00001;
      104571: inst = 32'hca0987f;
      104572: inst = 32'h13e00001;
      104573: inst = 32'hfe0d96a;
      104574: inst = 32'h5be00000;
      104575: inst = 32'h8c50000;
      104576: inst = 32'h24612800;
      104577: inst = 32'h10a00000;
      104578: inst = 32'hca00013;
      104579: inst = 32'h24822800;
      104580: inst = 32'h10a00000;
      104581: inst = 32'hca00004;
      104582: inst = 32'h38632800;
      104583: inst = 32'h38842800;
      104584: inst = 32'h10a00001;
      104585: inst = 32'hca0988d;
      104586: inst = 32'h13e00001;
      104587: inst = 32'hfe0d96a;
      104588: inst = 32'h5be00000;
      104589: inst = 32'h8c50000;
      104590: inst = 32'h24612800;
      104591: inst = 32'h10a00000;
      104592: inst = 32'hca00013;
      104593: inst = 32'h24822800;
      104594: inst = 32'h10a00000;
      104595: inst = 32'hca00004;
      104596: inst = 32'h38632800;
      104597: inst = 32'h38842800;
      104598: inst = 32'h10a00001;
      104599: inst = 32'hca0989b;
      104600: inst = 32'h13e00001;
      104601: inst = 32'hfe0d96a;
      104602: inst = 32'h5be00000;
      104603: inst = 32'h8c50000;
      104604: inst = 32'h24612800;
      104605: inst = 32'h10a00000;
      104606: inst = 32'hca00013;
      104607: inst = 32'h24822800;
      104608: inst = 32'h10a00000;
      104609: inst = 32'hca00004;
      104610: inst = 32'h38632800;
      104611: inst = 32'h38842800;
      104612: inst = 32'h10a00001;
      104613: inst = 32'hca098a9;
      104614: inst = 32'h13e00001;
      104615: inst = 32'hfe0d96a;
      104616: inst = 32'h5be00000;
      104617: inst = 32'h8c50000;
      104618: inst = 32'h24612800;
      104619: inst = 32'h10a00000;
      104620: inst = 32'hca00013;
      104621: inst = 32'h24822800;
      104622: inst = 32'h10a00000;
      104623: inst = 32'hca00004;
      104624: inst = 32'h38632800;
      104625: inst = 32'h38842800;
      104626: inst = 32'h10a00001;
      104627: inst = 32'hca098b7;
      104628: inst = 32'h13e00001;
      104629: inst = 32'hfe0d96a;
      104630: inst = 32'h5be00000;
      104631: inst = 32'h8c50000;
      104632: inst = 32'h24612800;
      104633: inst = 32'h10a00000;
      104634: inst = 32'hca00013;
      104635: inst = 32'h24822800;
      104636: inst = 32'h10a00000;
      104637: inst = 32'hca00004;
      104638: inst = 32'h38632800;
      104639: inst = 32'h38842800;
      104640: inst = 32'h10a00001;
      104641: inst = 32'hca098c5;
      104642: inst = 32'h13e00001;
      104643: inst = 32'hfe0d96a;
      104644: inst = 32'h5be00000;
      104645: inst = 32'h8c50000;
      104646: inst = 32'h24612800;
      104647: inst = 32'h10a00000;
      104648: inst = 32'hca00013;
      104649: inst = 32'h24822800;
      104650: inst = 32'h10a00000;
      104651: inst = 32'hca00004;
      104652: inst = 32'h38632800;
      104653: inst = 32'h38842800;
      104654: inst = 32'h10a00001;
      104655: inst = 32'hca098d3;
      104656: inst = 32'h13e00001;
      104657: inst = 32'hfe0d96a;
      104658: inst = 32'h5be00000;
      104659: inst = 32'h8c50000;
      104660: inst = 32'h24612800;
      104661: inst = 32'h10a00000;
      104662: inst = 32'hca00013;
      104663: inst = 32'h24822800;
      104664: inst = 32'h10a00000;
      104665: inst = 32'hca00004;
      104666: inst = 32'h38632800;
      104667: inst = 32'h38842800;
      104668: inst = 32'h10a00001;
      104669: inst = 32'hca098e1;
      104670: inst = 32'h13e00001;
      104671: inst = 32'hfe0d96a;
      104672: inst = 32'h5be00000;
      104673: inst = 32'h8c50000;
      104674: inst = 32'h24612800;
      104675: inst = 32'h10a00000;
      104676: inst = 32'hca00013;
      104677: inst = 32'h24822800;
      104678: inst = 32'h10a00000;
      104679: inst = 32'hca00004;
      104680: inst = 32'h38632800;
      104681: inst = 32'h38842800;
      104682: inst = 32'h10a00001;
      104683: inst = 32'hca098ef;
      104684: inst = 32'h13e00001;
      104685: inst = 32'hfe0d96a;
      104686: inst = 32'h5be00000;
      104687: inst = 32'h8c50000;
      104688: inst = 32'h24612800;
      104689: inst = 32'h10a00000;
      104690: inst = 32'hca00013;
      104691: inst = 32'h24822800;
      104692: inst = 32'h10a00000;
      104693: inst = 32'hca00004;
      104694: inst = 32'h38632800;
      104695: inst = 32'h38842800;
      104696: inst = 32'h10a00001;
      104697: inst = 32'hca098fd;
      104698: inst = 32'h13e00001;
      104699: inst = 32'hfe0d96a;
      104700: inst = 32'h5be00000;
      104701: inst = 32'h8c50000;
      104702: inst = 32'h24612800;
      104703: inst = 32'h10a00000;
      104704: inst = 32'hca00013;
      104705: inst = 32'h24822800;
      104706: inst = 32'h10a00000;
      104707: inst = 32'hca00004;
      104708: inst = 32'h38632800;
      104709: inst = 32'h38842800;
      104710: inst = 32'h10a00001;
      104711: inst = 32'hca0990b;
      104712: inst = 32'h13e00001;
      104713: inst = 32'hfe0d96a;
      104714: inst = 32'h5be00000;
      104715: inst = 32'h8c50000;
      104716: inst = 32'h24612800;
      104717: inst = 32'h10a00000;
      104718: inst = 32'hca00013;
      104719: inst = 32'h24822800;
      104720: inst = 32'h10a00000;
      104721: inst = 32'hca00004;
      104722: inst = 32'h38632800;
      104723: inst = 32'h38842800;
      104724: inst = 32'h10a00001;
      104725: inst = 32'hca09919;
      104726: inst = 32'h13e00001;
      104727: inst = 32'hfe0d96a;
      104728: inst = 32'h5be00000;
      104729: inst = 32'h8c50000;
      104730: inst = 32'h24612800;
      104731: inst = 32'h10a00000;
      104732: inst = 32'hca00013;
      104733: inst = 32'h24822800;
      104734: inst = 32'h10a00000;
      104735: inst = 32'hca00004;
      104736: inst = 32'h38632800;
      104737: inst = 32'h38842800;
      104738: inst = 32'h10a00001;
      104739: inst = 32'hca09927;
      104740: inst = 32'h13e00001;
      104741: inst = 32'hfe0d96a;
      104742: inst = 32'h5be00000;
      104743: inst = 32'h8c50000;
      104744: inst = 32'h24612800;
      104745: inst = 32'h10a00000;
      104746: inst = 32'hca00013;
      104747: inst = 32'h24822800;
      104748: inst = 32'h10a00000;
      104749: inst = 32'hca00004;
      104750: inst = 32'h38632800;
      104751: inst = 32'h38842800;
      104752: inst = 32'h10a00001;
      104753: inst = 32'hca09935;
      104754: inst = 32'h13e00001;
      104755: inst = 32'hfe0d96a;
      104756: inst = 32'h5be00000;
      104757: inst = 32'h8c50000;
      104758: inst = 32'h24612800;
      104759: inst = 32'h10a00000;
      104760: inst = 32'hca00013;
      104761: inst = 32'h24822800;
      104762: inst = 32'h10a00000;
      104763: inst = 32'hca00004;
      104764: inst = 32'h38632800;
      104765: inst = 32'h38842800;
      104766: inst = 32'h10a00001;
      104767: inst = 32'hca09943;
      104768: inst = 32'h13e00001;
      104769: inst = 32'hfe0d96a;
      104770: inst = 32'h5be00000;
      104771: inst = 32'h8c50000;
      104772: inst = 32'h24612800;
      104773: inst = 32'h10a00000;
      104774: inst = 32'hca00013;
      104775: inst = 32'h24822800;
      104776: inst = 32'h10a00000;
      104777: inst = 32'hca00004;
      104778: inst = 32'h38632800;
      104779: inst = 32'h38842800;
      104780: inst = 32'h10a00001;
      104781: inst = 32'hca09951;
      104782: inst = 32'h13e00001;
      104783: inst = 32'hfe0d96a;
      104784: inst = 32'h5be00000;
      104785: inst = 32'h8c50000;
      104786: inst = 32'h24612800;
      104787: inst = 32'h10a00000;
      104788: inst = 32'hca00013;
      104789: inst = 32'h24822800;
      104790: inst = 32'h10a00000;
      104791: inst = 32'hca00004;
      104792: inst = 32'h38632800;
      104793: inst = 32'h38842800;
      104794: inst = 32'h10a00001;
      104795: inst = 32'hca0995f;
      104796: inst = 32'h13e00001;
      104797: inst = 32'hfe0d96a;
      104798: inst = 32'h5be00000;
      104799: inst = 32'h8c50000;
      104800: inst = 32'h24612800;
      104801: inst = 32'h10a00000;
      104802: inst = 32'hca00013;
      104803: inst = 32'h24822800;
      104804: inst = 32'h10a00000;
      104805: inst = 32'hca00004;
      104806: inst = 32'h38632800;
      104807: inst = 32'h38842800;
      104808: inst = 32'h10a00001;
      104809: inst = 32'hca0996d;
      104810: inst = 32'h13e00001;
      104811: inst = 32'hfe0d96a;
      104812: inst = 32'h5be00000;
      104813: inst = 32'h8c50000;
      104814: inst = 32'h24612800;
      104815: inst = 32'h10a00000;
      104816: inst = 32'hca00013;
      104817: inst = 32'h24822800;
      104818: inst = 32'h10a00000;
      104819: inst = 32'hca00004;
      104820: inst = 32'h38632800;
      104821: inst = 32'h38842800;
      104822: inst = 32'h10a00001;
      104823: inst = 32'hca0997b;
      104824: inst = 32'h13e00001;
      104825: inst = 32'hfe0d96a;
      104826: inst = 32'h5be00000;
      104827: inst = 32'h8c50000;
      104828: inst = 32'h24612800;
      104829: inst = 32'h10a00000;
      104830: inst = 32'hca00013;
      104831: inst = 32'h24822800;
      104832: inst = 32'h10a00000;
      104833: inst = 32'hca00004;
      104834: inst = 32'h38632800;
      104835: inst = 32'h38842800;
      104836: inst = 32'h10a00001;
      104837: inst = 32'hca09989;
      104838: inst = 32'h13e00001;
      104839: inst = 32'hfe0d96a;
      104840: inst = 32'h5be00000;
      104841: inst = 32'h8c50000;
      104842: inst = 32'h24612800;
      104843: inst = 32'h10a00000;
      104844: inst = 32'hca00013;
      104845: inst = 32'h24822800;
      104846: inst = 32'h10a00000;
      104847: inst = 32'hca00004;
      104848: inst = 32'h38632800;
      104849: inst = 32'h38842800;
      104850: inst = 32'h10a00001;
      104851: inst = 32'hca09997;
      104852: inst = 32'h13e00001;
      104853: inst = 32'hfe0d96a;
      104854: inst = 32'h5be00000;
      104855: inst = 32'h8c50000;
      104856: inst = 32'h24612800;
      104857: inst = 32'h10a00000;
      104858: inst = 32'hca00013;
      104859: inst = 32'h24822800;
      104860: inst = 32'h10a00000;
      104861: inst = 32'hca00004;
      104862: inst = 32'h38632800;
      104863: inst = 32'h38842800;
      104864: inst = 32'h10a00001;
      104865: inst = 32'hca099a5;
      104866: inst = 32'h13e00001;
      104867: inst = 32'hfe0d96a;
      104868: inst = 32'h5be00000;
      104869: inst = 32'h8c50000;
      104870: inst = 32'h24612800;
      104871: inst = 32'h10a00000;
      104872: inst = 32'hca00013;
      104873: inst = 32'h24822800;
      104874: inst = 32'h10a00000;
      104875: inst = 32'hca00004;
      104876: inst = 32'h38632800;
      104877: inst = 32'h38842800;
      104878: inst = 32'h10a00001;
      104879: inst = 32'hca099b3;
      104880: inst = 32'h13e00001;
      104881: inst = 32'hfe0d96a;
      104882: inst = 32'h5be00000;
      104883: inst = 32'h8c50000;
      104884: inst = 32'h24612800;
      104885: inst = 32'h10a00000;
      104886: inst = 32'hca00013;
      104887: inst = 32'h24822800;
      104888: inst = 32'h10a00000;
      104889: inst = 32'hca00004;
      104890: inst = 32'h38632800;
      104891: inst = 32'h38842800;
      104892: inst = 32'h10a00001;
      104893: inst = 32'hca099c1;
      104894: inst = 32'h13e00001;
      104895: inst = 32'hfe0d96a;
      104896: inst = 32'h5be00000;
      104897: inst = 32'h8c50000;
      104898: inst = 32'h24612800;
      104899: inst = 32'h10a00000;
      104900: inst = 32'hca00013;
      104901: inst = 32'h24822800;
      104902: inst = 32'h10a00000;
      104903: inst = 32'hca00004;
      104904: inst = 32'h38632800;
      104905: inst = 32'h38842800;
      104906: inst = 32'h10a00001;
      104907: inst = 32'hca099cf;
      104908: inst = 32'h13e00001;
      104909: inst = 32'hfe0d96a;
      104910: inst = 32'h5be00000;
      104911: inst = 32'h8c50000;
      104912: inst = 32'h24612800;
      104913: inst = 32'h10a00000;
      104914: inst = 32'hca00013;
      104915: inst = 32'h24822800;
      104916: inst = 32'h10a00000;
      104917: inst = 32'hca00004;
      104918: inst = 32'h38632800;
      104919: inst = 32'h38842800;
      104920: inst = 32'h10a00001;
      104921: inst = 32'hca099dd;
      104922: inst = 32'h13e00001;
      104923: inst = 32'hfe0d96a;
      104924: inst = 32'h5be00000;
      104925: inst = 32'h8c50000;
      104926: inst = 32'h24612800;
      104927: inst = 32'h10a00000;
      104928: inst = 32'hca00013;
      104929: inst = 32'h24822800;
      104930: inst = 32'h10a00000;
      104931: inst = 32'hca00004;
      104932: inst = 32'h38632800;
      104933: inst = 32'h38842800;
      104934: inst = 32'h10a00001;
      104935: inst = 32'hca099eb;
      104936: inst = 32'h13e00001;
      104937: inst = 32'hfe0d96a;
      104938: inst = 32'h5be00000;
      104939: inst = 32'h8c50000;
      104940: inst = 32'h24612800;
      104941: inst = 32'h10a00000;
      104942: inst = 32'hca00013;
      104943: inst = 32'h24822800;
      104944: inst = 32'h10a00000;
      104945: inst = 32'hca00004;
      104946: inst = 32'h38632800;
      104947: inst = 32'h38842800;
      104948: inst = 32'h10a00001;
      104949: inst = 32'hca099f9;
      104950: inst = 32'h13e00001;
      104951: inst = 32'hfe0d96a;
      104952: inst = 32'h5be00000;
      104953: inst = 32'h8c50000;
      104954: inst = 32'h24612800;
      104955: inst = 32'h10a00000;
      104956: inst = 32'hca00013;
      104957: inst = 32'h24822800;
      104958: inst = 32'h10a00000;
      104959: inst = 32'hca00004;
      104960: inst = 32'h38632800;
      104961: inst = 32'h38842800;
      104962: inst = 32'h10a00001;
      104963: inst = 32'hca09a07;
      104964: inst = 32'h13e00001;
      104965: inst = 32'hfe0d96a;
      104966: inst = 32'h5be00000;
      104967: inst = 32'h8c50000;
      104968: inst = 32'h24612800;
      104969: inst = 32'h10a00000;
      104970: inst = 32'hca00013;
      104971: inst = 32'h24822800;
      104972: inst = 32'h10a00000;
      104973: inst = 32'hca00004;
      104974: inst = 32'h38632800;
      104975: inst = 32'h38842800;
      104976: inst = 32'h10a00001;
      104977: inst = 32'hca09a15;
      104978: inst = 32'h13e00001;
      104979: inst = 32'hfe0d96a;
      104980: inst = 32'h5be00000;
      104981: inst = 32'h8c50000;
      104982: inst = 32'h24612800;
      104983: inst = 32'h10a00000;
      104984: inst = 32'hca00013;
      104985: inst = 32'h24822800;
      104986: inst = 32'h10a00000;
      104987: inst = 32'hca00004;
      104988: inst = 32'h38632800;
      104989: inst = 32'h38842800;
      104990: inst = 32'h10a00001;
      104991: inst = 32'hca09a23;
      104992: inst = 32'h13e00001;
      104993: inst = 32'hfe0d96a;
      104994: inst = 32'h5be00000;
      104995: inst = 32'h8c50000;
      104996: inst = 32'h24612800;
      104997: inst = 32'h10a00000;
      104998: inst = 32'hca00013;
      104999: inst = 32'h24822800;
      105000: inst = 32'h10a00000;
      105001: inst = 32'hca00004;
      105002: inst = 32'h38632800;
      105003: inst = 32'h38842800;
      105004: inst = 32'h10a00001;
      105005: inst = 32'hca09a31;
      105006: inst = 32'h13e00001;
      105007: inst = 32'hfe0d96a;
      105008: inst = 32'h5be00000;
      105009: inst = 32'h8c50000;
      105010: inst = 32'h24612800;
      105011: inst = 32'h10a00000;
      105012: inst = 32'hca00013;
      105013: inst = 32'h24822800;
      105014: inst = 32'h10a00000;
      105015: inst = 32'hca00004;
      105016: inst = 32'h38632800;
      105017: inst = 32'h38842800;
      105018: inst = 32'h10a00001;
      105019: inst = 32'hca09a3f;
      105020: inst = 32'h13e00001;
      105021: inst = 32'hfe0d96a;
      105022: inst = 32'h5be00000;
      105023: inst = 32'h8c50000;
      105024: inst = 32'h24612800;
      105025: inst = 32'h10a00000;
      105026: inst = 32'hca00013;
      105027: inst = 32'h24822800;
      105028: inst = 32'h10a00000;
      105029: inst = 32'hca00004;
      105030: inst = 32'h38632800;
      105031: inst = 32'h38842800;
      105032: inst = 32'h10a00001;
      105033: inst = 32'hca09a4d;
      105034: inst = 32'h13e00001;
      105035: inst = 32'hfe0d96a;
      105036: inst = 32'h5be00000;
      105037: inst = 32'h8c50000;
      105038: inst = 32'h24612800;
      105039: inst = 32'h10a00000;
      105040: inst = 32'hca00013;
      105041: inst = 32'h24822800;
      105042: inst = 32'h10a00000;
      105043: inst = 32'hca00004;
      105044: inst = 32'h38632800;
      105045: inst = 32'h38842800;
      105046: inst = 32'h10a00001;
      105047: inst = 32'hca09a5b;
      105048: inst = 32'h13e00001;
      105049: inst = 32'hfe0d96a;
      105050: inst = 32'h5be00000;
      105051: inst = 32'h8c50000;
      105052: inst = 32'h24612800;
      105053: inst = 32'h10a00000;
      105054: inst = 32'hca00013;
      105055: inst = 32'h24822800;
      105056: inst = 32'h10a00000;
      105057: inst = 32'hca00004;
      105058: inst = 32'h38632800;
      105059: inst = 32'h38842800;
      105060: inst = 32'h10a00001;
      105061: inst = 32'hca09a69;
      105062: inst = 32'h13e00001;
      105063: inst = 32'hfe0d96a;
      105064: inst = 32'h5be00000;
      105065: inst = 32'h8c50000;
      105066: inst = 32'h24612800;
      105067: inst = 32'h10a00000;
      105068: inst = 32'hca00014;
      105069: inst = 32'h24822800;
      105070: inst = 32'h10a00000;
      105071: inst = 32'hca00004;
      105072: inst = 32'h38632800;
      105073: inst = 32'h38842800;
      105074: inst = 32'h10a00001;
      105075: inst = 32'hca09a77;
      105076: inst = 32'h13e00001;
      105077: inst = 32'hfe0d96a;
      105078: inst = 32'h5be00000;
      105079: inst = 32'h8c50000;
      105080: inst = 32'h24612800;
      105081: inst = 32'h10a00000;
      105082: inst = 32'hca00014;
      105083: inst = 32'h24822800;
      105084: inst = 32'h10a00000;
      105085: inst = 32'hca00004;
      105086: inst = 32'h38632800;
      105087: inst = 32'h38842800;
      105088: inst = 32'h10a00001;
      105089: inst = 32'hca09a85;
      105090: inst = 32'h13e00001;
      105091: inst = 32'hfe0d96a;
      105092: inst = 32'h5be00000;
      105093: inst = 32'h8c50000;
      105094: inst = 32'h24612800;
      105095: inst = 32'h10a00000;
      105096: inst = 32'hca00014;
      105097: inst = 32'h24822800;
      105098: inst = 32'h10a00000;
      105099: inst = 32'hca00004;
      105100: inst = 32'h38632800;
      105101: inst = 32'h38842800;
      105102: inst = 32'h10a00001;
      105103: inst = 32'hca09a93;
      105104: inst = 32'h13e00001;
      105105: inst = 32'hfe0d96a;
      105106: inst = 32'h5be00000;
      105107: inst = 32'h8c50000;
      105108: inst = 32'h24612800;
      105109: inst = 32'h10a00000;
      105110: inst = 32'hca00014;
      105111: inst = 32'h24822800;
      105112: inst = 32'h10a00000;
      105113: inst = 32'hca00004;
      105114: inst = 32'h38632800;
      105115: inst = 32'h38842800;
      105116: inst = 32'h10a00001;
      105117: inst = 32'hca09aa1;
      105118: inst = 32'h13e00001;
      105119: inst = 32'hfe0d96a;
      105120: inst = 32'h5be00000;
      105121: inst = 32'h8c50000;
      105122: inst = 32'h24612800;
      105123: inst = 32'h10a00000;
      105124: inst = 32'hca00014;
      105125: inst = 32'h24822800;
      105126: inst = 32'h10a00000;
      105127: inst = 32'hca00004;
      105128: inst = 32'h38632800;
      105129: inst = 32'h38842800;
      105130: inst = 32'h10a00001;
      105131: inst = 32'hca09aaf;
      105132: inst = 32'h13e00001;
      105133: inst = 32'hfe0d96a;
      105134: inst = 32'h5be00000;
      105135: inst = 32'h8c50000;
      105136: inst = 32'h24612800;
      105137: inst = 32'h10a00000;
      105138: inst = 32'hca00014;
      105139: inst = 32'h24822800;
      105140: inst = 32'h10a00000;
      105141: inst = 32'hca00004;
      105142: inst = 32'h38632800;
      105143: inst = 32'h38842800;
      105144: inst = 32'h10a00001;
      105145: inst = 32'hca09abd;
      105146: inst = 32'h13e00001;
      105147: inst = 32'hfe0d96a;
      105148: inst = 32'h5be00000;
      105149: inst = 32'h8c50000;
      105150: inst = 32'h24612800;
      105151: inst = 32'h10a00000;
      105152: inst = 32'hca00014;
      105153: inst = 32'h24822800;
      105154: inst = 32'h10a00000;
      105155: inst = 32'hca00004;
      105156: inst = 32'h38632800;
      105157: inst = 32'h38842800;
      105158: inst = 32'h10a00001;
      105159: inst = 32'hca09acb;
      105160: inst = 32'h13e00001;
      105161: inst = 32'hfe0d96a;
      105162: inst = 32'h5be00000;
      105163: inst = 32'h8c50000;
      105164: inst = 32'h24612800;
      105165: inst = 32'h10a00000;
      105166: inst = 32'hca00014;
      105167: inst = 32'h24822800;
      105168: inst = 32'h10a00000;
      105169: inst = 32'hca00004;
      105170: inst = 32'h38632800;
      105171: inst = 32'h38842800;
      105172: inst = 32'h10a00001;
      105173: inst = 32'hca09ad9;
      105174: inst = 32'h13e00001;
      105175: inst = 32'hfe0d96a;
      105176: inst = 32'h5be00000;
      105177: inst = 32'h8c50000;
      105178: inst = 32'h24612800;
      105179: inst = 32'h10a00000;
      105180: inst = 32'hca00014;
      105181: inst = 32'h24822800;
      105182: inst = 32'h10a00000;
      105183: inst = 32'hca00004;
      105184: inst = 32'h38632800;
      105185: inst = 32'h38842800;
      105186: inst = 32'h10a00001;
      105187: inst = 32'hca09ae7;
      105188: inst = 32'h13e00001;
      105189: inst = 32'hfe0d96a;
      105190: inst = 32'h5be00000;
      105191: inst = 32'h8c50000;
      105192: inst = 32'h24612800;
      105193: inst = 32'h10a00000;
      105194: inst = 32'hca00014;
      105195: inst = 32'h24822800;
      105196: inst = 32'h10a00000;
      105197: inst = 32'hca00004;
      105198: inst = 32'h38632800;
      105199: inst = 32'h38842800;
      105200: inst = 32'h10a00001;
      105201: inst = 32'hca09af5;
      105202: inst = 32'h13e00001;
      105203: inst = 32'hfe0d96a;
      105204: inst = 32'h5be00000;
      105205: inst = 32'h8c50000;
      105206: inst = 32'h24612800;
      105207: inst = 32'h10a00000;
      105208: inst = 32'hca00014;
      105209: inst = 32'h24822800;
      105210: inst = 32'h10a00000;
      105211: inst = 32'hca00004;
      105212: inst = 32'h38632800;
      105213: inst = 32'h38842800;
      105214: inst = 32'h10a00001;
      105215: inst = 32'hca09b03;
      105216: inst = 32'h13e00001;
      105217: inst = 32'hfe0d96a;
      105218: inst = 32'h5be00000;
      105219: inst = 32'h8c50000;
      105220: inst = 32'h24612800;
      105221: inst = 32'h10a00000;
      105222: inst = 32'hca00014;
      105223: inst = 32'h24822800;
      105224: inst = 32'h10a00000;
      105225: inst = 32'hca00004;
      105226: inst = 32'h38632800;
      105227: inst = 32'h38842800;
      105228: inst = 32'h10a00001;
      105229: inst = 32'hca09b11;
      105230: inst = 32'h13e00001;
      105231: inst = 32'hfe0d96a;
      105232: inst = 32'h5be00000;
      105233: inst = 32'h8c50000;
      105234: inst = 32'h24612800;
      105235: inst = 32'h10a00000;
      105236: inst = 32'hca00014;
      105237: inst = 32'h24822800;
      105238: inst = 32'h10a00000;
      105239: inst = 32'hca00004;
      105240: inst = 32'h38632800;
      105241: inst = 32'h38842800;
      105242: inst = 32'h10a00001;
      105243: inst = 32'hca09b1f;
      105244: inst = 32'h13e00001;
      105245: inst = 32'hfe0d96a;
      105246: inst = 32'h5be00000;
      105247: inst = 32'h8c50000;
      105248: inst = 32'h24612800;
      105249: inst = 32'h10a00000;
      105250: inst = 32'hca00014;
      105251: inst = 32'h24822800;
      105252: inst = 32'h10a00000;
      105253: inst = 32'hca00004;
      105254: inst = 32'h38632800;
      105255: inst = 32'h38842800;
      105256: inst = 32'h10a00001;
      105257: inst = 32'hca09b2d;
      105258: inst = 32'h13e00001;
      105259: inst = 32'hfe0d96a;
      105260: inst = 32'h5be00000;
      105261: inst = 32'h8c50000;
      105262: inst = 32'h24612800;
      105263: inst = 32'h10a00000;
      105264: inst = 32'hca00014;
      105265: inst = 32'h24822800;
      105266: inst = 32'h10a00000;
      105267: inst = 32'hca00004;
      105268: inst = 32'h38632800;
      105269: inst = 32'h38842800;
      105270: inst = 32'h10a00001;
      105271: inst = 32'hca09b3b;
      105272: inst = 32'h13e00001;
      105273: inst = 32'hfe0d96a;
      105274: inst = 32'h5be00000;
      105275: inst = 32'h8c50000;
      105276: inst = 32'h24612800;
      105277: inst = 32'h10a00000;
      105278: inst = 32'hca00014;
      105279: inst = 32'h24822800;
      105280: inst = 32'h10a00000;
      105281: inst = 32'hca00004;
      105282: inst = 32'h38632800;
      105283: inst = 32'h38842800;
      105284: inst = 32'h10a00001;
      105285: inst = 32'hca09b49;
      105286: inst = 32'h13e00001;
      105287: inst = 32'hfe0d96a;
      105288: inst = 32'h5be00000;
      105289: inst = 32'h8c50000;
      105290: inst = 32'h24612800;
      105291: inst = 32'h10a00000;
      105292: inst = 32'hca00014;
      105293: inst = 32'h24822800;
      105294: inst = 32'h10a00000;
      105295: inst = 32'hca00004;
      105296: inst = 32'h38632800;
      105297: inst = 32'h38842800;
      105298: inst = 32'h10a00001;
      105299: inst = 32'hca09b57;
      105300: inst = 32'h13e00001;
      105301: inst = 32'hfe0d96a;
      105302: inst = 32'h5be00000;
      105303: inst = 32'h8c50000;
      105304: inst = 32'h24612800;
      105305: inst = 32'h10a00000;
      105306: inst = 32'hca00014;
      105307: inst = 32'h24822800;
      105308: inst = 32'h10a00000;
      105309: inst = 32'hca00004;
      105310: inst = 32'h38632800;
      105311: inst = 32'h38842800;
      105312: inst = 32'h10a00001;
      105313: inst = 32'hca09b65;
      105314: inst = 32'h13e00001;
      105315: inst = 32'hfe0d96a;
      105316: inst = 32'h5be00000;
      105317: inst = 32'h8c50000;
      105318: inst = 32'h24612800;
      105319: inst = 32'h10a00000;
      105320: inst = 32'hca00014;
      105321: inst = 32'h24822800;
      105322: inst = 32'h10a00000;
      105323: inst = 32'hca00004;
      105324: inst = 32'h38632800;
      105325: inst = 32'h38842800;
      105326: inst = 32'h10a00001;
      105327: inst = 32'hca09b73;
      105328: inst = 32'h13e00001;
      105329: inst = 32'hfe0d96a;
      105330: inst = 32'h5be00000;
      105331: inst = 32'h8c50000;
      105332: inst = 32'h24612800;
      105333: inst = 32'h10a00000;
      105334: inst = 32'hca00014;
      105335: inst = 32'h24822800;
      105336: inst = 32'h10a00000;
      105337: inst = 32'hca00004;
      105338: inst = 32'h38632800;
      105339: inst = 32'h38842800;
      105340: inst = 32'h10a00001;
      105341: inst = 32'hca09b81;
      105342: inst = 32'h13e00001;
      105343: inst = 32'hfe0d96a;
      105344: inst = 32'h5be00000;
      105345: inst = 32'h8c50000;
      105346: inst = 32'h24612800;
      105347: inst = 32'h10a00000;
      105348: inst = 32'hca00014;
      105349: inst = 32'h24822800;
      105350: inst = 32'h10a00000;
      105351: inst = 32'hca00004;
      105352: inst = 32'h38632800;
      105353: inst = 32'h38842800;
      105354: inst = 32'h10a00001;
      105355: inst = 32'hca09b8f;
      105356: inst = 32'h13e00001;
      105357: inst = 32'hfe0d96a;
      105358: inst = 32'h5be00000;
      105359: inst = 32'h8c50000;
      105360: inst = 32'h24612800;
      105361: inst = 32'h10a00000;
      105362: inst = 32'hca00014;
      105363: inst = 32'h24822800;
      105364: inst = 32'h10a00000;
      105365: inst = 32'hca00004;
      105366: inst = 32'h38632800;
      105367: inst = 32'h38842800;
      105368: inst = 32'h10a00001;
      105369: inst = 32'hca09b9d;
      105370: inst = 32'h13e00001;
      105371: inst = 32'hfe0d96a;
      105372: inst = 32'h5be00000;
      105373: inst = 32'h8c50000;
      105374: inst = 32'h24612800;
      105375: inst = 32'h10a00000;
      105376: inst = 32'hca00014;
      105377: inst = 32'h24822800;
      105378: inst = 32'h10a00000;
      105379: inst = 32'hca00004;
      105380: inst = 32'h38632800;
      105381: inst = 32'h38842800;
      105382: inst = 32'h10a00001;
      105383: inst = 32'hca09bab;
      105384: inst = 32'h13e00001;
      105385: inst = 32'hfe0d96a;
      105386: inst = 32'h5be00000;
      105387: inst = 32'h8c50000;
      105388: inst = 32'h24612800;
      105389: inst = 32'h10a00000;
      105390: inst = 32'hca00014;
      105391: inst = 32'h24822800;
      105392: inst = 32'h10a00000;
      105393: inst = 32'hca00004;
      105394: inst = 32'h38632800;
      105395: inst = 32'h38842800;
      105396: inst = 32'h10a00001;
      105397: inst = 32'hca09bb9;
      105398: inst = 32'h13e00001;
      105399: inst = 32'hfe0d96a;
      105400: inst = 32'h5be00000;
      105401: inst = 32'h8c50000;
      105402: inst = 32'h24612800;
      105403: inst = 32'h10a00000;
      105404: inst = 32'hca00014;
      105405: inst = 32'h24822800;
      105406: inst = 32'h10a00000;
      105407: inst = 32'hca00004;
      105408: inst = 32'h38632800;
      105409: inst = 32'h38842800;
      105410: inst = 32'h10a00001;
      105411: inst = 32'hca09bc7;
      105412: inst = 32'h13e00001;
      105413: inst = 32'hfe0d96a;
      105414: inst = 32'h5be00000;
      105415: inst = 32'h8c50000;
      105416: inst = 32'h24612800;
      105417: inst = 32'h10a00000;
      105418: inst = 32'hca00014;
      105419: inst = 32'h24822800;
      105420: inst = 32'h10a00000;
      105421: inst = 32'hca00004;
      105422: inst = 32'h38632800;
      105423: inst = 32'h38842800;
      105424: inst = 32'h10a00001;
      105425: inst = 32'hca09bd5;
      105426: inst = 32'h13e00001;
      105427: inst = 32'hfe0d96a;
      105428: inst = 32'h5be00000;
      105429: inst = 32'h8c50000;
      105430: inst = 32'h24612800;
      105431: inst = 32'h10a00000;
      105432: inst = 32'hca00014;
      105433: inst = 32'h24822800;
      105434: inst = 32'h10a00000;
      105435: inst = 32'hca00004;
      105436: inst = 32'h38632800;
      105437: inst = 32'h38842800;
      105438: inst = 32'h10a00001;
      105439: inst = 32'hca09be3;
      105440: inst = 32'h13e00001;
      105441: inst = 32'hfe0d96a;
      105442: inst = 32'h5be00000;
      105443: inst = 32'h8c50000;
      105444: inst = 32'h24612800;
      105445: inst = 32'h10a00000;
      105446: inst = 32'hca00014;
      105447: inst = 32'h24822800;
      105448: inst = 32'h10a00000;
      105449: inst = 32'hca00004;
      105450: inst = 32'h38632800;
      105451: inst = 32'h38842800;
      105452: inst = 32'h10a00001;
      105453: inst = 32'hca09bf1;
      105454: inst = 32'h13e00001;
      105455: inst = 32'hfe0d96a;
      105456: inst = 32'h5be00000;
      105457: inst = 32'h8c50000;
      105458: inst = 32'h24612800;
      105459: inst = 32'h10a00000;
      105460: inst = 32'hca00014;
      105461: inst = 32'h24822800;
      105462: inst = 32'h10a00000;
      105463: inst = 32'hca00004;
      105464: inst = 32'h38632800;
      105465: inst = 32'h38842800;
      105466: inst = 32'h10a00001;
      105467: inst = 32'hca09bff;
      105468: inst = 32'h13e00001;
      105469: inst = 32'hfe0d96a;
      105470: inst = 32'h5be00000;
      105471: inst = 32'h8c50000;
      105472: inst = 32'h24612800;
      105473: inst = 32'h10a00000;
      105474: inst = 32'hca00014;
      105475: inst = 32'h24822800;
      105476: inst = 32'h10a00000;
      105477: inst = 32'hca00004;
      105478: inst = 32'h38632800;
      105479: inst = 32'h38842800;
      105480: inst = 32'h10a00001;
      105481: inst = 32'hca09c0d;
      105482: inst = 32'h13e00001;
      105483: inst = 32'hfe0d96a;
      105484: inst = 32'h5be00000;
      105485: inst = 32'h8c50000;
      105486: inst = 32'h24612800;
      105487: inst = 32'h10a00000;
      105488: inst = 32'hca00014;
      105489: inst = 32'h24822800;
      105490: inst = 32'h10a00000;
      105491: inst = 32'hca00004;
      105492: inst = 32'h38632800;
      105493: inst = 32'h38842800;
      105494: inst = 32'h10a00001;
      105495: inst = 32'hca09c1b;
      105496: inst = 32'h13e00001;
      105497: inst = 32'hfe0d96a;
      105498: inst = 32'h5be00000;
      105499: inst = 32'h8c50000;
      105500: inst = 32'h24612800;
      105501: inst = 32'h10a00000;
      105502: inst = 32'hca00014;
      105503: inst = 32'h24822800;
      105504: inst = 32'h10a00000;
      105505: inst = 32'hca00004;
      105506: inst = 32'h38632800;
      105507: inst = 32'h38842800;
      105508: inst = 32'h10a00001;
      105509: inst = 32'hca09c29;
      105510: inst = 32'h13e00001;
      105511: inst = 32'hfe0d96a;
      105512: inst = 32'h5be00000;
      105513: inst = 32'h8c50000;
      105514: inst = 32'h24612800;
      105515: inst = 32'h10a00000;
      105516: inst = 32'hca00014;
      105517: inst = 32'h24822800;
      105518: inst = 32'h10a00000;
      105519: inst = 32'hca00004;
      105520: inst = 32'h38632800;
      105521: inst = 32'h38842800;
      105522: inst = 32'h10a00001;
      105523: inst = 32'hca09c37;
      105524: inst = 32'h13e00001;
      105525: inst = 32'hfe0d96a;
      105526: inst = 32'h5be00000;
      105527: inst = 32'h8c50000;
      105528: inst = 32'h24612800;
      105529: inst = 32'h10a00000;
      105530: inst = 32'hca00014;
      105531: inst = 32'h24822800;
      105532: inst = 32'h10a00000;
      105533: inst = 32'hca00004;
      105534: inst = 32'h38632800;
      105535: inst = 32'h38842800;
      105536: inst = 32'h10a00001;
      105537: inst = 32'hca09c45;
      105538: inst = 32'h13e00001;
      105539: inst = 32'hfe0d96a;
      105540: inst = 32'h5be00000;
      105541: inst = 32'h8c50000;
      105542: inst = 32'h24612800;
      105543: inst = 32'h10a00000;
      105544: inst = 32'hca00014;
      105545: inst = 32'h24822800;
      105546: inst = 32'h10a00000;
      105547: inst = 32'hca00004;
      105548: inst = 32'h38632800;
      105549: inst = 32'h38842800;
      105550: inst = 32'h10a00001;
      105551: inst = 32'hca09c53;
      105552: inst = 32'h13e00001;
      105553: inst = 32'hfe0d96a;
      105554: inst = 32'h5be00000;
      105555: inst = 32'h8c50000;
      105556: inst = 32'h24612800;
      105557: inst = 32'h10a00000;
      105558: inst = 32'hca00014;
      105559: inst = 32'h24822800;
      105560: inst = 32'h10a00000;
      105561: inst = 32'hca00004;
      105562: inst = 32'h38632800;
      105563: inst = 32'h38842800;
      105564: inst = 32'h10a00001;
      105565: inst = 32'hca09c61;
      105566: inst = 32'h13e00001;
      105567: inst = 32'hfe0d96a;
      105568: inst = 32'h5be00000;
      105569: inst = 32'h8c50000;
      105570: inst = 32'h24612800;
      105571: inst = 32'h10a00000;
      105572: inst = 32'hca00014;
      105573: inst = 32'h24822800;
      105574: inst = 32'h10a00000;
      105575: inst = 32'hca00004;
      105576: inst = 32'h38632800;
      105577: inst = 32'h38842800;
      105578: inst = 32'h10a00001;
      105579: inst = 32'hca09c6f;
      105580: inst = 32'h13e00001;
      105581: inst = 32'hfe0d96a;
      105582: inst = 32'h5be00000;
      105583: inst = 32'h8c50000;
      105584: inst = 32'h24612800;
      105585: inst = 32'h10a00000;
      105586: inst = 32'hca00014;
      105587: inst = 32'h24822800;
      105588: inst = 32'h10a00000;
      105589: inst = 32'hca00004;
      105590: inst = 32'h38632800;
      105591: inst = 32'h38842800;
      105592: inst = 32'h10a00001;
      105593: inst = 32'hca09c7d;
      105594: inst = 32'h13e00001;
      105595: inst = 32'hfe0d96a;
      105596: inst = 32'h5be00000;
      105597: inst = 32'h8c50000;
      105598: inst = 32'h24612800;
      105599: inst = 32'h10a00000;
      105600: inst = 32'hca00014;
      105601: inst = 32'h24822800;
      105602: inst = 32'h10a00000;
      105603: inst = 32'hca00004;
      105604: inst = 32'h38632800;
      105605: inst = 32'h38842800;
      105606: inst = 32'h10a00001;
      105607: inst = 32'hca09c8b;
      105608: inst = 32'h13e00001;
      105609: inst = 32'hfe0d96a;
      105610: inst = 32'h5be00000;
      105611: inst = 32'h8c50000;
      105612: inst = 32'h24612800;
      105613: inst = 32'h10a00000;
      105614: inst = 32'hca00014;
      105615: inst = 32'h24822800;
      105616: inst = 32'h10a00000;
      105617: inst = 32'hca00004;
      105618: inst = 32'h38632800;
      105619: inst = 32'h38842800;
      105620: inst = 32'h10a00001;
      105621: inst = 32'hca09c99;
      105622: inst = 32'h13e00001;
      105623: inst = 32'hfe0d96a;
      105624: inst = 32'h5be00000;
      105625: inst = 32'h8c50000;
      105626: inst = 32'h24612800;
      105627: inst = 32'h10a00000;
      105628: inst = 32'hca00014;
      105629: inst = 32'h24822800;
      105630: inst = 32'h10a00000;
      105631: inst = 32'hca00004;
      105632: inst = 32'h38632800;
      105633: inst = 32'h38842800;
      105634: inst = 32'h10a00001;
      105635: inst = 32'hca09ca7;
      105636: inst = 32'h13e00001;
      105637: inst = 32'hfe0d96a;
      105638: inst = 32'h5be00000;
      105639: inst = 32'h8c50000;
      105640: inst = 32'h24612800;
      105641: inst = 32'h10a00000;
      105642: inst = 32'hca00014;
      105643: inst = 32'h24822800;
      105644: inst = 32'h10a00000;
      105645: inst = 32'hca00004;
      105646: inst = 32'h38632800;
      105647: inst = 32'h38842800;
      105648: inst = 32'h10a00001;
      105649: inst = 32'hca09cb5;
      105650: inst = 32'h13e00001;
      105651: inst = 32'hfe0d96a;
      105652: inst = 32'h5be00000;
      105653: inst = 32'h8c50000;
      105654: inst = 32'h24612800;
      105655: inst = 32'h10a00000;
      105656: inst = 32'hca00014;
      105657: inst = 32'h24822800;
      105658: inst = 32'h10a00000;
      105659: inst = 32'hca00004;
      105660: inst = 32'h38632800;
      105661: inst = 32'h38842800;
      105662: inst = 32'h10a00001;
      105663: inst = 32'hca09cc3;
      105664: inst = 32'h13e00001;
      105665: inst = 32'hfe0d96a;
      105666: inst = 32'h5be00000;
      105667: inst = 32'h8c50000;
      105668: inst = 32'h24612800;
      105669: inst = 32'h10a00000;
      105670: inst = 32'hca00014;
      105671: inst = 32'h24822800;
      105672: inst = 32'h10a00000;
      105673: inst = 32'hca00004;
      105674: inst = 32'h38632800;
      105675: inst = 32'h38842800;
      105676: inst = 32'h10a00001;
      105677: inst = 32'hca09cd1;
      105678: inst = 32'h13e00001;
      105679: inst = 32'hfe0d96a;
      105680: inst = 32'h5be00000;
      105681: inst = 32'h8c50000;
      105682: inst = 32'h24612800;
      105683: inst = 32'h10a00000;
      105684: inst = 32'hca00014;
      105685: inst = 32'h24822800;
      105686: inst = 32'h10a00000;
      105687: inst = 32'hca00004;
      105688: inst = 32'h38632800;
      105689: inst = 32'h38842800;
      105690: inst = 32'h10a00001;
      105691: inst = 32'hca09cdf;
      105692: inst = 32'h13e00001;
      105693: inst = 32'hfe0d96a;
      105694: inst = 32'h5be00000;
      105695: inst = 32'h8c50000;
      105696: inst = 32'h24612800;
      105697: inst = 32'h10a00000;
      105698: inst = 32'hca00014;
      105699: inst = 32'h24822800;
      105700: inst = 32'h10a00000;
      105701: inst = 32'hca00004;
      105702: inst = 32'h38632800;
      105703: inst = 32'h38842800;
      105704: inst = 32'h10a00001;
      105705: inst = 32'hca09ced;
      105706: inst = 32'h13e00001;
      105707: inst = 32'hfe0d96a;
      105708: inst = 32'h5be00000;
      105709: inst = 32'h8c50000;
      105710: inst = 32'h24612800;
      105711: inst = 32'h10a00000;
      105712: inst = 32'hca00014;
      105713: inst = 32'h24822800;
      105714: inst = 32'h10a00000;
      105715: inst = 32'hca00004;
      105716: inst = 32'h38632800;
      105717: inst = 32'h38842800;
      105718: inst = 32'h10a00001;
      105719: inst = 32'hca09cfb;
      105720: inst = 32'h13e00001;
      105721: inst = 32'hfe0d96a;
      105722: inst = 32'h5be00000;
      105723: inst = 32'h8c50000;
      105724: inst = 32'h24612800;
      105725: inst = 32'h10a00000;
      105726: inst = 32'hca00014;
      105727: inst = 32'h24822800;
      105728: inst = 32'h10a00000;
      105729: inst = 32'hca00004;
      105730: inst = 32'h38632800;
      105731: inst = 32'h38842800;
      105732: inst = 32'h10a00001;
      105733: inst = 32'hca09d09;
      105734: inst = 32'h13e00001;
      105735: inst = 32'hfe0d96a;
      105736: inst = 32'h5be00000;
      105737: inst = 32'h8c50000;
      105738: inst = 32'h24612800;
      105739: inst = 32'h10a00000;
      105740: inst = 32'hca00014;
      105741: inst = 32'h24822800;
      105742: inst = 32'h10a00000;
      105743: inst = 32'hca00004;
      105744: inst = 32'h38632800;
      105745: inst = 32'h38842800;
      105746: inst = 32'h10a00001;
      105747: inst = 32'hca09d17;
      105748: inst = 32'h13e00001;
      105749: inst = 32'hfe0d96a;
      105750: inst = 32'h5be00000;
      105751: inst = 32'h8c50000;
      105752: inst = 32'h24612800;
      105753: inst = 32'h10a00000;
      105754: inst = 32'hca00014;
      105755: inst = 32'h24822800;
      105756: inst = 32'h10a00000;
      105757: inst = 32'hca00004;
      105758: inst = 32'h38632800;
      105759: inst = 32'h38842800;
      105760: inst = 32'h10a00001;
      105761: inst = 32'hca09d25;
      105762: inst = 32'h13e00001;
      105763: inst = 32'hfe0d96a;
      105764: inst = 32'h5be00000;
      105765: inst = 32'h8c50000;
      105766: inst = 32'h24612800;
      105767: inst = 32'h10a00000;
      105768: inst = 32'hca00014;
      105769: inst = 32'h24822800;
      105770: inst = 32'h10a00000;
      105771: inst = 32'hca00004;
      105772: inst = 32'h38632800;
      105773: inst = 32'h38842800;
      105774: inst = 32'h10a00001;
      105775: inst = 32'hca09d33;
      105776: inst = 32'h13e00001;
      105777: inst = 32'hfe0d96a;
      105778: inst = 32'h5be00000;
      105779: inst = 32'h8c50000;
      105780: inst = 32'h24612800;
      105781: inst = 32'h10a00000;
      105782: inst = 32'hca00014;
      105783: inst = 32'h24822800;
      105784: inst = 32'h10a00000;
      105785: inst = 32'hca00004;
      105786: inst = 32'h38632800;
      105787: inst = 32'h38842800;
      105788: inst = 32'h10a00001;
      105789: inst = 32'hca09d41;
      105790: inst = 32'h13e00001;
      105791: inst = 32'hfe0d96a;
      105792: inst = 32'h5be00000;
      105793: inst = 32'h8c50000;
      105794: inst = 32'h24612800;
      105795: inst = 32'h10a00000;
      105796: inst = 32'hca00014;
      105797: inst = 32'h24822800;
      105798: inst = 32'h10a00000;
      105799: inst = 32'hca00004;
      105800: inst = 32'h38632800;
      105801: inst = 32'h38842800;
      105802: inst = 32'h10a00001;
      105803: inst = 32'hca09d4f;
      105804: inst = 32'h13e00001;
      105805: inst = 32'hfe0d96a;
      105806: inst = 32'h5be00000;
      105807: inst = 32'h8c50000;
      105808: inst = 32'h24612800;
      105809: inst = 32'h10a00000;
      105810: inst = 32'hca00014;
      105811: inst = 32'h24822800;
      105812: inst = 32'h10a00000;
      105813: inst = 32'hca00004;
      105814: inst = 32'h38632800;
      105815: inst = 32'h38842800;
      105816: inst = 32'h10a00001;
      105817: inst = 32'hca09d5d;
      105818: inst = 32'h13e00001;
      105819: inst = 32'hfe0d96a;
      105820: inst = 32'h5be00000;
      105821: inst = 32'h8c50000;
      105822: inst = 32'h24612800;
      105823: inst = 32'h10a00000;
      105824: inst = 32'hca00014;
      105825: inst = 32'h24822800;
      105826: inst = 32'h10a00000;
      105827: inst = 32'hca00004;
      105828: inst = 32'h38632800;
      105829: inst = 32'h38842800;
      105830: inst = 32'h10a00001;
      105831: inst = 32'hca09d6b;
      105832: inst = 32'h13e00001;
      105833: inst = 32'hfe0d96a;
      105834: inst = 32'h5be00000;
      105835: inst = 32'h8c50000;
      105836: inst = 32'h24612800;
      105837: inst = 32'h10a00000;
      105838: inst = 32'hca00014;
      105839: inst = 32'h24822800;
      105840: inst = 32'h10a00000;
      105841: inst = 32'hca00004;
      105842: inst = 32'h38632800;
      105843: inst = 32'h38842800;
      105844: inst = 32'h10a00001;
      105845: inst = 32'hca09d79;
      105846: inst = 32'h13e00001;
      105847: inst = 32'hfe0d96a;
      105848: inst = 32'h5be00000;
      105849: inst = 32'h8c50000;
      105850: inst = 32'h24612800;
      105851: inst = 32'h10a00000;
      105852: inst = 32'hca00014;
      105853: inst = 32'h24822800;
      105854: inst = 32'h10a00000;
      105855: inst = 32'hca00004;
      105856: inst = 32'h38632800;
      105857: inst = 32'h38842800;
      105858: inst = 32'h10a00001;
      105859: inst = 32'hca09d87;
      105860: inst = 32'h13e00001;
      105861: inst = 32'hfe0d96a;
      105862: inst = 32'h5be00000;
      105863: inst = 32'h8c50000;
      105864: inst = 32'h24612800;
      105865: inst = 32'h10a00000;
      105866: inst = 32'hca00014;
      105867: inst = 32'h24822800;
      105868: inst = 32'h10a00000;
      105869: inst = 32'hca00004;
      105870: inst = 32'h38632800;
      105871: inst = 32'h38842800;
      105872: inst = 32'h10a00001;
      105873: inst = 32'hca09d95;
      105874: inst = 32'h13e00001;
      105875: inst = 32'hfe0d96a;
      105876: inst = 32'h5be00000;
      105877: inst = 32'h8c50000;
      105878: inst = 32'h24612800;
      105879: inst = 32'h10a00000;
      105880: inst = 32'hca00014;
      105881: inst = 32'h24822800;
      105882: inst = 32'h10a00000;
      105883: inst = 32'hca00004;
      105884: inst = 32'h38632800;
      105885: inst = 32'h38842800;
      105886: inst = 32'h10a00001;
      105887: inst = 32'hca09da3;
      105888: inst = 32'h13e00001;
      105889: inst = 32'hfe0d96a;
      105890: inst = 32'h5be00000;
      105891: inst = 32'h8c50000;
      105892: inst = 32'h24612800;
      105893: inst = 32'h10a00000;
      105894: inst = 32'hca00014;
      105895: inst = 32'h24822800;
      105896: inst = 32'h10a00000;
      105897: inst = 32'hca00004;
      105898: inst = 32'h38632800;
      105899: inst = 32'h38842800;
      105900: inst = 32'h10a00001;
      105901: inst = 32'hca09db1;
      105902: inst = 32'h13e00001;
      105903: inst = 32'hfe0d96a;
      105904: inst = 32'h5be00000;
      105905: inst = 32'h8c50000;
      105906: inst = 32'h24612800;
      105907: inst = 32'h10a00000;
      105908: inst = 32'hca00014;
      105909: inst = 32'h24822800;
      105910: inst = 32'h10a00000;
      105911: inst = 32'hca00004;
      105912: inst = 32'h38632800;
      105913: inst = 32'h38842800;
      105914: inst = 32'h10a00001;
      105915: inst = 32'hca09dbf;
      105916: inst = 32'h13e00001;
      105917: inst = 32'hfe0d96a;
      105918: inst = 32'h5be00000;
      105919: inst = 32'h8c50000;
      105920: inst = 32'h24612800;
      105921: inst = 32'h10a00000;
      105922: inst = 32'hca00014;
      105923: inst = 32'h24822800;
      105924: inst = 32'h10a00000;
      105925: inst = 32'hca00004;
      105926: inst = 32'h38632800;
      105927: inst = 32'h38842800;
      105928: inst = 32'h10a00001;
      105929: inst = 32'hca09dcd;
      105930: inst = 32'h13e00001;
      105931: inst = 32'hfe0d96a;
      105932: inst = 32'h5be00000;
      105933: inst = 32'h8c50000;
      105934: inst = 32'h24612800;
      105935: inst = 32'h10a00000;
      105936: inst = 32'hca00014;
      105937: inst = 32'h24822800;
      105938: inst = 32'h10a00000;
      105939: inst = 32'hca00004;
      105940: inst = 32'h38632800;
      105941: inst = 32'h38842800;
      105942: inst = 32'h10a00001;
      105943: inst = 32'hca09ddb;
      105944: inst = 32'h13e00001;
      105945: inst = 32'hfe0d96a;
      105946: inst = 32'h5be00000;
      105947: inst = 32'h8c50000;
      105948: inst = 32'h24612800;
      105949: inst = 32'h10a00000;
      105950: inst = 32'hca00014;
      105951: inst = 32'h24822800;
      105952: inst = 32'h10a00000;
      105953: inst = 32'hca00004;
      105954: inst = 32'h38632800;
      105955: inst = 32'h38842800;
      105956: inst = 32'h10a00001;
      105957: inst = 32'hca09de9;
      105958: inst = 32'h13e00001;
      105959: inst = 32'hfe0d96a;
      105960: inst = 32'h5be00000;
      105961: inst = 32'h8c50000;
      105962: inst = 32'h24612800;
      105963: inst = 32'h10a00000;
      105964: inst = 32'hca00014;
      105965: inst = 32'h24822800;
      105966: inst = 32'h10a00000;
      105967: inst = 32'hca00004;
      105968: inst = 32'h38632800;
      105969: inst = 32'h38842800;
      105970: inst = 32'h10a00001;
      105971: inst = 32'hca09df7;
      105972: inst = 32'h13e00001;
      105973: inst = 32'hfe0d96a;
      105974: inst = 32'h5be00000;
      105975: inst = 32'h8c50000;
      105976: inst = 32'h24612800;
      105977: inst = 32'h10a00000;
      105978: inst = 32'hca00014;
      105979: inst = 32'h24822800;
      105980: inst = 32'h10a00000;
      105981: inst = 32'hca00004;
      105982: inst = 32'h38632800;
      105983: inst = 32'h38842800;
      105984: inst = 32'h10a00001;
      105985: inst = 32'hca09e05;
      105986: inst = 32'h13e00001;
      105987: inst = 32'hfe0d96a;
      105988: inst = 32'h5be00000;
      105989: inst = 32'h8c50000;
      105990: inst = 32'h24612800;
      105991: inst = 32'h10a00000;
      105992: inst = 32'hca00014;
      105993: inst = 32'h24822800;
      105994: inst = 32'h10a00000;
      105995: inst = 32'hca00004;
      105996: inst = 32'h38632800;
      105997: inst = 32'h38842800;
      105998: inst = 32'h10a00001;
      105999: inst = 32'hca09e13;
      106000: inst = 32'h13e00001;
      106001: inst = 32'hfe0d96a;
      106002: inst = 32'h5be00000;
      106003: inst = 32'h8c50000;
      106004: inst = 32'h24612800;
      106005: inst = 32'h10a00000;
      106006: inst = 32'hca00014;
      106007: inst = 32'h24822800;
      106008: inst = 32'h10a00000;
      106009: inst = 32'hca00004;
      106010: inst = 32'h38632800;
      106011: inst = 32'h38842800;
      106012: inst = 32'h10a00001;
      106013: inst = 32'hca09e21;
      106014: inst = 32'h13e00001;
      106015: inst = 32'hfe0d96a;
      106016: inst = 32'h5be00000;
      106017: inst = 32'h8c50000;
      106018: inst = 32'h24612800;
      106019: inst = 32'h10a00000;
      106020: inst = 32'hca00014;
      106021: inst = 32'h24822800;
      106022: inst = 32'h10a00000;
      106023: inst = 32'hca00004;
      106024: inst = 32'h38632800;
      106025: inst = 32'h38842800;
      106026: inst = 32'h10a00001;
      106027: inst = 32'hca09e2f;
      106028: inst = 32'h13e00001;
      106029: inst = 32'hfe0d96a;
      106030: inst = 32'h5be00000;
      106031: inst = 32'h8c50000;
      106032: inst = 32'h24612800;
      106033: inst = 32'h10a00000;
      106034: inst = 32'hca00014;
      106035: inst = 32'h24822800;
      106036: inst = 32'h10a00000;
      106037: inst = 32'hca00004;
      106038: inst = 32'h38632800;
      106039: inst = 32'h38842800;
      106040: inst = 32'h10a00001;
      106041: inst = 32'hca09e3d;
      106042: inst = 32'h13e00001;
      106043: inst = 32'hfe0d96a;
      106044: inst = 32'h5be00000;
      106045: inst = 32'h8c50000;
      106046: inst = 32'h24612800;
      106047: inst = 32'h10a00000;
      106048: inst = 32'hca00014;
      106049: inst = 32'h24822800;
      106050: inst = 32'h10a00000;
      106051: inst = 32'hca00004;
      106052: inst = 32'h38632800;
      106053: inst = 32'h38842800;
      106054: inst = 32'h10a00001;
      106055: inst = 32'hca09e4b;
      106056: inst = 32'h13e00001;
      106057: inst = 32'hfe0d96a;
      106058: inst = 32'h5be00000;
      106059: inst = 32'h8c50000;
      106060: inst = 32'h24612800;
      106061: inst = 32'h10a00000;
      106062: inst = 32'hca00014;
      106063: inst = 32'h24822800;
      106064: inst = 32'h10a00000;
      106065: inst = 32'hca00004;
      106066: inst = 32'h38632800;
      106067: inst = 32'h38842800;
      106068: inst = 32'h10a00001;
      106069: inst = 32'hca09e59;
      106070: inst = 32'h13e00001;
      106071: inst = 32'hfe0d96a;
      106072: inst = 32'h5be00000;
      106073: inst = 32'h8c50000;
      106074: inst = 32'h24612800;
      106075: inst = 32'h10a00000;
      106076: inst = 32'hca00014;
      106077: inst = 32'h24822800;
      106078: inst = 32'h10a00000;
      106079: inst = 32'hca00004;
      106080: inst = 32'h38632800;
      106081: inst = 32'h38842800;
      106082: inst = 32'h10a00001;
      106083: inst = 32'hca09e67;
      106084: inst = 32'h13e00001;
      106085: inst = 32'hfe0d96a;
      106086: inst = 32'h5be00000;
      106087: inst = 32'h8c50000;
      106088: inst = 32'h24612800;
      106089: inst = 32'h10a00000;
      106090: inst = 32'hca00014;
      106091: inst = 32'h24822800;
      106092: inst = 32'h10a00000;
      106093: inst = 32'hca00004;
      106094: inst = 32'h38632800;
      106095: inst = 32'h38842800;
      106096: inst = 32'h10a00001;
      106097: inst = 32'hca09e75;
      106098: inst = 32'h13e00001;
      106099: inst = 32'hfe0d96a;
      106100: inst = 32'h5be00000;
      106101: inst = 32'h8c50000;
      106102: inst = 32'h24612800;
      106103: inst = 32'h10a00000;
      106104: inst = 32'hca00014;
      106105: inst = 32'h24822800;
      106106: inst = 32'h10a00000;
      106107: inst = 32'hca00004;
      106108: inst = 32'h38632800;
      106109: inst = 32'h38842800;
      106110: inst = 32'h10a00001;
      106111: inst = 32'hca09e83;
      106112: inst = 32'h13e00001;
      106113: inst = 32'hfe0d96a;
      106114: inst = 32'h5be00000;
      106115: inst = 32'h8c50000;
      106116: inst = 32'h24612800;
      106117: inst = 32'h10a00000;
      106118: inst = 32'hca00014;
      106119: inst = 32'h24822800;
      106120: inst = 32'h10a00000;
      106121: inst = 32'hca00004;
      106122: inst = 32'h38632800;
      106123: inst = 32'h38842800;
      106124: inst = 32'h10a00001;
      106125: inst = 32'hca09e91;
      106126: inst = 32'h13e00001;
      106127: inst = 32'hfe0d96a;
      106128: inst = 32'h5be00000;
      106129: inst = 32'h8c50000;
      106130: inst = 32'h24612800;
      106131: inst = 32'h10a00000;
      106132: inst = 32'hca00014;
      106133: inst = 32'h24822800;
      106134: inst = 32'h10a00000;
      106135: inst = 32'hca00004;
      106136: inst = 32'h38632800;
      106137: inst = 32'h38842800;
      106138: inst = 32'h10a00001;
      106139: inst = 32'hca09e9f;
      106140: inst = 32'h13e00001;
      106141: inst = 32'hfe0d96a;
      106142: inst = 32'h5be00000;
      106143: inst = 32'h8c50000;
      106144: inst = 32'h24612800;
      106145: inst = 32'h10a00000;
      106146: inst = 32'hca00014;
      106147: inst = 32'h24822800;
      106148: inst = 32'h10a00000;
      106149: inst = 32'hca00004;
      106150: inst = 32'h38632800;
      106151: inst = 32'h38842800;
      106152: inst = 32'h10a00001;
      106153: inst = 32'hca09ead;
      106154: inst = 32'h13e00001;
      106155: inst = 32'hfe0d96a;
      106156: inst = 32'h5be00000;
      106157: inst = 32'h8c50000;
      106158: inst = 32'h24612800;
      106159: inst = 32'h10a00000;
      106160: inst = 32'hca00014;
      106161: inst = 32'h24822800;
      106162: inst = 32'h10a00000;
      106163: inst = 32'hca00004;
      106164: inst = 32'h38632800;
      106165: inst = 32'h38842800;
      106166: inst = 32'h10a00001;
      106167: inst = 32'hca09ebb;
      106168: inst = 32'h13e00001;
      106169: inst = 32'hfe0d96a;
      106170: inst = 32'h5be00000;
      106171: inst = 32'h8c50000;
      106172: inst = 32'h24612800;
      106173: inst = 32'h10a00000;
      106174: inst = 32'hca00014;
      106175: inst = 32'h24822800;
      106176: inst = 32'h10a00000;
      106177: inst = 32'hca00004;
      106178: inst = 32'h38632800;
      106179: inst = 32'h38842800;
      106180: inst = 32'h10a00001;
      106181: inst = 32'hca09ec9;
      106182: inst = 32'h13e00001;
      106183: inst = 32'hfe0d96a;
      106184: inst = 32'h5be00000;
      106185: inst = 32'h8c50000;
      106186: inst = 32'h24612800;
      106187: inst = 32'h10a00000;
      106188: inst = 32'hca00014;
      106189: inst = 32'h24822800;
      106190: inst = 32'h10a00000;
      106191: inst = 32'hca00004;
      106192: inst = 32'h38632800;
      106193: inst = 32'h38842800;
      106194: inst = 32'h10a00001;
      106195: inst = 32'hca09ed7;
      106196: inst = 32'h13e00001;
      106197: inst = 32'hfe0d96a;
      106198: inst = 32'h5be00000;
      106199: inst = 32'h8c50000;
      106200: inst = 32'h24612800;
      106201: inst = 32'h10a00000;
      106202: inst = 32'hca00014;
      106203: inst = 32'h24822800;
      106204: inst = 32'h10a00000;
      106205: inst = 32'hca00004;
      106206: inst = 32'h38632800;
      106207: inst = 32'h38842800;
      106208: inst = 32'h10a00001;
      106209: inst = 32'hca09ee5;
      106210: inst = 32'h13e00001;
      106211: inst = 32'hfe0d96a;
      106212: inst = 32'h5be00000;
      106213: inst = 32'h8c50000;
      106214: inst = 32'h24612800;
      106215: inst = 32'h10a00000;
      106216: inst = 32'hca00014;
      106217: inst = 32'h24822800;
      106218: inst = 32'h10a00000;
      106219: inst = 32'hca00004;
      106220: inst = 32'h38632800;
      106221: inst = 32'h38842800;
      106222: inst = 32'h10a00001;
      106223: inst = 32'hca09ef3;
      106224: inst = 32'h13e00001;
      106225: inst = 32'hfe0d96a;
      106226: inst = 32'h5be00000;
      106227: inst = 32'h8c50000;
      106228: inst = 32'h24612800;
      106229: inst = 32'h10a00000;
      106230: inst = 32'hca00014;
      106231: inst = 32'h24822800;
      106232: inst = 32'h10a00000;
      106233: inst = 32'hca00004;
      106234: inst = 32'h38632800;
      106235: inst = 32'h38842800;
      106236: inst = 32'h10a00001;
      106237: inst = 32'hca09f01;
      106238: inst = 32'h13e00001;
      106239: inst = 32'hfe0d96a;
      106240: inst = 32'h5be00000;
      106241: inst = 32'h8c50000;
      106242: inst = 32'h24612800;
      106243: inst = 32'h10a00000;
      106244: inst = 32'hca00014;
      106245: inst = 32'h24822800;
      106246: inst = 32'h10a00000;
      106247: inst = 32'hca00004;
      106248: inst = 32'h38632800;
      106249: inst = 32'h38842800;
      106250: inst = 32'h10a00001;
      106251: inst = 32'hca09f0f;
      106252: inst = 32'h13e00001;
      106253: inst = 32'hfe0d96a;
      106254: inst = 32'h5be00000;
      106255: inst = 32'h8c50000;
      106256: inst = 32'h24612800;
      106257: inst = 32'h10a00000;
      106258: inst = 32'hca00014;
      106259: inst = 32'h24822800;
      106260: inst = 32'h10a00000;
      106261: inst = 32'hca00004;
      106262: inst = 32'h38632800;
      106263: inst = 32'h38842800;
      106264: inst = 32'h10a00001;
      106265: inst = 32'hca09f1d;
      106266: inst = 32'h13e00001;
      106267: inst = 32'hfe0d96a;
      106268: inst = 32'h5be00000;
      106269: inst = 32'h8c50000;
      106270: inst = 32'h24612800;
      106271: inst = 32'h10a00000;
      106272: inst = 32'hca00014;
      106273: inst = 32'h24822800;
      106274: inst = 32'h10a00000;
      106275: inst = 32'hca00004;
      106276: inst = 32'h38632800;
      106277: inst = 32'h38842800;
      106278: inst = 32'h10a00001;
      106279: inst = 32'hca09f2b;
      106280: inst = 32'h13e00001;
      106281: inst = 32'hfe0d96a;
      106282: inst = 32'h5be00000;
      106283: inst = 32'h8c50000;
      106284: inst = 32'h24612800;
      106285: inst = 32'h10a00000;
      106286: inst = 32'hca00014;
      106287: inst = 32'h24822800;
      106288: inst = 32'h10a00000;
      106289: inst = 32'hca00004;
      106290: inst = 32'h38632800;
      106291: inst = 32'h38842800;
      106292: inst = 32'h10a00001;
      106293: inst = 32'hca09f39;
      106294: inst = 32'h13e00001;
      106295: inst = 32'hfe0d96a;
      106296: inst = 32'h5be00000;
      106297: inst = 32'h8c50000;
      106298: inst = 32'h24612800;
      106299: inst = 32'h10a00000;
      106300: inst = 32'hca00014;
      106301: inst = 32'h24822800;
      106302: inst = 32'h10a00000;
      106303: inst = 32'hca00004;
      106304: inst = 32'h38632800;
      106305: inst = 32'h38842800;
      106306: inst = 32'h10a00001;
      106307: inst = 32'hca09f47;
      106308: inst = 32'h13e00001;
      106309: inst = 32'hfe0d96a;
      106310: inst = 32'h5be00000;
      106311: inst = 32'h8c50000;
      106312: inst = 32'h24612800;
      106313: inst = 32'h10a00000;
      106314: inst = 32'hca00014;
      106315: inst = 32'h24822800;
      106316: inst = 32'h10a00000;
      106317: inst = 32'hca00004;
      106318: inst = 32'h38632800;
      106319: inst = 32'h38842800;
      106320: inst = 32'h10a00001;
      106321: inst = 32'hca09f55;
      106322: inst = 32'h13e00001;
      106323: inst = 32'hfe0d96a;
      106324: inst = 32'h5be00000;
      106325: inst = 32'h8c50000;
      106326: inst = 32'h24612800;
      106327: inst = 32'h10a00000;
      106328: inst = 32'hca00014;
      106329: inst = 32'h24822800;
      106330: inst = 32'h10a00000;
      106331: inst = 32'hca00004;
      106332: inst = 32'h38632800;
      106333: inst = 32'h38842800;
      106334: inst = 32'h10a00001;
      106335: inst = 32'hca09f63;
      106336: inst = 32'h13e00001;
      106337: inst = 32'hfe0d96a;
      106338: inst = 32'h5be00000;
      106339: inst = 32'h8c50000;
      106340: inst = 32'h24612800;
      106341: inst = 32'h10a00000;
      106342: inst = 32'hca00014;
      106343: inst = 32'h24822800;
      106344: inst = 32'h10a00000;
      106345: inst = 32'hca00004;
      106346: inst = 32'h38632800;
      106347: inst = 32'h38842800;
      106348: inst = 32'h10a00001;
      106349: inst = 32'hca09f71;
      106350: inst = 32'h13e00001;
      106351: inst = 32'hfe0d96a;
      106352: inst = 32'h5be00000;
      106353: inst = 32'h8c50000;
      106354: inst = 32'h24612800;
      106355: inst = 32'h10a00000;
      106356: inst = 32'hca00014;
      106357: inst = 32'h24822800;
      106358: inst = 32'h10a00000;
      106359: inst = 32'hca00004;
      106360: inst = 32'h38632800;
      106361: inst = 32'h38842800;
      106362: inst = 32'h10a00001;
      106363: inst = 32'hca09f7f;
      106364: inst = 32'h13e00001;
      106365: inst = 32'hfe0d96a;
      106366: inst = 32'h5be00000;
      106367: inst = 32'h8c50000;
      106368: inst = 32'h24612800;
      106369: inst = 32'h10a00000;
      106370: inst = 32'hca00014;
      106371: inst = 32'h24822800;
      106372: inst = 32'h10a00000;
      106373: inst = 32'hca00004;
      106374: inst = 32'h38632800;
      106375: inst = 32'h38842800;
      106376: inst = 32'h10a00001;
      106377: inst = 32'hca09f8d;
      106378: inst = 32'h13e00001;
      106379: inst = 32'hfe0d96a;
      106380: inst = 32'h5be00000;
      106381: inst = 32'h8c50000;
      106382: inst = 32'h24612800;
      106383: inst = 32'h10a00000;
      106384: inst = 32'hca00014;
      106385: inst = 32'h24822800;
      106386: inst = 32'h10a00000;
      106387: inst = 32'hca00004;
      106388: inst = 32'h38632800;
      106389: inst = 32'h38842800;
      106390: inst = 32'h10a00001;
      106391: inst = 32'hca09f9b;
      106392: inst = 32'h13e00001;
      106393: inst = 32'hfe0d96a;
      106394: inst = 32'h5be00000;
      106395: inst = 32'h8c50000;
      106396: inst = 32'h24612800;
      106397: inst = 32'h10a00000;
      106398: inst = 32'hca00014;
      106399: inst = 32'h24822800;
      106400: inst = 32'h10a00000;
      106401: inst = 32'hca00004;
      106402: inst = 32'h38632800;
      106403: inst = 32'h38842800;
      106404: inst = 32'h10a00001;
      106405: inst = 32'hca09fa9;
      106406: inst = 32'h13e00001;
      106407: inst = 32'hfe0d96a;
      106408: inst = 32'h5be00000;
      106409: inst = 32'h8c50000;
      106410: inst = 32'h24612800;
      106411: inst = 32'h10a00000;
      106412: inst = 32'hca00015;
      106413: inst = 32'h24822800;
      106414: inst = 32'h10a00000;
      106415: inst = 32'hca00004;
      106416: inst = 32'h38632800;
      106417: inst = 32'h38842800;
      106418: inst = 32'h10a00001;
      106419: inst = 32'hca09fb7;
      106420: inst = 32'h13e00001;
      106421: inst = 32'hfe0d96a;
      106422: inst = 32'h5be00000;
      106423: inst = 32'h8c50000;
      106424: inst = 32'h24612800;
      106425: inst = 32'h10a00000;
      106426: inst = 32'hca00015;
      106427: inst = 32'h24822800;
      106428: inst = 32'h10a00000;
      106429: inst = 32'hca00004;
      106430: inst = 32'h38632800;
      106431: inst = 32'h38842800;
      106432: inst = 32'h10a00001;
      106433: inst = 32'hca09fc5;
      106434: inst = 32'h13e00001;
      106435: inst = 32'hfe0d96a;
      106436: inst = 32'h5be00000;
      106437: inst = 32'h8c50000;
      106438: inst = 32'h24612800;
      106439: inst = 32'h10a00000;
      106440: inst = 32'hca00015;
      106441: inst = 32'h24822800;
      106442: inst = 32'h10a00000;
      106443: inst = 32'hca00004;
      106444: inst = 32'h38632800;
      106445: inst = 32'h38842800;
      106446: inst = 32'h10a00001;
      106447: inst = 32'hca09fd3;
      106448: inst = 32'h13e00001;
      106449: inst = 32'hfe0d96a;
      106450: inst = 32'h5be00000;
      106451: inst = 32'h8c50000;
      106452: inst = 32'h24612800;
      106453: inst = 32'h10a00000;
      106454: inst = 32'hca00015;
      106455: inst = 32'h24822800;
      106456: inst = 32'h10a00000;
      106457: inst = 32'hca00004;
      106458: inst = 32'h38632800;
      106459: inst = 32'h38842800;
      106460: inst = 32'h10a00001;
      106461: inst = 32'hca09fe1;
      106462: inst = 32'h13e00001;
      106463: inst = 32'hfe0d96a;
      106464: inst = 32'h5be00000;
      106465: inst = 32'h8c50000;
      106466: inst = 32'h24612800;
      106467: inst = 32'h10a00000;
      106468: inst = 32'hca00015;
      106469: inst = 32'h24822800;
      106470: inst = 32'h10a00000;
      106471: inst = 32'hca00004;
      106472: inst = 32'h38632800;
      106473: inst = 32'h38842800;
      106474: inst = 32'h10a00001;
      106475: inst = 32'hca09fef;
      106476: inst = 32'h13e00001;
      106477: inst = 32'hfe0d96a;
      106478: inst = 32'h5be00000;
      106479: inst = 32'h8c50000;
      106480: inst = 32'h24612800;
      106481: inst = 32'h10a00000;
      106482: inst = 32'hca00015;
      106483: inst = 32'h24822800;
      106484: inst = 32'h10a00000;
      106485: inst = 32'hca00004;
      106486: inst = 32'h38632800;
      106487: inst = 32'h38842800;
      106488: inst = 32'h10a00001;
      106489: inst = 32'hca09ffd;
      106490: inst = 32'h13e00001;
      106491: inst = 32'hfe0d96a;
      106492: inst = 32'h5be00000;
      106493: inst = 32'h8c50000;
      106494: inst = 32'h24612800;
      106495: inst = 32'h10a00000;
      106496: inst = 32'hca00015;
      106497: inst = 32'h24822800;
      106498: inst = 32'h10a00000;
      106499: inst = 32'hca00004;
      106500: inst = 32'h38632800;
      106501: inst = 32'h38842800;
      106502: inst = 32'h10a00001;
      106503: inst = 32'hca0a00b;
      106504: inst = 32'h13e00001;
      106505: inst = 32'hfe0d96a;
      106506: inst = 32'h5be00000;
      106507: inst = 32'h8c50000;
      106508: inst = 32'h24612800;
      106509: inst = 32'h10a00000;
      106510: inst = 32'hca00015;
      106511: inst = 32'h24822800;
      106512: inst = 32'h10a00000;
      106513: inst = 32'hca00004;
      106514: inst = 32'h38632800;
      106515: inst = 32'h38842800;
      106516: inst = 32'h10a00001;
      106517: inst = 32'hca0a019;
      106518: inst = 32'h13e00001;
      106519: inst = 32'hfe0d96a;
      106520: inst = 32'h5be00000;
      106521: inst = 32'h8c50000;
      106522: inst = 32'h24612800;
      106523: inst = 32'h10a00000;
      106524: inst = 32'hca00015;
      106525: inst = 32'h24822800;
      106526: inst = 32'h10a00000;
      106527: inst = 32'hca00004;
      106528: inst = 32'h38632800;
      106529: inst = 32'h38842800;
      106530: inst = 32'h10a00001;
      106531: inst = 32'hca0a027;
      106532: inst = 32'h13e00001;
      106533: inst = 32'hfe0d96a;
      106534: inst = 32'h5be00000;
      106535: inst = 32'h8c50000;
      106536: inst = 32'h24612800;
      106537: inst = 32'h10a00000;
      106538: inst = 32'hca00015;
      106539: inst = 32'h24822800;
      106540: inst = 32'h10a00000;
      106541: inst = 32'hca00004;
      106542: inst = 32'h38632800;
      106543: inst = 32'h38842800;
      106544: inst = 32'h10a00001;
      106545: inst = 32'hca0a035;
      106546: inst = 32'h13e00001;
      106547: inst = 32'hfe0d96a;
      106548: inst = 32'h5be00000;
      106549: inst = 32'h8c50000;
      106550: inst = 32'h24612800;
      106551: inst = 32'h10a00000;
      106552: inst = 32'hca00015;
      106553: inst = 32'h24822800;
      106554: inst = 32'h10a00000;
      106555: inst = 32'hca00004;
      106556: inst = 32'h38632800;
      106557: inst = 32'h38842800;
      106558: inst = 32'h10a00001;
      106559: inst = 32'hca0a043;
      106560: inst = 32'h13e00001;
      106561: inst = 32'hfe0d96a;
      106562: inst = 32'h5be00000;
      106563: inst = 32'h8c50000;
      106564: inst = 32'h24612800;
      106565: inst = 32'h10a00000;
      106566: inst = 32'hca00015;
      106567: inst = 32'h24822800;
      106568: inst = 32'h10a00000;
      106569: inst = 32'hca00004;
      106570: inst = 32'h38632800;
      106571: inst = 32'h38842800;
      106572: inst = 32'h10a00001;
      106573: inst = 32'hca0a051;
      106574: inst = 32'h13e00001;
      106575: inst = 32'hfe0d96a;
      106576: inst = 32'h5be00000;
      106577: inst = 32'h8c50000;
      106578: inst = 32'h24612800;
      106579: inst = 32'h10a00000;
      106580: inst = 32'hca00015;
      106581: inst = 32'h24822800;
      106582: inst = 32'h10a00000;
      106583: inst = 32'hca00004;
      106584: inst = 32'h38632800;
      106585: inst = 32'h38842800;
      106586: inst = 32'h10a00001;
      106587: inst = 32'hca0a05f;
      106588: inst = 32'h13e00001;
      106589: inst = 32'hfe0d96a;
      106590: inst = 32'h5be00000;
      106591: inst = 32'h8c50000;
      106592: inst = 32'h24612800;
      106593: inst = 32'h10a00000;
      106594: inst = 32'hca00015;
      106595: inst = 32'h24822800;
      106596: inst = 32'h10a00000;
      106597: inst = 32'hca00004;
      106598: inst = 32'h38632800;
      106599: inst = 32'h38842800;
      106600: inst = 32'h10a00001;
      106601: inst = 32'hca0a06d;
      106602: inst = 32'h13e00001;
      106603: inst = 32'hfe0d96a;
      106604: inst = 32'h5be00000;
      106605: inst = 32'h8c50000;
      106606: inst = 32'h24612800;
      106607: inst = 32'h10a00000;
      106608: inst = 32'hca00015;
      106609: inst = 32'h24822800;
      106610: inst = 32'h10a00000;
      106611: inst = 32'hca00004;
      106612: inst = 32'h38632800;
      106613: inst = 32'h38842800;
      106614: inst = 32'h10a00001;
      106615: inst = 32'hca0a07b;
      106616: inst = 32'h13e00001;
      106617: inst = 32'hfe0d96a;
      106618: inst = 32'h5be00000;
      106619: inst = 32'h8c50000;
      106620: inst = 32'h24612800;
      106621: inst = 32'h10a00000;
      106622: inst = 32'hca00015;
      106623: inst = 32'h24822800;
      106624: inst = 32'h10a00000;
      106625: inst = 32'hca00004;
      106626: inst = 32'h38632800;
      106627: inst = 32'h38842800;
      106628: inst = 32'h10a00001;
      106629: inst = 32'hca0a089;
      106630: inst = 32'h13e00001;
      106631: inst = 32'hfe0d96a;
      106632: inst = 32'h5be00000;
      106633: inst = 32'h8c50000;
      106634: inst = 32'h24612800;
      106635: inst = 32'h10a00000;
      106636: inst = 32'hca00015;
      106637: inst = 32'h24822800;
      106638: inst = 32'h10a00000;
      106639: inst = 32'hca00004;
      106640: inst = 32'h38632800;
      106641: inst = 32'h38842800;
      106642: inst = 32'h10a00001;
      106643: inst = 32'hca0a097;
      106644: inst = 32'h13e00001;
      106645: inst = 32'hfe0d96a;
      106646: inst = 32'h5be00000;
      106647: inst = 32'h8c50000;
      106648: inst = 32'h24612800;
      106649: inst = 32'h10a00000;
      106650: inst = 32'hca00015;
      106651: inst = 32'h24822800;
      106652: inst = 32'h10a00000;
      106653: inst = 32'hca00004;
      106654: inst = 32'h38632800;
      106655: inst = 32'h38842800;
      106656: inst = 32'h10a00001;
      106657: inst = 32'hca0a0a5;
      106658: inst = 32'h13e00001;
      106659: inst = 32'hfe0d96a;
      106660: inst = 32'h5be00000;
      106661: inst = 32'h8c50000;
      106662: inst = 32'h24612800;
      106663: inst = 32'h10a00000;
      106664: inst = 32'hca00015;
      106665: inst = 32'h24822800;
      106666: inst = 32'h10a00000;
      106667: inst = 32'hca00004;
      106668: inst = 32'h38632800;
      106669: inst = 32'h38842800;
      106670: inst = 32'h10a00001;
      106671: inst = 32'hca0a0b3;
      106672: inst = 32'h13e00001;
      106673: inst = 32'hfe0d96a;
      106674: inst = 32'h5be00000;
      106675: inst = 32'h8c50000;
      106676: inst = 32'h24612800;
      106677: inst = 32'h10a00000;
      106678: inst = 32'hca00015;
      106679: inst = 32'h24822800;
      106680: inst = 32'h10a00000;
      106681: inst = 32'hca00004;
      106682: inst = 32'h38632800;
      106683: inst = 32'h38842800;
      106684: inst = 32'h10a00001;
      106685: inst = 32'hca0a0c1;
      106686: inst = 32'h13e00001;
      106687: inst = 32'hfe0d96a;
      106688: inst = 32'h5be00000;
      106689: inst = 32'h8c50000;
      106690: inst = 32'h24612800;
      106691: inst = 32'h10a00000;
      106692: inst = 32'hca00015;
      106693: inst = 32'h24822800;
      106694: inst = 32'h10a00000;
      106695: inst = 32'hca00004;
      106696: inst = 32'h38632800;
      106697: inst = 32'h38842800;
      106698: inst = 32'h10a00001;
      106699: inst = 32'hca0a0cf;
      106700: inst = 32'h13e00001;
      106701: inst = 32'hfe0d96a;
      106702: inst = 32'h5be00000;
      106703: inst = 32'h8c50000;
      106704: inst = 32'h24612800;
      106705: inst = 32'h10a00000;
      106706: inst = 32'hca00015;
      106707: inst = 32'h24822800;
      106708: inst = 32'h10a00000;
      106709: inst = 32'hca00004;
      106710: inst = 32'h38632800;
      106711: inst = 32'h38842800;
      106712: inst = 32'h10a00001;
      106713: inst = 32'hca0a0dd;
      106714: inst = 32'h13e00001;
      106715: inst = 32'hfe0d96a;
      106716: inst = 32'h5be00000;
      106717: inst = 32'h8c50000;
      106718: inst = 32'h24612800;
      106719: inst = 32'h10a00000;
      106720: inst = 32'hca00015;
      106721: inst = 32'h24822800;
      106722: inst = 32'h10a00000;
      106723: inst = 32'hca00004;
      106724: inst = 32'h38632800;
      106725: inst = 32'h38842800;
      106726: inst = 32'h10a00001;
      106727: inst = 32'hca0a0eb;
      106728: inst = 32'h13e00001;
      106729: inst = 32'hfe0d96a;
      106730: inst = 32'h5be00000;
      106731: inst = 32'h8c50000;
      106732: inst = 32'h24612800;
      106733: inst = 32'h10a00000;
      106734: inst = 32'hca00015;
      106735: inst = 32'h24822800;
      106736: inst = 32'h10a00000;
      106737: inst = 32'hca00004;
      106738: inst = 32'h38632800;
      106739: inst = 32'h38842800;
      106740: inst = 32'h10a00001;
      106741: inst = 32'hca0a0f9;
      106742: inst = 32'h13e00001;
      106743: inst = 32'hfe0d96a;
      106744: inst = 32'h5be00000;
      106745: inst = 32'h8c50000;
      106746: inst = 32'h24612800;
      106747: inst = 32'h10a00000;
      106748: inst = 32'hca00015;
      106749: inst = 32'h24822800;
      106750: inst = 32'h10a00000;
      106751: inst = 32'hca00004;
      106752: inst = 32'h38632800;
      106753: inst = 32'h38842800;
      106754: inst = 32'h10a00001;
      106755: inst = 32'hca0a107;
      106756: inst = 32'h13e00001;
      106757: inst = 32'hfe0d96a;
      106758: inst = 32'h5be00000;
      106759: inst = 32'h8c50000;
      106760: inst = 32'h24612800;
      106761: inst = 32'h10a00000;
      106762: inst = 32'hca00015;
      106763: inst = 32'h24822800;
      106764: inst = 32'h10a00000;
      106765: inst = 32'hca00004;
      106766: inst = 32'h38632800;
      106767: inst = 32'h38842800;
      106768: inst = 32'h10a00001;
      106769: inst = 32'hca0a115;
      106770: inst = 32'h13e00001;
      106771: inst = 32'hfe0d96a;
      106772: inst = 32'h5be00000;
      106773: inst = 32'h8c50000;
      106774: inst = 32'h24612800;
      106775: inst = 32'h10a00000;
      106776: inst = 32'hca00015;
      106777: inst = 32'h24822800;
      106778: inst = 32'h10a00000;
      106779: inst = 32'hca00004;
      106780: inst = 32'h38632800;
      106781: inst = 32'h38842800;
      106782: inst = 32'h10a00001;
      106783: inst = 32'hca0a123;
      106784: inst = 32'h13e00001;
      106785: inst = 32'hfe0d96a;
      106786: inst = 32'h5be00000;
      106787: inst = 32'h8c50000;
      106788: inst = 32'h24612800;
      106789: inst = 32'h10a00000;
      106790: inst = 32'hca00015;
      106791: inst = 32'h24822800;
      106792: inst = 32'h10a00000;
      106793: inst = 32'hca00004;
      106794: inst = 32'h38632800;
      106795: inst = 32'h38842800;
      106796: inst = 32'h10a00001;
      106797: inst = 32'hca0a131;
      106798: inst = 32'h13e00001;
      106799: inst = 32'hfe0d96a;
      106800: inst = 32'h5be00000;
      106801: inst = 32'h8c50000;
      106802: inst = 32'h24612800;
      106803: inst = 32'h10a00000;
      106804: inst = 32'hca00015;
      106805: inst = 32'h24822800;
      106806: inst = 32'h10a00000;
      106807: inst = 32'hca00004;
      106808: inst = 32'h38632800;
      106809: inst = 32'h38842800;
      106810: inst = 32'h10a00001;
      106811: inst = 32'hca0a13f;
      106812: inst = 32'h13e00001;
      106813: inst = 32'hfe0d96a;
      106814: inst = 32'h5be00000;
      106815: inst = 32'h8c50000;
      106816: inst = 32'h24612800;
      106817: inst = 32'h10a00000;
      106818: inst = 32'hca00015;
      106819: inst = 32'h24822800;
      106820: inst = 32'h10a00000;
      106821: inst = 32'hca00004;
      106822: inst = 32'h38632800;
      106823: inst = 32'h38842800;
      106824: inst = 32'h10a00001;
      106825: inst = 32'hca0a14d;
      106826: inst = 32'h13e00001;
      106827: inst = 32'hfe0d96a;
      106828: inst = 32'h5be00000;
      106829: inst = 32'h8c50000;
      106830: inst = 32'h24612800;
      106831: inst = 32'h10a00000;
      106832: inst = 32'hca00015;
      106833: inst = 32'h24822800;
      106834: inst = 32'h10a00000;
      106835: inst = 32'hca00004;
      106836: inst = 32'h38632800;
      106837: inst = 32'h38842800;
      106838: inst = 32'h10a00001;
      106839: inst = 32'hca0a15b;
      106840: inst = 32'h13e00001;
      106841: inst = 32'hfe0d96a;
      106842: inst = 32'h5be00000;
      106843: inst = 32'h8c50000;
      106844: inst = 32'h24612800;
      106845: inst = 32'h10a00000;
      106846: inst = 32'hca00015;
      106847: inst = 32'h24822800;
      106848: inst = 32'h10a00000;
      106849: inst = 32'hca00004;
      106850: inst = 32'h38632800;
      106851: inst = 32'h38842800;
      106852: inst = 32'h10a00001;
      106853: inst = 32'hca0a169;
      106854: inst = 32'h13e00001;
      106855: inst = 32'hfe0d96a;
      106856: inst = 32'h5be00000;
      106857: inst = 32'h8c50000;
      106858: inst = 32'h24612800;
      106859: inst = 32'h10a00000;
      106860: inst = 32'hca00015;
      106861: inst = 32'h24822800;
      106862: inst = 32'h10a00000;
      106863: inst = 32'hca00004;
      106864: inst = 32'h38632800;
      106865: inst = 32'h38842800;
      106866: inst = 32'h10a00001;
      106867: inst = 32'hca0a177;
      106868: inst = 32'h13e00001;
      106869: inst = 32'hfe0d96a;
      106870: inst = 32'h5be00000;
      106871: inst = 32'h8c50000;
      106872: inst = 32'h24612800;
      106873: inst = 32'h10a00000;
      106874: inst = 32'hca00015;
      106875: inst = 32'h24822800;
      106876: inst = 32'h10a00000;
      106877: inst = 32'hca00004;
      106878: inst = 32'h38632800;
      106879: inst = 32'h38842800;
      106880: inst = 32'h10a00001;
      106881: inst = 32'hca0a185;
      106882: inst = 32'h13e00001;
      106883: inst = 32'hfe0d96a;
      106884: inst = 32'h5be00000;
      106885: inst = 32'h8c50000;
      106886: inst = 32'h24612800;
      106887: inst = 32'h10a00000;
      106888: inst = 32'hca00015;
      106889: inst = 32'h24822800;
      106890: inst = 32'h10a00000;
      106891: inst = 32'hca00004;
      106892: inst = 32'h38632800;
      106893: inst = 32'h38842800;
      106894: inst = 32'h10a00001;
      106895: inst = 32'hca0a193;
      106896: inst = 32'h13e00001;
      106897: inst = 32'hfe0d96a;
      106898: inst = 32'h5be00000;
      106899: inst = 32'h8c50000;
      106900: inst = 32'h24612800;
      106901: inst = 32'h10a00000;
      106902: inst = 32'hca00015;
      106903: inst = 32'h24822800;
      106904: inst = 32'h10a00000;
      106905: inst = 32'hca00004;
      106906: inst = 32'h38632800;
      106907: inst = 32'h38842800;
      106908: inst = 32'h10a00001;
      106909: inst = 32'hca0a1a1;
      106910: inst = 32'h13e00001;
      106911: inst = 32'hfe0d96a;
      106912: inst = 32'h5be00000;
      106913: inst = 32'h8c50000;
      106914: inst = 32'h24612800;
      106915: inst = 32'h10a00000;
      106916: inst = 32'hca00015;
      106917: inst = 32'h24822800;
      106918: inst = 32'h10a00000;
      106919: inst = 32'hca00004;
      106920: inst = 32'h38632800;
      106921: inst = 32'h38842800;
      106922: inst = 32'h10a00001;
      106923: inst = 32'hca0a1af;
      106924: inst = 32'h13e00001;
      106925: inst = 32'hfe0d96a;
      106926: inst = 32'h5be00000;
      106927: inst = 32'h8c50000;
      106928: inst = 32'h24612800;
      106929: inst = 32'h10a00000;
      106930: inst = 32'hca00015;
      106931: inst = 32'h24822800;
      106932: inst = 32'h10a00000;
      106933: inst = 32'hca00004;
      106934: inst = 32'h38632800;
      106935: inst = 32'h38842800;
      106936: inst = 32'h10a00001;
      106937: inst = 32'hca0a1bd;
      106938: inst = 32'h13e00001;
      106939: inst = 32'hfe0d96a;
      106940: inst = 32'h5be00000;
      106941: inst = 32'h8c50000;
      106942: inst = 32'h24612800;
      106943: inst = 32'h10a00000;
      106944: inst = 32'hca00015;
      106945: inst = 32'h24822800;
      106946: inst = 32'h10a00000;
      106947: inst = 32'hca00004;
      106948: inst = 32'h38632800;
      106949: inst = 32'h38842800;
      106950: inst = 32'h10a00001;
      106951: inst = 32'hca0a1cb;
      106952: inst = 32'h13e00001;
      106953: inst = 32'hfe0d96a;
      106954: inst = 32'h5be00000;
      106955: inst = 32'h8c50000;
      106956: inst = 32'h24612800;
      106957: inst = 32'h10a00000;
      106958: inst = 32'hca00015;
      106959: inst = 32'h24822800;
      106960: inst = 32'h10a00000;
      106961: inst = 32'hca00004;
      106962: inst = 32'h38632800;
      106963: inst = 32'h38842800;
      106964: inst = 32'h10a00001;
      106965: inst = 32'hca0a1d9;
      106966: inst = 32'h13e00001;
      106967: inst = 32'hfe0d96a;
      106968: inst = 32'h5be00000;
      106969: inst = 32'h8c50000;
      106970: inst = 32'h24612800;
      106971: inst = 32'h10a00000;
      106972: inst = 32'hca00015;
      106973: inst = 32'h24822800;
      106974: inst = 32'h10a00000;
      106975: inst = 32'hca00004;
      106976: inst = 32'h38632800;
      106977: inst = 32'h38842800;
      106978: inst = 32'h10a00001;
      106979: inst = 32'hca0a1e7;
      106980: inst = 32'h13e00001;
      106981: inst = 32'hfe0d96a;
      106982: inst = 32'h5be00000;
      106983: inst = 32'h8c50000;
      106984: inst = 32'h24612800;
      106985: inst = 32'h10a00000;
      106986: inst = 32'hca00015;
      106987: inst = 32'h24822800;
      106988: inst = 32'h10a00000;
      106989: inst = 32'hca00004;
      106990: inst = 32'h38632800;
      106991: inst = 32'h38842800;
      106992: inst = 32'h10a00001;
      106993: inst = 32'hca0a1f5;
      106994: inst = 32'h13e00001;
      106995: inst = 32'hfe0d96a;
      106996: inst = 32'h5be00000;
      106997: inst = 32'h8c50000;
      106998: inst = 32'h24612800;
      106999: inst = 32'h10a00000;
      107000: inst = 32'hca00015;
      107001: inst = 32'h24822800;
      107002: inst = 32'h10a00000;
      107003: inst = 32'hca00004;
      107004: inst = 32'h38632800;
      107005: inst = 32'h38842800;
      107006: inst = 32'h10a00001;
      107007: inst = 32'hca0a203;
      107008: inst = 32'h13e00001;
      107009: inst = 32'hfe0d96a;
      107010: inst = 32'h5be00000;
      107011: inst = 32'h8c50000;
      107012: inst = 32'h24612800;
      107013: inst = 32'h10a00000;
      107014: inst = 32'hca00015;
      107015: inst = 32'h24822800;
      107016: inst = 32'h10a00000;
      107017: inst = 32'hca00004;
      107018: inst = 32'h38632800;
      107019: inst = 32'h38842800;
      107020: inst = 32'h10a00001;
      107021: inst = 32'hca0a211;
      107022: inst = 32'h13e00001;
      107023: inst = 32'hfe0d96a;
      107024: inst = 32'h5be00000;
      107025: inst = 32'h8c50000;
      107026: inst = 32'h24612800;
      107027: inst = 32'h10a00000;
      107028: inst = 32'hca00015;
      107029: inst = 32'h24822800;
      107030: inst = 32'h10a00000;
      107031: inst = 32'hca00004;
      107032: inst = 32'h38632800;
      107033: inst = 32'h38842800;
      107034: inst = 32'h10a00001;
      107035: inst = 32'hca0a21f;
      107036: inst = 32'h13e00001;
      107037: inst = 32'hfe0d96a;
      107038: inst = 32'h5be00000;
      107039: inst = 32'h8c50000;
      107040: inst = 32'h24612800;
      107041: inst = 32'h10a00000;
      107042: inst = 32'hca00015;
      107043: inst = 32'h24822800;
      107044: inst = 32'h10a00000;
      107045: inst = 32'hca00004;
      107046: inst = 32'h38632800;
      107047: inst = 32'h38842800;
      107048: inst = 32'h10a00001;
      107049: inst = 32'hca0a22d;
      107050: inst = 32'h13e00001;
      107051: inst = 32'hfe0d96a;
      107052: inst = 32'h5be00000;
      107053: inst = 32'h8c50000;
      107054: inst = 32'h24612800;
      107055: inst = 32'h10a00000;
      107056: inst = 32'hca00015;
      107057: inst = 32'h24822800;
      107058: inst = 32'h10a00000;
      107059: inst = 32'hca00004;
      107060: inst = 32'h38632800;
      107061: inst = 32'h38842800;
      107062: inst = 32'h10a00001;
      107063: inst = 32'hca0a23b;
      107064: inst = 32'h13e00001;
      107065: inst = 32'hfe0d96a;
      107066: inst = 32'h5be00000;
      107067: inst = 32'h8c50000;
      107068: inst = 32'h24612800;
      107069: inst = 32'h10a00000;
      107070: inst = 32'hca00015;
      107071: inst = 32'h24822800;
      107072: inst = 32'h10a00000;
      107073: inst = 32'hca00004;
      107074: inst = 32'h38632800;
      107075: inst = 32'h38842800;
      107076: inst = 32'h10a00001;
      107077: inst = 32'hca0a249;
      107078: inst = 32'h13e00001;
      107079: inst = 32'hfe0d96a;
      107080: inst = 32'h5be00000;
      107081: inst = 32'h8c50000;
      107082: inst = 32'h24612800;
      107083: inst = 32'h10a00000;
      107084: inst = 32'hca00015;
      107085: inst = 32'h24822800;
      107086: inst = 32'h10a00000;
      107087: inst = 32'hca00004;
      107088: inst = 32'h38632800;
      107089: inst = 32'h38842800;
      107090: inst = 32'h10a00001;
      107091: inst = 32'hca0a257;
      107092: inst = 32'h13e00001;
      107093: inst = 32'hfe0d96a;
      107094: inst = 32'h5be00000;
      107095: inst = 32'h8c50000;
      107096: inst = 32'h24612800;
      107097: inst = 32'h10a00000;
      107098: inst = 32'hca00015;
      107099: inst = 32'h24822800;
      107100: inst = 32'h10a00000;
      107101: inst = 32'hca00004;
      107102: inst = 32'h38632800;
      107103: inst = 32'h38842800;
      107104: inst = 32'h10a00001;
      107105: inst = 32'hca0a265;
      107106: inst = 32'h13e00001;
      107107: inst = 32'hfe0d96a;
      107108: inst = 32'h5be00000;
      107109: inst = 32'h8c50000;
      107110: inst = 32'h24612800;
      107111: inst = 32'h10a00000;
      107112: inst = 32'hca00015;
      107113: inst = 32'h24822800;
      107114: inst = 32'h10a00000;
      107115: inst = 32'hca00004;
      107116: inst = 32'h38632800;
      107117: inst = 32'h38842800;
      107118: inst = 32'h10a00001;
      107119: inst = 32'hca0a273;
      107120: inst = 32'h13e00001;
      107121: inst = 32'hfe0d96a;
      107122: inst = 32'h5be00000;
      107123: inst = 32'h8c50000;
      107124: inst = 32'h24612800;
      107125: inst = 32'h10a00000;
      107126: inst = 32'hca00015;
      107127: inst = 32'h24822800;
      107128: inst = 32'h10a00000;
      107129: inst = 32'hca00004;
      107130: inst = 32'h38632800;
      107131: inst = 32'h38842800;
      107132: inst = 32'h10a00001;
      107133: inst = 32'hca0a281;
      107134: inst = 32'h13e00001;
      107135: inst = 32'hfe0d96a;
      107136: inst = 32'h5be00000;
      107137: inst = 32'h8c50000;
      107138: inst = 32'h24612800;
      107139: inst = 32'h10a00000;
      107140: inst = 32'hca00015;
      107141: inst = 32'h24822800;
      107142: inst = 32'h10a00000;
      107143: inst = 32'hca00004;
      107144: inst = 32'h38632800;
      107145: inst = 32'h38842800;
      107146: inst = 32'h10a00001;
      107147: inst = 32'hca0a28f;
      107148: inst = 32'h13e00001;
      107149: inst = 32'hfe0d96a;
      107150: inst = 32'h5be00000;
      107151: inst = 32'h8c50000;
      107152: inst = 32'h24612800;
      107153: inst = 32'h10a00000;
      107154: inst = 32'hca00015;
      107155: inst = 32'h24822800;
      107156: inst = 32'h10a00000;
      107157: inst = 32'hca00004;
      107158: inst = 32'h38632800;
      107159: inst = 32'h38842800;
      107160: inst = 32'h10a00001;
      107161: inst = 32'hca0a29d;
      107162: inst = 32'h13e00001;
      107163: inst = 32'hfe0d96a;
      107164: inst = 32'h5be00000;
      107165: inst = 32'h8c50000;
      107166: inst = 32'h24612800;
      107167: inst = 32'h10a00000;
      107168: inst = 32'hca00015;
      107169: inst = 32'h24822800;
      107170: inst = 32'h10a00000;
      107171: inst = 32'hca00004;
      107172: inst = 32'h38632800;
      107173: inst = 32'h38842800;
      107174: inst = 32'h10a00001;
      107175: inst = 32'hca0a2ab;
      107176: inst = 32'h13e00001;
      107177: inst = 32'hfe0d96a;
      107178: inst = 32'h5be00000;
      107179: inst = 32'h8c50000;
      107180: inst = 32'h24612800;
      107181: inst = 32'h10a00000;
      107182: inst = 32'hca00015;
      107183: inst = 32'h24822800;
      107184: inst = 32'h10a00000;
      107185: inst = 32'hca00004;
      107186: inst = 32'h38632800;
      107187: inst = 32'h38842800;
      107188: inst = 32'h10a00001;
      107189: inst = 32'hca0a2b9;
      107190: inst = 32'h13e00001;
      107191: inst = 32'hfe0d96a;
      107192: inst = 32'h5be00000;
      107193: inst = 32'h8c50000;
      107194: inst = 32'h24612800;
      107195: inst = 32'h10a00000;
      107196: inst = 32'hca00015;
      107197: inst = 32'h24822800;
      107198: inst = 32'h10a00000;
      107199: inst = 32'hca00004;
      107200: inst = 32'h38632800;
      107201: inst = 32'h38842800;
      107202: inst = 32'h10a00001;
      107203: inst = 32'hca0a2c7;
      107204: inst = 32'h13e00001;
      107205: inst = 32'hfe0d96a;
      107206: inst = 32'h5be00000;
      107207: inst = 32'h8c50000;
      107208: inst = 32'h24612800;
      107209: inst = 32'h10a00000;
      107210: inst = 32'hca00015;
      107211: inst = 32'h24822800;
      107212: inst = 32'h10a00000;
      107213: inst = 32'hca00004;
      107214: inst = 32'h38632800;
      107215: inst = 32'h38842800;
      107216: inst = 32'h10a00001;
      107217: inst = 32'hca0a2d5;
      107218: inst = 32'h13e00001;
      107219: inst = 32'hfe0d96a;
      107220: inst = 32'h5be00000;
      107221: inst = 32'h8c50000;
      107222: inst = 32'h24612800;
      107223: inst = 32'h10a00000;
      107224: inst = 32'hca00015;
      107225: inst = 32'h24822800;
      107226: inst = 32'h10a00000;
      107227: inst = 32'hca00004;
      107228: inst = 32'h38632800;
      107229: inst = 32'h38842800;
      107230: inst = 32'h10a00001;
      107231: inst = 32'hca0a2e3;
      107232: inst = 32'h13e00001;
      107233: inst = 32'hfe0d96a;
      107234: inst = 32'h5be00000;
      107235: inst = 32'h8c50000;
      107236: inst = 32'h24612800;
      107237: inst = 32'h10a00000;
      107238: inst = 32'hca00015;
      107239: inst = 32'h24822800;
      107240: inst = 32'h10a00000;
      107241: inst = 32'hca00004;
      107242: inst = 32'h38632800;
      107243: inst = 32'h38842800;
      107244: inst = 32'h10a00001;
      107245: inst = 32'hca0a2f1;
      107246: inst = 32'h13e00001;
      107247: inst = 32'hfe0d96a;
      107248: inst = 32'h5be00000;
      107249: inst = 32'h8c50000;
      107250: inst = 32'h24612800;
      107251: inst = 32'h10a00000;
      107252: inst = 32'hca00015;
      107253: inst = 32'h24822800;
      107254: inst = 32'h10a00000;
      107255: inst = 32'hca00004;
      107256: inst = 32'h38632800;
      107257: inst = 32'h38842800;
      107258: inst = 32'h10a00001;
      107259: inst = 32'hca0a2ff;
      107260: inst = 32'h13e00001;
      107261: inst = 32'hfe0d96a;
      107262: inst = 32'h5be00000;
      107263: inst = 32'h8c50000;
      107264: inst = 32'h24612800;
      107265: inst = 32'h10a00000;
      107266: inst = 32'hca00015;
      107267: inst = 32'h24822800;
      107268: inst = 32'h10a00000;
      107269: inst = 32'hca00004;
      107270: inst = 32'h38632800;
      107271: inst = 32'h38842800;
      107272: inst = 32'h10a00001;
      107273: inst = 32'hca0a30d;
      107274: inst = 32'h13e00001;
      107275: inst = 32'hfe0d96a;
      107276: inst = 32'h5be00000;
      107277: inst = 32'h8c50000;
      107278: inst = 32'h24612800;
      107279: inst = 32'h10a00000;
      107280: inst = 32'hca00015;
      107281: inst = 32'h24822800;
      107282: inst = 32'h10a00000;
      107283: inst = 32'hca00004;
      107284: inst = 32'h38632800;
      107285: inst = 32'h38842800;
      107286: inst = 32'h10a00001;
      107287: inst = 32'hca0a31b;
      107288: inst = 32'h13e00001;
      107289: inst = 32'hfe0d96a;
      107290: inst = 32'h5be00000;
      107291: inst = 32'h8c50000;
      107292: inst = 32'h24612800;
      107293: inst = 32'h10a00000;
      107294: inst = 32'hca00015;
      107295: inst = 32'h24822800;
      107296: inst = 32'h10a00000;
      107297: inst = 32'hca00004;
      107298: inst = 32'h38632800;
      107299: inst = 32'h38842800;
      107300: inst = 32'h10a00001;
      107301: inst = 32'hca0a329;
      107302: inst = 32'h13e00001;
      107303: inst = 32'hfe0d96a;
      107304: inst = 32'h5be00000;
      107305: inst = 32'h8c50000;
      107306: inst = 32'h24612800;
      107307: inst = 32'h10a00000;
      107308: inst = 32'hca00015;
      107309: inst = 32'h24822800;
      107310: inst = 32'h10a00000;
      107311: inst = 32'hca00004;
      107312: inst = 32'h38632800;
      107313: inst = 32'h38842800;
      107314: inst = 32'h10a00001;
      107315: inst = 32'hca0a337;
      107316: inst = 32'h13e00001;
      107317: inst = 32'hfe0d96a;
      107318: inst = 32'h5be00000;
      107319: inst = 32'h8c50000;
      107320: inst = 32'h24612800;
      107321: inst = 32'h10a00000;
      107322: inst = 32'hca00015;
      107323: inst = 32'h24822800;
      107324: inst = 32'h10a00000;
      107325: inst = 32'hca00004;
      107326: inst = 32'h38632800;
      107327: inst = 32'h38842800;
      107328: inst = 32'h10a00001;
      107329: inst = 32'hca0a345;
      107330: inst = 32'h13e00001;
      107331: inst = 32'hfe0d96a;
      107332: inst = 32'h5be00000;
      107333: inst = 32'h8c50000;
      107334: inst = 32'h24612800;
      107335: inst = 32'h10a00000;
      107336: inst = 32'hca00015;
      107337: inst = 32'h24822800;
      107338: inst = 32'h10a00000;
      107339: inst = 32'hca00004;
      107340: inst = 32'h38632800;
      107341: inst = 32'h38842800;
      107342: inst = 32'h10a00001;
      107343: inst = 32'hca0a353;
      107344: inst = 32'h13e00001;
      107345: inst = 32'hfe0d96a;
      107346: inst = 32'h5be00000;
      107347: inst = 32'h8c50000;
      107348: inst = 32'h24612800;
      107349: inst = 32'h10a00000;
      107350: inst = 32'hca00015;
      107351: inst = 32'h24822800;
      107352: inst = 32'h10a00000;
      107353: inst = 32'hca00004;
      107354: inst = 32'h38632800;
      107355: inst = 32'h38842800;
      107356: inst = 32'h10a00001;
      107357: inst = 32'hca0a361;
      107358: inst = 32'h13e00001;
      107359: inst = 32'hfe0d96a;
      107360: inst = 32'h5be00000;
      107361: inst = 32'h8c50000;
      107362: inst = 32'h24612800;
      107363: inst = 32'h10a00000;
      107364: inst = 32'hca00015;
      107365: inst = 32'h24822800;
      107366: inst = 32'h10a00000;
      107367: inst = 32'hca00004;
      107368: inst = 32'h38632800;
      107369: inst = 32'h38842800;
      107370: inst = 32'h10a00001;
      107371: inst = 32'hca0a36f;
      107372: inst = 32'h13e00001;
      107373: inst = 32'hfe0d96a;
      107374: inst = 32'h5be00000;
      107375: inst = 32'h8c50000;
      107376: inst = 32'h24612800;
      107377: inst = 32'h10a00000;
      107378: inst = 32'hca00015;
      107379: inst = 32'h24822800;
      107380: inst = 32'h10a00000;
      107381: inst = 32'hca00004;
      107382: inst = 32'h38632800;
      107383: inst = 32'h38842800;
      107384: inst = 32'h10a00001;
      107385: inst = 32'hca0a37d;
      107386: inst = 32'h13e00001;
      107387: inst = 32'hfe0d96a;
      107388: inst = 32'h5be00000;
      107389: inst = 32'h8c50000;
      107390: inst = 32'h24612800;
      107391: inst = 32'h10a00000;
      107392: inst = 32'hca00015;
      107393: inst = 32'h24822800;
      107394: inst = 32'h10a00000;
      107395: inst = 32'hca00004;
      107396: inst = 32'h38632800;
      107397: inst = 32'h38842800;
      107398: inst = 32'h10a00001;
      107399: inst = 32'hca0a38b;
      107400: inst = 32'h13e00001;
      107401: inst = 32'hfe0d96a;
      107402: inst = 32'h5be00000;
      107403: inst = 32'h8c50000;
      107404: inst = 32'h24612800;
      107405: inst = 32'h10a00000;
      107406: inst = 32'hca00015;
      107407: inst = 32'h24822800;
      107408: inst = 32'h10a00000;
      107409: inst = 32'hca00004;
      107410: inst = 32'h38632800;
      107411: inst = 32'h38842800;
      107412: inst = 32'h10a00001;
      107413: inst = 32'hca0a399;
      107414: inst = 32'h13e00001;
      107415: inst = 32'hfe0d96a;
      107416: inst = 32'h5be00000;
      107417: inst = 32'h8c50000;
      107418: inst = 32'h24612800;
      107419: inst = 32'h10a00000;
      107420: inst = 32'hca00015;
      107421: inst = 32'h24822800;
      107422: inst = 32'h10a00000;
      107423: inst = 32'hca00004;
      107424: inst = 32'h38632800;
      107425: inst = 32'h38842800;
      107426: inst = 32'h10a00001;
      107427: inst = 32'hca0a3a7;
      107428: inst = 32'h13e00001;
      107429: inst = 32'hfe0d96a;
      107430: inst = 32'h5be00000;
      107431: inst = 32'h8c50000;
      107432: inst = 32'h24612800;
      107433: inst = 32'h10a00000;
      107434: inst = 32'hca00015;
      107435: inst = 32'h24822800;
      107436: inst = 32'h10a00000;
      107437: inst = 32'hca00004;
      107438: inst = 32'h38632800;
      107439: inst = 32'h38842800;
      107440: inst = 32'h10a00001;
      107441: inst = 32'hca0a3b5;
      107442: inst = 32'h13e00001;
      107443: inst = 32'hfe0d96a;
      107444: inst = 32'h5be00000;
      107445: inst = 32'h8c50000;
      107446: inst = 32'h24612800;
      107447: inst = 32'h10a00000;
      107448: inst = 32'hca00015;
      107449: inst = 32'h24822800;
      107450: inst = 32'h10a00000;
      107451: inst = 32'hca00004;
      107452: inst = 32'h38632800;
      107453: inst = 32'h38842800;
      107454: inst = 32'h10a00001;
      107455: inst = 32'hca0a3c3;
      107456: inst = 32'h13e00001;
      107457: inst = 32'hfe0d96a;
      107458: inst = 32'h5be00000;
      107459: inst = 32'h8c50000;
      107460: inst = 32'h24612800;
      107461: inst = 32'h10a00000;
      107462: inst = 32'hca00015;
      107463: inst = 32'h24822800;
      107464: inst = 32'h10a00000;
      107465: inst = 32'hca00004;
      107466: inst = 32'h38632800;
      107467: inst = 32'h38842800;
      107468: inst = 32'h10a00001;
      107469: inst = 32'hca0a3d1;
      107470: inst = 32'h13e00001;
      107471: inst = 32'hfe0d96a;
      107472: inst = 32'h5be00000;
      107473: inst = 32'h8c50000;
      107474: inst = 32'h24612800;
      107475: inst = 32'h10a00000;
      107476: inst = 32'hca00015;
      107477: inst = 32'h24822800;
      107478: inst = 32'h10a00000;
      107479: inst = 32'hca00004;
      107480: inst = 32'h38632800;
      107481: inst = 32'h38842800;
      107482: inst = 32'h10a00001;
      107483: inst = 32'hca0a3df;
      107484: inst = 32'h13e00001;
      107485: inst = 32'hfe0d96a;
      107486: inst = 32'h5be00000;
      107487: inst = 32'h8c50000;
      107488: inst = 32'h24612800;
      107489: inst = 32'h10a00000;
      107490: inst = 32'hca00015;
      107491: inst = 32'h24822800;
      107492: inst = 32'h10a00000;
      107493: inst = 32'hca00004;
      107494: inst = 32'h38632800;
      107495: inst = 32'h38842800;
      107496: inst = 32'h10a00001;
      107497: inst = 32'hca0a3ed;
      107498: inst = 32'h13e00001;
      107499: inst = 32'hfe0d96a;
      107500: inst = 32'h5be00000;
      107501: inst = 32'h8c50000;
      107502: inst = 32'h24612800;
      107503: inst = 32'h10a00000;
      107504: inst = 32'hca00015;
      107505: inst = 32'h24822800;
      107506: inst = 32'h10a00000;
      107507: inst = 32'hca00004;
      107508: inst = 32'h38632800;
      107509: inst = 32'h38842800;
      107510: inst = 32'h10a00001;
      107511: inst = 32'hca0a3fb;
      107512: inst = 32'h13e00001;
      107513: inst = 32'hfe0d96a;
      107514: inst = 32'h5be00000;
      107515: inst = 32'h8c50000;
      107516: inst = 32'h24612800;
      107517: inst = 32'h10a00000;
      107518: inst = 32'hca00015;
      107519: inst = 32'h24822800;
      107520: inst = 32'h10a00000;
      107521: inst = 32'hca00004;
      107522: inst = 32'h38632800;
      107523: inst = 32'h38842800;
      107524: inst = 32'h10a00001;
      107525: inst = 32'hca0a409;
      107526: inst = 32'h13e00001;
      107527: inst = 32'hfe0d96a;
      107528: inst = 32'h5be00000;
      107529: inst = 32'h8c50000;
      107530: inst = 32'h24612800;
      107531: inst = 32'h10a00000;
      107532: inst = 32'hca00015;
      107533: inst = 32'h24822800;
      107534: inst = 32'h10a00000;
      107535: inst = 32'hca00004;
      107536: inst = 32'h38632800;
      107537: inst = 32'h38842800;
      107538: inst = 32'h10a00001;
      107539: inst = 32'hca0a417;
      107540: inst = 32'h13e00001;
      107541: inst = 32'hfe0d96a;
      107542: inst = 32'h5be00000;
      107543: inst = 32'h8c50000;
      107544: inst = 32'h24612800;
      107545: inst = 32'h10a00000;
      107546: inst = 32'hca00015;
      107547: inst = 32'h24822800;
      107548: inst = 32'h10a00000;
      107549: inst = 32'hca00004;
      107550: inst = 32'h38632800;
      107551: inst = 32'h38842800;
      107552: inst = 32'h10a00001;
      107553: inst = 32'hca0a425;
      107554: inst = 32'h13e00001;
      107555: inst = 32'hfe0d96a;
      107556: inst = 32'h5be00000;
      107557: inst = 32'h8c50000;
      107558: inst = 32'h24612800;
      107559: inst = 32'h10a00000;
      107560: inst = 32'hca00015;
      107561: inst = 32'h24822800;
      107562: inst = 32'h10a00000;
      107563: inst = 32'hca00004;
      107564: inst = 32'h38632800;
      107565: inst = 32'h38842800;
      107566: inst = 32'h10a00001;
      107567: inst = 32'hca0a433;
      107568: inst = 32'h13e00001;
      107569: inst = 32'hfe0d96a;
      107570: inst = 32'h5be00000;
      107571: inst = 32'h8c50000;
      107572: inst = 32'h24612800;
      107573: inst = 32'h10a00000;
      107574: inst = 32'hca00015;
      107575: inst = 32'h24822800;
      107576: inst = 32'h10a00000;
      107577: inst = 32'hca00004;
      107578: inst = 32'h38632800;
      107579: inst = 32'h38842800;
      107580: inst = 32'h10a00001;
      107581: inst = 32'hca0a441;
      107582: inst = 32'h13e00001;
      107583: inst = 32'hfe0d96a;
      107584: inst = 32'h5be00000;
      107585: inst = 32'h8c50000;
      107586: inst = 32'h24612800;
      107587: inst = 32'h10a00000;
      107588: inst = 32'hca00015;
      107589: inst = 32'h24822800;
      107590: inst = 32'h10a00000;
      107591: inst = 32'hca00004;
      107592: inst = 32'h38632800;
      107593: inst = 32'h38842800;
      107594: inst = 32'h10a00001;
      107595: inst = 32'hca0a44f;
      107596: inst = 32'h13e00001;
      107597: inst = 32'hfe0d96a;
      107598: inst = 32'h5be00000;
      107599: inst = 32'h8c50000;
      107600: inst = 32'h24612800;
      107601: inst = 32'h10a00000;
      107602: inst = 32'hca00015;
      107603: inst = 32'h24822800;
      107604: inst = 32'h10a00000;
      107605: inst = 32'hca00004;
      107606: inst = 32'h38632800;
      107607: inst = 32'h38842800;
      107608: inst = 32'h10a00001;
      107609: inst = 32'hca0a45d;
      107610: inst = 32'h13e00001;
      107611: inst = 32'hfe0d96a;
      107612: inst = 32'h5be00000;
      107613: inst = 32'h8c50000;
      107614: inst = 32'h24612800;
      107615: inst = 32'h10a00000;
      107616: inst = 32'hca00015;
      107617: inst = 32'h24822800;
      107618: inst = 32'h10a00000;
      107619: inst = 32'hca00004;
      107620: inst = 32'h38632800;
      107621: inst = 32'h38842800;
      107622: inst = 32'h10a00001;
      107623: inst = 32'hca0a46b;
      107624: inst = 32'h13e00001;
      107625: inst = 32'hfe0d96a;
      107626: inst = 32'h5be00000;
      107627: inst = 32'h8c50000;
      107628: inst = 32'h24612800;
      107629: inst = 32'h10a00000;
      107630: inst = 32'hca00015;
      107631: inst = 32'h24822800;
      107632: inst = 32'h10a00000;
      107633: inst = 32'hca00004;
      107634: inst = 32'h38632800;
      107635: inst = 32'h38842800;
      107636: inst = 32'h10a00001;
      107637: inst = 32'hca0a479;
      107638: inst = 32'h13e00001;
      107639: inst = 32'hfe0d96a;
      107640: inst = 32'h5be00000;
      107641: inst = 32'h8c50000;
      107642: inst = 32'h24612800;
      107643: inst = 32'h10a00000;
      107644: inst = 32'hca00015;
      107645: inst = 32'h24822800;
      107646: inst = 32'h10a00000;
      107647: inst = 32'hca00004;
      107648: inst = 32'h38632800;
      107649: inst = 32'h38842800;
      107650: inst = 32'h10a00001;
      107651: inst = 32'hca0a487;
      107652: inst = 32'h13e00001;
      107653: inst = 32'hfe0d96a;
      107654: inst = 32'h5be00000;
      107655: inst = 32'h8c50000;
      107656: inst = 32'h24612800;
      107657: inst = 32'h10a00000;
      107658: inst = 32'hca00015;
      107659: inst = 32'h24822800;
      107660: inst = 32'h10a00000;
      107661: inst = 32'hca00004;
      107662: inst = 32'h38632800;
      107663: inst = 32'h38842800;
      107664: inst = 32'h10a00001;
      107665: inst = 32'hca0a495;
      107666: inst = 32'h13e00001;
      107667: inst = 32'hfe0d96a;
      107668: inst = 32'h5be00000;
      107669: inst = 32'h8c50000;
      107670: inst = 32'h24612800;
      107671: inst = 32'h10a00000;
      107672: inst = 32'hca00015;
      107673: inst = 32'h24822800;
      107674: inst = 32'h10a00000;
      107675: inst = 32'hca00004;
      107676: inst = 32'h38632800;
      107677: inst = 32'h38842800;
      107678: inst = 32'h10a00001;
      107679: inst = 32'hca0a4a3;
      107680: inst = 32'h13e00001;
      107681: inst = 32'hfe0d96a;
      107682: inst = 32'h5be00000;
      107683: inst = 32'h8c50000;
      107684: inst = 32'h24612800;
      107685: inst = 32'h10a00000;
      107686: inst = 32'hca00015;
      107687: inst = 32'h24822800;
      107688: inst = 32'h10a00000;
      107689: inst = 32'hca00004;
      107690: inst = 32'h38632800;
      107691: inst = 32'h38842800;
      107692: inst = 32'h10a00001;
      107693: inst = 32'hca0a4b1;
      107694: inst = 32'h13e00001;
      107695: inst = 32'hfe0d96a;
      107696: inst = 32'h5be00000;
      107697: inst = 32'h8c50000;
      107698: inst = 32'h24612800;
      107699: inst = 32'h10a00000;
      107700: inst = 32'hca00015;
      107701: inst = 32'h24822800;
      107702: inst = 32'h10a00000;
      107703: inst = 32'hca00004;
      107704: inst = 32'h38632800;
      107705: inst = 32'h38842800;
      107706: inst = 32'h10a00001;
      107707: inst = 32'hca0a4bf;
      107708: inst = 32'h13e00001;
      107709: inst = 32'hfe0d96a;
      107710: inst = 32'h5be00000;
      107711: inst = 32'h8c50000;
      107712: inst = 32'h24612800;
      107713: inst = 32'h10a00000;
      107714: inst = 32'hca00015;
      107715: inst = 32'h24822800;
      107716: inst = 32'h10a00000;
      107717: inst = 32'hca00004;
      107718: inst = 32'h38632800;
      107719: inst = 32'h38842800;
      107720: inst = 32'h10a00001;
      107721: inst = 32'hca0a4cd;
      107722: inst = 32'h13e00001;
      107723: inst = 32'hfe0d96a;
      107724: inst = 32'h5be00000;
      107725: inst = 32'h8c50000;
      107726: inst = 32'h24612800;
      107727: inst = 32'h10a00000;
      107728: inst = 32'hca00015;
      107729: inst = 32'h24822800;
      107730: inst = 32'h10a00000;
      107731: inst = 32'hca00004;
      107732: inst = 32'h38632800;
      107733: inst = 32'h38842800;
      107734: inst = 32'h10a00001;
      107735: inst = 32'hca0a4db;
      107736: inst = 32'h13e00001;
      107737: inst = 32'hfe0d96a;
      107738: inst = 32'h5be00000;
      107739: inst = 32'h8c50000;
      107740: inst = 32'h24612800;
      107741: inst = 32'h10a00000;
      107742: inst = 32'hca00015;
      107743: inst = 32'h24822800;
      107744: inst = 32'h10a00000;
      107745: inst = 32'hca00004;
      107746: inst = 32'h38632800;
      107747: inst = 32'h38842800;
      107748: inst = 32'h10a00001;
      107749: inst = 32'hca0a4e9;
      107750: inst = 32'h13e00001;
      107751: inst = 32'hfe0d96a;
      107752: inst = 32'h5be00000;
      107753: inst = 32'h8c50000;
      107754: inst = 32'h24612800;
      107755: inst = 32'h10a00000;
      107756: inst = 32'hca00016;
      107757: inst = 32'h24822800;
      107758: inst = 32'h10a00000;
      107759: inst = 32'hca00004;
      107760: inst = 32'h38632800;
      107761: inst = 32'h38842800;
      107762: inst = 32'h10a00001;
      107763: inst = 32'hca0a4f7;
      107764: inst = 32'h13e00001;
      107765: inst = 32'hfe0d96a;
      107766: inst = 32'h5be00000;
      107767: inst = 32'h8c50000;
      107768: inst = 32'h24612800;
      107769: inst = 32'h10a00000;
      107770: inst = 32'hca00016;
      107771: inst = 32'h24822800;
      107772: inst = 32'h10a00000;
      107773: inst = 32'hca00004;
      107774: inst = 32'h38632800;
      107775: inst = 32'h38842800;
      107776: inst = 32'h10a00001;
      107777: inst = 32'hca0a505;
      107778: inst = 32'h13e00001;
      107779: inst = 32'hfe0d96a;
      107780: inst = 32'h5be00000;
      107781: inst = 32'h8c50000;
      107782: inst = 32'h24612800;
      107783: inst = 32'h10a00000;
      107784: inst = 32'hca00016;
      107785: inst = 32'h24822800;
      107786: inst = 32'h10a00000;
      107787: inst = 32'hca00004;
      107788: inst = 32'h38632800;
      107789: inst = 32'h38842800;
      107790: inst = 32'h10a00001;
      107791: inst = 32'hca0a513;
      107792: inst = 32'h13e00001;
      107793: inst = 32'hfe0d96a;
      107794: inst = 32'h5be00000;
      107795: inst = 32'h8c50000;
      107796: inst = 32'h24612800;
      107797: inst = 32'h10a00000;
      107798: inst = 32'hca00016;
      107799: inst = 32'h24822800;
      107800: inst = 32'h10a00000;
      107801: inst = 32'hca00004;
      107802: inst = 32'h38632800;
      107803: inst = 32'h38842800;
      107804: inst = 32'h10a00001;
      107805: inst = 32'hca0a521;
      107806: inst = 32'h13e00001;
      107807: inst = 32'hfe0d96a;
      107808: inst = 32'h5be00000;
      107809: inst = 32'h8c50000;
      107810: inst = 32'h24612800;
      107811: inst = 32'h10a00000;
      107812: inst = 32'hca00016;
      107813: inst = 32'h24822800;
      107814: inst = 32'h10a00000;
      107815: inst = 32'hca00004;
      107816: inst = 32'h38632800;
      107817: inst = 32'h38842800;
      107818: inst = 32'h10a00001;
      107819: inst = 32'hca0a52f;
      107820: inst = 32'h13e00001;
      107821: inst = 32'hfe0d96a;
      107822: inst = 32'h5be00000;
      107823: inst = 32'h8c50000;
      107824: inst = 32'h24612800;
      107825: inst = 32'h10a00000;
      107826: inst = 32'hca00016;
      107827: inst = 32'h24822800;
      107828: inst = 32'h10a00000;
      107829: inst = 32'hca00004;
      107830: inst = 32'h38632800;
      107831: inst = 32'h38842800;
      107832: inst = 32'h10a00001;
      107833: inst = 32'hca0a53d;
      107834: inst = 32'h13e00001;
      107835: inst = 32'hfe0d96a;
      107836: inst = 32'h5be00000;
      107837: inst = 32'h8c50000;
      107838: inst = 32'h24612800;
      107839: inst = 32'h10a00000;
      107840: inst = 32'hca00016;
      107841: inst = 32'h24822800;
      107842: inst = 32'h10a00000;
      107843: inst = 32'hca00004;
      107844: inst = 32'h38632800;
      107845: inst = 32'h38842800;
      107846: inst = 32'h10a00001;
      107847: inst = 32'hca0a54b;
      107848: inst = 32'h13e00001;
      107849: inst = 32'hfe0d96a;
      107850: inst = 32'h5be00000;
      107851: inst = 32'h8c50000;
      107852: inst = 32'h24612800;
      107853: inst = 32'h10a00000;
      107854: inst = 32'hca00016;
      107855: inst = 32'h24822800;
      107856: inst = 32'h10a00000;
      107857: inst = 32'hca00004;
      107858: inst = 32'h38632800;
      107859: inst = 32'h38842800;
      107860: inst = 32'h10a00001;
      107861: inst = 32'hca0a559;
      107862: inst = 32'h13e00001;
      107863: inst = 32'hfe0d96a;
      107864: inst = 32'h5be00000;
      107865: inst = 32'h8c50000;
      107866: inst = 32'h24612800;
      107867: inst = 32'h10a00000;
      107868: inst = 32'hca00016;
      107869: inst = 32'h24822800;
      107870: inst = 32'h10a00000;
      107871: inst = 32'hca00004;
      107872: inst = 32'h38632800;
      107873: inst = 32'h38842800;
      107874: inst = 32'h10a00001;
      107875: inst = 32'hca0a567;
      107876: inst = 32'h13e00001;
      107877: inst = 32'hfe0d96a;
      107878: inst = 32'h5be00000;
      107879: inst = 32'h8c50000;
      107880: inst = 32'h24612800;
      107881: inst = 32'h10a00000;
      107882: inst = 32'hca00016;
      107883: inst = 32'h24822800;
      107884: inst = 32'h10a00000;
      107885: inst = 32'hca00004;
      107886: inst = 32'h38632800;
      107887: inst = 32'h38842800;
      107888: inst = 32'h10a00001;
      107889: inst = 32'hca0a575;
      107890: inst = 32'h13e00001;
      107891: inst = 32'hfe0d96a;
      107892: inst = 32'h5be00000;
      107893: inst = 32'h8c50000;
      107894: inst = 32'h24612800;
      107895: inst = 32'h10a00000;
      107896: inst = 32'hca00016;
      107897: inst = 32'h24822800;
      107898: inst = 32'h10a00000;
      107899: inst = 32'hca00004;
      107900: inst = 32'h38632800;
      107901: inst = 32'h38842800;
      107902: inst = 32'h10a00001;
      107903: inst = 32'hca0a583;
      107904: inst = 32'h13e00001;
      107905: inst = 32'hfe0d96a;
      107906: inst = 32'h5be00000;
      107907: inst = 32'h8c50000;
      107908: inst = 32'h24612800;
      107909: inst = 32'h10a00000;
      107910: inst = 32'hca00016;
      107911: inst = 32'h24822800;
      107912: inst = 32'h10a00000;
      107913: inst = 32'hca00004;
      107914: inst = 32'h38632800;
      107915: inst = 32'h38842800;
      107916: inst = 32'h10a00001;
      107917: inst = 32'hca0a591;
      107918: inst = 32'h13e00001;
      107919: inst = 32'hfe0d96a;
      107920: inst = 32'h5be00000;
      107921: inst = 32'h8c50000;
      107922: inst = 32'h24612800;
      107923: inst = 32'h10a00000;
      107924: inst = 32'hca00016;
      107925: inst = 32'h24822800;
      107926: inst = 32'h10a00000;
      107927: inst = 32'hca00004;
      107928: inst = 32'h38632800;
      107929: inst = 32'h38842800;
      107930: inst = 32'h10a00001;
      107931: inst = 32'hca0a59f;
      107932: inst = 32'h13e00001;
      107933: inst = 32'hfe0d96a;
      107934: inst = 32'h5be00000;
      107935: inst = 32'h8c50000;
      107936: inst = 32'h24612800;
      107937: inst = 32'h10a00000;
      107938: inst = 32'hca00016;
      107939: inst = 32'h24822800;
      107940: inst = 32'h10a00000;
      107941: inst = 32'hca00004;
      107942: inst = 32'h38632800;
      107943: inst = 32'h38842800;
      107944: inst = 32'h10a00001;
      107945: inst = 32'hca0a5ad;
      107946: inst = 32'h13e00001;
      107947: inst = 32'hfe0d96a;
      107948: inst = 32'h5be00000;
      107949: inst = 32'h8c50000;
      107950: inst = 32'h24612800;
      107951: inst = 32'h10a00000;
      107952: inst = 32'hca00016;
      107953: inst = 32'h24822800;
      107954: inst = 32'h10a00000;
      107955: inst = 32'hca00004;
      107956: inst = 32'h38632800;
      107957: inst = 32'h38842800;
      107958: inst = 32'h10a00001;
      107959: inst = 32'hca0a5bb;
      107960: inst = 32'h13e00001;
      107961: inst = 32'hfe0d96a;
      107962: inst = 32'h5be00000;
      107963: inst = 32'h8c50000;
      107964: inst = 32'h24612800;
      107965: inst = 32'h10a00000;
      107966: inst = 32'hca00016;
      107967: inst = 32'h24822800;
      107968: inst = 32'h10a00000;
      107969: inst = 32'hca00004;
      107970: inst = 32'h38632800;
      107971: inst = 32'h38842800;
      107972: inst = 32'h10a00001;
      107973: inst = 32'hca0a5c9;
      107974: inst = 32'h13e00001;
      107975: inst = 32'hfe0d96a;
      107976: inst = 32'h5be00000;
      107977: inst = 32'h8c50000;
      107978: inst = 32'h24612800;
      107979: inst = 32'h10a00000;
      107980: inst = 32'hca00016;
      107981: inst = 32'h24822800;
      107982: inst = 32'h10a00000;
      107983: inst = 32'hca00004;
      107984: inst = 32'h38632800;
      107985: inst = 32'h38842800;
      107986: inst = 32'h10a00001;
      107987: inst = 32'hca0a5d7;
      107988: inst = 32'h13e00001;
      107989: inst = 32'hfe0d96a;
      107990: inst = 32'h5be00000;
      107991: inst = 32'h8c50000;
      107992: inst = 32'h24612800;
      107993: inst = 32'h10a00000;
      107994: inst = 32'hca00016;
      107995: inst = 32'h24822800;
      107996: inst = 32'h10a00000;
      107997: inst = 32'hca00004;
      107998: inst = 32'h38632800;
      107999: inst = 32'h38842800;
      108000: inst = 32'h10a00001;
      108001: inst = 32'hca0a5e5;
      108002: inst = 32'h13e00001;
      108003: inst = 32'hfe0d96a;
      108004: inst = 32'h5be00000;
      108005: inst = 32'h8c50000;
      108006: inst = 32'h24612800;
      108007: inst = 32'h10a00000;
      108008: inst = 32'hca00016;
      108009: inst = 32'h24822800;
      108010: inst = 32'h10a00000;
      108011: inst = 32'hca00004;
      108012: inst = 32'h38632800;
      108013: inst = 32'h38842800;
      108014: inst = 32'h10a00001;
      108015: inst = 32'hca0a5f3;
      108016: inst = 32'h13e00001;
      108017: inst = 32'hfe0d96a;
      108018: inst = 32'h5be00000;
      108019: inst = 32'h8c50000;
      108020: inst = 32'h24612800;
      108021: inst = 32'h10a00000;
      108022: inst = 32'hca00016;
      108023: inst = 32'h24822800;
      108024: inst = 32'h10a00000;
      108025: inst = 32'hca00004;
      108026: inst = 32'h38632800;
      108027: inst = 32'h38842800;
      108028: inst = 32'h10a00001;
      108029: inst = 32'hca0a601;
      108030: inst = 32'h13e00001;
      108031: inst = 32'hfe0d96a;
      108032: inst = 32'h5be00000;
      108033: inst = 32'h8c50000;
      108034: inst = 32'h24612800;
      108035: inst = 32'h10a00000;
      108036: inst = 32'hca00016;
      108037: inst = 32'h24822800;
      108038: inst = 32'h10a00000;
      108039: inst = 32'hca00004;
      108040: inst = 32'h38632800;
      108041: inst = 32'h38842800;
      108042: inst = 32'h10a00001;
      108043: inst = 32'hca0a60f;
      108044: inst = 32'h13e00001;
      108045: inst = 32'hfe0d96a;
      108046: inst = 32'h5be00000;
      108047: inst = 32'h8c50000;
      108048: inst = 32'h24612800;
      108049: inst = 32'h10a00000;
      108050: inst = 32'hca00016;
      108051: inst = 32'h24822800;
      108052: inst = 32'h10a00000;
      108053: inst = 32'hca00004;
      108054: inst = 32'h38632800;
      108055: inst = 32'h38842800;
      108056: inst = 32'h10a00001;
      108057: inst = 32'hca0a61d;
      108058: inst = 32'h13e00001;
      108059: inst = 32'hfe0d96a;
      108060: inst = 32'h5be00000;
      108061: inst = 32'h8c50000;
      108062: inst = 32'h24612800;
      108063: inst = 32'h10a00000;
      108064: inst = 32'hca00016;
      108065: inst = 32'h24822800;
      108066: inst = 32'h10a00000;
      108067: inst = 32'hca00004;
      108068: inst = 32'h38632800;
      108069: inst = 32'h38842800;
      108070: inst = 32'h10a00001;
      108071: inst = 32'hca0a62b;
      108072: inst = 32'h13e00001;
      108073: inst = 32'hfe0d96a;
      108074: inst = 32'h5be00000;
      108075: inst = 32'h8c50000;
      108076: inst = 32'h24612800;
      108077: inst = 32'h10a00000;
      108078: inst = 32'hca00016;
      108079: inst = 32'h24822800;
      108080: inst = 32'h10a00000;
      108081: inst = 32'hca00004;
      108082: inst = 32'h38632800;
      108083: inst = 32'h38842800;
      108084: inst = 32'h10a00001;
      108085: inst = 32'hca0a639;
      108086: inst = 32'h13e00001;
      108087: inst = 32'hfe0d96a;
      108088: inst = 32'h5be00000;
      108089: inst = 32'h8c50000;
      108090: inst = 32'h24612800;
      108091: inst = 32'h10a00000;
      108092: inst = 32'hca00016;
      108093: inst = 32'h24822800;
      108094: inst = 32'h10a00000;
      108095: inst = 32'hca00004;
      108096: inst = 32'h38632800;
      108097: inst = 32'h38842800;
      108098: inst = 32'h10a00001;
      108099: inst = 32'hca0a647;
      108100: inst = 32'h13e00001;
      108101: inst = 32'hfe0d96a;
      108102: inst = 32'h5be00000;
      108103: inst = 32'h8c50000;
      108104: inst = 32'h24612800;
      108105: inst = 32'h10a00000;
      108106: inst = 32'hca00016;
      108107: inst = 32'h24822800;
      108108: inst = 32'h10a00000;
      108109: inst = 32'hca00004;
      108110: inst = 32'h38632800;
      108111: inst = 32'h38842800;
      108112: inst = 32'h10a00001;
      108113: inst = 32'hca0a655;
      108114: inst = 32'h13e00001;
      108115: inst = 32'hfe0d96a;
      108116: inst = 32'h5be00000;
      108117: inst = 32'h8c50000;
      108118: inst = 32'h24612800;
      108119: inst = 32'h10a00000;
      108120: inst = 32'hca00016;
      108121: inst = 32'h24822800;
      108122: inst = 32'h10a00000;
      108123: inst = 32'hca00004;
      108124: inst = 32'h38632800;
      108125: inst = 32'h38842800;
      108126: inst = 32'h10a00001;
      108127: inst = 32'hca0a663;
      108128: inst = 32'h13e00001;
      108129: inst = 32'hfe0d96a;
      108130: inst = 32'h5be00000;
      108131: inst = 32'h8c50000;
      108132: inst = 32'h24612800;
      108133: inst = 32'h10a00000;
      108134: inst = 32'hca00016;
      108135: inst = 32'h24822800;
      108136: inst = 32'h10a00000;
      108137: inst = 32'hca00004;
      108138: inst = 32'h38632800;
      108139: inst = 32'h38842800;
      108140: inst = 32'h10a00001;
      108141: inst = 32'hca0a671;
      108142: inst = 32'h13e00001;
      108143: inst = 32'hfe0d96a;
      108144: inst = 32'h5be00000;
      108145: inst = 32'h8c50000;
      108146: inst = 32'h24612800;
      108147: inst = 32'h10a00000;
      108148: inst = 32'hca00016;
      108149: inst = 32'h24822800;
      108150: inst = 32'h10a00000;
      108151: inst = 32'hca00004;
      108152: inst = 32'h38632800;
      108153: inst = 32'h38842800;
      108154: inst = 32'h10a00001;
      108155: inst = 32'hca0a67f;
      108156: inst = 32'h13e00001;
      108157: inst = 32'hfe0d96a;
      108158: inst = 32'h5be00000;
      108159: inst = 32'h8c50000;
      108160: inst = 32'h24612800;
      108161: inst = 32'h10a00000;
      108162: inst = 32'hca00016;
      108163: inst = 32'h24822800;
      108164: inst = 32'h10a00000;
      108165: inst = 32'hca00004;
      108166: inst = 32'h38632800;
      108167: inst = 32'h38842800;
      108168: inst = 32'h10a00001;
      108169: inst = 32'hca0a68d;
      108170: inst = 32'h13e00001;
      108171: inst = 32'hfe0d96a;
      108172: inst = 32'h5be00000;
      108173: inst = 32'h8c50000;
      108174: inst = 32'h24612800;
      108175: inst = 32'h10a00000;
      108176: inst = 32'hca00016;
      108177: inst = 32'h24822800;
      108178: inst = 32'h10a00000;
      108179: inst = 32'hca00004;
      108180: inst = 32'h38632800;
      108181: inst = 32'h38842800;
      108182: inst = 32'h10a00001;
      108183: inst = 32'hca0a69b;
      108184: inst = 32'h13e00001;
      108185: inst = 32'hfe0d96a;
      108186: inst = 32'h5be00000;
      108187: inst = 32'h8c50000;
      108188: inst = 32'h24612800;
      108189: inst = 32'h10a00000;
      108190: inst = 32'hca00016;
      108191: inst = 32'h24822800;
      108192: inst = 32'h10a00000;
      108193: inst = 32'hca00004;
      108194: inst = 32'h38632800;
      108195: inst = 32'h38842800;
      108196: inst = 32'h10a00001;
      108197: inst = 32'hca0a6a9;
      108198: inst = 32'h13e00001;
      108199: inst = 32'hfe0d96a;
      108200: inst = 32'h5be00000;
      108201: inst = 32'h8c50000;
      108202: inst = 32'h24612800;
      108203: inst = 32'h10a00000;
      108204: inst = 32'hca00016;
      108205: inst = 32'h24822800;
      108206: inst = 32'h10a00000;
      108207: inst = 32'hca00004;
      108208: inst = 32'h38632800;
      108209: inst = 32'h38842800;
      108210: inst = 32'h10a00001;
      108211: inst = 32'hca0a6b7;
      108212: inst = 32'h13e00001;
      108213: inst = 32'hfe0d96a;
      108214: inst = 32'h5be00000;
      108215: inst = 32'h8c50000;
      108216: inst = 32'h24612800;
      108217: inst = 32'h10a00000;
      108218: inst = 32'hca00016;
      108219: inst = 32'h24822800;
      108220: inst = 32'h10a00000;
      108221: inst = 32'hca00004;
      108222: inst = 32'h38632800;
      108223: inst = 32'h38842800;
      108224: inst = 32'h10a00001;
      108225: inst = 32'hca0a6c5;
      108226: inst = 32'h13e00001;
      108227: inst = 32'hfe0d96a;
      108228: inst = 32'h5be00000;
      108229: inst = 32'h8c50000;
      108230: inst = 32'h24612800;
      108231: inst = 32'h10a00000;
      108232: inst = 32'hca00016;
      108233: inst = 32'h24822800;
      108234: inst = 32'h10a00000;
      108235: inst = 32'hca00004;
      108236: inst = 32'h38632800;
      108237: inst = 32'h38842800;
      108238: inst = 32'h10a00001;
      108239: inst = 32'hca0a6d3;
      108240: inst = 32'h13e00001;
      108241: inst = 32'hfe0d96a;
      108242: inst = 32'h5be00000;
      108243: inst = 32'h8c50000;
      108244: inst = 32'h24612800;
      108245: inst = 32'h10a00000;
      108246: inst = 32'hca00016;
      108247: inst = 32'h24822800;
      108248: inst = 32'h10a00000;
      108249: inst = 32'hca00004;
      108250: inst = 32'h38632800;
      108251: inst = 32'h38842800;
      108252: inst = 32'h10a00001;
      108253: inst = 32'hca0a6e1;
      108254: inst = 32'h13e00001;
      108255: inst = 32'hfe0d96a;
      108256: inst = 32'h5be00000;
      108257: inst = 32'h8c50000;
      108258: inst = 32'h24612800;
      108259: inst = 32'h10a00000;
      108260: inst = 32'hca00016;
      108261: inst = 32'h24822800;
      108262: inst = 32'h10a00000;
      108263: inst = 32'hca00004;
      108264: inst = 32'h38632800;
      108265: inst = 32'h38842800;
      108266: inst = 32'h10a00001;
      108267: inst = 32'hca0a6ef;
      108268: inst = 32'h13e00001;
      108269: inst = 32'hfe0d96a;
      108270: inst = 32'h5be00000;
      108271: inst = 32'h8c50000;
      108272: inst = 32'h24612800;
      108273: inst = 32'h10a00000;
      108274: inst = 32'hca00016;
      108275: inst = 32'h24822800;
      108276: inst = 32'h10a00000;
      108277: inst = 32'hca00004;
      108278: inst = 32'h38632800;
      108279: inst = 32'h38842800;
      108280: inst = 32'h10a00001;
      108281: inst = 32'hca0a6fd;
      108282: inst = 32'h13e00001;
      108283: inst = 32'hfe0d96a;
      108284: inst = 32'h5be00000;
      108285: inst = 32'h8c50000;
      108286: inst = 32'h24612800;
      108287: inst = 32'h10a00000;
      108288: inst = 32'hca00016;
      108289: inst = 32'h24822800;
      108290: inst = 32'h10a00000;
      108291: inst = 32'hca00004;
      108292: inst = 32'h38632800;
      108293: inst = 32'h38842800;
      108294: inst = 32'h10a00001;
      108295: inst = 32'hca0a70b;
      108296: inst = 32'h13e00001;
      108297: inst = 32'hfe0d96a;
      108298: inst = 32'h5be00000;
      108299: inst = 32'h8c50000;
      108300: inst = 32'h24612800;
      108301: inst = 32'h10a00000;
      108302: inst = 32'hca00016;
      108303: inst = 32'h24822800;
      108304: inst = 32'h10a00000;
      108305: inst = 32'hca00004;
      108306: inst = 32'h38632800;
      108307: inst = 32'h38842800;
      108308: inst = 32'h10a00001;
      108309: inst = 32'hca0a719;
      108310: inst = 32'h13e00001;
      108311: inst = 32'hfe0d96a;
      108312: inst = 32'h5be00000;
      108313: inst = 32'h8c50000;
      108314: inst = 32'h24612800;
      108315: inst = 32'h10a00000;
      108316: inst = 32'hca00016;
      108317: inst = 32'h24822800;
      108318: inst = 32'h10a00000;
      108319: inst = 32'hca00004;
      108320: inst = 32'h38632800;
      108321: inst = 32'h38842800;
      108322: inst = 32'h10a00001;
      108323: inst = 32'hca0a727;
      108324: inst = 32'h13e00001;
      108325: inst = 32'hfe0d96a;
      108326: inst = 32'h5be00000;
      108327: inst = 32'h8c50000;
      108328: inst = 32'h24612800;
      108329: inst = 32'h10a00000;
      108330: inst = 32'hca00016;
      108331: inst = 32'h24822800;
      108332: inst = 32'h10a00000;
      108333: inst = 32'hca00004;
      108334: inst = 32'h38632800;
      108335: inst = 32'h38842800;
      108336: inst = 32'h10a00001;
      108337: inst = 32'hca0a735;
      108338: inst = 32'h13e00001;
      108339: inst = 32'hfe0d96a;
      108340: inst = 32'h5be00000;
      108341: inst = 32'h8c50000;
      108342: inst = 32'h24612800;
      108343: inst = 32'h10a00000;
      108344: inst = 32'hca00016;
      108345: inst = 32'h24822800;
      108346: inst = 32'h10a00000;
      108347: inst = 32'hca00004;
      108348: inst = 32'h38632800;
      108349: inst = 32'h38842800;
      108350: inst = 32'h10a00001;
      108351: inst = 32'hca0a743;
      108352: inst = 32'h13e00001;
      108353: inst = 32'hfe0d96a;
      108354: inst = 32'h5be00000;
      108355: inst = 32'h8c50000;
      108356: inst = 32'h24612800;
      108357: inst = 32'h10a00000;
      108358: inst = 32'hca00016;
      108359: inst = 32'h24822800;
      108360: inst = 32'h10a00000;
      108361: inst = 32'hca00004;
      108362: inst = 32'h38632800;
      108363: inst = 32'h38842800;
      108364: inst = 32'h10a00001;
      108365: inst = 32'hca0a751;
      108366: inst = 32'h13e00001;
      108367: inst = 32'hfe0d96a;
      108368: inst = 32'h5be00000;
      108369: inst = 32'h8c50000;
      108370: inst = 32'h24612800;
      108371: inst = 32'h10a00000;
      108372: inst = 32'hca00016;
      108373: inst = 32'h24822800;
      108374: inst = 32'h10a00000;
      108375: inst = 32'hca00004;
      108376: inst = 32'h38632800;
      108377: inst = 32'h38842800;
      108378: inst = 32'h10a00001;
      108379: inst = 32'hca0a75f;
      108380: inst = 32'h13e00001;
      108381: inst = 32'hfe0d96a;
      108382: inst = 32'h5be00000;
      108383: inst = 32'h8c50000;
      108384: inst = 32'h24612800;
      108385: inst = 32'h10a00000;
      108386: inst = 32'hca00016;
      108387: inst = 32'h24822800;
      108388: inst = 32'h10a00000;
      108389: inst = 32'hca00004;
      108390: inst = 32'h38632800;
      108391: inst = 32'h38842800;
      108392: inst = 32'h10a00001;
      108393: inst = 32'hca0a76d;
      108394: inst = 32'h13e00001;
      108395: inst = 32'hfe0d96a;
      108396: inst = 32'h5be00000;
      108397: inst = 32'h8c50000;
      108398: inst = 32'h24612800;
      108399: inst = 32'h10a00000;
      108400: inst = 32'hca00016;
      108401: inst = 32'h24822800;
      108402: inst = 32'h10a00000;
      108403: inst = 32'hca00004;
      108404: inst = 32'h38632800;
      108405: inst = 32'h38842800;
      108406: inst = 32'h10a00001;
      108407: inst = 32'hca0a77b;
      108408: inst = 32'h13e00001;
      108409: inst = 32'hfe0d96a;
      108410: inst = 32'h5be00000;
      108411: inst = 32'h8c50000;
      108412: inst = 32'h24612800;
      108413: inst = 32'h10a00000;
      108414: inst = 32'hca00016;
      108415: inst = 32'h24822800;
      108416: inst = 32'h10a00000;
      108417: inst = 32'hca00004;
      108418: inst = 32'h38632800;
      108419: inst = 32'h38842800;
      108420: inst = 32'h10a00001;
      108421: inst = 32'hca0a789;
      108422: inst = 32'h13e00001;
      108423: inst = 32'hfe0d96a;
      108424: inst = 32'h5be00000;
      108425: inst = 32'h8c50000;
      108426: inst = 32'h24612800;
      108427: inst = 32'h10a00000;
      108428: inst = 32'hca00016;
      108429: inst = 32'h24822800;
      108430: inst = 32'h10a00000;
      108431: inst = 32'hca00004;
      108432: inst = 32'h38632800;
      108433: inst = 32'h38842800;
      108434: inst = 32'h10a00001;
      108435: inst = 32'hca0a797;
      108436: inst = 32'h13e00001;
      108437: inst = 32'hfe0d96a;
      108438: inst = 32'h5be00000;
      108439: inst = 32'h8c50000;
      108440: inst = 32'h24612800;
      108441: inst = 32'h10a00000;
      108442: inst = 32'hca00016;
      108443: inst = 32'h24822800;
      108444: inst = 32'h10a00000;
      108445: inst = 32'hca00004;
      108446: inst = 32'h38632800;
      108447: inst = 32'h38842800;
      108448: inst = 32'h10a00001;
      108449: inst = 32'hca0a7a5;
      108450: inst = 32'h13e00001;
      108451: inst = 32'hfe0d96a;
      108452: inst = 32'h5be00000;
      108453: inst = 32'h8c50000;
      108454: inst = 32'h24612800;
      108455: inst = 32'h10a00000;
      108456: inst = 32'hca00016;
      108457: inst = 32'h24822800;
      108458: inst = 32'h10a00000;
      108459: inst = 32'hca00004;
      108460: inst = 32'h38632800;
      108461: inst = 32'h38842800;
      108462: inst = 32'h10a00001;
      108463: inst = 32'hca0a7b3;
      108464: inst = 32'h13e00001;
      108465: inst = 32'hfe0d96a;
      108466: inst = 32'h5be00000;
      108467: inst = 32'h8c50000;
      108468: inst = 32'h24612800;
      108469: inst = 32'h10a00000;
      108470: inst = 32'hca00016;
      108471: inst = 32'h24822800;
      108472: inst = 32'h10a00000;
      108473: inst = 32'hca00004;
      108474: inst = 32'h38632800;
      108475: inst = 32'h38842800;
      108476: inst = 32'h10a00001;
      108477: inst = 32'hca0a7c1;
      108478: inst = 32'h13e00001;
      108479: inst = 32'hfe0d96a;
      108480: inst = 32'h5be00000;
      108481: inst = 32'h8c50000;
      108482: inst = 32'h24612800;
      108483: inst = 32'h10a00000;
      108484: inst = 32'hca00016;
      108485: inst = 32'h24822800;
      108486: inst = 32'h10a00000;
      108487: inst = 32'hca00004;
      108488: inst = 32'h38632800;
      108489: inst = 32'h38842800;
      108490: inst = 32'h10a00001;
      108491: inst = 32'hca0a7cf;
      108492: inst = 32'h13e00001;
      108493: inst = 32'hfe0d96a;
      108494: inst = 32'h5be00000;
      108495: inst = 32'h8c50000;
      108496: inst = 32'h24612800;
      108497: inst = 32'h10a00000;
      108498: inst = 32'hca00016;
      108499: inst = 32'h24822800;
      108500: inst = 32'h10a00000;
      108501: inst = 32'hca00004;
      108502: inst = 32'h38632800;
      108503: inst = 32'h38842800;
      108504: inst = 32'h10a00001;
      108505: inst = 32'hca0a7dd;
      108506: inst = 32'h13e00001;
      108507: inst = 32'hfe0d96a;
      108508: inst = 32'h5be00000;
      108509: inst = 32'h8c50000;
      108510: inst = 32'h24612800;
      108511: inst = 32'h10a00000;
      108512: inst = 32'hca00016;
      108513: inst = 32'h24822800;
      108514: inst = 32'h10a00000;
      108515: inst = 32'hca00004;
      108516: inst = 32'h38632800;
      108517: inst = 32'h38842800;
      108518: inst = 32'h10a00001;
      108519: inst = 32'hca0a7eb;
      108520: inst = 32'h13e00001;
      108521: inst = 32'hfe0d96a;
      108522: inst = 32'h5be00000;
      108523: inst = 32'h8c50000;
      108524: inst = 32'h24612800;
      108525: inst = 32'h10a00000;
      108526: inst = 32'hca00016;
      108527: inst = 32'h24822800;
      108528: inst = 32'h10a00000;
      108529: inst = 32'hca00004;
      108530: inst = 32'h38632800;
      108531: inst = 32'h38842800;
      108532: inst = 32'h10a00001;
      108533: inst = 32'hca0a7f9;
      108534: inst = 32'h13e00001;
      108535: inst = 32'hfe0d96a;
      108536: inst = 32'h5be00000;
      108537: inst = 32'h8c50000;
      108538: inst = 32'h24612800;
      108539: inst = 32'h10a00000;
      108540: inst = 32'hca00016;
      108541: inst = 32'h24822800;
      108542: inst = 32'h10a00000;
      108543: inst = 32'hca00004;
      108544: inst = 32'h38632800;
      108545: inst = 32'h38842800;
      108546: inst = 32'h10a00001;
      108547: inst = 32'hca0a807;
      108548: inst = 32'h13e00001;
      108549: inst = 32'hfe0d96a;
      108550: inst = 32'h5be00000;
      108551: inst = 32'h8c50000;
      108552: inst = 32'h24612800;
      108553: inst = 32'h10a00000;
      108554: inst = 32'hca00016;
      108555: inst = 32'h24822800;
      108556: inst = 32'h10a00000;
      108557: inst = 32'hca00004;
      108558: inst = 32'h38632800;
      108559: inst = 32'h38842800;
      108560: inst = 32'h10a00001;
      108561: inst = 32'hca0a815;
      108562: inst = 32'h13e00001;
      108563: inst = 32'hfe0d96a;
      108564: inst = 32'h5be00000;
      108565: inst = 32'h8c50000;
      108566: inst = 32'h24612800;
      108567: inst = 32'h10a00000;
      108568: inst = 32'hca00016;
      108569: inst = 32'h24822800;
      108570: inst = 32'h10a00000;
      108571: inst = 32'hca00004;
      108572: inst = 32'h38632800;
      108573: inst = 32'h38842800;
      108574: inst = 32'h10a00001;
      108575: inst = 32'hca0a823;
      108576: inst = 32'h13e00001;
      108577: inst = 32'hfe0d96a;
      108578: inst = 32'h5be00000;
      108579: inst = 32'h8c50000;
      108580: inst = 32'h24612800;
      108581: inst = 32'h10a00000;
      108582: inst = 32'hca00016;
      108583: inst = 32'h24822800;
      108584: inst = 32'h10a00000;
      108585: inst = 32'hca00004;
      108586: inst = 32'h38632800;
      108587: inst = 32'h38842800;
      108588: inst = 32'h10a00001;
      108589: inst = 32'hca0a831;
      108590: inst = 32'h13e00001;
      108591: inst = 32'hfe0d96a;
      108592: inst = 32'h5be00000;
      108593: inst = 32'h8c50000;
      108594: inst = 32'h24612800;
      108595: inst = 32'h10a00000;
      108596: inst = 32'hca00016;
      108597: inst = 32'h24822800;
      108598: inst = 32'h10a00000;
      108599: inst = 32'hca00004;
      108600: inst = 32'h38632800;
      108601: inst = 32'h38842800;
      108602: inst = 32'h10a00001;
      108603: inst = 32'hca0a83f;
      108604: inst = 32'h13e00001;
      108605: inst = 32'hfe0d96a;
      108606: inst = 32'h5be00000;
      108607: inst = 32'h8c50000;
      108608: inst = 32'h24612800;
      108609: inst = 32'h10a00000;
      108610: inst = 32'hca00016;
      108611: inst = 32'h24822800;
      108612: inst = 32'h10a00000;
      108613: inst = 32'hca00004;
      108614: inst = 32'h38632800;
      108615: inst = 32'h38842800;
      108616: inst = 32'h10a00001;
      108617: inst = 32'hca0a84d;
      108618: inst = 32'h13e00001;
      108619: inst = 32'hfe0d96a;
      108620: inst = 32'h5be00000;
      108621: inst = 32'h8c50000;
      108622: inst = 32'h24612800;
      108623: inst = 32'h10a00000;
      108624: inst = 32'hca00016;
      108625: inst = 32'h24822800;
      108626: inst = 32'h10a00000;
      108627: inst = 32'hca00004;
      108628: inst = 32'h38632800;
      108629: inst = 32'h38842800;
      108630: inst = 32'h10a00001;
      108631: inst = 32'hca0a85b;
      108632: inst = 32'h13e00001;
      108633: inst = 32'hfe0d96a;
      108634: inst = 32'h5be00000;
      108635: inst = 32'h8c50000;
      108636: inst = 32'h24612800;
      108637: inst = 32'h10a00000;
      108638: inst = 32'hca00016;
      108639: inst = 32'h24822800;
      108640: inst = 32'h10a00000;
      108641: inst = 32'hca00004;
      108642: inst = 32'h38632800;
      108643: inst = 32'h38842800;
      108644: inst = 32'h10a00001;
      108645: inst = 32'hca0a869;
      108646: inst = 32'h13e00001;
      108647: inst = 32'hfe0d96a;
      108648: inst = 32'h5be00000;
      108649: inst = 32'h8c50000;
      108650: inst = 32'h24612800;
      108651: inst = 32'h10a00000;
      108652: inst = 32'hca00016;
      108653: inst = 32'h24822800;
      108654: inst = 32'h10a00000;
      108655: inst = 32'hca00004;
      108656: inst = 32'h38632800;
      108657: inst = 32'h38842800;
      108658: inst = 32'h10a00001;
      108659: inst = 32'hca0a877;
      108660: inst = 32'h13e00001;
      108661: inst = 32'hfe0d96a;
      108662: inst = 32'h5be00000;
      108663: inst = 32'h8c50000;
      108664: inst = 32'h24612800;
      108665: inst = 32'h10a00000;
      108666: inst = 32'hca00016;
      108667: inst = 32'h24822800;
      108668: inst = 32'h10a00000;
      108669: inst = 32'hca00004;
      108670: inst = 32'h38632800;
      108671: inst = 32'h38842800;
      108672: inst = 32'h10a00001;
      108673: inst = 32'hca0a885;
      108674: inst = 32'h13e00001;
      108675: inst = 32'hfe0d96a;
      108676: inst = 32'h5be00000;
      108677: inst = 32'h8c50000;
      108678: inst = 32'h24612800;
      108679: inst = 32'h10a00000;
      108680: inst = 32'hca00016;
      108681: inst = 32'h24822800;
      108682: inst = 32'h10a00000;
      108683: inst = 32'hca00004;
      108684: inst = 32'h38632800;
      108685: inst = 32'h38842800;
      108686: inst = 32'h10a00001;
      108687: inst = 32'hca0a893;
      108688: inst = 32'h13e00001;
      108689: inst = 32'hfe0d96a;
      108690: inst = 32'h5be00000;
      108691: inst = 32'h8c50000;
      108692: inst = 32'h24612800;
      108693: inst = 32'h10a00000;
      108694: inst = 32'hca00016;
      108695: inst = 32'h24822800;
      108696: inst = 32'h10a00000;
      108697: inst = 32'hca00004;
      108698: inst = 32'h38632800;
      108699: inst = 32'h38842800;
      108700: inst = 32'h10a00001;
      108701: inst = 32'hca0a8a1;
      108702: inst = 32'h13e00001;
      108703: inst = 32'hfe0d96a;
      108704: inst = 32'h5be00000;
      108705: inst = 32'h8c50000;
      108706: inst = 32'h24612800;
      108707: inst = 32'h10a00000;
      108708: inst = 32'hca00016;
      108709: inst = 32'h24822800;
      108710: inst = 32'h10a00000;
      108711: inst = 32'hca00004;
      108712: inst = 32'h38632800;
      108713: inst = 32'h38842800;
      108714: inst = 32'h10a00001;
      108715: inst = 32'hca0a8af;
      108716: inst = 32'h13e00001;
      108717: inst = 32'hfe0d96a;
      108718: inst = 32'h5be00000;
      108719: inst = 32'h8c50000;
      108720: inst = 32'h24612800;
      108721: inst = 32'h10a00000;
      108722: inst = 32'hca00016;
      108723: inst = 32'h24822800;
      108724: inst = 32'h10a00000;
      108725: inst = 32'hca00004;
      108726: inst = 32'h38632800;
      108727: inst = 32'h38842800;
      108728: inst = 32'h10a00001;
      108729: inst = 32'hca0a8bd;
      108730: inst = 32'h13e00001;
      108731: inst = 32'hfe0d96a;
      108732: inst = 32'h5be00000;
      108733: inst = 32'h8c50000;
      108734: inst = 32'h24612800;
      108735: inst = 32'h10a00000;
      108736: inst = 32'hca00016;
      108737: inst = 32'h24822800;
      108738: inst = 32'h10a00000;
      108739: inst = 32'hca00004;
      108740: inst = 32'h38632800;
      108741: inst = 32'h38842800;
      108742: inst = 32'h10a00001;
      108743: inst = 32'hca0a8cb;
      108744: inst = 32'h13e00001;
      108745: inst = 32'hfe0d96a;
      108746: inst = 32'h5be00000;
      108747: inst = 32'h8c50000;
      108748: inst = 32'h24612800;
      108749: inst = 32'h10a00000;
      108750: inst = 32'hca00016;
      108751: inst = 32'h24822800;
      108752: inst = 32'h10a00000;
      108753: inst = 32'hca00004;
      108754: inst = 32'h38632800;
      108755: inst = 32'h38842800;
      108756: inst = 32'h10a00001;
      108757: inst = 32'hca0a8d9;
      108758: inst = 32'h13e00001;
      108759: inst = 32'hfe0d96a;
      108760: inst = 32'h5be00000;
      108761: inst = 32'h8c50000;
      108762: inst = 32'h24612800;
      108763: inst = 32'h10a00000;
      108764: inst = 32'hca00016;
      108765: inst = 32'h24822800;
      108766: inst = 32'h10a00000;
      108767: inst = 32'hca00004;
      108768: inst = 32'h38632800;
      108769: inst = 32'h38842800;
      108770: inst = 32'h10a00001;
      108771: inst = 32'hca0a8e7;
      108772: inst = 32'h13e00001;
      108773: inst = 32'hfe0d96a;
      108774: inst = 32'h5be00000;
      108775: inst = 32'h8c50000;
      108776: inst = 32'h24612800;
      108777: inst = 32'h10a00000;
      108778: inst = 32'hca00016;
      108779: inst = 32'h24822800;
      108780: inst = 32'h10a00000;
      108781: inst = 32'hca00004;
      108782: inst = 32'h38632800;
      108783: inst = 32'h38842800;
      108784: inst = 32'h10a00001;
      108785: inst = 32'hca0a8f5;
      108786: inst = 32'h13e00001;
      108787: inst = 32'hfe0d96a;
      108788: inst = 32'h5be00000;
      108789: inst = 32'h8c50000;
      108790: inst = 32'h24612800;
      108791: inst = 32'h10a00000;
      108792: inst = 32'hca00016;
      108793: inst = 32'h24822800;
      108794: inst = 32'h10a00000;
      108795: inst = 32'hca00004;
      108796: inst = 32'h38632800;
      108797: inst = 32'h38842800;
      108798: inst = 32'h10a00001;
      108799: inst = 32'hca0a903;
      108800: inst = 32'h13e00001;
      108801: inst = 32'hfe0d96a;
      108802: inst = 32'h5be00000;
      108803: inst = 32'h8c50000;
      108804: inst = 32'h24612800;
      108805: inst = 32'h10a00000;
      108806: inst = 32'hca00016;
      108807: inst = 32'h24822800;
      108808: inst = 32'h10a00000;
      108809: inst = 32'hca00004;
      108810: inst = 32'h38632800;
      108811: inst = 32'h38842800;
      108812: inst = 32'h10a00001;
      108813: inst = 32'hca0a911;
      108814: inst = 32'h13e00001;
      108815: inst = 32'hfe0d96a;
      108816: inst = 32'h5be00000;
      108817: inst = 32'h8c50000;
      108818: inst = 32'h24612800;
      108819: inst = 32'h10a00000;
      108820: inst = 32'hca00016;
      108821: inst = 32'h24822800;
      108822: inst = 32'h10a00000;
      108823: inst = 32'hca00004;
      108824: inst = 32'h38632800;
      108825: inst = 32'h38842800;
      108826: inst = 32'h10a00001;
      108827: inst = 32'hca0a91f;
      108828: inst = 32'h13e00001;
      108829: inst = 32'hfe0d96a;
      108830: inst = 32'h5be00000;
      108831: inst = 32'h8c50000;
      108832: inst = 32'h24612800;
      108833: inst = 32'h10a00000;
      108834: inst = 32'hca00016;
      108835: inst = 32'h24822800;
      108836: inst = 32'h10a00000;
      108837: inst = 32'hca00004;
      108838: inst = 32'h38632800;
      108839: inst = 32'h38842800;
      108840: inst = 32'h10a00001;
      108841: inst = 32'hca0a92d;
      108842: inst = 32'h13e00001;
      108843: inst = 32'hfe0d96a;
      108844: inst = 32'h5be00000;
      108845: inst = 32'h8c50000;
      108846: inst = 32'h24612800;
      108847: inst = 32'h10a00000;
      108848: inst = 32'hca00016;
      108849: inst = 32'h24822800;
      108850: inst = 32'h10a00000;
      108851: inst = 32'hca00004;
      108852: inst = 32'h38632800;
      108853: inst = 32'h38842800;
      108854: inst = 32'h10a00001;
      108855: inst = 32'hca0a93b;
      108856: inst = 32'h13e00001;
      108857: inst = 32'hfe0d96a;
      108858: inst = 32'h5be00000;
      108859: inst = 32'h8c50000;
      108860: inst = 32'h24612800;
      108861: inst = 32'h10a00000;
      108862: inst = 32'hca00016;
      108863: inst = 32'h24822800;
      108864: inst = 32'h10a00000;
      108865: inst = 32'hca00004;
      108866: inst = 32'h38632800;
      108867: inst = 32'h38842800;
      108868: inst = 32'h10a00001;
      108869: inst = 32'hca0a949;
      108870: inst = 32'h13e00001;
      108871: inst = 32'hfe0d96a;
      108872: inst = 32'h5be00000;
      108873: inst = 32'h8c50000;
      108874: inst = 32'h24612800;
      108875: inst = 32'h10a00000;
      108876: inst = 32'hca00016;
      108877: inst = 32'h24822800;
      108878: inst = 32'h10a00000;
      108879: inst = 32'hca00004;
      108880: inst = 32'h38632800;
      108881: inst = 32'h38842800;
      108882: inst = 32'h10a00001;
      108883: inst = 32'hca0a957;
      108884: inst = 32'h13e00001;
      108885: inst = 32'hfe0d96a;
      108886: inst = 32'h5be00000;
      108887: inst = 32'h8c50000;
      108888: inst = 32'h24612800;
      108889: inst = 32'h10a00000;
      108890: inst = 32'hca00016;
      108891: inst = 32'h24822800;
      108892: inst = 32'h10a00000;
      108893: inst = 32'hca00004;
      108894: inst = 32'h38632800;
      108895: inst = 32'h38842800;
      108896: inst = 32'h10a00001;
      108897: inst = 32'hca0a965;
      108898: inst = 32'h13e00001;
      108899: inst = 32'hfe0d96a;
      108900: inst = 32'h5be00000;
      108901: inst = 32'h8c50000;
      108902: inst = 32'h24612800;
      108903: inst = 32'h10a00000;
      108904: inst = 32'hca00016;
      108905: inst = 32'h24822800;
      108906: inst = 32'h10a00000;
      108907: inst = 32'hca00004;
      108908: inst = 32'h38632800;
      108909: inst = 32'h38842800;
      108910: inst = 32'h10a00001;
      108911: inst = 32'hca0a973;
      108912: inst = 32'h13e00001;
      108913: inst = 32'hfe0d96a;
      108914: inst = 32'h5be00000;
      108915: inst = 32'h8c50000;
      108916: inst = 32'h24612800;
      108917: inst = 32'h10a00000;
      108918: inst = 32'hca00016;
      108919: inst = 32'h24822800;
      108920: inst = 32'h10a00000;
      108921: inst = 32'hca00004;
      108922: inst = 32'h38632800;
      108923: inst = 32'h38842800;
      108924: inst = 32'h10a00001;
      108925: inst = 32'hca0a981;
      108926: inst = 32'h13e00001;
      108927: inst = 32'hfe0d96a;
      108928: inst = 32'h5be00000;
      108929: inst = 32'h8c50000;
      108930: inst = 32'h24612800;
      108931: inst = 32'h10a00000;
      108932: inst = 32'hca00016;
      108933: inst = 32'h24822800;
      108934: inst = 32'h10a00000;
      108935: inst = 32'hca00004;
      108936: inst = 32'h38632800;
      108937: inst = 32'h38842800;
      108938: inst = 32'h10a00001;
      108939: inst = 32'hca0a98f;
      108940: inst = 32'h13e00001;
      108941: inst = 32'hfe0d96a;
      108942: inst = 32'h5be00000;
      108943: inst = 32'h8c50000;
      108944: inst = 32'h24612800;
      108945: inst = 32'h10a00000;
      108946: inst = 32'hca00016;
      108947: inst = 32'h24822800;
      108948: inst = 32'h10a00000;
      108949: inst = 32'hca00004;
      108950: inst = 32'h38632800;
      108951: inst = 32'h38842800;
      108952: inst = 32'h10a00001;
      108953: inst = 32'hca0a99d;
      108954: inst = 32'h13e00001;
      108955: inst = 32'hfe0d96a;
      108956: inst = 32'h5be00000;
      108957: inst = 32'h8c50000;
      108958: inst = 32'h24612800;
      108959: inst = 32'h10a00000;
      108960: inst = 32'hca00016;
      108961: inst = 32'h24822800;
      108962: inst = 32'h10a00000;
      108963: inst = 32'hca00004;
      108964: inst = 32'h38632800;
      108965: inst = 32'h38842800;
      108966: inst = 32'h10a00001;
      108967: inst = 32'hca0a9ab;
      108968: inst = 32'h13e00001;
      108969: inst = 32'hfe0d96a;
      108970: inst = 32'h5be00000;
      108971: inst = 32'h8c50000;
      108972: inst = 32'h24612800;
      108973: inst = 32'h10a00000;
      108974: inst = 32'hca00016;
      108975: inst = 32'h24822800;
      108976: inst = 32'h10a00000;
      108977: inst = 32'hca00004;
      108978: inst = 32'h38632800;
      108979: inst = 32'h38842800;
      108980: inst = 32'h10a00001;
      108981: inst = 32'hca0a9b9;
      108982: inst = 32'h13e00001;
      108983: inst = 32'hfe0d96a;
      108984: inst = 32'h5be00000;
      108985: inst = 32'h8c50000;
      108986: inst = 32'h24612800;
      108987: inst = 32'h10a00000;
      108988: inst = 32'hca00016;
      108989: inst = 32'h24822800;
      108990: inst = 32'h10a00000;
      108991: inst = 32'hca00004;
      108992: inst = 32'h38632800;
      108993: inst = 32'h38842800;
      108994: inst = 32'h10a00001;
      108995: inst = 32'hca0a9c7;
      108996: inst = 32'h13e00001;
      108997: inst = 32'hfe0d96a;
      108998: inst = 32'h5be00000;
      108999: inst = 32'h8c50000;
      109000: inst = 32'h24612800;
      109001: inst = 32'h10a00000;
      109002: inst = 32'hca00016;
      109003: inst = 32'h24822800;
      109004: inst = 32'h10a00000;
      109005: inst = 32'hca00004;
      109006: inst = 32'h38632800;
      109007: inst = 32'h38842800;
      109008: inst = 32'h10a00001;
      109009: inst = 32'hca0a9d5;
      109010: inst = 32'h13e00001;
      109011: inst = 32'hfe0d96a;
      109012: inst = 32'h5be00000;
      109013: inst = 32'h8c50000;
      109014: inst = 32'h24612800;
      109015: inst = 32'h10a00000;
      109016: inst = 32'hca00016;
      109017: inst = 32'h24822800;
      109018: inst = 32'h10a00000;
      109019: inst = 32'hca00004;
      109020: inst = 32'h38632800;
      109021: inst = 32'h38842800;
      109022: inst = 32'h10a00001;
      109023: inst = 32'hca0a9e3;
      109024: inst = 32'h13e00001;
      109025: inst = 32'hfe0d96a;
      109026: inst = 32'h5be00000;
      109027: inst = 32'h8c50000;
      109028: inst = 32'h24612800;
      109029: inst = 32'h10a00000;
      109030: inst = 32'hca00016;
      109031: inst = 32'h24822800;
      109032: inst = 32'h10a00000;
      109033: inst = 32'hca00004;
      109034: inst = 32'h38632800;
      109035: inst = 32'h38842800;
      109036: inst = 32'h10a00001;
      109037: inst = 32'hca0a9f1;
      109038: inst = 32'h13e00001;
      109039: inst = 32'hfe0d96a;
      109040: inst = 32'h5be00000;
      109041: inst = 32'h8c50000;
      109042: inst = 32'h24612800;
      109043: inst = 32'h10a00000;
      109044: inst = 32'hca00016;
      109045: inst = 32'h24822800;
      109046: inst = 32'h10a00000;
      109047: inst = 32'hca00004;
      109048: inst = 32'h38632800;
      109049: inst = 32'h38842800;
      109050: inst = 32'h10a00001;
      109051: inst = 32'hca0a9ff;
      109052: inst = 32'h13e00001;
      109053: inst = 32'hfe0d96a;
      109054: inst = 32'h5be00000;
      109055: inst = 32'h8c50000;
      109056: inst = 32'h24612800;
      109057: inst = 32'h10a00000;
      109058: inst = 32'hca00016;
      109059: inst = 32'h24822800;
      109060: inst = 32'h10a00000;
      109061: inst = 32'hca00004;
      109062: inst = 32'h38632800;
      109063: inst = 32'h38842800;
      109064: inst = 32'h10a00001;
      109065: inst = 32'hca0aa0d;
      109066: inst = 32'h13e00001;
      109067: inst = 32'hfe0d96a;
      109068: inst = 32'h5be00000;
      109069: inst = 32'h8c50000;
      109070: inst = 32'h24612800;
      109071: inst = 32'h10a00000;
      109072: inst = 32'hca00016;
      109073: inst = 32'h24822800;
      109074: inst = 32'h10a00000;
      109075: inst = 32'hca00004;
      109076: inst = 32'h38632800;
      109077: inst = 32'h38842800;
      109078: inst = 32'h10a00001;
      109079: inst = 32'hca0aa1b;
      109080: inst = 32'h13e00001;
      109081: inst = 32'hfe0d96a;
      109082: inst = 32'h5be00000;
      109083: inst = 32'h8c50000;
      109084: inst = 32'h24612800;
      109085: inst = 32'h10a00000;
      109086: inst = 32'hca00016;
      109087: inst = 32'h24822800;
      109088: inst = 32'h10a00000;
      109089: inst = 32'hca00004;
      109090: inst = 32'h38632800;
      109091: inst = 32'h38842800;
      109092: inst = 32'h10a00001;
      109093: inst = 32'hca0aa29;
      109094: inst = 32'h13e00001;
      109095: inst = 32'hfe0d96a;
      109096: inst = 32'h5be00000;
      109097: inst = 32'h8c50000;
      109098: inst = 32'h24612800;
      109099: inst = 32'h10a00000;
      109100: inst = 32'hca00017;
      109101: inst = 32'h24822800;
      109102: inst = 32'h10a00000;
      109103: inst = 32'hca00004;
      109104: inst = 32'h38632800;
      109105: inst = 32'h38842800;
      109106: inst = 32'h10a00001;
      109107: inst = 32'hca0aa37;
      109108: inst = 32'h13e00001;
      109109: inst = 32'hfe0d96a;
      109110: inst = 32'h5be00000;
      109111: inst = 32'h8c50000;
      109112: inst = 32'h24612800;
      109113: inst = 32'h10a00000;
      109114: inst = 32'hca00017;
      109115: inst = 32'h24822800;
      109116: inst = 32'h10a00000;
      109117: inst = 32'hca00004;
      109118: inst = 32'h38632800;
      109119: inst = 32'h38842800;
      109120: inst = 32'h10a00001;
      109121: inst = 32'hca0aa45;
      109122: inst = 32'h13e00001;
      109123: inst = 32'hfe0d96a;
      109124: inst = 32'h5be00000;
      109125: inst = 32'h8c50000;
      109126: inst = 32'h24612800;
      109127: inst = 32'h10a00000;
      109128: inst = 32'hca00017;
      109129: inst = 32'h24822800;
      109130: inst = 32'h10a00000;
      109131: inst = 32'hca00004;
      109132: inst = 32'h38632800;
      109133: inst = 32'h38842800;
      109134: inst = 32'h10a00001;
      109135: inst = 32'hca0aa53;
      109136: inst = 32'h13e00001;
      109137: inst = 32'hfe0d96a;
      109138: inst = 32'h5be00000;
      109139: inst = 32'h8c50000;
      109140: inst = 32'h24612800;
      109141: inst = 32'h10a00000;
      109142: inst = 32'hca00017;
      109143: inst = 32'h24822800;
      109144: inst = 32'h10a00000;
      109145: inst = 32'hca00004;
      109146: inst = 32'h38632800;
      109147: inst = 32'h38842800;
      109148: inst = 32'h10a00001;
      109149: inst = 32'hca0aa61;
      109150: inst = 32'h13e00001;
      109151: inst = 32'hfe0d96a;
      109152: inst = 32'h5be00000;
      109153: inst = 32'h8c50000;
      109154: inst = 32'h24612800;
      109155: inst = 32'h10a00000;
      109156: inst = 32'hca00017;
      109157: inst = 32'h24822800;
      109158: inst = 32'h10a00000;
      109159: inst = 32'hca00004;
      109160: inst = 32'h38632800;
      109161: inst = 32'h38842800;
      109162: inst = 32'h10a00001;
      109163: inst = 32'hca0aa6f;
      109164: inst = 32'h13e00001;
      109165: inst = 32'hfe0d96a;
      109166: inst = 32'h5be00000;
      109167: inst = 32'h8c50000;
      109168: inst = 32'h24612800;
      109169: inst = 32'h10a00000;
      109170: inst = 32'hca00017;
      109171: inst = 32'h24822800;
      109172: inst = 32'h10a00000;
      109173: inst = 32'hca00004;
      109174: inst = 32'h38632800;
      109175: inst = 32'h38842800;
      109176: inst = 32'h10a00001;
      109177: inst = 32'hca0aa7d;
      109178: inst = 32'h13e00001;
      109179: inst = 32'hfe0d96a;
      109180: inst = 32'h5be00000;
      109181: inst = 32'h8c50000;
      109182: inst = 32'h24612800;
      109183: inst = 32'h10a00000;
      109184: inst = 32'hca00017;
      109185: inst = 32'h24822800;
      109186: inst = 32'h10a00000;
      109187: inst = 32'hca00004;
      109188: inst = 32'h38632800;
      109189: inst = 32'h38842800;
      109190: inst = 32'h10a00001;
      109191: inst = 32'hca0aa8b;
      109192: inst = 32'h13e00001;
      109193: inst = 32'hfe0d96a;
      109194: inst = 32'h5be00000;
      109195: inst = 32'h8c50000;
      109196: inst = 32'h24612800;
      109197: inst = 32'h10a00000;
      109198: inst = 32'hca00017;
      109199: inst = 32'h24822800;
      109200: inst = 32'h10a00000;
      109201: inst = 32'hca00004;
      109202: inst = 32'h38632800;
      109203: inst = 32'h38842800;
      109204: inst = 32'h10a00001;
      109205: inst = 32'hca0aa99;
      109206: inst = 32'h13e00001;
      109207: inst = 32'hfe0d96a;
      109208: inst = 32'h5be00000;
      109209: inst = 32'h8c50000;
      109210: inst = 32'h24612800;
      109211: inst = 32'h10a00000;
      109212: inst = 32'hca00017;
      109213: inst = 32'h24822800;
      109214: inst = 32'h10a00000;
      109215: inst = 32'hca00004;
      109216: inst = 32'h38632800;
      109217: inst = 32'h38842800;
      109218: inst = 32'h10a00001;
      109219: inst = 32'hca0aaa7;
      109220: inst = 32'h13e00001;
      109221: inst = 32'hfe0d96a;
      109222: inst = 32'h5be00000;
      109223: inst = 32'h8c50000;
      109224: inst = 32'h24612800;
      109225: inst = 32'h10a00000;
      109226: inst = 32'hca00017;
      109227: inst = 32'h24822800;
      109228: inst = 32'h10a00000;
      109229: inst = 32'hca00004;
      109230: inst = 32'h38632800;
      109231: inst = 32'h38842800;
      109232: inst = 32'h10a00001;
      109233: inst = 32'hca0aab5;
      109234: inst = 32'h13e00001;
      109235: inst = 32'hfe0d96a;
      109236: inst = 32'h5be00000;
      109237: inst = 32'h8c50000;
      109238: inst = 32'h24612800;
      109239: inst = 32'h10a00000;
      109240: inst = 32'hca00017;
      109241: inst = 32'h24822800;
      109242: inst = 32'h10a00000;
      109243: inst = 32'hca00004;
      109244: inst = 32'h38632800;
      109245: inst = 32'h38842800;
      109246: inst = 32'h10a00001;
      109247: inst = 32'hca0aac3;
      109248: inst = 32'h13e00001;
      109249: inst = 32'hfe0d96a;
      109250: inst = 32'h5be00000;
      109251: inst = 32'h8c50000;
      109252: inst = 32'h24612800;
      109253: inst = 32'h10a00000;
      109254: inst = 32'hca00017;
      109255: inst = 32'h24822800;
      109256: inst = 32'h10a00000;
      109257: inst = 32'hca00004;
      109258: inst = 32'h38632800;
      109259: inst = 32'h38842800;
      109260: inst = 32'h10a00001;
      109261: inst = 32'hca0aad1;
      109262: inst = 32'h13e00001;
      109263: inst = 32'hfe0d96a;
      109264: inst = 32'h5be00000;
      109265: inst = 32'h8c50000;
      109266: inst = 32'h24612800;
      109267: inst = 32'h10a00000;
      109268: inst = 32'hca00017;
      109269: inst = 32'h24822800;
      109270: inst = 32'h10a00000;
      109271: inst = 32'hca00004;
      109272: inst = 32'h38632800;
      109273: inst = 32'h38842800;
      109274: inst = 32'h10a00001;
      109275: inst = 32'hca0aadf;
      109276: inst = 32'h13e00001;
      109277: inst = 32'hfe0d96a;
      109278: inst = 32'h5be00000;
      109279: inst = 32'h8c50000;
      109280: inst = 32'h24612800;
      109281: inst = 32'h10a00000;
      109282: inst = 32'hca00017;
      109283: inst = 32'h24822800;
      109284: inst = 32'h10a00000;
      109285: inst = 32'hca00004;
      109286: inst = 32'h38632800;
      109287: inst = 32'h38842800;
      109288: inst = 32'h10a00001;
      109289: inst = 32'hca0aaed;
      109290: inst = 32'h13e00001;
      109291: inst = 32'hfe0d96a;
      109292: inst = 32'h5be00000;
      109293: inst = 32'h8c50000;
      109294: inst = 32'h24612800;
      109295: inst = 32'h10a00000;
      109296: inst = 32'hca00017;
      109297: inst = 32'h24822800;
      109298: inst = 32'h10a00000;
      109299: inst = 32'hca00004;
      109300: inst = 32'h38632800;
      109301: inst = 32'h38842800;
      109302: inst = 32'h10a00001;
      109303: inst = 32'hca0aafb;
      109304: inst = 32'h13e00001;
      109305: inst = 32'hfe0d96a;
      109306: inst = 32'h5be00000;
      109307: inst = 32'h8c50000;
      109308: inst = 32'h24612800;
      109309: inst = 32'h10a00000;
      109310: inst = 32'hca00017;
      109311: inst = 32'h24822800;
      109312: inst = 32'h10a00000;
      109313: inst = 32'hca00004;
      109314: inst = 32'h38632800;
      109315: inst = 32'h38842800;
      109316: inst = 32'h10a00001;
      109317: inst = 32'hca0ab09;
      109318: inst = 32'h13e00001;
      109319: inst = 32'hfe0d96a;
      109320: inst = 32'h5be00000;
      109321: inst = 32'h8c50000;
      109322: inst = 32'h24612800;
      109323: inst = 32'h10a00000;
      109324: inst = 32'hca00017;
      109325: inst = 32'h24822800;
      109326: inst = 32'h10a00000;
      109327: inst = 32'hca00004;
      109328: inst = 32'h38632800;
      109329: inst = 32'h38842800;
      109330: inst = 32'h10a00001;
      109331: inst = 32'hca0ab17;
      109332: inst = 32'h13e00001;
      109333: inst = 32'hfe0d96a;
      109334: inst = 32'h5be00000;
      109335: inst = 32'h8c50000;
      109336: inst = 32'h24612800;
      109337: inst = 32'h10a00000;
      109338: inst = 32'hca00017;
      109339: inst = 32'h24822800;
      109340: inst = 32'h10a00000;
      109341: inst = 32'hca00004;
      109342: inst = 32'h38632800;
      109343: inst = 32'h38842800;
      109344: inst = 32'h10a00001;
      109345: inst = 32'hca0ab25;
      109346: inst = 32'h13e00001;
      109347: inst = 32'hfe0d96a;
      109348: inst = 32'h5be00000;
      109349: inst = 32'h8c50000;
      109350: inst = 32'h24612800;
      109351: inst = 32'h10a00000;
      109352: inst = 32'hca00017;
      109353: inst = 32'h24822800;
      109354: inst = 32'h10a00000;
      109355: inst = 32'hca00004;
      109356: inst = 32'h38632800;
      109357: inst = 32'h38842800;
      109358: inst = 32'h10a00001;
      109359: inst = 32'hca0ab33;
      109360: inst = 32'h13e00001;
      109361: inst = 32'hfe0d96a;
      109362: inst = 32'h5be00000;
      109363: inst = 32'h8c50000;
      109364: inst = 32'h24612800;
      109365: inst = 32'h10a00000;
      109366: inst = 32'hca00017;
      109367: inst = 32'h24822800;
      109368: inst = 32'h10a00000;
      109369: inst = 32'hca00004;
      109370: inst = 32'h38632800;
      109371: inst = 32'h38842800;
      109372: inst = 32'h10a00001;
      109373: inst = 32'hca0ab41;
      109374: inst = 32'h13e00001;
      109375: inst = 32'hfe0d96a;
      109376: inst = 32'h5be00000;
      109377: inst = 32'h8c50000;
      109378: inst = 32'h24612800;
      109379: inst = 32'h10a00000;
      109380: inst = 32'hca00017;
      109381: inst = 32'h24822800;
      109382: inst = 32'h10a00000;
      109383: inst = 32'hca00004;
      109384: inst = 32'h38632800;
      109385: inst = 32'h38842800;
      109386: inst = 32'h10a00001;
      109387: inst = 32'hca0ab4f;
      109388: inst = 32'h13e00001;
      109389: inst = 32'hfe0d96a;
      109390: inst = 32'h5be00000;
      109391: inst = 32'h8c50000;
      109392: inst = 32'h24612800;
      109393: inst = 32'h10a00000;
      109394: inst = 32'hca00017;
      109395: inst = 32'h24822800;
      109396: inst = 32'h10a00000;
      109397: inst = 32'hca00004;
      109398: inst = 32'h38632800;
      109399: inst = 32'h38842800;
      109400: inst = 32'h10a00001;
      109401: inst = 32'hca0ab5d;
      109402: inst = 32'h13e00001;
      109403: inst = 32'hfe0d96a;
      109404: inst = 32'h5be00000;
      109405: inst = 32'h8c50000;
      109406: inst = 32'h24612800;
      109407: inst = 32'h10a00000;
      109408: inst = 32'hca00017;
      109409: inst = 32'h24822800;
      109410: inst = 32'h10a00000;
      109411: inst = 32'hca00004;
      109412: inst = 32'h38632800;
      109413: inst = 32'h38842800;
      109414: inst = 32'h10a00001;
      109415: inst = 32'hca0ab6b;
      109416: inst = 32'h13e00001;
      109417: inst = 32'hfe0d96a;
      109418: inst = 32'h5be00000;
      109419: inst = 32'h8c50000;
      109420: inst = 32'h24612800;
      109421: inst = 32'h10a00000;
      109422: inst = 32'hca00017;
      109423: inst = 32'h24822800;
      109424: inst = 32'h10a00000;
      109425: inst = 32'hca00004;
      109426: inst = 32'h38632800;
      109427: inst = 32'h38842800;
      109428: inst = 32'h10a00001;
      109429: inst = 32'hca0ab79;
      109430: inst = 32'h13e00001;
      109431: inst = 32'hfe0d96a;
      109432: inst = 32'h5be00000;
      109433: inst = 32'h8c50000;
      109434: inst = 32'h24612800;
      109435: inst = 32'h10a00000;
      109436: inst = 32'hca00017;
      109437: inst = 32'h24822800;
      109438: inst = 32'h10a00000;
      109439: inst = 32'hca00004;
      109440: inst = 32'h38632800;
      109441: inst = 32'h38842800;
      109442: inst = 32'h10a00001;
      109443: inst = 32'hca0ab87;
      109444: inst = 32'h13e00001;
      109445: inst = 32'hfe0d96a;
      109446: inst = 32'h5be00000;
      109447: inst = 32'h8c50000;
      109448: inst = 32'h24612800;
      109449: inst = 32'h10a00000;
      109450: inst = 32'hca00017;
      109451: inst = 32'h24822800;
      109452: inst = 32'h10a00000;
      109453: inst = 32'hca00004;
      109454: inst = 32'h38632800;
      109455: inst = 32'h38842800;
      109456: inst = 32'h10a00001;
      109457: inst = 32'hca0ab95;
      109458: inst = 32'h13e00001;
      109459: inst = 32'hfe0d96a;
      109460: inst = 32'h5be00000;
      109461: inst = 32'h8c50000;
      109462: inst = 32'h24612800;
      109463: inst = 32'h10a00000;
      109464: inst = 32'hca00017;
      109465: inst = 32'h24822800;
      109466: inst = 32'h10a00000;
      109467: inst = 32'hca00004;
      109468: inst = 32'h38632800;
      109469: inst = 32'h38842800;
      109470: inst = 32'h10a00001;
      109471: inst = 32'hca0aba3;
      109472: inst = 32'h13e00001;
      109473: inst = 32'hfe0d96a;
      109474: inst = 32'h5be00000;
      109475: inst = 32'h8c50000;
      109476: inst = 32'h24612800;
      109477: inst = 32'h10a00000;
      109478: inst = 32'hca00017;
      109479: inst = 32'h24822800;
      109480: inst = 32'h10a00000;
      109481: inst = 32'hca00004;
      109482: inst = 32'h38632800;
      109483: inst = 32'h38842800;
      109484: inst = 32'h10a00001;
      109485: inst = 32'hca0abb1;
      109486: inst = 32'h13e00001;
      109487: inst = 32'hfe0d96a;
      109488: inst = 32'h5be00000;
      109489: inst = 32'h8c50000;
      109490: inst = 32'h24612800;
      109491: inst = 32'h10a00000;
      109492: inst = 32'hca00017;
      109493: inst = 32'h24822800;
      109494: inst = 32'h10a00000;
      109495: inst = 32'hca00004;
      109496: inst = 32'h38632800;
      109497: inst = 32'h38842800;
      109498: inst = 32'h10a00001;
      109499: inst = 32'hca0abbf;
      109500: inst = 32'h13e00001;
      109501: inst = 32'hfe0d96a;
      109502: inst = 32'h5be00000;
      109503: inst = 32'h8c50000;
      109504: inst = 32'h24612800;
      109505: inst = 32'h10a00000;
      109506: inst = 32'hca00017;
      109507: inst = 32'h24822800;
      109508: inst = 32'h10a00000;
      109509: inst = 32'hca00004;
      109510: inst = 32'h38632800;
      109511: inst = 32'h38842800;
      109512: inst = 32'h10a00001;
      109513: inst = 32'hca0abcd;
      109514: inst = 32'h13e00001;
      109515: inst = 32'hfe0d96a;
      109516: inst = 32'h5be00000;
      109517: inst = 32'h8c50000;
      109518: inst = 32'h24612800;
      109519: inst = 32'h10a00000;
      109520: inst = 32'hca00017;
      109521: inst = 32'h24822800;
      109522: inst = 32'h10a00000;
      109523: inst = 32'hca00004;
      109524: inst = 32'h38632800;
      109525: inst = 32'h38842800;
      109526: inst = 32'h10a00001;
      109527: inst = 32'hca0abdb;
      109528: inst = 32'h13e00001;
      109529: inst = 32'hfe0d96a;
      109530: inst = 32'h5be00000;
      109531: inst = 32'h8c50000;
      109532: inst = 32'h24612800;
      109533: inst = 32'h10a00000;
      109534: inst = 32'hca00017;
      109535: inst = 32'h24822800;
      109536: inst = 32'h10a00000;
      109537: inst = 32'hca00004;
      109538: inst = 32'h38632800;
      109539: inst = 32'h38842800;
      109540: inst = 32'h10a00001;
      109541: inst = 32'hca0abe9;
      109542: inst = 32'h13e00001;
      109543: inst = 32'hfe0d96a;
      109544: inst = 32'h5be00000;
      109545: inst = 32'h8c50000;
      109546: inst = 32'h24612800;
      109547: inst = 32'h10a00000;
      109548: inst = 32'hca00017;
      109549: inst = 32'h24822800;
      109550: inst = 32'h10a00000;
      109551: inst = 32'hca00004;
      109552: inst = 32'h38632800;
      109553: inst = 32'h38842800;
      109554: inst = 32'h10a00001;
      109555: inst = 32'hca0abf7;
      109556: inst = 32'h13e00001;
      109557: inst = 32'hfe0d96a;
      109558: inst = 32'h5be00000;
      109559: inst = 32'h8c50000;
      109560: inst = 32'h24612800;
      109561: inst = 32'h10a00000;
      109562: inst = 32'hca00017;
      109563: inst = 32'h24822800;
      109564: inst = 32'h10a00000;
      109565: inst = 32'hca00004;
      109566: inst = 32'h38632800;
      109567: inst = 32'h38842800;
      109568: inst = 32'h10a00001;
      109569: inst = 32'hca0ac05;
      109570: inst = 32'h13e00001;
      109571: inst = 32'hfe0d96a;
      109572: inst = 32'h5be00000;
      109573: inst = 32'h8c50000;
      109574: inst = 32'h24612800;
      109575: inst = 32'h10a00000;
      109576: inst = 32'hca00017;
      109577: inst = 32'h24822800;
      109578: inst = 32'h10a00000;
      109579: inst = 32'hca00004;
      109580: inst = 32'h38632800;
      109581: inst = 32'h38842800;
      109582: inst = 32'h10a00001;
      109583: inst = 32'hca0ac13;
      109584: inst = 32'h13e00001;
      109585: inst = 32'hfe0d96a;
      109586: inst = 32'h5be00000;
      109587: inst = 32'h8c50000;
      109588: inst = 32'h24612800;
      109589: inst = 32'h10a00000;
      109590: inst = 32'hca00017;
      109591: inst = 32'h24822800;
      109592: inst = 32'h10a00000;
      109593: inst = 32'hca00004;
      109594: inst = 32'h38632800;
      109595: inst = 32'h38842800;
      109596: inst = 32'h10a00001;
      109597: inst = 32'hca0ac21;
      109598: inst = 32'h13e00001;
      109599: inst = 32'hfe0d96a;
      109600: inst = 32'h5be00000;
      109601: inst = 32'h8c50000;
      109602: inst = 32'h24612800;
      109603: inst = 32'h10a00000;
      109604: inst = 32'hca00017;
      109605: inst = 32'h24822800;
      109606: inst = 32'h10a00000;
      109607: inst = 32'hca00004;
      109608: inst = 32'h38632800;
      109609: inst = 32'h38842800;
      109610: inst = 32'h10a00001;
      109611: inst = 32'hca0ac2f;
      109612: inst = 32'h13e00001;
      109613: inst = 32'hfe0d96a;
      109614: inst = 32'h5be00000;
      109615: inst = 32'h8c50000;
      109616: inst = 32'h24612800;
      109617: inst = 32'h10a00000;
      109618: inst = 32'hca00017;
      109619: inst = 32'h24822800;
      109620: inst = 32'h10a00000;
      109621: inst = 32'hca00004;
      109622: inst = 32'h38632800;
      109623: inst = 32'h38842800;
      109624: inst = 32'h10a00001;
      109625: inst = 32'hca0ac3d;
      109626: inst = 32'h13e00001;
      109627: inst = 32'hfe0d96a;
      109628: inst = 32'h5be00000;
      109629: inst = 32'h8c50000;
      109630: inst = 32'h24612800;
      109631: inst = 32'h10a00000;
      109632: inst = 32'hca00017;
      109633: inst = 32'h24822800;
      109634: inst = 32'h10a00000;
      109635: inst = 32'hca00004;
      109636: inst = 32'h38632800;
      109637: inst = 32'h38842800;
      109638: inst = 32'h10a00001;
      109639: inst = 32'hca0ac4b;
      109640: inst = 32'h13e00001;
      109641: inst = 32'hfe0d96a;
      109642: inst = 32'h5be00000;
      109643: inst = 32'h8c50000;
      109644: inst = 32'h24612800;
      109645: inst = 32'h10a00000;
      109646: inst = 32'hca00017;
      109647: inst = 32'h24822800;
      109648: inst = 32'h10a00000;
      109649: inst = 32'hca00004;
      109650: inst = 32'h38632800;
      109651: inst = 32'h38842800;
      109652: inst = 32'h10a00001;
      109653: inst = 32'hca0ac59;
      109654: inst = 32'h13e00001;
      109655: inst = 32'hfe0d96a;
      109656: inst = 32'h5be00000;
      109657: inst = 32'h8c50000;
      109658: inst = 32'h24612800;
      109659: inst = 32'h10a00000;
      109660: inst = 32'hca00017;
      109661: inst = 32'h24822800;
      109662: inst = 32'h10a00000;
      109663: inst = 32'hca00004;
      109664: inst = 32'h38632800;
      109665: inst = 32'h38842800;
      109666: inst = 32'h10a00001;
      109667: inst = 32'hca0ac67;
      109668: inst = 32'h13e00001;
      109669: inst = 32'hfe0d96a;
      109670: inst = 32'h5be00000;
      109671: inst = 32'h8c50000;
      109672: inst = 32'h24612800;
      109673: inst = 32'h10a00000;
      109674: inst = 32'hca00017;
      109675: inst = 32'h24822800;
      109676: inst = 32'h10a00000;
      109677: inst = 32'hca00004;
      109678: inst = 32'h38632800;
      109679: inst = 32'h38842800;
      109680: inst = 32'h10a00001;
      109681: inst = 32'hca0ac75;
      109682: inst = 32'h13e00001;
      109683: inst = 32'hfe0d96a;
      109684: inst = 32'h5be00000;
      109685: inst = 32'h8c50000;
      109686: inst = 32'h24612800;
      109687: inst = 32'h10a00000;
      109688: inst = 32'hca00017;
      109689: inst = 32'h24822800;
      109690: inst = 32'h10a00000;
      109691: inst = 32'hca00004;
      109692: inst = 32'h38632800;
      109693: inst = 32'h38842800;
      109694: inst = 32'h10a00001;
      109695: inst = 32'hca0ac83;
      109696: inst = 32'h13e00001;
      109697: inst = 32'hfe0d96a;
      109698: inst = 32'h5be00000;
      109699: inst = 32'h8c50000;
      109700: inst = 32'h24612800;
      109701: inst = 32'h10a00000;
      109702: inst = 32'hca00017;
      109703: inst = 32'h24822800;
      109704: inst = 32'h10a00000;
      109705: inst = 32'hca00004;
      109706: inst = 32'h38632800;
      109707: inst = 32'h38842800;
      109708: inst = 32'h10a00001;
      109709: inst = 32'hca0ac91;
      109710: inst = 32'h13e00001;
      109711: inst = 32'hfe0d96a;
      109712: inst = 32'h5be00000;
      109713: inst = 32'h8c50000;
      109714: inst = 32'h24612800;
      109715: inst = 32'h10a00000;
      109716: inst = 32'hca00017;
      109717: inst = 32'h24822800;
      109718: inst = 32'h10a00000;
      109719: inst = 32'hca00004;
      109720: inst = 32'h38632800;
      109721: inst = 32'h38842800;
      109722: inst = 32'h10a00001;
      109723: inst = 32'hca0ac9f;
      109724: inst = 32'h13e00001;
      109725: inst = 32'hfe0d96a;
      109726: inst = 32'h5be00000;
      109727: inst = 32'h8c50000;
      109728: inst = 32'h24612800;
      109729: inst = 32'h10a00000;
      109730: inst = 32'hca00017;
      109731: inst = 32'h24822800;
      109732: inst = 32'h10a00000;
      109733: inst = 32'hca00004;
      109734: inst = 32'h38632800;
      109735: inst = 32'h38842800;
      109736: inst = 32'h10a00001;
      109737: inst = 32'hca0acad;
      109738: inst = 32'h13e00001;
      109739: inst = 32'hfe0d96a;
      109740: inst = 32'h5be00000;
      109741: inst = 32'h8c50000;
      109742: inst = 32'h24612800;
      109743: inst = 32'h10a00000;
      109744: inst = 32'hca00017;
      109745: inst = 32'h24822800;
      109746: inst = 32'h10a00000;
      109747: inst = 32'hca00004;
      109748: inst = 32'h38632800;
      109749: inst = 32'h38842800;
      109750: inst = 32'h10a00001;
      109751: inst = 32'hca0acbb;
      109752: inst = 32'h13e00001;
      109753: inst = 32'hfe0d96a;
      109754: inst = 32'h5be00000;
      109755: inst = 32'h8c50000;
      109756: inst = 32'h24612800;
      109757: inst = 32'h10a00000;
      109758: inst = 32'hca00017;
      109759: inst = 32'h24822800;
      109760: inst = 32'h10a00000;
      109761: inst = 32'hca00004;
      109762: inst = 32'h38632800;
      109763: inst = 32'h38842800;
      109764: inst = 32'h10a00001;
      109765: inst = 32'hca0acc9;
      109766: inst = 32'h13e00001;
      109767: inst = 32'hfe0d96a;
      109768: inst = 32'h5be00000;
      109769: inst = 32'h8c50000;
      109770: inst = 32'h24612800;
      109771: inst = 32'h10a00000;
      109772: inst = 32'hca00017;
      109773: inst = 32'h24822800;
      109774: inst = 32'h10a00000;
      109775: inst = 32'hca00004;
      109776: inst = 32'h38632800;
      109777: inst = 32'h38842800;
      109778: inst = 32'h10a00001;
      109779: inst = 32'hca0acd7;
      109780: inst = 32'h13e00001;
      109781: inst = 32'hfe0d96a;
      109782: inst = 32'h5be00000;
      109783: inst = 32'h8c50000;
      109784: inst = 32'h24612800;
      109785: inst = 32'h10a00000;
      109786: inst = 32'hca00017;
      109787: inst = 32'h24822800;
      109788: inst = 32'h10a00000;
      109789: inst = 32'hca00004;
      109790: inst = 32'h38632800;
      109791: inst = 32'h38842800;
      109792: inst = 32'h10a00001;
      109793: inst = 32'hca0ace5;
      109794: inst = 32'h13e00001;
      109795: inst = 32'hfe0d96a;
      109796: inst = 32'h5be00000;
      109797: inst = 32'h8c50000;
      109798: inst = 32'h24612800;
      109799: inst = 32'h10a00000;
      109800: inst = 32'hca00017;
      109801: inst = 32'h24822800;
      109802: inst = 32'h10a00000;
      109803: inst = 32'hca00004;
      109804: inst = 32'h38632800;
      109805: inst = 32'h38842800;
      109806: inst = 32'h10a00001;
      109807: inst = 32'hca0acf3;
      109808: inst = 32'h13e00001;
      109809: inst = 32'hfe0d96a;
      109810: inst = 32'h5be00000;
      109811: inst = 32'h8c50000;
      109812: inst = 32'h24612800;
      109813: inst = 32'h10a00000;
      109814: inst = 32'hca00017;
      109815: inst = 32'h24822800;
      109816: inst = 32'h10a00000;
      109817: inst = 32'hca00004;
      109818: inst = 32'h38632800;
      109819: inst = 32'h38842800;
      109820: inst = 32'h10a00001;
      109821: inst = 32'hca0ad01;
      109822: inst = 32'h13e00001;
      109823: inst = 32'hfe0d96a;
      109824: inst = 32'h5be00000;
      109825: inst = 32'h8c50000;
      109826: inst = 32'h24612800;
      109827: inst = 32'h10a00000;
      109828: inst = 32'hca00017;
      109829: inst = 32'h24822800;
      109830: inst = 32'h10a00000;
      109831: inst = 32'hca00004;
      109832: inst = 32'h38632800;
      109833: inst = 32'h38842800;
      109834: inst = 32'h10a00001;
      109835: inst = 32'hca0ad0f;
      109836: inst = 32'h13e00001;
      109837: inst = 32'hfe0d96a;
      109838: inst = 32'h5be00000;
      109839: inst = 32'h8c50000;
      109840: inst = 32'h24612800;
      109841: inst = 32'h10a00000;
      109842: inst = 32'hca00017;
      109843: inst = 32'h24822800;
      109844: inst = 32'h10a00000;
      109845: inst = 32'hca00004;
      109846: inst = 32'h38632800;
      109847: inst = 32'h38842800;
      109848: inst = 32'h10a00001;
      109849: inst = 32'hca0ad1d;
      109850: inst = 32'h13e00001;
      109851: inst = 32'hfe0d96a;
      109852: inst = 32'h5be00000;
      109853: inst = 32'h8c50000;
      109854: inst = 32'h24612800;
      109855: inst = 32'h10a00000;
      109856: inst = 32'hca00017;
      109857: inst = 32'h24822800;
      109858: inst = 32'h10a00000;
      109859: inst = 32'hca00004;
      109860: inst = 32'h38632800;
      109861: inst = 32'h38842800;
      109862: inst = 32'h10a00001;
      109863: inst = 32'hca0ad2b;
      109864: inst = 32'h13e00001;
      109865: inst = 32'hfe0d96a;
      109866: inst = 32'h5be00000;
      109867: inst = 32'h8c50000;
      109868: inst = 32'h24612800;
      109869: inst = 32'h10a00000;
      109870: inst = 32'hca00017;
      109871: inst = 32'h24822800;
      109872: inst = 32'h10a00000;
      109873: inst = 32'hca00004;
      109874: inst = 32'h38632800;
      109875: inst = 32'h38842800;
      109876: inst = 32'h10a00001;
      109877: inst = 32'hca0ad39;
      109878: inst = 32'h13e00001;
      109879: inst = 32'hfe0d96a;
      109880: inst = 32'h5be00000;
      109881: inst = 32'h8c50000;
      109882: inst = 32'h24612800;
      109883: inst = 32'h10a00000;
      109884: inst = 32'hca00017;
      109885: inst = 32'h24822800;
      109886: inst = 32'h10a00000;
      109887: inst = 32'hca00004;
      109888: inst = 32'h38632800;
      109889: inst = 32'h38842800;
      109890: inst = 32'h10a00001;
      109891: inst = 32'hca0ad47;
      109892: inst = 32'h13e00001;
      109893: inst = 32'hfe0d96a;
      109894: inst = 32'h5be00000;
      109895: inst = 32'h8c50000;
      109896: inst = 32'h24612800;
      109897: inst = 32'h10a00000;
      109898: inst = 32'hca00017;
      109899: inst = 32'h24822800;
      109900: inst = 32'h10a00000;
      109901: inst = 32'hca00004;
      109902: inst = 32'h38632800;
      109903: inst = 32'h38842800;
      109904: inst = 32'h10a00001;
      109905: inst = 32'hca0ad55;
      109906: inst = 32'h13e00001;
      109907: inst = 32'hfe0d96a;
      109908: inst = 32'h5be00000;
      109909: inst = 32'h8c50000;
      109910: inst = 32'h24612800;
      109911: inst = 32'h10a00000;
      109912: inst = 32'hca00017;
      109913: inst = 32'h24822800;
      109914: inst = 32'h10a00000;
      109915: inst = 32'hca00004;
      109916: inst = 32'h38632800;
      109917: inst = 32'h38842800;
      109918: inst = 32'h10a00001;
      109919: inst = 32'hca0ad63;
      109920: inst = 32'h13e00001;
      109921: inst = 32'hfe0d96a;
      109922: inst = 32'h5be00000;
      109923: inst = 32'h8c50000;
      109924: inst = 32'h24612800;
      109925: inst = 32'h10a00000;
      109926: inst = 32'hca00017;
      109927: inst = 32'h24822800;
      109928: inst = 32'h10a00000;
      109929: inst = 32'hca00004;
      109930: inst = 32'h38632800;
      109931: inst = 32'h38842800;
      109932: inst = 32'h10a00001;
      109933: inst = 32'hca0ad71;
      109934: inst = 32'h13e00001;
      109935: inst = 32'hfe0d96a;
      109936: inst = 32'h5be00000;
      109937: inst = 32'h8c50000;
      109938: inst = 32'h24612800;
      109939: inst = 32'h10a00000;
      109940: inst = 32'hca00017;
      109941: inst = 32'h24822800;
      109942: inst = 32'h10a00000;
      109943: inst = 32'hca00004;
      109944: inst = 32'h38632800;
      109945: inst = 32'h38842800;
      109946: inst = 32'h10a00001;
      109947: inst = 32'hca0ad7f;
      109948: inst = 32'h13e00001;
      109949: inst = 32'hfe0d96a;
      109950: inst = 32'h5be00000;
      109951: inst = 32'h8c50000;
      109952: inst = 32'h24612800;
      109953: inst = 32'h10a00000;
      109954: inst = 32'hca00017;
      109955: inst = 32'h24822800;
      109956: inst = 32'h10a00000;
      109957: inst = 32'hca00004;
      109958: inst = 32'h38632800;
      109959: inst = 32'h38842800;
      109960: inst = 32'h10a00001;
      109961: inst = 32'hca0ad8d;
      109962: inst = 32'h13e00001;
      109963: inst = 32'hfe0d96a;
      109964: inst = 32'h5be00000;
      109965: inst = 32'h8c50000;
      109966: inst = 32'h24612800;
      109967: inst = 32'h10a00000;
      109968: inst = 32'hca00017;
      109969: inst = 32'h24822800;
      109970: inst = 32'h10a00000;
      109971: inst = 32'hca00004;
      109972: inst = 32'h38632800;
      109973: inst = 32'h38842800;
      109974: inst = 32'h10a00001;
      109975: inst = 32'hca0ad9b;
      109976: inst = 32'h13e00001;
      109977: inst = 32'hfe0d96a;
      109978: inst = 32'h5be00000;
      109979: inst = 32'h8c50000;
      109980: inst = 32'h24612800;
      109981: inst = 32'h10a00000;
      109982: inst = 32'hca00017;
      109983: inst = 32'h24822800;
      109984: inst = 32'h10a00000;
      109985: inst = 32'hca00004;
      109986: inst = 32'h38632800;
      109987: inst = 32'h38842800;
      109988: inst = 32'h10a00001;
      109989: inst = 32'hca0ada9;
      109990: inst = 32'h13e00001;
      109991: inst = 32'hfe0d96a;
      109992: inst = 32'h5be00000;
      109993: inst = 32'h8c50000;
      109994: inst = 32'h24612800;
      109995: inst = 32'h10a00000;
      109996: inst = 32'hca00017;
      109997: inst = 32'h24822800;
      109998: inst = 32'h10a00000;
      109999: inst = 32'hca00004;
      110000: inst = 32'h38632800;
      110001: inst = 32'h38842800;
      110002: inst = 32'h10a00001;
      110003: inst = 32'hca0adb7;
      110004: inst = 32'h13e00001;
      110005: inst = 32'hfe0d96a;
      110006: inst = 32'h5be00000;
      110007: inst = 32'h8c50000;
      110008: inst = 32'h24612800;
      110009: inst = 32'h10a00000;
      110010: inst = 32'hca00017;
      110011: inst = 32'h24822800;
      110012: inst = 32'h10a00000;
      110013: inst = 32'hca00004;
      110014: inst = 32'h38632800;
      110015: inst = 32'h38842800;
      110016: inst = 32'h10a00001;
      110017: inst = 32'hca0adc5;
      110018: inst = 32'h13e00001;
      110019: inst = 32'hfe0d96a;
      110020: inst = 32'h5be00000;
      110021: inst = 32'h8c50000;
      110022: inst = 32'h24612800;
      110023: inst = 32'h10a00000;
      110024: inst = 32'hca00017;
      110025: inst = 32'h24822800;
      110026: inst = 32'h10a00000;
      110027: inst = 32'hca00004;
      110028: inst = 32'h38632800;
      110029: inst = 32'h38842800;
      110030: inst = 32'h10a00001;
      110031: inst = 32'hca0add3;
      110032: inst = 32'h13e00001;
      110033: inst = 32'hfe0d96a;
      110034: inst = 32'h5be00000;
      110035: inst = 32'h8c50000;
      110036: inst = 32'h24612800;
      110037: inst = 32'h10a00000;
      110038: inst = 32'hca00017;
      110039: inst = 32'h24822800;
      110040: inst = 32'h10a00000;
      110041: inst = 32'hca00004;
      110042: inst = 32'h38632800;
      110043: inst = 32'h38842800;
      110044: inst = 32'h10a00001;
      110045: inst = 32'hca0ade1;
      110046: inst = 32'h13e00001;
      110047: inst = 32'hfe0d96a;
      110048: inst = 32'h5be00000;
      110049: inst = 32'h8c50000;
      110050: inst = 32'h24612800;
      110051: inst = 32'h10a00000;
      110052: inst = 32'hca00017;
      110053: inst = 32'h24822800;
      110054: inst = 32'h10a00000;
      110055: inst = 32'hca00004;
      110056: inst = 32'h38632800;
      110057: inst = 32'h38842800;
      110058: inst = 32'h10a00001;
      110059: inst = 32'hca0adef;
      110060: inst = 32'h13e00001;
      110061: inst = 32'hfe0d96a;
      110062: inst = 32'h5be00000;
      110063: inst = 32'h8c50000;
      110064: inst = 32'h24612800;
      110065: inst = 32'h10a00000;
      110066: inst = 32'hca00017;
      110067: inst = 32'h24822800;
      110068: inst = 32'h10a00000;
      110069: inst = 32'hca00004;
      110070: inst = 32'h38632800;
      110071: inst = 32'h38842800;
      110072: inst = 32'h10a00001;
      110073: inst = 32'hca0adfd;
      110074: inst = 32'h13e00001;
      110075: inst = 32'hfe0d96a;
      110076: inst = 32'h5be00000;
      110077: inst = 32'h8c50000;
      110078: inst = 32'h24612800;
      110079: inst = 32'h10a00000;
      110080: inst = 32'hca00017;
      110081: inst = 32'h24822800;
      110082: inst = 32'h10a00000;
      110083: inst = 32'hca00004;
      110084: inst = 32'h38632800;
      110085: inst = 32'h38842800;
      110086: inst = 32'h10a00001;
      110087: inst = 32'hca0ae0b;
      110088: inst = 32'h13e00001;
      110089: inst = 32'hfe0d96a;
      110090: inst = 32'h5be00000;
      110091: inst = 32'h8c50000;
      110092: inst = 32'h24612800;
      110093: inst = 32'h10a00000;
      110094: inst = 32'hca00017;
      110095: inst = 32'h24822800;
      110096: inst = 32'h10a00000;
      110097: inst = 32'hca00004;
      110098: inst = 32'h38632800;
      110099: inst = 32'h38842800;
      110100: inst = 32'h10a00001;
      110101: inst = 32'hca0ae19;
      110102: inst = 32'h13e00001;
      110103: inst = 32'hfe0d96a;
      110104: inst = 32'h5be00000;
      110105: inst = 32'h8c50000;
      110106: inst = 32'h24612800;
      110107: inst = 32'h10a00000;
      110108: inst = 32'hca00017;
      110109: inst = 32'h24822800;
      110110: inst = 32'h10a00000;
      110111: inst = 32'hca00004;
      110112: inst = 32'h38632800;
      110113: inst = 32'h38842800;
      110114: inst = 32'h10a00001;
      110115: inst = 32'hca0ae27;
      110116: inst = 32'h13e00001;
      110117: inst = 32'hfe0d96a;
      110118: inst = 32'h5be00000;
      110119: inst = 32'h8c50000;
      110120: inst = 32'h24612800;
      110121: inst = 32'h10a00000;
      110122: inst = 32'hca00017;
      110123: inst = 32'h24822800;
      110124: inst = 32'h10a00000;
      110125: inst = 32'hca00004;
      110126: inst = 32'h38632800;
      110127: inst = 32'h38842800;
      110128: inst = 32'h10a00001;
      110129: inst = 32'hca0ae35;
      110130: inst = 32'h13e00001;
      110131: inst = 32'hfe0d96a;
      110132: inst = 32'h5be00000;
      110133: inst = 32'h8c50000;
      110134: inst = 32'h24612800;
      110135: inst = 32'h10a00000;
      110136: inst = 32'hca00017;
      110137: inst = 32'h24822800;
      110138: inst = 32'h10a00000;
      110139: inst = 32'hca00004;
      110140: inst = 32'h38632800;
      110141: inst = 32'h38842800;
      110142: inst = 32'h10a00001;
      110143: inst = 32'hca0ae43;
      110144: inst = 32'h13e00001;
      110145: inst = 32'hfe0d96a;
      110146: inst = 32'h5be00000;
      110147: inst = 32'h8c50000;
      110148: inst = 32'h24612800;
      110149: inst = 32'h10a00000;
      110150: inst = 32'hca00017;
      110151: inst = 32'h24822800;
      110152: inst = 32'h10a00000;
      110153: inst = 32'hca00004;
      110154: inst = 32'h38632800;
      110155: inst = 32'h38842800;
      110156: inst = 32'h10a00001;
      110157: inst = 32'hca0ae51;
      110158: inst = 32'h13e00001;
      110159: inst = 32'hfe0d96a;
      110160: inst = 32'h5be00000;
      110161: inst = 32'h8c50000;
      110162: inst = 32'h24612800;
      110163: inst = 32'h10a00000;
      110164: inst = 32'hca00017;
      110165: inst = 32'h24822800;
      110166: inst = 32'h10a00000;
      110167: inst = 32'hca00004;
      110168: inst = 32'h38632800;
      110169: inst = 32'h38842800;
      110170: inst = 32'h10a00001;
      110171: inst = 32'hca0ae5f;
      110172: inst = 32'h13e00001;
      110173: inst = 32'hfe0d96a;
      110174: inst = 32'h5be00000;
      110175: inst = 32'h8c50000;
      110176: inst = 32'h24612800;
      110177: inst = 32'h10a00000;
      110178: inst = 32'hca00017;
      110179: inst = 32'h24822800;
      110180: inst = 32'h10a00000;
      110181: inst = 32'hca00004;
      110182: inst = 32'h38632800;
      110183: inst = 32'h38842800;
      110184: inst = 32'h10a00001;
      110185: inst = 32'hca0ae6d;
      110186: inst = 32'h13e00001;
      110187: inst = 32'hfe0d96a;
      110188: inst = 32'h5be00000;
      110189: inst = 32'h8c50000;
      110190: inst = 32'h24612800;
      110191: inst = 32'h10a00000;
      110192: inst = 32'hca00017;
      110193: inst = 32'h24822800;
      110194: inst = 32'h10a00000;
      110195: inst = 32'hca00004;
      110196: inst = 32'h38632800;
      110197: inst = 32'h38842800;
      110198: inst = 32'h10a00001;
      110199: inst = 32'hca0ae7b;
      110200: inst = 32'h13e00001;
      110201: inst = 32'hfe0d96a;
      110202: inst = 32'h5be00000;
      110203: inst = 32'h8c50000;
      110204: inst = 32'h24612800;
      110205: inst = 32'h10a00000;
      110206: inst = 32'hca00017;
      110207: inst = 32'h24822800;
      110208: inst = 32'h10a00000;
      110209: inst = 32'hca00004;
      110210: inst = 32'h38632800;
      110211: inst = 32'h38842800;
      110212: inst = 32'h10a00001;
      110213: inst = 32'hca0ae89;
      110214: inst = 32'h13e00001;
      110215: inst = 32'hfe0d96a;
      110216: inst = 32'h5be00000;
      110217: inst = 32'h8c50000;
      110218: inst = 32'h24612800;
      110219: inst = 32'h10a00000;
      110220: inst = 32'hca00017;
      110221: inst = 32'h24822800;
      110222: inst = 32'h10a00000;
      110223: inst = 32'hca00004;
      110224: inst = 32'h38632800;
      110225: inst = 32'h38842800;
      110226: inst = 32'h10a00001;
      110227: inst = 32'hca0ae97;
      110228: inst = 32'h13e00001;
      110229: inst = 32'hfe0d96a;
      110230: inst = 32'h5be00000;
      110231: inst = 32'h8c50000;
      110232: inst = 32'h24612800;
      110233: inst = 32'h10a00000;
      110234: inst = 32'hca00017;
      110235: inst = 32'h24822800;
      110236: inst = 32'h10a00000;
      110237: inst = 32'hca00004;
      110238: inst = 32'h38632800;
      110239: inst = 32'h38842800;
      110240: inst = 32'h10a00001;
      110241: inst = 32'hca0aea5;
      110242: inst = 32'h13e00001;
      110243: inst = 32'hfe0d96a;
      110244: inst = 32'h5be00000;
      110245: inst = 32'h8c50000;
      110246: inst = 32'h24612800;
      110247: inst = 32'h10a00000;
      110248: inst = 32'hca00017;
      110249: inst = 32'h24822800;
      110250: inst = 32'h10a00000;
      110251: inst = 32'hca00004;
      110252: inst = 32'h38632800;
      110253: inst = 32'h38842800;
      110254: inst = 32'h10a00001;
      110255: inst = 32'hca0aeb3;
      110256: inst = 32'h13e00001;
      110257: inst = 32'hfe0d96a;
      110258: inst = 32'h5be00000;
      110259: inst = 32'h8c50000;
      110260: inst = 32'h24612800;
      110261: inst = 32'h10a00000;
      110262: inst = 32'hca00017;
      110263: inst = 32'h24822800;
      110264: inst = 32'h10a00000;
      110265: inst = 32'hca00004;
      110266: inst = 32'h38632800;
      110267: inst = 32'h38842800;
      110268: inst = 32'h10a00001;
      110269: inst = 32'hca0aec1;
      110270: inst = 32'h13e00001;
      110271: inst = 32'hfe0d96a;
      110272: inst = 32'h5be00000;
      110273: inst = 32'h8c50000;
      110274: inst = 32'h24612800;
      110275: inst = 32'h10a00000;
      110276: inst = 32'hca00017;
      110277: inst = 32'h24822800;
      110278: inst = 32'h10a00000;
      110279: inst = 32'hca00004;
      110280: inst = 32'h38632800;
      110281: inst = 32'h38842800;
      110282: inst = 32'h10a00001;
      110283: inst = 32'hca0aecf;
      110284: inst = 32'h13e00001;
      110285: inst = 32'hfe0d96a;
      110286: inst = 32'h5be00000;
      110287: inst = 32'h8c50000;
      110288: inst = 32'h24612800;
      110289: inst = 32'h10a00000;
      110290: inst = 32'hca00017;
      110291: inst = 32'h24822800;
      110292: inst = 32'h10a00000;
      110293: inst = 32'hca00004;
      110294: inst = 32'h38632800;
      110295: inst = 32'h38842800;
      110296: inst = 32'h10a00001;
      110297: inst = 32'hca0aedd;
      110298: inst = 32'h13e00001;
      110299: inst = 32'hfe0d96a;
      110300: inst = 32'h5be00000;
      110301: inst = 32'h8c50000;
      110302: inst = 32'h24612800;
      110303: inst = 32'h10a00000;
      110304: inst = 32'hca00017;
      110305: inst = 32'h24822800;
      110306: inst = 32'h10a00000;
      110307: inst = 32'hca00004;
      110308: inst = 32'h38632800;
      110309: inst = 32'h38842800;
      110310: inst = 32'h10a00001;
      110311: inst = 32'hca0aeeb;
      110312: inst = 32'h13e00001;
      110313: inst = 32'hfe0d96a;
      110314: inst = 32'h5be00000;
      110315: inst = 32'h8c50000;
      110316: inst = 32'h24612800;
      110317: inst = 32'h10a00000;
      110318: inst = 32'hca00017;
      110319: inst = 32'h24822800;
      110320: inst = 32'h10a00000;
      110321: inst = 32'hca00004;
      110322: inst = 32'h38632800;
      110323: inst = 32'h38842800;
      110324: inst = 32'h10a00001;
      110325: inst = 32'hca0aef9;
      110326: inst = 32'h13e00001;
      110327: inst = 32'hfe0d96a;
      110328: inst = 32'h5be00000;
      110329: inst = 32'h8c50000;
      110330: inst = 32'h24612800;
      110331: inst = 32'h10a00000;
      110332: inst = 32'hca00017;
      110333: inst = 32'h24822800;
      110334: inst = 32'h10a00000;
      110335: inst = 32'hca00004;
      110336: inst = 32'h38632800;
      110337: inst = 32'h38842800;
      110338: inst = 32'h10a00001;
      110339: inst = 32'hca0af07;
      110340: inst = 32'h13e00001;
      110341: inst = 32'hfe0d96a;
      110342: inst = 32'h5be00000;
      110343: inst = 32'h8c50000;
      110344: inst = 32'h24612800;
      110345: inst = 32'h10a00000;
      110346: inst = 32'hca00017;
      110347: inst = 32'h24822800;
      110348: inst = 32'h10a00000;
      110349: inst = 32'hca00004;
      110350: inst = 32'h38632800;
      110351: inst = 32'h38842800;
      110352: inst = 32'h10a00001;
      110353: inst = 32'hca0af15;
      110354: inst = 32'h13e00001;
      110355: inst = 32'hfe0d96a;
      110356: inst = 32'h5be00000;
      110357: inst = 32'h8c50000;
      110358: inst = 32'h24612800;
      110359: inst = 32'h10a00000;
      110360: inst = 32'hca00017;
      110361: inst = 32'h24822800;
      110362: inst = 32'h10a00000;
      110363: inst = 32'hca00004;
      110364: inst = 32'h38632800;
      110365: inst = 32'h38842800;
      110366: inst = 32'h10a00001;
      110367: inst = 32'hca0af23;
      110368: inst = 32'h13e00001;
      110369: inst = 32'hfe0d96a;
      110370: inst = 32'h5be00000;
      110371: inst = 32'h8c50000;
      110372: inst = 32'h24612800;
      110373: inst = 32'h10a00000;
      110374: inst = 32'hca00017;
      110375: inst = 32'h24822800;
      110376: inst = 32'h10a00000;
      110377: inst = 32'hca00004;
      110378: inst = 32'h38632800;
      110379: inst = 32'h38842800;
      110380: inst = 32'h10a00001;
      110381: inst = 32'hca0af31;
      110382: inst = 32'h13e00001;
      110383: inst = 32'hfe0d96a;
      110384: inst = 32'h5be00000;
      110385: inst = 32'h8c50000;
      110386: inst = 32'h24612800;
      110387: inst = 32'h10a00000;
      110388: inst = 32'hca00017;
      110389: inst = 32'h24822800;
      110390: inst = 32'h10a00000;
      110391: inst = 32'hca00004;
      110392: inst = 32'h38632800;
      110393: inst = 32'h38842800;
      110394: inst = 32'h10a00001;
      110395: inst = 32'hca0af3f;
      110396: inst = 32'h13e00001;
      110397: inst = 32'hfe0d96a;
      110398: inst = 32'h5be00000;
      110399: inst = 32'h8c50000;
      110400: inst = 32'h24612800;
      110401: inst = 32'h10a00000;
      110402: inst = 32'hca00017;
      110403: inst = 32'h24822800;
      110404: inst = 32'h10a00000;
      110405: inst = 32'hca00004;
      110406: inst = 32'h38632800;
      110407: inst = 32'h38842800;
      110408: inst = 32'h10a00001;
      110409: inst = 32'hca0af4d;
      110410: inst = 32'h13e00001;
      110411: inst = 32'hfe0d96a;
      110412: inst = 32'h5be00000;
      110413: inst = 32'h8c50000;
      110414: inst = 32'h24612800;
      110415: inst = 32'h10a00000;
      110416: inst = 32'hca00017;
      110417: inst = 32'h24822800;
      110418: inst = 32'h10a00000;
      110419: inst = 32'hca00004;
      110420: inst = 32'h38632800;
      110421: inst = 32'h38842800;
      110422: inst = 32'h10a00001;
      110423: inst = 32'hca0af5b;
      110424: inst = 32'h13e00001;
      110425: inst = 32'hfe0d96a;
      110426: inst = 32'h5be00000;
      110427: inst = 32'h8c50000;
      110428: inst = 32'h24612800;
      110429: inst = 32'h10a00000;
      110430: inst = 32'hca00017;
      110431: inst = 32'h24822800;
      110432: inst = 32'h10a00000;
      110433: inst = 32'hca00004;
      110434: inst = 32'h38632800;
      110435: inst = 32'h38842800;
      110436: inst = 32'h10a00001;
      110437: inst = 32'hca0af69;
      110438: inst = 32'h13e00001;
      110439: inst = 32'hfe0d96a;
      110440: inst = 32'h5be00000;
      110441: inst = 32'h8c50000;
      110442: inst = 32'h24612800;
      110443: inst = 32'h10a00000;
      110444: inst = 32'hca00018;
      110445: inst = 32'h24822800;
      110446: inst = 32'h10a00000;
      110447: inst = 32'hca00004;
      110448: inst = 32'h38632800;
      110449: inst = 32'h38842800;
      110450: inst = 32'h10a00001;
      110451: inst = 32'hca0af77;
      110452: inst = 32'h13e00001;
      110453: inst = 32'hfe0d96a;
      110454: inst = 32'h5be00000;
      110455: inst = 32'h8c50000;
      110456: inst = 32'h24612800;
      110457: inst = 32'h10a00000;
      110458: inst = 32'hca00018;
      110459: inst = 32'h24822800;
      110460: inst = 32'h10a00000;
      110461: inst = 32'hca00004;
      110462: inst = 32'h38632800;
      110463: inst = 32'h38842800;
      110464: inst = 32'h10a00001;
      110465: inst = 32'hca0af85;
      110466: inst = 32'h13e00001;
      110467: inst = 32'hfe0d96a;
      110468: inst = 32'h5be00000;
      110469: inst = 32'h8c50000;
      110470: inst = 32'h24612800;
      110471: inst = 32'h10a00000;
      110472: inst = 32'hca00018;
      110473: inst = 32'h24822800;
      110474: inst = 32'h10a00000;
      110475: inst = 32'hca00004;
      110476: inst = 32'h38632800;
      110477: inst = 32'h38842800;
      110478: inst = 32'h10a00001;
      110479: inst = 32'hca0af93;
      110480: inst = 32'h13e00001;
      110481: inst = 32'hfe0d96a;
      110482: inst = 32'h5be00000;
      110483: inst = 32'h8c50000;
      110484: inst = 32'h24612800;
      110485: inst = 32'h10a00000;
      110486: inst = 32'hca00018;
      110487: inst = 32'h24822800;
      110488: inst = 32'h10a00000;
      110489: inst = 32'hca00004;
      110490: inst = 32'h38632800;
      110491: inst = 32'h38842800;
      110492: inst = 32'h10a00001;
      110493: inst = 32'hca0afa1;
      110494: inst = 32'h13e00001;
      110495: inst = 32'hfe0d96a;
      110496: inst = 32'h5be00000;
      110497: inst = 32'h8c50000;
      110498: inst = 32'h24612800;
      110499: inst = 32'h10a00000;
      110500: inst = 32'hca00018;
      110501: inst = 32'h24822800;
      110502: inst = 32'h10a00000;
      110503: inst = 32'hca00004;
      110504: inst = 32'h38632800;
      110505: inst = 32'h38842800;
      110506: inst = 32'h10a00001;
      110507: inst = 32'hca0afaf;
      110508: inst = 32'h13e00001;
      110509: inst = 32'hfe0d96a;
      110510: inst = 32'h5be00000;
      110511: inst = 32'h8c50000;
      110512: inst = 32'h24612800;
      110513: inst = 32'h10a00000;
      110514: inst = 32'hca00018;
      110515: inst = 32'h24822800;
      110516: inst = 32'h10a00000;
      110517: inst = 32'hca00004;
      110518: inst = 32'h38632800;
      110519: inst = 32'h38842800;
      110520: inst = 32'h10a00001;
      110521: inst = 32'hca0afbd;
      110522: inst = 32'h13e00001;
      110523: inst = 32'hfe0d96a;
      110524: inst = 32'h5be00000;
      110525: inst = 32'h8c50000;
      110526: inst = 32'h24612800;
      110527: inst = 32'h10a00000;
      110528: inst = 32'hca00018;
      110529: inst = 32'h24822800;
      110530: inst = 32'h10a00000;
      110531: inst = 32'hca00004;
      110532: inst = 32'h38632800;
      110533: inst = 32'h38842800;
      110534: inst = 32'h10a00001;
      110535: inst = 32'hca0afcb;
      110536: inst = 32'h13e00001;
      110537: inst = 32'hfe0d96a;
      110538: inst = 32'h5be00000;
      110539: inst = 32'h8c50000;
      110540: inst = 32'h24612800;
      110541: inst = 32'h10a00000;
      110542: inst = 32'hca00018;
      110543: inst = 32'h24822800;
      110544: inst = 32'h10a00000;
      110545: inst = 32'hca00004;
      110546: inst = 32'h38632800;
      110547: inst = 32'h38842800;
      110548: inst = 32'h10a00001;
      110549: inst = 32'hca0afd9;
      110550: inst = 32'h13e00001;
      110551: inst = 32'hfe0d96a;
      110552: inst = 32'h5be00000;
      110553: inst = 32'h8c50000;
      110554: inst = 32'h24612800;
      110555: inst = 32'h10a00000;
      110556: inst = 32'hca00018;
      110557: inst = 32'h24822800;
      110558: inst = 32'h10a00000;
      110559: inst = 32'hca00004;
      110560: inst = 32'h38632800;
      110561: inst = 32'h38842800;
      110562: inst = 32'h10a00001;
      110563: inst = 32'hca0afe7;
      110564: inst = 32'h13e00001;
      110565: inst = 32'hfe0d96a;
      110566: inst = 32'h5be00000;
      110567: inst = 32'h8c50000;
      110568: inst = 32'h24612800;
      110569: inst = 32'h10a00000;
      110570: inst = 32'hca00018;
      110571: inst = 32'h24822800;
      110572: inst = 32'h10a00000;
      110573: inst = 32'hca00004;
      110574: inst = 32'h38632800;
      110575: inst = 32'h38842800;
      110576: inst = 32'h10a00001;
      110577: inst = 32'hca0aff5;
      110578: inst = 32'h13e00001;
      110579: inst = 32'hfe0d96a;
      110580: inst = 32'h5be00000;
      110581: inst = 32'h8c50000;
      110582: inst = 32'h24612800;
      110583: inst = 32'h10a00000;
      110584: inst = 32'hca00018;
      110585: inst = 32'h24822800;
      110586: inst = 32'h10a00000;
      110587: inst = 32'hca00004;
      110588: inst = 32'h38632800;
      110589: inst = 32'h38842800;
      110590: inst = 32'h10a00001;
      110591: inst = 32'hca0b003;
      110592: inst = 32'h13e00001;
      110593: inst = 32'hfe0d96a;
      110594: inst = 32'h5be00000;
      110595: inst = 32'h8c50000;
      110596: inst = 32'h24612800;
      110597: inst = 32'h10a00000;
      110598: inst = 32'hca00018;
      110599: inst = 32'h24822800;
      110600: inst = 32'h10a00000;
      110601: inst = 32'hca00004;
      110602: inst = 32'h38632800;
      110603: inst = 32'h38842800;
      110604: inst = 32'h10a00001;
      110605: inst = 32'hca0b011;
      110606: inst = 32'h13e00001;
      110607: inst = 32'hfe0d96a;
      110608: inst = 32'h5be00000;
      110609: inst = 32'h8c50000;
      110610: inst = 32'h24612800;
      110611: inst = 32'h10a00000;
      110612: inst = 32'hca00018;
      110613: inst = 32'h24822800;
      110614: inst = 32'h10a00000;
      110615: inst = 32'hca00004;
      110616: inst = 32'h38632800;
      110617: inst = 32'h38842800;
      110618: inst = 32'h10a00001;
      110619: inst = 32'hca0b01f;
      110620: inst = 32'h13e00001;
      110621: inst = 32'hfe0d96a;
      110622: inst = 32'h5be00000;
      110623: inst = 32'h8c50000;
      110624: inst = 32'h24612800;
      110625: inst = 32'h10a00000;
      110626: inst = 32'hca00018;
      110627: inst = 32'h24822800;
      110628: inst = 32'h10a00000;
      110629: inst = 32'hca00004;
      110630: inst = 32'h38632800;
      110631: inst = 32'h38842800;
      110632: inst = 32'h10a00001;
      110633: inst = 32'hca0b02d;
      110634: inst = 32'h13e00001;
      110635: inst = 32'hfe0d96a;
      110636: inst = 32'h5be00000;
      110637: inst = 32'h8c50000;
      110638: inst = 32'h24612800;
      110639: inst = 32'h10a00000;
      110640: inst = 32'hca00018;
      110641: inst = 32'h24822800;
      110642: inst = 32'h10a00000;
      110643: inst = 32'hca00004;
      110644: inst = 32'h38632800;
      110645: inst = 32'h38842800;
      110646: inst = 32'h10a00001;
      110647: inst = 32'hca0b03b;
      110648: inst = 32'h13e00001;
      110649: inst = 32'hfe0d96a;
      110650: inst = 32'h5be00000;
      110651: inst = 32'h8c50000;
      110652: inst = 32'h24612800;
      110653: inst = 32'h10a00000;
      110654: inst = 32'hca00018;
      110655: inst = 32'h24822800;
      110656: inst = 32'h10a00000;
      110657: inst = 32'hca00004;
      110658: inst = 32'h38632800;
      110659: inst = 32'h38842800;
      110660: inst = 32'h10a00001;
      110661: inst = 32'hca0b049;
      110662: inst = 32'h13e00001;
      110663: inst = 32'hfe0d96a;
      110664: inst = 32'h5be00000;
      110665: inst = 32'h8c50000;
      110666: inst = 32'h24612800;
      110667: inst = 32'h10a00000;
      110668: inst = 32'hca00018;
      110669: inst = 32'h24822800;
      110670: inst = 32'h10a00000;
      110671: inst = 32'hca00004;
      110672: inst = 32'h38632800;
      110673: inst = 32'h38842800;
      110674: inst = 32'h10a00001;
      110675: inst = 32'hca0b057;
      110676: inst = 32'h13e00001;
      110677: inst = 32'hfe0d96a;
      110678: inst = 32'h5be00000;
      110679: inst = 32'h8c50000;
      110680: inst = 32'h24612800;
      110681: inst = 32'h10a00000;
      110682: inst = 32'hca00018;
      110683: inst = 32'h24822800;
      110684: inst = 32'h10a00000;
      110685: inst = 32'hca00004;
      110686: inst = 32'h38632800;
      110687: inst = 32'h38842800;
      110688: inst = 32'h10a00001;
      110689: inst = 32'hca0b065;
      110690: inst = 32'h13e00001;
      110691: inst = 32'hfe0d96a;
      110692: inst = 32'h5be00000;
      110693: inst = 32'h8c50000;
      110694: inst = 32'h24612800;
      110695: inst = 32'h10a00000;
      110696: inst = 32'hca00018;
      110697: inst = 32'h24822800;
      110698: inst = 32'h10a00000;
      110699: inst = 32'hca00004;
      110700: inst = 32'h38632800;
      110701: inst = 32'h38842800;
      110702: inst = 32'h10a00001;
      110703: inst = 32'hca0b073;
      110704: inst = 32'h13e00001;
      110705: inst = 32'hfe0d96a;
      110706: inst = 32'h5be00000;
      110707: inst = 32'h8c50000;
      110708: inst = 32'h24612800;
      110709: inst = 32'h10a00000;
      110710: inst = 32'hca00018;
      110711: inst = 32'h24822800;
      110712: inst = 32'h10a00000;
      110713: inst = 32'hca00004;
      110714: inst = 32'h38632800;
      110715: inst = 32'h38842800;
      110716: inst = 32'h10a00001;
      110717: inst = 32'hca0b081;
      110718: inst = 32'h13e00001;
      110719: inst = 32'hfe0d96a;
      110720: inst = 32'h5be00000;
      110721: inst = 32'h8c50000;
      110722: inst = 32'h24612800;
      110723: inst = 32'h10a00000;
      110724: inst = 32'hca00018;
      110725: inst = 32'h24822800;
      110726: inst = 32'h10a00000;
      110727: inst = 32'hca00004;
      110728: inst = 32'h38632800;
      110729: inst = 32'h38842800;
      110730: inst = 32'h10a00001;
      110731: inst = 32'hca0b08f;
      110732: inst = 32'h13e00001;
      110733: inst = 32'hfe0d96a;
      110734: inst = 32'h5be00000;
      110735: inst = 32'h8c50000;
      110736: inst = 32'h24612800;
      110737: inst = 32'h10a00000;
      110738: inst = 32'hca00018;
      110739: inst = 32'h24822800;
      110740: inst = 32'h10a00000;
      110741: inst = 32'hca00004;
      110742: inst = 32'h38632800;
      110743: inst = 32'h38842800;
      110744: inst = 32'h10a00001;
      110745: inst = 32'hca0b09d;
      110746: inst = 32'h13e00001;
      110747: inst = 32'hfe0d96a;
      110748: inst = 32'h5be00000;
      110749: inst = 32'h8c50000;
      110750: inst = 32'h24612800;
      110751: inst = 32'h10a00000;
      110752: inst = 32'hca00018;
      110753: inst = 32'h24822800;
      110754: inst = 32'h10a00000;
      110755: inst = 32'hca00004;
      110756: inst = 32'h38632800;
      110757: inst = 32'h38842800;
      110758: inst = 32'h10a00001;
      110759: inst = 32'hca0b0ab;
      110760: inst = 32'h13e00001;
      110761: inst = 32'hfe0d96a;
      110762: inst = 32'h5be00000;
      110763: inst = 32'h8c50000;
      110764: inst = 32'h24612800;
      110765: inst = 32'h10a00000;
      110766: inst = 32'hca00018;
      110767: inst = 32'h24822800;
      110768: inst = 32'h10a00000;
      110769: inst = 32'hca00004;
      110770: inst = 32'h38632800;
      110771: inst = 32'h38842800;
      110772: inst = 32'h10a00001;
      110773: inst = 32'hca0b0b9;
      110774: inst = 32'h13e00001;
      110775: inst = 32'hfe0d96a;
      110776: inst = 32'h5be00000;
      110777: inst = 32'h8c50000;
      110778: inst = 32'h24612800;
      110779: inst = 32'h10a00000;
      110780: inst = 32'hca00018;
      110781: inst = 32'h24822800;
      110782: inst = 32'h10a00000;
      110783: inst = 32'hca00004;
      110784: inst = 32'h38632800;
      110785: inst = 32'h38842800;
      110786: inst = 32'h10a00001;
      110787: inst = 32'hca0b0c7;
      110788: inst = 32'h13e00001;
      110789: inst = 32'hfe0d96a;
      110790: inst = 32'h5be00000;
      110791: inst = 32'h8c50000;
      110792: inst = 32'h24612800;
      110793: inst = 32'h10a00000;
      110794: inst = 32'hca00018;
      110795: inst = 32'h24822800;
      110796: inst = 32'h10a00000;
      110797: inst = 32'hca00004;
      110798: inst = 32'h38632800;
      110799: inst = 32'h38842800;
      110800: inst = 32'h10a00001;
      110801: inst = 32'hca0b0d5;
      110802: inst = 32'h13e00001;
      110803: inst = 32'hfe0d96a;
      110804: inst = 32'h5be00000;
      110805: inst = 32'h8c50000;
      110806: inst = 32'h24612800;
      110807: inst = 32'h10a00000;
      110808: inst = 32'hca00018;
      110809: inst = 32'h24822800;
      110810: inst = 32'h10a00000;
      110811: inst = 32'hca00004;
      110812: inst = 32'h38632800;
      110813: inst = 32'h38842800;
      110814: inst = 32'h10a00001;
      110815: inst = 32'hca0b0e3;
      110816: inst = 32'h13e00001;
      110817: inst = 32'hfe0d96a;
      110818: inst = 32'h5be00000;
      110819: inst = 32'h8c50000;
      110820: inst = 32'h24612800;
      110821: inst = 32'h10a00000;
      110822: inst = 32'hca00018;
      110823: inst = 32'h24822800;
      110824: inst = 32'h10a00000;
      110825: inst = 32'hca00004;
      110826: inst = 32'h38632800;
      110827: inst = 32'h38842800;
      110828: inst = 32'h10a00001;
      110829: inst = 32'hca0b0f1;
      110830: inst = 32'h13e00001;
      110831: inst = 32'hfe0d96a;
      110832: inst = 32'h5be00000;
      110833: inst = 32'h8c50000;
      110834: inst = 32'h24612800;
      110835: inst = 32'h10a00000;
      110836: inst = 32'hca00018;
      110837: inst = 32'h24822800;
      110838: inst = 32'h10a00000;
      110839: inst = 32'hca00004;
      110840: inst = 32'h38632800;
      110841: inst = 32'h38842800;
      110842: inst = 32'h10a00001;
      110843: inst = 32'hca0b0ff;
      110844: inst = 32'h13e00001;
      110845: inst = 32'hfe0d96a;
      110846: inst = 32'h5be00000;
      110847: inst = 32'h8c50000;
      110848: inst = 32'h24612800;
      110849: inst = 32'h10a00000;
      110850: inst = 32'hca00018;
      110851: inst = 32'h24822800;
      110852: inst = 32'h10a00000;
      110853: inst = 32'hca00004;
      110854: inst = 32'h38632800;
      110855: inst = 32'h38842800;
      110856: inst = 32'h10a00001;
      110857: inst = 32'hca0b10d;
      110858: inst = 32'h13e00001;
      110859: inst = 32'hfe0d96a;
      110860: inst = 32'h5be00000;
      110861: inst = 32'h8c50000;
      110862: inst = 32'h24612800;
      110863: inst = 32'h10a00000;
      110864: inst = 32'hca00018;
      110865: inst = 32'h24822800;
      110866: inst = 32'h10a00000;
      110867: inst = 32'hca00004;
      110868: inst = 32'h38632800;
      110869: inst = 32'h38842800;
      110870: inst = 32'h10a00001;
      110871: inst = 32'hca0b11b;
      110872: inst = 32'h13e00001;
      110873: inst = 32'hfe0d96a;
      110874: inst = 32'h5be00000;
      110875: inst = 32'h8c50000;
      110876: inst = 32'h24612800;
      110877: inst = 32'h10a00000;
      110878: inst = 32'hca00018;
      110879: inst = 32'h24822800;
      110880: inst = 32'h10a00000;
      110881: inst = 32'hca00004;
      110882: inst = 32'h38632800;
      110883: inst = 32'h38842800;
      110884: inst = 32'h10a00001;
      110885: inst = 32'hca0b129;
      110886: inst = 32'h13e00001;
      110887: inst = 32'hfe0d96a;
      110888: inst = 32'h5be00000;
      110889: inst = 32'h8c50000;
      110890: inst = 32'h24612800;
      110891: inst = 32'h10a00000;
      110892: inst = 32'hca00018;
      110893: inst = 32'h24822800;
      110894: inst = 32'h10a00000;
      110895: inst = 32'hca00004;
      110896: inst = 32'h38632800;
      110897: inst = 32'h38842800;
      110898: inst = 32'h10a00001;
      110899: inst = 32'hca0b137;
      110900: inst = 32'h13e00001;
      110901: inst = 32'hfe0d96a;
      110902: inst = 32'h5be00000;
      110903: inst = 32'h8c50000;
      110904: inst = 32'h24612800;
      110905: inst = 32'h10a00000;
      110906: inst = 32'hca00018;
      110907: inst = 32'h24822800;
      110908: inst = 32'h10a00000;
      110909: inst = 32'hca00004;
      110910: inst = 32'h38632800;
      110911: inst = 32'h38842800;
      110912: inst = 32'h10a00001;
      110913: inst = 32'hca0b145;
      110914: inst = 32'h13e00001;
      110915: inst = 32'hfe0d96a;
      110916: inst = 32'h5be00000;
      110917: inst = 32'h8c50000;
      110918: inst = 32'h24612800;
      110919: inst = 32'h10a00000;
      110920: inst = 32'hca00018;
      110921: inst = 32'h24822800;
      110922: inst = 32'h10a00000;
      110923: inst = 32'hca00004;
      110924: inst = 32'h38632800;
      110925: inst = 32'h38842800;
      110926: inst = 32'h10a00001;
      110927: inst = 32'hca0b153;
      110928: inst = 32'h13e00001;
      110929: inst = 32'hfe0d96a;
      110930: inst = 32'h5be00000;
      110931: inst = 32'h8c50000;
      110932: inst = 32'h24612800;
      110933: inst = 32'h10a00000;
      110934: inst = 32'hca00018;
      110935: inst = 32'h24822800;
      110936: inst = 32'h10a00000;
      110937: inst = 32'hca00004;
      110938: inst = 32'h38632800;
      110939: inst = 32'h38842800;
      110940: inst = 32'h10a00001;
      110941: inst = 32'hca0b161;
      110942: inst = 32'h13e00001;
      110943: inst = 32'hfe0d96a;
      110944: inst = 32'h5be00000;
      110945: inst = 32'h8c50000;
      110946: inst = 32'h24612800;
      110947: inst = 32'h10a00000;
      110948: inst = 32'hca00018;
      110949: inst = 32'h24822800;
      110950: inst = 32'h10a00000;
      110951: inst = 32'hca00004;
      110952: inst = 32'h38632800;
      110953: inst = 32'h38842800;
      110954: inst = 32'h10a00001;
      110955: inst = 32'hca0b16f;
      110956: inst = 32'h13e00001;
      110957: inst = 32'hfe0d96a;
      110958: inst = 32'h5be00000;
      110959: inst = 32'h8c50000;
      110960: inst = 32'h24612800;
      110961: inst = 32'h10a00000;
      110962: inst = 32'hca00018;
      110963: inst = 32'h24822800;
      110964: inst = 32'h10a00000;
      110965: inst = 32'hca00004;
      110966: inst = 32'h38632800;
      110967: inst = 32'h38842800;
      110968: inst = 32'h10a00001;
      110969: inst = 32'hca0b17d;
      110970: inst = 32'h13e00001;
      110971: inst = 32'hfe0d96a;
      110972: inst = 32'h5be00000;
      110973: inst = 32'h8c50000;
      110974: inst = 32'h24612800;
      110975: inst = 32'h10a00000;
      110976: inst = 32'hca00018;
      110977: inst = 32'h24822800;
      110978: inst = 32'h10a00000;
      110979: inst = 32'hca00004;
      110980: inst = 32'h38632800;
      110981: inst = 32'h38842800;
      110982: inst = 32'h10a00001;
      110983: inst = 32'hca0b18b;
      110984: inst = 32'h13e00001;
      110985: inst = 32'hfe0d96a;
      110986: inst = 32'h5be00000;
      110987: inst = 32'h8c50000;
      110988: inst = 32'h24612800;
      110989: inst = 32'h10a00000;
      110990: inst = 32'hca00018;
      110991: inst = 32'h24822800;
      110992: inst = 32'h10a00000;
      110993: inst = 32'hca00004;
      110994: inst = 32'h38632800;
      110995: inst = 32'h38842800;
      110996: inst = 32'h10a00001;
      110997: inst = 32'hca0b199;
      110998: inst = 32'h13e00001;
      110999: inst = 32'hfe0d96a;
      111000: inst = 32'h5be00000;
      111001: inst = 32'h8c50000;
      111002: inst = 32'h24612800;
      111003: inst = 32'h10a00000;
      111004: inst = 32'hca00018;
      111005: inst = 32'h24822800;
      111006: inst = 32'h10a00000;
      111007: inst = 32'hca00004;
      111008: inst = 32'h38632800;
      111009: inst = 32'h38842800;
      111010: inst = 32'h10a00001;
      111011: inst = 32'hca0b1a7;
      111012: inst = 32'h13e00001;
      111013: inst = 32'hfe0d96a;
      111014: inst = 32'h5be00000;
      111015: inst = 32'h8c50000;
      111016: inst = 32'h24612800;
      111017: inst = 32'h10a00000;
      111018: inst = 32'hca00018;
      111019: inst = 32'h24822800;
      111020: inst = 32'h10a00000;
      111021: inst = 32'hca00004;
      111022: inst = 32'h38632800;
      111023: inst = 32'h38842800;
      111024: inst = 32'h10a00001;
      111025: inst = 32'hca0b1b5;
      111026: inst = 32'h13e00001;
      111027: inst = 32'hfe0d96a;
      111028: inst = 32'h5be00000;
      111029: inst = 32'h8c50000;
      111030: inst = 32'h24612800;
      111031: inst = 32'h10a00000;
      111032: inst = 32'hca00018;
      111033: inst = 32'h24822800;
      111034: inst = 32'h10a00000;
      111035: inst = 32'hca00004;
      111036: inst = 32'h38632800;
      111037: inst = 32'h38842800;
      111038: inst = 32'h10a00001;
      111039: inst = 32'hca0b1c3;
      111040: inst = 32'h13e00001;
      111041: inst = 32'hfe0d96a;
      111042: inst = 32'h5be00000;
      111043: inst = 32'h8c50000;
      111044: inst = 32'h24612800;
      111045: inst = 32'h10a00000;
      111046: inst = 32'hca00018;
      111047: inst = 32'h24822800;
      111048: inst = 32'h10a00000;
      111049: inst = 32'hca00004;
      111050: inst = 32'h38632800;
      111051: inst = 32'h38842800;
      111052: inst = 32'h10a00001;
      111053: inst = 32'hca0b1d1;
      111054: inst = 32'h13e00001;
      111055: inst = 32'hfe0d96a;
      111056: inst = 32'h5be00000;
      111057: inst = 32'h8c50000;
      111058: inst = 32'h24612800;
      111059: inst = 32'h10a00000;
      111060: inst = 32'hca00018;
      111061: inst = 32'h24822800;
      111062: inst = 32'h10a00000;
      111063: inst = 32'hca00004;
      111064: inst = 32'h38632800;
      111065: inst = 32'h38842800;
      111066: inst = 32'h10a00001;
      111067: inst = 32'hca0b1df;
      111068: inst = 32'h13e00001;
      111069: inst = 32'hfe0d96a;
      111070: inst = 32'h5be00000;
      111071: inst = 32'h8c50000;
      111072: inst = 32'h24612800;
      111073: inst = 32'h10a00000;
      111074: inst = 32'hca00018;
      111075: inst = 32'h24822800;
      111076: inst = 32'h10a00000;
      111077: inst = 32'hca00004;
      111078: inst = 32'h38632800;
      111079: inst = 32'h38842800;
      111080: inst = 32'h10a00001;
      111081: inst = 32'hca0b1ed;
      111082: inst = 32'h13e00001;
      111083: inst = 32'hfe0d96a;
      111084: inst = 32'h5be00000;
      111085: inst = 32'h8c50000;
      111086: inst = 32'h24612800;
      111087: inst = 32'h10a00000;
      111088: inst = 32'hca00018;
      111089: inst = 32'h24822800;
      111090: inst = 32'h10a00000;
      111091: inst = 32'hca00004;
      111092: inst = 32'h38632800;
      111093: inst = 32'h38842800;
      111094: inst = 32'h10a00001;
      111095: inst = 32'hca0b1fb;
      111096: inst = 32'h13e00001;
      111097: inst = 32'hfe0d96a;
      111098: inst = 32'h5be00000;
      111099: inst = 32'h8c50000;
      111100: inst = 32'h24612800;
      111101: inst = 32'h10a00000;
      111102: inst = 32'hca00018;
      111103: inst = 32'h24822800;
      111104: inst = 32'h10a00000;
      111105: inst = 32'hca00004;
      111106: inst = 32'h38632800;
      111107: inst = 32'h38842800;
      111108: inst = 32'h10a00001;
      111109: inst = 32'hca0b209;
      111110: inst = 32'h13e00001;
      111111: inst = 32'hfe0d96a;
      111112: inst = 32'h5be00000;
      111113: inst = 32'h8c50000;
      111114: inst = 32'h24612800;
      111115: inst = 32'h10a00000;
      111116: inst = 32'hca00018;
      111117: inst = 32'h24822800;
      111118: inst = 32'h10a00000;
      111119: inst = 32'hca00004;
      111120: inst = 32'h38632800;
      111121: inst = 32'h38842800;
      111122: inst = 32'h10a00001;
      111123: inst = 32'hca0b217;
      111124: inst = 32'h13e00001;
      111125: inst = 32'hfe0d96a;
      111126: inst = 32'h5be00000;
      111127: inst = 32'h8c50000;
      111128: inst = 32'h24612800;
      111129: inst = 32'h10a00000;
      111130: inst = 32'hca00018;
      111131: inst = 32'h24822800;
      111132: inst = 32'h10a00000;
      111133: inst = 32'hca00004;
      111134: inst = 32'h38632800;
      111135: inst = 32'h38842800;
      111136: inst = 32'h10a00001;
      111137: inst = 32'hca0b225;
      111138: inst = 32'h13e00001;
      111139: inst = 32'hfe0d96a;
      111140: inst = 32'h5be00000;
      111141: inst = 32'h8c50000;
      111142: inst = 32'h24612800;
      111143: inst = 32'h10a00000;
      111144: inst = 32'hca00018;
      111145: inst = 32'h24822800;
      111146: inst = 32'h10a00000;
      111147: inst = 32'hca00004;
      111148: inst = 32'h38632800;
      111149: inst = 32'h38842800;
      111150: inst = 32'h10a00001;
      111151: inst = 32'hca0b233;
      111152: inst = 32'h13e00001;
      111153: inst = 32'hfe0d96a;
      111154: inst = 32'h5be00000;
      111155: inst = 32'h8c50000;
      111156: inst = 32'h24612800;
      111157: inst = 32'h10a00000;
      111158: inst = 32'hca00018;
      111159: inst = 32'h24822800;
      111160: inst = 32'h10a00000;
      111161: inst = 32'hca00004;
      111162: inst = 32'h38632800;
      111163: inst = 32'h38842800;
      111164: inst = 32'h10a00001;
      111165: inst = 32'hca0b241;
      111166: inst = 32'h13e00001;
      111167: inst = 32'hfe0d96a;
      111168: inst = 32'h5be00000;
      111169: inst = 32'h8c50000;
      111170: inst = 32'h24612800;
      111171: inst = 32'h10a00000;
      111172: inst = 32'hca00018;
      111173: inst = 32'h24822800;
      111174: inst = 32'h10a00000;
      111175: inst = 32'hca00004;
      111176: inst = 32'h38632800;
      111177: inst = 32'h38842800;
      111178: inst = 32'h10a00001;
      111179: inst = 32'hca0b24f;
      111180: inst = 32'h13e00001;
      111181: inst = 32'hfe0d96a;
      111182: inst = 32'h5be00000;
      111183: inst = 32'h8c50000;
      111184: inst = 32'h24612800;
      111185: inst = 32'h10a00000;
      111186: inst = 32'hca00018;
      111187: inst = 32'h24822800;
      111188: inst = 32'h10a00000;
      111189: inst = 32'hca00004;
      111190: inst = 32'h38632800;
      111191: inst = 32'h38842800;
      111192: inst = 32'h10a00001;
      111193: inst = 32'hca0b25d;
      111194: inst = 32'h13e00001;
      111195: inst = 32'hfe0d96a;
      111196: inst = 32'h5be00000;
      111197: inst = 32'h8c50000;
      111198: inst = 32'h24612800;
      111199: inst = 32'h10a00000;
      111200: inst = 32'hca00018;
      111201: inst = 32'h24822800;
      111202: inst = 32'h10a00000;
      111203: inst = 32'hca00004;
      111204: inst = 32'h38632800;
      111205: inst = 32'h38842800;
      111206: inst = 32'h10a00001;
      111207: inst = 32'hca0b26b;
      111208: inst = 32'h13e00001;
      111209: inst = 32'hfe0d96a;
      111210: inst = 32'h5be00000;
      111211: inst = 32'h8c50000;
      111212: inst = 32'h24612800;
      111213: inst = 32'h10a00000;
      111214: inst = 32'hca00018;
      111215: inst = 32'h24822800;
      111216: inst = 32'h10a00000;
      111217: inst = 32'hca00004;
      111218: inst = 32'h38632800;
      111219: inst = 32'h38842800;
      111220: inst = 32'h10a00001;
      111221: inst = 32'hca0b279;
      111222: inst = 32'h13e00001;
      111223: inst = 32'hfe0d96a;
      111224: inst = 32'h5be00000;
      111225: inst = 32'h8c50000;
      111226: inst = 32'h24612800;
      111227: inst = 32'h10a00000;
      111228: inst = 32'hca00018;
      111229: inst = 32'h24822800;
      111230: inst = 32'h10a00000;
      111231: inst = 32'hca00004;
      111232: inst = 32'h38632800;
      111233: inst = 32'h38842800;
      111234: inst = 32'h10a00001;
      111235: inst = 32'hca0b287;
      111236: inst = 32'h13e00001;
      111237: inst = 32'hfe0d96a;
      111238: inst = 32'h5be00000;
      111239: inst = 32'h8c50000;
      111240: inst = 32'h24612800;
      111241: inst = 32'h10a00000;
      111242: inst = 32'hca00018;
      111243: inst = 32'h24822800;
      111244: inst = 32'h10a00000;
      111245: inst = 32'hca00004;
      111246: inst = 32'h38632800;
      111247: inst = 32'h38842800;
      111248: inst = 32'h10a00001;
      111249: inst = 32'hca0b295;
      111250: inst = 32'h13e00001;
      111251: inst = 32'hfe0d96a;
      111252: inst = 32'h5be00000;
      111253: inst = 32'h8c50000;
      111254: inst = 32'h24612800;
      111255: inst = 32'h10a00000;
      111256: inst = 32'hca00018;
      111257: inst = 32'h24822800;
      111258: inst = 32'h10a00000;
      111259: inst = 32'hca00004;
      111260: inst = 32'h38632800;
      111261: inst = 32'h38842800;
      111262: inst = 32'h10a00001;
      111263: inst = 32'hca0b2a3;
      111264: inst = 32'h13e00001;
      111265: inst = 32'hfe0d96a;
      111266: inst = 32'h5be00000;
      111267: inst = 32'h8c50000;
      111268: inst = 32'h24612800;
      111269: inst = 32'h10a00000;
      111270: inst = 32'hca00018;
      111271: inst = 32'h24822800;
      111272: inst = 32'h10a00000;
      111273: inst = 32'hca00004;
      111274: inst = 32'h38632800;
      111275: inst = 32'h38842800;
      111276: inst = 32'h10a00001;
      111277: inst = 32'hca0b2b1;
      111278: inst = 32'h13e00001;
      111279: inst = 32'hfe0d96a;
      111280: inst = 32'h5be00000;
      111281: inst = 32'h8c50000;
      111282: inst = 32'h24612800;
      111283: inst = 32'h10a00000;
      111284: inst = 32'hca00018;
      111285: inst = 32'h24822800;
      111286: inst = 32'h10a00000;
      111287: inst = 32'hca00004;
      111288: inst = 32'h38632800;
      111289: inst = 32'h38842800;
      111290: inst = 32'h10a00001;
      111291: inst = 32'hca0b2bf;
      111292: inst = 32'h13e00001;
      111293: inst = 32'hfe0d96a;
      111294: inst = 32'h5be00000;
      111295: inst = 32'h8c50000;
      111296: inst = 32'h24612800;
      111297: inst = 32'h10a00000;
      111298: inst = 32'hca00018;
      111299: inst = 32'h24822800;
      111300: inst = 32'h10a00000;
      111301: inst = 32'hca00004;
      111302: inst = 32'h38632800;
      111303: inst = 32'h38842800;
      111304: inst = 32'h10a00001;
      111305: inst = 32'hca0b2cd;
      111306: inst = 32'h13e00001;
      111307: inst = 32'hfe0d96a;
      111308: inst = 32'h5be00000;
      111309: inst = 32'h8c50000;
      111310: inst = 32'h24612800;
      111311: inst = 32'h10a00000;
      111312: inst = 32'hca00018;
      111313: inst = 32'h24822800;
      111314: inst = 32'h10a00000;
      111315: inst = 32'hca00004;
      111316: inst = 32'h38632800;
      111317: inst = 32'h38842800;
      111318: inst = 32'h10a00001;
      111319: inst = 32'hca0b2db;
      111320: inst = 32'h13e00001;
      111321: inst = 32'hfe0d96a;
      111322: inst = 32'h5be00000;
      111323: inst = 32'h8c50000;
      111324: inst = 32'h24612800;
      111325: inst = 32'h10a00000;
      111326: inst = 32'hca00018;
      111327: inst = 32'h24822800;
      111328: inst = 32'h10a00000;
      111329: inst = 32'hca00004;
      111330: inst = 32'h38632800;
      111331: inst = 32'h38842800;
      111332: inst = 32'h10a00001;
      111333: inst = 32'hca0b2e9;
      111334: inst = 32'h13e00001;
      111335: inst = 32'hfe0d96a;
      111336: inst = 32'h5be00000;
      111337: inst = 32'h8c50000;
      111338: inst = 32'h24612800;
      111339: inst = 32'h10a00000;
      111340: inst = 32'hca00018;
      111341: inst = 32'h24822800;
      111342: inst = 32'h10a00000;
      111343: inst = 32'hca00004;
      111344: inst = 32'h38632800;
      111345: inst = 32'h38842800;
      111346: inst = 32'h10a00001;
      111347: inst = 32'hca0b2f7;
      111348: inst = 32'h13e00001;
      111349: inst = 32'hfe0d96a;
      111350: inst = 32'h5be00000;
      111351: inst = 32'h8c50000;
      111352: inst = 32'h24612800;
      111353: inst = 32'h10a00000;
      111354: inst = 32'hca00018;
      111355: inst = 32'h24822800;
      111356: inst = 32'h10a00000;
      111357: inst = 32'hca00004;
      111358: inst = 32'h38632800;
      111359: inst = 32'h38842800;
      111360: inst = 32'h10a00001;
      111361: inst = 32'hca0b305;
      111362: inst = 32'h13e00001;
      111363: inst = 32'hfe0d96a;
      111364: inst = 32'h5be00000;
      111365: inst = 32'h8c50000;
      111366: inst = 32'h24612800;
      111367: inst = 32'h10a00000;
      111368: inst = 32'hca00018;
      111369: inst = 32'h24822800;
      111370: inst = 32'h10a00000;
      111371: inst = 32'hca00004;
      111372: inst = 32'h38632800;
      111373: inst = 32'h38842800;
      111374: inst = 32'h10a00001;
      111375: inst = 32'hca0b313;
      111376: inst = 32'h13e00001;
      111377: inst = 32'hfe0d96a;
      111378: inst = 32'h5be00000;
      111379: inst = 32'h8c50000;
      111380: inst = 32'h24612800;
      111381: inst = 32'h10a00000;
      111382: inst = 32'hca00018;
      111383: inst = 32'h24822800;
      111384: inst = 32'h10a00000;
      111385: inst = 32'hca00004;
      111386: inst = 32'h38632800;
      111387: inst = 32'h38842800;
      111388: inst = 32'h10a00001;
      111389: inst = 32'hca0b321;
      111390: inst = 32'h13e00001;
      111391: inst = 32'hfe0d96a;
      111392: inst = 32'h5be00000;
      111393: inst = 32'h8c50000;
      111394: inst = 32'h24612800;
      111395: inst = 32'h10a00000;
      111396: inst = 32'hca00018;
      111397: inst = 32'h24822800;
      111398: inst = 32'h10a00000;
      111399: inst = 32'hca00004;
      111400: inst = 32'h38632800;
      111401: inst = 32'h38842800;
      111402: inst = 32'h10a00001;
      111403: inst = 32'hca0b32f;
      111404: inst = 32'h13e00001;
      111405: inst = 32'hfe0d96a;
      111406: inst = 32'h5be00000;
      111407: inst = 32'h8c50000;
      111408: inst = 32'h24612800;
      111409: inst = 32'h10a00000;
      111410: inst = 32'hca00018;
      111411: inst = 32'h24822800;
      111412: inst = 32'h10a00000;
      111413: inst = 32'hca00004;
      111414: inst = 32'h38632800;
      111415: inst = 32'h38842800;
      111416: inst = 32'h10a00001;
      111417: inst = 32'hca0b33d;
      111418: inst = 32'h13e00001;
      111419: inst = 32'hfe0d96a;
      111420: inst = 32'h5be00000;
      111421: inst = 32'h8c50000;
      111422: inst = 32'h24612800;
      111423: inst = 32'h10a00000;
      111424: inst = 32'hca00018;
      111425: inst = 32'h24822800;
      111426: inst = 32'h10a00000;
      111427: inst = 32'hca00004;
      111428: inst = 32'h38632800;
      111429: inst = 32'h38842800;
      111430: inst = 32'h10a00001;
      111431: inst = 32'hca0b34b;
      111432: inst = 32'h13e00001;
      111433: inst = 32'hfe0d96a;
      111434: inst = 32'h5be00000;
      111435: inst = 32'h8c50000;
      111436: inst = 32'h24612800;
      111437: inst = 32'h10a00000;
      111438: inst = 32'hca00018;
      111439: inst = 32'h24822800;
      111440: inst = 32'h10a00000;
      111441: inst = 32'hca00004;
      111442: inst = 32'h38632800;
      111443: inst = 32'h38842800;
      111444: inst = 32'h10a00001;
      111445: inst = 32'hca0b359;
      111446: inst = 32'h13e00001;
      111447: inst = 32'hfe0d96a;
      111448: inst = 32'h5be00000;
      111449: inst = 32'h8c50000;
      111450: inst = 32'h24612800;
      111451: inst = 32'h10a00000;
      111452: inst = 32'hca00018;
      111453: inst = 32'h24822800;
      111454: inst = 32'h10a00000;
      111455: inst = 32'hca00004;
      111456: inst = 32'h38632800;
      111457: inst = 32'h38842800;
      111458: inst = 32'h10a00001;
      111459: inst = 32'hca0b367;
      111460: inst = 32'h13e00001;
      111461: inst = 32'hfe0d96a;
      111462: inst = 32'h5be00000;
      111463: inst = 32'h8c50000;
      111464: inst = 32'h24612800;
      111465: inst = 32'h10a00000;
      111466: inst = 32'hca00018;
      111467: inst = 32'h24822800;
      111468: inst = 32'h10a00000;
      111469: inst = 32'hca00004;
      111470: inst = 32'h38632800;
      111471: inst = 32'h38842800;
      111472: inst = 32'h10a00001;
      111473: inst = 32'hca0b375;
      111474: inst = 32'h13e00001;
      111475: inst = 32'hfe0d96a;
      111476: inst = 32'h5be00000;
      111477: inst = 32'h8c50000;
      111478: inst = 32'h24612800;
      111479: inst = 32'h10a00000;
      111480: inst = 32'hca00018;
      111481: inst = 32'h24822800;
      111482: inst = 32'h10a00000;
      111483: inst = 32'hca00004;
      111484: inst = 32'h38632800;
      111485: inst = 32'h38842800;
      111486: inst = 32'h10a00001;
      111487: inst = 32'hca0b383;
      111488: inst = 32'h13e00001;
      111489: inst = 32'hfe0d96a;
      111490: inst = 32'h5be00000;
      111491: inst = 32'h8c50000;
      111492: inst = 32'h24612800;
      111493: inst = 32'h10a00000;
      111494: inst = 32'hca00018;
      111495: inst = 32'h24822800;
      111496: inst = 32'h10a00000;
      111497: inst = 32'hca00004;
      111498: inst = 32'h38632800;
      111499: inst = 32'h38842800;
      111500: inst = 32'h10a00001;
      111501: inst = 32'hca0b391;
      111502: inst = 32'h13e00001;
      111503: inst = 32'hfe0d96a;
      111504: inst = 32'h5be00000;
      111505: inst = 32'h8c50000;
      111506: inst = 32'h24612800;
      111507: inst = 32'h10a00000;
      111508: inst = 32'hca00018;
      111509: inst = 32'h24822800;
      111510: inst = 32'h10a00000;
      111511: inst = 32'hca00004;
      111512: inst = 32'h38632800;
      111513: inst = 32'h38842800;
      111514: inst = 32'h10a00001;
      111515: inst = 32'hca0b39f;
      111516: inst = 32'h13e00001;
      111517: inst = 32'hfe0d96a;
      111518: inst = 32'h5be00000;
      111519: inst = 32'h8c50000;
      111520: inst = 32'h24612800;
      111521: inst = 32'h10a00000;
      111522: inst = 32'hca00018;
      111523: inst = 32'h24822800;
      111524: inst = 32'h10a00000;
      111525: inst = 32'hca00004;
      111526: inst = 32'h38632800;
      111527: inst = 32'h38842800;
      111528: inst = 32'h10a00001;
      111529: inst = 32'hca0b3ad;
      111530: inst = 32'h13e00001;
      111531: inst = 32'hfe0d96a;
      111532: inst = 32'h5be00000;
      111533: inst = 32'h8c50000;
      111534: inst = 32'h24612800;
      111535: inst = 32'h10a00000;
      111536: inst = 32'hca00018;
      111537: inst = 32'h24822800;
      111538: inst = 32'h10a00000;
      111539: inst = 32'hca00004;
      111540: inst = 32'h38632800;
      111541: inst = 32'h38842800;
      111542: inst = 32'h10a00001;
      111543: inst = 32'hca0b3bb;
      111544: inst = 32'h13e00001;
      111545: inst = 32'hfe0d96a;
      111546: inst = 32'h5be00000;
      111547: inst = 32'h8c50000;
      111548: inst = 32'h24612800;
      111549: inst = 32'h10a00000;
      111550: inst = 32'hca00018;
      111551: inst = 32'h24822800;
      111552: inst = 32'h10a00000;
      111553: inst = 32'hca00004;
      111554: inst = 32'h38632800;
      111555: inst = 32'h38842800;
      111556: inst = 32'h10a00001;
      111557: inst = 32'hca0b3c9;
      111558: inst = 32'h13e00001;
      111559: inst = 32'hfe0d96a;
      111560: inst = 32'h5be00000;
      111561: inst = 32'h8c50000;
      111562: inst = 32'h24612800;
      111563: inst = 32'h10a00000;
      111564: inst = 32'hca00018;
      111565: inst = 32'h24822800;
      111566: inst = 32'h10a00000;
      111567: inst = 32'hca00004;
      111568: inst = 32'h38632800;
      111569: inst = 32'h38842800;
      111570: inst = 32'h10a00001;
      111571: inst = 32'hca0b3d7;
      111572: inst = 32'h13e00001;
      111573: inst = 32'hfe0d96a;
      111574: inst = 32'h5be00000;
      111575: inst = 32'h8c50000;
      111576: inst = 32'h24612800;
      111577: inst = 32'h10a00000;
      111578: inst = 32'hca00018;
      111579: inst = 32'h24822800;
      111580: inst = 32'h10a00000;
      111581: inst = 32'hca00004;
      111582: inst = 32'h38632800;
      111583: inst = 32'h38842800;
      111584: inst = 32'h10a00001;
      111585: inst = 32'hca0b3e5;
      111586: inst = 32'h13e00001;
      111587: inst = 32'hfe0d96a;
      111588: inst = 32'h5be00000;
      111589: inst = 32'h8c50000;
      111590: inst = 32'h24612800;
      111591: inst = 32'h10a00000;
      111592: inst = 32'hca00018;
      111593: inst = 32'h24822800;
      111594: inst = 32'h10a00000;
      111595: inst = 32'hca00004;
      111596: inst = 32'h38632800;
      111597: inst = 32'h38842800;
      111598: inst = 32'h10a00001;
      111599: inst = 32'hca0b3f3;
      111600: inst = 32'h13e00001;
      111601: inst = 32'hfe0d96a;
      111602: inst = 32'h5be00000;
      111603: inst = 32'h8c50000;
      111604: inst = 32'h24612800;
      111605: inst = 32'h10a00000;
      111606: inst = 32'hca00018;
      111607: inst = 32'h24822800;
      111608: inst = 32'h10a00000;
      111609: inst = 32'hca00004;
      111610: inst = 32'h38632800;
      111611: inst = 32'h38842800;
      111612: inst = 32'h10a00001;
      111613: inst = 32'hca0b401;
      111614: inst = 32'h13e00001;
      111615: inst = 32'hfe0d96a;
      111616: inst = 32'h5be00000;
      111617: inst = 32'h8c50000;
      111618: inst = 32'h24612800;
      111619: inst = 32'h10a00000;
      111620: inst = 32'hca00018;
      111621: inst = 32'h24822800;
      111622: inst = 32'h10a00000;
      111623: inst = 32'hca00004;
      111624: inst = 32'h38632800;
      111625: inst = 32'h38842800;
      111626: inst = 32'h10a00001;
      111627: inst = 32'hca0b40f;
      111628: inst = 32'h13e00001;
      111629: inst = 32'hfe0d96a;
      111630: inst = 32'h5be00000;
      111631: inst = 32'h8c50000;
      111632: inst = 32'h24612800;
      111633: inst = 32'h10a00000;
      111634: inst = 32'hca00018;
      111635: inst = 32'h24822800;
      111636: inst = 32'h10a00000;
      111637: inst = 32'hca00004;
      111638: inst = 32'h38632800;
      111639: inst = 32'h38842800;
      111640: inst = 32'h10a00001;
      111641: inst = 32'hca0b41d;
      111642: inst = 32'h13e00001;
      111643: inst = 32'hfe0d96a;
      111644: inst = 32'h5be00000;
      111645: inst = 32'h8c50000;
      111646: inst = 32'h24612800;
      111647: inst = 32'h10a00000;
      111648: inst = 32'hca00018;
      111649: inst = 32'h24822800;
      111650: inst = 32'h10a00000;
      111651: inst = 32'hca00004;
      111652: inst = 32'h38632800;
      111653: inst = 32'h38842800;
      111654: inst = 32'h10a00001;
      111655: inst = 32'hca0b42b;
      111656: inst = 32'h13e00001;
      111657: inst = 32'hfe0d96a;
      111658: inst = 32'h5be00000;
      111659: inst = 32'h8c50000;
      111660: inst = 32'h24612800;
      111661: inst = 32'h10a00000;
      111662: inst = 32'hca00018;
      111663: inst = 32'h24822800;
      111664: inst = 32'h10a00000;
      111665: inst = 32'hca00004;
      111666: inst = 32'h38632800;
      111667: inst = 32'h38842800;
      111668: inst = 32'h10a00001;
      111669: inst = 32'hca0b439;
      111670: inst = 32'h13e00001;
      111671: inst = 32'hfe0d96a;
      111672: inst = 32'h5be00000;
      111673: inst = 32'h8c50000;
      111674: inst = 32'h24612800;
      111675: inst = 32'h10a00000;
      111676: inst = 32'hca00018;
      111677: inst = 32'h24822800;
      111678: inst = 32'h10a00000;
      111679: inst = 32'hca00004;
      111680: inst = 32'h38632800;
      111681: inst = 32'h38842800;
      111682: inst = 32'h10a00001;
      111683: inst = 32'hca0b447;
      111684: inst = 32'h13e00001;
      111685: inst = 32'hfe0d96a;
      111686: inst = 32'h5be00000;
      111687: inst = 32'h8c50000;
      111688: inst = 32'h24612800;
      111689: inst = 32'h10a00000;
      111690: inst = 32'hca00018;
      111691: inst = 32'h24822800;
      111692: inst = 32'h10a00000;
      111693: inst = 32'hca00004;
      111694: inst = 32'h38632800;
      111695: inst = 32'h38842800;
      111696: inst = 32'h10a00001;
      111697: inst = 32'hca0b455;
      111698: inst = 32'h13e00001;
      111699: inst = 32'hfe0d96a;
      111700: inst = 32'h5be00000;
      111701: inst = 32'h8c50000;
      111702: inst = 32'h24612800;
      111703: inst = 32'h10a00000;
      111704: inst = 32'hca00018;
      111705: inst = 32'h24822800;
      111706: inst = 32'h10a00000;
      111707: inst = 32'hca00004;
      111708: inst = 32'h38632800;
      111709: inst = 32'h38842800;
      111710: inst = 32'h10a00001;
      111711: inst = 32'hca0b463;
      111712: inst = 32'h13e00001;
      111713: inst = 32'hfe0d96a;
      111714: inst = 32'h5be00000;
      111715: inst = 32'h8c50000;
      111716: inst = 32'h24612800;
      111717: inst = 32'h10a00000;
      111718: inst = 32'hca00018;
      111719: inst = 32'h24822800;
      111720: inst = 32'h10a00000;
      111721: inst = 32'hca00004;
      111722: inst = 32'h38632800;
      111723: inst = 32'h38842800;
      111724: inst = 32'h10a00001;
      111725: inst = 32'hca0b471;
      111726: inst = 32'h13e00001;
      111727: inst = 32'hfe0d96a;
      111728: inst = 32'h5be00000;
      111729: inst = 32'h8c50000;
      111730: inst = 32'h24612800;
      111731: inst = 32'h10a00000;
      111732: inst = 32'hca00018;
      111733: inst = 32'h24822800;
      111734: inst = 32'h10a00000;
      111735: inst = 32'hca00004;
      111736: inst = 32'h38632800;
      111737: inst = 32'h38842800;
      111738: inst = 32'h10a00001;
      111739: inst = 32'hca0b47f;
      111740: inst = 32'h13e00001;
      111741: inst = 32'hfe0d96a;
      111742: inst = 32'h5be00000;
      111743: inst = 32'h8c50000;
      111744: inst = 32'h24612800;
      111745: inst = 32'h10a00000;
      111746: inst = 32'hca00018;
      111747: inst = 32'h24822800;
      111748: inst = 32'h10a00000;
      111749: inst = 32'hca00004;
      111750: inst = 32'h38632800;
      111751: inst = 32'h38842800;
      111752: inst = 32'h10a00001;
      111753: inst = 32'hca0b48d;
      111754: inst = 32'h13e00001;
      111755: inst = 32'hfe0d96a;
      111756: inst = 32'h5be00000;
      111757: inst = 32'h8c50000;
      111758: inst = 32'h24612800;
      111759: inst = 32'h10a00000;
      111760: inst = 32'hca00018;
      111761: inst = 32'h24822800;
      111762: inst = 32'h10a00000;
      111763: inst = 32'hca00004;
      111764: inst = 32'h38632800;
      111765: inst = 32'h38842800;
      111766: inst = 32'h10a00001;
      111767: inst = 32'hca0b49b;
      111768: inst = 32'h13e00001;
      111769: inst = 32'hfe0d96a;
      111770: inst = 32'h5be00000;
      111771: inst = 32'h8c50000;
      111772: inst = 32'h24612800;
      111773: inst = 32'h10a00000;
      111774: inst = 32'hca00018;
      111775: inst = 32'h24822800;
      111776: inst = 32'h10a00000;
      111777: inst = 32'hca00004;
      111778: inst = 32'h38632800;
      111779: inst = 32'h38842800;
      111780: inst = 32'h10a00001;
      111781: inst = 32'hca0b4a9;
      111782: inst = 32'h13e00001;
      111783: inst = 32'hfe0d96a;
      111784: inst = 32'h5be00000;
      111785: inst = 32'h8c50000;
      111786: inst = 32'h24612800;
      111787: inst = 32'h10a00000;
      111788: inst = 32'hca00019;
      111789: inst = 32'h24822800;
      111790: inst = 32'h10a00000;
      111791: inst = 32'hca00004;
      111792: inst = 32'h38632800;
      111793: inst = 32'h38842800;
      111794: inst = 32'h10a00001;
      111795: inst = 32'hca0b4b7;
      111796: inst = 32'h13e00001;
      111797: inst = 32'hfe0d96a;
      111798: inst = 32'h5be00000;
      111799: inst = 32'h8c50000;
      111800: inst = 32'h24612800;
      111801: inst = 32'h10a00000;
      111802: inst = 32'hca00019;
      111803: inst = 32'h24822800;
      111804: inst = 32'h10a00000;
      111805: inst = 32'hca00004;
      111806: inst = 32'h38632800;
      111807: inst = 32'h38842800;
      111808: inst = 32'h10a00001;
      111809: inst = 32'hca0b4c5;
      111810: inst = 32'h13e00001;
      111811: inst = 32'hfe0d96a;
      111812: inst = 32'h5be00000;
      111813: inst = 32'h8c50000;
      111814: inst = 32'h24612800;
      111815: inst = 32'h10a00000;
      111816: inst = 32'hca00019;
      111817: inst = 32'h24822800;
      111818: inst = 32'h10a00000;
      111819: inst = 32'hca00004;
      111820: inst = 32'h38632800;
      111821: inst = 32'h38842800;
      111822: inst = 32'h10a00001;
      111823: inst = 32'hca0b4d3;
      111824: inst = 32'h13e00001;
      111825: inst = 32'hfe0d96a;
      111826: inst = 32'h5be00000;
      111827: inst = 32'h8c50000;
      111828: inst = 32'h24612800;
      111829: inst = 32'h10a00000;
      111830: inst = 32'hca00019;
      111831: inst = 32'h24822800;
      111832: inst = 32'h10a00000;
      111833: inst = 32'hca00004;
      111834: inst = 32'h38632800;
      111835: inst = 32'h38842800;
      111836: inst = 32'h10a00001;
      111837: inst = 32'hca0b4e1;
      111838: inst = 32'h13e00001;
      111839: inst = 32'hfe0d96a;
      111840: inst = 32'h5be00000;
      111841: inst = 32'h8c50000;
      111842: inst = 32'h24612800;
      111843: inst = 32'h10a00000;
      111844: inst = 32'hca00019;
      111845: inst = 32'h24822800;
      111846: inst = 32'h10a00000;
      111847: inst = 32'hca00004;
      111848: inst = 32'h38632800;
      111849: inst = 32'h38842800;
      111850: inst = 32'h10a00001;
      111851: inst = 32'hca0b4ef;
      111852: inst = 32'h13e00001;
      111853: inst = 32'hfe0d96a;
      111854: inst = 32'h5be00000;
      111855: inst = 32'h8c50000;
      111856: inst = 32'h24612800;
      111857: inst = 32'h10a00000;
      111858: inst = 32'hca00019;
      111859: inst = 32'h24822800;
      111860: inst = 32'h10a00000;
      111861: inst = 32'hca00004;
      111862: inst = 32'h38632800;
      111863: inst = 32'h38842800;
      111864: inst = 32'h10a00001;
      111865: inst = 32'hca0b4fd;
      111866: inst = 32'h13e00001;
      111867: inst = 32'hfe0d96a;
      111868: inst = 32'h5be00000;
      111869: inst = 32'h8c50000;
      111870: inst = 32'h24612800;
      111871: inst = 32'h10a00000;
      111872: inst = 32'hca00019;
      111873: inst = 32'h24822800;
      111874: inst = 32'h10a00000;
      111875: inst = 32'hca00004;
      111876: inst = 32'h38632800;
      111877: inst = 32'h38842800;
      111878: inst = 32'h10a00001;
      111879: inst = 32'hca0b50b;
      111880: inst = 32'h13e00001;
      111881: inst = 32'hfe0d96a;
      111882: inst = 32'h5be00000;
      111883: inst = 32'h8c50000;
      111884: inst = 32'h24612800;
      111885: inst = 32'h10a00000;
      111886: inst = 32'hca00019;
      111887: inst = 32'h24822800;
      111888: inst = 32'h10a00000;
      111889: inst = 32'hca00004;
      111890: inst = 32'h38632800;
      111891: inst = 32'h38842800;
      111892: inst = 32'h10a00001;
      111893: inst = 32'hca0b519;
      111894: inst = 32'h13e00001;
      111895: inst = 32'hfe0d96a;
      111896: inst = 32'h5be00000;
      111897: inst = 32'h8c50000;
      111898: inst = 32'h24612800;
      111899: inst = 32'h10a00000;
      111900: inst = 32'hca00019;
      111901: inst = 32'h24822800;
      111902: inst = 32'h10a00000;
      111903: inst = 32'hca00004;
      111904: inst = 32'h38632800;
      111905: inst = 32'h38842800;
      111906: inst = 32'h10a00001;
      111907: inst = 32'hca0b527;
      111908: inst = 32'h13e00001;
      111909: inst = 32'hfe0d96a;
      111910: inst = 32'h5be00000;
      111911: inst = 32'h8c50000;
      111912: inst = 32'h24612800;
      111913: inst = 32'h10a00000;
      111914: inst = 32'hca00019;
      111915: inst = 32'h24822800;
      111916: inst = 32'h10a00000;
      111917: inst = 32'hca00004;
      111918: inst = 32'h38632800;
      111919: inst = 32'h38842800;
      111920: inst = 32'h10a00001;
      111921: inst = 32'hca0b535;
      111922: inst = 32'h13e00001;
      111923: inst = 32'hfe0d96a;
      111924: inst = 32'h5be00000;
      111925: inst = 32'h8c50000;
      111926: inst = 32'h24612800;
      111927: inst = 32'h10a00000;
      111928: inst = 32'hca00019;
      111929: inst = 32'h24822800;
      111930: inst = 32'h10a00000;
      111931: inst = 32'hca00004;
      111932: inst = 32'h38632800;
      111933: inst = 32'h38842800;
      111934: inst = 32'h10a00001;
      111935: inst = 32'hca0b543;
      111936: inst = 32'h13e00001;
      111937: inst = 32'hfe0d96a;
      111938: inst = 32'h5be00000;
      111939: inst = 32'h8c50000;
      111940: inst = 32'h24612800;
      111941: inst = 32'h10a00000;
      111942: inst = 32'hca00019;
      111943: inst = 32'h24822800;
      111944: inst = 32'h10a00000;
      111945: inst = 32'hca00004;
      111946: inst = 32'h38632800;
      111947: inst = 32'h38842800;
      111948: inst = 32'h10a00001;
      111949: inst = 32'hca0b551;
      111950: inst = 32'h13e00001;
      111951: inst = 32'hfe0d96a;
      111952: inst = 32'h5be00000;
      111953: inst = 32'h8c50000;
      111954: inst = 32'h24612800;
      111955: inst = 32'h10a00000;
      111956: inst = 32'hca00019;
      111957: inst = 32'h24822800;
      111958: inst = 32'h10a00000;
      111959: inst = 32'hca00004;
      111960: inst = 32'h38632800;
      111961: inst = 32'h38842800;
      111962: inst = 32'h10a00001;
      111963: inst = 32'hca0b55f;
      111964: inst = 32'h13e00001;
      111965: inst = 32'hfe0d96a;
      111966: inst = 32'h5be00000;
      111967: inst = 32'h8c50000;
      111968: inst = 32'h24612800;
      111969: inst = 32'h10a00000;
      111970: inst = 32'hca00019;
      111971: inst = 32'h24822800;
      111972: inst = 32'h10a00000;
      111973: inst = 32'hca00004;
      111974: inst = 32'h38632800;
      111975: inst = 32'h38842800;
      111976: inst = 32'h10a00001;
      111977: inst = 32'hca0b56d;
      111978: inst = 32'h13e00001;
      111979: inst = 32'hfe0d96a;
      111980: inst = 32'h5be00000;
      111981: inst = 32'h8c50000;
      111982: inst = 32'h24612800;
      111983: inst = 32'h10a00000;
      111984: inst = 32'hca00019;
      111985: inst = 32'h24822800;
      111986: inst = 32'h10a00000;
      111987: inst = 32'hca00004;
      111988: inst = 32'h38632800;
      111989: inst = 32'h38842800;
      111990: inst = 32'h10a00001;
      111991: inst = 32'hca0b57b;
      111992: inst = 32'h13e00001;
      111993: inst = 32'hfe0d96a;
      111994: inst = 32'h5be00000;
      111995: inst = 32'h8c50000;
      111996: inst = 32'h24612800;
      111997: inst = 32'h10a00000;
      111998: inst = 32'hca00019;
      111999: inst = 32'h24822800;
      112000: inst = 32'h10a00000;
      112001: inst = 32'hca00004;
      112002: inst = 32'h38632800;
      112003: inst = 32'h38842800;
      112004: inst = 32'h10a00001;
      112005: inst = 32'hca0b589;
      112006: inst = 32'h13e00001;
      112007: inst = 32'hfe0d96a;
      112008: inst = 32'h5be00000;
      112009: inst = 32'h8c50000;
      112010: inst = 32'h24612800;
      112011: inst = 32'h10a00000;
      112012: inst = 32'hca00019;
      112013: inst = 32'h24822800;
      112014: inst = 32'h10a00000;
      112015: inst = 32'hca00004;
      112016: inst = 32'h38632800;
      112017: inst = 32'h38842800;
      112018: inst = 32'h10a00001;
      112019: inst = 32'hca0b597;
      112020: inst = 32'h13e00001;
      112021: inst = 32'hfe0d96a;
      112022: inst = 32'h5be00000;
      112023: inst = 32'h8c50000;
      112024: inst = 32'h24612800;
      112025: inst = 32'h10a00000;
      112026: inst = 32'hca00019;
      112027: inst = 32'h24822800;
      112028: inst = 32'h10a00000;
      112029: inst = 32'hca00004;
      112030: inst = 32'h38632800;
      112031: inst = 32'h38842800;
      112032: inst = 32'h10a00001;
      112033: inst = 32'hca0b5a5;
      112034: inst = 32'h13e00001;
      112035: inst = 32'hfe0d96a;
      112036: inst = 32'h5be00000;
      112037: inst = 32'h8c50000;
      112038: inst = 32'h24612800;
      112039: inst = 32'h10a00000;
      112040: inst = 32'hca00019;
      112041: inst = 32'h24822800;
      112042: inst = 32'h10a00000;
      112043: inst = 32'hca00004;
      112044: inst = 32'h38632800;
      112045: inst = 32'h38842800;
      112046: inst = 32'h10a00001;
      112047: inst = 32'hca0b5b3;
      112048: inst = 32'h13e00001;
      112049: inst = 32'hfe0d96a;
      112050: inst = 32'h5be00000;
      112051: inst = 32'h8c50000;
      112052: inst = 32'h24612800;
      112053: inst = 32'h10a00000;
      112054: inst = 32'hca00019;
      112055: inst = 32'h24822800;
      112056: inst = 32'h10a00000;
      112057: inst = 32'hca00004;
      112058: inst = 32'h38632800;
      112059: inst = 32'h38842800;
      112060: inst = 32'h10a00001;
      112061: inst = 32'hca0b5c1;
      112062: inst = 32'h13e00001;
      112063: inst = 32'hfe0d96a;
      112064: inst = 32'h5be00000;
      112065: inst = 32'h8c50000;
      112066: inst = 32'h24612800;
      112067: inst = 32'h10a00000;
      112068: inst = 32'hca00019;
      112069: inst = 32'h24822800;
      112070: inst = 32'h10a00000;
      112071: inst = 32'hca00004;
      112072: inst = 32'h38632800;
      112073: inst = 32'h38842800;
      112074: inst = 32'h10a00001;
      112075: inst = 32'hca0b5cf;
      112076: inst = 32'h13e00001;
      112077: inst = 32'hfe0d96a;
      112078: inst = 32'h5be00000;
      112079: inst = 32'h8c50000;
      112080: inst = 32'h24612800;
      112081: inst = 32'h10a00000;
      112082: inst = 32'hca00019;
      112083: inst = 32'h24822800;
      112084: inst = 32'h10a00000;
      112085: inst = 32'hca00004;
      112086: inst = 32'h38632800;
      112087: inst = 32'h38842800;
      112088: inst = 32'h10a00001;
      112089: inst = 32'hca0b5dd;
      112090: inst = 32'h13e00001;
      112091: inst = 32'hfe0d96a;
      112092: inst = 32'h5be00000;
      112093: inst = 32'h8c50000;
      112094: inst = 32'h24612800;
      112095: inst = 32'h10a00000;
      112096: inst = 32'hca00019;
      112097: inst = 32'h24822800;
      112098: inst = 32'h10a00000;
      112099: inst = 32'hca00004;
      112100: inst = 32'h38632800;
      112101: inst = 32'h38842800;
      112102: inst = 32'h10a00001;
      112103: inst = 32'hca0b5eb;
      112104: inst = 32'h13e00001;
      112105: inst = 32'hfe0d96a;
      112106: inst = 32'h5be00000;
      112107: inst = 32'h8c50000;
      112108: inst = 32'h24612800;
      112109: inst = 32'h10a00000;
      112110: inst = 32'hca00019;
      112111: inst = 32'h24822800;
      112112: inst = 32'h10a00000;
      112113: inst = 32'hca00004;
      112114: inst = 32'h38632800;
      112115: inst = 32'h38842800;
      112116: inst = 32'h10a00001;
      112117: inst = 32'hca0b5f9;
      112118: inst = 32'h13e00001;
      112119: inst = 32'hfe0d96a;
      112120: inst = 32'h5be00000;
      112121: inst = 32'h8c50000;
      112122: inst = 32'h24612800;
      112123: inst = 32'h10a00000;
      112124: inst = 32'hca00019;
      112125: inst = 32'h24822800;
      112126: inst = 32'h10a00000;
      112127: inst = 32'hca00004;
      112128: inst = 32'h38632800;
      112129: inst = 32'h38842800;
      112130: inst = 32'h10a00001;
      112131: inst = 32'hca0b607;
      112132: inst = 32'h13e00001;
      112133: inst = 32'hfe0d96a;
      112134: inst = 32'h5be00000;
      112135: inst = 32'h8c50000;
      112136: inst = 32'h24612800;
      112137: inst = 32'h10a00000;
      112138: inst = 32'hca00019;
      112139: inst = 32'h24822800;
      112140: inst = 32'h10a00000;
      112141: inst = 32'hca00004;
      112142: inst = 32'h38632800;
      112143: inst = 32'h38842800;
      112144: inst = 32'h10a00001;
      112145: inst = 32'hca0b615;
      112146: inst = 32'h13e00001;
      112147: inst = 32'hfe0d96a;
      112148: inst = 32'h5be00000;
      112149: inst = 32'h8c50000;
      112150: inst = 32'h24612800;
      112151: inst = 32'h10a00000;
      112152: inst = 32'hca00019;
      112153: inst = 32'h24822800;
      112154: inst = 32'h10a00000;
      112155: inst = 32'hca00004;
      112156: inst = 32'h38632800;
      112157: inst = 32'h38842800;
      112158: inst = 32'h10a00001;
      112159: inst = 32'hca0b623;
      112160: inst = 32'h13e00001;
      112161: inst = 32'hfe0d96a;
      112162: inst = 32'h5be00000;
      112163: inst = 32'h8c50000;
      112164: inst = 32'h24612800;
      112165: inst = 32'h10a00000;
      112166: inst = 32'hca00019;
      112167: inst = 32'h24822800;
      112168: inst = 32'h10a00000;
      112169: inst = 32'hca00004;
      112170: inst = 32'h38632800;
      112171: inst = 32'h38842800;
      112172: inst = 32'h10a00001;
      112173: inst = 32'hca0b631;
      112174: inst = 32'h13e00001;
      112175: inst = 32'hfe0d96a;
      112176: inst = 32'h5be00000;
      112177: inst = 32'h8c50000;
      112178: inst = 32'h24612800;
      112179: inst = 32'h10a00000;
      112180: inst = 32'hca00019;
      112181: inst = 32'h24822800;
      112182: inst = 32'h10a00000;
      112183: inst = 32'hca00004;
      112184: inst = 32'h38632800;
      112185: inst = 32'h38842800;
      112186: inst = 32'h10a00001;
      112187: inst = 32'hca0b63f;
      112188: inst = 32'h13e00001;
      112189: inst = 32'hfe0d96a;
      112190: inst = 32'h5be00000;
      112191: inst = 32'h8c50000;
      112192: inst = 32'h24612800;
      112193: inst = 32'h10a00000;
      112194: inst = 32'hca00019;
      112195: inst = 32'h24822800;
      112196: inst = 32'h10a00000;
      112197: inst = 32'hca00004;
      112198: inst = 32'h38632800;
      112199: inst = 32'h38842800;
      112200: inst = 32'h10a00001;
      112201: inst = 32'hca0b64d;
      112202: inst = 32'h13e00001;
      112203: inst = 32'hfe0d96a;
      112204: inst = 32'h5be00000;
      112205: inst = 32'h8c50000;
      112206: inst = 32'h24612800;
      112207: inst = 32'h10a00000;
      112208: inst = 32'hca00019;
      112209: inst = 32'h24822800;
      112210: inst = 32'h10a00000;
      112211: inst = 32'hca00004;
      112212: inst = 32'h38632800;
      112213: inst = 32'h38842800;
      112214: inst = 32'h10a00001;
      112215: inst = 32'hca0b65b;
      112216: inst = 32'h13e00001;
      112217: inst = 32'hfe0d96a;
      112218: inst = 32'h5be00000;
      112219: inst = 32'h8c50000;
      112220: inst = 32'h24612800;
      112221: inst = 32'h10a00000;
      112222: inst = 32'hca00019;
      112223: inst = 32'h24822800;
      112224: inst = 32'h10a00000;
      112225: inst = 32'hca00004;
      112226: inst = 32'h38632800;
      112227: inst = 32'h38842800;
      112228: inst = 32'h10a00001;
      112229: inst = 32'hca0b669;
      112230: inst = 32'h13e00001;
      112231: inst = 32'hfe0d96a;
      112232: inst = 32'h5be00000;
      112233: inst = 32'h8c50000;
      112234: inst = 32'h24612800;
      112235: inst = 32'h10a00000;
      112236: inst = 32'hca00019;
      112237: inst = 32'h24822800;
      112238: inst = 32'h10a00000;
      112239: inst = 32'hca00004;
      112240: inst = 32'h38632800;
      112241: inst = 32'h38842800;
      112242: inst = 32'h10a00001;
      112243: inst = 32'hca0b677;
      112244: inst = 32'h13e00001;
      112245: inst = 32'hfe0d96a;
      112246: inst = 32'h5be00000;
      112247: inst = 32'h8c50000;
      112248: inst = 32'h24612800;
      112249: inst = 32'h10a00000;
      112250: inst = 32'hca00019;
      112251: inst = 32'h24822800;
      112252: inst = 32'h10a00000;
      112253: inst = 32'hca00004;
      112254: inst = 32'h38632800;
      112255: inst = 32'h38842800;
      112256: inst = 32'h10a00001;
      112257: inst = 32'hca0b685;
      112258: inst = 32'h13e00001;
      112259: inst = 32'hfe0d96a;
      112260: inst = 32'h5be00000;
      112261: inst = 32'h8c50000;
      112262: inst = 32'h24612800;
      112263: inst = 32'h10a00000;
      112264: inst = 32'hca00019;
      112265: inst = 32'h24822800;
      112266: inst = 32'h10a00000;
      112267: inst = 32'hca00004;
      112268: inst = 32'h38632800;
      112269: inst = 32'h38842800;
      112270: inst = 32'h10a00001;
      112271: inst = 32'hca0b693;
      112272: inst = 32'h13e00001;
      112273: inst = 32'hfe0d96a;
      112274: inst = 32'h5be00000;
      112275: inst = 32'h8c50000;
      112276: inst = 32'h24612800;
      112277: inst = 32'h10a00000;
      112278: inst = 32'hca00019;
      112279: inst = 32'h24822800;
      112280: inst = 32'h10a00000;
      112281: inst = 32'hca00004;
      112282: inst = 32'h38632800;
      112283: inst = 32'h38842800;
      112284: inst = 32'h10a00001;
      112285: inst = 32'hca0b6a1;
      112286: inst = 32'h13e00001;
      112287: inst = 32'hfe0d96a;
      112288: inst = 32'h5be00000;
      112289: inst = 32'h8c50000;
      112290: inst = 32'h24612800;
      112291: inst = 32'h10a00000;
      112292: inst = 32'hca00019;
      112293: inst = 32'h24822800;
      112294: inst = 32'h10a00000;
      112295: inst = 32'hca00004;
      112296: inst = 32'h38632800;
      112297: inst = 32'h38842800;
      112298: inst = 32'h10a00001;
      112299: inst = 32'hca0b6af;
      112300: inst = 32'h13e00001;
      112301: inst = 32'hfe0d96a;
      112302: inst = 32'h5be00000;
      112303: inst = 32'h8c50000;
      112304: inst = 32'h24612800;
      112305: inst = 32'h10a00000;
      112306: inst = 32'hca00019;
      112307: inst = 32'h24822800;
      112308: inst = 32'h10a00000;
      112309: inst = 32'hca00004;
      112310: inst = 32'h38632800;
      112311: inst = 32'h38842800;
      112312: inst = 32'h10a00001;
      112313: inst = 32'hca0b6bd;
      112314: inst = 32'h13e00001;
      112315: inst = 32'hfe0d96a;
      112316: inst = 32'h5be00000;
      112317: inst = 32'h8c50000;
      112318: inst = 32'h24612800;
      112319: inst = 32'h10a00000;
      112320: inst = 32'hca00019;
      112321: inst = 32'h24822800;
      112322: inst = 32'h10a00000;
      112323: inst = 32'hca00004;
      112324: inst = 32'h38632800;
      112325: inst = 32'h38842800;
      112326: inst = 32'h10a00001;
      112327: inst = 32'hca0b6cb;
      112328: inst = 32'h13e00001;
      112329: inst = 32'hfe0d96a;
      112330: inst = 32'h5be00000;
      112331: inst = 32'h8c50000;
      112332: inst = 32'h24612800;
      112333: inst = 32'h10a00000;
      112334: inst = 32'hca00019;
      112335: inst = 32'h24822800;
      112336: inst = 32'h10a00000;
      112337: inst = 32'hca00004;
      112338: inst = 32'h38632800;
      112339: inst = 32'h38842800;
      112340: inst = 32'h10a00001;
      112341: inst = 32'hca0b6d9;
      112342: inst = 32'h13e00001;
      112343: inst = 32'hfe0d96a;
      112344: inst = 32'h5be00000;
      112345: inst = 32'h8c50000;
      112346: inst = 32'h24612800;
      112347: inst = 32'h10a00000;
      112348: inst = 32'hca00019;
      112349: inst = 32'h24822800;
      112350: inst = 32'h10a00000;
      112351: inst = 32'hca00004;
      112352: inst = 32'h38632800;
      112353: inst = 32'h38842800;
      112354: inst = 32'h10a00001;
      112355: inst = 32'hca0b6e7;
      112356: inst = 32'h13e00001;
      112357: inst = 32'hfe0d96a;
      112358: inst = 32'h5be00000;
      112359: inst = 32'h8c50000;
      112360: inst = 32'h24612800;
      112361: inst = 32'h10a00000;
      112362: inst = 32'hca00019;
      112363: inst = 32'h24822800;
      112364: inst = 32'h10a00000;
      112365: inst = 32'hca00004;
      112366: inst = 32'h38632800;
      112367: inst = 32'h38842800;
      112368: inst = 32'h10a00001;
      112369: inst = 32'hca0b6f5;
      112370: inst = 32'h13e00001;
      112371: inst = 32'hfe0d96a;
      112372: inst = 32'h5be00000;
      112373: inst = 32'h8c50000;
      112374: inst = 32'h24612800;
      112375: inst = 32'h10a00000;
      112376: inst = 32'hca00019;
      112377: inst = 32'h24822800;
      112378: inst = 32'h10a00000;
      112379: inst = 32'hca00004;
      112380: inst = 32'h38632800;
      112381: inst = 32'h38842800;
      112382: inst = 32'h10a00001;
      112383: inst = 32'hca0b703;
      112384: inst = 32'h13e00001;
      112385: inst = 32'hfe0d96a;
      112386: inst = 32'h5be00000;
      112387: inst = 32'h8c50000;
      112388: inst = 32'h24612800;
      112389: inst = 32'h10a00000;
      112390: inst = 32'hca00019;
      112391: inst = 32'h24822800;
      112392: inst = 32'h10a00000;
      112393: inst = 32'hca00004;
      112394: inst = 32'h38632800;
      112395: inst = 32'h38842800;
      112396: inst = 32'h10a00001;
      112397: inst = 32'hca0b711;
      112398: inst = 32'h13e00001;
      112399: inst = 32'hfe0d96a;
      112400: inst = 32'h5be00000;
      112401: inst = 32'h8c50000;
      112402: inst = 32'h24612800;
      112403: inst = 32'h10a00000;
      112404: inst = 32'hca00019;
      112405: inst = 32'h24822800;
      112406: inst = 32'h10a00000;
      112407: inst = 32'hca00004;
      112408: inst = 32'h38632800;
      112409: inst = 32'h38842800;
      112410: inst = 32'h10a00001;
      112411: inst = 32'hca0b71f;
      112412: inst = 32'h13e00001;
      112413: inst = 32'hfe0d96a;
      112414: inst = 32'h5be00000;
      112415: inst = 32'h8c50000;
      112416: inst = 32'h24612800;
      112417: inst = 32'h10a00000;
      112418: inst = 32'hca00019;
      112419: inst = 32'h24822800;
      112420: inst = 32'h10a00000;
      112421: inst = 32'hca00004;
      112422: inst = 32'h38632800;
      112423: inst = 32'h38842800;
      112424: inst = 32'h10a00001;
      112425: inst = 32'hca0b72d;
      112426: inst = 32'h13e00001;
      112427: inst = 32'hfe0d96a;
      112428: inst = 32'h5be00000;
      112429: inst = 32'h8c50000;
      112430: inst = 32'h24612800;
      112431: inst = 32'h10a00000;
      112432: inst = 32'hca00019;
      112433: inst = 32'h24822800;
      112434: inst = 32'h10a00000;
      112435: inst = 32'hca00004;
      112436: inst = 32'h38632800;
      112437: inst = 32'h38842800;
      112438: inst = 32'h10a00001;
      112439: inst = 32'hca0b73b;
      112440: inst = 32'h13e00001;
      112441: inst = 32'hfe0d96a;
      112442: inst = 32'h5be00000;
      112443: inst = 32'h8c50000;
      112444: inst = 32'h24612800;
      112445: inst = 32'h10a00000;
      112446: inst = 32'hca00019;
      112447: inst = 32'h24822800;
      112448: inst = 32'h10a00000;
      112449: inst = 32'hca00004;
      112450: inst = 32'h38632800;
      112451: inst = 32'h38842800;
      112452: inst = 32'h10a00001;
      112453: inst = 32'hca0b749;
      112454: inst = 32'h13e00001;
      112455: inst = 32'hfe0d96a;
      112456: inst = 32'h5be00000;
      112457: inst = 32'h8c50000;
      112458: inst = 32'h24612800;
      112459: inst = 32'h10a00000;
      112460: inst = 32'hca00019;
      112461: inst = 32'h24822800;
      112462: inst = 32'h10a00000;
      112463: inst = 32'hca00004;
      112464: inst = 32'h38632800;
      112465: inst = 32'h38842800;
      112466: inst = 32'h10a00001;
      112467: inst = 32'hca0b757;
      112468: inst = 32'h13e00001;
      112469: inst = 32'hfe0d96a;
      112470: inst = 32'h5be00000;
      112471: inst = 32'h8c50000;
      112472: inst = 32'h24612800;
      112473: inst = 32'h10a00000;
      112474: inst = 32'hca00019;
      112475: inst = 32'h24822800;
      112476: inst = 32'h10a00000;
      112477: inst = 32'hca00004;
      112478: inst = 32'h38632800;
      112479: inst = 32'h38842800;
      112480: inst = 32'h10a00001;
      112481: inst = 32'hca0b765;
      112482: inst = 32'h13e00001;
      112483: inst = 32'hfe0d96a;
      112484: inst = 32'h5be00000;
      112485: inst = 32'h8c50000;
      112486: inst = 32'h24612800;
      112487: inst = 32'h10a00000;
      112488: inst = 32'hca00019;
      112489: inst = 32'h24822800;
      112490: inst = 32'h10a00000;
      112491: inst = 32'hca00004;
      112492: inst = 32'h38632800;
      112493: inst = 32'h38842800;
      112494: inst = 32'h10a00001;
      112495: inst = 32'hca0b773;
      112496: inst = 32'h13e00001;
      112497: inst = 32'hfe0d96a;
      112498: inst = 32'h5be00000;
      112499: inst = 32'h8c50000;
      112500: inst = 32'h24612800;
      112501: inst = 32'h10a00000;
      112502: inst = 32'hca00019;
      112503: inst = 32'h24822800;
      112504: inst = 32'h10a00000;
      112505: inst = 32'hca00004;
      112506: inst = 32'h38632800;
      112507: inst = 32'h38842800;
      112508: inst = 32'h10a00001;
      112509: inst = 32'hca0b781;
      112510: inst = 32'h13e00001;
      112511: inst = 32'hfe0d96a;
      112512: inst = 32'h5be00000;
      112513: inst = 32'h8c50000;
      112514: inst = 32'h24612800;
      112515: inst = 32'h10a00000;
      112516: inst = 32'hca00019;
      112517: inst = 32'h24822800;
      112518: inst = 32'h10a00000;
      112519: inst = 32'hca00004;
      112520: inst = 32'h38632800;
      112521: inst = 32'h38842800;
      112522: inst = 32'h10a00001;
      112523: inst = 32'hca0b78f;
      112524: inst = 32'h13e00001;
      112525: inst = 32'hfe0d96a;
      112526: inst = 32'h5be00000;
      112527: inst = 32'h8c50000;
      112528: inst = 32'h24612800;
      112529: inst = 32'h10a00000;
      112530: inst = 32'hca00019;
      112531: inst = 32'h24822800;
      112532: inst = 32'h10a00000;
      112533: inst = 32'hca00004;
      112534: inst = 32'h38632800;
      112535: inst = 32'h38842800;
      112536: inst = 32'h10a00001;
      112537: inst = 32'hca0b79d;
      112538: inst = 32'h13e00001;
      112539: inst = 32'hfe0d96a;
      112540: inst = 32'h5be00000;
      112541: inst = 32'h8c50000;
      112542: inst = 32'h24612800;
      112543: inst = 32'h10a00000;
      112544: inst = 32'hca00019;
      112545: inst = 32'h24822800;
      112546: inst = 32'h10a00000;
      112547: inst = 32'hca00004;
      112548: inst = 32'h38632800;
      112549: inst = 32'h38842800;
      112550: inst = 32'h10a00001;
      112551: inst = 32'hca0b7ab;
      112552: inst = 32'h13e00001;
      112553: inst = 32'hfe0d96a;
      112554: inst = 32'h5be00000;
      112555: inst = 32'h8c50000;
      112556: inst = 32'h24612800;
      112557: inst = 32'h10a00000;
      112558: inst = 32'hca00019;
      112559: inst = 32'h24822800;
      112560: inst = 32'h10a00000;
      112561: inst = 32'hca00004;
      112562: inst = 32'h38632800;
      112563: inst = 32'h38842800;
      112564: inst = 32'h10a00001;
      112565: inst = 32'hca0b7b9;
      112566: inst = 32'h13e00001;
      112567: inst = 32'hfe0d96a;
      112568: inst = 32'h5be00000;
      112569: inst = 32'h8c50000;
      112570: inst = 32'h24612800;
      112571: inst = 32'h10a00000;
      112572: inst = 32'hca00019;
      112573: inst = 32'h24822800;
      112574: inst = 32'h10a00000;
      112575: inst = 32'hca00004;
      112576: inst = 32'h38632800;
      112577: inst = 32'h38842800;
      112578: inst = 32'h10a00001;
      112579: inst = 32'hca0b7c7;
      112580: inst = 32'h13e00001;
      112581: inst = 32'hfe0d96a;
      112582: inst = 32'h5be00000;
      112583: inst = 32'h8c50000;
      112584: inst = 32'h24612800;
      112585: inst = 32'h10a00000;
      112586: inst = 32'hca00019;
      112587: inst = 32'h24822800;
      112588: inst = 32'h10a00000;
      112589: inst = 32'hca00004;
      112590: inst = 32'h38632800;
      112591: inst = 32'h38842800;
      112592: inst = 32'h10a00001;
      112593: inst = 32'hca0b7d5;
      112594: inst = 32'h13e00001;
      112595: inst = 32'hfe0d96a;
      112596: inst = 32'h5be00000;
      112597: inst = 32'h8c50000;
      112598: inst = 32'h24612800;
      112599: inst = 32'h10a00000;
      112600: inst = 32'hca00019;
      112601: inst = 32'h24822800;
      112602: inst = 32'h10a00000;
      112603: inst = 32'hca00004;
      112604: inst = 32'h38632800;
      112605: inst = 32'h38842800;
      112606: inst = 32'h10a00001;
      112607: inst = 32'hca0b7e3;
      112608: inst = 32'h13e00001;
      112609: inst = 32'hfe0d96a;
      112610: inst = 32'h5be00000;
      112611: inst = 32'h8c50000;
      112612: inst = 32'h24612800;
      112613: inst = 32'h10a00000;
      112614: inst = 32'hca00019;
      112615: inst = 32'h24822800;
      112616: inst = 32'h10a00000;
      112617: inst = 32'hca00004;
      112618: inst = 32'h38632800;
      112619: inst = 32'h38842800;
      112620: inst = 32'h10a00001;
      112621: inst = 32'hca0b7f1;
      112622: inst = 32'h13e00001;
      112623: inst = 32'hfe0d96a;
      112624: inst = 32'h5be00000;
      112625: inst = 32'h8c50000;
      112626: inst = 32'h24612800;
      112627: inst = 32'h10a00000;
      112628: inst = 32'hca00019;
      112629: inst = 32'h24822800;
      112630: inst = 32'h10a00000;
      112631: inst = 32'hca00004;
      112632: inst = 32'h38632800;
      112633: inst = 32'h38842800;
      112634: inst = 32'h10a00001;
      112635: inst = 32'hca0b7ff;
      112636: inst = 32'h13e00001;
      112637: inst = 32'hfe0d96a;
      112638: inst = 32'h5be00000;
      112639: inst = 32'h8c50000;
      112640: inst = 32'h24612800;
      112641: inst = 32'h10a00000;
      112642: inst = 32'hca00019;
      112643: inst = 32'h24822800;
      112644: inst = 32'h10a00000;
      112645: inst = 32'hca00004;
      112646: inst = 32'h38632800;
      112647: inst = 32'h38842800;
      112648: inst = 32'h10a00001;
      112649: inst = 32'hca0b80d;
      112650: inst = 32'h13e00001;
      112651: inst = 32'hfe0d96a;
      112652: inst = 32'h5be00000;
      112653: inst = 32'h8c50000;
      112654: inst = 32'h24612800;
      112655: inst = 32'h10a00000;
      112656: inst = 32'hca00019;
      112657: inst = 32'h24822800;
      112658: inst = 32'h10a00000;
      112659: inst = 32'hca00004;
      112660: inst = 32'h38632800;
      112661: inst = 32'h38842800;
      112662: inst = 32'h10a00001;
      112663: inst = 32'hca0b81b;
      112664: inst = 32'h13e00001;
      112665: inst = 32'hfe0d96a;
      112666: inst = 32'h5be00000;
      112667: inst = 32'h8c50000;
      112668: inst = 32'h24612800;
      112669: inst = 32'h10a00000;
      112670: inst = 32'hca00019;
      112671: inst = 32'h24822800;
      112672: inst = 32'h10a00000;
      112673: inst = 32'hca00004;
      112674: inst = 32'h38632800;
      112675: inst = 32'h38842800;
      112676: inst = 32'h10a00001;
      112677: inst = 32'hca0b829;
      112678: inst = 32'h13e00001;
      112679: inst = 32'hfe0d96a;
      112680: inst = 32'h5be00000;
      112681: inst = 32'h8c50000;
      112682: inst = 32'h24612800;
      112683: inst = 32'h10a00000;
      112684: inst = 32'hca00019;
      112685: inst = 32'h24822800;
      112686: inst = 32'h10a00000;
      112687: inst = 32'hca00004;
      112688: inst = 32'h38632800;
      112689: inst = 32'h38842800;
      112690: inst = 32'h10a00001;
      112691: inst = 32'hca0b837;
      112692: inst = 32'h13e00001;
      112693: inst = 32'hfe0d96a;
      112694: inst = 32'h5be00000;
      112695: inst = 32'h8c50000;
      112696: inst = 32'h24612800;
      112697: inst = 32'h10a00000;
      112698: inst = 32'hca00019;
      112699: inst = 32'h24822800;
      112700: inst = 32'h10a00000;
      112701: inst = 32'hca00004;
      112702: inst = 32'h38632800;
      112703: inst = 32'h38842800;
      112704: inst = 32'h10a00001;
      112705: inst = 32'hca0b845;
      112706: inst = 32'h13e00001;
      112707: inst = 32'hfe0d96a;
      112708: inst = 32'h5be00000;
      112709: inst = 32'h8c50000;
      112710: inst = 32'h24612800;
      112711: inst = 32'h10a00000;
      112712: inst = 32'hca00019;
      112713: inst = 32'h24822800;
      112714: inst = 32'h10a00000;
      112715: inst = 32'hca00004;
      112716: inst = 32'h38632800;
      112717: inst = 32'h38842800;
      112718: inst = 32'h10a00001;
      112719: inst = 32'hca0b853;
      112720: inst = 32'h13e00001;
      112721: inst = 32'hfe0d96a;
      112722: inst = 32'h5be00000;
      112723: inst = 32'h8c50000;
      112724: inst = 32'h24612800;
      112725: inst = 32'h10a00000;
      112726: inst = 32'hca00019;
      112727: inst = 32'h24822800;
      112728: inst = 32'h10a00000;
      112729: inst = 32'hca00004;
      112730: inst = 32'h38632800;
      112731: inst = 32'h38842800;
      112732: inst = 32'h10a00001;
      112733: inst = 32'hca0b861;
      112734: inst = 32'h13e00001;
      112735: inst = 32'hfe0d96a;
      112736: inst = 32'h5be00000;
      112737: inst = 32'h8c50000;
      112738: inst = 32'h24612800;
      112739: inst = 32'h10a00000;
      112740: inst = 32'hca00019;
      112741: inst = 32'h24822800;
      112742: inst = 32'h10a00000;
      112743: inst = 32'hca00004;
      112744: inst = 32'h38632800;
      112745: inst = 32'h38842800;
      112746: inst = 32'h10a00001;
      112747: inst = 32'hca0b86f;
      112748: inst = 32'h13e00001;
      112749: inst = 32'hfe0d96a;
      112750: inst = 32'h5be00000;
      112751: inst = 32'h8c50000;
      112752: inst = 32'h24612800;
      112753: inst = 32'h10a00000;
      112754: inst = 32'hca00019;
      112755: inst = 32'h24822800;
      112756: inst = 32'h10a00000;
      112757: inst = 32'hca00004;
      112758: inst = 32'h38632800;
      112759: inst = 32'h38842800;
      112760: inst = 32'h10a00001;
      112761: inst = 32'hca0b87d;
      112762: inst = 32'h13e00001;
      112763: inst = 32'hfe0d96a;
      112764: inst = 32'h5be00000;
      112765: inst = 32'h8c50000;
      112766: inst = 32'h24612800;
      112767: inst = 32'h10a00000;
      112768: inst = 32'hca00019;
      112769: inst = 32'h24822800;
      112770: inst = 32'h10a00000;
      112771: inst = 32'hca00004;
      112772: inst = 32'h38632800;
      112773: inst = 32'h38842800;
      112774: inst = 32'h10a00001;
      112775: inst = 32'hca0b88b;
      112776: inst = 32'h13e00001;
      112777: inst = 32'hfe0d96a;
      112778: inst = 32'h5be00000;
      112779: inst = 32'h8c50000;
      112780: inst = 32'h24612800;
      112781: inst = 32'h10a00000;
      112782: inst = 32'hca00019;
      112783: inst = 32'h24822800;
      112784: inst = 32'h10a00000;
      112785: inst = 32'hca00004;
      112786: inst = 32'h38632800;
      112787: inst = 32'h38842800;
      112788: inst = 32'h10a00001;
      112789: inst = 32'hca0b899;
      112790: inst = 32'h13e00001;
      112791: inst = 32'hfe0d96a;
      112792: inst = 32'h5be00000;
      112793: inst = 32'h8c50000;
      112794: inst = 32'h24612800;
      112795: inst = 32'h10a00000;
      112796: inst = 32'hca00019;
      112797: inst = 32'h24822800;
      112798: inst = 32'h10a00000;
      112799: inst = 32'hca00004;
      112800: inst = 32'h38632800;
      112801: inst = 32'h38842800;
      112802: inst = 32'h10a00001;
      112803: inst = 32'hca0b8a7;
      112804: inst = 32'h13e00001;
      112805: inst = 32'hfe0d96a;
      112806: inst = 32'h5be00000;
      112807: inst = 32'h8c50000;
      112808: inst = 32'h24612800;
      112809: inst = 32'h10a00000;
      112810: inst = 32'hca00019;
      112811: inst = 32'h24822800;
      112812: inst = 32'h10a00000;
      112813: inst = 32'hca00004;
      112814: inst = 32'h38632800;
      112815: inst = 32'h38842800;
      112816: inst = 32'h10a00001;
      112817: inst = 32'hca0b8b5;
      112818: inst = 32'h13e00001;
      112819: inst = 32'hfe0d96a;
      112820: inst = 32'h5be00000;
      112821: inst = 32'h8c50000;
      112822: inst = 32'h24612800;
      112823: inst = 32'h10a00000;
      112824: inst = 32'hca00019;
      112825: inst = 32'h24822800;
      112826: inst = 32'h10a00000;
      112827: inst = 32'hca00004;
      112828: inst = 32'h38632800;
      112829: inst = 32'h38842800;
      112830: inst = 32'h10a00001;
      112831: inst = 32'hca0b8c3;
      112832: inst = 32'h13e00001;
      112833: inst = 32'hfe0d96a;
      112834: inst = 32'h5be00000;
      112835: inst = 32'h8c50000;
      112836: inst = 32'h24612800;
      112837: inst = 32'h10a00000;
      112838: inst = 32'hca00019;
      112839: inst = 32'h24822800;
      112840: inst = 32'h10a00000;
      112841: inst = 32'hca00004;
      112842: inst = 32'h38632800;
      112843: inst = 32'h38842800;
      112844: inst = 32'h10a00001;
      112845: inst = 32'hca0b8d1;
      112846: inst = 32'h13e00001;
      112847: inst = 32'hfe0d96a;
      112848: inst = 32'h5be00000;
      112849: inst = 32'h8c50000;
      112850: inst = 32'h24612800;
      112851: inst = 32'h10a00000;
      112852: inst = 32'hca00019;
      112853: inst = 32'h24822800;
      112854: inst = 32'h10a00000;
      112855: inst = 32'hca00004;
      112856: inst = 32'h38632800;
      112857: inst = 32'h38842800;
      112858: inst = 32'h10a00001;
      112859: inst = 32'hca0b8df;
      112860: inst = 32'h13e00001;
      112861: inst = 32'hfe0d96a;
      112862: inst = 32'h5be00000;
      112863: inst = 32'h8c50000;
      112864: inst = 32'h24612800;
      112865: inst = 32'h10a00000;
      112866: inst = 32'hca00019;
      112867: inst = 32'h24822800;
      112868: inst = 32'h10a00000;
      112869: inst = 32'hca00004;
      112870: inst = 32'h38632800;
      112871: inst = 32'h38842800;
      112872: inst = 32'h10a00001;
      112873: inst = 32'hca0b8ed;
      112874: inst = 32'h13e00001;
      112875: inst = 32'hfe0d96a;
      112876: inst = 32'h5be00000;
      112877: inst = 32'h8c50000;
      112878: inst = 32'h24612800;
      112879: inst = 32'h10a00000;
      112880: inst = 32'hca00019;
      112881: inst = 32'h24822800;
      112882: inst = 32'h10a00000;
      112883: inst = 32'hca00004;
      112884: inst = 32'h38632800;
      112885: inst = 32'h38842800;
      112886: inst = 32'h10a00001;
      112887: inst = 32'hca0b8fb;
      112888: inst = 32'h13e00001;
      112889: inst = 32'hfe0d96a;
      112890: inst = 32'h5be00000;
      112891: inst = 32'h8c50000;
      112892: inst = 32'h24612800;
      112893: inst = 32'h10a00000;
      112894: inst = 32'hca00019;
      112895: inst = 32'h24822800;
      112896: inst = 32'h10a00000;
      112897: inst = 32'hca00004;
      112898: inst = 32'h38632800;
      112899: inst = 32'h38842800;
      112900: inst = 32'h10a00001;
      112901: inst = 32'hca0b909;
      112902: inst = 32'h13e00001;
      112903: inst = 32'hfe0d96a;
      112904: inst = 32'h5be00000;
      112905: inst = 32'h8c50000;
      112906: inst = 32'h24612800;
      112907: inst = 32'h10a00000;
      112908: inst = 32'hca00019;
      112909: inst = 32'h24822800;
      112910: inst = 32'h10a00000;
      112911: inst = 32'hca00004;
      112912: inst = 32'h38632800;
      112913: inst = 32'h38842800;
      112914: inst = 32'h10a00001;
      112915: inst = 32'hca0b917;
      112916: inst = 32'h13e00001;
      112917: inst = 32'hfe0d96a;
      112918: inst = 32'h5be00000;
      112919: inst = 32'h8c50000;
      112920: inst = 32'h24612800;
      112921: inst = 32'h10a00000;
      112922: inst = 32'hca00019;
      112923: inst = 32'h24822800;
      112924: inst = 32'h10a00000;
      112925: inst = 32'hca00004;
      112926: inst = 32'h38632800;
      112927: inst = 32'h38842800;
      112928: inst = 32'h10a00001;
      112929: inst = 32'hca0b925;
      112930: inst = 32'h13e00001;
      112931: inst = 32'hfe0d96a;
      112932: inst = 32'h5be00000;
      112933: inst = 32'h8c50000;
      112934: inst = 32'h24612800;
      112935: inst = 32'h10a00000;
      112936: inst = 32'hca00019;
      112937: inst = 32'h24822800;
      112938: inst = 32'h10a00000;
      112939: inst = 32'hca00004;
      112940: inst = 32'h38632800;
      112941: inst = 32'h38842800;
      112942: inst = 32'h10a00001;
      112943: inst = 32'hca0b933;
      112944: inst = 32'h13e00001;
      112945: inst = 32'hfe0d96a;
      112946: inst = 32'h5be00000;
      112947: inst = 32'h8c50000;
      112948: inst = 32'h24612800;
      112949: inst = 32'h10a00000;
      112950: inst = 32'hca00019;
      112951: inst = 32'h24822800;
      112952: inst = 32'h10a00000;
      112953: inst = 32'hca00004;
      112954: inst = 32'h38632800;
      112955: inst = 32'h38842800;
      112956: inst = 32'h10a00001;
      112957: inst = 32'hca0b941;
      112958: inst = 32'h13e00001;
      112959: inst = 32'hfe0d96a;
      112960: inst = 32'h5be00000;
      112961: inst = 32'h8c50000;
      112962: inst = 32'h24612800;
      112963: inst = 32'h10a00000;
      112964: inst = 32'hca00019;
      112965: inst = 32'h24822800;
      112966: inst = 32'h10a00000;
      112967: inst = 32'hca00004;
      112968: inst = 32'h38632800;
      112969: inst = 32'h38842800;
      112970: inst = 32'h10a00001;
      112971: inst = 32'hca0b94f;
      112972: inst = 32'h13e00001;
      112973: inst = 32'hfe0d96a;
      112974: inst = 32'h5be00000;
      112975: inst = 32'h8c50000;
      112976: inst = 32'h24612800;
      112977: inst = 32'h10a00000;
      112978: inst = 32'hca00019;
      112979: inst = 32'h24822800;
      112980: inst = 32'h10a00000;
      112981: inst = 32'hca00004;
      112982: inst = 32'h38632800;
      112983: inst = 32'h38842800;
      112984: inst = 32'h10a00001;
      112985: inst = 32'hca0b95d;
      112986: inst = 32'h13e00001;
      112987: inst = 32'hfe0d96a;
      112988: inst = 32'h5be00000;
      112989: inst = 32'h8c50000;
      112990: inst = 32'h24612800;
      112991: inst = 32'h10a00000;
      112992: inst = 32'hca00019;
      112993: inst = 32'h24822800;
      112994: inst = 32'h10a00000;
      112995: inst = 32'hca00004;
      112996: inst = 32'h38632800;
      112997: inst = 32'h38842800;
      112998: inst = 32'h10a00001;
      112999: inst = 32'hca0b96b;
      113000: inst = 32'h13e00001;
      113001: inst = 32'hfe0d96a;
      113002: inst = 32'h5be00000;
      113003: inst = 32'h8c50000;
      113004: inst = 32'h24612800;
      113005: inst = 32'h10a00000;
      113006: inst = 32'hca00019;
      113007: inst = 32'h24822800;
      113008: inst = 32'h10a00000;
      113009: inst = 32'hca00004;
      113010: inst = 32'h38632800;
      113011: inst = 32'h38842800;
      113012: inst = 32'h10a00001;
      113013: inst = 32'hca0b979;
      113014: inst = 32'h13e00001;
      113015: inst = 32'hfe0d96a;
      113016: inst = 32'h5be00000;
      113017: inst = 32'h8c50000;
      113018: inst = 32'h24612800;
      113019: inst = 32'h10a00000;
      113020: inst = 32'hca00019;
      113021: inst = 32'h24822800;
      113022: inst = 32'h10a00000;
      113023: inst = 32'hca00004;
      113024: inst = 32'h38632800;
      113025: inst = 32'h38842800;
      113026: inst = 32'h10a00001;
      113027: inst = 32'hca0b987;
      113028: inst = 32'h13e00001;
      113029: inst = 32'hfe0d96a;
      113030: inst = 32'h5be00000;
      113031: inst = 32'h8c50000;
      113032: inst = 32'h24612800;
      113033: inst = 32'h10a00000;
      113034: inst = 32'hca00019;
      113035: inst = 32'h24822800;
      113036: inst = 32'h10a00000;
      113037: inst = 32'hca00004;
      113038: inst = 32'h38632800;
      113039: inst = 32'h38842800;
      113040: inst = 32'h10a00001;
      113041: inst = 32'hca0b995;
      113042: inst = 32'h13e00001;
      113043: inst = 32'hfe0d96a;
      113044: inst = 32'h5be00000;
      113045: inst = 32'h8c50000;
      113046: inst = 32'h24612800;
      113047: inst = 32'h10a00000;
      113048: inst = 32'hca00019;
      113049: inst = 32'h24822800;
      113050: inst = 32'h10a00000;
      113051: inst = 32'hca00004;
      113052: inst = 32'h38632800;
      113053: inst = 32'h38842800;
      113054: inst = 32'h10a00001;
      113055: inst = 32'hca0b9a3;
      113056: inst = 32'h13e00001;
      113057: inst = 32'hfe0d96a;
      113058: inst = 32'h5be00000;
      113059: inst = 32'h8c50000;
      113060: inst = 32'h24612800;
      113061: inst = 32'h10a00000;
      113062: inst = 32'hca00019;
      113063: inst = 32'h24822800;
      113064: inst = 32'h10a00000;
      113065: inst = 32'hca00004;
      113066: inst = 32'h38632800;
      113067: inst = 32'h38842800;
      113068: inst = 32'h10a00001;
      113069: inst = 32'hca0b9b1;
      113070: inst = 32'h13e00001;
      113071: inst = 32'hfe0d96a;
      113072: inst = 32'h5be00000;
      113073: inst = 32'h8c50000;
      113074: inst = 32'h24612800;
      113075: inst = 32'h10a00000;
      113076: inst = 32'hca00019;
      113077: inst = 32'h24822800;
      113078: inst = 32'h10a00000;
      113079: inst = 32'hca00004;
      113080: inst = 32'h38632800;
      113081: inst = 32'h38842800;
      113082: inst = 32'h10a00001;
      113083: inst = 32'hca0b9bf;
      113084: inst = 32'h13e00001;
      113085: inst = 32'hfe0d96a;
      113086: inst = 32'h5be00000;
      113087: inst = 32'h8c50000;
      113088: inst = 32'h24612800;
      113089: inst = 32'h10a00000;
      113090: inst = 32'hca00019;
      113091: inst = 32'h24822800;
      113092: inst = 32'h10a00000;
      113093: inst = 32'hca00004;
      113094: inst = 32'h38632800;
      113095: inst = 32'h38842800;
      113096: inst = 32'h10a00001;
      113097: inst = 32'hca0b9cd;
      113098: inst = 32'h13e00001;
      113099: inst = 32'hfe0d96a;
      113100: inst = 32'h5be00000;
      113101: inst = 32'h8c50000;
      113102: inst = 32'h24612800;
      113103: inst = 32'h10a00000;
      113104: inst = 32'hca00019;
      113105: inst = 32'h24822800;
      113106: inst = 32'h10a00000;
      113107: inst = 32'hca00004;
      113108: inst = 32'h38632800;
      113109: inst = 32'h38842800;
      113110: inst = 32'h10a00001;
      113111: inst = 32'hca0b9db;
      113112: inst = 32'h13e00001;
      113113: inst = 32'hfe0d96a;
      113114: inst = 32'h5be00000;
      113115: inst = 32'h8c50000;
      113116: inst = 32'h24612800;
      113117: inst = 32'h10a00000;
      113118: inst = 32'hca00019;
      113119: inst = 32'h24822800;
      113120: inst = 32'h10a00000;
      113121: inst = 32'hca00004;
      113122: inst = 32'h38632800;
      113123: inst = 32'h38842800;
      113124: inst = 32'h10a00001;
      113125: inst = 32'hca0b9e9;
      113126: inst = 32'h13e00001;
      113127: inst = 32'hfe0d96a;
      113128: inst = 32'h5be00000;
      113129: inst = 32'h8c50000;
      113130: inst = 32'h24612800;
      113131: inst = 32'h10a00000;
      113132: inst = 32'hca0001a;
      113133: inst = 32'h24822800;
      113134: inst = 32'h10a00000;
      113135: inst = 32'hca00004;
      113136: inst = 32'h38632800;
      113137: inst = 32'h38842800;
      113138: inst = 32'h10a00001;
      113139: inst = 32'hca0b9f7;
      113140: inst = 32'h13e00001;
      113141: inst = 32'hfe0d96a;
      113142: inst = 32'h5be00000;
      113143: inst = 32'h8c50000;
      113144: inst = 32'h24612800;
      113145: inst = 32'h10a00000;
      113146: inst = 32'hca0001a;
      113147: inst = 32'h24822800;
      113148: inst = 32'h10a00000;
      113149: inst = 32'hca00004;
      113150: inst = 32'h38632800;
      113151: inst = 32'h38842800;
      113152: inst = 32'h10a00001;
      113153: inst = 32'hca0ba05;
      113154: inst = 32'h13e00001;
      113155: inst = 32'hfe0d96a;
      113156: inst = 32'h5be00000;
      113157: inst = 32'h8c50000;
      113158: inst = 32'h24612800;
      113159: inst = 32'h10a00000;
      113160: inst = 32'hca0001a;
      113161: inst = 32'h24822800;
      113162: inst = 32'h10a00000;
      113163: inst = 32'hca00004;
      113164: inst = 32'h38632800;
      113165: inst = 32'h38842800;
      113166: inst = 32'h10a00001;
      113167: inst = 32'hca0ba13;
      113168: inst = 32'h13e00001;
      113169: inst = 32'hfe0d96a;
      113170: inst = 32'h5be00000;
      113171: inst = 32'h8c50000;
      113172: inst = 32'h24612800;
      113173: inst = 32'h10a00000;
      113174: inst = 32'hca0001a;
      113175: inst = 32'h24822800;
      113176: inst = 32'h10a00000;
      113177: inst = 32'hca00004;
      113178: inst = 32'h38632800;
      113179: inst = 32'h38842800;
      113180: inst = 32'h10a00001;
      113181: inst = 32'hca0ba21;
      113182: inst = 32'h13e00001;
      113183: inst = 32'hfe0d96a;
      113184: inst = 32'h5be00000;
      113185: inst = 32'h8c50000;
      113186: inst = 32'h24612800;
      113187: inst = 32'h10a00000;
      113188: inst = 32'hca0001a;
      113189: inst = 32'h24822800;
      113190: inst = 32'h10a00000;
      113191: inst = 32'hca00004;
      113192: inst = 32'h38632800;
      113193: inst = 32'h38842800;
      113194: inst = 32'h10a00001;
      113195: inst = 32'hca0ba2f;
      113196: inst = 32'h13e00001;
      113197: inst = 32'hfe0d96a;
      113198: inst = 32'h5be00000;
      113199: inst = 32'h8c50000;
      113200: inst = 32'h24612800;
      113201: inst = 32'h10a00000;
      113202: inst = 32'hca0001a;
      113203: inst = 32'h24822800;
      113204: inst = 32'h10a00000;
      113205: inst = 32'hca00004;
      113206: inst = 32'h38632800;
      113207: inst = 32'h38842800;
      113208: inst = 32'h10a00001;
      113209: inst = 32'hca0ba3d;
      113210: inst = 32'h13e00001;
      113211: inst = 32'hfe0d96a;
      113212: inst = 32'h5be00000;
      113213: inst = 32'h8c50000;
      113214: inst = 32'h24612800;
      113215: inst = 32'h10a00000;
      113216: inst = 32'hca0001a;
      113217: inst = 32'h24822800;
      113218: inst = 32'h10a00000;
      113219: inst = 32'hca00004;
      113220: inst = 32'h38632800;
      113221: inst = 32'h38842800;
      113222: inst = 32'h10a00001;
      113223: inst = 32'hca0ba4b;
      113224: inst = 32'h13e00001;
      113225: inst = 32'hfe0d96a;
      113226: inst = 32'h5be00000;
      113227: inst = 32'h8c50000;
      113228: inst = 32'h24612800;
      113229: inst = 32'h10a00000;
      113230: inst = 32'hca0001a;
      113231: inst = 32'h24822800;
      113232: inst = 32'h10a00000;
      113233: inst = 32'hca00004;
      113234: inst = 32'h38632800;
      113235: inst = 32'h38842800;
      113236: inst = 32'h10a00001;
      113237: inst = 32'hca0ba59;
      113238: inst = 32'h13e00001;
      113239: inst = 32'hfe0d96a;
      113240: inst = 32'h5be00000;
      113241: inst = 32'h8c50000;
      113242: inst = 32'h24612800;
      113243: inst = 32'h10a00000;
      113244: inst = 32'hca0001a;
      113245: inst = 32'h24822800;
      113246: inst = 32'h10a00000;
      113247: inst = 32'hca00004;
      113248: inst = 32'h38632800;
      113249: inst = 32'h38842800;
      113250: inst = 32'h10a00001;
      113251: inst = 32'hca0ba67;
      113252: inst = 32'h13e00001;
      113253: inst = 32'hfe0d96a;
      113254: inst = 32'h5be00000;
      113255: inst = 32'h8c50000;
      113256: inst = 32'h24612800;
      113257: inst = 32'h10a00000;
      113258: inst = 32'hca0001a;
      113259: inst = 32'h24822800;
      113260: inst = 32'h10a00000;
      113261: inst = 32'hca00004;
      113262: inst = 32'h38632800;
      113263: inst = 32'h38842800;
      113264: inst = 32'h10a00001;
      113265: inst = 32'hca0ba75;
      113266: inst = 32'h13e00001;
      113267: inst = 32'hfe0d96a;
      113268: inst = 32'h5be00000;
      113269: inst = 32'h8c50000;
      113270: inst = 32'h24612800;
      113271: inst = 32'h10a00000;
      113272: inst = 32'hca0001a;
      113273: inst = 32'h24822800;
      113274: inst = 32'h10a00000;
      113275: inst = 32'hca00004;
      113276: inst = 32'h38632800;
      113277: inst = 32'h38842800;
      113278: inst = 32'h10a00001;
      113279: inst = 32'hca0ba83;
      113280: inst = 32'h13e00001;
      113281: inst = 32'hfe0d96a;
      113282: inst = 32'h5be00000;
      113283: inst = 32'h8c50000;
      113284: inst = 32'h24612800;
      113285: inst = 32'h10a00000;
      113286: inst = 32'hca0001a;
      113287: inst = 32'h24822800;
      113288: inst = 32'h10a00000;
      113289: inst = 32'hca00004;
      113290: inst = 32'h38632800;
      113291: inst = 32'h38842800;
      113292: inst = 32'h10a00001;
      113293: inst = 32'hca0ba91;
      113294: inst = 32'h13e00001;
      113295: inst = 32'hfe0d96a;
      113296: inst = 32'h5be00000;
      113297: inst = 32'h8c50000;
      113298: inst = 32'h24612800;
      113299: inst = 32'h10a00000;
      113300: inst = 32'hca0001a;
      113301: inst = 32'h24822800;
      113302: inst = 32'h10a00000;
      113303: inst = 32'hca00004;
      113304: inst = 32'h38632800;
      113305: inst = 32'h38842800;
      113306: inst = 32'h10a00001;
      113307: inst = 32'hca0ba9f;
      113308: inst = 32'h13e00001;
      113309: inst = 32'hfe0d96a;
      113310: inst = 32'h5be00000;
      113311: inst = 32'h8c50000;
      113312: inst = 32'h24612800;
      113313: inst = 32'h10a00000;
      113314: inst = 32'hca0001a;
      113315: inst = 32'h24822800;
      113316: inst = 32'h10a00000;
      113317: inst = 32'hca00004;
      113318: inst = 32'h38632800;
      113319: inst = 32'h38842800;
      113320: inst = 32'h10a00001;
      113321: inst = 32'hca0baad;
      113322: inst = 32'h13e00001;
      113323: inst = 32'hfe0d96a;
      113324: inst = 32'h5be00000;
      113325: inst = 32'h8c50000;
      113326: inst = 32'h24612800;
      113327: inst = 32'h10a00000;
      113328: inst = 32'hca0001a;
      113329: inst = 32'h24822800;
      113330: inst = 32'h10a00000;
      113331: inst = 32'hca00004;
      113332: inst = 32'h38632800;
      113333: inst = 32'h38842800;
      113334: inst = 32'h10a00001;
      113335: inst = 32'hca0babb;
      113336: inst = 32'h13e00001;
      113337: inst = 32'hfe0d96a;
      113338: inst = 32'h5be00000;
      113339: inst = 32'h8c50000;
      113340: inst = 32'h24612800;
      113341: inst = 32'h10a00000;
      113342: inst = 32'hca0001a;
      113343: inst = 32'h24822800;
      113344: inst = 32'h10a00000;
      113345: inst = 32'hca00004;
      113346: inst = 32'h38632800;
      113347: inst = 32'h38842800;
      113348: inst = 32'h10a00001;
      113349: inst = 32'hca0bac9;
      113350: inst = 32'h13e00001;
      113351: inst = 32'hfe0d96a;
      113352: inst = 32'h5be00000;
      113353: inst = 32'h8c50000;
      113354: inst = 32'h24612800;
      113355: inst = 32'h10a00000;
      113356: inst = 32'hca0001a;
      113357: inst = 32'h24822800;
      113358: inst = 32'h10a00000;
      113359: inst = 32'hca00004;
      113360: inst = 32'h38632800;
      113361: inst = 32'h38842800;
      113362: inst = 32'h10a00001;
      113363: inst = 32'hca0bad7;
      113364: inst = 32'h13e00001;
      113365: inst = 32'hfe0d96a;
      113366: inst = 32'h5be00000;
      113367: inst = 32'h8c50000;
      113368: inst = 32'h24612800;
      113369: inst = 32'h10a00000;
      113370: inst = 32'hca0001a;
      113371: inst = 32'h24822800;
      113372: inst = 32'h10a00000;
      113373: inst = 32'hca00004;
      113374: inst = 32'h38632800;
      113375: inst = 32'h38842800;
      113376: inst = 32'h10a00001;
      113377: inst = 32'hca0bae5;
      113378: inst = 32'h13e00001;
      113379: inst = 32'hfe0d96a;
      113380: inst = 32'h5be00000;
      113381: inst = 32'h8c50000;
      113382: inst = 32'h24612800;
      113383: inst = 32'h10a00000;
      113384: inst = 32'hca0001a;
      113385: inst = 32'h24822800;
      113386: inst = 32'h10a00000;
      113387: inst = 32'hca00004;
      113388: inst = 32'h38632800;
      113389: inst = 32'h38842800;
      113390: inst = 32'h10a00001;
      113391: inst = 32'hca0baf3;
      113392: inst = 32'h13e00001;
      113393: inst = 32'hfe0d96a;
      113394: inst = 32'h5be00000;
      113395: inst = 32'h8c50000;
      113396: inst = 32'h24612800;
      113397: inst = 32'h10a00000;
      113398: inst = 32'hca0001a;
      113399: inst = 32'h24822800;
      113400: inst = 32'h10a00000;
      113401: inst = 32'hca00004;
      113402: inst = 32'h38632800;
      113403: inst = 32'h38842800;
      113404: inst = 32'h10a00001;
      113405: inst = 32'hca0bb01;
      113406: inst = 32'h13e00001;
      113407: inst = 32'hfe0d96a;
      113408: inst = 32'h5be00000;
      113409: inst = 32'h8c50000;
      113410: inst = 32'h24612800;
      113411: inst = 32'h10a00000;
      113412: inst = 32'hca0001a;
      113413: inst = 32'h24822800;
      113414: inst = 32'h10a00000;
      113415: inst = 32'hca00004;
      113416: inst = 32'h38632800;
      113417: inst = 32'h38842800;
      113418: inst = 32'h10a00001;
      113419: inst = 32'hca0bb0f;
      113420: inst = 32'h13e00001;
      113421: inst = 32'hfe0d96a;
      113422: inst = 32'h5be00000;
      113423: inst = 32'h8c50000;
      113424: inst = 32'h24612800;
      113425: inst = 32'h10a00000;
      113426: inst = 32'hca0001a;
      113427: inst = 32'h24822800;
      113428: inst = 32'h10a00000;
      113429: inst = 32'hca00004;
      113430: inst = 32'h38632800;
      113431: inst = 32'h38842800;
      113432: inst = 32'h10a00001;
      113433: inst = 32'hca0bb1d;
      113434: inst = 32'h13e00001;
      113435: inst = 32'hfe0d96a;
      113436: inst = 32'h5be00000;
      113437: inst = 32'h8c50000;
      113438: inst = 32'h24612800;
      113439: inst = 32'h10a00000;
      113440: inst = 32'hca0001a;
      113441: inst = 32'h24822800;
      113442: inst = 32'h10a00000;
      113443: inst = 32'hca00004;
      113444: inst = 32'h38632800;
      113445: inst = 32'h38842800;
      113446: inst = 32'h10a00001;
      113447: inst = 32'hca0bb2b;
      113448: inst = 32'h13e00001;
      113449: inst = 32'hfe0d96a;
      113450: inst = 32'h5be00000;
      113451: inst = 32'h8c50000;
      113452: inst = 32'h24612800;
      113453: inst = 32'h10a00000;
      113454: inst = 32'hca0001a;
      113455: inst = 32'h24822800;
      113456: inst = 32'h10a00000;
      113457: inst = 32'hca00004;
      113458: inst = 32'h38632800;
      113459: inst = 32'h38842800;
      113460: inst = 32'h10a00001;
      113461: inst = 32'hca0bb39;
      113462: inst = 32'h13e00001;
      113463: inst = 32'hfe0d96a;
      113464: inst = 32'h5be00000;
      113465: inst = 32'h8c50000;
      113466: inst = 32'h24612800;
      113467: inst = 32'h10a00000;
      113468: inst = 32'hca0001a;
      113469: inst = 32'h24822800;
      113470: inst = 32'h10a00000;
      113471: inst = 32'hca00004;
      113472: inst = 32'h38632800;
      113473: inst = 32'h38842800;
      113474: inst = 32'h10a00001;
      113475: inst = 32'hca0bb47;
      113476: inst = 32'h13e00001;
      113477: inst = 32'hfe0d96a;
      113478: inst = 32'h5be00000;
      113479: inst = 32'h8c50000;
      113480: inst = 32'h24612800;
      113481: inst = 32'h10a00000;
      113482: inst = 32'hca0001a;
      113483: inst = 32'h24822800;
      113484: inst = 32'h10a00000;
      113485: inst = 32'hca00004;
      113486: inst = 32'h38632800;
      113487: inst = 32'h38842800;
      113488: inst = 32'h10a00001;
      113489: inst = 32'hca0bb55;
      113490: inst = 32'h13e00001;
      113491: inst = 32'hfe0d96a;
      113492: inst = 32'h5be00000;
      113493: inst = 32'h8c50000;
      113494: inst = 32'h24612800;
      113495: inst = 32'h10a00000;
      113496: inst = 32'hca0001a;
      113497: inst = 32'h24822800;
      113498: inst = 32'h10a00000;
      113499: inst = 32'hca00004;
      113500: inst = 32'h38632800;
      113501: inst = 32'h38842800;
      113502: inst = 32'h10a00001;
      113503: inst = 32'hca0bb63;
      113504: inst = 32'h13e00001;
      113505: inst = 32'hfe0d96a;
      113506: inst = 32'h5be00000;
      113507: inst = 32'h8c50000;
      113508: inst = 32'h24612800;
      113509: inst = 32'h10a00000;
      113510: inst = 32'hca0001a;
      113511: inst = 32'h24822800;
      113512: inst = 32'h10a00000;
      113513: inst = 32'hca00004;
      113514: inst = 32'h38632800;
      113515: inst = 32'h38842800;
      113516: inst = 32'h10a00001;
      113517: inst = 32'hca0bb71;
      113518: inst = 32'h13e00001;
      113519: inst = 32'hfe0d96a;
      113520: inst = 32'h5be00000;
      113521: inst = 32'h8c50000;
      113522: inst = 32'h24612800;
      113523: inst = 32'h10a00000;
      113524: inst = 32'hca0001a;
      113525: inst = 32'h24822800;
      113526: inst = 32'h10a00000;
      113527: inst = 32'hca00004;
      113528: inst = 32'h38632800;
      113529: inst = 32'h38842800;
      113530: inst = 32'h10a00001;
      113531: inst = 32'hca0bb7f;
      113532: inst = 32'h13e00001;
      113533: inst = 32'hfe0d96a;
      113534: inst = 32'h5be00000;
      113535: inst = 32'h8c50000;
      113536: inst = 32'h24612800;
      113537: inst = 32'h10a00000;
      113538: inst = 32'hca0001a;
      113539: inst = 32'h24822800;
      113540: inst = 32'h10a00000;
      113541: inst = 32'hca00004;
      113542: inst = 32'h38632800;
      113543: inst = 32'h38842800;
      113544: inst = 32'h10a00001;
      113545: inst = 32'hca0bb8d;
      113546: inst = 32'h13e00001;
      113547: inst = 32'hfe0d96a;
      113548: inst = 32'h5be00000;
      113549: inst = 32'h8c50000;
      113550: inst = 32'h24612800;
      113551: inst = 32'h10a00000;
      113552: inst = 32'hca0001a;
      113553: inst = 32'h24822800;
      113554: inst = 32'h10a00000;
      113555: inst = 32'hca00004;
      113556: inst = 32'h38632800;
      113557: inst = 32'h38842800;
      113558: inst = 32'h10a00001;
      113559: inst = 32'hca0bb9b;
      113560: inst = 32'h13e00001;
      113561: inst = 32'hfe0d96a;
      113562: inst = 32'h5be00000;
      113563: inst = 32'h8c50000;
      113564: inst = 32'h24612800;
      113565: inst = 32'h10a00000;
      113566: inst = 32'hca0001a;
      113567: inst = 32'h24822800;
      113568: inst = 32'h10a00000;
      113569: inst = 32'hca00004;
      113570: inst = 32'h38632800;
      113571: inst = 32'h38842800;
      113572: inst = 32'h10a00001;
      113573: inst = 32'hca0bba9;
      113574: inst = 32'h13e00001;
      113575: inst = 32'hfe0d96a;
      113576: inst = 32'h5be00000;
      113577: inst = 32'h8c50000;
      113578: inst = 32'h24612800;
      113579: inst = 32'h10a00000;
      113580: inst = 32'hca0001a;
      113581: inst = 32'h24822800;
      113582: inst = 32'h10a00000;
      113583: inst = 32'hca00004;
      113584: inst = 32'h38632800;
      113585: inst = 32'h38842800;
      113586: inst = 32'h10a00001;
      113587: inst = 32'hca0bbb7;
      113588: inst = 32'h13e00001;
      113589: inst = 32'hfe0d96a;
      113590: inst = 32'h5be00000;
      113591: inst = 32'h8c50000;
      113592: inst = 32'h24612800;
      113593: inst = 32'h10a00000;
      113594: inst = 32'hca0001a;
      113595: inst = 32'h24822800;
      113596: inst = 32'h10a00000;
      113597: inst = 32'hca00004;
      113598: inst = 32'h38632800;
      113599: inst = 32'h38842800;
      113600: inst = 32'h10a00001;
      113601: inst = 32'hca0bbc5;
      113602: inst = 32'h13e00001;
      113603: inst = 32'hfe0d96a;
      113604: inst = 32'h5be00000;
      113605: inst = 32'h8c50000;
      113606: inst = 32'h24612800;
      113607: inst = 32'h10a00000;
      113608: inst = 32'hca0001a;
      113609: inst = 32'h24822800;
      113610: inst = 32'h10a00000;
      113611: inst = 32'hca00004;
      113612: inst = 32'h38632800;
      113613: inst = 32'h38842800;
      113614: inst = 32'h10a00001;
      113615: inst = 32'hca0bbd3;
      113616: inst = 32'h13e00001;
      113617: inst = 32'hfe0d96a;
      113618: inst = 32'h5be00000;
      113619: inst = 32'h8c50000;
      113620: inst = 32'h24612800;
      113621: inst = 32'h10a00000;
      113622: inst = 32'hca0001a;
      113623: inst = 32'h24822800;
      113624: inst = 32'h10a00000;
      113625: inst = 32'hca00004;
      113626: inst = 32'h38632800;
      113627: inst = 32'h38842800;
      113628: inst = 32'h10a00001;
      113629: inst = 32'hca0bbe1;
      113630: inst = 32'h13e00001;
      113631: inst = 32'hfe0d96a;
      113632: inst = 32'h5be00000;
      113633: inst = 32'h8c50000;
      113634: inst = 32'h24612800;
      113635: inst = 32'h10a00000;
      113636: inst = 32'hca0001a;
      113637: inst = 32'h24822800;
      113638: inst = 32'h10a00000;
      113639: inst = 32'hca00004;
      113640: inst = 32'h38632800;
      113641: inst = 32'h38842800;
      113642: inst = 32'h10a00001;
      113643: inst = 32'hca0bbef;
      113644: inst = 32'h13e00001;
      113645: inst = 32'hfe0d96a;
      113646: inst = 32'h5be00000;
      113647: inst = 32'h8c50000;
      113648: inst = 32'h24612800;
      113649: inst = 32'h10a00000;
      113650: inst = 32'hca0001a;
      113651: inst = 32'h24822800;
      113652: inst = 32'h10a00000;
      113653: inst = 32'hca00004;
      113654: inst = 32'h38632800;
      113655: inst = 32'h38842800;
      113656: inst = 32'h10a00001;
      113657: inst = 32'hca0bbfd;
      113658: inst = 32'h13e00001;
      113659: inst = 32'hfe0d96a;
      113660: inst = 32'h5be00000;
      113661: inst = 32'h8c50000;
      113662: inst = 32'h24612800;
      113663: inst = 32'h10a00000;
      113664: inst = 32'hca0001a;
      113665: inst = 32'h24822800;
      113666: inst = 32'h10a00000;
      113667: inst = 32'hca00004;
      113668: inst = 32'h38632800;
      113669: inst = 32'h38842800;
      113670: inst = 32'h10a00001;
      113671: inst = 32'hca0bc0b;
      113672: inst = 32'h13e00001;
      113673: inst = 32'hfe0d96a;
      113674: inst = 32'h5be00000;
      113675: inst = 32'h8c50000;
      113676: inst = 32'h24612800;
      113677: inst = 32'h10a00000;
      113678: inst = 32'hca0001a;
      113679: inst = 32'h24822800;
      113680: inst = 32'h10a00000;
      113681: inst = 32'hca00004;
      113682: inst = 32'h38632800;
      113683: inst = 32'h38842800;
      113684: inst = 32'h10a00001;
      113685: inst = 32'hca0bc19;
      113686: inst = 32'h13e00001;
      113687: inst = 32'hfe0d96a;
      113688: inst = 32'h5be00000;
      113689: inst = 32'h8c50000;
      113690: inst = 32'h24612800;
      113691: inst = 32'h10a00000;
      113692: inst = 32'hca0001a;
      113693: inst = 32'h24822800;
      113694: inst = 32'h10a00000;
      113695: inst = 32'hca00004;
      113696: inst = 32'h38632800;
      113697: inst = 32'h38842800;
      113698: inst = 32'h10a00001;
      113699: inst = 32'hca0bc27;
      113700: inst = 32'h13e00001;
      113701: inst = 32'hfe0d96a;
      113702: inst = 32'h5be00000;
      113703: inst = 32'h8c50000;
      113704: inst = 32'h24612800;
      113705: inst = 32'h10a00000;
      113706: inst = 32'hca0001a;
      113707: inst = 32'h24822800;
      113708: inst = 32'h10a00000;
      113709: inst = 32'hca00004;
      113710: inst = 32'h38632800;
      113711: inst = 32'h38842800;
      113712: inst = 32'h10a00001;
      113713: inst = 32'hca0bc35;
      113714: inst = 32'h13e00001;
      113715: inst = 32'hfe0d96a;
      113716: inst = 32'h5be00000;
      113717: inst = 32'h8c50000;
      113718: inst = 32'h24612800;
      113719: inst = 32'h10a00000;
      113720: inst = 32'hca0001a;
      113721: inst = 32'h24822800;
      113722: inst = 32'h10a00000;
      113723: inst = 32'hca00004;
      113724: inst = 32'h38632800;
      113725: inst = 32'h38842800;
      113726: inst = 32'h10a00001;
      113727: inst = 32'hca0bc43;
      113728: inst = 32'h13e00001;
      113729: inst = 32'hfe0d96a;
      113730: inst = 32'h5be00000;
      113731: inst = 32'h8c50000;
      113732: inst = 32'h24612800;
      113733: inst = 32'h10a00000;
      113734: inst = 32'hca0001a;
      113735: inst = 32'h24822800;
      113736: inst = 32'h10a00000;
      113737: inst = 32'hca00004;
      113738: inst = 32'h38632800;
      113739: inst = 32'h38842800;
      113740: inst = 32'h10a00001;
      113741: inst = 32'hca0bc51;
      113742: inst = 32'h13e00001;
      113743: inst = 32'hfe0d96a;
      113744: inst = 32'h5be00000;
      113745: inst = 32'h8c50000;
      113746: inst = 32'h24612800;
      113747: inst = 32'h10a00000;
      113748: inst = 32'hca0001a;
      113749: inst = 32'h24822800;
      113750: inst = 32'h10a00000;
      113751: inst = 32'hca00004;
      113752: inst = 32'h38632800;
      113753: inst = 32'h38842800;
      113754: inst = 32'h10a00001;
      113755: inst = 32'hca0bc5f;
      113756: inst = 32'h13e00001;
      113757: inst = 32'hfe0d96a;
      113758: inst = 32'h5be00000;
      113759: inst = 32'h8c50000;
      113760: inst = 32'h24612800;
      113761: inst = 32'h10a00000;
      113762: inst = 32'hca0001a;
      113763: inst = 32'h24822800;
      113764: inst = 32'h10a00000;
      113765: inst = 32'hca00004;
      113766: inst = 32'h38632800;
      113767: inst = 32'h38842800;
      113768: inst = 32'h10a00001;
      113769: inst = 32'hca0bc6d;
      113770: inst = 32'h13e00001;
      113771: inst = 32'hfe0d96a;
      113772: inst = 32'h5be00000;
      113773: inst = 32'h8c50000;
      113774: inst = 32'h24612800;
      113775: inst = 32'h10a00000;
      113776: inst = 32'hca0001a;
      113777: inst = 32'h24822800;
      113778: inst = 32'h10a00000;
      113779: inst = 32'hca00004;
      113780: inst = 32'h38632800;
      113781: inst = 32'h38842800;
      113782: inst = 32'h10a00001;
      113783: inst = 32'hca0bc7b;
      113784: inst = 32'h13e00001;
      113785: inst = 32'hfe0d96a;
      113786: inst = 32'h5be00000;
      113787: inst = 32'h8c50000;
      113788: inst = 32'h24612800;
      113789: inst = 32'h10a00000;
      113790: inst = 32'hca0001a;
      113791: inst = 32'h24822800;
      113792: inst = 32'h10a00000;
      113793: inst = 32'hca00004;
      113794: inst = 32'h38632800;
      113795: inst = 32'h38842800;
      113796: inst = 32'h10a00001;
      113797: inst = 32'hca0bc89;
      113798: inst = 32'h13e00001;
      113799: inst = 32'hfe0d96a;
      113800: inst = 32'h5be00000;
      113801: inst = 32'h8c50000;
      113802: inst = 32'h24612800;
      113803: inst = 32'h10a00000;
      113804: inst = 32'hca0001a;
      113805: inst = 32'h24822800;
      113806: inst = 32'h10a00000;
      113807: inst = 32'hca00004;
      113808: inst = 32'h38632800;
      113809: inst = 32'h38842800;
      113810: inst = 32'h10a00001;
      113811: inst = 32'hca0bc97;
      113812: inst = 32'h13e00001;
      113813: inst = 32'hfe0d96a;
      113814: inst = 32'h5be00000;
      113815: inst = 32'h8c50000;
      113816: inst = 32'h24612800;
      113817: inst = 32'h10a00000;
      113818: inst = 32'hca0001a;
      113819: inst = 32'h24822800;
      113820: inst = 32'h10a00000;
      113821: inst = 32'hca00004;
      113822: inst = 32'h38632800;
      113823: inst = 32'h38842800;
      113824: inst = 32'h10a00001;
      113825: inst = 32'hca0bca5;
      113826: inst = 32'h13e00001;
      113827: inst = 32'hfe0d96a;
      113828: inst = 32'h5be00000;
      113829: inst = 32'h8c50000;
      113830: inst = 32'h24612800;
      113831: inst = 32'h10a00000;
      113832: inst = 32'hca0001a;
      113833: inst = 32'h24822800;
      113834: inst = 32'h10a00000;
      113835: inst = 32'hca00004;
      113836: inst = 32'h38632800;
      113837: inst = 32'h38842800;
      113838: inst = 32'h10a00001;
      113839: inst = 32'hca0bcb3;
      113840: inst = 32'h13e00001;
      113841: inst = 32'hfe0d96a;
      113842: inst = 32'h5be00000;
      113843: inst = 32'h8c50000;
      113844: inst = 32'h24612800;
      113845: inst = 32'h10a00000;
      113846: inst = 32'hca0001a;
      113847: inst = 32'h24822800;
      113848: inst = 32'h10a00000;
      113849: inst = 32'hca00004;
      113850: inst = 32'h38632800;
      113851: inst = 32'h38842800;
      113852: inst = 32'h10a00001;
      113853: inst = 32'hca0bcc1;
      113854: inst = 32'h13e00001;
      113855: inst = 32'hfe0d96a;
      113856: inst = 32'h5be00000;
      113857: inst = 32'h8c50000;
      113858: inst = 32'h24612800;
      113859: inst = 32'h10a00000;
      113860: inst = 32'hca0001a;
      113861: inst = 32'h24822800;
      113862: inst = 32'h10a00000;
      113863: inst = 32'hca00004;
      113864: inst = 32'h38632800;
      113865: inst = 32'h38842800;
      113866: inst = 32'h10a00001;
      113867: inst = 32'hca0bccf;
      113868: inst = 32'h13e00001;
      113869: inst = 32'hfe0d96a;
      113870: inst = 32'h5be00000;
      113871: inst = 32'h8c50000;
      113872: inst = 32'h24612800;
      113873: inst = 32'h10a00000;
      113874: inst = 32'hca0001a;
      113875: inst = 32'h24822800;
      113876: inst = 32'h10a00000;
      113877: inst = 32'hca00004;
      113878: inst = 32'h38632800;
      113879: inst = 32'h38842800;
      113880: inst = 32'h10a00001;
      113881: inst = 32'hca0bcdd;
      113882: inst = 32'h13e00001;
      113883: inst = 32'hfe0d96a;
      113884: inst = 32'h5be00000;
      113885: inst = 32'h8c50000;
      113886: inst = 32'h24612800;
      113887: inst = 32'h10a00000;
      113888: inst = 32'hca0001a;
      113889: inst = 32'h24822800;
      113890: inst = 32'h10a00000;
      113891: inst = 32'hca00004;
      113892: inst = 32'h38632800;
      113893: inst = 32'h38842800;
      113894: inst = 32'h10a00001;
      113895: inst = 32'hca0bceb;
      113896: inst = 32'h13e00001;
      113897: inst = 32'hfe0d96a;
      113898: inst = 32'h5be00000;
      113899: inst = 32'h8c50000;
      113900: inst = 32'h24612800;
      113901: inst = 32'h10a00000;
      113902: inst = 32'hca0001a;
      113903: inst = 32'h24822800;
      113904: inst = 32'h10a00000;
      113905: inst = 32'hca00004;
      113906: inst = 32'h38632800;
      113907: inst = 32'h38842800;
      113908: inst = 32'h10a00001;
      113909: inst = 32'hca0bcf9;
      113910: inst = 32'h13e00001;
      113911: inst = 32'hfe0d96a;
      113912: inst = 32'h5be00000;
      113913: inst = 32'h8c50000;
      113914: inst = 32'h24612800;
      113915: inst = 32'h10a00000;
      113916: inst = 32'hca0001a;
      113917: inst = 32'h24822800;
      113918: inst = 32'h10a00000;
      113919: inst = 32'hca00004;
      113920: inst = 32'h38632800;
      113921: inst = 32'h38842800;
      113922: inst = 32'h10a00001;
      113923: inst = 32'hca0bd07;
      113924: inst = 32'h13e00001;
      113925: inst = 32'hfe0d96a;
      113926: inst = 32'h5be00000;
      113927: inst = 32'h8c50000;
      113928: inst = 32'h24612800;
      113929: inst = 32'h10a00000;
      113930: inst = 32'hca0001a;
      113931: inst = 32'h24822800;
      113932: inst = 32'h10a00000;
      113933: inst = 32'hca00004;
      113934: inst = 32'h38632800;
      113935: inst = 32'h38842800;
      113936: inst = 32'h10a00001;
      113937: inst = 32'hca0bd15;
      113938: inst = 32'h13e00001;
      113939: inst = 32'hfe0d96a;
      113940: inst = 32'h5be00000;
      113941: inst = 32'h8c50000;
      113942: inst = 32'h24612800;
      113943: inst = 32'h10a00000;
      113944: inst = 32'hca0001a;
      113945: inst = 32'h24822800;
      113946: inst = 32'h10a00000;
      113947: inst = 32'hca00004;
      113948: inst = 32'h38632800;
      113949: inst = 32'h38842800;
      113950: inst = 32'h10a00001;
      113951: inst = 32'hca0bd23;
      113952: inst = 32'h13e00001;
      113953: inst = 32'hfe0d96a;
      113954: inst = 32'h5be00000;
      113955: inst = 32'h8c50000;
      113956: inst = 32'h24612800;
      113957: inst = 32'h10a00000;
      113958: inst = 32'hca0001a;
      113959: inst = 32'h24822800;
      113960: inst = 32'h10a00000;
      113961: inst = 32'hca00004;
      113962: inst = 32'h38632800;
      113963: inst = 32'h38842800;
      113964: inst = 32'h10a00001;
      113965: inst = 32'hca0bd31;
      113966: inst = 32'h13e00001;
      113967: inst = 32'hfe0d96a;
      113968: inst = 32'h5be00000;
      113969: inst = 32'h8c50000;
      113970: inst = 32'h24612800;
      113971: inst = 32'h10a00000;
      113972: inst = 32'hca0001a;
      113973: inst = 32'h24822800;
      113974: inst = 32'h10a00000;
      113975: inst = 32'hca00004;
      113976: inst = 32'h38632800;
      113977: inst = 32'h38842800;
      113978: inst = 32'h10a00001;
      113979: inst = 32'hca0bd3f;
      113980: inst = 32'h13e00001;
      113981: inst = 32'hfe0d96a;
      113982: inst = 32'h5be00000;
      113983: inst = 32'h8c50000;
      113984: inst = 32'h24612800;
      113985: inst = 32'h10a00000;
      113986: inst = 32'hca0001a;
      113987: inst = 32'h24822800;
      113988: inst = 32'h10a00000;
      113989: inst = 32'hca00004;
      113990: inst = 32'h38632800;
      113991: inst = 32'h38842800;
      113992: inst = 32'h10a00001;
      113993: inst = 32'hca0bd4d;
      113994: inst = 32'h13e00001;
      113995: inst = 32'hfe0d96a;
      113996: inst = 32'h5be00000;
      113997: inst = 32'h8c50000;
      113998: inst = 32'h24612800;
      113999: inst = 32'h10a00000;
      114000: inst = 32'hca0001a;
      114001: inst = 32'h24822800;
      114002: inst = 32'h10a00000;
      114003: inst = 32'hca00004;
      114004: inst = 32'h38632800;
      114005: inst = 32'h38842800;
      114006: inst = 32'h10a00001;
      114007: inst = 32'hca0bd5b;
      114008: inst = 32'h13e00001;
      114009: inst = 32'hfe0d96a;
      114010: inst = 32'h5be00000;
      114011: inst = 32'h8c50000;
      114012: inst = 32'h24612800;
      114013: inst = 32'h10a00000;
      114014: inst = 32'hca0001a;
      114015: inst = 32'h24822800;
      114016: inst = 32'h10a00000;
      114017: inst = 32'hca00004;
      114018: inst = 32'h38632800;
      114019: inst = 32'h38842800;
      114020: inst = 32'h10a00001;
      114021: inst = 32'hca0bd69;
      114022: inst = 32'h13e00001;
      114023: inst = 32'hfe0d96a;
      114024: inst = 32'h5be00000;
      114025: inst = 32'h8c50000;
      114026: inst = 32'h24612800;
      114027: inst = 32'h10a00000;
      114028: inst = 32'hca0001a;
      114029: inst = 32'h24822800;
      114030: inst = 32'h10a00000;
      114031: inst = 32'hca00004;
      114032: inst = 32'h38632800;
      114033: inst = 32'h38842800;
      114034: inst = 32'h10a00001;
      114035: inst = 32'hca0bd77;
      114036: inst = 32'h13e00001;
      114037: inst = 32'hfe0d96a;
      114038: inst = 32'h5be00000;
      114039: inst = 32'h8c50000;
      114040: inst = 32'h24612800;
      114041: inst = 32'h10a00000;
      114042: inst = 32'hca0001a;
      114043: inst = 32'h24822800;
      114044: inst = 32'h10a00000;
      114045: inst = 32'hca00004;
      114046: inst = 32'h38632800;
      114047: inst = 32'h38842800;
      114048: inst = 32'h10a00001;
      114049: inst = 32'hca0bd85;
      114050: inst = 32'h13e00001;
      114051: inst = 32'hfe0d96a;
      114052: inst = 32'h5be00000;
      114053: inst = 32'h8c50000;
      114054: inst = 32'h24612800;
      114055: inst = 32'h10a00000;
      114056: inst = 32'hca0001a;
      114057: inst = 32'h24822800;
      114058: inst = 32'h10a00000;
      114059: inst = 32'hca00004;
      114060: inst = 32'h38632800;
      114061: inst = 32'h38842800;
      114062: inst = 32'h10a00001;
      114063: inst = 32'hca0bd93;
      114064: inst = 32'h13e00001;
      114065: inst = 32'hfe0d96a;
      114066: inst = 32'h5be00000;
      114067: inst = 32'h8c50000;
      114068: inst = 32'h24612800;
      114069: inst = 32'h10a00000;
      114070: inst = 32'hca0001a;
      114071: inst = 32'h24822800;
      114072: inst = 32'h10a00000;
      114073: inst = 32'hca00004;
      114074: inst = 32'h38632800;
      114075: inst = 32'h38842800;
      114076: inst = 32'h10a00001;
      114077: inst = 32'hca0bda1;
      114078: inst = 32'h13e00001;
      114079: inst = 32'hfe0d96a;
      114080: inst = 32'h5be00000;
      114081: inst = 32'h8c50000;
      114082: inst = 32'h24612800;
      114083: inst = 32'h10a00000;
      114084: inst = 32'hca0001a;
      114085: inst = 32'h24822800;
      114086: inst = 32'h10a00000;
      114087: inst = 32'hca00004;
      114088: inst = 32'h38632800;
      114089: inst = 32'h38842800;
      114090: inst = 32'h10a00001;
      114091: inst = 32'hca0bdaf;
      114092: inst = 32'h13e00001;
      114093: inst = 32'hfe0d96a;
      114094: inst = 32'h5be00000;
      114095: inst = 32'h8c50000;
      114096: inst = 32'h24612800;
      114097: inst = 32'h10a00000;
      114098: inst = 32'hca0001a;
      114099: inst = 32'h24822800;
      114100: inst = 32'h10a00000;
      114101: inst = 32'hca00004;
      114102: inst = 32'h38632800;
      114103: inst = 32'h38842800;
      114104: inst = 32'h10a00001;
      114105: inst = 32'hca0bdbd;
      114106: inst = 32'h13e00001;
      114107: inst = 32'hfe0d96a;
      114108: inst = 32'h5be00000;
      114109: inst = 32'h8c50000;
      114110: inst = 32'h24612800;
      114111: inst = 32'h10a00000;
      114112: inst = 32'hca0001a;
      114113: inst = 32'h24822800;
      114114: inst = 32'h10a00000;
      114115: inst = 32'hca00004;
      114116: inst = 32'h38632800;
      114117: inst = 32'h38842800;
      114118: inst = 32'h10a00001;
      114119: inst = 32'hca0bdcb;
      114120: inst = 32'h13e00001;
      114121: inst = 32'hfe0d96a;
      114122: inst = 32'h5be00000;
      114123: inst = 32'h8c50000;
      114124: inst = 32'h24612800;
      114125: inst = 32'h10a00000;
      114126: inst = 32'hca0001a;
      114127: inst = 32'h24822800;
      114128: inst = 32'h10a00000;
      114129: inst = 32'hca00004;
      114130: inst = 32'h38632800;
      114131: inst = 32'h38842800;
      114132: inst = 32'h10a00001;
      114133: inst = 32'hca0bdd9;
      114134: inst = 32'h13e00001;
      114135: inst = 32'hfe0d96a;
      114136: inst = 32'h5be00000;
      114137: inst = 32'h8c50000;
      114138: inst = 32'h24612800;
      114139: inst = 32'h10a00000;
      114140: inst = 32'hca0001a;
      114141: inst = 32'h24822800;
      114142: inst = 32'h10a00000;
      114143: inst = 32'hca00004;
      114144: inst = 32'h38632800;
      114145: inst = 32'h38842800;
      114146: inst = 32'h10a00001;
      114147: inst = 32'hca0bde7;
      114148: inst = 32'h13e00001;
      114149: inst = 32'hfe0d96a;
      114150: inst = 32'h5be00000;
      114151: inst = 32'h8c50000;
      114152: inst = 32'h24612800;
      114153: inst = 32'h10a00000;
      114154: inst = 32'hca0001a;
      114155: inst = 32'h24822800;
      114156: inst = 32'h10a00000;
      114157: inst = 32'hca00004;
      114158: inst = 32'h38632800;
      114159: inst = 32'h38842800;
      114160: inst = 32'h10a00001;
      114161: inst = 32'hca0bdf5;
      114162: inst = 32'h13e00001;
      114163: inst = 32'hfe0d96a;
      114164: inst = 32'h5be00000;
      114165: inst = 32'h8c50000;
      114166: inst = 32'h24612800;
      114167: inst = 32'h10a00000;
      114168: inst = 32'hca0001a;
      114169: inst = 32'h24822800;
      114170: inst = 32'h10a00000;
      114171: inst = 32'hca00004;
      114172: inst = 32'h38632800;
      114173: inst = 32'h38842800;
      114174: inst = 32'h10a00001;
      114175: inst = 32'hca0be03;
      114176: inst = 32'h13e00001;
      114177: inst = 32'hfe0d96a;
      114178: inst = 32'h5be00000;
      114179: inst = 32'h8c50000;
      114180: inst = 32'h24612800;
      114181: inst = 32'h10a00000;
      114182: inst = 32'hca0001a;
      114183: inst = 32'h24822800;
      114184: inst = 32'h10a00000;
      114185: inst = 32'hca00004;
      114186: inst = 32'h38632800;
      114187: inst = 32'h38842800;
      114188: inst = 32'h10a00001;
      114189: inst = 32'hca0be11;
      114190: inst = 32'h13e00001;
      114191: inst = 32'hfe0d96a;
      114192: inst = 32'h5be00000;
      114193: inst = 32'h8c50000;
      114194: inst = 32'h24612800;
      114195: inst = 32'h10a00000;
      114196: inst = 32'hca0001a;
      114197: inst = 32'h24822800;
      114198: inst = 32'h10a00000;
      114199: inst = 32'hca00004;
      114200: inst = 32'h38632800;
      114201: inst = 32'h38842800;
      114202: inst = 32'h10a00001;
      114203: inst = 32'hca0be1f;
      114204: inst = 32'h13e00001;
      114205: inst = 32'hfe0d96a;
      114206: inst = 32'h5be00000;
      114207: inst = 32'h8c50000;
      114208: inst = 32'h24612800;
      114209: inst = 32'h10a00000;
      114210: inst = 32'hca0001a;
      114211: inst = 32'h24822800;
      114212: inst = 32'h10a00000;
      114213: inst = 32'hca00004;
      114214: inst = 32'h38632800;
      114215: inst = 32'h38842800;
      114216: inst = 32'h10a00001;
      114217: inst = 32'hca0be2d;
      114218: inst = 32'h13e00001;
      114219: inst = 32'hfe0d96a;
      114220: inst = 32'h5be00000;
      114221: inst = 32'h8c50000;
      114222: inst = 32'h24612800;
      114223: inst = 32'h10a00000;
      114224: inst = 32'hca0001a;
      114225: inst = 32'h24822800;
      114226: inst = 32'h10a00000;
      114227: inst = 32'hca00004;
      114228: inst = 32'h38632800;
      114229: inst = 32'h38842800;
      114230: inst = 32'h10a00001;
      114231: inst = 32'hca0be3b;
      114232: inst = 32'h13e00001;
      114233: inst = 32'hfe0d96a;
      114234: inst = 32'h5be00000;
      114235: inst = 32'h8c50000;
      114236: inst = 32'h24612800;
      114237: inst = 32'h10a00000;
      114238: inst = 32'hca0001a;
      114239: inst = 32'h24822800;
      114240: inst = 32'h10a00000;
      114241: inst = 32'hca00004;
      114242: inst = 32'h38632800;
      114243: inst = 32'h38842800;
      114244: inst = 32'h10a00001;
      114245: inst = 32'hca0be49;
      114246: inst = 32'h13e00001;
      114247: inst = 32'hfe0d96a;
      114248: inst = 32'h5be00000;
      114249: inst = 32'h8c50000;
      114250: inst = 32'h24612800;
      114251: inst = 32'h10a00000;
      114252: inst = 32'hca0001a;
      114253: inst = 32'h24822800;
      114254: inst = 32'h10a00000;
      114255: inst = 32'hca00004;
      114256: inst = 32'h38632800;
      114257: inst = 32'h38842800;
      114258: inst = 32'h10a00001;
      114259: inst = 32'hca0be57;
      114260: inst = 32'h13e00001;
      114261: inst = 32'hfe0d96a;
      114262: inst = 32'h5be00000;
      114263: inst = 32'h8c50000;
      114264: inst = 32'h24612800;
      114265: inst = 32'h10a00000;
      114266: inst = 32'hca0001a;
      114267: inst = 32'h24822800;
      114268: inst = 32'h10a00000;
      114269: inst = 32'hca00004;
      114270: inst = 32'h38632800;
      114271: inst = 32'h38842800;
      114272: inst = 32'h10a00001;
      114273: inst = 32'hca0be65;
      114274: inst = 32'h13e00001;
      114275: inst = 32'hfe0d96a;
      114276: inst = 32'h5be00000;
      114277: inst = 32'h8c50000;
      114278: inst = 32'h24612800;
      114279: inst = 32'h10a00000;
      114280: inst = 32'hca0001a;
      114281: inst = 32'h24822800;
      114282: inst = 32'h10a00000;
      114283: inst = 32'hca00004;
      114284: inst = 32'h38632800;
      114285: inst = 32'h38842800;
      114286: inst = 32'h10a00001;
      114287: inst = 32'hca0be73;
      114288: inst = 32'h13e00001;
      114289: inst = 32'hfe0d96a;
      114290: inst = 32'h5be00000;
      114291: inst = 32'h8c50000;
      114292: inst = 32'h24612800;
      114293: inst = 32'h10a00000;
      114294: inst = 32'hca0001a;
      114295: inst = 32'h24822800;
      114296: inst = 32'h10a00000;
      114297: inst = 32'hca00004;
      114298: inst = 32'h38632800;
      114299: inst = 32'h38842800;
      114300: inst = 32'h10a00001;
      114301: inst = 32'hca0be81;
      114302: inst = 32'h13e00001;
      114303: inst = 32'hfe0d96a;
      114304: inst = 32'h5be00000;
      114305: inst = 32'h8c50000;
      114306: inst = 32'h24612800;
      114307: inst = 32'h10a00000;
      114308: inst = 32'hca0001a;
      114309: inst = 32'h24822800;
      114310: inst = 32'h10a00000;
      114311: inst = 32'hca00004;
      114312: inst = 32'h38632800;
      114313: inst = 32'h38842800;
      114314: inst = 32'h10a00001;
      114315: inst = 32'hca0be8f;
      114316: inst = 32'h13e00001;
      114317: inst = 32'hfe0d96a;
      114318: inst = 32'h5be00000;
      114319: inst = 32'h8c50000;
      114320: inst = 32'h24612800;
      114321: inst = 32'h10a00000;
      114322: inst = 32'hca0001a;
      114323: inst = 32'h24822800;
      114324: inst = 32'h10a00000;
      114325: inst = 32'hca00004;
      114326: inst = 32'h38632800;
      114327: inst = 32'h38842800;
      114328: inst = 32'h10a00001;
      114329: inst = 32'hca0be9d;
      114330: inst = 32'h13e00001;
      114331: inst = 32'hfe0d96a;
      114332: inst = 32'h5be00000;
      114333: inst = 32'h8c50000;
      114334: inst = 32'h24612800;
      114335: inst = 32'h10a00000;
      114336: inst = 32'hca0001a;
      114337: inst = 32'h24822800;
      114338: inst = 32'h10a00000;
      114339: inst = 32'hca00004;
      114340: inst = 32'h38632800;
      114341: inst = 32'h38842800;
      114342: inst = 32'h10a00001;
      114343: inst = 32'hca0beab;
      114344: inst = 32'h13e00001;
      114345: inst = 32'hfe0d96a;
      114346: inst = 32'h5be00000;
      114347: inst = 32'h8c50000;
      114348: inst = 32'h24612800;
      114349: inst = 32'h10a00000;
      114350: inst = 32'hca0001a;
      114351: inst = 32'h24822800;
      114352: inst = 32'h10a00000;
      114353: inst = 32'hca00004;
      114354: inst = 32'h38632800;
      114355: inst = 32'h38842800;
      114356: inst = 32'h10a00001;
      114357: inst = 32'hca0beb9;
      114358: inst = 32'h13e00001;
      114359: inst = 32'hfe0d96a;
      114360: inst = 32'h5be00000;
      114361: inst = 32'h8c50000;
      114362: inst = 32'h24612800;
      114363: inst = 32'h10a00000;
      114364: inst = 32'hca0001a;
      114365: inst = 32'h24822800;
      114366: inst = 32'h10a00000;
      114367: inst = 32'hca00004;
      114368: inst = 32'h38632800;
      114369: inst = 32'h38842800;
      114370: inst = 32'h10a00001;
      114371: inst = 32'hca0bec7;
      114372: inst = 32'h13e00001;
      114373: inst = 32'hfe0d96a;
      114374: inst = 32'h5be00000;
      114375: inst = 32'h8c50000;
      114376: inst = 32'h24612800;
      114377: inst = 32'h10a00000;
      114378: inst = 32'hca0001a;
      114379: inst = 32'h24822800;
      114380: inst = 32'h10a00000;
      114381: inst = 32'hca00004;
      114382: inst = 32'h38632800;
      114383: inst = 32'h38842800;
      114384: inst = 32'h10a00001;
      114385: inst = 32'hca0bed5;
      114386: inst = 32'h13e00001;
      114387: inst = 32'hfe0d96a;
      114388: inst = 32'h5be00000;
      114389: inst = 32'h8c50000;
      114390: inst = 32'h24612800;
      114391: inst = 32'h10a00000;
      114392: inst = 32'hca0001a;
      114393: inst = 32'h24822800;
      114394: inst = 32'h10a00000;
      114395: inst = 32'hca00004;
      114396: inst = 32'h38632800;
      114397: inst = 32'h38842800;
      114398: inst = 32'h10a00001;
      114399: inst = 32'hca0bee3;
      114400: inst = 32'h13e00001;
      114401: inst = 32'hfe0d96a;
      114402: inst = 32'h5be00000;
      114403: inst = 32'h8c50000;
      114404: inst = 32'h24612800;
      114405: inst = 32'h10a00000;
      114406: inst = 32'hca0001a;
      114407: inst = 32'h24822800;
      114408: inst = 32'h10a00000;
      114409: inst = 32'hca00004;
      114410: inst = 32'h38632800;
      114411: inst = 32'h38842800;
      114412: inst = 32'h10a00001;
      114413: inst = 32'hca0bef1;
      114414: inst = 32'h13e00001;
      114415: inst = 32'hfe0d96a;
      114416: inst = 32'h5be00000;
      114417: inst = 32'h8c50000;
      114418: inst = 32'h24612800;
      114419: inst = 32'h10a00000;
      114420: inst = 32'hca0001a;
      114421: inst = 32'h24822800;
      114422: inst = 32'h10a00000;
      114423: inst = 32'hca00004;
      114424: inst = 32'h38632800;
      114425: inst = 32'h38842800;
      114426: inst = 32'h10a00001;
      114427: inst = 32'hca0beff;
      114428: inst = 32'h13e00001;
      114429: inst = 32'hfe0d96a;
      114430: inst = 32'h5be00000;
      114431: inst = 32'h8c50000;
      114432: inst = 32'h24612800;
      114433: inst = 32'h10a00000;
      114434: inst = 32'hca0001a;
      114435: inst = 32'h24822800;
      114436: inst = 32'h10a00000;
      114437: inst = 32'hca00004;
      114438: inst = 32'h38632800;
      114439: inst = 32'h38842800;
      114440: inst = 32'h10a00001;
      114441: inst = 32'hca0bf0d;
      114442: inst = 32'h13e00001;
      114443: inst = 32'hfe0d96a;
      114444: inst = 32'h5be00000;
      114445: inst = 32'h8c50000;
      114446: inst = 32'h24612800;
      114447: inst = 32'h10a00000;
      114448: inst = 32'hca0001a;
      114449: inst = 32'h24822800;
      114450: inst = 32'h10a00000;
      114451: inst = 32'hca00004;
      114452: inst = 32'h38632800;
      114453: inst = 32'h38842800;
      114454: inst = 32'h10a00001;
      114455: inst = 32'hca0bf1b;
      114456: inst = 32'h13e00001;
      114457: inst = 32'hfe0d96a;
      114458: inst = 32'h5be00000;
      114459: inst = 32'h8c50000;
      114460: inst = 32'h24612800;
      114461: inst = 32'h10a00000;
      114462: inst = 32'hca0001a;
      114463: inst = 32'h24822800;
      114464: inst = 32'h10a00000;
      114465: inst = 32'hca00004;
      114466: inst = 32'h38632800;
      114467: inst = 32'h38842800;
      114468: inst = 32'h10a00001;
      114469: inst = 32'hca0bf29;
      114470: inst = 32'h13e00001;
      114471: inst = 32'hfe0d96a;
      114472: inst = 32'h5be00000;
      114473: inst = 32'h8c50000;
      114474: inst = 32'h24612800;
      114475: inst = 32'h10a00000;
      114476: inst = 32'hca0001b;
      114477: inst = 32'h24822800;
      114478: inst = 32'h10a00000;
      114479: inst = 32'hca00004;
      114480: inst = 32'h38632800;
      114481: inst = 32'h38842800;
      114482: inst = 32'h10a00001;
      114483: inst = 32'hca0bf37;
      114484: inst = 32'h13e00001;
      114485: inst = 32'hfe0d96a;
      114486: inst = 32'h5be00000;
      114487: inst = 32'h8c50000;
      114488: inst = 32'h24612800;
      114489: inst = 32'h10a00000;
      114490: inst = 32'hca0001b;
      114491: inst = 32'h24822800;
      114492: inst = 32'h10a00000;
      114493: inst = 32'hca00004;
      114494: inst = 32'h38632800;
      114495: inst = 32'h38842800;
      114496: inst = 32'h10a00001;
      114497: inst = 32'hca0bf45;
      114498: inst = 32'h13e00001;
      114499: inst = 32'hfe0d96a;
      114500: inst = 32'h5be00000;
      114501: inst = 32'h8c50000;
      114502: inst = 32'h24612800;
      114503: inst = 32'h10a00000;
      114504: inst = 32'hca0001b;
      114505: inst = 32'h24822800;
      114506: inst = 32'h10a00000;
      114507: inst = 32'hca00004;
      114508: inst = 32'h38632800;
      114509: inst = 32'h38842800;
      114510: inst = 32'h10a00001;
      114511: inst = 32'hca0bf53;
      114512: inst = 32'h13e00001;
      114513: inst = 32'hfe0d96a;
      114514: inst = 32'h5be00000;
      114515: inst = 32'h8c50000;
      114516: inst = 32'h24612800;
      114517: inst = 32'h10a00000;
      114518: inst = 32'hca0001b;
      114519: inst = 32'h24822800;
      114520: inst = 32'h10a00000;
      114521: inst = 32'hca00004;
      114522: inst = 32'h38632800;
      114523: inst = 32'h38842800;
      114524: inst = 32'h10a00001;
      114525: inst = 32'hca0bf61;
      114526: inst = 32'h13e00001;
      114527: inst = 32'hfe0d96a;
      114528: inst = 32'h5be00000;
      114529: inst = 32'h8c50000;
      114530: inst = 32'h24612800;
      114531: inst = 32'h10a00000;
      114532: inst = 32'hca0001b;
      114533: inst = 32'h24822800;
      114534: inst = 32'h10a00000;
      114535: inst = 32'hca00004;
      114536: inst = 32'h38632800;
      114537: inst = 32'h38842800;
      114538: inst = 32'h10a00001;
      114539: inst = 32'hca0bf6f;
      114540: inst = 32'h13e00001;
      114541: inst = 32'hfe0d96a;
      114542: inst = 32'h5be00000;
      114543: inst = 32'h8c50000;
      114544: inst = 32'h24612800;
      114545: inst = 32'h10a00000;
      114546: inst = 32'hca0001b;
      114547: inst = 32'h24822800;
      114548: inst = 32'h10a00000;
      114549: inst = 32'hca00004;
      114550: inst = 32'h38632800;
      114551: inst = 32'h38842800;
      114552: inst = 32'h10a00001;
      114553: inst = 32'hca0bf7d;
      114554: inst = 32'h13e00001;
      114555: inst = 32'hfe0d96a;
      114556: inst = 32'h5be00000;
      114557: inst = 32'h8c50000;
      114558: inst = 32'h24612800;
      114559: inst = 32'h10a00000;
      114560: inst = 32'hca0001b;
      114561: inst = 32'h24822800;
      114562: inst = 32'h10a00000;
      114563: inst = 32'hca00004;
      114564: inst = 32'h38632800;
      114565: inst = 32'h38842800;
      114566: inst = 32'h10a00001;
      114567: inst = 32'hca0bf8b;
      114568: inst = 32'h13e00001;
      114569: inst = 32'hfe0d96a;
      114570: inst = 32'h5be00000;
      114571: inst = 32'h8c50000;
      114572: inst = 32'h24612800;
      114573: inst = 32'h10a00000;
      114574: inst = 32'hca0001b;
      114575: inst = 32'h24822800;
      114576: inst = 32'h10a00000;
      114577: inst = 32'hca00004;
      114578: inst = 32'h38632800;
      114579: inst = 32'h38842800;
      114580: inst = 32'h10a00001;
      114581: inst = 32'hca0bf99;
      114582: inst = 32'h13e00001;
      114583: inst = 32'hfe0d96a;
      114584: inst = 32'h5be00000;
      114585: inst = 32'h8c50000;
      114586: inst = 32'h24612800;
      114587: inst = 32'h10a00000;
      114588: inst = 32'hca0001b;
      114589: inst = 32'h24822800;
      114590: inst = 32'h10a00000;
      114591: inst = 32'hca00004;
      114592: inst = 32'h38632800;
      114593: inst = 32'h38842800;
      114594: inst = 32'h10a00001;
      114595: inst = 32'hca0bfa7;
      114596: inst = 32'h13e00001;
      114597: inst = 32'hfe0d96a;
      114598: inst = 32'h5be00000;
      114599: inst = 32'h8c50000;
      114600: inst = 32'h24612800;
      114601: inst = 32'h10a00000;
      114602: inst = 32'hca0001b;
      114603: inst = 32'h24822800;
      114604: inst = 32'h10a00000;
      114605: inst = 32'hca00004;
      114606: inst = 32'h38632800;
      114607: inst = 32'h38842800;
      114608: inst = 32'h10a00001;
      114609: inst = 32'hca0bfb5;
      114610: inst = 32'h13e00001;
      114611: inst = 32'hfe0d96a;
      114612: inst = 32'h5be00000;
      114613: inst = 32'h8c50000;
      114614: inst = 32'h24612800;
      114615: inst = 32'h10a00000;
      114616: inst = 32'hca0001b;
      114617: inst = 32'h24822800;
      114618: inst = 32'h10a00000;
      114619: inst = 32'hca00004;
      114620: inst = 32'h38632800;
      114621: inst = 32'h38842800;
      114622: inst = 32'h10a00001;
      114623: inst = 32'hca0bfc3;
      114624: inst = 32'h13e00001;
      114625: inst = 32'hfe0d96a;
      114626: inst = 32'h5be00000;
      114627: inst = 32'h8c50000;
      114628: inst = 32'h24612800;
      114629: inst = 32'h10a00000;
      114630: inst = 32'hca0001b;
      114631: inst = 32'h24822800;
      114632: inst = 32'h10a00000;
      114633: inst = 32'hca00004;
      114634: inst = 32'h38632800;
      114635: inst = 32'h38842800;
      114636: inst = 32'h10a00001;
      114637: inst = 32'hca0bfd1;
      114638: inst = 32'h13e00001;
      114639: inst = 32'hfe0d96a;
      114640: inst = 32'h5be00000;
      114641: inst = 32'h8c50000;
      114642: inst = 32'h24612800;
      114643: inst = 32'h10a00000;
      114644: inst = 32'hca0001b;
      114645: inst = 32'h24822800;
      114646: inst = 32'h10a00000;
      114647: inst = 32'hca00004;
      114648: inst = 32'h38632800;
      114649: inst = 32'h38842800;
      114650: inst = 32'h10a00001;
      114651: inst = 32'hca0bfdf;
      114652: inst = 32'h13e00001;
      114653: inst = 32'hfe0d96a;
      114654: inst = 32'h5be00000;
      114655: inst = 32'h8c50000;
      114656: inst = 32'h24612800;
      114657: inst = 32'h10a00000;
      114658: inst = 32'hca0001b;
      114659: inst = 32'h24822800;
      114660: inst = 32'h10a00000;
      114661: inst = 32'hca00004;
      114662: inst = 32'h38632800;
      114663: inst = 32'h38842800;
      114664: inst = 32'h10a00001;
      114665: inst = 32'hca0bfed;
      114666: inst = 32'h13e00001;
      114667: inst = 32'hfe0d96a;
      114668: inst = 32'h5be00000;
      114669: inst = 32'h8c50000;
      114670: inst = 32'h24612800;
      114671: inst = 32'h10a00000;
      114672: inst = 32'hca0001b;
      114673: inst = 32'h24822800;
      114674: inst = 32'h10a00000;
      114675: inst = 32'hca00004;
      114676: inst = 32'h38632800;
      114677: inst = 32'h38842800;
      114678: inst = 32'h10a00001;
      114679: inst = 32'hca0bffb;
      114680: inst = 32'h13e00001;
      114681: inst = 32'hfe0d96a;
      114682: inst = 32'h5be00000;
      114683: inst = 32'h8c50000;
      114684: inst = 32'h24612800;
      114685: inst = 32'h10a00000;
      114686: inst = 32'hca0001b;
      114687: inst = 32'h24822800;
      114688: inst = 32'h10a00000;
      114689: inst = 32'hca00004;
      114690: inst = 32'h38632800;
      114691: inst = 32'h38842800;
      114692: inst = 32'h10a00001;
      114693: inst = 32'hca0c009;
      114694: inst = 32'h13e00001;
      114695: inst = 32'hfe0d96a;
      114696: inst = 32'h5be00000;
      114697: inst = 32'h8c50000;
      114698: inst = 32'h24612800;
      114699: inst = 32'h10a00000;
      114700: inst = 32'hca0001b;
      114701: inst = 32'h24822800;
      114702: inst = 32'h10a00000;
      114703: inst = 32'hca00004;
      114704: inst = 32'h38632800;
      114705: inst = 32'h38842800;
      114706: inst = 32'h10a00001;
      114707: inst = 32'hca0c017;
      114708: inst = 32'h13e00001;
      114709: inst = 32'hfe0d96a;
      114710: inst = 32'h5be00000;
      114711: inst = 32'h8c50000;
      114712: inst = 32'h24612800;
      114713: inst = 32'h10a00000;
      114714: inst = 32'hca0001b;
      114715: inst = 32'h24822800;
      114716: inst = 32'h10a00000;
      114717: inst = 32'hca00004;
      114718: inst = 32'h38632800;
      114719: inst = 32'h38842800;
      114720: inst = 32'h10a00001;
      114721: inst = 32'hca0c025;
      114722: inst = 32'h13e00001;
      114723: inst = 32'hfe0d96a;
      114724: inst = 32'h5be00000;
      114725: inst = 32'h8c50000;
      114726: inst = 32'h24612800;
      114727: inst = 32'h10a00000;
      114728: inst = 32'hca0001b;
      114729: inst = 32'h24822800;
      114730: inst = 32'h10a00000;
      114731: inst = 32'hca00004;
      114732: inst = 32'h38632800;
      114733: inst = 32'h38842800;
      114734: inst = 32'h10a00001;
      114735: inst = 32'hca0c033;
      114736: inst = 32'h13e00001;
      114737: inst = 32'hfe0d96a;
      114738: inst = 32'h5be00000;
      114739: inst = 32'h8c50000;
      114740: inst = 32'h24612800;
      114741: inst = 32'h10a00000;
      114742: inst = 32'hca0001b;
      114743: inst = 32'h24822800;
      114744: inst = 32'h10a00000;
      114745: inst = 32'hca00004;
      114746: inst = 32'h38632800;
      114747: inst = 32'h38842800;
      114748: inst = 32'h10a00001;
      114749: inst = 32'hca0c041;
      114750: inst = 32'h13e00001;
      114751: inst = 32'hfe0d96a;
      114752: inst = 32'h5be00000;
      114753: inst = 32'h8c50000;
      114754: inst = 32'h24612800;
      114755: inst = 32'h10a00000;
      114756: inst = 32'hca0001b;
      114757: inst = 32'h24822800;
      114758: inst = 32'h10a00000;
      114759: inst = 32'hca00004;
      114760: inst = 32'h38632800;
      114761: inst = 32'h38842800;
      114762: inst = 32'h10a00001;
      114763: inst = 32'hca0c04f;
      114764: inst = 32'h13e00001;
      114765: inst = 32'hfe0d96a;
      114766: inst = 32'h5be00000;
      114767: inst = 32'h8c50000;
      114768: inst = 32'h24612800;
      114769: inst = 32'h10a00000;
      114770: inst = 32'hca0001b;
      114771: inst = 32'h24822800;
      114772: inst = 32'h10a00000;
      114773: inst = 32'hca00004;
      114774: inst = 32'h38632800;
      114775: inst = 32'h38842800;
      114776: inst = 32'h10a00001;
      114777: inst = 32'hca0c05d;
      114778: inst = 32'h13e00001;
      114779: inst = 32'hfe0d96a;
      114780: inst = 32'h5be00000;
      114781: inst = 32'h8c50000;
      114782: inst = 32'h24612800;
      114783: inst = 32'h10a00000;
      114784: inst = 32'hca0001b;
      114785: inst = 32'h24822800;
      114786: inst = 32'h10a00000;
      114787: inst = 32'hca00004;
      114788: inst = 32'h38632800;
      114789: inst = 32'h38842800;
      114790: inst = 32'h10a00001;
      114791: inst = 32'hca0c06b;
      114792: inst = 32'h13e00001;
      114793: inst = 32'hfe0d96a;
      114794: inst = 32'h5be00000;
      114795: inst = 32'h8c50000;
      114796: inst = 32'h24612800;
      114797: inst = 32'h10a00000;
      114798: inst = 32'hca0001b;
      114799: inst = 32'h24822800;
      114800: inst = 32'h10a00000;
      114801: inst = 32'hca00004;
      114802: inst = 32'h38632800;
      114803: inst = 32'h38842800;
      114804: inst = 32'h10a00001;
      114805: inst = 32'hca0c079;
      114806: inst = 32'h13e00001;
      114807: inst = 32'hfe0d96a;
      114808: inst = 32'h5be00000;
      114809: inst = 32'h8c50000;
      114810: inst = 32'h24612800;
      114811: inst = 32'h10a00000;
      114812: inst = 32'hca0001b;
      114813: inst = 32'h24822800;
      114814: inst = 32'h10a00000;
      114815: inst = 32'hca00004;
      114816: inst = 32'h38632800;
      114817: inst = 32'h38842800;
      114818: inst = 32'h10a00001;
      114819: inst = 32'hca0c087;
      114820: inst = 32'h13e00001;
      114821: inst = 32'hfe0d96a;
      114822: inst = 32'h5be00000;
      114823: inst = 32'h8c50000;
      114824: inst = 32'h24612800;
      114825: inst = 32'h10a00000;
      114826: inst = 32'hca0001b;
      114827: inst = 32'h24822800;
      114828: inst = 32'h10a00000;
      114829: inst = 32'hca00004;
      114830: inst = 32'h38632800;
      114831: inst = 32'h38842800;
      114832: inst = 32'h10a00001;
      114833: inst = 32'hca0c095;
      114834: inst = 32'h13e00001;
      114835: inst = 32'hfe0d96a;
      114836: inst = 32'h5be00000;
      114837: inst = 32'h8c50000;
      114838: inst = 32'h24612800;
      114839: inst = 32'h10a00000;
      114840: inst = 32'hca0001b;
      114841: inst = 32'h24822800;
      114842: inst = 32'h10a00000;
      114843: inst = 32'hca00004;
      114844: inst = 32'h38632800;
      114845: inst = 32'h38842800;
      114846: inst = 32'h10a00001;
      114847: inst = 32'hca0c0a3;
      114848: inst = 32'h13e00001;
      114849: inst = 32'hfe0d96a;
      114850: inst = 32'h5be00000;
      114851: inst = 32'h8c50000;
      114852: inst = 32'h24612800;
      114853: inst = 32'h10a00000;
      114854: inst = 32'hca0001b;
      114855: inst = 32'h24822800;
      114856: inst = 32'h10a00000;
      114857: inst = 32'hca00004;
      114858: inst = 32'h38632800;
      114859: inst = 32'h38842800;
      114860: inst = 32'h10a00001;
      114861: inst = 32'hca0c0b1;
      114862: inst = 32'h13e00001;
      114863: inst = 32'hfe0d96a;
      114864: inst = 32'h5be00000;
      114865: inst = 32'h8c50000;
      114866: inst = 32'h24612800;
      114867: inst = 32'h10a00000;
      114868: inst = 32'hca0001b;
      114869: inst = 32'h24822800;
      114870: inst = 32'h10a00000;
      114871: inst = 32'hca00004;
      114872: inst = 32'h38632800;
      114873: inst = 32'h38842800;
      114874: inst = 32'h10a00001;
      114875: inst = 32'hca0c0bf;
      114876: inst = 32'h13e00001;
      114877: inst = 32'hfe0d96a;
      114878: inst = 32'h5be00000;
      114879: inst = 32'h8c50000;
      114880: inst = 32'h24612800;
      114881: inst = 32'h10a00000;
      114882: inst = 32'hca0001b;
      114883: inst = 32'h24822800;
      114884: inst = 32'h10a00000;
      114885: inst = 32'hca00004;
      114886: inst = 32'h38632800;
      114887: inst = 32'h38842800;
      114888: inst = 32'h10a00001;
      114889: inst = 32'hca0c0cd;
      114890: inst = 32'h13e00001;
      114891: inst = 32'hfe0d96a;
      114892: inst = 32'h5be00000;
      114893: inst = 32'h8c50000;
      114894: inst = 32'h24612800;
      114895: inst = 32'h10a00000;
      114896: inst = 32'hca0001b;
      114897: inst = 32'h24822800;
      114898: inst = 32'h10a00000;
      114899: inst = 32'hca00004;
      114900: inst = 32'h38632800;
      114901: inst = 32'h38842800;
      114902: inst = 32'h10a00001;
      114903: inst = 32'hca0c0db;
      114904: inst = 32'h13e00001;
      114905: inst = 32'hfe0d96a;
      114906: inst = 32'h5be00000;
      114907: inst = 32'h8c50000;
      114908: inst = 32'h24612800;
      114909: inst = 32'h10a00000;
      114910: inst = 32'hca0001b;
      114911: inst = 32'h24822800;
      114912: inst = 32'h10a00000;
      114913: inst = 32'hca00004;
      114914: inst = 32'h38632800;
      114915: inst = 32'h38842800;
      114916: inst = 32'h10a00001;
      114917: inst = 32'hca0c0e9;
      114918: inst = 32'h13e00001;
      114919: inst = 32'hfe0d96a;
      114920: inst = 32'h5be00000;
      114921: inst = 32'h8c50000;
      114922: inst = 32'h24612800;
      114923: inst = 32'h10a00000;
      114924: inst = 32'hca0001b;
      114925: inst = 32'h24822800;
      114926: inst = 32'h10a00000;
      114927: inst = 32'hca00004;
      114928: inst = 32'h38632800;
      114929: inst = 32'h38842800;
      114930: inst = 32'h10a00001;
      114931: inst = 32'hca0c0f7;
      114932: inst = 32'h13e00001;
      114933: inst = 32'hfe0d96a;
      114934: inst = 32'h5be00000;
      114935: inst = 32'h8c50000;
      114936: inst = 32'h24612800;
      114937: inst = 32'h10a00000;
      114938: inst = 32'hca0001b;
      114939: inst = 32'h24822800;
      114940: inst = 32'h10a00000;
      114941: inst = 32'hca00004;
      114942: inst = 32'h38632800;
      114943: inst = 32'h38842800;
      114944: inst = 32'h10a00001;
      114945: inst = 32'hca0c105;
      114946: inst = 32'h13e00001;
      114947: inst = 32'hfe0d96a;
      114948: inst = 32'h5be00000;
      114949: inst = 32'h8c50000;
      114950: inst = 32'h24612800;
      114951: inst = 32'h10a00000;
      114952: inst = 32'hca0001b;
      114953: inst = 32'h24822800;
      114954: inst = 32'h10a00000;
      114955: inst = 32'hca00004;
      114956: inst = 32'h38632800;
      114957: inst = 32'h38842800;
      114958: inst = 32'h10a00001;
      114959: inst = 32'hca0c113;
      114960: inst = 32'h13e00001;
      114961: inst = 32'hfe0d96a;
      114962: inst = 32'h5be00000;
      114963: inst = 32'h8c50000;
      114964: inst = 32'h24612800;
      114965: inst = 32'h10a00000;
      114966: inst = 32'hca0001b;
      114967: inst = 32'h24822800;
      114968: inst = 32'h10a00000;
      114969: inst = 32'hca00004;
      114970: inst = 32'h38632800;
      114971: inst = 32'h38842800;
      114972: inst = 32'h10a00001;
      114973: inst = 32'hca0c121;
      114974: inst = 32'h13e00001;
      114975: inst = 32'hfe0d96a;
      114976: inst = 32'h5be00000;
      114977: inst = 32'h8c50000;
      114978: inst = 32'h24612800;
      114979: inst = 32'h10a00000;
      114980: inst = 32'hca0001b;
      114981: inst = 32'h24822800;
      114982: inst = 32'h10a00000;
      114983: inst = 32'hca00004;
      114984: inst = 32'h38632800;
      114985: inst = 32'h38842800;
      114986: inst = 32'h10a00001;
      114987: inst = 32'hca0c12f;
      114988: inst = 32'h13e00001;
      114989: inst = 32'hfe0d96a;
      114990: inst = 32'h5be00000;
      114991: inst = 32'h8c50000;
      114992: inst = 32'h24612800;
      114993: inst = 32'h10a00000;
      114994: inst = 32'hca0001b;
      114995: inst = 32'h24822800;
      114996: inst = 32'h10a00000;
      114997: inst = 32'hca00004;
      114998: inst = 32'h38632800;
      114999: inst = 32'h38842800;
      115000: inst = 32'h10a00001;
      115001: inst = 32'hca0c13d;
      115002: inst = 32'h13e00001;
      115003: inst = 32'hfe0d96a;
      115004: inst = 32'h5be00000;
      115005: inst = 32'h8c50000;
      115006: inst = 32'h24612800;
      115007: inst = 32'h10a00000;
      115008: inst = 32'hca0001b;
      115009: inst = 32'h24822800;
      115010: inst = 32'h10a00000;
      115011: inst = 32'hca00004;
      115012: inst = 32'h38632800;
      115013: inst = 32'h38842800;
      115014: inst = 32'h10a00001;
      115015: inst = 32'hca0c14b;
      115016: inst = 32'h13e00001;
      115017: inst = 32'hfe0d96a;
      115018: inst = 32'h5be00000;
      115019: inst = 32'h8c50000;
      115020: inst = 32'h24612800;
      115021: inst = 32'h10a00000;
      115022: inst = 32'hca0001b;
      115023: inst = 32'h24822800;
      115024: inst = 32'h10a00000;
      115025: inst = 32'hca00004;
      115026: inst = 32'h38632800;
      115027: inst = 32'h38842800;
      115028: inst = 32'h10a00001;
      115029: inst = 32'hca0c159;
      115030: inst = 32'h13e00001;
      115031: inst = 32'hfe0d96a;
      115032: inst = 32'h5be00000;
      115033: inst = 32'h8c50000;
      115034: inst = 32'h24612800;
      115035: inst = 32'h10a00000;
      115036: inst = 32'hca0001b;
      115037: inst = 32'h24822800;
      115038: inst = 32'h10a00000;
      115039: inst = 32'hca00004;
      115040: inst = 32'h38632800;
      115041: inst = 32'h38842800;
      115042: inst = 32'h10a00001;
      115043: inst = 32'hca0c167;
      115044: inst = 32'h13e00001;
      115045: inst = 32'hfe0d96a;
      115046: inst = 32'h5be00000;
      115047: inst = 32'h8c50000;
      115048: inst = 32'h24612800;
      115049: inst = 32'h10a00000;
      115050: inst = 32'hca0001b;
      115051: inst = 32'h24822800;
      115052: inst = 32'h10a00000;
      115053: inst = 32'hca00004;
      115054: inst = 32'h38632800;
      115055: inst = 32'h38842800;
      115056: inst = 32'h10a00001;
      115057: inst = 32'hca0c175;
      115058: inst = 32'h13e00001;
      115059: inst = 32'hfe0d96a;
      115060: inst = 32'h5be00000;
      115061: inst = 32'h8c50000;
      115062: inst = 32'h24612800;
      115063: inst = 32'h10a00000;
      115064: inst = 32'hca0001b;
      115065: inst = 32'h24822800;
      115066: inst = 32'h10a00000;
      115067: inst = 32'hca00004;
      115068: inst = 32'h38632800;
      115069: inst = 32'h38842800;
      115070: inst = 32'h10a00001;
      115071: inst = 32'hca0c183;
      115072: inst = 32'h13e00001;
      115073: inst = 32'hfe0d96a;
      115074: inst = 32'h5be00000;
      115075: inst = 32'h8c50000;
      115076: inst = 32'h24612800;
      115077: inst = 32'h10a00000;
      115078: inst = 32'hca0001b;
      115079: inst = 32'h24822800;
      115080: inst = 32'h10a00000;
      115081: inst = 32'hca00004;
      115082: inst = 32'h38632800;
      115083: inst = 32'h38842800;
      115084: inst = 32'h10a00001;
      115085: inst = 32'hca0c191;
      115086: inst = 32'h13e00001;
      115087: inst = 32'hfe0d96a;
      115088: inst = 32'h5be00000;
      115089: inst = 32'h8c50000;
      115090: inst = 32'h24612800;
      115091: inst = 32'h10a00000;
      115092: inst = 32'hca0001b;
      115093: inst = 32'h24822800;
      115094: inst = 32'h10a00000;
      115095: inst = 32'hca00004;
      115096: inst = 32'h38632800;
      115097: inst = 32'h38842800;
      115098: inst = 32'h10a00001;
      115099: inst = 32'hca0c19f;
      115100: inst = 32'h13e00001;
      115101: inst = 32'hfe0d96a;
      115102: inst = 32'h5be00000;
      115103: inst = 32'h8c50000;
      115104: inst = 32'h24612800;
      115105: inst = 32'h10a00000;
      115106: inst = 32'hca0001b;
      115107: inst = 32'h24822800;
      115108: inst = 32'h10a00000;
      115109: inst = 32'hca00004;
      115110: inst = 32'h38632800;
      115111: inst = 32'h38842800;
      115112: inst = 32'h10a00001;
      115113: inst = 32'hca0c1ad;
      115114: inst = 32'h13e00001;
      115115: inst = 32'hfe0d96a;
      115116: inst = 32'h5be00000;
      115117: inst = 32'h8c50000;
      115118: inst = 32'h24612800;
      115119: inst = 32'h10a00000;
      115120: inst = 32'hca0001b;
      115121: inst = 32'h24822800;
      115122: inst = 32'h10a00000;
      115123: inst = 32'hca00004;
      115124: inst = 32'h38632800;
      115125: inst = 32'h38842800;
      115126: inst = 32'h10a00001;
      115127: inst = 32'hca0c1bb;
      115128: inst = 32'h13e00001;
      115129: inst = 32'hfe0d96a;
      115130: inst = 32'h5be00000;
      115131: inst = 32'h8c50000;
      115132: inst = 32'h24612800;
      115133: inst = 32'h10a00000;
      115134: inst = 32'hca0001b;
      115135: inst = 32'h24822800;
      115136: inst = 32'h10a00000;
      115137: inst = 32'hca00004;
      115138: inst = 32'h38632800;
      115139: inst = 32'h38842800;
      115140: inst = 32'h10a00001;
      115141: inst = 32'hca0c1c9;
      115142: inst = 32'h13e00001;
      115143: inst = 32'hfe0d96a;
      115144: inst = 32'h5be00000;
      115145: inst = 32'h8c50000;
      115146: inst = 32'h24612800;
      115147: inst = 32'h10a00000;
      115148: inst = 32'hca0001b;
      115149: inst = 32'h24822800;
      115150: inst = 32'h10a00000;
      115151: inst = 32'hca00004;
      115152: inst = 32'h38632800;
      115153: inst = 32'h38842800;
      115154: inst = 32'h10a00001;
      115155: inst = 32'hca0c1d7;
      115156: inst = 32'h13e00001;
      115157: inst = 32'hfe0d96a;
      115158: inst = 32'h5be00000;
      115159: inst = 32'h8c50000;
      115160: inst = 32'h24612800;
      115161: inst = 32'h10a00000;
      115162: inst = 32'hca0001b;
      115163: inst = 32'h24822800;
      115164: inst = 32'h10a00000;
      115165: inst = 32'hca00004;
      115166: inst = 32'h38632800;
      115167: inst = 32'h38842800;
      115168: inst = 32'h10a00001;
      115169: inst = 32'hca0c1e5;
      115170: inst = 32'h13e00001;
      115171: inst = 32'hfe0d96a;
      115172: inst = 32'h5be00000;
      115173: inst = 32'h8c50000;
      115174: inst = 32'h24612800;
      115175: inst = 32'h10a00000;
      115176: inst = 32'hca0001b;
      115177: inst = 32'h24822800;
      115178: inst = 32'h10a00000;
      115179: inst = 32'hca00004;
      115180: inst = 32'h38632800;
      115181: inst = 32'h38842800;
      115182: inst = 32'h10a00001;
      115183: inst = 32'hca0c1f3;
      115184: inst = 32'h13e00001;
      115185: inst = 32'hfe0d96a;
      115186: inst = 32'h5be00000;
      115187: inst = 32'h8c50000;
      115188: inst = 32'h24612800;
      115189: inst = 32'h10a00000;
      115190: inst = 32'hca0001b;
      115191: inst = 32'h24822800;
      115192: inst = 32'h10a00000;
      115193: inst = 32'hca00004;
      115194: inst = 32'h38632800;
      115195: inst = 32'h38842800;
      115196: inst = 32'h10a00001;
      115197: inst = 32'hca0c201;
      115198: inst = 32'h13e00001;
      115199: inst = 32'hfe0d96a;
      115200: inst = 32'h5be00000;
      115201: inst = 32'h8c50000;
      115202: inst = 32'h24612800;
      115203: inst = 32'h10a00000;
      115204: inst = 32'hca0001b;
      115205: inst = 32'h24822800;
      115206: inst = 32'h10a00000;
      115207: inst = 32'hca00004;
      115208: inst = 32'h38632800;
      115209: inst = 32'h38842800;
      115210: inst = 32'h10a00001;
      115211: inst = 32'hca0c20f;
      115212: inst = 32'h13e00001;
      115213: inst = 32'hfe0d96a;
      115214: inst = 32'h5be00000;
      115215: inst = 32'h8c50000;
      115216: inst = 32'h24612800;
      115217: inst = 32'h10a00000;
      115218: inst = 32'hca0001b;
      115219: inst = 32'h24822800;
      115220: inst = 32'h10a00000;
      115221: inst = 32'hca00004;
      115222: inst = 32'h38632800;
      115223: inst = 32'h38842800;
      115224: inst = 32'h10a00001;
      115225: inst = 32'hca0c21d;
      115226: inst = 32'h13e00001;
      115227: inst = 32'hfe0d96a;
      115228: inst = 32'h5be00000;
      115229: inst = 32'h8c50000;
      115230: inst = 32'h24612800;
      115231: inst = 32'h10a00000;
      115232: inst = 32'hca0001b;
      115233: inst = 32'h24822800;
      115234: inst = 32'h10a00000;
      115235: inst = 32'hca00004;
      115236: inst = 32'h38632800;
      115237: inst = 32'h38842800;
      115238: inst = 32'h10a00001;
      115239: inst = 32'hca0c22b;
      115240: inst = 32'h13e00001;
      115241: inst = 32'hfe0d96a;
      115242: inst = 32'h5be00000;
      115243: inst = 32'h8c50000;
      115244: inst = 32'h24612800;
      115245: inst = 32'h10a00000;
      115246: inst = 32'hca0001b;
      115247: inst = 32'h24822800;
      115248: inst = 32'h10a00000;
      115249: inst = 32'hca00004;
      115250: inst = 32'h38632800;
      115251: inst = 32'h38842800;
      115252: inst = 32'h10a00001;
      115253: inst = 32'hca0c239;
      115254: inst = 32'h13e00001;
      115255: inst = 32'hfe0d96a;
      115256: inst = 32'h5be00000;
      115257: inst = 32'h8c50000;
      115258: inst = 32'h24612800;
      115259: inst = 32'h10a00000;
      115260: inst = 32'hca0001b;
      115261: inst = 32'h24822800;
      115262: inst = 32'h10a00000;
      115263: inst = 32'hca00004;
      115264: inst = 32'h38632800;
      115265: inst = 32'h38842800;
      115266: inst = 32'h10a00001;
      115267: inst = 32'hca0c247;
      115268: inst = 32'h13e00001;
      115269: inst = 32'hfe0d96a;
      115270: inst = 32'h5be00000;
      115271: inst = 32'h8c50000;
      115272: inst = 32'h24612800;
      115273: inst = 32'h10a00000;
      115274: inst = 32'hca0001b;
      115275: inst = 32'h24822800;
      115276: inst = 32'h10a00000;
      115277: inst = 32'hca00004;
      115278: inst = 32'h38632800;
      115279: inst = 32'h38842800;
      115280: inst = 32'h10a00001;
      115281: inst = 32'hca0c255;
      115282: inst = 32'h13e00001;
      115283: inst = 32'hfe0d96a;
      115284: inst = 32'h5be00000;
      115285: inst = 32'h8c50000;
      115286: inst = 32'h24612800;
      115287: inst = 32'h10a00000;
      115288: inst = 32'hca0001b;
      115289: inst = 32'h24822800;
      115290: inst = 32'h10a00000;
      115291: inst = 32'hca00004;
      115292: inst = 32'h38632800;
      115293: inst = 32'h38842800;
      115294: inst = 32'h10a00001;
      115295: inst = 32'hca0c263;
      115296: inst = 32'h13e00001;
      115297: inst = 32'hfe0d96a;
      115298: inst = 32'h5be00000;
      115299: inst = 32'h8c50000;
      115300: inst = 32'h24612800;
      115301: inst = 32'h10a00000;
      115302: inst = 32'hca0001b;
      115303: inst = 32'h24822800;
      115304: inst = 32'h10a00000;
      115305: inst = 32'hca00004;
      115306: inst = 32'h38632800;
      115307: inst = 32'h38842800;
      115308: inst = 32'h10a00001;
      115309: inst = 32'hca0c271;
      115310: inst = 32'h13e00001;
      115311: inst = 32'hfe0d96a;
      115312: inst = 32'h5be00000;
      115313: inst = 32'h8c50000;
      115314: inst = 32'h24612800;
      115315: inst = 32'h10a00000;
      115316: inst = 32'hca0001b;
      115317: inst = 32'h24822800;
      115318: inst = 32'h10a00000;
      115319: inst = 32'hca00004;
      115320: inst = 32'h38632800;
      115321: inst = 32'h38842800;
      115322: inst = 32'h10a00001;
      115323: inst = 32'hca0c27f;
      115324: inst = 32'h13e00001;
      115325: inst = 32'hfe0d96a;
      115326: inst = 32'h5be00000;
      115327: inst = 32'h8c50000;
      115328: inst = 32'h24612800;
      115329: inst = 32'h10a00000;
      115330: inst = 32'hca0001b;
      115331: inst = 32'h24822800;
      115332: inst = 32'h10a00000;
      115333: inst = 32'hca00004;
      115334: inst = 32'h38632800;
      115335: inst = 32'h38842800;
      115336: inst = 32'h10a00001;
      115337: inst = 32'hca0c28d;
      115338: inst = 32'h13e00001;
      115339: inst = 32'hfe0d96a;
      115340: inst = 32'h5be00000;
      115341: inst = 32'h8c50000;
      115342: inst = 32'h24612800;
      115343: inst = 32'h10a00000;
      115344: inst = 32'hca0001b;
      115345: inst = 32'h24822800;
      115346: inst = 32'h10a00000;
      115347: inst = 32'hca00004;
      115348: inst = 32'h38632800;
      115349: inst = 32'h38842800;
      115350: inst = 32'h10a00001;
      115351: inst = 32'hca0c29b;
      115352: inst = 32'h13e00001;
      115353: inst = 32'hfe0d96a;
      115354: inst = 32'h5be00000;
      115355: inst = 32'h8c50000;
      115356: inst = 32'h24612800;
      115357: inst = 32'h10a00000;
      115358: inst = 32'hca0001b;
      115359: inst = 32'h24822800;
      115360: inst = 32'h10a00000;
      115361: inst = 32'hca00004;
      115362: inst = 32'h38632800;
      115363: inst = 32'h38842800;
      115364: inst = 32'h10a00001;
      115365: inst = 32'hca0c2a9;
      115366: inst = 32'h13e00001;
      115367: inst = 32'hfe0d96a;
      115368: inst = 32'h5be00000;
      115369: inst = 32'h8c50000;
      115370: inst = 32'h24612800;
      115371: inst = 32'h10a00000;
      115372: inst = 32'hca0001b;
      115373: inst = 32'h24822800;
      115374: inst = 32'h10a00000;
      115375: inst = 32'hca00004;
      115376: inst = 32'h38632800;
      115377: inst = 32'h38842800;
      115378: inst = 32'h10a00001;
      115379: inst = 32'hca0c2b7;
      115380: inst = 32'h13e00001;
      115381: inst = 32'hfe0d96a;
      115382: inst = 32'h5be00000;
      115383: inst = 32'h8c50000;
      115384: inst = 32'h24612800;
      115385: inst = 32'h10a00000;
      115386: inst = 32'hca0001b;
      115387: inst = 32'h24822800;
      115388: inst = 32'h10a00000;
      115389: inst = 32'hca00004;
      115390: inst = 32'h38632800;
      115391: inst = 32'h38842800;
      115392: inst = 32'h10a00001;
      115393: inst = 32'hca0c2c5;
      115394: inst = 32'h13e00001;
      115395: inst = 32'hfe0d96a;
      115396: inst = 32'h5be00000;
      115397: inst = 32'h8c50000;
      115398: inst = 32'h24612800;
      115399: inst = 32'h10a00000;
      115400: inst = 32'hca0001b;
      115401: inst = 32'h24822800;
      115402: inst = 32'h10a00000;
      115403: inst = 32'hca00004;
      115404: inst = 32'h38632800;
      115405: inst = 32'h38842800;
      115406: inst = 32'h10a00001;
      115407: inst = 32'hca0c2d3;
      115408: inst = 32'h13e00001;
      115409: inst = 32'hfe0d96a;
      115410: inst = 32'h5be00000;
      115411: inst = 32'h8c50000;
      115412: inst = 32'h24612800;
      115413: inst = 32'h10a00000;
      115414: inst = 32'hca0001b;
      115415: inst = 32'h24822800;
      115416: inst = 32'h10a00000;
      115417: inst = 32'hca00004;
      115418: inst = 32'h38632800;
      115419: inst = 32'h38842800;
      115420: inst = 32'h10a00001;
      115421: inst = 32'hca0c2e1;
      115422: inst = 32'h13e00001;
      115423: inst = 32'hfe0d96a;
      115424: inst = 32'h5be00000;
      115425: inst = 32'h8c50000;
      115426: inst = 32'h24612800;
      115427: inst = 32'h10a00000;
      115428: inst = 32'hca0001b;
      115429: inst = 32'h24822800;
      115430: inst = 32'h10a00000;
      115431: inst = 32'hca00004;
      115432: inst = 32'h38632800;
      115433: inst = 32'h38842800;
      115434: inst = 32'h10a00001;
      115435: inst = 32'hca0c2ef;
      115436: inst = 32'h13e00001;
      115437: inst = 32'hfe0d96a;
      115438: inst = 32'h5be00000;
      115439: inst = 32'h8c50000;
      115440: inst = 32'h24612800;
      115441: inst = 32'h10a00000;
      115442: inst = 32'hca0001b;
      115443: inst = 32'h24822800;
      115444: inst = 32'h10a00000;
      115445: inst = 32'hca00004;
      115446: inst = 32'h38632800;
      115447: inst = 32'h38842800;
      115448: inst = 32'h10a00001;
      115449: inst = 32'hca0c2fd;
      115450: inst = 32'h13e00001;
      115451: inst = 32'hfe0d96a;
      115452: inst = 32'h5be00000;
      115453: inst = 32'h8c50000;
      115454: inst = 32'h24612800;
      115455: inst = 32'h10a00000;
      115456: inst = 32'hca0001b;
      115457: inst = 32'h24822800;
      115458: inst = 32'h10a00000;
      115459: inst = 32'hca00004;
      115460: inst = 32'h38632800;
      115461: inst = 32'h38842800;
      115462: inst = 32'h10a00001;
      115463: inst = 32'hca0c30b;
      115464: inst = 32'h13e00001;
      115465: inst = 32'hfe0d96a;
      115466: inst = 32'h5be00000;
      115467: inst = 32'h8c50000;
      115468: inst = 32'h24612800;
      115469: inst = 32'h10a00000;
      115470: inst = 32'hca0001b;
      115471: inst = 32'h24822800;
      115472: inst = 32'h10a00000;
      115473: inst = 32'hca00004;
      115474: inst = 32'h38632800;
      115475: inst = 32'h38842800;
      115476: inst = 32'h10a00001;
      115477: inst = 32'hca0c319;
      115478: inst = 32'h13e00001;
      115479: inst = 32'hfe0d96a;
      115480: inst = 32'h5be00000;
      115481: inst = 32'h8c50000;
      115482: inst = 32'h24612800;
      115483: inst = 32'h10a00000;
      115484: inst = 32'hca0001b;
      115485: inst = 32'h24822800;
      115486: inst = 32'h10a00000;
      115487: inst = 32'hca00004;
      115488: inst = 32'h38632800;
      115489: inst = 32'h38842800;
      115490: inst = 32'h10a00001;
      115491: inst = 32'hca0c327;
      115492: inst = 32'h13e00001;
      115493: inst = 32'hfe0d96a;
      115494: inst = 32'h5be00000;
      115495: inst = 32'h8c50000;
      115496: inst = 32'h24612800;
      115497: inst = 32'h10a00000;
      115498: inst = 32'hca0001b;
      115499: inst = 32'h24822800;
      115500: inst = 32'h10a00000;
      115501: inst = 32'hca00004;
      115502: inst = 32'h38632800;
      115503: inst = 32'h38842800;
      115504: inst = 32'h10a00001;
      115505: inst = 32'hca0c335;
      115506: inst = 32'h13e00001;
      115507: inst = 32'hfe0d96a;
      115508: inst = 32'h5be00000;
      115509: inst = 32'h8c50000;
      115510: inst = 32'h24612800;
      115511: inst = 32'h10a00000;
      115512: inst = 32'hca0001b;
      115513: inst = 32'h24822800;
      115514: inst = 32'h10a00000;
      115515: inst = 32'hca00004;
      115516: inst = 32'h38632800;
      115517: inst = 32'h38842800;
      115518: inst = 32'h10a00001;
      115519: inst = 32'hca0c343;
      115520: inst = 32'h13e00001;
      115521: inst = 32'hfe0d96a;
      115522: inst = 32'h5be00000;
      115523: inst = 32'h8c50000;
      115524: inst = 32'h24612800;
      115525: inst = 32'h10a00000;
      115526: inst = 32'hca0001b;
      115527: inst = 32'h24822800;
      115528: inst = 32'h10a00000;
      115529: inst = 32'hca00004;
      115530: inst = 32'h38632800;
      115531: inst = 32'h38842800;
      115532: inst = 32'h10a00001;
      115533: inst = 32'hca0c351;
      115534: inst = 32'h13e00001;
      115535: inst = 32'hfe0d96a;
      115536: inst = 32'h5be00000;
      115537: inst = 32'h8c50000;
      115538: inst = 32'h24612800;
      115539: inst = 32'h10a00000;
      115540: inst = 32'hca0001b;
      115541: inst = 32'h24822800;
      115542: inst = 32'h10a00000;
      115543: inst = 32'hca00004;
      115544: inst = 32'h38632800;
      115545: inst = 32'h38842800;
      115546: inst = 32'h10a00001;
      115547: inst = 32'hca0c35f;
      115548: inst = 32'h13e00001;
      115549: inst = 32'hfe0d96a;
      115550: inst = 32'h5be00000;
      115551: inst = 32'h8c50000;
      115552: inst = 32'h24612800;
      115553: inst = 32'h10a00000;
      115554: inst = 32'hca0001b;
      115555: inst = 32'h24822800;
      115556: inst = 32'h10a00000;
      115557: inst = 32'hca00004;
      115558: inst = 32'h38632800;
      115559: inst = 32'h38842800;
      115560: inst = 32'h10a00001;
      115561: inst = 32'hca0c36d;
      115562: inst = 32'h13e00001;
      115563: inst = 32'hfe0d96a;
      115564: inst = 32'h5be00000;
      115565: inst = 32'h8c50000;
      115566: inst = 32'h24612800;
      115567: inst = 32'h10a00000;
      115568: inst = 32'hca0001b;
      115569: inst = 32'h24822800;
      115570: inst = 32'h10a00000;
      115571: inst = 32'hca00004;
      115572: inst = 32'h38632800;
      115573: inst = 32'h38842800;
      115574: inst = 32'h10a00001;
      115575: inst = 32'hca0c37b;
      115576: inst = 32'h13e00001;
      115577: inst = 32'hfe0d96a;
      115578: inst = 32'h5be00000;
      115579: inst = 32'h8c50000;
      115580: inst = 32'h24612800;
      115581: inst = 32'h10a00000;
      115582: inst = 32'hca0001b;
      115583: inst = 32'h24822800;
      115584: inst = 32'h10a00000;
      115585: inst = 32'hca00004;
      115586: inst = 32'h38632800;
      115587: inst = 32'h38842800;
      115588: inst = 32'h10a00001;
      115589: inst = 32'hca0c389;
      115590: inst = 32'h13e00001;
      115591: inst = 32'hfe0d96a;
      115592: inst = 32'h5be00000;
      115593: inst = 32'h8c50000;
      115594: inst = 32'h24612800;
      115595: inst = 32'h10a00000;
      115596: inst = 32'hca0001b;
      115597: inst = 32'h24822800;
      115598: inst = 32'h10a00000;
      115599: inst = 32'hca00004;
      115600: inst = 32'h38632800;
      115601: inst = 32'h38842800;
      115602: inst = 32'h10a00001;
      115603: inst = 32'hca0c397;
      115604: inst = 32'h13e00001;
      115605: inst = 32'hfe0d96a;
      115606: inst = 32'h5be00000;
      115607: inst = 32'h8c50000;
      115608: inst = 32'h24612800;
      115609: inst = 32'h10a00000;
      115610: inst = 32'hca0001b;
      115611: inst = 32'h24822800;
      115612: inst = 32'h10a00000;
      115613: inst = 32'hca00004;
      115614: inst = 32'h38632800;
      115615: inst = 32'h38842800;
      115616: inst = 32'h10a00001;
      115617: inst = 32'hca0c3a5;
      115618: inst = 32'h13e00001;
      115619: inst = 32'hfe0d96a;
      115620: inst = 32'h5be00000;
      115621: inst = 32'h8c50000;
      115622: inst = 32'h24612800;
      115623: inst = 32'h10a00000;
      115624: inst = 32'hca0001b;
      115625: inst = 32'h24822800;
      115626: inst = 32'h10a00000;
      115627: inst = 32'hca00004;
      115628: inst = 32'h38632800;
      115629: inst = 32'h38842800;
      115630: inst = 32'h10a00001;
      115631: inst = 32'hca0c3b3;
      115632: inst = 32'h13e00001;
      115633: inst = 32'hfe0d96a;
      115634: inst = 32'h5be00000;
      115635: inst = 32'h8c50000;
      115636: inst = 32'h24612800;
      115637: inst = 32'h10a00000;
      115638: inst = 32'hca0001b;
      115639: inst = 32'h24822800;
      115640: inst = 32'h10a00000;
      115641: inst = 32'hca00004;
      115642: inst = 32'h38632800;
      115643: inst = 32'h38842800;
      115644: inst = 32'h10a00001;
      115645: inst = 32'hca0c3c1;
      115646: inst = 32'h13e00001;
      115647: inst = 32'hfe0d96a;
      115648: inst = 32'h5be00000;
      115649: inst = 32'h8c50000;
      115650: inst = 32'h24612800;
      115651: inst = 32'h10a00000;
      115652: inst = 32'hca0001b;
      115653: inst = 32'h24822800;
      115654: inst = 32'h10a00000;
      115655: inst = 32'hca00004;
      115656: inst = 32'h38632800;
      115657: inst = 32'h38842800;
      115658: inst = 32'h10a00001;
      115659: inst = 32'hca0c3cf;
      115660: inst = 32'h13e00001;
      115661: inst = 32'hfe0d96a;
      115662: inst = 32'h5be00000;
      115663: inst = 32'h8c50000;
      115664: inst = 32'h24612800;
      115665: inst = 32'h10a00000;
      115666: inst = 32'hca0001b;
      115667: inst = 32'h24822800;
      115668: inst = 32'h10a00000;
      115669: inst = 32'hca00004;
      115670: inst = 32'h38632800;
      115671: inst = 32'h38842800;
      115672: inst = 32'h10a00001;
      115673: inst = 32'hca0c3dd;
      115674: inst = 32'h13e00001;
      115675: inst = 32'hfe0d96a;
      115676: inst = 32'h5be00000;
      115677: inst = 32'h8c50000;
      115678: inst = 32'h24612800;
      115679: inst = 32'h10a00000;
      115680: inst = 32'hca0001b;
      115681: inst = 32'h24822800;
      115682: inst = 32'h10a00000;
      115683: inst = 32'hca00004;
      115684: inst = 32'h38632800;
      115685: inst = 32'h38842800;
      115686: inst = 32'h10a00001;
      115687: inst = 32'hca0c3eb;
      115688: inst = 32'h13e00001;
      115689: inst = 32'hfe0d96a;
      115690: inst = 32'h5be00000;
      115691: inst = 32'h8c50000;
      115692: inst = 32'h24612800;
      115693: inst = 32'h10a00000;
      115694: inst = 32'hca0001b;
      115695: inst = 32'h24822800;
      115696: inst = 32'h10a00000;
      115697: inst = 32'hca00004;
      115698: inst = 32'h38632800;
      115699: inst = 32'h38842800;
      115700: inst = 32'h10a00001;
      115701: inst = 32'hca0c3f9;
      115702: inst = 32'h13e00001;
      115703: inst = 32'hfe0d96a;
      115704: inst = 32'h5be00000;
      115705: inst = 32'h8c50000;
      115706: inst = 32'h24612800;
      115707: inst = 32'h10a00000;
      115708: inst = 32'hca0001b;
      115709: inst = 32'h24822800;
      115710: inst = 32'h10a00000;
      115711: inst = 32'hca00004;
      115712: inst = 32'h38632800;
      115713: inst = 32'h38842800;
      115714: inst = 32'h10a00001;
      115715: inst = 32'hca0c407;
      115716: inst = 32'h13e00001;
      115717: inst = 32'hfe0d96a;
      115718: inst = 32'h5be00000;
      115719: inst = 32'h8c50000;
      115720: inst = 32'h24612800;
      115721: inst = 32'h10a00000;
      115722: inst = 32'hca0001b;
      115723: inst = 32'h24822800;
      115724: inst = 32'h10a00000;
      115725: inst = 32'hca00004;
      115726: inst = 32'h38632800;
      115727: inst = 32'h38842800;
      115728: inst = 32'h10a00001;
      115729: inst = 32'hca0c415;
      115730: inst = 32'h13e00001;
      115731: inst = 32'hfe0d96a;
      115732: inst = 32'h5be00000;
      115733: inst = 32'h8c50000;
      115734: inst = 32'h24612800;
      115735: inst = 32'h10a00000;
      115736: inst = 32'hca0001b;
      115737: inst = 32'h24822800;
      115738: inst = 32'h10a00000;
      115739: inst = 32'hca00004;
      115740: inst = 32'h38632800;
      115741: inst = 32'h38842800;
      115742: inst = 32'h10a00001;
      115743: inst = 32'hca0c423;
      115744: inst = 32'h13e00001;
      115745: inst = 32'hfe0d96a;
      115746: inst = 32'h5be00000;
      115747: inst = 32'h8c50000;
      115748: inst = 32'h24612800;
      115749: inst = 32'h10a00000;
      115750: inst = 32'hca0001b;
      115751: inst = 32'h24822800;
      115752: inst = 32'h10a00000;
      115753: inst = 32'hca00004;
      115754: inst = 32'h38632800;
      115755: inst = 32'h38842800;
      115756: inst = 32'h10a00001;
      115757: inst = 32'hca0c431;
      115758: inst = 32'h13e00001;
      115759: inst = 32'hfe0d96a;
      115760: inst = 32'h5be00000;
      115761: inst = 32'h8c50000;
      115762: inst = 32'h24612800;
      115763: inst = 32'h10a00000;
      115764: inst = 32'hca0001b;
      115765: inst = 32'h24822800;
      115766: inst = 32'h10a00000;
      115767: inst = 32'hca00004;
      115768: inst = 32'h38632800;
      115769: inst = 32'h38842800;
      115770: inst = 32'h10a00001;
      115771: inst = 32'hca0c43f;
      115772: inst = 32'h13e00001;
      115773: inst = 32'hfe0d96a;
      115774: inst = 32'h5be00000;
      115775: inst = 32'h8c50000;
      115776: inst = 32'h24612800;
      115777: inst = 32'h10a00000;
      115778: inst = 32'hca0001b;
      115779: inst = 32'h24822800;
      115780: inst = 32'h10a00000;
      115781: inst = 32'hca00004;
      115782: inst = 32'h38632800;
      115783: inst = 32'h38842800;
      115784: inst = 32'h10a00001;
      115785: inst = 32'hca0c44d;
      115786: inst = 32'h13e00001;
      115787: inst = 32'hfe0d96a;
      115788: inst = 32'h5be00000;
      115789: inst = 32'h8c50000;
      115790: inst = 32'h24612800;
      115791: inst = 32'h10a00000;
      115792: inst = 32'hca0001b;
      115793: inst = 32'h24822800;
      115794: inst = 32'h10a00000;
      115795: inst = 32'hca00004;
      115796: inst = 32'h38632800;
      115797: inst = 32'h38842800;
      115798: inst = 32'h10a00001;
      115799: inst = 32'hca0c45b;
      115800: inst = 32'h13e00001;
      115801: inst = 32'hfe0d96a;
      115802: inst = 32'h5be00000;
      115803: inst = 32'h8c50000;
      115804: inst = 32'h24612800;
      115805: inst = 32'h10a00000;
      115806: inst = 32'hca0001b;
      115807: inst = 32'h24822800;
      115808: inst = 32'h10a00000;
      115809: inst = 32'hca00004;
      115810: inst = 32'h38632800;
      115811: inst = 32'h38842800;
      115812: inst = 32'h10a00001;
      115813: inst = 32'hca0c469;
      115814: inst = 32'h13e00001;
      115815: inst = 32'hfe0d96a;
      115816: inst = 32'h5be00000;
      115817: inst = 32'h8c50000;
      115818: inst = 32'h24612800;
      115819: inst = 32'h10a00000;
      115820: inst = 32'hca0001c;
      115821: inst = 32'h24822800;
      115822: inst = 32'h10a00000;
      115823: inst = 32'hca00004;
      115824: inst = 32'h38632800;
      115825: inst = 32'h38842800;
      115826: inst = 32'h10a00001;
      115827: inst = 32'hca0c477;
      115828: inst = 32'h13e00001;
      115829: inst = 32'hfe0d96a;
      115830: inst = 32'h5be00000;
      115831: inst = 32'h8c50000;
      115832: inst = 32'h24612800;
      115833: inst = 32'h10a00000;
      115834: inst = 32'hca0001c;
      115835: inst = 32'h24822800;
      115836: inst = 32'h10a00000;
      115837: inst = 32'hca00004;
      115838: inst = 32'h38632800;
      115839: inst = 32'h38842800;
      115840: inst = 32'h10a00001;
      115841: inst = 32'hca0c485;
      115842: inst = 32'h13e00001;
      115843: inst = 32'hfe0d96a;
      115844: inst = 32'h5be00000;
      115845: inst = 32'h8c50000;
      115846: inst = 32'h24612800;
      115847: inst = 32'h10a00000;
      115848: inst = 32'hca0001c;
      115849: inst = 32'h24822800;
      115850: inst = 32'h10a00000;
      115851: inst = 32'hca00004;
      115852: inst = 32'h38632800;
      115853: inst = 32'h38842800;
      115854: inst = 32'h10a00001;
      115855: inst = 32'hca0c493;
      115856: inst = 32'h13e00001;
      115857: inst = 32'hfe0d96a;
      115858: inst = 32'h5be00000;
      115859: inst = 32'h8c50000;
      115860: inst = 32'h24612800;
      115861: inst = 32'h10a00000;
      115862: inst = 32'hca0001c;
      115863: inst = 32'h24822800;
      115864: inst = 32'h10a00000;
      115865: inst = 32'hca00004;
      115866: inst = 32'h38632800;
      115867: inst = 32'h38842800;
      115868: inst = 32'h10a00001;
      115869: inst = 32'hca0c4a1;
      115870: inst = 32'h13e00001;
      115871: inst = 32'hfe0d96a;
      115872: inst = 32'h5be00000;
      115873: inst = 32'h8c50000;
      115874: inst = 32'h24612800;
      115875: inst = 32'h10a00000;
      115876: inst = 32'hca0001c;
      115877: inst = 32'h24822800;
      115878: inst = 32'h10a00000;
      115879: inst = 32'hca00004;
      115880: inst = 32'h38632800;
      115881: inst = 32'h38842800;
      115882: inst = 32'h10a00001;
      115883: inst = 32'hca0c4af;
      115884: inst = 32'h13e00001;
      115885: inst = 32'hfe0d96a;
      115886: inst = 32'h5be00000;
      115887: inst = 32'h8c50000;
      115888: inst = 32'h24612800;
      115889: inst = 32'h10a00000;
      115890: inst = 32'hca0001c;
      115891: inst = 32'h24822800;
      115892: inst = 32'h10a00000;
      115893: inst = 32'hca00004;
      115894: inst = 32'h38632800;
      115895: inst = 32'h38842800;
      115896: inst = 32'h10a00001;
      115897: inst = 32'hca0c4bd;
      115898: inst = 32'h13e00001;
      115899: inst = 32'hfe0d96a;
      115900: inst = 32'h5be00000;
      115901: inst = 32'h8c50000;
      115902: inst = 32'h24612800;
      115903: inst = 32'h10a00000;
      115904: inst = 32'hca0001c;
      115905: inst = 32'h24822800;
      115906: inst = 32'h10a00000;
      115907: inst = 32'hca00004;
      115908: inst = 32'h38632800;
      115909: inst = 32'h38842800;
      115910: inst = 32'h10a00001;
      115911: inst = 32'hca0c4cb;
      115912: inst = 32'h13e00001;
      115913: inst = 32'hfe0d96a;
      115914: inst = 32'h5be00000;
      115915: inst = 32'h8c50000;
      115916: inst = 32'h24612800;
      115917: inst = 32'h10a00000;
      115918: inst = 32'hca0001c;
      115919: inst = 32'h24822800;
      115920: inst = 32'h10a00000;
      115921: inst = 32'hca00004;
      115922: inst = 32'h38632800;
      115923: inst = 32'h38842800;
      115924: inst = 32'h10a00001;
      115925: inst = 32'hca0c4d9;
      115926: inst = 32'h13e00001;
      115927: inst = 32'hfe0d96a;
      115928: inst = 32'h5be00000;
      115929: inst = 32'h8c50000;
      115930: inst = 32'h24612800;
      115931: inst = 32'h10a00000;
      115932: inst = 32'hca0001c;
      115933: inst = 32'h24822800;
      115934: inst = 32'h10a00000;
      115935: inst = 32'hca00004;
      115936: inst = 32'h38632800;
      115937: inst = 32'h38842800;
      115938: inst = 32'h10a00001;
      115939: inst = 32'hca0c4e7;
      115940: inst = 32'h13e00001;
      115941: inst = 32'hfe0d96a;
      115942: inst = 32'h5be00000;
      115943: inst = 32'h8c50000;
      115944: inst = 32'h24612800;
      115945: inst = 32'h10a00000;
      115946: inst = 32'hca0001c;
      115947: inst = 32'h24822800;
      115948: inst = 32'h10a00000;
      115949: inst = 32'hca00004;
      115950: inst = 32'h38632800;
      115951: inst = 32'h38842800;
      115952: inst = 32'h10a00001;
      115953: inst = 32'hca0c4f5;
      115954: inst = 32'h13e00001;
      115955: inst = 32'hfe0d96a;
      115956: inst = 32'h5be00000;
      115957: inst = 32'h8c50000;
      115958: inst = 32'h24612800;
      115959: inst = 32'h10a00000;
      115960: inst = 32'hca0001c;
      115961: inst = 32'h24822800;
      115962: inst = 32'h10a00000;
      115963: inst = 32'hca00004;
      115964: inst = 32'h38632800;
      115965: inst = 32'h38842800;
      115966: inst = 32'h10a00001;
      115967: inst = 32'hca0c503;
      115968: inst = 32'h13e00001;
      115969: inst = 32'hfe0d96a;
      115970: inst = 32'h5be00000;
      115971: inst = 32'h8c50000;
      115972: inst = 32'h24612800;
      115973: inst = 32'h10a00000;
      115974: inst = 32'hca0001c;
      115975: inst = 32'h24822800;
      115976: inst = 32'h10a00000;
      115977: inst = 32'hca00004;
      115978: inst = 32'h38632800;
      115979: inst = 32'h38842800;
      115980: inst = 32'h10a00001;
      115981: inst = 32'hca0c511;
      115982: inst = 32'h13e00001;
      115983: inst = 32'hfe0d96a;
      115984: inst = 32'h5be00000;
      115985: inst = 32'h8c50000;
      115986: inst = 32'h24612800;
      115987: inst = 32'h10a00000;
      115988: inst = 32'hca0001c;
      115989: inst = 32'h24822800;
      115990: inst = 32'h10a00000;
      115991: inst = 32'hca00004;
      115992: inst = 32'h38632800;
      115993: inst = 32'h38842800;
      115994: inst = 32'h10a00001;
      115995: inst = 32'hca0c51f;
      115996: inst = 32'h13e00001;
      115997: inst = 32'hfe0d96a;
      115998: inst = 32'h5be00000;
      115999: inst = 32'h8c50000;
      116000: inst = 32'h24612800;
      116001: inst = 32'h10a00000;
      116002: inst = 32'hca0001c;
      116003: inst = 32'h24822800;
      116004: inst = 32'h10a00000;
      116005: inst = 32'hca00004;
      116006: inst = 32'h38632800;
      116007: inst = 32'h38842800;
      116008: inst = 32'h10a00001;
      116009: inst = 32'hca0c52d;
      116010: inst = 32'h13e00001;
      116011: inst = 32'hfe0d96a;
      116012: inst = 32'h5be00000;
      116013: inst = 32'h8c50000;
      116014: inst = 32'h24612800;
      116015: inst = 32'h10a00000;
      116016: inst = 32'hca0001c;
      116017: inst = 32'h24822800;
      116018: inst = 32'h10a00000;
      116019: inst = 32'hca00004;
      116020: inst = 32'h38632800;
      116021: inst = 32'h38842800;
      116022: inst = 32'h10a00001;
      116023: inst = 32'hca0c53b;
      116024: inst = 32'h13e00001;
      116025: inst = 32'hfe0d96a;
      116026: inst = 32'h5be00000;
      116027: inst = 32'h8c50000;
      116028: inst = 32'h24612800;
      116029: inst = 32'h10a00000;
      116030: inst = 32'hca0001c;
      116031: inst = 32'h24822800;
      116032: inst = 32'h10a00000;
      116033: inst = 32'hca00004;
      116034: inst = 32'h38632800;
      116035: inst = 32'h38842800;
      116036: inst = 32'h10a00001;
      116037: inst = 32'hca0c549;
      116038: inst = 32'h13e00001;
      116039: inst = 32'hfe0d96a;
      116040: inst = 32'h5be00000;
      116041: inst = 32'h8c50000;
      116042: inst = 32'h24612800;
      116043: inst = 32'h10a00000;
      116044: inst = 32'hca0001c;
      116045: inst = 32'h24822800;
      116046: inst = 32'h10a00000;
      116047: inst = 32'hca00004;
      116048: inst = 32'h38632800;
      116049: inst = 32'h38842800;
      116050: inst = 32'h10a00001;
      116051: inst = 32'hca0c557;
      116052: inst = 32'h13e00001;
      116053: inst = 32'hfe0d96a;
      116054: inst = 32'h5be00000;
      116055: inst = 32'h8c50000;
      116056: inst = 32'h24612800;
      116057: inst = 32'h10a00000;
      116058: inst = 32'hca0001c;
      116059: inst = 32'h24822800;
      116060: inst = 32'h10a00000;
      116061: inst = 32'hca00004;
      116062: inst = 32'h38632800;
      116063: inst = 32'h38842800;
      116064: inst = 32'h10a00001;
      116065: inst = 32'hca0c565;
      116066: inst = 32'h13e00001;
      116067: inst = 32'hfe0d96a;
      116068: inst = 32'h5be00000;
      116069: inst = 32'h8c50000;
      116070: inst = 32'h24612800;
      116071: inst = 32'h10a00000;
      116072: inst = 32'hca0001c;
      116073: inst = 32'h24822800;
      116074: inst = 32'h10a00000;
      116075: inst = 32'hca00004;
      116076: inst = 32'h38632800;
      116077: inst = 32'h38842800;
      116078: inst = 32'h10a00001;
      116079: inst = 32'hca0c573;
      116080: inst = 32'h13e00001;
      116081: inst = 32'hfe0d96a;
      116082: inst = 32'h5be00000;
      116083: inst = 32'h8c50000;
      116084: inst = 32'h24612800;
      116085: inst = 32'h10a00000;
      116086: inst = 32'hca0001c;
      116087: inst = 32'h24822800;
      116088: inst = 32'h10a00000;
      116089: inst = 32'hca00004;
      116090: inst = 32'h38632800;
      116091: inst = 32'h38842800;
      116092: inst = 32'h10a00001;
      116093: inst = 32'hca0c581;
      116094: inst = 32'h13e00001;
      116095: inst = 32'hfe0d96a;
      116096: inst = 32'h5be00000;
      116097: inst = 32'h8c50000;
      116098: inst = 32'h24612800;
      116099: inst = 32'h10a00000;
      116100: inst = 32'hca0001c;
      116101: inst = 32'h24822800;
      116102: inst = 32'h10a00000;
      116103: inst = 32'hca00004;
      116104: inst = 32'h38632800;
      116105: inst = 32'h38842800;
      116106: inst = 32'h10a00001;
      116107: inst = 32'hca0c58f;
      116108: inst = 32'h13e00001;
      116109: inst = 32'hfe0d96a;
      116110: inst = 32'h5be00000;
      116111: inst = 32'h8c50000;
      116112: inst = 32'h24612800;
      116113: inst = 32'h10a00000;
      116114: inst = 32'hca0001c;
      116115: inst = 32'h24822800;
      116116: inst = 32'h10a00000;
      116117: inst = 32'hca00004;
      116118: inst = 32'h38632800;
      116119: inst = 32'h38842800;
      116120: inst = 32'h10a00001;
      116121: inst = 32'hca0c59d;
      116122: inst = 32'h13e00001;
      116123: inst = 32'hfe0d96a;
      116124: inst = 32'h5be00000;
      116125: inst = 32'h8c50000;
      116126: inst = 32'h24612800;
      116127: inst = 32'h10a00000;
      116128: inst = 32'hca0001c;
      116129: inst = 32'h24822800;
      116130: inst = 32'h10a00000;
      116131: inst = 32'hca00004;
      116132: inst = 32'h38632800;
      116133: inst = 32'h38842800;
      116134: inst = 32'h10a00001;
      116135: inst = 32'hca0c5ab;
      116136: inst = 32'h13e00001;
      116137: inst = 32'hfe0d96a;
      116138: inst = 32'h5be00000;
      116139: inst = 32'h8c50000;
      116140: inst = 32'h24612800;
      116141: inst = 32'h10a00000;
      116142: inst = 32'hca0001c;
      116143: inst = 32'h24822800;
      116144: inst = 32'h10a00000;
      116145: inst = 32'hca00004;
      116146: inst = 32'h38632800;
      116147: inst = 32'h38842800;
      116148: inst = 32'h10a00001;
      116149: inst = 32'hca0c5b9;
      116150: inst = 32'h13e00001;
      116151: inst = 32'hfe0d96a;
      116152: inst = 32'h5be00000;
      116153: inst = 32'h8c50000;
      116154: inst = 32'h24612800;
      116155: inst = 32'h10a00000;
      116156: inst = 32'hca0001c;
      116157: inst = 32'h24822800;
      116158: inst = 32'h10a00000;
      116159: inst = 32'hca00004;
      116160: inst = 32'h38632800;
      116161: inst = 32'h38842800;
      116162: inst = 32'h10a00001;
      116163: inst = 32'hca0c5c7;
      116164: inst = 32'h13e00001;
      116165: inst = 32'hfe0d96a;
      116166: inst = 32'h5be00000;
      116167: inst = 32'h8c50000;
      116168: inst = 32'h24612800;
      116169: inst = 32'h10a00000;
      116170: inst = 32'hca0001c;
      116171: inst = 32'h24822800;
      116172: inst = 32'h10a00000;
      116173: inst = 32'hca00004;
      116174: inst = 32'h38632800;
      116175: inst = 32'h38842800;
      116176: inst = 32'h10a00001;
      116177: inst = 32'hca0c5d5;
      116178: inst = 32'h13e00001;
      116179: inst = 32'hfe0d96a;
      116180: inst = 32'h5be00000;
      116181: inst = 32'h8c50000;
      116182: inst = 32'h24612800;
      116183: inst = 32'h10a00000;
      116184: inst = 32'hca0001c;
      116185: inst = 32'h24822800;
      116186: inst = 32'h10a00000;
      116187: inst = 32'hca00004;
      116188: inst = 32'h38632800;
      116189: inst = 32'h38842800;
      116190: inst = 32'h10a00001;
      116191: inst = 32'hca0c5e3;
      116192: inst = 32'h13e00001;
      116193: inst = 32'hfe0d96a;
      116194: inst = 32'h5be00000;
      116195: inst = 32'h8c50000;
      116196: inst = 32'h24612800;
      116197: inst = 32'h10a00000;
      116198: inst = 32'hca0001c;
      116199: inst = 32'h24822800;
      116200: inst = 32'h10a00000;
      116201: inst = 32'hca00004;
      116202: inst = 32'h38632800;
      116203: inst = 32'h38842800;
      116204: inst = 32'h10a00001;
      116205: inst = 32'hca0c5f1;
      116206: inst = 32'h13e00001;
      116207: inst = 32'hfe0d96a;
      116208: inst = 32'h5be00000;
      116209: inst = 32'h8c50000;
      116210: inst = 32'h24612800;
      116211: inst = 32'h10a00000;
      116212: inst = 32'hca0001c;
      116213: inst = 32'h24822800;
      116214: inst = 32'h10a00000;
      116215: inst = 32'hca00004;
      116216: inst = 32'h38632800;
      116217: inst = 32'h38842800;
      116218: inst = 32'h10a00001;
      116219: inst = 32'hca0c5ff;
      116220: inst = 32'h13e00001;
      116221: inst = 32'hfe0d96a;
      116222: inst = 32'h5be00000;
      116223: inst = 32'h8c50000;
      116224: inst = 32'h24612800;
      116225: inst = 32'h10a00000;
      116226: inst = 32'hca0001c;
      116227: inst = 32'h24822800;
      116228: inst = 32'h10a00000;
      116229: inst = 32'hca00004;
      116230: inst = 32'h38632800;
      116231: inst = 32'h38842800;
      116232: inst = 32'h10a00001;
      116233: inst = 32'hca0c60d;
      116234: inst = 32'h13e00001;
      116235: inst = 32'hfe0d96a;
      116236: inst = 32'h5be00000;
      116237: inst = 32'h8c50000;
      116238: inst = 32'h24612800;
      116239: inst = 32'h10a00000;
      116240: inst = 32'hca0001c;
      116241: inst = 32'h24822800;
      116242: inst = 32'h10a00000;
      116243: inst = 32'hca00004;
      116244: inst = 32'h38632800;
      116245: inst = 32'h38842800;
      116246: inst = 32'h10a00001;
      116247: inst = 32'hca0c61b;
      116248: inst = 32'h13e00001;
      116249: inst = 32'hfe0d96a;
      116250: inst = 32'h5be00000;
      116251: inst = 32'h8c50000;
      116252: inst = 32'h24612800;
      116253: inst = 32'h10a00000;
      116254: inst = 32'hca0001c;
      116255: inst = 32'h24822800;
      116256: inst = 32'h10a00000;
      116257: inst = 32'hca00004;
      116258: inst = 32'h38632800;
      116259: inst = 32'h38842800;
      116260: inst = 32'h10a00001;
      116261: inst = 32'hca0c629;
      116262: inst = 32'h13e00001;
      116263: inst = 32'hfe0d96a;
      116264: inst = 32'h5be00000;
      116265: inst = 32'h8c50000;
      116266: inst = 32'h24612800;
      116267: inst = 32'h10a00000;
      116268: inst = 32'hca0001c;
      116269: inst = 32'h24822800;
      116270: inst = 32'h10a00000;
      116271: inst = 32'hca00004;
      116272: inst = 32'h38632800;
      116273: inst = 32'h38842800;
      116274: inst = 32'h10a00001;
      116275: inst = 32'hca0c637;
      116276: inst = 32'h13e00001;
      116277: inst = 32'hfe0d96a;
      116278: inst = 32'h5be00000;
      116279: inst = 32'h8c50000;
      116280: inst = 32'h24612800;
      116281: inst = 32'h10a00000;
      116282: inst = 32'hca0001c;
      116283: inst = 32'h24822800;
      116284: inst = 32'h10a00000;
      116285: inst = 32'hca00004;
      116286: inst = 32'h38632800;
      116287: inst = 32'h38842800;
      116288: inst = 32'h10a00001;
      116289: inst = 32'hca0c645;
      116290: inst = 32'h13e00001;
      116291: inst = 32'hfe0d96a;
      116292: inst = 32'h5be00000;
      116293: inst = 32'h8c50000;
      116294: inst = 32'h24612800;
      116295: inst = 32'h10a00000;
      116296: inst = 32'hca0001c;
      116297: inst = 32'h24822800;
      116298: inst = 32'h10a00000;
      116299: inst = 32'hca00004;
      116300: inst = 32'h38632800;
      116301: inst = 32'h38842800;
      116302: inst = 32'h10a00001;
      116303: inst = 32'hca0c653;
      116304: inst = 32'h13e00001;
      116305: inst = 32'hfe0d96a;
      116306: inst = 32'h5be00000;
      116307: inst = 32'h8c50000;
      116308: inst = 32'h24612800;
      116309: inst = 32'h10a00000;
      116310: inst = 32'hca0001c;
      116311: inst = 32'h24822800;
      116312: inst = 32'h10a00000;
      116313: inst = 32'hca00004;
      116314: inst = 32'h38632800;
      116315: inst = 32'h38842800;
      116316: inst = 32'h10a00001;
      116317: inst = 32'hca0c661;
      116318: inst = 32'h13e00001;
      116319: inst = 32'hfe0d96a;
      116320: inst = 32'h5be00000;
      116321: inst = 32'h8c50000;
      116322: inst = 32'h24612800;
      116323: inst = 32'h10a00000;
      116324: inst = 32'hca0001c;
      116325: inst = 32'h24822800;
      116326: inst = 32'h10a00000;
      116327: inst = 32'hca00004;
      116328: inst = 32'h38632800;
      116329: inst = 32'h38842800;
      116330: inst = 32'h10a00001;
      116331: inst = 32'hca0c66f;
      116332: inst = 32'h13e00001;
      116333: inst = 32'hfe0d96a;
      116334: inst = 32'h5be00000;
      116335: inst = 32'h8c50000;
      116336: inst = 32'h24612800;
      116337: inst = 32'h10a00000;
      116338: inst = 32'hca0001c;
      116339: inst = 32'h24822800;
      116340: inst = 32'h10a00000;
      116341: inst = 32'hca00004;
      116342: inst = 32'h38632800;
      116343: inst = 32'h38842800;
      116344: inst = 32'h10a00001;
      116345: inst = 32'hca0c67d;
      116346: inst = 32'h13e00001;
      116347: inst = 32'hfe0d96a;
      116348: inst = 32'h5be00000;
      116349: inst = 32'h8c50000;
      116350: inst = 32'h24612800;
      116351: inst = 32'h10a00000;
      116352: inst = 32'hca0001c;
      116353: inst = 32'h24822800;
      116354: inst = 32'h10a00000;
      116355: inst = 32'hca00004;
      116356: inst = 32'h38632800;
      116357: inst = 32'h38842800;
      116358: inst = 32'h10a00001;
      116359: inst = 32'hca0c68b;
      116360: inst = 32'h13e00001;
      116361: inst = 32'hfe0d96a;
      116362: inst = 32'h5be00000;
      116363: inst = 32'h8c50000;
      116364: inst = 32'h24612800;
      116365: inst = 32'h10a00000;
      116366: inst = 32'hca0001c;
      116367: inst = 32'h24822800;
      116368: inst = 32'h10a00000;
      116369: inst = 32'hca00004;
      116370: inst = 32'h38632800;
      116371: inst = 32'h38842800;
      116372: inst = 32'h10a00001;
      116373: inst = 32'hca0c699;
      116374: inst = 32'h13e00001;
      116375: inst = 32'hfe0d96a;
      116376: inst = 32'h5be00000;
      116377: inst = 32'h8c50000;
      116378: inst = 32'h24612800;
      116379: inst = 32'h10a00000;
      116380: inst = 32'hca0001c;
      116381: inst = 32'h24822800;
      116382: inst = 32'h10a00000;
      116383: inst = 32'hca00004;
      116384: inst = 32'h38632800;
      116385: inst = 32'h38842800;
      116386: inst = 32'h10a00001;
      116387: inst = 32'hca0c6a7;
      116388: inst = 32'h13e00001;
      116389: inst = 32'hfe0d96a;
      116390: inst = 32'h5be00000;
      116391: inst = 32'h8c50000;
      116392: inst = 32'h24612800;
      116393: inst = 32'h10a00000;
      116394: inst = 32'hca0001c;
      116395: inst = 32'h24822800;
      116396: inst = 32'h10a00000;
      116397: inst = 32'hca00004;
      116398: inst = 32'h38632800;
      116399: inst = 32'h38842800;
      116400: inst = 32'h10a00001;
      116401: inst = 32'hca0c6b5;
      116402: inst = 32'h13e00001;
      116403: inst = 32'hfe0d96a;
      116404: inst = 32'h5be00000;
      116405: inst = 32'h8c50000;
      116406: inst = 32'h24612800;
      116407: inst = 32'h10a00000;
      116408: inst = 32'hca0001c;
      116409: inst = 32'h24822800;
      116410: inst = 32'h10a00000;
      116411: inst = 32'hca00004;
      116412: inst = 32'h38632800;
      116413: inst = 32'h38842800;
      116414: inst = 32'h10a00001;
      116415: inst = 32'hca0c6c3;
      116416: inst = 32'h13e00001;
      116417: inst = 32'hfe0d96a;
      116418: inst = 32'h5be00000;
      116419: inst = 32'h8c50000;
      116420: inst = 32'h24612800;
      116421: inst = 32'h10a00000;
      116422: inst = 32'hca0001c;
      116423: inst = 32'h24822800;
      116424: inst = 32'h10a00000;
      116425: inst = 32'hca00004;
      116426: inst = 32'h38632800;
      116427: inst = 32'h38842800;
      116428: inst = 32'h10a00001;
      116429: inst = 32'hca0c6d1;
      116430: inst = 32'h13e00001;
      116431: inst = 32'hfe0d96a;
      116432: inst = 32'h5be00000;
      116433: inst = 32'h8c50000;
      116434: inst = 32'h24612800;
      116435: inst = 32'h10a00000;
      116436: inst = 32'hca0001c;
      116437: inst = 32'h24822800;
      116438: inst = 32'h10a00000;
      116439: inst = 32'hca00004;
      116440: inst = 32'h38632800;
      116441: inst = 32'h38842800;
      116442: inst = 32'h10a00001;
      116443: inst = 32'hca0c6df;
      116444: inst = 32'h13e00001;
      116445: inst = 32'hfe0d96a;
      116446: inst = 32'h5be00000;
      116447: inst = 32'h8c50000;
      116448: inst = 32'h24612800;
      116449: inst = 32'h10a00000;
      116450: inst = 32'hca0001c;
      116451: inst = 32'h24822800;
      116452: inst = 32'h10a00000;
      116453: inst = 32'hca00004;
      116454: inst = 32'h38632800;
      116455: inst = 32'h38842800;
      116456: inst = 32'h10a00001;
      116457: inst = 32'hca0c6ed;
      116458: inst = 32'h13e00001;
      116459: inst = 32'hfe0d96a;
      116460: inst = 32'h5be00000;
      116461: inst = 32'h8c50000;
      116462: inst = 32'h24612800;
      116463: inst = 32'h10a00000;
      116464: inst = 32'hca0001c;
      116465: inst = 32'h24822800;
      116466: inst = 32'h10a00000;
      116467: inst = 32'hca00004;
      116468: inst = 32'h38632800;
      116469: inst = 32'h38842800;
      116470: inst = 32'h10a00001;
      116471: inst = 32'hca0c6fb;
      116472: inst = 32'h13e00001;
      116473: inst = 32'hfe0d96a;
      116474: inst = 32'h5be00000;
      116475: inst = 32'h8c50000;
      116476: inst = 32'h24612800;
      116477: inst = 32'h10a00000;
      116478: inst = 32'hca0001c;
      116479: inst = 32'h24822800;
      116480: inst = 32'h10a00000;
      116481: inst = 32'hca00004;
      116482: inst = 32'h38632800;
      116483: inst = 32'h38842800;
      116484: inst = 32'h10a00001;
      116485: inst = 32'hca0c709;
      116486: inst = 32'h13e00001;
      116487: inst = 32'hfe0d96a;
      116488: inst = 32'h5be00000;
      116489: inst = 32'h8c50000;
      116490: inst = 32'h24612800;
      116491: inst = 32'h10a00000;
      116492: inst = 32'hca0001c;
      116493: inst = 32'h24822800;
      116494: inst = 32'h10a00000;
      116495: inst = 32'hca00004;
      116496: inst = 32'h38632800;
      116497: inst = 32'h38842800;
      116498: inst = 32'h10a00001;
      116499: inst = 32'hca0c717;
      116500: inst = 32'h13e00001;
      116501: inst = 32'hfe0d96a;
      116502: inst = 32'h5be00000;
      116503: inst = 32'h8c50000;
      116504: inst = 32'h24612800;
      116505: inst = 32'h10a00000;
      116506: inst = 32'hca0001c;
      116507: inst = 32'h24822800;
      116508: inst = 32'h10a00000;
      116509: inst = 32'hca00004;
      116510: inst = 32'h38632800;
      116511: inst = 32'h38842800;
      116512: inst = 32'h10a00001;
      116513: inst = 32'hca0c725;
      116514: inst = 32'h13e00001;
      116515: inst = 32'hfe0d96a;
      116516: inst = 32'h5be00000;
      116517: inst = 32'h8c50000;
      116518: inst = 32'h24612800;
      116519: inst = 32'h10a00000;
      116520: inst = 32'hca0001c;
      116521: inst = 32'h24822800;
      116522: inst = 32'h10a00000;
      116523: inst = 32'hca00004;
      116524: inst = 32'h38632800;
      116525: inst = 32'h38842800;
      116526: inst = 32'h10a00001;
      116527: inst = 32'hca0c733;
      116528: inst = 32'h13e00001;
      116529: inst = 32'hfe0d96a;
      116530: inst = 32'h5be00000;
      116531: inst = 32'h8c50000;
      116532: inst = 32'h24612800;
      116533: inst = 32'h10a00000;
      116534: inst = 32'hca0001c;
      116535: inst = 32'h24822800;
      116536: inst = 32'h10a00000;
      116537: inst = 32'hca00004;
      116538: inst = 32'h38632800;
      116539: inst = 32'h38842800;
      116540: inst = 32'h10a00001;
      116541: inst = 32'hca0c741;
      116542: inst = 32'h13e00001;
      116543: inst = 32'hfe0d96a;
      116544: inst = 32'h5be00000;
      116545: inst = 32'h8c50000;
      116546: inst = 32'h24612800;
      116547: inst = 32'h10a00000;
      116548: inst = 32'hca0001c;
      116549: inst = 32'h24822800;
      116550: inst = 32'h10a00000;
      116551: inst = 32'hca00004;
      116552: inst = 32'h38632800;
      116553: inst = 32'h38842800;
      116554: inst = 32'h10a00001;
      116555: inst = 32'hca0c74f;
      116556: inst = 32'h13e00001;
      116557: inst = 32'hfe0d96a;
      116558: inst = 32'h5be00000;
      116559: inst = 32'h8c50000;
      116560: inst = 32'h24612800;
      116561: inst = 32'h10a00000;
      116562: inst = 32'hca0001c;
      116563: inst = 32'h24822800;
      116564: inst = 32'h10a00000;
      116565: inst = 32'hca00004;
      116566: inst = 32'h38632800;
      116567: inst = 32'h38842800;
      116568: inst = 32'h10a00001;
      116569: inst = 32'hca0c75d;
      116570: inst = 32'h13e00001;
      116571: inst = 32'hfe0d96a;
      116572: inst = 32'h5be00000;
      116573: inst = 32'h8c50000;
      116574: inst = 32'h24612800;
      116575: inst = 32'h10a00000;
      116576: inst = 32'hca0001c;
      116577: inst = 32'h24822800;
      116578: inst = 32'h10a00000;
      116579: inst = 32'hca00004;
      116580: inst = 32'h38632800;
      116581: inst = 32'h38842800;
      116582: inst = 32'h10a00001;
      116583: inst = 32'hca0c76b;
      116584: inst = 32'h13e00001;
      116585: inst = 32'hfe0d96a;
      116586: inst = 32'h5be00000;
      116587: inst = 32'h8c50000;
      116588: inst = 32'h24612800;
      116589: inst = 32'h10a00000;
      116590: inst = 32'hca0001c;
      116591: inst = 32'h24822800;
      116592: inst = 32'h10a00000;
      116593: inst = 32'hca00004;
      116594: inst = 32'h38632800;
      116595: inst = 32'h38842800;
      116596: inst = 32'h10a00001;
      116597: inst = 32'hca0c779;
      116598: inst = 32'h13e00001;
      116599: inst = 32'hfe0d96a;
      116600: inst = 32'h5be00000;
      116601: inst = 32'h8c50000;
      116602: inst = 32'h24612800;
      116603: inst = 32'h10a00000;
      116604: inst = 32'hca0001c;
      116605: inst = 32'h24822800;
      116606: inst = 32'h10a00000;
      116607: inst = 32'hca00004;
      116608: inst = 32'h38632800;
      116609: inst = 32'h38842800;
      116610: inst = 32'h10a00001;
      116611: inst = 32'hca0c787;
      116612: inst = 32'h13e00001;
      116613: inst = 32'hfe0d96a;
      116614: inst = 32'h5be00000;
      116615: inst = 32'h8c50000;
      116616: inst = 32'h24612800;
      116617: inst = 32'h10a00000;
      116618: inst = 32'hca0001c;
      116619: inst = 32'h24822800;
      116620: inst = 32'h10a00000;
      116621: inst = 32'hca00004;
      116622: inst = 32'h38632800;
      116623: inst = 32'h38842800;
      116624: inst = 32'h10a00001;
      116625: inst = 32'hca0c795;
      116626: inst = 32'h13e00001;
      116627: inst = 32'hfe0d96a;
      116628: inst = 32'h5be00000;
      116629: inst = 32'h8c50000;
      116630: inst = 32'h24612800;
      116631: inst = 32'h10a00000;
      116632: inst = 32'hca0001c;
      116633: inst = 32'h24822800;
      116634: inst = 32'h10a00000;
      116635: inst = 32'hca00004;
      116636: inst = 32'h38632800;
      116637: inst = 32'h38842800;
      116638: inst = 32'h10a00001;
      116639: inst = 32'hca0c7a3;
      116640: inst = 32'h13e00001;
      116641: inst = 32'hfe0d96a;
      116642: inst = 32'h5be00000;
      116643: inst = 32'h8c50000;
      116644: inst = 32'h24612800;
      116645: inst = 32'h10a00000;
      116646: inst = 32'hca0001c;
      116647: inst = 32'h24822800;
      116648: inst = 32'h10a00000;
      116649: inst = 32'hca00004;
      116650: inst = 32'h38632800;
      116651: inst = 32'h38842800;
      116652: inst = 32'h10a00001;
      116653: inst = 32'hca0c7b1;
      116654: inst = 32'h13e00001;
      116655: inst = 32'hfe0d96a;
      116656: inst = 32'h5be00000;
      116657: inst = 32'h8c50000;
      116658: inst = 32'h24612800;
      116659: inst = 32'h10a00000;
      116660: inst = 32'hca0001c;
      116661: inst = 32'h24822800;
      116662: inst = 32'h10a00000;
      116663: inst = 32'hca00004;
      116664: inst = 32'h38632800;
      116665: inst = 32'h38842800;
      116666: inst = 32'h10a00001;
      116667: inst = 32'hca0c7bf;
      116668: inst = 32'h13e00001;
      116669: inst = 32'hfe0d96a;
      116670: inst = 32'h5be00000;
      116671: inst = 32'h8c50000;
      116672: inst = 32'h24612800;
      116673: inst = 32'h10a00000;
      116674: inst = 32'hca0001c;
      116675: inst = 32'h24822800;
      116676: inst = 32'h10a00000;
      116677: inst = 32'hca00004;
      116678: inst = 32'h38632800;
      116679: inst = 32'h38842800;
      116680: inst = 32'h10a00001;
      116681: inst = 32'hca0c7cd;
      116682: inst = 32'h13e00001;
      116683: inst = 32'hfe0d96a;
      116684: inst = 32'h5be00000;
      116685: inst = 32'h8c50000;
      116686: inst = 32'h24612800;
      116687: inst = 32'h10a00000;
      116688: inst = 32'hca0001c;
      116689: inst = 32'h24822800;
      116690: inst = 32'h10a00000;
      116691: inst = 32'hca00004;
      116692: inst = 32'h38632800;
      116693: inst = 32'h38842800;
      116694: inst = 32'h10a00001;
      116695: inst = 32'hca0c7db;
      116696: inst = 32'h13e00001;
      116697: inst = 32'hfe0d96a;
      116698: inst = 32'h5be00000;
      116699: inst = 32'h8c50000;
      116700: inst = 32'h24612800;
      116701: inst = 32'h10a00000;
      116702: inst = 32'hca0001c;
      116703: inst = 32'h24822800;
      116704: inst = 32'h10a00000;
      116705: inst = 32'hca00004;
      116706: inst = 32'h38632800;
      116707: inst = 32'h38842800;
      116708: inst = 32'h10a00001;
      116709: inst = 32'hca0c7e9;
      116710: inst = 32'h13e00001;
      116711: inst = 32'hfe0d96a;
      116712: inst = 32'h5be00000;
      116713: inst = 32'h8c50000;
      116714: inst = 32'h24612800;
      116715: inst = 32'h10a00000;
      116716: inst = 32'hca0001c;
      116717: inst = 32'h24822800;
      116718: inst = 32'h10a00000;
      116719: inst = 32'hca00004;
      116720: inst = 32'h38632800;
      116721: inst = 32'h38842800;
      116722: inst = 32'h10a00001;
      116723: inst = 32'hca0c7f7;
      116724: inst = 32'h13e00001;
      116725: inst = 32'hfe0d96a;
      116726: inst = 32'h5be00000;
      116727: inst = 32'h8c50000;
      116728: inst = 32'h24612800;
      116729: inst = 32'h10a00000;
      116730: inst = 32'hca0001c;
      116731: inst = 32'h24822800;
      116732: inst = 32'h10a00000;
      116733: inst = 32'hca00004;
      116734: inst = 32'h38632800;
      116735: inst = 32'h38842800;
      116736: inst = 32'h10a00001;
      116737: inst = 32'hca0c805;
      116738: inst = 32'h13e00001;
      116739: inst = 32'hfe0d96a;
      116740: inst = 32'h5be00000;
      116741: inst = 32'h8c50000;
      116742: inst = 32'h24612800;
      116743: inst = 32'h10a00000;
      116744: inst = 32'hca0001c;
      116745: inst = 32'h24822800;
      116746: inst = 32'h10a00000;
      116747: inst = 32'hca00004;
      116748: inst = 32'h38632800;
      116749: inst = 32'h38842800;
      116750: inst = 32'h10a00001;
      116751: inst = 32'hca0c813;
      116752: inst = 32'h13e00001;
      116753: inst = 32'hfe0d96a;
      116754: inst = 32'h5be00000;
      116755: inst = 32'h8c50000;
      116756: inst = 32'h24612800;
      116757: inst = 32'h10a00000;
      116758: inst = 32'hca0001c;
      116759: inst = 32'h24822800;
      116760: inst = 32'h10a00000;
      116761: inst = 32'hca00004;
      116762: inst = 32'h38632800;
      116763: inst = 32'h38842800;
      116764: inst = 32'h10a00001;
      116765: inst = 32'hca0c821;
      116766: inst = 32'h13e00001;
      116767: inst = 32'hfe0d96a;
      116768: inst = 32'h5be00000;
      116769: inst = 32'h8c50000;
      116770: inst = 32'h24612800;
      116771: inst = 32'h10a00000;
      116772: inst = 32'hca0001c;
      116773: inst = 32'h24822800;
      116774: inst = 32'h10a00000;
      116775: inst = 32'hca00004;
      116776: inst = 32'h38632800;
      116777: inst = 32'h38842800;
      116778: inst = 32'h10a00001;
      116779: inst = 32'hca0c82f;
      116780: inst = 32'h13e00001;
      116781: inst = 32'hfe0d96a;
      116782: inst = 32'h5be00000;
      116783: inst = 32'h8c50000;
      116784: inst = 32'h24612800;
      116785: inst = 32'h10a00000;
      116786: inst = 32'hca0001c;
      116787: inst = 32'h24822800;
      116788: inst = 32'h10a00000;
      116789: inst = 32'hca00004;
      116790: inst = 32'h38632800;
      116791: inst = 32'h38842800;
      116792: inst = 32'h10a00001;
      116793: inst = 32'hca0c83d;
      116794: inst = 32'h13e00001;
      116795: inst = 32'hfe0d96a;
      116796: inst = 32'h5be00000;
      116797: inst = 32'h8c50000;
      116798: inst = 32'h24612800;
      116799: inst = 32'h10a00000;
      116800: inst = 32'hca0001c;
      116801: inst = 32'h24822800;
      116802: inst = 32'h10a00000;
      116803: inst = 32'hca00004;
      116804: inst = 32'h38632800;
      116805: inst = 32'h38842800;
      116806: inst = 32'h10a00001;
      116807: inst = 32'hca0c84b;
      116808: inst = 32'h13e00001;
      116809: inst = 32'hfe0d96a;
      116810: inst = 32'h5be00000;
      116811: inst = 32'h8c50000;
      116812: inst = 32'h24612800;
      116813: inst = 32'h10a00000;
      116814: inst = 32'hca0001c;
      116815: inst = 32'h24822800;
      116816: inst = 32'h10a00000;
      116817: inst = 32'hca00004;
      116818: inst = 32'h38632800;
      116819: inst = 32'h38842800;
      116820: inst = 32'h10a00001;
      116821: inst = 32'hca0c859;
      116822: inst = 32'h13e00001;
      116823: inst = 32'hfe0d96a;
      116824: inst = 32'h5be00000;
      116825: inst = 32'h8c50000;
      116826: inst = 32'h24612800;
      116827: inst = 32'h10a00000;
      116828: inst = 32'hca0001c;
      116829: inst = 32'h24822800;
      116830: inst = 32'h10a00000;
      116831: inst = 32'hca00004;
      116832: inst = 32'h38632800;
      116833: inst = 32'h38842800;
      116834: inst = 32'h10a00001;
      116835: inst = 32'hca0c867;
      116836: inst = 32'h13e00001;
      116837: inst = 32'hfe0d96a;
      116838: inst = 32'h5be00000;
      116839: inst = 32'h8c50000;
      116840: inst = 32'h24612800;
      116841: inst = 32'h10a00000;
      116842: inst = 32'hca0001c;
      116843: inst = 32'h24822800;
      116844: inst = 32'h10a00000;
      116845: inst = 32'hca00004;
      116846: inst = 32'h38632800;
      116847: inst = 32'h38842800;
      116848: inst = 32'h10a00001;
      116849: inst = 32'hca0c875;
      116850: inst = 32'h13e00001;
      116851: inst = 32'hfe0d96a;
      116852: inst = 32'h5be00000;
      116853: inst = 32'h8c50000;
      116854: inst = 32'h24612800;
      116855: inst = 32'h10a00000;
      116856: inst = 32'hca0001c;
      116857: inst = 32'h24822800;
      116858: inst = 32'h10a00000;
      116859: inst = 32'hca00004;
      116860: inst = 32'h38632800;
      116861: inst = 32'h38842800;
      116862: inst = 32'h10a00001;
      116863: inst = 32'hca0c883;
      116864: inst = 32'h13e00001;
      116865: inst = 32'hfe0d96a;
      116866: inst = 32'h5be00000;
      116867: inst = 32'h8c50000;
      116868: inst = 32'h24612800;
      116869: inst = 32'h10a00000;
      116870: inst = 32'hca0001c;
      116871: inst = 32'h24822800;
      116872: inst = 32'h10a00000;
      116873: inst = 32'hca00004;
      116874: inst = 32'h38632800;
      116875: inst = 32'h38842800;
      116876: inst = 32'h10a00001;
      116877: inst = 32'hca0c891;
      116878: inst = 32'h13e00001;
      116879: inst = 32'hfe0d96a;
      116880: inst = 32'h5be00000;
      116881: inst = 32'h8c50000;
      116882: inst = 32'h24612800;
      116883: inst = 32'h10a00000;
      116884: inst = 32'hca0001c;
      116885: inst = 32'h24822800;
      116886: inst = 32'h10a00000;
      116887: inst = 32'hca00004;
      116888: inst = 32'h38632800;
      116889: inst = 32'h38842800;
      116890: inst = 32'h10a00001;
      116891: inst = 32'hca0c89f;
      116892: inst = 32'h13e00001;
      116893: inst = 32'hfe0d96a;
      116894: inst = 32'h5be00000;
      116895: inst = 32'h8c50000;
      116896: inst = 32'h24612800;
      116897: inst = 32'h10a00000;
      116898: inst = 32'hca0001c;
      116899: inst = 32'h24822800;
      116900: inst = 32'h10a00000;
      116901: inst = 32'hca00004;
      116902: inst = 32'h38632800;
      116903: inst = 32'h38842800;
      116904: inst = 32'h10a00001;
      116905: inst = 32'hca0c8ad;
      116906: inst = 32'h13e00001;
      116907: inst = 32'hfe0d96a;
      116908: inst = 32'h5be00000;
      116909: inst = 32'h8c50000;
      116910: inst = 32'h24612800;
      116911: inst = 32'h10a00000;
      116912: inst = 32'hca0001c;
      116913: inst = 32'h24822800;
      116914: inst = 32'h10a00000;
      116915: inst = 32'hca00004;
      116916: inst = 32'h38632800;
      116917: inst = 32'h38842800;
      116918: inst = 32'h10a00001;
      116919: inst = 32'hca0c8bb;
      116920: inst = 32'h13e00001;
      116921: inst = 32'hfe0d96a;
      116922: inst = 32'h5be00000;
      116923: inst = 32'h8c50000;
      116924: inst = 32'h24612800;
      116925: inst = 32'h10a00000;
      116926: inst = 32'hca0001c;
      116927: inst = 32'h24822800;
      116928: inst = 32'h10a00000;
      116929: inst = 32'hca00004;
      116930: inst = 32'h38632800;
      116931: inst = 32'h38842800;
      116932: inst = 32'h10a00001;
      116933: inst = 32'hca0c8c9;
      116934: inst = 32'h13e00001;
      116935: inst = 32'hfe0d96a;
      116936: inst = 32'h5be00000;
      116937: inst = 32'h8c50000;
      116938: inst = 32'h24612800;
      116939: inst = 32'h10a00000;
      116940: inst = 32'hca0001c;
      116941: inst = 32'h24822800;
      116942: inst = 32'h10a00000;
      116943: inst = 32'hca00004;
      116944: inst = 32'h38632800;
      116945: inst = 32'h38842800;
      116946: inst = 32'h10a00001;
      116947: inst = 32'hca0c8d7;
      116948: inst = 32'h13e00001;
      116949: inst = 32'hfe0d96a;
      116950: inst = 32'h5be00000;
      116951: inst = 32'h8c50000;
      116952: inst = 32'h24612800;
      116953: inst = 32'h10a00000;
      116954: inst = 32'hca0001c;
      116955: inst = 32'h24822800;
      116956: inst = 32'h10a00000;
      116957: inst = 32'hca00004;
      116958: inst = 32'h38632800;
      116959: inst = 32'h38842800;
      116960: inst = 32'h10a00001;
      116961: inst = 32'hca0c8e5;
      116962: inst = 32'h13e00001;
      116963: inst = 32'hfe0d96a;
      116964: inst = 32'h5be00000;
      116965: inst = 32'h8c50000;
      116966: inst = 32'h24612800;
      116967: inst = 32'h10a00000;
      116968: inst = 32'hca0001c;
      116969: inst = 32'h24822800;
      116970: inst = 32'h10a00000;
      116971: inst = 32'hca00004;
      116972: inst = 32'h38632800;
      116973: inst = 32'h38842800;
      116974: inst = 32'h10a00001;
      116975: inst = 32'hca0c8f3;
      116976: inst = 32'h13e00001;
      116977: inst = 32'hfe0d96a;
      116978: inst = 32'h5be00000;
      116979: inst = 32'h8c50000;
      116980: inst = 32'h24612800;
      116981: inst = 32'h10a00000;
      116982: inst = 32'hca0001c;
      116983: inst = 32'h24822800;
      116984: inst = 32'h10a00000;
      116985: inst = 32'hca00004;
      116986: inst = 32'h38632800;
      116987: inst = 32'h38842800;
      116988: inst = 32'h10a00001;
      116989: inst = 32'hca0c901;
      116990: inst = 32'h13e00001;
      116991: inst = 32'hfe0d96a;
      116992: inst = 32'h5be00000;
      116993: inst = 32'h8c50000;
      116994: inst = 32'h24612800;
      116995: inst = 32'h10a00000;
      116996: inst = 32'hca0001c;
      116997: inst = 32'h24822800;
      116998: inst = 32'h10a00000;
      116999: inst = 32'hca00004;
      117000: inst = 32'h38632800;
      117001: inst = 32'h38842800;
      117002: inst = 32'h10a00001;
      117003: inst = 32'hca0c90f;
      117004: inst = 32'h13e00001;
      117005: inst = 32'hfe0d96a;
      117006: inst = 32'h5be00000;
      117007: inst = 32'h8c50000;
      117008: inst = 32'h24612800;
      117009: inst = 32'h10a00000;
      117010: inst = 32'hca0001c;
      117011: inst = 32'h24822800;
      117012: inst = 32'h10a00000;
      117013: inst = 32'hca00004;
      117014: inst = 32'h38632800;
      117015: inst = 32'h38842800;
      117016: inst = 32'h10a00001;
      117017: inst = 32'hca0c91d;
      117018: inst = 32'h13e00001;
      117019: inst = 32'hfe0d96a;
      117020: inst = 32'h5be00000;
      117021: inst = 32'h8c50000;
      117022: inst = 32'h24612800;
      117023: inst = 32'h10a00000;
      117024: inst = 32'hca0001c;
      117025: inst = 32'h24822800;
      117026: inst = 32'h10a00000;
      117027: inst = 32'hca00004;
      117028: inst = 32'h38632800;
      117029: inst = 32'h38842800;
      117030: inst = 32'h10a00001;
      117031: inst = 32'hca0c92b;
      117032: inst = 32'h13e00001;
      117033: inst = 32'hfe0d96a;
      117034: inst = 32'h5be00000;
      117035: inst = 32'h8c50000;
      117036: inst = 32'h24612800;
      117037: inst = 32'h10a00000;
      117038: inst = 32'hca0001c;
      117039: inst = 32'h24822800;
      117040: inst = 32'h10a00000;
      117041: inst = 32'hca00004;
      117042: inst = 32'h38632800;
      117043: inst = 32'h38842800;
      117044: inst = 32'h10a00001;
      117045: inst = 32'hca0c939;
      117046: inst = 32'h13e00001;
      117047: inst = 32'hfe0d96a;
      117048: inst = 32'h5be00000;
      117049: inst = 32'h8c50000;
      117050: inst = 32'h24612800;
      117051: inst = 32'h10a00000;
      117052: inst = 32'hca0001c;
      117053: inst = 32'h24822800;
      117054: inst = 32'h10a00000;
      117055: inst = 32'hca00004;
      117056: inst = 32'h38632800;
      117057: inst = 32'h38842800;
      117058: inst = 32'h10a00001;
      117059: inst = 32'hca0c947;
      117060: inst = 32'h13e00001;
      117061: inst = 32'hfe0d96a;
      117062: inst = 32'h5be00000;
      117063: inst = 32'h8c50000;
      117064: inst = 32'h24612800;
      117065: inst = 32'h10a00000;
      117066: inst = 32'hca0001c;
      117067: inst = 32'h24822800;
      117068: inst = 32'h10a00000;
      117069: inst = 32'hca00004;
      117070: inst = 32'h38632800;
      117071: inst = 32'h38842800;
      117072: inst = 32'h10a00001;
      117073: inst = 32'hca0c955;
      117074: inst = 32'h13e00001;
      117075: inst = 32'hfe0d96a;
      117076: inst = 32'h5be00000;
      117077: inst = 32'h8c50000;
      117078: inst = 32'h24612800;
      117079: inst = 32'h10a00000;
      117080: inst = 32'hca0001c;
      117081: inst = 32'h24822800;
      117082: inst = 32'h10a00000;
      117083: inst = 32'hca00004;
      117084: inst = 32'h38632800;
      117085: inst = 32'h38842800;
      117086: inst = 32'h10a00001;
      117087: inst = 32'hca0c963;
      117088: inst = 32'h13e00001;
      117089: inst = 32'hfe0d96a;
      117090: inst = 32'h5be00000;
      117091: inst = 32'h8c50000;
      117092: inst = 32'h24612800;
      117093: inst = 32'h10a00000;
      117094: inst = 32'hca0001c;
      117095: inst = 32'h24822800;
      117096: inst = 32'h10a00000;
      117097: inst = 32'hca00004;
      117098: inst = 32'h38632800;
      117099: inst = 32'h38842800;
      117100: inst = 32'h10a00001;
      117101: inst = 32'hca0c971;
      117102: inst = 32'h13e00001;
      117103: inst = 32'hfe0d96a;
      117104: inst = 32'h5be00000;
      117105: inst = 32'h8c50000;
      117106: inst = 32'h24612800;
      117107: inst = 32'h10a00000;
      117108: inst = 32'hca0001c;
      117109: inst = 32'h24822800;
      117110: inst = 32'h10a00000;
      117111: inst = 32'hca00004;
      117112: inst = 32'h38632800;
      117113: inst = 32'h38842800;
      117114: inst = 32'h10a00001;
      117115: inst = 32'hca0c97f;
      117116: inst = 32'h13e00001;
      117117: inst = 32'hfe0d96a;
      117118: inst = 32'h5be00000;
      117119: inst = 32'h8c50000;
      117120: inst = 32'h24612800;
      117121: inst = 32'h10a00000;
      117122: inst = 32'hca0001c;
      117123: inst = 32'h24822800;
      117124: inst = 32'h10a00000;
      117125: inst = 32'hca00004;
      117126: inst = 32'h38632800;
      117127: inst = 32'h38842800;
      117128: inst = 32'h10a00001;
      117129: inst = 32'hca0c98d;
      117130: inst = 32'h13e00001;
      117131: inst = 32'hfe0d96a;
      117132: inst = 32'h5be00000;
      117133: inst = 32'h8c50000;
      117134: inst = 32'h24612800;
      117135: inst = 32'h10a00000;
      117136: inst = 32'hca0001c;
      117137: inst = 32'h24822800;
      117138: inst = 32'h10a00000;
      117139: inst = 32'hca00004;
      117140: inst = 32'h38632800;
      117141: inst = 32'h38842800;
      117142: inst = 32'h10a00001;
      117143: inst = 32'hca0c99b;
      117144: inst = 32'h13e00001;
      117145: inst = 32'hfe0d96a;
      117146: inst = 32'h5be00000;
      117147: inst = 32'h8c50000;
      117148: inst = 32'h24612800;
      117149: inst = 32'h10a00000;
      117150: inst = 32'hca0001c;
      117151: inst = 32'h24822800;
      117152: inst = 32'h10a00000;
      117153: inst = 32'hca00004;
      117154: inst = 32'h38632800;
      117155: inst = 32'h38842800;
      117156: inst = 32'h10a00001;
      117157: inst = 32'hca0c9a9;
      117158: inst = 32'h13e00001;
      117159: inst = 32'hfe0d96a;
      117160: inst = 32'h5be00000;
      117161: inst = 32'h8c50000;
      117162: inst = 32'h24612800;
      117163: inst = 32'h10a00000;
      117164: inst = 32'hca0001d;
      117165: inst = 32'h24822800;
      117166: inst = 32'h10a00000;
      117167: inst = 32'hca00004;
      117168: inst = 32'h38632800;
      117169: inst = 32'h38842800;
      117170: inst = 32'h10a00001;
      117171: inst = 32'hca0c9b7;
      117172: inst = 32'h13e00001;
      117173: inst = 32'hfe0d96a;
      117174: inst = 32'h5be00000;
      117175: inst = 32'h8c50000;
      117176: inst = 32'h24612800;
      117177: inst = 32'h10a00000;
      117178: inst = 32'hca0001d;
      117179: inst = 32'h24822800;
      117180: inst = 32'h10a00000;
      117181: inst = 32'hca00004;
      117182: inst = 32'h38632800;
      117183: inst = 32'h38842800;
      117184: inst = 32'h10a00001;
      117185: inst = 32'hca0c9c5;
      117186: inst = 32'h13e00001;
      117187: inst = 32'hfe0d96a;
      117188: inst = 32'h5be00000;
      117189: inst = 32'h8c50000;
      117190: inst = 32'h24612800;
      117191: inst = 32'h10a00000;
      117192: inst = 32'hca0001d;
      117193: inst = 32'h24822800;
      117194: inst = 32'h10a00000;
      117195: inst = 32'hca00004;
      117196: inst = 32'h38632800;
      117197: inst = 32'h38842800;
      117198: inst = 32'h10a00001;
      117199: inst = 32'hca0c9d3;
      117200: inst = 32'h13e00001;
      117201: inst = 32'hfe0d96a;
      117202: inst = 32'h5be00000;
      117203: inst = 32'h8c50000;
      117204: inst = 32'h24612800;
      117205: inst = 32'h10a00000;
      117206: inst = 32'hca0001d;
      117207: inst = 32'h24822800;
      117208: inst = 32'h10a00000;
      117209: inst = 32'hca00004;
      117210: inst = 32'h38632800;
      117211: inst = 32'h38842800;
      117212: inst = 32'h10a00001;
      117213: inst = 32'hca0c9e1;
      117214: inst = 32'h13e00001;
      117215: inst = 32'hfe0d96a;
      117216: inst = 32'h5be00000;
      117217: inst = 32'h8c50000;
      117218: inst = 32'h24612800;
      117219: inst = 32'h10a00000;
      117220: inst = 32'hca0001d;
      117221: inst = 32'h24822800;
      117222: inst = 32'h10a00000;
      117223: inst = 32'hca00004;
      117224: inst = 32'h38632800;
      117225: inst = 32'h38842800;
      117226: inst = 32'h10a00001;
      117227: inst = 32'hca0c9ef;
      117228: inst = 32'h13e00001;
      117229: inst = 32'hfe0d96a;
      117230: inst = 32'h5be00000;
      117231: inst = 32'h8c50000;
      117232: inst = 32'h24612800;
      117233: inst = 32'h10a00000;
      117234: inst = 32'hca0001d;
      117235: inst = 32'h24822800;
      117236: inst = 32'h10a00000;
      117237: inst = 32'hca00004;
      117238: inst = 32'h38632800;
      117239: inst = 32'h38842800;
      117240: inst = 32'h10a00001;
      117241: inst = 32'hca0c9fd;
      117242: inst = 32'h13e00001;
      117243: inst = 32'hfe0d96a;
      117244: inst = 32'h5be00000;
      117245: inst = 32'h8c50000;
      117246: inst = 32'h24612800;
      117247: inst = 32'h10a00000;
      117248: inst = 32'hca0001d;
      117249: inst = 32'h24822800;
      117250: inst = 32'h10a00000;
      117251: inst = 32'hca00004;
      117252: inst = 32'h38632800;
      117253: inst = 32'h38842800;
      117254: inst = 32'h10a00001;
      117255: inst = 32'hca0ca0b;
      117256: inst = 32'h13e00001;
      117257: inst = 32'hfe0d96a;
      117258: inst = 32'h5be00000;
      117259: inst = 32'h8c50000;
      117260: inst = 32'h24612800;
      117261: inst = 32'h10a00000;
      117262: inst = 32'hca0001d;
      117263: inst = 32'h24822800;
      117264: inst = 32'h10a00000;
      117265: inst = 32'hca00004;
      117266: inst = 32'h38632800;
      117267: inst = 32'h38842800;
      117268: inst = 32'h10a00001;
      117269: inst = 32'hca0ca19;
      117270: inst = 32'h13e00001;
      117271: inst = 32'hfe0d96a;
      117272: inst = 32'h5be00000;
      117273: inst = 32'h8c50000;
      117274: inst = 32'h24612800;
      117275: inst = 32'h10a00000;
      117276: inst = 32'hca0001d;
      117277: inst = 32'h24822800;
      117278: inst = 32'h10a00000;
      117279: inst = 32'hca00004;
      117280: inst = 32'h38632800;
      117281: inst = 32'h38842800;
      117282: inst = 32'h10a00001;
      117283: inst = 32'hca0ca27;
      117284: inst = 32'h13e00001;
      117285: inst = 32'hfe0d96a;
      117286: inst = 32'h5be00000;
      117287: inst = 32'h8c50000;
      117288: inst = 32'h24612800;
      117289: inst = 32'h10a00000;
      117290: inst = 32'hca0001d;
      117291: inst = 32'h24822800;
      117292: inst = 32'h10a00000;
      117293: inst = 32'hca00004;
      117294: inst = 32'h38632800;
      117295: inst = 32'h38842800;
      117296: inst = 32'h10a00001;
      117297: inst = 32'hca0ca35;
      117298: inst = 32'h13e00001;
      117299: inst = 32'hfe0d96a;
      117300: inst = 32'h5be00000;
      117301: inst = 32'h8c50000;
      117302: inst = 32'h24612800;
      117303: inst = 32'h10a00000;
      117304: inst = 32'hca0001d;
      117305: inst = 32'h24822800;
      117306: inst = 32'h10a00000;
      117307: inst = 32'hca00004;
      117308: inst = 32'h38632800;
      117309: inst = 32'h38842800;
      117310: inst = 32'h10a00001;
      117311: inst = 32'hca0ca43;
      117312: inst = 32'h13e00001;
      117313: inst = 32'hfe0d96a;
      117314: inst = 32'h5be00000;
      117315: inst = 32'h8c50000;
      117316: inst = 32'h24612800;
      117317: inst = 32'h10a00000;
      117318: inst = 32'hca0001d;
      117319: inst = 32'h24822800;
      117320: inst = 32'h10a00000;
      117321: inst = 32'hca00004;
      117322: inst = 32'h38632800;
      117323: inst = 32'h38842800;
      117324: inst = 32'h10a00001;
      117325: inst = 32'hca0ca51;
      117326: inst = 32'h13e00001;
      117327: inst = 32'hfe0d96a;
      117328: inst = 32'h5be00000;
      117329: inst = 32'h8c50000;
      117330: inst = 32'h24612800;
      117331: inst = 32'h10a00000;
      117332: inst = 32'hca0001d;
      117333: inst = 32'h24822800;
      117334: inst = 32'h10a00000;
      117335: inst = 32'hca00004;
      117336: inst = 32'h38632800;
      117337: inst = 32'h38842800;
      117338: inst = 32'h10a00001;
      117339: inst = 32'hca0ca5f;
      117340: inst = 32'h13e00001;
      117341: inst = 32'hfe0d96a;
      117342: inst = 32'h5be00000;
      117343: inst = 32'h8c50000;
      117344: inst = 32'h24612800;
      117345: inst = 32'h10a00000;
      117346: inst = 32'hca0001d;
      117347: inst = 32'h24822800;
      117348: inst = 32'h10a00000;
      117349: inst = 32'hca00004;
      117350: inst = 32'h38632800;
      117351: inst = 32'h38842800;
      117352: inst = 32'h10a00001;
      117353: inst = 32'hca0ca6d;
      117354: inst = 32'h13e00001;
      117355: inst = 32'hfe0d96a;
      117356: inst = 32'h5be00000;
      117357: inst = 32'h8c50000;
      117358: inst = 32'h24612800;
      117359: inst = 32'h10a00000;
      117360: inst = 32'hca0001d;
      117361: inst = 32'h24822800;
      117362: inst = 32'h10a00000;
      117363: inst = 32'hca00004;
      117364: inst = 32'h38632800;
      117365: inst = 32'h38842800;
      117366: inst = 32'h10a00001;
      117367: inst = 32'hca0ca7b;
      117368: inst = 32'h13e00001;
      117369: inst = 32'hfe0d96a;
      117370: inst = 32'h5be00000;
      117371: inst = 32'h8c50000;
      117372: inst = 32'h24612800;
      117373: inst = 32'h10a00000;
      117374: inst = 32'hca0001d;
      117375: inst = 32'h24822800;
      117376: inst = 32'h10a00000;
      117377: inst = 32'hca00004;
      117378: inst = 32'h38632800;
      117379: inst = 32'h38842800;
      117380: inst = 32'h10a00001;
      117381: inst = 32'hca0ca89;
      117382: inst = 32'h13e00001;
      117383: inst = 32'hfe0d96a;
      117384: inst = 32'h5be00000;
      117385: inst = 32'h8c50000;
      117386: inst = 32'h24612800;
      117387: inst = 32'h10a00000;
      117388: inst = 32'hca0001d;
      117389: inst = 32'h24822800;
      117390: inst = 32'h10a00000;
      117391: inst = 32'hca00004;
      117392: inst = 32'h38632800;
      117393: inst = 32'h38842800;
      117394: inst = 32'h10a00001;
      117395: inst = 32'hca0ca97;
      117396: inst = 32'h13e00001;
      117397: inst = 32'hfe0d96a;
      117398: inst = 32'h5be00000;
      117399: inst = 32'h8c50000;
      117400: inst = 32'h24612800;
      117401: inst = 32'h10a00000;
      117402: inst = 32'hca0001d;
      117403: inst = 32'h24822800;
      117404: inst = 32'h10a00000;
      117405: inst = 32'hca00004;
      117406: inst = 32'h38632800;
      117407: inst = 32'h38842800;
      117408: inst = 32'h10a00001;
      117409: inst = 32'hca0caa5;
      117410: inst = 32'h13e00001;
      117411: inst = 32'hfe0d96a;
      117412: inst = 32'h5be00000;
      117413: inst = 32'h8c50000;
      117414: inst = 32'h24612800;
      117415: inst = 32'h10a00000;
      117416: inst = 32'hca0001d;
      117417: inst = 32'h24822800;
      117418: inst = 32'h10a00000;
      117419: inst = 32'hca00004;
      117420: inst = 32'h38632800;
      117421: inst = 32'h38842800;
      117422: inst = 32'h10a00001;
      117423: inst = 32'hca0cab3;
      117424: inst = 32'h13e00001;
      117425: inst = 32'hfe0d96a;
      117426: inst = 32'h5be00000;
      117427: inst = 32'h8c50000;
      117428: inst = 32'h24612800;
      117429: inst = 32'h10a00000;
      117430: inst = 32'hca0001d;
      117431: inst = 32'h24822800;
      117432: inst = 32'h10a00000;
      117433: inst = 32'hca00004;
      117434: inst = 32'h38632800;
      117435: inst = 32'h38842800;
      117436: inst = 32'h10a00001;
      117437: inst = 32'hca0cac1;
      117438: inst = 32'h13e00001;
      117439: inst = 32'hfe0d96a;
      117440: inst = 32'h5be00000;
      117441: inst = 32'h8c50000;
      117442: inst = 32'h24612800;
      117443: inst = 32'h10a00000;
      117444: inst = 32'hca0001d;
      117445: inst = 32'h24822800;
      117446: inst = 32'h10a00000;
      117447: inst = 32'hca00004;
      117448: inst = 32'h38632800;
      117449: inst = 32'h38842800;
      117450: inst = 32'h10a00001;
      117451: inst = 32'hca0cacf;
      117452: inst = 32'h13e00001;
      117453: inst = 32'hfe0d96a;
      117454: inst = 32'h5be00000;
      117455: inst = 32'h8c50000;
      117456: inst = 32'h24612800;
      117457: inst = 32'h10a00000;
      117458: inst = 32'hca0001d;
      117459: inst = 32'h24822800;
      117460: inst = 32'h10a00000;
      117461: inst = 32'hca00004;
      117462: inst = 32'h38632800;
      117463: inst = 32'h38842800;
      117464: inst = 32'h10a00001;
      117465: inst = 32'hca0cadd;
      117466: inst = 32'h13e00001;
      117467: inst = 32'hfe0d96a;
      117468: inst = 32'h5be00000;
      117469: inst = 32'h8c50000;
      117470: inst = 32'h24612800;
      117471: inst = 32'h10a00000;
      117472: inst = 32'hca0001d;
      117473: inst = 32'h24822800;
      117474: inst = 32'h10a00000;
      117475: inst = 32'hca00004;
      117476: inst = 32'h38632800;
      117477: inst = 32'h38842800;
      117478: inst = 32'h10a00001;
      117479: inst = 32'hca0caeb;
      117480: inst = 32'h13e00001;
      117481: inst = 32'hfe0d96a;
      117482: inst = 32'h5be00000;
      117483: inst = 32'h8c50000;
      117484: inst = 32'h24612800;
      117485: inst = 32'h10a00000;
      117486: inst = 32'hca0001d;
      117487: inst = 32'h24822800;
      117488: inst = 32'h10a00000;
      117489: inst = 32'hca00004;
      117490: inst = 32'h38632800;
      117491: inst = 32'h38842800;
      117492: inst = 32'h10a00001;
      117493: inst = 32'hca0caf9;
      117494: inst = 32'h13e00001;
      117495: inst = 32'hfe0d96a;
      117496: inst = 32'h5be00000;
      117497: inst = 32'h8c50000;
      117498: inst = 32'h24612800;
      117499: inst = 32'h10a00000;
      117500: inst = 32'hca0001d;
      117501: inst = 32'h24822800;
      117502: inst = 32'h10a00000;
      117503: inst = 32'hca00004;
      117504: inst = 32'h38632800;
      117505: inst = 32'h38842800;
      117506: inst = 32'h10a00001;
      117507: inst = 32'hca0cb07;
      117508: inst = 32'h13e00001;
      117509: inst = 32'hfe0d96a;
      117510: inst = 32'h5be00000;
      117511: inst = 32'h8c50000;
      117512: inst = 32'h24612800;
      117513: inst = 32'h10a00000;
      117514: inst = 32'hca0001d;
      117515: inst = 32'h24822800;
      117516: inst = 32'h10a00000;
      117517: inst = 32'hca00004;
      117518: inst = 32'h38632800;
      117519: inst = 32'h38842800;
      117520: inst = 32'h10a00001;
      117521: inst = 32'hca0cb15;
      117522: inst = 32'h13e00001;
      117523: inst = 32'hfe0d96a;
      117524: inst = 32'h5be00000;
      117525: inst = 32'h8c50000;
      117526: inst = 32'h24612800;
      117527: inst = 32'h10a00000;
      117528: inst = 32'hca0001d;
      117529: inst = 32'h24822800;
      117530: inst = 32'h10a00000;
      117531: inst = 32'hca00004;
      117532: inst = 32'h38632800;
      117533: inst = 32'h38842800;
      117534: inst = 32'h10a00001;
      117535: inst = 32'hca0cb23;
      117536: inst = 32'h13e00001;
      117537: inst = 32'hfe0d96a;
      117538: inst = 32'h5be00000;
      117539: inst = 32'h8c50000;
      117540: inst = 32'h24612800;
      117541: inst = 32'h10a00000;
      117542: inst = 32'hca0001d;
      117543: inst = 32'h24822800;
      117544: inst = 32'h10a00000;
      117545: inst = 32'hca00004;
      117546: inst = 32'h38632800;
      117547: inst = 32'h38842800;
      117548: inst = 32'h10a00001;
      117549: inst = 32'hca0cb31;
      117550: inst = 32'h13e00001;
      117551: inst = 32'hfe0d96a;
      117552: inst = 32'h5be00000;
      117553: inst = 32'h8c50000;
      117554: inst = 32'h24612800;
      117555: inst = 32'h10a00000;
      117556: inst = 32'hca0001d;
      117557: inst = 32'h24822800;
      117558: inst = 32'h10a00000;
      117559: inst = 32'hca00004;
      117560: inst = 32'h38632800;
      117561: inst = 32'h38842800;
      117562: inst = 32'h10a00001;
      117563: inst = 32'hca0cb3f;
      117564: inst = 32'h13e00001;
      117565: inst = 32'hfe0d96a;
      117566: inst = 32'h5be00000;
      117567: inst = 32'h8c50000;
      117568: inst = 32'h24612800;
      117569: inst = 32'h10a00000;
      117570: inst = 32'hca0001d;
      117571: inst = 32'h24822800;
      117572: inst = 32'h10a00000;
      117573: inst = 32'hca00004;
      117574: inst = 32'h38632800;
      117575: inst = 32'h38842800;
      117576: inst = 32'h10a00001;
      117577: inst = 32'hca0cb4d;
      117578: inst = 32'h13e00001;
      117579: inst = 32'hfe0d96a;
      117580: inst = 32'h5be00000;
      117581: inst = 32'h8c50000;
      117582: inst = 32'h24612800;
      117583: inst = 32'h10a00000;
      117584: inst = 32'hca0001d;
      117585: inst = 32'h24822800;
      117586: inst = 32'h10a00000;
      117587: inst = 32'hca00004;
      117588: inst = 32'h38632800;
      117589: inst = 32'h38842800;
      117590: inst = 32'h10a00001;
      117591: inst = 32'hca0cb5b;
      117592: inst = 32'h13e00001;
      117593: inst = 32'hfe0d96a;
      117594: inst = 32'h5be00000;
      117595: inst = 32'h8c50000;
      117596: inst = 32'h24612800;
      117597: inst = 32'h10a00000;
      117598: inst = 32'hca0001d;
      117599: inst = 32'h24822800;
      117600: inst = 32'h10a00000;
      117601: inst = 32'hca00004;
      117602: inst = 32'h38632800;
      117603: inst = 32'h38842800;
      117604: inst = 32'h10a00001;
      117605: inst = 32'hca0cb69;
      117606: inst = 32'h13e00001;
      117607: inst = 32'hfe0d96a;
      117608: inst = 32'h5be00000;
      117609: inst = 32'h8c50000;
      117610: inst = 32'h24612800;
      117611: inst = 32'h10a00000;
      117612: inst = 32'hca0001d;
      117613: inst = 32'h24822800;
      117614: inst = 32'h10a00000;
      117615: inst = 32'hca00004;
      117616: inst = 32'h38632800;
      117617: inst = 32'h38842800;
      117618: inst = 32'h10a00001;
      117619: inst = 32'hca0cb77;
      117620: inst = 32'h13e00001;
      117621: inst = 32'hfe0d96a;
      117622: inst = 32'h5be00000;
      117623: inst = 32'h8c50000;
      117624: inst = 32'h24612800;
      117625: inst = 32'h10a00000;
      117626: inst = 32'hca0001d;
      117627: inst = 32'h24822800;
      117628: inst = 32'h10a00000;
      117629: inst = 32'hca00004;
      117630: inst = 32'h38632800;
      117631: inst = 32'h38842800;
      117632: inst = 32'h10a00001;
      117633: inst = 32'hca0cb85;
      117634: inst = 32'h13e00001;
      117635: inst = 32'hfe0d96a;
      117636: inst = 32'h5be00000;
      117637: inst = 32'h8c50000;
      117638: inst = 32'h24612800;
      117639: inst = 32'h10a00000;
      117640: inst = 32'hca0001d;
      117641: inst = 32'h24822800;
      117642: inst = 32'h10a00000;
      117643: inst = 32'hca00004;
      117644: inst = 32'h38632800;
      117645: inst = 32'h38842800;
      117646: inst = 32'h10a00001;
      117647: inst = 32'hca0cb93;
      117648: inst = 32'h13e00001;
      117649: inst = 32'hfe0d96a;
      117650: inst = 32'h5be00000;
      117651: inst = 32'h8c50000;
      117652: inst = 32'h24612800;
      117653: inst = 32'h10a00000;
      117654: inst = 32'hca0001d;
      117655: inst = 32'h24822800;
      117656: inst = 32'h10a00000;
      117657: inst = 32'hca00004;
      117658: inst = 32'h38632800;
      117659: inst = 32'h38842800;
      117660: inst = 32'h10a00001;
      117661: inst = 32'hca0cba1;
      117662: inst = 32'h13e00001;
      117663: inst = 32'hfe0d96a;
      117664: inst = 32'h5be00000;
      117665: inst = 32'h8c50000;
      117666: inst = 32'h24612800;
      117667: inst = 32'h10a00000;
      117668: inst = 32'hca0001d;
      117669: inst = 32'h24822800;
      117670: inst = 32'h10a00000;
      117671: inst = 32'hca00004;
      117672: inst = 32'h38632800;
      117673: inst = 32'h38842800;
      117674: inst = 32'h10a00001;
      117675: inst = 32'hca0cbaf;
      117676: inst = 32'h13e00001;
      117677: inst = 32'hfe0d96a;
      117678: inst = 32'h5be00000;
      117679: inst = 32'h8c50000;
      117680: inst = 32'h24612800;
      117681: inst = 32'h10a00000;
      117682: inst = 32'hca0001d;
      117683: inst = 32'h24822800;
      117684: inst = 32'h10a00000;
      117685: inst = 32'hca00004;
      117686: inst = 32'h38632800;
      117687: inst = 32'h38842800;
      117688: inst = 32'h10a00001;
      117689: inst = 32'hca0cbbd;
      117690: inst = 32'h13e00001;
      117691: inst = 32'hfe0d96a;
      117692: inst = 32'h5be00000;
      117693: inst = 32'h8c50000;
      117694: inst = 32'h24612800;
      117695: inst = 32'h10a00000;
      117696: inst = 32'hca0001d;
      117697: inst = 32'h24822800;
      117698: inst = 32'h10a00000;
      117699: inst = 32'hca00004;
      117700: inst = 32'h38632800;
      117701: inst = 32'h38842800;
      117702: inst = 32'h10a00001;
      117703: inst = 32'hca0cbcb;
      117704: inst = 32'h13e00001;
      117705: inst = 32'hfe0d96a;
      117706: inst = 32'h5be00000;
      117707: inst = 32'h8c50000;
      117708: inst = 32'h24612800;
      117709: inst = 32'h10a00000;
      117710: inst = 32'hca0001d;
      117711: inst = 32'h24822800;
      117712: inst = 32'h10a00000;
      117713: inst = 32'hca00004;
      117714: inst = 32'h38632800;
      117715: inst = 32'h38842800;
      117716: inst = 32'h10a00001;
      117717: inst = 32'hca0cbd9;
      117718: inst = 32'h13e00001;
      117719: inst = 32'hfe0d96a;
      117720: inst = 32'h5be00000;
      117721: inst = 32'h8c50000;
      117722: inst = 32'h24612800;
      117723: inst = 32'h10a00000;
      117724: inst = 32'hca0001d;
      117725: inst = 32'h24822800;
      117726: inst = 32'h10a00000;
      117727: inst = 32'hca00004;
      117728: inst = 32'h38632800;
      117729: inst = 32'h38842800;
      117730: inst = 32'h10a00001;
      117731: inst = 32'hca0cbe7;
      117732: inst = 32'h13e00001;
      117733: inst = 32'hfe0d96a;
      117734: inst = 32'h5be00000;
      117735: inst = 32'h8c50000;
      117736: inst = 32'h24612800;
      117737: inst = 32'h10a00000;
      117738: inst = 32'hca0001d;
      117739: inst = 32'h24822800;
      117740: inst = 32'h10a00000;
      117741: inst = 32'hca00004;
      117742: inst = 32'h38632800;
      117743: inst = 32'h38842800;
      117744: inst = 32'h10a00001;
      117745: inst = 32'hca0cbf5;
      117746: inst = 32'h13e00001;
      117747: inst = 32'hfe0d96a;
      117748: inst = 32'h5be00000;
      117749: inst = 32'h8c50000;
      117750: inst = 32'h24612800;
      117751: inst = 32'h10a00000;
      117752: inst = 32'hca0001d;
      117753: inst = 32'h24822800;
      117754: inst = 32'h10a00000;
      117755: inst = 32'hca00004;
      117756: inst = 32'h38632800;
      117757: inst = 32'h38842800;
      117758: inst = 32'h10a00001;
      117759: inst = 32'hca0cc03;
      117760: inst = 32'h13e00001;
      117761: inst = 32'hfe0d96a;
      117762: inst = 32'h5be00000;
      117763: inst = 32'h8c50000;
      117764: inst = 32'h24612800;
      117765: inst = 32'h10a00000;
      117766: inst = 32'hca0001d;
      117767: inst = 32'h24822800;
      117768: inst = 32'h10a00000;
      117769: inst = 32'hca00004;
      117770: inst = 32'h38632800;
      117771: inst = 32'h38842800;
      117772: inst = 32'h10a00001;
      117773: inst = 32'hca0cc11;
      117774: inst = 32'h13e00001;
      117775: inst = 32'hfe0d96a;
      117776: inst = 32'h5be00000;
      117777: inst = 32'h8c50000;
      117778: inst = 32'h24612800;
      117779: inst = 32'h10a00000;
      117780: inst = 32'hca0001d;
      117781: inst = 32'h24822800;
      117782: inst = 32'h10a00000;
      117783: inst = 32'hca00004;
      117784: inst = 32'h38632800;
      117785: inst = 32'h38842800;
      117786: inst = 32'h10a00001;
      117787: inst = 32'hca0cc1f;
      117788: inst = 32'h13e00001;
      117789: inst = 32'hfe0d96a;
      117790: inst = 32'h5be00000;
      117791: inst = 32'h8c50000;
      117792: inst = 32'h24612800;
      117793: inst = 32'h10a00000;
      117794: inst = 32'hca0001d;
      117795: inst = 32'h24822800;
      117796: inst = 32'h10a00000;
      117797: inst = 32'hca00004;
      117798: inst = 32'h38632800;
      117799: inst = 32'h38842800;
      117800: inst = 32'h10a00001;
      117801: inst = 32'hca0cc2d;
      117802: inst = 32'h13e00001;
      117803: inst = 32'hfe0d96a;
      117804: inst = 32'h5be00000;
      117805: inst = 32'h8c50000;
      117806: inst = 32'h24612800;
      117807: inst = 32'h10a00000;
      117808: inst = 32'hca0001d;
      117809: inst = 32'h24822800;
      117810: inst = 32'h10a00000;
      117811: inst = 32'hca00004;
      117812: inst = 32'h38632800;
      117813: inst = 32'h38842800;
      117814: inst = 32'h10a00001;
      117815: inst = 32'hca0cc3b;
      117816: inst = 32'h13e00001;
      117817: inst = 32'hfe0d96a;
      117818: inst = 32'h5be00000;
      117819: inst = 32'h8c50000;
      117820: inst = 32'h24612800;
      117821: inst = 32'h10a00000;
      117822: inst = 32'hca0001d;
      117823: inst = 32'h24822800;
      117824: inst = 32'h10a00000;
      117825: inst = 32'hca00004;
      117826: inst = 32'h38632800;
      117827: inst = 32'h38842800;
      117828: inst = 32'h10a00001;
      117829: inst = 32'hca0cc49;
      117830: inst = 32'h13e00001;
      117831: inst = 32'hfe0d96a;
      117832: inst = 32'h5be00000;
      117833: inst = 32'h8c50000;
      117834: inst = 32'h24612800;
      117835: inst = 32'h10a00000;
      117836: inst = 32'hca0001d;
      117837: inst = 32'h24822800;
      117838: inst = 32'h10a00000;
      117839: inst = 32'hca00004;
      117840: inst = 32'h38632800;
      117841: inst = 32'h38842800;
      117842: inst = 32'h10a00001;
      117843: inst = 32'hca0cc57;
      117844: inst = 32'h13e00001;
      117845: inst = 32'hfe0d96a;
      117846: inst = 32'h5be00000;
      117847: inst = 32'h8c50000;
      117848: inst = 32'h24612800;
      117849: inst = 32'h10a00000;
      117850: inst = 32'hca0001d;
      117851: inst = 32'h24822800;
      117852: inst = 32'h10a00000;
      117853: inst = 32'hca00004;
      117854: inst = 32'h38632800;
      117855: inst = 32'h38842800;
      117856: inst = 32'h10a00001;
      117857: inst = 32'hca0cc65;
      117858: inst = 32'h13e00001;
      117859: inst = 32'hfe0d96a;
      117860: inst = 32'h5be00000;
      117861: inst = 32'h8c50000;
      117862: inst = 32'h24612800;
      117863: inst = 32'h10a00000;
      117864: inst = 32'hca0001d;
      117865: inst = 32'h24822800;
      117866: inst = 32'h10a00000;
      117867: inst = 32'hca00004;
      117868: inst = 32'h38632800;
      117869: inst = 32'h38842800;
      117870: inst = 32'h10a00001;
      117871: inst = 32'hca0cc73;
      117872: inst = 32'h13e00001;
      117873: inst = 32'hfe0d96a;
      117874: inst = 32'h5be00000;
      117875: inst = 32'h8c50000;
      117876: inst = 32'h24612800;
      117877: inst = 32'h10a00000;
      117878: inst = 32'hca0001d;
      117879: inst = 32'h24822800;
      117880: inst = 32'h10a00000;
      117881: inst = 32'hca00004;
      117882: inst = 32'h38632800;
      117883: inst = 32'h38842800;
      117884: inst = 32'h10a00001;
      117885: inst = 32'hca0cc81;
      117886: inst = 32'h13e00001;
      117887: inst = 32'hfe0d96a;
      117888: inst = 32'h5be00000;
      117889: inst = 32'h8c50000;
      117890: inst = 32'h24612800;
      117891: inst = 32'h10a00000;
      117892: inst = 32'hca0001d;
      117893: inst = 32'h24822800;
      117894: inst = 32'h10a00000;
      117895: inst = 32'hca00004;
      117896: inst = 32'h38632800;
      117897: inst = 32'h38842800;
      117898: inst = 32'h10a00001;
      117899: inst = 32'hca0cc8f;
      117900: inst = 32'h13e00001;
      117901: inst = 32'hfe0d96a;
      117902: inst = 32'h5be00000;
      117903: inst = 32'h8c50000;
      117904: inst = 32'h24612800;
      117905: inst = 32'h10a00000;
      117906: inst = 32'hca0001d;
      117907: inst = 32'h24822800;
      117908: inst = 32'h10a00000;
      117909: inst = 32'hca00004;
      117910: inst = 32'h38632800;
      117911: inst = 32'h38842800;
      117912: inst = 32'h10a00001;
      117913: inst = 32'hca0cc9d;
      117914: inst = 32'h13e00001;
      117915: inst = 32'hfe0d96a;
      117916: inst = 32'h5be00000;
      117917: inst = 32'h8c50000;
      117918: inst = 32'h24612800;
      117919: inst = 32'h10a00000;
      117920: inst = 32'hca0001d;
      117921: inst = 32'h24822800;
      117922: inst = 32'h10a00000;
      117923: inst = 32'hca00004;
      117924: inst = 32'h38632800;
      117925: inst = 32'h38842800;
      117926: inst = 32'h10a00001;
      117927: inst = 32'hca0ccab;
      117928: inst = 32'h13e00001;
      117929: inst = 32'hfe0d96a;
      117930: inst = 32'h5be00000;
      117931: inst = 32'h8c50000;
      117932: inst = 32'h24612800;
      117933: inst = 32'h10a00000;
      117934: inst = 32'hca0001d;
      117935: inst = 32'h24822800;
      117936: inst = 32'h10a00000;
      117937: inst = 32'hca00004;
      117938: inst = 32'h38632800;
      117939: inst = 32'h38842800;
      117940: inst = 32'h10a00001;
      117941: inst = 32'hca0ccb9;
      117942: inst = 32'h13e00001;
      117943: inst = 32'hfe0d96a;
      117944: inst = 32'h5be00000;
      117945: inst = 32'h8c50000;
      117946: inst = 32'h24612800;
      117947: inst = 32'h10a00000;
      117948: inst = 32'hca0001d;
      117949: inst = 32'h24822800;
      117950: inst = 32'h10a00000;
      117951: inst = 32'hca00004;
      117952: inst = 32'h38632800;
      117953: inst = 32'h38842800;
      117954: inst = 32'h10a00001;
      117955: inst = 32'hca0ccc7;
      117956: inst = 32'h13e00001;
      117957: inst = 32'hfe0d96a;
      117958: inst = 32'h5be00000;
      117959: inst = 32'h8c50000;
      117960: inst = 32'h24612800;
      117961: inst = 32'h10a00000;
      117962: inst = 32'hca0001d;
      117963: inst = 32'h24822800;
      117964: inst = 32'h10a00000;
      117965: inst = 32'hca00004;
      117966: inst = 32'h38632800;
      117967: inst = 32'h38842800;
      117968: inst = 32'h10a00001;
      117969: inst = 32'hca0ccd5;
      117970: inst = 32'h13e00001;
      117971: inst = 32'hfe0d96a;
      117972: inst = 32'h5be00000;
      117973: inst = 32'h8c50000;
      117974: inst = 32'h24612800;
      117975: inst = 32'h10a00000;
      117976: inst = 32'hca0001d;
      117977: inst = 32'h24822800;
      117978: inst = 32'h10a00000;
      117979: inst = 32'hca00004;
      117980: inst = 32'h38632800;
      117981: inst = 32'h38842800;
      117982: inst = 32'h10a00001;
      117983: inst = 32'hca0cce3;
      117984: inst = 32'h13e00001;
      117985: inst = 32'hfe0d96a;
      117986: inst = 32'h5be00000;
      117987: inst = 32'h8c50000;
      117988: inst = 32'h24612800;
      117989: inst = 32'h10a00000;
      117990: inst = 32'hca0001d;
      117991: inst = 32'h24822800;
      117992: inst = 32'h10a00000;
      117993: inst = 32'hca00004;
      117994: inst = 32'h38632800;
      117995: inst = 32'h38842800;
      117996: inst = 32'h10a00001;
      117997: inst = 32'hca0ccf1;
      117998: inst = 32'h13e00001;
      117999: inst = 32'hfe0d96a;
      118000: inst = 32'h5be00000;
      118001: inst = 32'h8c50000;
      118002: inst = 32'h24612800;
      118003: inst = 32'h10a00000;
      118004: inst = 32'hca0001d;
      118005: inst = 32'h24822800;
      118006: inst = 32'h10a00000;
      118007: inst = 32'hca00004;
      118008: inst = 32'h38632800;
      118009: inst = 32'h38842800;
      118010: inst = 32'h10a00001;
      118011: inst = 32'hca0ccff;
      118012: inst = 32'h13e00001;
      118013: inst = 32'hfe0d96a;
      118014: inst = 32'h5be00000;
      118015: inst = 32'h8c50000;
      118016: inst = 32'h24612800;
      118017: inst = 32'h10a00000;
      118018: inst = 32'hca0001d;
      118019: inst = 32'h24822800;
      118020: inst = 32'h10a00000;
      118021: inst = 32'hca00004;
      118022: inst = 32'h38632800;
      118023: inst = 32'h38842800;
      118024: inst = 32'h10a00001;
      118025: inst = 32'hca0cd0d;
      118026: inst = 32'h13e00001;
      118027: inst = 32'hfe0d96a;
      118028: inst = 32'h5be00000;
      118029: inst = 32'h8c50000;
      118030: inst = 32'h24612800;
      118031: inst = 32'h10a00000;
      118032: inst = 32'hca0001d;
      118033: inst = 32'h24822800;
      118034: inst = 32'h10a00000;
      118035: inst = 32'hca00004;
      118036: inst = 32'h38632800;
      118037: inst = 32'h38842800;
      118038: inst = 32'h10a00001;
      118039: inst = 32'hca0cd1b;
      118040: inst = 32'h13e00001;
      118041: inst = 32'hfe0d96a;
      118042: inst = 32'h5be00000;
      118043: inst = 32'h8c50000;
      118044: inst = 32'h24612800;
      118045: inst = 32'h10a00000;
      118046: inst = 32'hca0001d;
      118047: inst = 32'h24822800;
      118048: inst = 32'h10a00000;
      118049: inst = 32'hca00004;
      118050: inst = 32'h38632800;
      118051: inst = 32'h38842800;
      118052: inst = 32'h10a00001;
      118053: inst = 32'hca0cd29;
      118054: inst = 32'h13e00001;
      118055: inst = 32'hfe0d96a;
      118056: inst = 32'h5be00000;
      118057: inst = 32'h8c50000;
      118058: inst = 32'h24612800;
      118059: inst = 32'h10a00000;
      118060: inst = 32'hca0001d;
      118061: inst = 32'h24822800;
      118062: inst = 32'h10a00000;
      118063: inst = 32'hca00004;
      118064: inst = 32'h38632800;
      118065: inst = 32'h38842800;
      118066: inst = 32'h10a00001;
      118067: inst = 32'hca0cd37;
      118068: inst = 32'h13e00001;
      118069: inst = 32'hfe0d96a;
      118070: inst = 32'h5be00000;
      118071: inst = 32'h8c50000;
      118072: inst = 32'h24612800;
      118073: inst = 32'h10a00000;
      118074: inst = 32'hca0001d;
      118075: inst = 32'h24822800;
      118076: inst = 32'h10a00000;
      118077: inst = 32'hca00004;
      118078: inst = 32'h38632800;
      118079: inst = 32'h38842800;
      118080: inst = 32'h10a00001;
      118081: inst = 32'hca0cd45;
      118082: inst = 32'h13e00001;
      118083: inst = 32'hfe0d96a;
      118084: inst = 32'h5be00000;
      118085: inst = 32'h8c50000;
      118086: inst = 32'h24612800;
      118087: inst = 32'h10a00000;
      118088: inst = 32'hca0001d;
      118089: inst = 32'h24822800;
      118090: inst = 32'h10a00000;
      118091: inst = 32'hca00004;
      118092: inst = 32'h38632800;
      118093: inst = 32'h38842800;
      118094: inst = 32'h10a00001;
      118095: inst = 32'hca0cd53;
      118096: inst = 32'h13e00001;
      118097: inst = 32'hfe0d96a;
      118098: inst = 32'h5be00000;
      118099: inst = 32'h8c50000;
      118100: inst = 32'h24612800;
      118101: inst = 32'h10a00000;
      118102: inst = 32'hca0001d;
      118103: inst = 32'h24822800;
      118104: inst = 32'h10a00000;
      118105: inst = 32'hca00004;
      118106: inst = 32'h38632800;
      118107: inst = 32'h38842800;
      118108: inst = 32'h10a00001;
      118109: inst = 32'hca0cd61;
      118110: inst = 32'h13e00001;
      118111: inst = 32'hfe0d96a;
      118112: inst = 32'h5be00000;
      118113: inst = 32'h8c50000;
      118114: inst = 32'h24612800;
      118115: inst = 32'h10a00000;
      118116: inst = 32'hca0001d;
      118117: inst = 32'h24822800;
      118118: inst = 32'h10a00000;
      118119: inst = 32'hca00004;
      118120: inst = 32'h38632800;
      118121: inst = 32'h38842800;
      118122: inst = 32'h10a00001;
      118123: inst = 32'hca0cd6f;
      118124: inst = 32'h13e00001;
      118125: inst = 32'hfe0d96a;
      118126: inst = 32'h5be00000;
      118127: inst = 32'h8c50000;
      118128: inst = 32'h24612800;
      118129: inst = 32'h10a00000;
      118130: inst = 32'hca0001d;
      118131: inst = 32'h24822800;
      118132: inst = 32'h10a00000;
      118133: inst = 32'hca00004;
      118134: inst = 32'h38632800;
      118135: inst = 32'h38842800;
      118136: inst = 32'h10a00001;
      118137: inst = 32'hca0cd7d;
      118138: inst = 32'h13e00001;
      118139: inst = 32'hfe0d96a;
      118140: inst = 32'h5be00000;
      118141: inst = 32'h8c50000;
      118142: inst = 32'h24612800;
      118143: inst = 32'h10a00000;
      118144: inst = 32'hca0001d;
      118145: inst = 32'h24822800;
      118146: inst = 32'h10a00000;
      118147: inst = 32'hca00004;
      118148: inst = 32'h38632800;
      118149: inst = 32'h38842800;
      118150: inst = 32'h10a00001;
      118151: inst = 32'hca0cd8b;
      118152: inst = 32'h13e00001;
      118153: inst = 32'hfe0d96a;
      118154: inst = 32'h5be00000;
      118155: inst = 32'h8c50000;
      118156: inst = 32'h24612800;
      118157: inst = 32'h10a00000;
      118158: inst = 32'hca0001d;
      118159: inst = 32'h24822800;
      118160: inst = 32'h10a00000;
      118161: inst = 32'hca00004;
      118162: inst = 32'h38632800;
      118163: inst = 32'h38842800;
      118164: inst = 32'h10a00001;
      118165: inst = 32'hca0cd99;
      118166: inst = 32'h13e00001;
      118167: inst = 32'hfe0d96a;
      118168: inst = 32'h5be00000;
      118169: inst = 32'h8c50000;
      118170: inst = 32'h24612800;
      118171: inst = 32'h10a00000;
      118172: inst = 32'hca0001d;
      118173: inst = 32'h24822800;
      118174: inst = 32'h10a00000;
      118175: inst = 32'hca00004;
      118176: inst = 32'h38632800;
      118177: inst = 32'h38842800;
      118178: inst = 32'h10a00001;
      118179: inst = 32'hca0cda7;
      118180: inst = 32'h13e00001;
      118181: inst = 32'hfe0d96a;
      118182: inst = 32'h5be00000;
      118183: inst = 32'h8c50000;
      118184: inst = 32'h24612800;
      118185: inst = 32'h10a00000;
      118186: inst = 32'hca0001d;
      118187: inst = 32'h24822800;
      118188: inst = 32'h10a00000;
      118189: inst = 32'hca00004;
      118190: inst = 32'h38632800;
      118191: inst = 32'h38842800;
      118192: inst = 32'h10a00001;
      118193: inst = 32'hca0cdb5;
      118194: inst = 32'h13e00001;
      118195: inst = 32'hfe0d96a;
      118196: inst = 32'h5be00000;
      118197: inst = 32'h8c50000;
      118198: inst = 32'h24612800;
      118199: inst = 32'h10a00000;
      118200: inst = 32'hca0001d;
      118201: inst = 32'h24822800;
      118202: inst = 32'h10a00000;
      118203: inst = 32'hca00004;
      118204: inst = 32'h38632800;
      118205: inst = 32'h38842800;
      118206: inst = 32'h10a00001;
      118207: inst = 32'hca0cdc3;
      118208: inst = 32'h13e00001;
      118209: inst = 32'hfe0d96a;
      118210: inst = 32'h5be00000;
      118211: inst = 32'h8c50000;
      118212: inst = 32'h24612800;
      118213: inst = 32'h10a00000;
      118214: inst = 32'hca0001d;
      118215: inst = 32'h24822800;
      118216: inst = 32'h10a00000;
      118217: inst = 32'hca00004;
      118218: inst = 32'h38632800;
      118219: inst = 32'h38842800;
      118220: inst = 32'h10a00001;
      118221: inst = 32'hca0cdd1;
      118222: inst = 32'h13e00001;
      118223: inst = 32'hfe0d96a;
      118224: inst = 32'h5be00000;
      118225: inst = 32'h8c50000;
      118226: inst = 32'h24612800;
      118227: inst = 32'h10a00000;
      118228: inst = 32'hca0001d;
      118229: inst = 32'h24822800;
      118230: inst = 32'h10a00000;
      118231: inst = 32'hca00004;
      118232: inst = 32'h38632800;
      118233: inst = 32'h38842800;
      118234: inst = 32'h10a00001;
      118235: inst = 32'hca0cddf;
      118236: inst = 32'h13e00001;
      118237: inst = 32'hfe0d96a;
      118238: inst = 32'h5be00000;
      118239: inst = 32'h8c50000;
      118240: inst = 32'h24612800;
      118241: inst = 32'h10a00000;
      118242: inst = 32'hca0001d;
      118243: inst = 32'h24822800;
      118244: inst = 32'h10a00000;
      118245: inst = 32'hca00004;
      118246: inst = 32'h38632800;
      118247: inst = 32'h38842800;
      118248: inst = 32'h10a00001;
      118249: inst = 32'hca0cded;
      118250: inst = 32'h13e00001;
      118251: inst = 32'hfe0d96a;
      118252: inst = 32'h5be00000;
      118253: inst = 32'h8c50000;
      118254: inst = 32'h24612800;
      118255: inst = 32'h10a00000;
      118256: inst = 32'hca0001d;
      118257: inst = 32'h24822800;
      118258: inst = 32'h10a00000;
      118259: inst = 32'hca00004;
      118260: inst = 32'h38632800;
      118261: inst = 32'h38842800;
      118262: inst = 32'h10a00001;
      118263: inst = 32'hca0cdfb;
      118264: inst = 32'h13e00001;
      118265: inst = 32'hfe0d96a;
      118266: inst = 32'h5be00000;
      118267: inst = 32'h8c50000;
      118268: inst = 32'h24612800;
      118269: inst = 32'h10a00000;
      118270: inst = 32'hca0001d;
      118271: inst = 32'h24822800;
      118272: inst = 32'h10a00000;
      118273: inst = 32'hca00004;
      118274: inst = 32'h38632800;
      118275: inst = 32'h38842800;
      118276: inst = 32'h10a00001;
      118277: inst = 32'hca0ce09;
      118278: inst = 32'h13e00001;
      118279: inst = 32'hfe0d96a;
      118280: inst = 32'h5be00000;
      118281: inst = 32'h8c50000;
      118282: inst = 32'h24612800;
      118283: inst = 32'h10a00000;
      118284: inst = 32'hca0001d;
      118285: inst = 32'h24822800;
      118286: inst = 32'h10a00000;
      118287: inst = 32'hca00004;
      118288: inst = 32'h38632800;
      118289: inst = 32'h38842800;
      118290: inst = 32'h10a00001;
      118291: inst = 32'hca0ce17;
      118292: inst = 32'h13e00001;
      118293: inst = 32'hfe0d96a;
      118294: inst = 32'h5be00000;
      118295: inst = 32'h8c50000;
      118296: inst = 32'h24612800;
      118297: inst = 32'h10a00000;
      118298: inst = 32'hca0001d;
      118299: inst = 32'h24822800;
      118300: inst = 32'h10a00000;
      118301: inst = 32'hca00004;
      118302: inst = 32'h38632800;
      118303: inst = 32'h38842800;
      118304: inst = 32'h10a00001;
      118305: inst = 32'hca0ce25;
      118306: inst = 32'h13e00001;
      118307: inst = 32'hfe0d96a;
      118308: inst = 32'h5be00000;
      118309: inst = 32'h8c50000;
      118310: inst = 32'h24612800;
      118311: inst = 32'h10a00000;
      118312: inst = 32'hca0001d;
      118313: inst = 32'h24822800;
      118314: inst = 32'h10a00000;
      118315: inst = 32'hca00004;
      118316: inst = 32'h38632800;
      118317: inst = 32'h38842800;
      118318: inst = 32'h10a00001;
      118319: inst = 32'hca0ce33;
      118320: inst = 32'h13e00001;
      118321: inst = 32'hfe0d96a;
      118322: inst = 32'h5be00000;
      118323: inst = 32'h8c50000;
      118324: inst = 32'h24612800;
      118325: inst = 32'h10a00000;
      118326: inst = 32'hca0001d;
      118327: inst = 32'h24822800;
      118328: inst = 32'h10a00000;
      118329: inst = 32'hca00004;
      118330: inst = 32'h38632800;
      118331: inst = 32'h38842800;
      118332: inst = 32'h10a00001;
      118333: inst = 32'hca0ce41;
      118334: inst = 32'h13e00001;
      118335: inst = 32'hfe0d96a;
      118336: inst = 32'h5be00000;
      118337: inst = 32'h8c50000;
      118338: inst = 32'h24612800;
      118339: inst = 32'h10a00000;
      118340: inst = 32'hca0001d;
      118341: inst = 32'h24822800;
      118342: inst = 32'h10a00000;
      118343: inst = 32'hca00004;
      118344: inst = 32'h38632800;
      118345: inst = 32'h38842800;
      118346: inst = 32'h10a00001;
      118347: inst = 32'hca0ce4f;
      118348: inst = 32'h13e00001;
      118349: inst = 32'hfe0d96a;
      118350: inst = 32'h5be00000;
      118351: inst = 32'h8c50000;
      118352: inst = 32'h24612800;
      118353: inst = 32'h10a00000;
      118354: inst = 32'hca0001d;
      118355: inst = 32'h24822800;
      118356: inst = 32'h10a00000;
      118357: inst = 32'hca00004;
      118358: inst = 32'h38632800;
      118359: inst = 32'h38842800;
      118360: inst = 32'h10a00001;
      118361: inst = 32'hca0ce5d;
      118362: inst = 32'h13e00001;
      118363: inst = 32'hfe0d96a;
      118364: inst = 32'h5be00000;
      118365: inst = 32'h8c50000;
      118366: inst = 32'h24612800;
      118367: inst = 32'h10a00000;
      118368: inst = 32'hca0001d;
      118369: inst = 32'h24822800;
      118370: inst = 32'h10a00000;
      118371: inst = 32'hca00004;
      118372: inst = 32'h38632800;
      118373: inst = 32'h38842800;
      118374: inst = 32'h10a00001;
      118375: inst = 32'hca0ce6b;
      118376: inst = 32'h13e00001;
      118377: inst = 32'hfe0d96a;
      118378: inst = 32'h5be00000;
      118379: inst = 32'h8c50000;
      118380: inst = 32'h24612800;
      118381: inst = 32'h10a00000;
      118382: inst = 32'hca0001d;
      118383: inst = 32'h24822800;
      118384: inst = 32'h10a00000;
      118385: inst = 32'hca00004;
      118386: inst = 32'h38632800;
      118387: inst = 32'h38842800;
      118388: inst = 32'h10a00001;
      118389: inst = 32'hca0ce79;
      118390: inst = 32'h13e00001;
      118391: inst = 32'hfe0d96a;
      118392: inst = 32'h5be00000;
      118393: inst = 32'h8c50000;
      118394: inst = 32'h24612800;
      118395: inst = 32'h10a00000;
      118396: inst = 32'hca0001d;
      118397: inst = 32'h24822800;
      118398: inst = 32'h10a00000;
      118399: inst = 32'hca00004;
      118400: inst = 32'h38632800;
      118401: inst = 32'h38842800;
      118402: inst = 32'h10a00001;
      118403: inst = 32'hca0ce87;
      118404: inst = 32'h13e00001;
      118405: inst = 32'hfe0d96a;
      118406: inst = 32'h5be00000;
      118407: inst = 32'h8c50000;
      118408: inst = 32'h24612800;
      118409: inst = 32'h10a00000;
      118410: inst = 32'hca0001d;
      118411: inst = 32'h24822800;
      118412: inst = 32'h10a00000;
      118413: inst = 32'hca00004;
      118414: inst = 32'h38632800;
      118415: inst = 32'h38842800;
      118416: inst = 32'h10a00001;
      118417: inst = 32'hca0ce95;
      118418: inst = 32'h13e00001;
      118419: inst = 32'hfe0d96a;
      118420: inst = 32'h5be00000;
      118421: inst = 32'h8c50000;
      118422: inst = 32'h24612800;
      118423: inst = 32'h10a00000;
      118424: inst = 32'hca0001d;
      118425: inst = 32'h24822800;
      118426: inst = 32'h10a00000;
      118427: inst = 32'hca00004;
      118428: inst = 32'h38632800;
      118429: inst = 32'h38842800;
      118430: inst = 32'h10a00001;
      118431: inst = 32'hca0cea3;
      118432: inst = 32'h13e00001;
      118433: inst = 32'hfe0d96a;
      118434: inst = 32'h5be00000;
      118435: inst = 32'h8c50000;
      118436: inst = 32'h24612800;
      118437: inst = 32'h10a00000;
      118438: inst = 32'hca0001d;
      118439: inst = 32'h24822800;
      118440: inst = 32'h10a00000;
      118441: inst = 32'hca00004;
      118442: inst = 32'h38632800;
      118443: inst = 32'h38842800;
      118444: inst = 32'h10a00001;
      118445: inst = 32'hca0ceb1;
      118446: inst = 32'h13e00001;
      118447: inst = 32'hfe0d96a;
      118448: inst = 32'h5be00000;
      118449: inst = 32'h8c50000;
      118450: inst = 32'h24612800;
      118451: inst = 32'h10a00000;
      118452: inst = 32'hca0001d;
      118453: inst = 32'h24822800;
      118454: inst = 32'h10a00000;
      118455: inst = 32'hca00004;
      118456: inst = 32'h38632800;
      118457: inst = 32'h38842800;
      118458: inst = 32'h10a00001;
      118459: inst = 32'hca0cebf;
      118460: inst = 32'h13e00001;
      118461: inst = 32'hfe0d96a;
      118462: inst = 32'h5be00000;
      118463: inst = 32'h8c50000;
      118464: inst = 32'h24612800;
      118465: inst = 32'h10a00000;
      118466: inst = 32'hca0001d;
      118467: inst = 32'h24822800;
      118468: inst = 32'h10a00000;
      118469: inst = 32'hca00004;
      118470: inst = 32'h38632800;
      118471: inst = 32'h38842800;
      118472: inst = 32'h10a00001;
      118473: inst = 32'hca0cecd;
      118474: inst = 32'h13e00001;
      118475: inst = 32'hfe0d96a;
      118476: inst = 32'h5be00000;
      118477: inst = 32'h8c50000;
      118478: inst = 32'h24612800;
      118479: inst = 32'h10a00000;
      118480: inst = 32'hca0001d;
      118481: inst = 32'h24822800;
      118482: inst = 32'h10a00000;
      118483: inst = 32'hca00004;
      118484: inst = 32'h38632800;
      118485: inst = 32'h38842800;
      118486: inst = 32'h10a00001;
      118487: inst = 32'hca0cedb;
      118488: inst = 32'h13e00001;
      118489: inst = 32'hfe0d96a;
      118490: inst = 32'h5be00000;
      118491: inst = 32'h8c50000;
      118492: inst = 32'h24612800;
      118493: inst = 32'h10a00000;
      118494: inst = 32'hca0001d;
      118495: inst = 32'h24822800;
      118496: inst = 32'h10a00000;
      118497: inst = 32'hca00004;
      118498: inst = 32'h38632800;
      118499: inst = 32'h38842800;
      118500: inst = 32'h10a00001;
      118501: inst = 32'hca0cee9;
      118502: inst = 32'h13e00001;
      118503: inst = 32'hfe0d96a;
      118504: inst = 32'h5be00000;
      118505: inst = 32'h8c50000;
      118506: inst = 32'h24612800;
      118507: inst = 32'h10a00000;
      118508: inst = 32'hca0001e;
      118509: inst = 32'h24822800;
      118510: inst = 32'h10a00000;
      118511: inst = 32'hca00004;
      118512: inst = 32'h38632800;
      118513: inst = 32'h38842800;
      118514: inst = 32'h10a00001;
      118515: inst = 32'hca0cef7;
      118516: inst = 32'h13e00001;
      118517: inst = 32'hfe0d96a;
      118518: inst = 32'h5be00000;
      118519: inst = 32'h8c50000;
      118520: inst = 32'h24612800;
      118521: inst = 32'h10a00000;
      118522: inst = 32'hca0001e;
      118523: inst = 32'h24822800;
      118524: inst = 32'h10a00000;
      118525: inst = 32'hca00004;
      118526: inst = 32'h38632800;
      118527: inst = 32'h38842800;
      118528: inst = 32'h10a00001;
      118529: inst = 32'hca0cf05;
      118530: inst = 32'h13e00001;
      118531: inst = 32'hfe0d96a;
      118532: inst = 32'h5be00000;
      118533: inst = 32'h8c50000;
      118534: inst = 32'h24612800;
      118535: inst = 32'h10a00000;
      118536: inst = 32'hca0001e;
      118537: inst = 32'h24822800;
      118538: inst = 32'h10a00000;
      118539: inst = 32'hca00004;
      118540: inst = 32'h38632800;
      118541: inst = 32'h38842800;
      118542: inst = 32'h10a00001;
      118543: inst = 32'hca0cf13;
      118544: inst = 32'h13e00001;
      118545: inst = 32'hfe0d96a;
      118546: inst = 32'h5be00000;
      118547: inst = 32'h8c50000;
      118548: inst = 32'h24612800;
      118549: inst = 32'h10a00000;
      118550: inst = 32'hca0001e;
      118551: inst = 32'h24822800;
      118552: inst = 32'h10a00000;
      118553: inst = 32'hca00004;
      118554: inst = 32'h38632800;
      118555: inst = 32'h38842800;
      118556: inst = 32'h10a00001;
      118557: inst = 32'hca0cf21;
      118558: inst = 32'h13e00001;
      118559: inst = 32'hfe0d96a;
      118560: inst = 32'h5be00000;
      118561: inst = 32'h8c50000;
      118562: inst = 32'h24612800;
      118563: inst = 32'h10a00000;
      118564: inst = 32'hca0001e;
      118565: inst = 32'h24822800;
      118566: inst = 32'h10a00000;
      118567: inst = 32'hca00004;
      118568: inst = 32'h38632800;
      118569: inst = 32'h38842800;
      118570: inst = 32'h10a00001;
      118571: inst = 32'hca0cf2f;
      118572: inst = 32'h13e00001;
      118573: inst = 32'hfe0d96a;
      118574: inst = 32'h5be00000;
      118575: inst = 32'h8c50000;
      118576: inst = 32'h24612800;
      118577: inst = 32'h10a00000;
      118578: inst = 32'hca0001e;
      118579: inst = 32'h24822800;
      118580: inst = 32'h10a00000;
      118581: inst = 32'hca00004;
      118582: inst = 32'h38632800;
      118583: inst = 32'h38842800;
      118584: inst = 32'h10a00001;
      118585: inst = 32'hca0cf3d;
      118586: inst = 32'h13e00001;
      118587: inst = 32'hfe0d96a;
      118588: inst = 32'h5be00000;
      118589: inst = 32'h8c50000;
      118590: inst = 32'h24612800;
      118591: inst = 32'h10a00000;
      118592: inst = 32'hca0001e;
      118593: inst = 32'h24822800;
      118594: inst = 32'h10a00000;
      118595: inst = 32'hca00004;
      118596: inst = 32'h38632800;
      118597: inst = 32'h38842800;
      118598: inst = 32'h10a00001;
      118599: inst = 32'hca0cf4b;
      118600: inst = 32'h13e00001;
      118601: inst = 32'hfe0d96a;
      118602: inst = 32'h5be00000;
      118603: inst = 32'h8c50000;
      118604: inst = 32'h24612800;
      118605: inst = 32'h10a00000;
      118606: inst = 32'hca0001e;
      118607: inst = 32'h24822800;
      118608: inst = 32'h10a00000;
      118609: inst = 32'hca00004;
      118610: inst = 32'h38632800;
      118611: inst = 32'h38842800;
      118612: inst = 32'h10a00001;
      118613: inst = 32'hca0cf59;
      118614: inst = 32'h13e00001;
      118615: inst = 32'hfe0d96a;
      118616: inst = 32'h5be00000;
      118617: inst = 32'h8c50000;
      118618: inst = 32'h24612800;
      118619: inst = 32'h10a00000;
      118620: inst = 32'hca0001e;
      118621: inst = 32'h24822800;
      118622: inst = 32'h10a00000;
      118623: inst = 32'hca00004;
      118624: inst = 32'h38632800;
      118625: inst = 32'h38842800;
      118626: inst = 32'h10a00001;
      118627: inst = 32'hca0cf67;
      118628: inst = 32'h13e00001;
      118629: inst = 32'hfe0d96a;
      118630: inst = 32'h5be00000;
      118631: inst = 32'h8c50000;
      118632: inst = 32'h24612800;
      118633: inst = 32'h10a00000;
      118634: inst = 32'hca0001e;
      118635: inst = 32'h24822800;
      118636: inst = 32'h10a00000;
      118637: inst = 32'hca00004;
      118638: inst = 32'h38632800;
      118639: inst = 32'h38842800;
      118640: inst = 32'h10a00001;
      118641: inst = 32'hca0cf75;
      118642: inst = 32'h13e00001;
      118643: inst = 32'hfe0d96a;
      118644: inst = 32'h5be00000;
      118645: inst = 32'h8c50000;
      118646: inst = 32'h24612800;
      118647: inst = 32'h10a00000;
      118648: inst = 32'hca0001e;
      118649: inst = 32'h24822800;
      118650: inst = 32'h10a00000;
      118651: inst = 32'hca00004;
      118652: inst = 32'h38632800;
      118653: inst = 32'h38842800;
      118654: inst = 32'h10a00001;
      118655: inst = 32'hca0cf83;
      118656: inst = 32'h13e00001;
      118657: inst = 32'hfe0d96a;
      118658: inst = 32'h5be00000;
      118659: inst = 32'h8c50000;
      118660: inst = 32'h24612800;
      118661: inst = 32'h10a00000;
      118662: inst = 32'hca0001e;
      118663: inst = 32'h24822800;
      118664: inst = 32'h10a00000;
      118665: inst = 32'hca00004;
      118666: inst = 32'h38632800;
      118667: inst = 32'h38842800;
      118668: inst = 32'h10a00001;
      118669: inst = 32'hca0cf91;
      118670: inst = 32'h13e00001;
      118671: inst = 32'hfe0d96a;
      118672: inst = 32'h5be00000;
      118673: inst = 32'h8c50000;
      118674: inst = 32'h24612800;
      118675: inst = 32'h10a00000;
      118676: inst = 32'hca0001e;
      118677: inst = 32'h24822800;
      118678: inst = 32'h10a00000;
      118679: inst = 32'hca00004;
      118680: inst = 32'h38632800;
      118681: inst = 32'h38842800;
      118682: inst = 32'h10a00001;
      118683: inst = 32'hca0cf9f;
      118684: inst = 32'h13e00001;
      118685: inst = 32'hfe0d96a;
      118686: inst = 32'h5be00000;
      118687: inst = 32'h8c50000;
      118688: inst = 32'h24612800;
      118689: inst = 32'h10a00000;
      118690: inst = 32'hca0001e;
      118691: inst = 32'h24822800;
      118692: inst = 32'h10a00000;
      118693: inst = 32'hca00004;
      118694: inst = 32'h38632800;
      118695: inst = 32'h38842800;
      118696: inst = 32'h10a00001;
      118697: inst = 32'hca0cfad;
      118698: inst = 32'h13e00001;
      118699: inst = 32'hfe0d96a;
      118700: inst = 32'h5be00000;
      118701: inst = 32'h8c50000;
      118702: inst = 32'h24612800;
      118703: inst = 32'h10a00000;
      118704: inst = 32'hca0001e;
      118705: inst = 32'h24822800;
      118706: inst = 32'h10a00000;
      118707: inst = 32'hca00004;
      118708: inst = 32'h38632800;
      118709: inst = 32'h38842800;
      118710: inst = 32'h10a00001;
      118711: inst = 32'hca0cfbb;
      118712: inst = 32'h13e00001;
      118713: inst = 32'hfe0d96a;
      118714: inst = 32'h5be00000;
      118715: inst = 32'h8c50000;
      118716: inst = 32'h24612800;
      118717: inst = 32'h10a00000;
      118718: inst = 32'hca0001e;
      118719: inst = 32'h24822800;
      118720: inst = 32'h10a00000;
      118721: inst = 32'hca00004;
      118722: inst = 32'h38632800;
      118723: inst = 32'h38842800;
      118724: inst = 32'h10a00001;
      118725: inst = 32'hca0cfc9;
      118726: inst = 32'h13e00001;
      118727: inst = 32'hfe0d96a;
      118728: inst = 32'h5be00000;
      118729: inst = 32'h8c50000;
      118730: inst = 32'h24612800;
      118731: inst = 32'h10a00000;
      118732: inst = 32'hca0001e;
      118733: inst = 32'h24822800;
      118734: inst = 32'h10a00000;
      118735: inst = 32'hca00004;
      118736: inst = 32'h38632800;
      118737: inst = 32'h38842800;
      118738: inst = 32'h10a00001;
      118739: inst = 32'hca0cfd7;
      118740: inst = 32'h13e00001;
      118741: inst = 32'hfe0d96a;
      118742: inst = 32'h5be00000;
      118743: inst = 32'h8c50000;
      118744: inst = 32'h24612800;
      118745: inst = 32'h10a00000;
      118746: inst = 32'hca0001e;
      118747: inst = 32'h24822800;
      118748: inst = 32'h10a00000;
      118749: inst = 32'hca00004;
      118750: inst = 32'h38632800;
      118751: inst = 32'h38842800;
      118752: inst = 32'h10a00001;
      118753: inst = 32'hca0cfe5;
      118754: inst = 32'h13e00001;
      118755: inst = 32'hfe0d96a;
      118756: inst = 32'h5be00000;
      118757: inst = 32'h8c50000;
      118758: inst = 32'h24612800;
      118759: inst = 32'h10a00000;
      118760: inst = 32'hca0001e;
      118761: inst = 32'h24822800;
      118762: inst = 32'h10a00000;
      118763: inst = 32'hca00004;
      118764: inst = 32'h38632800;
      118765: inst = 32'h38842800;
      118766: inst = 32'h10a00001;
      118767: inst = 32'hca0cff3;
      118768: inst = 32'h13e00001;
      118769: inst = 32'hfe0d96a;
      118770: inst = 32'h5be00000;
      118771: inst = 32'h8c50000;
      118772: inst = 32'h24612800;
      118773: inst = 32'h10a00000;
      118774: inst = 32'hca0001e;
      118775: inst = 32'h24822800;
      118776: inst = 32'h10a00000;
      118777: inst = 32'hca00004;
      118778: inst = 32'h38632800;
      118779: inst = 32'h38842800;
      118780: inst = 32'h10a00001;
      118781: inst = 32'hca0d001;
      118782: inst = 32'h13e00001;
      118783: inst = 32'hfe0d96a;
      118784: inst = 32'h5be00000;
      118785: inst = 32'h8c50000;
      118786: inst = 32'h24612800;
      118787: inst = 32'h10a00000;
      118788: inst = 32'hca0001e;
      118789: inst = 32'h24822800;
      118790: inst = 32'h10a00000;
      118791: inst = 32'hca00004;
      118792: inst = 32'h38632800;
      118793: inst = 32'h38842800;
      118794: inst = 32'h10a00001;
      118795: inst = 32'hca0d00f;
      118796: inst = 32'h13e00001;
      118797: inst = 32'hfe0d96a;
      118798: inst = 32'h5be00000;
      118799: inst = 32'h8c50000;
      118800: inst = 32'h24612800;
      118801: inst = 32'h10a00000;
      118802: inst = 32'hca0001e;
      118803: inst = 32'h24822800;
      118804: inst = 32'h10a00000;
      118805: inst = 32'hca00004;
      118806: inst = 32'h38632800;
      118807: inst = 32'h38842800;
      118808: inst = 32'h10a00001;
      118809: inst = 32'hca0d01d;
      118810: inst = 32'h13e00001;
      118811: inst = 32'hfe0d96a;
      118812: inst = 32'h5be00000;
      118813: inst = 32'h8c50000;
      118814: inst = 32'h24612800;
      118815: inst = 32'h10a00000;
      118816: inst = 32'hca0001e;
      118817: inst = 32'h24822800;
      118818: inst = 32'h10a00000;
      118819: inst = 32'hca00004;
      118820: inst = 32'h38632800;
      118821: inst = 32'h38842800;
      118822: inst = 32'h10a00001;
      118823: inst = 32'hca0d02b;
      118824: inst = 32'h13e00001;
      118825: inst = 32'hfe0d96a;
      118826: inst = 32'h5be00000;
      118827: inst = 32'h8c50000;
      118828: inst = 32'h24612800;
      118829: inst = 32'h10a00000;
      118830: inst = 32'hca0001e;
      118831: inst = 32'h24822800;
      118832: inst = 32'h10a00000;
      118833: inst = 32'hca00004;
      118834: inst = 32'h38632800;
      118835: inst = 32'h38842800;
      118836: inst = 32'h10a00001;
      118837: inst = 32'hca0d039;
      118838: inst = 32'h13e00001;
      118839: inst = 32'hfe0d96a;
      118840: inst = 32'h5be00000;
      118841: inst = 32'h8c50000;
      118842: inst = 32'h24612800;
      118843: inst = 32'h10a00000;
      118844: inst = 32'hca0001e;
      118845: inst = 32'h24822800;
      118846: inst = 32'h10a00000;
      118847: inst = 32'hca00004;
      118848: inst = 32'h38632800;
      118849: inst = 32'h38842800;
      118850: inst = 32'h10a00001;
      118851: inst = 32'hca0d047;
      118852: inst = 32'h13e00001;
      118853: inst = 32'hfe0d96a;
      118854: inst = 32'h5be00000;
      118855: inst = 32'h8c50000;
      118856: inst = 32'h24612800;
      118857: inst = 32'h10a00000;
      118858: inst = 32'hca0001e;
      118859: inst = 32'h24822800;
      118860: inst = 32'h10a00000;
      118861: inst = 32'hca00004;
      118862: inst = 32'h38632800;
      118863: inst = 32'h38842800;
      118864: inst = 32'h10a00001;
      118865: inst = 32'hca0d055;
      118866: inst = 32'h13e00001;
      118867: inst = 32'hfe0d96a;
      118868: inst = 32'h5be00000;
      118869: inst = 32'h8c50000;
      118870: inst = 32'h24612800;
      118871: inst = 32'h10a00000;
      118872: inst = 32'hca0001e;
      118873: inst = 32'h24822800;
      118874: inst = 32'h10a00000;
      118875: inst = 32'hca00004;
      118876: inst = 32'h38632800;
      118877: inst = 32'h38842800;
      118878: inst = 32'h10a00001;
      118879: inst = 32'hca0d063;
      118880: inst = 32'h13e00001;
      118881: inst = 32'hfe0d96a;
      118882: inst = 32'h5be00000;
      118883: inst = 32'h8c50000;
      118884: inst = 32'h24612800;
      118885: inst = 32'h10a00000;
      118886: inst = 32'hca0001e;
      118887: inst = 32'h24822800;
      118888: inst = 32'h10a00000;
      118889: inst = 32'hca00004;
      118890: inst = 32'h38632800;
      118891: inst = 32'h38842800;
      118892: inst = 32'h10a00001;
      118893: inst = 32'hca0d071;
      118894: inst = 32'h13e00001;
      118895: inst = 32'hfe0d96a;
      118896: inst = 32'h5be00000;
      118897: inst = 32'h8c50000;
      118898: inst = 32'h24612800;
      118899: inst = 32'h10a00000;
      118900: inst = 32'hca0001e;
      118901: inst = 32'h24822800;
      118902: inst = 32'h10a00000;
      118903: inst = 32'hca00004;
      118904: inst = 32'h38632800;
      118905: inst = 32'h38842800;
      118906: inst = 32'h10a00001;
      118907: inst = 32'hca0d07f;
      118908: inst = 32'h13e00001;
      118909: inst = 32'hfe0d96a;
      118910: inst = 32'h5be00000;
      118911: inst = 32'h8c50000;
      118912: inst = 32'h24612800;
      118913: inst = 32'h10a00000;
      118914: inst = 32'hca0001e;
      118915: inst = 32'h24822800;
      118916: inst = 32'h10a00000;
      118917: inst = 32'hca00004;
      118918: inst = 32'h38632800;
      118919: inst = 32'h38842800;
      118920: inst = 32'h10a00001;
      118921: inst = 32'hca0d08d;
      118922: inst = 32'h13e00001;
      118923: inst = 32'hfe0d96a;
      118924: inst = 32'h5be00000;
      118925: inst = 32'h8c50000;
      118926: inst = 32'h24612800;
      118927: inst = 32'h10a00000;
      118928: inst = 32'hca0001e;
      118929: inst = 32'h24822800;
      118930: inst = 32'h10a00000;
      118931: inst = 32'hca00004;
      118932: inst = 32'h38632800;
      118933: inst = 32'h38842800;
      118934: inst = 32'h10a00001;
      118935: inst = 32'hca0d09b;
      118936: inst = 32'h13e00001;
      118937: inst = 32'hfe0d96a;
      118938: inst = 32'h5be00000;
      118939: inst = 32'h8c50000;
      118940: inst = 32'h24612800;
      118941: inst = 32'h10a00000;
      118942: inst = 32'hca0001e;
      118943: inst = 32'h24822800;
      118944: inst = 32'h10a00000;
      118945: inst = 32'hca00004;
      118946: inst = 32'h38632800;
      118947: inst = 32'h38842800;
      118948: inst = 32'h10a00001;
      118949: inst = 32'hca0d0a9;
      118950: inst = 32'h13e00001;
      118951: inst = 32'hfe0d96a;
      118952: inst = 32'h5be00000;
      118953: inst = 32'h8c50000;
      118954: inst = 32'h24612800;
      118955: inst = 32'h10a00000;
      118956: inst = 32'hca0001e;
      118957: inst = 32'h24822800;
      118958: inst = 32'h10a00000;
      118959: inst = 32'hca00004;
      118960: inst = 32'h38632800;
      118961: inst = 32'h38842800;
      118962: inst = 32'h10a00001;
      118963: inst = 32'hca0d0b7;
      118964: inst = 32'h13e00001;
      118965: inst = 32'hfe0d96a;
      118966: inst = 32'h5be00000;
      118967: inst = 32'h8c50000;
      118968: inst = 32'h24612800;
      118969: inst = 32'h10a00000;
      118970: inst = 32'hca0001e;
      118971: inst = 32'h24822800;
      118972: inst = 32'h10a00000;
      118973: inst = 32'hca00004;
      118974: inst = 32'h38632800;
      118975: inst = 32'h38842800;
      118976: inst = 32'h10a00001;
      118977: inst = 32'hca0d0c5;
      118978: inst = 32'h13e00001;
      118979: inst = 32'hfe0d96a;
      118980: inst = 32'h5be00000;
      118981: inst = 32'h8c50000;
      118982: inst = 32'h24612800;
      118983: inst = 32'h10a00000;
      118984: inst = 32'hca0001e;
      118985: inst = 32'h24822800;
      118986: inst = 32'h10a00000;
      118987: inst = 32'hca00004;
      118988: inst = 32'h38632800;
      118989: inst = 32'h38842800;
      118990: inst = 32'h10a00001;
      118991: inst = 32'hca0d0d3;
      118992: inst = 32'h13e00001;
      118993: inst = 32'hfe0d96a;
      118994: inst = 32'h5be00000;
      118995: inst = 32'h8c50000;
      118996: inst = 32'h24612800;
      118997: inst = 32'h10a00000;
      118998: inst = 32'hca0001e;
      118999: inst = 32'h24822800;
      119000: inst = 32'h10a00000;
      119001: inst = 32'hca00004;
      119002: inst = 32'h38632800;
      119003: inst = 32'h38842800;
      119004: inst = 32'h10a00001;
      119005: inst = 32'hca0d0e1;
      119006: inst = 32'h13e00001;
      119007: inst = 32'hfe0d96a;
      119008: inst = 32'h5be00000;
      119009: inst = 32'h8c50000;
      119010: inst = 32'h24612800;
      119011: inst = 32'h10a00000;
      119012: inst = 32'hca0001e;
      119013: inst = 32'h24822800;
      119014: inst = 32'h10a00000;
      119015: inst = 32'hca00004;
      119016: inst = 32'h38632800;
      119017: inst = 32'h38842800;
      119018: inst = 32'h10a00001;
      119019: inst = 32'hca0d0ef;
      119020: inst = 32'h13e00001;
      119021: inst = 32'hfe0d96a;
      119022: inst = 32'h5be00000;
      119023: inst = 32'h8c50000;
      119024: inst = 32'h24612800;
      119025: inst = 32'h10a00000;
      119026: inst = 32'hca0001e;
      119027: inst = 32'h24822800;
      119028: inst = 32'h10a00000;
      119029: inst = 32'hca00004;
      119030: inst = 32'h38632800;
      119031: inst = 32'h38842800;
      119032: inst = 32'h10a00001;
      119033: inst = 32'hca0d0fd;
      119034: inst = 32'h13e00001;
      119035: inst = 32'hfe0d96a;
      119036: inst = 32'h5be00000;
      119037: inst = 32'h8c50000;
      119038: inst = 32'h24612800;
      119039: inst = 32'h10a00000;
      119040: inst = 32'hca0001e;
      119041: inst = 32'h24822800;
      119042: inst = 32'h10a00000;
      119043: inst = 32'hca00004;
      119044: inst = 32'h38632800;
      119045: inst = 32'h38842800;
      119046: inst = 32'h10a00001;
      119047: inst = 32'hca0d10b;
      119048: inst = 32'h13e00001;
      119049: inst = 32'hfe0d96a;
      119050: inst = 32'h5be00000;
      119051: inst = 32'h8c50000;
      119052: inst = 32'h24612800;
      119053: inst = 32'h10a00000;
      119054: inst = 32'hca0001e;
      119055: inst = 32'h24822800;
      119056: inst = 32'h10a00000;
      119057: inst = 32'hca00004;
      119058: inst = 32'h38632800;
      119059: inst = 32'h38842800;
      119060: inst = 32'h10a00001;
      119061: inst = 32'hca0d119;
      119062: inst = 32'h13e00001;
      119063: inst = 32'hfe0d96a;
      119064: inst = 32'h5be00000;
      119065: inst = 32'h8c50000;
      119066: inst = 32'h24612800;
      119067: inst = 32'h10a00000;
      119068: inst = 32'hca0001e;
      119069: inst = 32'h24822800;
      119070: inst = 32'h10a00000;
      119071: inst = 32'hca00004;
      119072: inst = 32'h38632800;
      119073: inst = 32'h38842800;
      119074: inst = 32'h10a00001;
      119075: inst = 32'hca0d127;
      119076: inst = 32'h13e00001;
      119077: inst = 32'hfe0d96a;
      119078: inst = 32'h5be00000;
      119079: inst = 32'h8c50000;
      119080: inst = 32'h24612800;
      119081: inst = 32'h10a00000;
      119082: inst = 32'hca0001e;
      119083: inst = 32'h24822800;
      119084: inst = 32'h10a00000;
      119085: inst = 32'hca00004;
      119086: inst = 32'h38632800;
      119087: inst = 32'h38842800;
      119088: inst = 32'h10a00001;
      119089: inst = 32'hca0d135;
      119090: inst = 32'h13e00001;
      119091: inst = 32'hfe0d96a;
      119092: inst = 32'h5be00000;
      119093: inst = 32'h8c50000;
      119094: inst = 32'h24612800;
      119095: inst = 32'h10a00000;
      119096: inst = 32'hca0001e;
      119097: inst = 32'h24822800;
      119098: inst = 32'h10a00000;
      119099: inst = 32'hca00004;
      119100: inst = 32'h38632800;
      119101: inst = 32'h38842800;
      119102: inst = 32'h10a00001;
      119103: inst = 32'hca0d143;
      119104: inst = 32'h13e00001;
      119105: inst = 32'hfe0d96a;
      119106: inst = 32'h5be00000;
      119107: inst = 32'h8c50000;
      119108: inst = 32'h24612800;
      119109: inst = 32'h10a00000;
      119110: inst = 32'hca0001e;
      119111: inst = 32'h24822800;
      119112: inst = 32'h10a00000;
      119113: inst = 32'hca00004;
      119114: inst = 32'h38632800;
      119115: inst = 32'h38842800;
      119116: inst = 32'h10a00001;
      119117: inst = 32'hca0d151;
      119118: inst = 32'h13e00001;
      119119: inst = 32'hfe0d96a;
      119120: inst = 32'h5be00000;
      119121: inst = 32'h8c50000;
      119122: inst = 32'h24612800;
      119123: inst = 32'h10a00000;
      119124: inst = 32'hca0001e;
      119125: inst = 32'h24822800;
      119126: inst = 32'h10a00000;
      119127: inst = 32'hca00004;
      119128: inst = 32'h38632800;
      119129: inst = 32'h38842800;
      119130: inst = 32'h10a00001;
      119131: inst = 32'hca0d15f;
      119132: inst = 32'h13e00001;
      119133: inst = 32'hfe0d96a;
      119134: inst = 32'h5be00000;
      119135: inst = 32'h8c50000;
      119136: inst = 32'h24612800;
      119137: inst = 32'h10a00000;
      119138: inst = 32'hca0001e;
      119139: inst = 32'h24822800;
      119140: inst = 32'h10a00000;
      119141: inst = 32'hca00004;
      119142: inst = 32'h38632800;
      119143: inst = 32'h38842800;
      119144: inst = 32'h10a00001;
      119145: inst = 32'hca0d16d;
      119146: inst = 32'h13e00001;
      119147: inst = 32'hfe0d96a;
      119148: inst = 32'h5be00000;
      119149: inst = 32'h8c50000;
      119150: inst = 32'h24612800;
      119151: inst = 32'h10a00000;
      119152: inst = 32'hca0001e;
      119153: inst = 32'h24822800;
      119154: inst = 32'h10a00000;
      119155: inst = 32'hca00004;
      119156: inst = 32'h38632800;
      119157: inst = 32'h38842800;
      119158: inst = 32'h10a00001;
      119159: inst = 32'hca0d17b;
      119160: inst = 32'h13e00001;
      119161: inst = 32'hfe0d96a;
      119162: inst = 32'h5be00000;
      119163: inst = 32'h8c50000;
      119164: inst = 32'h24612800;
      119165: inst = 32'h10a00000;
      119166: inst = 32'hca0001e;
      119167: inst = 32'h24822800;
      119168: inst = 32'h10a00000;
      119169: inst = 32'hca00004;
      119170: inst = 32'h38632800;
      119171: inst = 32'h38842800;
      119172: inst = 32'h10a00001;
      119173: inst = 32'hca0d189;
      119174: inst = 32'h13e00001;
      119175: inst = 32'hfe0d96a;
      119176: inst = 32'h5be00000;
      119177: inst = 32'h8c50000;
      119178: inst = 32'h24612800;
      119179: inst = 32'h10a00000;
      119180: inst = 32'hca0001e;
      119181: inst = 32'h24822800;
      119182: inst = 32'h10a00000;
      119183: inst = 32'hca00004;
      119184: inst = 32'h38632800;
      119185: inst = 32'h38842800;
      119186: inst = 32'h10a00001;
      119187: inst = 32'hca0d197;
      119188: inst = 32'h13e00001;
      119189: inst = 32'hfe0d96a;
      119190: inst = 32'h5be00000;
      119191: inst = 32'h8c50000;
      119192: inst = 32'h24612800;
      119193: inst = 32'h10a00000;
      119194: inst = 32'hca0001e;
      119195: inst = 32'h24822800;
      119196: inst = 32'h10a00000;
      119197: inst = 32'hca00004;
      119198: inst = 32'h38632800;
      119199: inst = 32'h38842800;
      119200: inst = 32'h10a00001;
      119201: inst = 32'hca0d1a5;
      119202: inst = 32'h13e00001;
      119203: inst = 32'hfe0d96a;
      119204: inst = 32'h5be00000;
      119205: inst = 32'h8c50000;
      119206: inst = 32'h24612800;
      119207: inst = 32'h10a00000;
      119208: inst = 32'hca0001e;
      119209: inst = 32'h24822800;
      119210: inst = 32'h10a00000;
      119211: inst = 32'hca00004;
      119212: inst = 32'h38632800;
      119213: inst = 32'h38842800;
      119214: inst = 32'h10a00001;
      119215: inst = 32'hca0d1b3;
      119216: inst = 32'h13e00001;
      119217: inst = 32'hfe0d96a;
      119218: inst = 32'h5be00000;
      119219: inst = 32'h8c50000;
      119220: inst = 32'h24612800;
      119221: inst = 32'h10a00000;
      119222: inst = 32'hca0001e;
      119223: inst = 32'h24822800;
      119224: inst = 32'h10a00000;
      119225: inst = 32'hca00004;
      119226: inst = 32'h38632800;
      119227: inst = 32'h38842800;
      119228: inst = 32'h10a00001;
      119229: inst = 32'hca0d1c1;
      119230: inst = 32'h13e00001;
      119231: inst = 32'hfe0d96a;
      119232: inst = 32'h5be00000;
      119233: inst = 32'h8c50000;
      119234: inst = 32'h24612800;
      119235: inst = 32'h10a00000;
      119236: inst = 32'hca0001e;
      119237: inst = 32'h24822800;
      119238: inst = 32'h10a00000;
      119239: inst = 32'hca00004;
      119240: inst = 32'h38632800;
      119241: inst = 32'h38842800;
      119242: inst = 32'h10a00001;
      119243: inst = 32'hca0d1cf;
      119244: inst = 32'h13e00001;
      119245: inst = 32'hfe0d96a;
      119246: inst = 32'h5be00000;
      119247: inst = 32'h8c50000;
      119248: inst = 32'h24612800;
      119249: inst = 32'h10a00000;
      119250: inst = 32'hca0001e;
      119251: inst = 32'h24822800;
      119252: inst = 32'h10a00000;
      119253: inst = 32'hca00004;
      119254: inst = 32'h38632800;
      119255: inst = 32'h38842800;
      119256: inst = 32'h10a00001;
      119257: inst = 32'hca0d1dd;
      119258: inst = 32'h13e00001;
      119259: inst = 32'hfe0d96a;
      119260: inst = 32'h5be00000;
      119261: inst = 32'h8c50000;
      119262: inst = 32'h24612800;
      119263: inst = 32'h10a00000;
      119264: inst = 32'hca0001e;
      119265: inst = 32'h24822800;
      119266: inst = 32'h10a00000;
      119267: inst = 32'hca00004;
      119268: inst = 32'h38632800;
      119269: inst = 32'h38842800;
      119270: inst = 32'h10a00001;
      119271: inst = 32'hca0d1eb;
      119272: inst = 32'h13e00001;
      119273: inst = 32'hfe0d96a;
      119274: inst = 32'h5be00000;
      119275: inst = 32'h8c50000;
      119276: inst = 32'h24612800;
      119277: inst = 32'h10a00000;
      119278: inst = 32'hca0001e;
      119279: inst = 32'h24822800;
      119280: inst = 32'h10a00000;
      119281: inst = 32'hca00004;
      119282: inst = 32'h38632800;
      119283: inst = 32'h38842800;
      119284: inst = 32'h10a00001;
      119285: inst = 32'hca0d1f9;
      119286: inst = 32'h13e00001;
      119287: inst = 32'hfe0d96a;
      119288: inst = 32'h5be00000;
      119289: inst = 32'h8c50000;
      119290: inst = 32'h24612800;
      119291: inst = 32'h10a00000;
      119292: inst = 32'hca0001e;
      119293: inst = 32'h24822800;
      119294: inst = 32'h10a00000;
      119295: inst = 32'hca00004;
      119296: inst = 32'h38632800;
      119297: inst = 32'h38842800;
      119298: inst = 32'h10a00001;
      119299: inst = 32'hca0d207;
      119300: inst = 32'h13e00001;
      119301: inst = 32'hfe0d96a;
      119302: inst = 32'h5be00000;
      119303: inst = 32'h8c50000;
      119304: inst = 32'h24612800;
      119305: inst = 32'h10a00000;
      119306: inst = 32'hca0001e;
      119307: inst = 32'h24822800;
      119308: inst = 32'h10a00000;
      119309: inst = 32'hca00004;
      119310: inst = 32'h38632800;
      119311: inst = 32'h38842800;
      119312: inst = 32'h10a00001;
      119313: inst = 32'hca0d215;
      119314: inst = 32'h13e00001;
      119315: inst = 32'hfe0d96a;
      119316: inst = 32'h5be00000;
      119317: inst = 32'h8c50000;
      119318: inst = 32'h24612800;
      119319: inst = 32'h10a00000;
      119320: inst = 32'hca0001e;
      119321: inst = 32'h24822800;
      119322: inst = 32'h10a00000;
      119323: inst = 32'hca00004;
      119324: inst = 32'h38632800;
      119325: inst = 32'h38842800;
      119326: inst = 32'h10a00001;
      119327: inst = 32'hca0d223;
      119328: inst = 32'h13e00001;
      119329: inst = 32'hfe0d96a;
      119330: inst = 32'h5be00000;
      119331: inst = 32'h8c50000;
      119332: inst = 32'h24612800;
      119333: inst = 32'h10a00000;
      119334: inst = 32'hca0001e;
      119335: inst = 32'h24822800;
      119336: inst = 32'h10a00000;
      119337: inst = 32'hca00004;
      119338: inst = 32'h38632800;
      119339: inst = 32'h38842800;
      119340: inst = 32'h10a00001;
      119341: inst = 32'hca0d231;
      119342: inst = 32'h13e00001;
      119343: inst = 32'hfe0d96a;
      119344: inst = 32'h5be00000;
      119345: inst = 32'h8c50000;
      119346: inst = 32'h24612800;
      119347: inst = 32'h10a00000;
      119348: inst = 32'hca0001e;
      119349: inst = 32'h24822800;
      119350: inst = 32'h10a00000;
      119351: inst = 32'hca00004;
      119352: inst = 32'h38632800;
      119353: inst = 32'h38842800;
      119354: inst = 32'h10a00001;
      119355: inst = 32'hca0d23f;
      119356: inst = 32'h13e00001;
      119357: inst = 32'hfe0d96a;
      119358: inst = 32'h5be00000;
      119359: inst = 32'h8c50000;
      119360: inst = 32'h24612800;
      119361: inst = 32'h10a00000;
      119362: inst = 32'hca0001e;
      119363: inst = 32'h24822800;
      119364: inst = 32'h10a00000;
      119365: inst = 32'hca00004;
      119366: inst = 32'h38632800;
      119367: inst = 32'h38842800;
      119368: inst = 32'h10a00001;
      119369: inst = 32'hca0d24d;
      119370: inst = 32'h13e00001;
      119371: inst = 32'hfe0d96a;
      119372: inst = 32'h5be00000;
      119373: inst = 32'h8c50000;
      119374: inst = 32'h24612800;
      119375: inst = 32'h10a00000;
      119376: inst = 32'hca0001e;
      119377: inst = 32'h24822800;
      119378: inst = 32'h10a00000;
      119379: inst = 32'hca00004;
      119380: inst = 32'h38632800;
      119381: inst = 32'h38842800;
      119382: inst = 32'h10a00001;
      119383: inst = 32'hca0d25b;
      119384: inst = 32'h13e00001;
      119385: inst = 32'hfe0d96a;
      119386: inst = 32'h5be00000;
      119387: inst = 32'h8c50000;
      119388: inst = 32'h24612800;
      119389: inst = 32'h10a00000;
      119390: inst = 32'hca0001e;
      119391: inst = 32'h24822800;
      119392: inst = 32'h10a00000;
      119393: inst = 32'hca00004;
      119394: inst = 32'h38632800;
      119395: inst = 32'h38842800;
      119396: inst = 32'h10a00001;
      119397: inst = 32'hca0d269;
      119398: inst = 32'h13e00001;
      119399: inst = 32'hfe0d96a;
      119400: inst = 32'h5be00000;
      119401: inst = 32'h8c50000;
      119402: inst = 32'h24612800;
      119403: inst = 32'h10a00000;
      119404: inst = 32'hca0001e;
      119405: inst = 32'h24822800;
      119406: inst = 32'h10a00000;
      119407: inst = 32'hca00004;
      119408: inst = 32'h38632800;
      119409: inst = 32'h38842800;
      119410: inst = 32'h10a00001;
      119411: inst = 32'hca0d277;
      119412: inst = 32'h13e00001;
      119413: inst = 32'hfe0d96a;
      119414: inst = 32'h5be00000;
      119415: inst = 32'h8c50000;
      119416: inst = 32'h24612800;
      119417: inst = 32'h10a00000;
      119418: inst = 32'hca0001e;
      119419: inst = 32'h24822800;
      119420: inst = 32'h10a00000;
      119421: inst = 32'hca00004;
      119422: inst = 32'h38632800;
      119423: inst = 32'h38842800;
      119424: inst = 32'h10a00001;
      119425: inst = 32'hca0d285;
      119426: inst = 32'h13e00001;
      119427: inst = 32'hfe0d96a;
      119428: inst = 32'h5be00000;
      119429: inst = 32'h8c50000;
      119430: inst = 32'h24612800;
      119431: inst = 32'h10a00000;
      119432: inst = 32'hca0001e;
      119433: inst = 32'h24822800;
      119434: inst = 32'h10a00000;
      119435: inst = 32'hca00004;
      119436: inst = 32'h38632800;
      119437: inst = 32'h38842800;
      119438: inst = 32'h10a00001;
      119439: inst = 32'hca0d293;
      119440: inst = 32'h13e00001;
      119441: inst = 32'hfe0d96a;
      119442: inst = 32'h5be00000;
      119443: inst = 32'h8c50000;
      119444: inst = 32'h24612800;
      119445: inst = 32'h10a00000;
      119446: inst = 32'hca0001e;
      119447: inst = 32'h24822800;
      119448: inst = 32'h10a00000;
      119449: inst = 32'hca00004;
      119450: inst = 32'h38632800;
      119451: inst = 32'h38842800;
      119452: inst = 32'h10a00001;
      119453: inst = 32'hca0d2a1;
      119454: inst = 32'h13e00001;
      119455: inst = 32'hfe0d96a;
      119456: inst = 32'h5be00000;
      119457: inst = 32'h8c50000;
      119458: inst = 32'h24612800;
      119459: inst = 32'h10a00000;
      119460: inst = 32'hca0001e;
      119461: inst = 32'h24822800;
      119462: inst = 32'h10a00000;
      119463: inst = 32'hca00004;
      119464: inst = 32'h38632800;
      119465: inst = 32'h38842800;
      119466: inst = 32'h10a00001;
      119467: inst = 32'hca0d2af;
      119468: inst = 32'h13e00001;
      119469: inst = 32'hfe0d96a;
      119470: inst = 32'h5be00000;
      119471: inst = 32'h8c50000;
      119472: inst = 32'h24612800;
      119473: inst = 32'h10a00000;
      119474: inst = 32'hca0001e;
      119475: inst = 32'h24822800;
      119476: inst = 32'h10a00000;
      119477: inst = 32'hca00004;
      119478: inst = 32'h38632800;
      119479: inst = 32'h38842800;
      119480: inst = 32'h10a00001;
      119481: inst = 32'hca0d2bd;
      119482: inst = 32'h13e00001;
      119483: inst = 32'hfe0d96a;
      119484: inst = 32'h5be00000;
      119485: inst = 32'h8c50000;
      119486: inst = 32'h24612800;
      119487: inst = 32'h10a00000;
      119488: inst = 32'hca0001e;
      119489: inst = 32'h24822800;
      119490: inst = 32'h10a00000;
      119491: inst = 32'hca00004;
      119492: inst = 32'h38632800;
      119493: inst = 32'h38842800;
      119494: inst = 32'h10a00001;
      119495: inst = 32'hca0d2cb;
      119496: inst = 32'h13e00001;
      119497: inst = 32'hfe0d96a;
      119498: inst = 32'h5be00000;
      119499: inst = 32'h8c50000;
      119500: inst = 32'h24612800;
      119501: inst = 32'h10a00000;
      119502: inst = 32'hca0001e;
      119503: inst = 32'h24822800;
      119504: inst = 32'h10a00000;
      119505: inst = 32'hca00004;
      119506: inst = 32'h38632800;
      119507: inst = 32'h38842800;
      119508: inst = 32'h10a00001;
      119509: inst = 32'hca0d2d9;
      119510: inst = 32'h13e00001;
      119511: inst = 32'hfe0d96a;
      119512: inst = 32'h5be00000;
      119513: inst = 32'h8c50000;
      119514: inst = 32'h24612800;
      119515: inst = 32'h10a00000;
      119516: inst = 32'hca0001e;
      119517: inst = 32'h24822800;
      119518: inst = 32'h10a00000;
      119519: inst = 32'hca00004;
      119520: inst = 32'h38632800;
      119521: inst = 32'h38842800;
      119522: inst = 32'h10a00001;
      119523: inst = 32'hca0d2e7;
      119524: inst = 32'h13e00001;
      119525: inst = 32'hfe0d96a;
      119526: inst = 32'h5be00000;
      119527: inst = 32'h8c50000;
      119528: inst = 32'h24612800;
      119529: inst = 32'h10a00000;
      119530: inst = 32'hca0001e;
      119531: inst = 32'h24822800;
      119532: inst = 32'h10a00000;
      119533: inst = 32'hca00004;
      119534: inst = 32'h38632800;
      119535: inst = 32'h38842800;
      119536: inst = 32'h10a00001;
      119537: inst = 32'hca0d2f5;
      119538: inst = 32'h13e00001;
      119539: inst = 32'hfe0d96a;
      119540: inst = 32'h5be00000;
      119541: inst = 32'h8c50000;
      119542: inst = 32'h24612800;
      119543: inst = 32'h10a00000;
      119544: inst = 32'hca0001e;
      119545: inst = 32'h24822800;
      119546: inst = 32'h10a00000;
      119547: inst = 32'hca00004;
      119548: inst = 32'h38632800;
      119549: inst = 32'h38842800;
      119550: inst = 32'h10a00001;
      119551: inst = 32'hca0d303;
      119552: inst = 32'h13e00001;
      119553: inst = 32'hfe0d96a;
      119554: inst = 32'h5be00000;
      119555: inst = 32'h8c50000;
      119556: inst = 32'h24612800;
      119557: inst = 32'h10a00000;
      119558: inst = 32'hca0001e;
      119559: inst = 32'h24822800;
      119560: inst = 32'h10a00000;
      119561: inst = 32'hca00004;
      119562: inst = 32'h38632800;
      119563: inst = 32'h38842800;
      119564: inst = 32'h10a00001;
      119565: inst = 32'hca0d311;
      119566: inst = 32'h13e00001;
      119567: inst = 32'hfe0d96a;
      119568: inst = 32'h5be00000;
      119569: inst = 32'h8c50000;
      119570: inst = 32'h24612800;
      119571: inst = 32'h10a00000;
      119572: inst = 32'hca0001e;
      119573: inst = 32'h24822800;
      119574: inst = 32'h10a00000;
      119575: inst = 32'hca00004;
      119576: inst = 32'h38632800;
      119577: inst = 32'h38842800;
      119578: inst = 32'h10a00001;
      119579: inst = 32'hca0d31f;
      119580: inst = 32'h13e00001;
      119581: inst = 32'hfe0d96a;
      119582: inst = 32'h5be00000;
      119583: inst = 32'h8c50000;
      119584: inst = 32'h24612800;
      119585: inst = 32'h10a00000;
      119586: inst = 32'hca0001e;
      119587: inst = 32'h24822800;
      119588: inst = 32'h10a00000;
      119589: inst = 32'hca00004;
      119590: inst = 32'h38632800;
      119591: inst = 32'h38842800;
      119592: inst = 32'h10a00001;
      119593: inst = 32'hca0d32d;
      119594: inst = 32'h13e00001;
      119595: inst = 32'hfe0d96a;
      119596: inst = 32'h5be00000;
      119597: inst = 32'h8c50000;
      119598: inst = 32'h24612800;
      119599: inst = 32'h10a00000;
      119600: inst = 32'hca0001e;
      119601: inst = 32'h24822800;
      119602: inst = 32'h10a00000;
      119603: inst = 32'hca00004;
      119604: inst = 32'h38632800;
      119605: inst = 32'h38842800;
      119606: inst = 32'h10a00001;
      119607: inst = 32'hca0d33b;
      119608: inst = 32'h13e00001;
      119609: inst = 32'hfe0d96a;
      119610: inst = 32'h5be00000;
      119611: inst = 32'h8c50000;
      119612: inst = 32'h24612800;
      119613: inst = 32'h10a00000;
      119614: inst = 32'hca0001e;
      119615: inst = 32'h24822800;
      119616: inst = 32'h10a00000;
      119617: inst = 32'hca00004;
      119618: inst = 32'h38632800;
      119619: inst = 32'h38842800;
      119620: inst = 32'h10a00001;
      119621: inst = 32'hca0d349;
      119622: inst = 32'h13e00001;
      119623: inst = 32'hfe0d96a;
      119624: inst = 32'h5be00000;
      119625: inst = 32'h8c50000;
      119626: inst = 32'h24612800;
      119627: inst = 32'h10a00000;
      119628: inst = 32'hca0001e;
      119629: inst = 32'h24822800;
      119630: inst = 32'h10a00000;
      119631: inst = 32'hca00004;
      119632: inst = 32'h38632800;
      119633: inst = 32'h38842800;
      119634: inst = 32'h10a00001;
      119635: inst = 32'hca0d357;
      119636: inst = 32'h13e00001;
      119637: inst = 32'hfe0d96a;
      119638: inst = 32'h5be00000;
      119639: inst = 32'h8c50000;
      119640: inst = 32'h24612800;
      119641: inst = 32'h10a00000;
      119642: inst = 32'hca0001e;
      119643: inst = 32'h24822800;
      119644: inst = 32'h10a00000;
      119645: inst = 32'hca00004;
      119646: inst = 32'h38632800;
      119647: inst = 32'h38842800;
      119648: inst = 32'h10a00001;
      119649: inst = 32'hca0d365;
      119650: inst = 32'h13e00001;
      119651: inst = 32'hfe0d96a;
      119652: inst = 32'h5be00000;
      119653: inst = 32'h8c50000;
      119654: inst = 32'h24612800;
      119655: inst = 32'h10a00000;
      119656: inst = 32'hca0001e;
      119657: inst = 32'h24822800;
      119658: inst = 32'h10a00000;
      119659: inst = 32'hca00004;
      119660: inst = 32'h38632800;
      119661: inst = 32'h38842800;
      119662: inst = 32'h10a00001;
      119663: inst = 32'hca0d373;
      119664: inst = 32'h13e00001;
      119665: inst = 32'hfe0d96a;
      119666: inst = 32'h5be00000;
      119667: inst = 32'h8c50000;
      119668: inst = 32'h24612800;
      119669: inst = 32'h10a00000;
      119670: inst = 32'hca0001e;
      119671: inst = 32'h24822800;
      119672: inst = 32'h10a00000;
      119673: inst = 32'hca00004;
      119674: inst = 32'h38632800;
      119675: inst = 32'h38842800;
      119676: inst = 32'h10a00001;
      119677: inst = 32'hca0d381;
      119678: inst = 32'h13e00001;
      119679: inst = 32'hfe0d96a;
      119680: inst = 32'h5be00000;
      119681: inst = 32'h8c50000;
      119682: inst = 32'h24612800;
      119683: inst = 32'h10a00000;
      119684: inst = 32'hca0001e;
      119685: inst = 32'h24822800;
      119686: inst = 32'h10a00000;
      119687: inst = 32'hca00004;
      119688: inst = 32'h38632800;
      119689: inst = 32'h38842800;
      119690: inst = 32'h10a00001;
      119691: inst = 32'hca0d38f;
      119692: inst = 32'h13e00001;
      119693: inst = 32'hfe0d96a;
      119694: inst = 32'h5be00000;
      119695: inst = 32'h8c50000;
      119696: inst = 32'h24612800;
      119697: inst = 32'h10a00000;
      119698: inst = 32'hca0001e;
      119699: inst = 32'h24822800;
      119700: inst = 32'h10a00000;
      119701: inst = 32'hca00004;
      119702: inst = 32'h38632800;
      119703: inst = 32'h38842800;
      119704: inst = 32'h10a00001;
      119705: inst = 32'hca0d39d;
      119706: inst = 32'h13e00001;
      119707: inst = 32'hfe0d96a;
      119708: inst = 32'h5be00000;
      119709: inst = 32'h8c50000;
      119710: inst = 32'h24612800;
      119711: inst = 32'h10a00000;
      119712: inst = 32'hca0001e;
      119713: inst = 32'h24822800;
      119714: inst = 32'h10a00000;
      119715: inst = 32'hca00004;
      119716: inst = 32'h38632800;
      119717: inst = 32'h38842800;
      119718: inst = 32'h10a00001;
      119719: inst = 32'hca0d3ab;
      119720: inst = 32'h13e00001;
      119721: inst = 32'hfe0d96a;
      119722: inst = 32'h5be00000;
      119723: inst = 32'h8c50000;
      119724: inst = 32'h24612800;
      119725: inst = 32'h10a00000;
      119726: inst = 32'hca0001e;
      119727: inst = 32'h24822800;
      119728: inst = 32'h10a00000;
      119729: inst = 32'hca00004;
      119730: inst = 32'h38632800;
      119731: inst = 32'h38842800;
      119732: inst = 32'h10a00001;
      119733: inst = 32'hca0d3b9;
      119734: inst = 32'h13e00001;
      119735: inst = 32'hfe0d96a;
      119736: inst = 32'h5be00000;
      119737: inst = 32'h8c50000;
      119738: inst = 32'h24612800;
      119739: inst = 32'h10a00000;
      119740: inst = 32'hca0001e;
      119741: inst = 32'h24822800;
      119742: inst = 32'h10a00000;
      119743: inst = 32'hca00004;
      119744: inst = 32'h38632800;
      119745: inst = 32'h38842800;
      119746: inst = 32'h10a00001;
      119747: inst = 32'hca0d3c7;
      119748: inst = 32'h13e00001;
      119749: inst = 32'hfe0d96a;
      119750: inst = 32'h5be00000;
      119751: inst = 32'h8c50000;
      119752: inst = 32'h24612800;
      119753: inst = 32'h10a00000;
      119754: inst = 32'hca0001e;
      119755: inst = 32'h24822800;
      119756: inst = 32'h10a00000;
      119757: inst = 32'hca00004;
      119758: inst = 32'h38632800;
      119759: inst = 32'h38842800;
      119760: inst = 32'h10a00001;
      119761: inst = 32'hca0d3d5;
      119762: inst = 32'h13e00001;
      119763: inst = 32'hfe0d96a;
      119764: inst = 32'h5be00000;
      119765: inst = 32'h8c50000;
      119766: inst = 32'h24612800;
      119767: inst = 32'h10a00000;
      119768: inst = 32'hca0001e;
      119769: inst = 32'h24822800;
      119770: inst = 32'h10a00000;
      119771: inst = 32'hca00004;
      119772: inst = 32'h38632800;
      119773: inst = 32'h38842800;
      119774: inst = 32'h10a00001;
      119775: inst = 32'hca0d3e3;
      119776: inst = 32'h13e00001;
      119777: inst = 32'hfe0d96a;
      119778: inst = 32'h5be00000;
      119779: inst = 32'h8c50000;
      119780: inst = 32'h24612800;
      119781: inst = 32'h10a00000;
      119782: inst = 32'hca0001e;
      119783: inst = 32'h24822800;
      119784: inst = 32'h10a00000;
      119785: inst = 32'hca00004;
      119786: inst = 32'h38632800;
      119787: inst = 32'h38842800;
      119788: inst = 32'h10a00001;
      119789: inst = 32'hca0d3f1;
      119790: inst = 32'h13e00001;
      119791: inst = 32'hfe0d96a;
      119792: inst = 32'h5be00000;
      119793: inst = 32'h8c50000;
      119794: inst = 32'h24612800;
      119795: inst = 32'h10a00000;
      119796: inst = 32'hca0001e;
      119797: inst = 32'h24822800;
      119798: inst = 32'h10a00000;
      119799: inst = 32'hca00004;
      119800: inst = 32'h38632800;
      119801: inst = 32'h38842800;
      119802: inst = 32'h10a00001;
      119803: inst = 32'hca0d3ff;
      119804: inst = 32'h13e00001;
      119805: inst = 32'hfe0d96a;
      119806: inst = 32'h5be00000;
      119807: inst = 32'h8c50000;
      119808: inst = 32'h24612800;
      119809: inst = 32'h10a00000;
      119810: inst = 32'hca0001e;
      119811: inst = 32'h24822800;
      119812: inst = 32'h10a00000;
      119813: inst = 32'hca00004;
      119814: inst = 32'h38632800;
      119815: inst = 32'h38842800;
      119816: inst = 32'h10a00001;
      119817: inst = 32'hca0d40d;
      119818: inst = 32'h13e00001;
      119819: inst = 32'hfe0d96a;
      119820: inst = 32'h5be00000;
      119821: inst = 32'h8c50000;
      119822: inst = 32'h24612800;
      119823: inst = 32'h10a00000;
      119824: inst = 32'hca0001e;
      119825: inst = 32'h24822800;
      119826: inst = 32'h10a00000;
      119827: inst = 32'hca00004;
      119828: inst = 32'h38632800;
      119829: inst = 32'h38842800;
      119830: inst = 32'h10a00001;
      119831: inst = 32'hca0d41b;
      119832: inst = 32'h13e00001;
      119833: inst = 32'hfe0d96a;
      119834: inst = 32'h5be00000;
      119835: inst = 32'h8c50000;
      119836: inst = 32'h24612800;
      119837: inst = 32'h10a00000;
      119838: inst = 32'hca0001e;
      119839: inst = 32'h24822800;
      119840: inst = 32'h10a00000;
      119841: inst = 32'hca00004;
      119842: inst = 32'h38632800;
      119843: inst = 32'h38842800;
      119844: inst = 32'h10a00001;
      119845: inst = 32'hca0d429;
      119846: inst = 32'h13e00001;
      119847: inst = 32'hfe0d96a;
      119848: inst = 32'h5be00000;
      119849: inst = 32'h8c50000;
      119850: inst = 32'h24612800;
      119851: inst = 32'h10a00000;
      119852: inst = 32'hca0001f;
      119853: inst = 32'h24822800;
      119854: inst = 32'h10a00000;
      119855: inst = 32'hca00004;
      119856: inst = 32'h38632800;
      119857: inst = 32'h38842800;
      119858: inst = 32'h10a00001;
      119859: inst = 32'hca0d437;
      119860: inst = 32'h13e00001;
      119861: inst = 32'hfe0d96a;
      119862: inst = 32'h5be00000;
      119863: inst = 32'h8c50000;
      119864: inst = 32'h24612800;
      119865: inst = 32'h10a00000;
      119866: inst = 32'hca0001f;
      119867: inst = 32'h24822800;
      119868: inst = 32'h10a00000;
      119869: inst = 32'hca00004;
      119870: inst = 32'h38632800;
      119871: inst = 32'h38842800;
      119872: inst = 32'h10a00001;
      119873: inst = 32'hca0d445;
      119874: inst = 32'h13e00001;
      119875: inst = 32'hfe0d96a;
      119876: inst = 32'h5be00000;
      119877: inst = 32'h8c50000;
      119878: inst = 32'h24612800;
      119879: inst = 32'h10a00000;
      119880: inst = 32'hca0001f;
      119881: inst = 32'h24822800;
      119882: inst = 32'h10a00000;
      119883: inst = 32'hca00004;
      119884: inst = 32'h38632800;
      119885: inst = 32'h38842800;
      119886: inst = 32'h10a00001;
      119887: inst = 32'hca0d453;
      119888: inst = 32'h13e00001;
      119889: inst = 32'hfe0d96a;
      119890: inst = 32'h5be00000;
      119891: inst = 32'h8c50000;
      119892: inst = 32'h24612800;
      119893: inst = 32'h10a00000;
      119894: inst = 32'hca0001f;
      119895: inst = 32'h24822800;
      119896: inst = 32'h10a00000;
      119897: inst = 32'hca00004;
      119898: inst = 32'h38632800;
      119899: inst = 32'h38842800;
      119900: inst = 32'h10a00001;
      119901: inst = 32'hca0d461;
      119902: inst = 32'h13e00001;
      119903: inst = 32'hfe0d96a;
      119904: inst = 32'h5be00000;
      119905: inst = 32'h8c50000;
      119906: inst = 32'h24612800;
      119907: inst = 32'h10a00000;
      119908: inst = 32'hca0001f;
      119909: inst = 32'h24822800;
      119910: inst = 32'h10a00000;
      119911: inst = 32'hca00004;
      119912: inst = 32'h38632800;
      119913: inst = 32'h38842800;
      119914: inst = 32'h10a00001;
      119915: inst = 32'hca0d46f;
      119916: inst = 32'h13e00001;
      119917: inst = 32'hfe0d96a;
      119918: inst = 32'h5be00000;
      119919: inst = 32'h8c50000;
      119920: inst = 32'h24612800;
      119921: inst = 32'h10a00000;
      119922: inst = 32'hca0001f;
      119923: inst = 32'h24822800;
      119924: inst = 32'h10a00000;
      119925: inst = 32'hca00004;
      119926: inst = 32'h38632800;
      119927: inst = 32'h38842800;
      119928: inst = 32'h10a00001;
      119929: inst = 32'hca0d47d;
      119930: inst = 32'h13e00001;
      119931: inst = 32'hfe0d96a;
      119932: inst = 32'h5be00000;
      119933: inst = 32'h8c50000;
      119934: inst = 32'h24612800;
      119935: inst = 32'h10a00000;
      119936: inst = 32'hca0001f;
      119937: inst = 32'h24822800;
      119938: inst = 32'h10a00000;
      119939: inst = 32'hca00004;
      119940: inst = 32'h38632800;
      119941: inst = 32'h38842800;
      119942: inst = 32'h10a00001;
      119943: inst = 32'hca0d48b;
      119944: inst = 32'h13e00001;
      119945: inst = 32'hfe0d96a;
      119946: inst = 32'h5be00000;
      119947: inst = 32'h8c50000;
      119948: inst = 32'h24612800;
      119949: inst = 32'h10a00000;
      119950: inst = 32'hca0001f;
      119951: inst = 32'h24822800;
      119952: inst = 32'h10a00000;
      119953: inst = 32'hca00004;
      119954: inst = 32'h38632800;
      119955: inst = 32'h38842800;
      119956: inst = 32'h10a00001;
      119957: inst = 32'hca0d499;
      119958: inst = 32'h13e00001;
      119959: inst = 32'hfe0d96a;
      119960: inst = 32'h5be00000;
      119961: inst = 32'h8c50000;
      119962: inst = 32'h24612800;
      119963: inst = 32'h10a00000;
      119964: inst = 32'hca0001f;
      119965: inst = 32'h24822800;
      119966: inst = 32'h10a00000;
      119967: inst = 32'hca00004;
      119968: inst = 32'h38632800;
      119969: inst = 32'h38842800;
      119970: inst = 32'h10a00001;
      119971: inst = 32'hca0d4a7;
      119972: inst = 32'h13e00001;
      119973: inst = 32'hfe0d96a;
      119974: inst = 32'h5be00000;
      119975: inst = 32'h8c50000;
      119976: inst = 32'h24612800;
      119977: inst = 32'h10a00000;
      119978: inst = 32'hca0001f;
      119979: inst = 32'h24822800;
      119980: inst = 32'h10a00000;
      119981: inst = 32'hca00004;
      119982: inst = 32'h38632800;
      119983: inst = 32'h38842800;
      119984: inst = 32'h10a00001;
      119985: inst = 32'hca0d4b5;
      119986: inst = 32'h13e00001;
      119987: inst = 32'hfe0d96a;
      119988: inst = 32'h5be00000;
      119989: inst = 32'h8c50000;
      119990: inst = 32'h24612800;
      119991: inst = 32'h10a00000;
      119992: inst = 32'hca0001f;
      119993: inst = 32'h24822800;
      119994: inst = 32'h10a00000;
      119995: inst = 32'hca00004;
      119996: inst = 32'h38632800;
      119997: inst = 32'h38842800;
      119998: inst = 32'h10a00001;
      119999: inst = 32'hca0d4c3;
      120000: inst = 32'h13e00001;
      120001: inst = 32'hfe0d96a;
      120002: inst = 32'h5be00000;
      120003: inst = 32'h8c50000;
      120004: inst = 32'h24612800;
      120005: inst = 32'h10a00000;
      120006: inst = 32'hca0001f;
      120007: inst = 32'h24822800;
      120008: inst = 32'h10a00000;
      120009: inst = 32'hca00004;
      120010: inst = 32'h38632800;
      120011: inst = 32'h38842800;
      120012: inst = 32'h10a00001;
      120013: inst = 32'hca0d4d1;
      120014: inst = 32'h13e00001;
      120015: inst = 32'hfe0d96a;
      120016: inst = 32'h5be00000;
      120017: inst = 32'h8c50000;
      120018: inst = 32'h24612800;
      120019: inst = 32'h10a00000;
      120020: inst = 32'hca0001f;
      120021: inst = 32'h24822800;
      120022: inst = 32'h10a00000;
      120023: inst = 32'hca00004;
      120024: inst = 32'h38632800;
      120025: inst = 32'h38842800;
      120026: inst = 32'h10a00001;
      120027: inst = 32'hca0d4df;
      120028: inst = 32'h13e00001;
      120029: inst = 32'hfe0d96a;
      120030: inst = 32'h5be00000;
      120031: inst = 32'h8c50000;
      120032: inst = 32'h24612800;
      120033: inst = 32'h10a00000;
      120034: inst = 32'hca0001f;
      120035: inst = 32'h24822800;
      120036: inst = 32'h10a00000;
      120037: inst = 32'hca00004;
      120038: inst = 32'h38632800;
      120039: inst = 32'h38842800;
      120040: inst = 32'h10a00001;
      120041: inst = 32'hca0d4ed;
      120042: inst = 32'h13e00001;
      120043: inst = 32'hfe0d96a;
      120044: inst = 32'h5be00000;
      120045: inst = 32'h8c50000;
      120046: inst = 32'h24612800;
      120047: inst = 32'h10a00000;
      120048: inst = 32'hca0001f;
      120049: inst = 32'h24822800;
      120050: inst = 32'h10a00000;
      120051: inst = 32'hca00004;
      120052: inst = 32'h38632800;
      120053: inst = 32'h38842800;
      120054: inst = 32'h10a00001;
      120055: inst = 32'hca0d4fb;
      120056: inst = 32'h13e00001;
      120057: inst = 32'hfe0d96a;
      120058: inst = 32'h5be00000;
      120059: inst = 32'h8c50000;
      120060: inst = 32'h24612800;
      120061: inst = 32'h10a00000;
      120062: inst = 32'hca0001f;
      120063: inst = 32'h24822800;
      120064: inst = 32'h10a00000;
      120065: inst = 32'hca00004;
      120066: inst = 32'h38632800;
      120067: inst = 32'h38842800;
      120068: inst = 32'h10a00001;
      120069: inst = 32'hca0d509;
      120070: inst = 32'h13e00001;
      120071: inst = 32'hfe0d96a;
      120072: inst = 32'h5be00000;
      120073: inst = 32'h8c50000;
      120074: inst = 32'h24612800;
      120075: inst = 32'h10a00000;
      120076: inst = 32'hca0001f;
      120077: inst = 32'h24822800;
      120078: inst = 32'h10a00000;
      120079: inst = 32'hca00004;
      120080: inst = 32'h38632800;
      120081: inst = 32'h38842800;
      120082: inst = 32'h10a00001;
      120083: inst = 32'hca0d517;
      120084: inst = 32'h13e00001;
      120085: inst = 32'hfe0d96a;
      120086: inst = 32'h5be00000;
      120087: inst = 32'h8c50000;
      120088: inst = 32'h24612800;
      120089: inst = 32'h10a00000;
      120090: inst = 32'hca0001f;
      120091: inst = 32'h24822800;
      120092: inst = 32'h10a00000;
      120093: inst = 32'hca00004;
      120094: inst = 32'h38632800;
      120095: inst = 32'h38842800;
      120096: inst = 32'h10a00001;
      120097: inst = 32'hca0d525;
      120098: inst = 32'h13e00001;
      120099: inst = 32'hfe0d96a;
      120100: inst = 32'h5be00000;
      120101: inst = 32'h8c50000;
      120102: inst = 32'h24612800;
      120103: inst = 32'h10a00000;
      120104: inst = 32'hca0001f;
      120105: inst = 32'h24822800;
      120106: inst = 32'h10a00000;
      120107: inst = 32'hca00004;
      120108: inst = 32'h38632800;
      120109: inst = 32'h38842800;
      120110: inst = 32'h10a00001;
      120111: inst = 32'hca0d533;
      120112: inst = 32'h13e00001;
      120113: inst = 32'hfe0d96a;
      120114: inst = 32'h5be00000;
      120115: inst = 32'h8c50000;
      120116: inst = 32'h24612800;
      120117: inst = 32'h10a00000;
      120118: inst = 32'hca0001f;
      120119: inst = 32'h24822800;
      120120: inst = 32'h10a00000;
      120121: inst = 32'hca00004;
      120122: inst = 32'h38632800;
      120123: inst = 32'h38842800;
      120124: inst = 32'h10a00001;
      120125: inst = 32'hca0d541;
      120126: inst = 32'h13e00001;
      120127: inst = 32'hfe0d96a;
      120128: inst = 32'h5be00000;
      120129: inst = 32'h8c50000;
      120130: inst = 32'h24612800;
      120131: inst = 32'h10a00000;
      120132: inst = 32'hca0001f;
      120133: inst = 32'h24822800;
      120134: inst = 32'h10a00000;
      120135: inst = 32'hca00004;
      120136: inst = 32'h38632800;
      120137: inst = 32'h38842800;
      120138: inst = 32'h10a00001;
      120139: inst = 32'hca0d54f;
      120140: inst = 32'h13e00001;
      120141: inst = 32'hfe0d96a;
      120142: inst = 32'h5be00000;
      120143: inst = 32'h8c50000;
      120144: inst = 32'h24612800;
      120145: inst = 32'h10a00000;
      120146: inst = 32'hca0001f;
      120147: inst = 32'h24822800;
      120148: inst = 32'h10a00000;
      120149: inst = 32'hca00004;
      120150: inst = 32'h38632800;
      120151: inst = 32'h38842800;
      120152: inst = 32'h10a00001;
      120153: inst = 32'hca0d55d;
      120154: inst = 32'h13e00001;
      120155: inst = 32'hfe0d96a;
      120156: inst = 32'h5be00000;
      120157: inst = 32'h8c50000;
      120158: inst = 32'h24612800;
      120159: inst = 32'h10a00000;
      120160: inst = 32'hca0001f;
      120161: inst = 32'h24822800;
      120162: inst = 32'h10a00000;
      120163: inst = 32'hca00004;
      120164: inst = 32'h38632800;
      120165: inst = 32'h38842800;
      120166: inst = 32'h10a00001;
      120167: inst = 32'hca0d56b;
      120168: inst = 32'h13e00001;
      120169: inst = 32'hfe0d96a;
      120170: inst = 32'h5be00000;
      120171: inst = 32'h8c50000;
      120172: inst = 32'h24612800;
      120173: inst = 32'h10a00000;
      120174: inst = 32'hca0001f;
      120175: inst = 32'h24822800;
      120176: inst = 32'h10a00000;
      120177: inst = 32'hca00004;
      120178: inst = 32'h38632800;
      120179: inst = 32'h38842800;
      120180: inst = 32'h10a00001;
      120181: inst = 32'hca0d579;
      120182: inst = 32'h13e00001;
      120183: inst = 32'hfe0d96a;
      120184: inst = 32'h5be00000;
      120185: inst = 32'h8c50000;
      120186: inst = 32'h24612800;
      120187: inst = 32'h10a00000;
      120188: inst = 32'hca0001f;
      120189: inst = 32'h24822800;
      120190: inst = 32'h10a00000;
      120191: inst = 32'hca00004;
      120192: inst = 32'h38632800;
      120193: inst = 32'h38842800;
      120194: inst = 32'h10a00001;
      120195: inst = 32'hca0d587;
      120196: inst = 32'h13e00001;
      120197: inst = 32'hfe0d96a;
      120198: inst = 32'h5be00000;
      120199: inst = 32'h8c50000;
      120200: inst = 32'h24612800;
      120201: inst = 32'h10a00000;
      120202: inst = 32'hca0001f;
      120203: inst = 32'h24822800;
      120204: inst = 32'h10a00000;
      120205: inst = 32'hca00004;
      120206: inst = 32'h38632800;
      120207: inst = 32'h38842800;
      120208: inst = 32'h10a00001;
      120209: inst = 32'hca0d595;
      120210: inst = 32'h13e00001;
      120211: inst = 32'hfe0d96a;
      120212: inst = 32'h5be00000;
      120213: inst = 32'h8c50000;
      120214: inst = 32'h24612800;
      120215: inst = 32'h10a00000;
      120216: inst = 32'hca0001f;
      120217: inst = 32'h24822800;
      120218: inst = 32'h10a00000;
      120219: inst = 32'hca00004;
      120220: inst = 32'h38632800;
      120221: inst = 32'h38842800;
      120222: inst = 32'h10a00001;
      120223: inst = 32'hca0d5a3;
      120224: inst = 32'h13e00001;
      120225: inst = 32'hfe0d96a;
      120226: inst = 32'h5be00000;
      120227: inst = 32'h8c50000;
      120228: inst = 32'h24612800;
      120229: inst = 32'h10a00000;
      120230: inst = 32'hca0001f;
      120231: inst = 32'h24822800;
      120232: inst = 32'h10a00000;
      120233: inst = 32'hca00004;
      120234: inst = 32'h38632800;
      120235: inst = 32'h38842800;
      120236: inst = 32'h10a00001;
      120237: inst = 32'hca0d5b1;
      120238: inst = 32'h13e00001;
      120239: inst = 32'hfe0d96a;
      120240: inst = 32'h5be00000;
      120241: inst = 32'h8c50000;
      120242: inst = 32'h24612800;
      120243: inst = 32'h10a00000;
      120244: inst = 32'hca0001f;
      120245: inst = 32'h24822800;
      120246: inst = 32'h10a00000;
      120247: inst = 32'hca00004;
      120248: inst = 32'h38632800;
      120249: inst = 32'h38842800;
      120250: inst = 32'h10a00001;
      120251: inst = 32'hca0d5bf;
      120252: inst = 32'h13e00001;
      120253: inst = 32'hfe0d96a;
      120254: inst = 32'h5be00000;
      120255: inst = 32'h8c50000;
      120256: inst = 32'h24612800;
      120257: inst = 32'h10a00000;
      120258: inst = 32'hca0001f;
      120259: inst = 32'h24822800;
      120260: inst = 32'h10a00000;
      120261: inst = 32'hca00004;
      120262: inst = 32'h38632800;
      120263: inst = 32'h38842800;
      120264: inst = 32'h10a00001;
      120265: inst = 32'hca0d5cd;
      120266: inst = 32'h13e00001;
      120267: inst = 32'hfe0d96a;
      120268: inst = 32'h5be00000;
      120269: inst = 32'h8c50000;
      120270: inst = 32'h24612800;
      120271: inst = 32'h10a00000;
      120272: inst = 32'hca0001f;
      120273: inst = 32'h24822800;
      120274: inst = 32'h10a00000;
      120275: inst = 32'hca00004;
      120276: inst = 32'h38632800;
      120277: inst = 32'h38842800;
      120278: inst = 32'h10a00001;
      120279: inst = 32'hca0d5db;
      120280: inst = 32'h13e00001;
      120281: inst = 32'hfe0d96a;
      120282: inst = 32'h5be00000;
      120283: inst = 32'h8c50000;
      120284: inst = 32'h24612800;
      120285: inst = 32'h10a00000;
      120286: inst = 32'hca0001f;
      120287: inst = 32'h24822800;
      120288: inst = 32'h10a00000;
      120289: inst = 32'hca00004;
      120290: inst = 32'h38632800;
      120291: inst = 32'h38842800;
      120292: inst = 32'h10a00001;
      120293: inst = 32'hca0d5e9;
      120294: inst = 32'h13e00001;
      120295: inst = 32'hfe0d96a;
      120296: inst = 32'h5be00000;
      120297: inst = 32'h8c50000;
      120298: inst = 32'h24612800;
      120299: inst = 32'h10a00000;
      120300: inst = 32'hca0001f;
      120301: inst = 32'h24822800;
      120302: inst = 32'h10a00000;
      120303: inst = 32'hca00004;
      120304: inst = 32'h38632800;
      120305: inst = 32'h38842800;
      120306: inst = 32'h10a00001;
      120307: inst = 32'hca0d5f7;
      120308: inst = 32'h13e00001;
      120309: inst = 32'hfe0d96a;
      120310: inst = 32'h5be00000;
      120311: inst = 32'h8c50000;
      120312: inst = 32'h24612800;
      120313: inst = 32'h10a00000;
      120314: inst = 32'hca0001f;
      120315: inst = 32'h24822800;
      120316: inst = 32'h10a00000;
      120317: inst = 32'hca00004;
      120318: inst = 32'h38632800;
      120319: inst = 32'h38842800;
      120320: inst = 32'h10a00001;
      120321: inst = 32'hca0d605;
      120322: inst = 32'h13e00001;
      120323: inst = 32'hfe0d96a;
      120324: inst = 32'h5be00000;
      120325: inst = 32'h8c50000;
      120326: inst = 32'h24612800;
      120327: inst = 32'h10a00000;
      120328: inst = 32'hca0001f;
      120329: inst = 32'h24822800;
      120330: inst = 32'h10a00000;
      120331: inst = 32'hca00004;
      120332: inst = 32'h38632800;
      120333: inst = 32'h38842800;
      120334: inst = 32'h10a00001;
      120335: inst = 32'hca0d613;
      120336: inst = 32'h13e00001;
      120337: inst = 32'hfe0d96a;
      120338: inst = 32'h5be00000;
      120339: inst = 32'h8c50000;
      120340: inst = 32'h24612800;
      120341: inst = 32'h10a00000;
      120342: inst = 32'hca0001f;
      120343: inst = 32'h24822800;
      120344: inst = 32'h10a00000;
      120345: inst = 32'hca00004;
      120346: inst = 32'h38632800;
      120347: inst = 32'h38842800;
      120348: inst = 32'h10a00001;
      120349: inst = 32'hca0d621;
      120350: inst = 32'h13e00001;
      120351: inst = 32'hfe0d96a;
      120352: inst = 32'h5be00000;
      120353: inst = 32'h8c50000;
      120354: inst = 32'h24612800;
      120355: inst = 32'h10a00000;
      120356: inst = 32'hca0001f;
      120357: inst = 32'h24822800;
      120358: inst = 32'h10a00000;
      120359: inst = 32'hca00004;
      120360: inst = 32'h38632800;
      120361: inst = 32'h38842800;
      120362: inst = 32'h10a00001;
      120363: inst = 32'hca0d62f;
      120364: inst = 32'h13e00001;
      120365: inst = 32'hfe0d96a;
      120366: inst = 32'h5be00000;
      120367: inst = 32'h8c50000;
      120368: inst = 32'h24612800;
      120369: inst = 32'h10a00000;
      120370: inst = 32'hca0001f;
      120371: inst = 32'h24822800;
      120372: inst = 32'h10a00000;
      120373: inst = 32'hca00004;
      120374: inst = 32'h38632800;
      120375: inst = 32'h38842800;
      120376: inst = 32'h10a00001;
      120377: inst = 32'hca0d63d;
      120378: inst = 32'h13e00001;
      120379: inst = 32'hfe0d96a;
      120380: inst = 32'h5be00000;
      120381: inst = 32'h8c50000;
      120382: inst = 32'h24612800;
      120383: inst = 32'h10a00000;
      120384: inst = 32'hca0001f;
      120385: inst = 32'h24822800;
      120386: inst = 32'h10a00000;
      120387: inst = 32'hca00004;
      120388: inst = 32'h38632800;
      120389: inst = 32'h38842800;
      120390: inst = 32'h10a00001;
      120391: inst = 32'hca0d64b;
      120392: inst = 32'h13e00001;
      120393: inst = 32'hfe0d96a;
      120394: inst = 32'h5be00000;
      120395: inst = 32'h8c50000;
      120396: inst = 32'h24612800;
      120397: inst = 32'h10a00000;
      120398: inst = 32'hca0001f;
      120399: inst = 32'h24822800;
      120400: inst = 32'h10a00000;
      120401: inst = 32'hca00004;
      120402: inst = 32'h38632800;
      120403: inst = 32'h38842800;
      120404: inst = 32'h10a00001;
      120405: inst = 32'hca0d659;
      120406: inst = 32'h13e00001;
      120407: inst = 32'hfe0d96a;
      120408: inst = 32'h5be00000;
      120409: inst = 32'h8c50000;
      120410: inst = 32'h24612800;
      120411: inst = 32'h10a00000;
      120412: inst = 32'hca0001f;
      120413: inst = 32'h24822800;
      120414: inst = 32'h10a00000;
      120415: inst = 32'hca00004;
      120416: inst = 32'h38632800;
      120417: inst = 32'h38842800;
      120418: inst = 32'h10a00001;
      120419: inst = 32'hca0d667;
      120420: inst = 32'h13e00001;
      120421: inst = 32'hfe0d96a;
      120422: inst = 32'h5be00000;
      120423: inst = 32'h8c50000;
      120424: inst = 32'h24612800;
      120425: inst = 32'h10a00000;
      120426: inst = 32'hca0001f;
      120427: inst = 32'h24822800;
      120428: inst = 32'h10a00000;
      120429: inst = 32'hca00004;
      120430: inst = 32'h38632800;
      120431: inst = 32'h38842800;
      120432: inst = 32'h10a00001;
      120433: inst = 32'hca0d675;
      120434: inst = 32'h13e00001;
      120435: inst = 32'hfe0d96a;
      120436: inst = 32'h5be00000;
      120437: inst = 32'h8c50000;
      120438: inst = 32'h24612800;
      120439: inst = 32'h10a00000;
      120440: inst = 32'hca0001f;
      120441: inst = 32'h24822800;
      120442: inst = 32'h10a00000;
      120443: inst = 32'hca00004;
      120444: inst = 32'h38632800;
      120445: inst = 32'h38842800;
      120446: inst = 32'h10a00001;
      120447: inst = 32'hca0d683;
      120448: inst = 32'h13e00001;
      120449: inst = 32'hfe0d96a;
      120450: inst = 32'h5be00000;
      120451: inst = 32'h8c50000;
      120452: inst = 32'h24612800;
      120453: inst = 32'h10a00000;
      120454: inst = 32'hca0001f;
      120455: inst = 32'h24822800;
      120456: inst = 32'h10a00000;
      120457: inst = 32'hca00004;
      120458: inst = 32'h38632800;
      120459: inst = 32'h38842800;
      120460: inst = 32'h10a00001;
      120461: inst = 32'hca0d691;
      120462: inst = 32'h13e00001;
      120463: inst = 32'hfe0d96a;
      120464: inst = 32'h5be00000;
      120465: inst = 32'h8c50000;
      120466: inst = 32'h24612800;
      120467: inst = 32'h10a00000;
      120468: inst = 32'hca0001f;
      120469: inst = 32'h24822800;
      120470: inst = 32'h10a00000;
      120471: inst = 32'hca00004;
      120472: inst = 32'h38632800;
      120473: inst = 32'h38842800;
      120474: inst = 32'h10a00001;
      120475: inst = 32'hca0d69f;
      120476: inst = 32'h13e00001;
      120477: inst = 32'hfe0d96a;
      120478: inst = 32'h5be00000;
      120479: inst = 32'h8c50000;
      120480: inst = 32'h24612800;
      120481: inst = 32'h10a00000;
      120482: inst = 32'hca0001f;
      120483: inst = 32'h24822800;
      120484: inst = 32'h10a00000;
      120485: inst = 32'hca00004;
      120486: inst = 32'h38632800;
      120487: inst = 32'h38842800;
      120488: inst = 32'h10a00001;
      120489: inst = 32'hca0d6ad;
      120490: inst = 32'h13e00001;
      120491: inst = 32'hfe0d96a;
      120492: inst = 32'h5be00000;
      120493: inst = 32'h8c50000;
      120494: inst = 32'h24612800;
      120495: inst = 32'h10a00000;
      120496: inst = 32'hca0001f;
      120497: inst = 32'h24822800;
      120498: inst = 32'h10a00000;
      120499: inst = 32'hca00004;
      120500: inst = 32'h38632800;
      120501: inst = 32'h38842800;
      120502: inst = 32'h10a00001;
      120503: inst = 32'hca0d6bb;
      120504: inst = 32'h13e00001;
      120505: inst = 32'hfe0d96a;
      120506: inst = 32'h5be00000;
      120507: inst = 32'h8c50000;
      120508: inst = 32'h24612800;
      120509: inst = 32'h10a00000;
      120510: inst = 32'hca0001f;
      120511: inst = 32'h24822800;
      120512: inst = 32'h10a00000;
      120513: inst = 32'hca00004;
      120514: inst = 32'h38632800;
      120515: inst = 32'h38842800;
      120516: inst = 32'h10a00001;
      120517: inst = 32'hca0d6c9;
      120518: inst = 32'h13e00001;
      120519: inst = 32'hfe0d96a;
      120520: inst = 32'h5be00000;
      120521: inst = 32'h8c50000;
      120522: inst = 32'h24612800;
      120523: inst = 32'h10a00000;
      120524: inst = 32'hca0001f;
      120525: inst = 32'h24822800;
      120526: inst = 32'h10a00000;
      120527: inst = 32'hca00004;
      120528: inst = 32'h38632800;
      120529: inst = 32'h38842800;
      120530: inst = 32'h10a00001;
      120531: inst = 32'hca0d6d7;
      120532: inst = 32'h13e00001;
      120533: inst = 32'hfe0d96a;
      120534: inst = 32'h5be00000;
      120535: inst = 32'h8c50000;
      120536: inst = 32'h24612800;
      120537: inst = 32'h10a00000;
      120538: inst = 32'hca0001f;
      120539: inst = 32'h24822800;
      120540: inst = 32'h10a00000;
      120541: inst = 32'hca00004;
      120542: inst = 32'h38632800;
      120543: inst = 32'h38842800;
      120544: inst = 32'h10a00001;
      120545: inst = 32'hca0d6e5;
      120546: inst = 32'h13e00001;
      120547: inst = 32'hfe0d96a;
      120548: inst = 32'h5be00000;
      120549: inst = 32'h8c50000;
      120550: inst = 32'h24612800;
      120551: inst = 32'h10a00000;
      120552: inst = 32'hca0001f;
      120553: inst = 32'h24822800;
      120554: inst = 32'h10a00000;
      120555: inst = 32'hca00004;
      120556: inst = 32'h38632800;
      120557: inst = 32'h38842800;
      120558: inst = 32'h10a00001;
      120559: inst = 32'hca0d6f3;
      120560: inst = 32'h13e00001;
      120561: inst = 32'hfe0d96a;
      120562: inst = 32'h5be00000;
      120563: inst = 32'h8c50000;
      120564: inst = 32'h24612800;
      120565: inst = 32'h10a00000;
      120566: inst = 32'hca0001f;
      120567: inst = 32'h24822800;
      120568: inst = 32'h10a00000;
      120569: inst = 32'hca00004;
      120570: inst = 32'h38632800;
      120571: inst = 32'h38842800;
      120572: inst = 32'h10a00001;
      120573: inst = 32'hca0d701;
      120574: inst = 32'h13e00001;
      120575: inst = 32'hfe0d96a;
      120576: inst = 32'h5be00000;
      120577: inst = 32'h8c50000;
      120578: inst = 32'h24612800;
      120579: inst = 32'h10a00000;
      120580: inst = 32'hca0001f;
      120581: inst = 32'h24822800;
      120582: inst = 32'h10a00000;
      120583: inst = 32'hca00004;
      120584: inst = 32'h38632800;
      120585: inst = 32'h38842800;
      120586: inst = 32'h10a00001;
      120587: inst = 32'hca0d70f;
      120588: inst = 32'h13e00001;
      120589: inst = 32'hfe0d96a;
      120590: inst = 32'h5be00000;
      120591: inst = 32'h8c50000;
      120592: inst = 32'h24612800;
      120593: inst = 32'h10a00000;
      120594: inst = 32'hca0001f;
      120595: inst = 32'h24822800;
      120596: inst = 32'h10a00000;
      120597: inst = 32'hca00004;
      120598: inst = 32'h38632800;
      120599: inst = 32'h38842800;
      120600: inst = 32'h10a00001;
      120601: inst = 32'hca0d71d;
      120602: inst = 32'h13e00001;
      120603: inst = 32'hfe0d96a;
      120604: inst = 32'h5be00000;
      120605: inst = 32'h8c50000;
      120606: inst = 32'h24612800;
      120607: inst = 32'h10a00000;
      120608: inst = 32'hca0001f;
      120609: inst = 32'h24822800;
      120610: inst = 32'h10a00000;
      120611: inst = 32'hca00004;
      120612: inst = 32'h38632800;
      120613: inst = 32'h38842800;
      120614: inst = 32'h10a00001;
      120615: inst = 32'hca0d72b;
      120616: inst = 32'h13e00001;
      120617: inst = 32'hfe0d96a;
      120618: inst = 32'h5be00000;
      120619: inst = 32'h8c50000;
      120620: inst = 32'h24612800;
      120621: inst = 32'h10a00000;
      120622: inst = 32'hca0001f;
      120623: inst = 32'h24822800;
      120624: inst = 32'h10a00000;
      120625: inst = 32'hca00004;
      120626: inst = 32'h38632800;
      120627: inst = 32'h38842800;
      120628: inst = 32'h10a00001;
      120629: inst = 32'hca0d739;
      120630: inst = 32'h13e00001;
      120631: inst = 32'hfe0d96a;
      120632: inst = 32'h5be00000;
      120633: inst = 32'h8c50000;
      120634: inst = 32'h24612800;
      120635: inst = 32'h10a00000;
      120636: inst = 32'hca0001f;
      120637: inst = 32'h24822800;
      120638: inst = 32'h10a00000;
      120639: inst = 32'hca00004;
      120640: inst = 32'h38632800;
      120641: inst = 32'h38842800;
      120642: inst = 32'h10a00001;
      120643: inst = 32'hca0d747;
      120644: inst = 32'h13e00001;
      120645: inst = 32'hfe0d96a;
      120646: inst = 32'h5be00000;
      120647: inst = 32'h8c50000;
      120648: inst = 32'h24612800;
      120649: inst = 32'h10a00000;
      120650: inst = 32'hca0001f;
      120651: inst = 32'h24822800;
      120652: inst = 32'h10a00000;
      120653: inst = 32'hca00004;
      120654: inst = 32'h38632800;
      120655: inst = 32'h38842800;
      120656: inst = 32'h10a00001;
      120657: inst = 32'hca0d755;
      120658: inst = 32'h13e00001;
      120659: inst = 32'hfe0d96a;
      120660: inst = 32'h5be00000;
      120661: inst = 32'h8c50000;
      120662: inst = 32'h24612800;
      120663: inst = 32'h10a00000;
      120664: inst = 32'hca0001f;
      120665: inst = 32'h24822800;
      120666: inst = 32'h10a00000;
      120667: inst = 32'hca00004;
      120668: inst = 32'h38632800;
      120669: inst = 32'h38842800;
      120670: inst = 32'h10a00001;
      120671: inst = 32'hca0d763;
      120672: inst = 32'h13e00001;
      120673: inst = 32'hfe0d96a;
      120674: inst = 32'h5be00000;
      120675: inst = 32'h8c50000;
      120676: inst = 32'h24612800;
      120677: inst = 32'h10a00000;
      120678: inst = 32'hca0001f;
      120679: inst = 32'h24822800;
      120680: inst = 32'h10a00000;
      120681: inst = 32'hca00004;
      120682: inst = 32'h38632800;
      120683: inst = 32'h38842800;
      120684: inst = 32'h10a00001;
      120685: inst = 32'hca0d771;
      120686: inst = 32'h13e00001;
      120687: inst = 32'hfe0d96a;
      120688: inst = 32'h5be00000;
      120689: inst = 32'h8c50000;
      120690: inst = 32'h24612800;
      120691: inst = 32'h10a00000;
      120692: inst = 32'hca0001f;
      120693: inst = 32'h24822800;
      120694: inst = 32'h10a00000;
      120695: inst = 32'hca00004;
      120696: inst = 32'h38632800;
      120697: inst = 32'h38842800;
      120698: inst = 32'h10a00001;
      120699: inst = 32'hca0d77f;
      120700: inst = 32'h13e00001;
      120701: inst = 32'hfe0d96a;
      120702: inst = 32'h5be00000;
      120703: inst = 32'h8c50000;
      120704: inst = 32'h24612800;
      120705: inst = 32'h10a00000;
      120706: inst = 32'hca0001f;
      120707: inst = 32'h24822800;
      120708: inst = 32'h10a00000;
      120709: inst = 32'hca00004;
      120710: inst = 32'h38632800;
      120711: inst = 32'h38842800;
      120712: inst = 32'h10a00001;
      120713: inst = 32'hca0d78d;
      120714: inst = 32'h13e00001;
      120715: inst = 32'hfe0d96a;
      120716: inst = 32'h5be00000;
      120717: inst = 32'h8c50000;
      120718: inst = 32'h24612800;
      120719: inst = 32'h10a00000;
      120720: inst = 32'hca0001f;
      120721: inst = 32'h24822800;
      120722: inst = 32'h10a00000;
      120723: inst = 32'hca00004;
      120724: inst = 32'h38632800;
      120725: inst = 32'h38842800;
      120726: inst = 32'h10a00001;
      120727: inst = 32'hca0d79b;
      120728: inst = 32'h13e00001;
      120729: inst = 32'hfe0d96a;
      120730: inst = 32'h5be00000;
      120731: inst = 32'h8c50000;
      120732: inst = 32'h24612800;
      120733: inst = 32'h10a00000;
      120734: inst = 32'hca0001f;
      120735: inst = 32'h24822800;
      120736: inst = 32'h10a00000;
      120737: inst = 32'hca00004;
      120738: inst = 32'h38632800;
      120739: inst = 32'h38842800;
      120740: inst = 32'h10a00001;
      120741: inst = 32'hca0d7a9;
      120742: inst = 32'h13e00001;
      120743: inst = 32'hfe0d96a;
      120744: inst = 32'h5be00000;
      120745: inst = 32'h8c50000;
      120746: inst = 32'h24612800;
      120747: inst = 32'h10a00000;
      120748: inst = 32'hca0001f;
      120749: inst = 32'h24822800;
      120750: inst = 32'h10a00000;
      120751: inst = 32'hca00004;
      120752: inst = 32'h38632800;
      120753: inst = 32'h38842800;
      120754: inst = 32'h10a00001;
      120755: inst = 32'hca0d7b7;
      120756: inst = 32'h13e00001;
      120757: inst = 32'hfe0d96a;
      120758: inst = 32'h5be00000;
      120759: inst = 32'h8c50000;
      120760: inst = 32'h24612800;
      120761: inst = 32'h10a00000;
      120762: inst = 32'hca0001f;
      120763: inst = 32'h24822800;
      120764: inst = 32'h10a00000;
      120765: inst = 32'hca00004;
      120766: inst = 32'h38632800;
      120767: inst = 32'h38842800;
      120768: inst = 32'h10a00001;
      120769: inst = 32'hca0d7c5;
      120770: inst = 32'h13e00001;
      120771: inst = 32'hfe0d96a;
      120772: inst = 32'h5be00000;
      120773: inst = 32'h8c50000;
      120774: inst = 32'h24612800;
      120775: inst = 32'h10a00000;
      120776: inst = 32'hca0001f;
      120777: inst = 32'h24822800;
      120778: inst = 32'h10a00000;
      120779: inst = 32'hca00004;
      120780: inst = 32'h38632800;
      120781: inst = 32'h38842800;
      120782: inst = 32'h10a00001;
      120783: inst = 32'hca0d7d3;
      120784: inst = 32'h13e00001;
      120785: inst = 32'hfe0d96a;
      120786: inst = 32'h5be00000;
      120787: inst = 32'h8c50000;
      120788: inst = 32'h24612800;
      120789: inst = 32'h10a00000;
      120790: inst = 32'hca0001f;
      120791: inst = 32'h24822800;
      120792: inst = 32'h10a00000;
      120793: inst = 32'hca00004;
      120794: inst = 32'h38632800;
      120795: inst = 32'h38842800;
      120796: inst = 32'h10a00001;
      120797: inst = 32'hca0d7e1;
      120798: inst = 32'h13e00001;
      120799: inst = 32'hfe0d96a;
      120800: inst = 32'h5be00000;
      120801: inst = 32'h8c50000;
      120802: inst = 32'h24612800;
      120803: inst = 32'h10a00000;
      120804: inst = 32'hca0001f;
      120805: inst = 32'h24822800;
      120806: inst = 32'h10a00000;
      120807: inst = 32'hca00004;
      120808: inst = 32'h38632800;
      120809: inst = 32'h38842800;
      120810: inst = 32'h10a00001;
      120811: inst = 32'hca0d7ef;
      120812: inst = 32'h13e00001;
      120813: inst = 32'hfe0d96a;
      120814: inst = 32'h5be00000;
      120815: inst = 32'h8c50000;
      120816: inst = 32'h24612800;
      120817: inst = 32'h10a00000;
      120818: inst = 32'hca0001f;
      120819: inst = 32'h24822800;
      120820: inst = 32'h10a00000;
      120821: inst = 32'hca00004;
      120822: inst = 32'h38632800;
      120823: inst = 32'h38842800;
      120824: inst = 32'h10a00001;
      120825: inst = 32'hca0d7fd;
      120826: inst = 32'h13e00001;
      120827: inst = 32'hfe0d96a;
      120828: inst = 32'h5be00000;
      120829: inst = 32'h8c50000;
      120830: inst = 32'h24612800;
      120831: inst = 32'h10a00000;
      120832: inst = 32'hca0001f;
      120833: inst = 32'h24822800;
      120834: inst = 32'h10a00000;
      120835: inst = 32'hca00004;
      120836: inst = 32'h38632800;
      120837: inst = 32'h38842800;
      120838: inst = 32'h10a00001;
      120839: inst = 32'hca0d80b;
      120840: inst = 32'h13e00001;
      120841: inst = 32'hfe0d96a;
      120842: inst = 32'h5be00000;
      120843: inst = 32'h8c50000;
      120844: inst = 32'h24612800;
      120845: inst = 32'h10a00000;
      120846: inst = 32'hca0001f;
      120847: inst = 32'h24822800;
      120848: inst = 32'h10a00000;
      120849: inst = 32'hca00004;
      120850: inst = 32'h38632800;
      120851: inst = 32'h38842800;
      120852: inst = 32'h10a00001;
      120853: inst = 32'hca0d819;
      120854: inst = 32'h13e00001;
      120855: inst = 32'hfe0d96a;
      120856: inst = 32'h5be00000;
      120857: inst = 32'h8c50000;
      120858: inst = 32'h24612800;
      120859: inst = 32'h10a00000;
      120860: inst = 32'hca0001f;
      120861: inst = 32'h24822800;
      120862: inst = 32'h10a00000;
      120863: inst = 32'hca00004;
      120864: inst = 32'h38632800;
      120865: inst = 32'h38842800;
      120866: inst = 32'h10a00001;
      120867: inst = 32'hca0d827;
      120868: inst = 32'h13e00001;
      120869: inst = 32'hfe0d96a;
      120870: inst = 32'h5be00000;
      120871: inst = 32'h8c50000;
      120872: inst = 32'h24612800;
      120873: inst = 32'h10a00000;
      120874: inst = 32'hca0001f;
      120875: inst = 32'h24822800;
      120876: inst = 32'h10a00000;
      120877: inst = 32'hca00004;
      120878: inst = 32'h38632800;
      120879: inst = 32'h38842800;
      120880: inst = 32'h10a00001;
      120881: inst = 32'hca0d835;
      120882: inst = 32'h13e00001;
      120883: inst = 32'hfe0d96a;
      120884: inst = 32'h5be00000;
      120885: inst = 32'h8c50000;
      120886: inst = 32'h24612800;
      120887: inst = 32'h10a00000;
      120888: inst = 32'hca0001f;
      120889: inst = 32'h24822800;
      120890: inst = 32'h10a00000;
      120891: inst = 32'hca00004;
      120892: inst = 32'h38632800;
      120893: inst = 32'h38842800;
      120894: inst = 32'h10a00001;
      120895: inst = 32'hca0d843;
      120896: inst = 32'h13e00001;
      120897: inst = 32'hfe0d96a;
      120898: inst = 32'h5be00000;
      120899: inst = 32'h8c50000;
      120900: inst = 32'h24612800;
      120901: inst = 32'h10a00000;
      120902: inst = 32'hca0001f;
      120903: inst = 32'h24822800;
      120904: inst = 32'h10a00000;
      120905: inst = 32'hca00004;
      120906: inst = 32'h38632800;
      120907: inst = 32'h38842800;
      120908: inst = 32'h10a00001;
      120909: inst = 32'hca0d851;
      120910: inst = 32'h13e00001;
      120911: inst = 32'hfe0d96a;
      120912: inst = 32'h5be00000;
      120913: inst = 32'h8c50000;
      120914: inst = 32'h24612800;
      120915: inst = 32'h10a00000;
      120916: inst = 32'hca0001f;
      120917: inst = 32'h24822800;
      120918: inst = 32'h10a00000;
      120919: inst = 32'hca00004;
      120920: inst = 32'h38632800;
      120921: inst = 32'h38842800;
      120922: inst = 32'h10a00001;
      120923: inst = 32'hca0d85f;
      120924: inst = 32'h13e00001;
      120925: inst = 32'hfe0d96a;
      120926: inst = 32'h5be00000;
      120927: inst = 32'h8c50000;
      120928: inst = 32'h24612800;
      120929: inst = 32'h10a00000;
      120930: inst = 32'hca0001f;
      120931: inst = 32'h24822800;
      120932: inst = 32'h10a00000;
      120933: inst = 32'hca00004;
      120934: inst = 32'h38632800;
      120935: inst = 32'h38842800;
      120936: inst = 32'h10a00001;
      120937: inst = 32'hca0d86d;
      120938: inst = 32'h13e00001;
      120939: inst = 32'hfe0d96a;
      120940: inst = 32'h5be00000;
      120941: inst = 32'h8c50000;
      120942: inst = 32'h24612800;
      120943: inst = 32'h10a00000;
      120944: inst = 32'hca0001f;
      120945: inst = 32'h24822800;
      120946: inst = 32'h10a00000;
      120947: inst = 32'hca00004;
      120948: inst = 32'h38632800;
      120949: inst = 32'h38842800;
      120950: inst = 32'h10a00001;
      120951: inst = 32'hca0d87b;
      120952: inst = 32'h13e00001;
      120953: inst = 32'hfe0d96a;
      120954: inst = 32'h5be00000;
      120955: inst = 32'h8c50000;
      120956: inst = 32'h24612800;
      120957: inst = 32'h10a00000;
      120958: inst = 32'hca0001f;
      120959: inst = 32'h24822800;
      120960: inst = 32'h10a00000;
      120961: inst = 32'hca00004;
      120962: inst = 32'h38632800;
      120963: inst = 32'h38842800;
      120964: inst = 32'h10a00001;
      120965: inst = 32'hca0d889;
      120966: inst = 32'h13e00001;
      120967: inst = 32'hfe0d96a;
      120968: inst = 32'h5be00000;
      120969: inst = 32'h8c50000;
      120970: inst = 32'h24612800;
      120971: inst = 32'h10a00000;
      120972: inst = 32'hca0001f;
      120973: inst = 32'h24822800;
      120974: inst = 32'h10a00000;
      120975: inst = 32'hca00004;
      120976: inst = 32'h38632800;
      120977: inst = 32'h38842800;
      120978: inst = 32'h10a00001;
      120979: inst = 32'hca0d897;
      120980: inst = 32'h13e00001;
      120981: inst = 32'hfe0d96a;
      120982: inst = 32'h5be00000;
      120983: inst = 32'h8c50000;
      120984: inst = 32'h24612800;
      120985: inst = 32'h10a00000;
      120986: inst = 32'hca0001f;
      120987: inst = 32'h24822800;
      120988: inst = 32'h10a00000;
      120989: inst = 32'hca00004;
      120990: inst = 32'h38632800;
      120991: inst = 32'h38842800;
      120992: inst = 32'h10a00001;
      120993: inst = 32'hca0d8a5;
      120994: inst = 32'h13e00001;
      120995: inst = 32'hfe0d96a;
      120996: inst = 32'h5be00000;
      120997: inst = 32'h8c50000;
      120998: inst = 32'h24612800;
      120999: inst = 32'h10a00000;
      121000: inst = 32'hca0001f;
      121001: inst = 32'h24822800;
      121002: inst = 32'h10a00000;
      121003: inst = 32'hca00004;
      121004: inst = 32'h38632800;
      121005: inst = 32'h38842800;
      121006: inst = 32'h10a00001;
      121007: inst = 32'hca0d8b3;
      121008: inst = 32'h13e00001;
      121009: inst = 32'hfe0d96a;
      121010: inst = 32'h5be00000;
      121011: inst = 32'h8c50000;
      121012: inst = 32'h24612800;
      121013: inst = 32'h10a00000;
      121014: inst = 32'hca0001f;
      121015: inst = 32'h24822800;
      121016: inst = 32'h10a00000;
      121017: inst = 32'hca00004;
      121018: inst = 32'h38632800;
      121019: inst = 32'h38842800;
      121020: inst = 32'h10a00001;
      121021: inst = 32'hca0d8c1;
      121022: inst = 32'h13e00001;
      121023: inst = 32'hfe0d96a;
      121024: inst = 32'h5be00000;
      121025: inst = 32'h8c50000;
      121026: inst = 32'h24612800;
      121027: inst = 32'h10a00000;
      121028: inst = 32'hca0001f;
      121029: inst = 32'h24822800;
      121030: inst = 32'h10a00000;
      121031: inst = 32'hca00004;
      121032: inst = 32'h38632800;
      121033: inst = 32'h38842800;
      121034: inst = 32'h10a00001;
      121035: inst = 32'hca0d8cf;
      121036: inst = 32'h13e00001;
      121037: inst = 32'hfe0d96a;
      121038: inst = 32'h5be00000;
      121039: inst = 32'h8c50000;
      121040: inst = 32'h24612800;
      121041: inst = 32'h10a00000;
      121042: inst = 32'hca0001f;
      121043: inst = 32'h24822800;
      121044: inst = 32'h10a00000;
      121045: inst = 32'hca00004;
      121046: inst = 32'h38632800;
      121047: inst = 32'h38842800;
      121048: inst = 32'h10a00001;
      121049: inst = 32'hca0d8dd;
      121050: inst = 32'h13e00001;
      121051: inst = 32'hfe0d96a;
      121052: inst = 32'h5be00000;
      121053: inst = 32'h8c50000;
      121054: inst = 32'h24612800;
      121055: inst = 32'h10a00000;
      121056: inst = 32'hca0001f;
      121057: inst = 32'h24822800;
      121058: inst = 32'h10a00000;
      121059: inst = 32'hca00004;
      121060: inst = 32'h38632800;
      121061: inst = 32'h38842800;
      121062: inst = 32'h10a00001;
      121063: inst = 32'hca0d8eb;
      121064: inst = 32'h13e00001;
      121065: inst = 32'hfe0d96a;
      121066: inst = 32'h5be00000;
      121067: inst = 32'h8c50000;
      121068: inst = 32'h24612800;
      121069: inst = 32'h10a00000;
      121070: inst = 32'hca0001f;
      121071: inst = 32'h24822800;
      121072: inst = 32'h10a00000;
      121073: inst = 32'hca00004;
      121074: inst = 32'h38632800;
      121075: inst = 32'h38842800;
      121076: inst = 32'h10a00001;
      121077: inst = 32'hca0d8f9;
      121078: inst = 32'h13e00001;
      121079: inst = 32'hfe0d96a;
      121080: inst = 32'h5be00000;
      121081: inst = 32'h8c50000;
      121082: inst = 32'h24612800;
      121083: inst = 32'h10a00000;
      121084: inst = 32'hca0001f;
      121085: inst = 32'h24822800;
      121086: inst = 32'h10a00000;
      121087: inst = 32'hca00004;
      121088: inst = 32'h38632800;
      121089: inst = 32'h38842800;
      121090: inst = 32'h10a00001;
      121091: inst = 32'hca0d907;
      121092: inst = 32'h13e00001;
      121093: inst = 32'hfe0d96a;
      121094: inst = 32'h5be00000;
      121095: inst = 32'h8c50000;
      121096: inst = 32'h24612800;
      121097: inst = 32'h10a00000;
      121098: inst = 32'hca0001f;
      121099: inst = 32'h24822800;
      121100: inst = 32'h10a00000;
      121101: inst = 32'hca00004;
      121102: inst = 32'h38632800;
      121103: inst = 32'h38842800;
      121104: inst = 32'h10a00001;
      121105: inst = 32'hca0d915;
      121106: inst = 32'h13e00001;
      121107: inst = 32'hfe0d96a;
      121108: inst = 32'h5be00000;
      121109: inst = 32'h8c50000;
      121110: inst = 32'h24612800;
      121111: inst = 32'h10a00000;
      121112: inst = 32'hca0001f;
      121113: inst = 32'h24822800;
      121114: inst = 32'h10a00000;
      121115: inst = 32'hca00004;
      121116: inst = 32'h38632800;
      121117: inst = 32'h38842800;
      121118: inst = 32'h10a00001;
      121119: inst = 32'hca0d923;
      121120: inst = 32'h13e00001;
      121121: inst = 32'hfe0d96a;
      121122: inst = 32'h5be00000;
      121123: inst = 32'h8c50000;
      121124: inst = 32'h24612800;
      121125: inst = 32'h10a00000;
      121126: inst = 32'hca0001f;
      121127: inst = 32'h24822800;
      121128: inst = 32'h10a00000;
      121129: inst = 32'hca00004;
      121130: inst = 32'h38632800;
      121131: inst = 32'h38842800;
      121132: inst = 32'h10a00001;
      121133: inst = 32'hca0d931;
      121134: inst = 32'h13e00001;
      121135: inst = 32'hfe0d96a;
      121136: inst = 32'h5be00000;
      121137: inst = 32'h8c50000;
      121138: inst = 32'h24612800;
      121139: inst = 32'h10a00000;
      121140: inst = 32'hca0001f;
      121141: inst = 32'h24822800;
      121142: inst = 32'h10a00000;
      121143: inst = 32'hca00004;
      121144: inst = 32'h38632800;
      121145: inst = 32'h38842800;
      121146: inst = 32'h10a00001;
      121147: inst = 32'hca0d93f;
      121148: inst = 32'h13e00001;
      121149: inst = 32'hfe0d96a;
      121150: inst = 32'h5be00000;
      121151: inst = 32'h8c50000;
      121152: inst = 32'h24612800;
      121153: inst = 32'h10a00000;
      121154: inst = 32'hca0001f;
      121155: inst = 32'h24822800;
      121156: inst = 32'h10a00000;
      121157: inst = 32'hca00004;
      121158: inst = 32'h38632800;
      121159: inst = 32'h38842800;
      121160: inst = 32'h10a00001;
      121161: inst = 32'hca0d94d;
      121162: inst = 32'h13e00001;
      121163: inst = 32'hfe0d96a;
      121164: inst = 32'h5be00000;
      121165: inst = 32'h8c50000;
      121166: inst = 32'h24612800;
      121167: inst = 32'h10a00000;
      121168: inst = 32'hca0001f;
      121169: inst = 32'h24822800;
      121170: inst = 32'h10a00000;
      121171: inst = 32'hca00004;
      121172: inst = 32'h38632800;
      121173: inst = 32'h38842800;
      121174: inst = 32'h10a00001;
      121175: inst = 32'hca0d95b;
      121176: inst = 32'h13e00001;
      121177: inst = 32'hfe0d96a;
      121178: inst = 32'h5be00000;
      121179: inst = 32'h8c50000;
      121180: inst = 32'h24612800;
      121181: inst = 32'h10a00000;
      121182: inst = 32'hca0001f;
      121183: inst = 32'h24822800;
      121184: inst = 32'h10a00000;
      121185: inst = 32'hca00004;
      121186: inst = 32'h38632800;
      121187: inst = 32'h38842800;
      121188: inst = 32'h10a00001;
      121189: inst = 32'hca0d969;
      121190: inst = 32'h13e00001;
      121191: inst = 32'hfe0d96a;
      121192: inst = 32'h5be00000;
      121193: inst = 32'h8c50000;
      121194: inst = 32'h13e0ffff;
      121195: inst = 32'h13e00001;
      121196: inst = 32'hfe0d9b7;
      121197: inst = 32'h5be00000;
      121198: inst = 32'h13e00001;
      121199: inst = 32'hfe0d9ed;
      121200: inst = 32'h5be00000;
      121201: inst = 32'h13e00001;
      121202: inst = 32'hfe0da23;
      121203: inst = 32'h5be00000;
      121204: inst = 32'h13e00001;
      121205: inst = 32'hfe0da59;
      121206: inst = 32'h5be00000;
      121207: inst = 32'h13e00001;
      121208: inst = 32'hfe0da8f;
      121209: inst = 32'h5be00000;
      121210: inst = 32'h13e00001;
      121211: inst = 32'hfe0dac5;
      121212: inst = 32'h5be00000;
      121213: inst = 32'h13e00001;
      121214: inst = 32'hfe0dafb;
      121215: inst = 32'h5be00000;
      121216: inst = 32'h13e00001;
      121217: inst = 32'hfe0db31;
      121218: inst = 32'h5be00000;
      121219: inst = 32'h13e00001;
      121220: inst = 32'hfe0db67;
      121221: inst = 32'h5be00000;
      121222: inst = 32'h13e00001;
      121223: inst = 32'hfe0db9d;
      121224: inst = 32'h5be00000;
      121225: inst = 32'h13e00001;
      121226: inst = 32'hfe0dbd3;
      121227: inst = 32'h5be00000;
      121228: inst = 32'h13e00001;
      121229: inst = 32'hfe0dc09;
      121230: inst = 32'h5be00000;
      121231: inst = 32'h13e00001;
      121232: inst = 32'hfe0dc3f;
      121233: inst = 32'h5be00000;
      121234: inst = 32'h13e00001;
      121235: inst = 32'hfe0dc75;
      121236: inst = 32'h5be00000;
      121237: inst = 32'h13e00001;
      121238: inst = 32'hfe0dcab;
      121239: inst = 32'h5be00000;
      121240: inst = 32'h13e00001;
      121241: inst = 32'hfe0dce1;
      121242: inst = 32'h5be00000;
      121243: inst = 32'h13e00001;
      121244: inst = 32'hfe0dd17;
      121245: inst = 32'h5be00000;
      121246: inst = 32'h13e00001;
      121247: inst = 32'hfe0dd4d;
      121248: inst = 32'h5be00000;
      121249: inst = 32'h13e00001;
      121250: inst = 32'hfe0dd83;
      121251: inst = 32'h5be00000;
      121252: inst = 32'h13e00001;
      121253: inst = 32'hfe0ddb9;
      121254: inst = 32'h5be00000;
      121255: inst = 32'h13e00001;
      121256: inst = 32'hfe0ddef;
      121257: inst = 32'h5be00000;
      121258: inst = 32'h13e00001;
      121259: inst = 32'hfe0de25;
      121260: inst = 32'h5be00000;
      121261: inst = 32'h13e00001;
      121262: inst = 32'hfe0de5b;
      121263: inst = 32'h5be00000;
      121264: inst = 32'h13e00001;
      121265: inst = 32'hfe0de91;
      121266: inst = 32'h5be00000;
      121267: inst = 32'h13e00001;
      121268: inst = 32'hfe0dec7;
      121269: inst = 32'h5be00000;
      121270: inst = 32'h58a00000;
      121271: inst = 32'h20800000;
      121272: inst = 32'h10c00000;
      121273: inst = 32'hcc06b50;
      121274: inst = 32'h20800001;
      121275: inst = 32'h10c00000;
      121276: inst = 32'hcc06b50;
      121277: inst = 32'h20800002;
      121278: inst = 32'h10c00000;
      121279: inst = 32'hcc06b50;
      121280: inst = 32'h20800003;
      121281: inst = 32'h10c00000;
      121282: inst = 32'hcc06b50;
      121283: inst = 32'h20800004;
      121284: inst = 32'h10c00000;
      121285: inst = 32'hcc06b50;
      121286: inst = 32'h20800005;
      121287: inst = 32'h10c00000;
      121288: inst = 32'hcc06b50;
      121289: inst = 32'h20800006;
      121290: inst = 32'h10c00000;
      121291: inst = 32'hcc06b50;
      121292: inst = 32'h20800007;
      121293: inst = 32'h10c00000;
      121294: inst = 32'hcc06b50;
      121295: inst = 32'h20800008;
      121296: inst = 32'h10c00000;
      121297: inst = 32'hcc06b50;
      121298: inst = 32'h20800009;
      121299: inst = 32'h10c00000;
      121300: inst = 32'hcc06b50;
      121301: inst = 32'h2080000a;
      121302: inst = 32'h10c00000;
      121303: inst = 32'hcc06b50;
      121304: inst = 32'h2080000b;
      121305: inst = 32'h10c00000;
      121306: inst = 32'hcc06b50;
      121307: inst = 32'h2080000c;
      121308: inst = 32'h10c00000;
      121309: inst = 32'hcc06b50;
      121310: inst = 32'h2080000d;
      121311: inst = 32'h10c00000;
      121312: inst = 32'hcc06b50;
      121313: inst = 32'h2080000e;
      121314: inst = 32'h10c00000;
      121315: inst = 32'hcc06b50;
      121316: inst = 32'h2080000f;
      121317: inst = 32'h10c00000;
      121318: inst = 32'hcc06b50;
      121319: inst = 32'h20800010;
      121320: inst = 32'h10c00000;
      121321: inst = 32'hcc06b50;
      121322: inst = 32'h20800011;
      121323: inst = 32'h10c00000;
      121324: inst = 32'hcc06b50;
      121325: inst = 32'h20800000;
      121326: inst = 32'h10c00000;
      121327: inst = 32'hcc06b50;
      121328: inst = 32'h20800001;
      121329: inst = 32'h10c00000;
      121330: inst = 32'hcc06b50;
      121331: inst = 32'h20800002;
      121332: inst = 32'h10c00000;
      121333: inst = 32'hcc06b50;
      121334: inst = 32'h20800003;
      121335: inst = 32'h10c00000;
      121336: inst = 32'hcc06b50;
      121337: inst = 32'h20800004;
      121338: inst = 32'h10c00000;
      121339: inst = 32'hcc06b50;
      121340: inst = 32'h20800005;
      121341: inst = 32'h10c00000;
      121342: inst = 32'hcc06b50;
      121343: inst = 32'h20800006;
      121344: inst = 32'h10c00000;
      121345: inst = 32'hcc06b50;
      121346: inst = 32'h20800007;
      121347: inst = 32'h10c00000;
      121348: inst = 32'hcc06b50;
      121349: inst = 32'h20800008;
      121350: inst = 32'h10c00000;
      121351: inst = 32'hcc06b50;
      121352: inst = 32'h20800009;
      121353: inst = 32'h10c00000;
      121354: inst = 32'hcc06b50;
      121355: inst = 32'h2080000a;
      121356: inst = 32'h10c00000;
      121357: inst = 32'hcc06b50;
      121358: inst = 32'h2080000b;
      121359: inst = 32'h10c00000;
      121360: inst = 32'hcc06b50;
      121361: inst = 32'h2080000c;
      121362: inst = 32'h10c00000;
      121363: inst = 32'hcc06b50;
      121364: inst = 32'h2080000d;
      121365: inst = 32'h10c00000;
      121366: inst = 32'hcc06b50;
      121367: inst = 32'h2080000e;
      121368: inst = 32'h10c00000;
      121369: inst = 32'hcc06b50;
      121370: inst = 32'h2080000f;
      121371: inst = 32'h10c00000;
      121372: inst = 32'hcc06b50;
      121373: inst = 32'h20800010;
      121374: inst = 32'h10c00000;
      121375: inst = 32'hcc06b50;
      121376: inst = 32'h20800011;
      121377: inst = 32'h10c00000;
      121378: inst = 32'hcc06b50;
      121379: inst = 32'h20800000;
      121380: inst = 32'h10c00000;
      121381: inst = 32'hcc06b50;
      121382: inst = 32'h20800001;
      121383: inst = 32'h10c00000;
      121384: inst = 32'hcc06b50;
      121385: inst = 32'h20800002;
      121386: inst = 32'h10c00000;
      121387: inst = 32'hcc06b50;
      121388: inst = 32'h20800003;
      121389: inst = 32'h10c00000;
      121390: inst = 32'hcc06b50;
      121391: inst = 32'h20800004;
      121392: inst = 32'h10c00000;
      121393: inst = 32'hcc06b50;
      121394: inst = 32'h20800005;
      121395: inst = 32'h10c00000;
      121396: inst = 32'hcc06b50;
      121397: inst = 32'h20800006;
      121398: inst = 32'h10c00000;
      121399: inst = 32'hcc06b50;
      121400: inst = 32'h20800007;
      121401: inst = 32'h10c00000;
      121402: inst = 32'hcc06b50;
      121403: inst = 32'h20800008;
      121404: inst = 32'h10c00000;
      121405: inst = 32'hcc06b50;
      121406: inst = 32'h20800009;
      121407: inst = 32'h10c00000;
      121408: inst = 32'hcc06b50;
      121409: inst = 32'h2080000a;
      121410: inst = 32'h10c00000;
      121411: inst = 32'hcc06b50;
      121412: inst = 32'h2080000b;
      121413: inst = 32'h10c00000;
      121414: inst = 32'hcc06b50;
      121415: inst = 32'h2080000c;
      121416: inst = 32'h10c00000;
      121417: inst = 32'hcc06b50;
      121418: inst = 32'h2080000d;
      121419: inst = 32'h10c00000;
      121420: inst = 32'hcc06b50;
      121421: inst = 32'h2080000e;
      121422: inst = 32'h10c00000;
      121423: inst = 32'hcc06b50;
      121424: inst = 32'h2080000f;
      121425: inst = 32'h10c00000;
      121426: inst = 32'hcc06b50;
      121427: inst = 32'h20800010;
      121428: inst = 32'h10c00000;
      121429: inst = 32'hcc06b50;
      121430: inst = 32'h20800011;
      121431: inst = 32'h10c00000;
      121432: inst = 32'hcc06b50;
      121433: inst = 32'h20800000;
      121434: inst = 32'h10c00000;
      121435: inst = 32'hcc06b50;
      121436: inst = 32'h20800001;
      121437: inst = 32'h10c00000;
      121438: inst = 32'hcc06b50;
      121439: inst = 32'h20800002;
      121440: inst = 32'h10c00000;
      121441: inst = 32'hcc06b50;
      121442: inst = 32'h20800003;
      121443: inst = 32'h10c00000;
      121444: inst = 32'hcc06b50;
      121445: inst = 32'h20800004;
      121446: inst = 32'h10c00000;
      121447: inst = 32'hcc06b50;
      121448: inst = 32'h20800005;
      121449: inst = 32'h10c00000;
      121450: inst = 32'hcc06b50;
      121451: inst = 32'h20800006;
      121452: inst = 32'h10c00000;
      121453: inst = 32'hcc06b50;
      121454: inst = 32'h20800007;
      121455: inst = 32'h10c00000;
      121456: inst = 32'hcc06b50;
      121457: inst = 32'h20800008;
      121458: inst = 32'h10c00000;
      121459: inst = 32'hcc06b50;
      121460: inst = 32'h20800009;
      121461: inst = 32'h10c00000;
      121462: inst = 32'hcc06b50;
      121463: inst = 32'h2080000a;
      121464: inst = 32'h10c00000;
      121465: inst = 32'hcc06b50;
      121466: inst = 32'h2080000b;
      121467: inst = 32'h10c00000;
      121468: inst = 32'hcc06b50;
      121469: inst = 32'h2080000c;
      121470: inst = 32'h10c00000;
      121471: inst = 32'hcc06b50;
      121472: inst = 32'h2080000d;
      121473: inst = 32'h10c00000;
      121474: inst = 32'hcc06b50;
      121475: inst = 32'h2080000e;
      121476: inst = 32'h10c00000;
      121477: inst = 32'hcc06b50;
      121478: inst = 32'h2080000f;
      121479: inst = 32'h10c00000;
      121480: inst = 32'hcc06b50;
      121481: inst = 32'h20800010;
      121482: inst = 32'h10c00000;
      121483: inst = 32'hcc06b50;
      121484: inst = 32'h20800011;
      121485: inst = 32'h10c00000;
      121486: inst = 32'hcc06b50;
      121487: inst = 32'h20800000;
      121488: inst = 32'h10c00000;
      121489: inst = 32'hcc06b50;
      121490: inst = 32'h20800001;
      121491: inst = 32'h10c00000;
      121492: inst = 32'hcc06b50;
      121493: inst = 32'h20800002;
      121494: inst = 32'h10c00000;
      121495: inst = 32'hcc06b50;
      121496: inst = 32'h20800003;
      121497: inst = 32'h10c00000;
      121498: inst = 32'hcc06b50;
      121499: inst = 32'h20800004;
      121500: inst = 32'h10c00000;
      121501: inst = 32'hcc06b50;
      121502: inst = 32'h20800005;
      121503: inst = 32'h10c00000;
      121504: inst = 32'hcc06b50;
      121505: inst = 32'h20800006;
      121506: inst = 32'h10c00000;
      121507: inst = 32'hcc06b50;
      121508: inst = 32'h20800007;
      121509: inst = 32'h10c00000;
      121510: inst = 32'hcc06b50;
      121511: inst = 32'h20800008;
      121512: inst = 32'h10c00000;
      121513: inst = 32'hcc06b50;
      121514: inst = 32'h20800009;
      121515: inst = 32'h10c00000;
      121516: inst = 32'hcc06b50;
      121517: inst = 32'h2080000a;
      121518: inst = 32'h10c00000;
      121519: inst = 32'hcc0eeb6;
      121520: inst = 32'h2080000b;
      121521: inst = 32'h10c00000;
      121522: inst = 32'hcc0eeb6;
      121523: inst = 32'h2080000c;
      121524: inst = 32'h10c00000;
      121525: inst = 32'hcc0eeb6;
      121526: inst = 32'h2080000d;
      121527: inst = 32'h10c00000;
      121528: inst = 32'hcc06b50;
      121529: inst = 32'h2080000e;
      121530: inst = 32'h10c00000;
      121531: inst = 32'hcc06b50;
      121532: inst = 32'h2080000f;
      121533: inst = 32'h10c00000;
      121534: inst = 32'hcc06b50;
      121535: inst = 32'h20800010;
      121536: inst = 32'h10c00000;
      121537: inst = 32'hcc06b50;
      121538: inst = 32'h20800011;
      121539: inst = 32'h10c00000;
      121540: inst = 32'hcc06b50;
      121541: inst = 32'h20800000;
      121542: inst = 32'h10c00000;
      121543: inst = 32'hcc06b50;
      121544: inst = 32'h20800001;
      121545: inst = 32'h10c00000;
      121546: inst = 32'hcc06b50;
      121547: inst = 32'h20800002;
      121548: inst = 32'h10c00000;
      121549: inst = 32'hcc06b50;
      121550: inst = 32'h20800003;
      121551: inst = 32'h10c00000;
      121552: inst = 32'hcc06b50;
      121553: inst = 32'h20800004;
      121554: inst = 32'h10c00000;
      121555: inst = 32'hcc06b50;
      121556: inst = 32'h20800005;
      121557: inst = 32'h10c00000;
      121558: inst = 32'hcc06b50;
      121559: inst = 32'h20800006;
      121560: inst = 32'h10c00000;
      121561: inst = 32'hcc06b50;
      121562: inst = 32'h20800007;
      121563: inst = 32'h10c00000;
      121564: inst = 32'hcc06b50;
      121565: inst = 32'h20800008;
      121566: inst = 32'h10c00000;
      121567: inst = 32'hcc06b50;
      121568: inst = 32'h20800009;
      121569: inst = 32'h10c00000;
      121570: inst = 32'hcc06b50;
      121571: inst = 32'h2080000a;
      121572: inst = 32'h10c00000;
      121573: inst = 32'hcc0eeb6;
      121574: inst = 32'h2080000b;
      121575: inst = 32'h10c00000;
      121576: inst = 32'hcc0eeb6;
      121577: inst = 32'h2080000c;
      121578: inst = 32'h10c00000;
      121579: inst = 32'hcc0eeb6;
      121580: inst = 32'h2080000d;
      121581: inst = 32'h10c00000;
      121582: inst = 32'hcc06b50;
      121583: inst = 32'h2080000e;
      121584: inst = 32'h10c00000;
      121585: inst = 32'hcc06b50;
      121586: inst = 32'h2080000f;
      121587: inst = 32'h10c00000;
      121588: inst = 32'hcc06b50;
      121589: inst = 32'h20800010;
      121590: inst = 32'h10c00000;
      121591: inst = 32'hcc06b50;
      121592: inst = 32'h20800011;
      121593: inst = 32'h10c00000;
      121594: inst = 32'hcc06b50;
      121595: inst = 32'h20800000;
      121596: inst = 32'h10c00000;
      121597: inst = 32'hcc06b50;
      121598: inst = 32'h20800001;
      121599: inst = 32'h10c00000;
      121600: inst = 32'hcc06b50;
      121601: inst = 32'h20800002;
      121602: inst = 32'h10c00000;
      121603: inst = 32'hcc06b50;
      121604: inst = 32'h20800003;
      121605: inst = 32'h10c00000;
      121606: inst = 32'hcc06b50;
      121607: inst = 32'h20800004;
      121608: inst = 32'h10c00000;
      121609: inst = 32'hcc06b50;
      121610: inst = 32'h20800005;
      121611: inst = 32'h10c00000;
      121612: inst = 32'hcc0eeb6;
      121613: inst = 32'h20800006;
      121614: inst = 32'h10c00000;
      121615: inst = 32'hcc0eeb6;
      121616: inst = 32'h20800007;
      121617: inst = 32'h10c00000;
      121618: inst = 32'hcc0eeb6;
      121619: inst = 32'h20800008;
      121620: inst = 32'h10c00000;
      121621: inst = 32'hcc06b50;
      121622: inst = 32'h20800009;
      121623: inst = 32'h10c00000;
      121624: inst = 32'hcc06b50;
      121625: inst = 32'h2080000a;
      121626: inst = 32'h10c00000;
      121627: inst = 32'hcc0eeb6;
      121628: inst = 32'h2080000b;
      121629: inst = 32'h10c00000;
      121630: inst = 32'hcc0eeb6;
      121631: inst = 32'h2080000c;
      121632: inst = 32'h10c00000;
      121633: inst = 32'hcc0eeb6;
      121634: inst = 32'h2080000d;
      121635: inst = 32'h10c00000;
      121636: inst = 32'hcc06b50;
      121637: inst = 32'h2080000e;
      121638: inst = 32'h10c00000;
      121639: inst = 32'hcc06b50;
      121640: inst = 32'h2080000f;
      121641: inst = 32'h10c00000;
      121642: inst = 32'hcc06b50;
      121643: inst = 32'h20800010;
      121644: inst = 32'h10c00000;
      121645: inst = 32'hcc06b50;
      121646: inst = 32'h20800011;
      121647: inst = 32'h10c00000;
      121648: inst = 32'hcc06b50;
      121649: inst = 32'h20800000;
      121650: inst = 32'h10c00000;
      121651: inst = 32'hcc06b50;
      121652: inst = 32'h20800001;
      121653: inst = 32'h10c00000;
      121654: inst = 32'hcc06b50;
      121655: inst = 32'h20800002;
      121656: inst = 32'h10c00000;
      121657: inst = 32'hcc06b50;
      121658: inst = 32'h20800003;
      121659: inst = 32'h10c00000;
      121660: inst = 32'hcc06b50;
      121661: inst = 32'h20800004;
      121662: inst = 32'h10c00000;
      121663: inst = 32'hcc06b50;
      121664: inst = 32'h20800005;
      121665: inst = 32'h10c00000;
      121666: inst = 32'hcc0eeb6;
      121667: inst = 32'h20800006;
      121668: inst = 32'h10c00000;
      121669: inst = 32'hcc0eeb6;
      121670: inst = 32'h20800007;
      121671: inst = 32'h10c00000;
      121672: inst = 32'hcc0eeb6;
      121673: inst = 32'h20800008;
      121674: inst = 32'h10c00000;
      121675: inst = 32'hcc06b50;
      121676: inst = 32'h20800009;
      121677: inst = 32'h10c00000;
      121678: inst = 32'hcc06b50;
      121679: inst = 32'h2080000a;
      121680: inst = 32'h10c00000;
      121681: inst = 32'hcc0eeb6;
      121682: inst = 32'h2080000b;
      121683: inst = 32'h10c00000;
      121684: inst = 32'hcc0eeb6;
      121685: inst = 32'h2080000c;
      121686: inst = 32'h10c00000;
      121687: inst = 32'hcc06b50;
      121688: inst = 32'h2080000d;
      121689: inst = 32'h10c00000;
      121690: inst = 32'hcc06b50;
      121691: inst = 32'h2080000e;
      121692: inst = 32'h10c00000;
      121693: inst = 32'hcc06b50;
      121694: inst = 32'h2080000f;
      121695: inst = 32'h10c00000;
      121696: inst = 32'hcc06b50;
      121697: inst = 32'h20800010;
      121698: inst = 32'h10c00000;
      121699: inst = 32'hcc06b50;
      121700: inst = 32'h20800011;
      121701: inst = 32'h10c00000;
      121702: inst = 32'hcc06b50;
      121703: inst = 32'h20800000;
      121704: inst = 32'h10c00000;
      121705: inst = 32'hcc06b50;
      121706: inst = 32'h20800001;
      121707: inst = 32'h10c00000;
      121708: inst = 32'hcc06b50;
      121709: inst = 32'h20800002;
      121710: inst = 32'h10c00000;
      121711: inst = 32'hcc06b50;
      121712: inst = 32'h20800003;
      121713: inst = 32'h10c00000;
      121714: inst = 32'hcc06b50;
      121715: inst = 32'h20800004;
      121716: inst = 32'h10c00000;
      121717: inst = 32'hcc06b50;
      121718: inst = 32'h20800005;
      121719: inst = 32'h10c00000;
      121720: inst = 32'hcc0eeb6;
      121721: inst = 32'h20800006;
      121722: inst = 32'h10c00000;
      121723: inst = 32'hcc0eeb6;
      121724: inst = 32'h20800007;
      121725: inst = 32'h10c00000;
      121726: inst = 32'hcc0eeb6;
      121727: inst = 32'h20800008;
      121728: inst = 32'h10c00000;
      121729: inst = 32'hcc0eeb6;
      121730: inst = 32'h20800009;
      121731: inst = 32'h10c00000;
      121732: inst = 32'hcc06b50;
      121733: inst = 32'h2080000a;
      121734: inst = 32'h10c00000;
      121735: inst = 32'hcc0eeb6;
      121736: inst = 32'h2080000b;
      121737: inst = 32'h10c00000;
      121738: inst = 32'hcc0eeb6;
      121739: inst = 32'h2080000c;
      121740: inst = 32'h10c00000;
      121741: inst = 32'hcc06b50;
      121742: inst = 32'h2080000d;
      121743: inst = 32'h10c00000;
      121744: inst = 32'hcc06b50;
      121745: inst = 32'h2080000e;
      121746: inst = 32'h10c00000;
      121747: inst = 32'hcc06b50;
      121748: inst = 32'h2080000f;
      121749: inst = 32'h10c00000;
      121750: inst = 32'hcc06b50;
      121751: inst = 32'h20800010;
      121752: inst = 32'h10c00000;
      121753: inst = 32'hcc06b50;
      121754: inst = 32'h20800011;
      121755: inst = 32'h10c00000;
      121756: inst = 32'hcc06b50;
      121757: inst = 32'h20800000;
      121758: inst = 32'h10c00000;
      121759: inst = 32'hcc06b50;
      121760: inst = 32'h20800001;
      121761: inst = 32'h10c00000;
      121762: inst = 32'hcc06b50;
      121763: inst = 32'h20800002;
      121764: inst = 32'h10c00000;
      121765: inst = 32'hcc06b50;
      121766: inst = 32'h20800003;
      121767: inst = 32'h10c00000;
      121768: inst = 32'hcc06b50;
      121769: inst = 32'h20800004;
      121770: inst = 32'h10c00000;
      121771: inst = 32'hcc06b50;
      121772: inst = 32'h20800005;
      121773: inst = 32'h10c00000;
      121774: inst = 32'hcc0eeb6;
      121775: inst = 32'h20800006;
      121776: inst = 32'h10c00000;
      121777: inst = 32'hcc0eeb6;
      121778: inst = 32'h20800007;
      121779: inst = 32'h10c00000;
      121780: inst = 32'hcc06b50;
      121781: inst = 32'h20800008;
      121782: inst = 32'h10c00000;
      121783: inst = 32'hcc0eeb6;
      121784: inst = 32'h20800009;
      121785: inst = 32'h10c00000;
      121786: inst = 32'hcc06b50;
      121787: inst = 32'h2080000a;
      121788: inst = 32'h10c00000;
      121789: inst = 32'hcc0eeb6;
      121790: inst = 32'h2080000b;
      121791: inst = 32'h10c00000;
      121792: inst = 32'hcc0eeb6;
      121793: inst = 32'h2080000c;
      121794: inst = 32'h10c00000;
      121795: inst = 32'hcc06b50;
      121796: inst = 32'h2080000d;
      121797: inst = 32'h10c00000;
      121798: inst = 32'hcc06b50;
      121799: inst = 32'h2080000e;
      121800: inst = 32'h10c00000;
      121801: inst = 32'hcc06b50;
      121802: inst = 32'h2080000f;
      121803: inst = 32'h10c00000;
      121804: inst = 32'hcc06b50;
      121805: inst = 32'h20800010;
      121806: inst = 32'h10c00000;
      121807: inst = 32'hcc06b50;
      121808: inst = 32'h20800011;
      121809: inst = 32'h10c00000;
      121810: inst = 32'hcc06b50;
      121811: inst = 32'h20800000;
      121812: inst = 32'h10c00000;
      121813: inst = 32'hcc06b50;
      121814: inst = 32'h20800001;
      121815: inst = 32'h10c00000;
      121816: inst = 32'hcc06b50;
      121817: inst = 32'h20800002;
      121818: inst = 32'h10c00000;
      121819: inst = 32'hcc06b50;
      121820: inst = 32'h20800003;
      121821: inst = 32'h10c00000;
      121822: inst = 32'hcc06b50;
      121823: inst = 32'h20800004;
      121824: inst = 32'h10c00000;
      121825: inst = 32'hcc06b50;
      121826: inst = 32'h20800005;
      121827: inst = 32'h10c00000;
      121828: inst = 32'hcc06b50;
      121829: inst = 32'h20800006;
      121830: inst = 32'h10c00000;
      121831: inst = 32'hcc0eeb6;
      121832: inst = 32'h20800007;
      121833: inst = 32'h10c00000;
      121834: inst = 32'hcc06b50;
      121835: inst = 32'h20800008;
      121836: inst = 32'h10c00000;
      121837: inst = 32'hcc0eeb6;
      121838: inst = 32'h20800009;
      121839: inst = 32'h10c00000;
      121840: inst = 32'hcc0eeb6;
      121841: inst = 32'h2080000a;
      121842: inst = 32'h10c00000;
      121843: inst = 32'hcc0eeb6;
      121844: inst = 32'h2080000b;
      121845: inst = 32'h10c00000;
      121846: inst = 32'hcc0eeb6;
      121847: inst = 32'h2080000c;
      121848: inst = 32'h10c00000;
      121849: inst = 32'hcc0eeb6;
      121850: inst = 32'h2080000d;
      121851: inst = 32'h10c00000;
      121852: inst = 32'hcc06b50;
      121853: inst = 32'h2080000e;
      121854: inst = 32'h10c00000;
      121855: inst = 32'hcc06b50;
      121856: inst = 32'h2080000f;
      121857: inst = 32'h10c00000;
      121858: inst = 32'hcc06b50;
      121859: inst = 32'h20800010;
      121860: inst = 32'h10c00000;
      121861: inst = 32'hcc06b50;
      121862: inst = 32'h20800011;
      121863: inst = 32'h10c00000;
      121864: inst = 32'hcc06b50;
      121865: inst = 32'h20800000;
      121866: inst = 32'h10c00000;
      121867: inst = 32'hcc06b50;
      121868: inst = 32'h20800001;
      121869: inst = 32'h10c00000;
      121870: inst = 32'hcc06b50;
      121871: inst = 32'h20800002;
      121872: inst = 32'h10c00000;
      121873: inst = 32'hcc06b50;
      121874: inst = 32'h20800003;
      121875: inst = 32'h10c00000;
      121876: inst = 32'hcc06b50;
      121877: inst = 32'h20800004;
      121878: inst = 32'h10c00000;
      121879: inst = 32'hcc06b50;
      121880: inst = 32'h20800005;
      121881: inst = 32'h10c00000;
      121882: inst = 32'hcc06b50;
      121883: inst = 32'h20800006;
      121884: inst = 32'h10c00000;
      121885: inst = 32'hcc0eeb6;
      121886: inst = 32'h20800007;
      121887: inst = 32'h10c00000;
      121888: inst = 32'hcc06b50;
      121889: inst = 32'h20800008;
      121890: inst = 32'h10c00000;
      121891: inst = 32'hcc0eeb6;
      121892: inst = 32'h20800009;
      121893: inst = 32'h10c00000;
      121894: inst = 32'hcc0eeb6;
      121895: inst = 32'h2080000a;
      121896: inst = 32'h10c00000;
      121897: inst = 32'hcc06b50;
      121898: inst = 32'h2080000b;
      121899: inst = 32'h10c00000;
      121900: inst = 32'hcc0eeb6;
      121901: inst = 32'h2080000c;
      121902: inst = 32'h10c00000;
      121903: inst = 32'hcc0eeb6;
      121904: inst = 32'h2080000d;
      121905: inst = 32'h10c00000;
      121906: inst = 32'hcc06b50;
      121907: inst = 32'h2080000e;
      121908: inst = 32'h10c00000;
      121909: inst = 32'hcc06b50;
      121910: inst = 32'h2080000f;
      121911: inst = 32'h10c00000;
      121912: inst = 32'hcc06b50;
      121913: inst = 32'h20800010;
      121914: inst = 32'h10c00000;
      121915: inst = 32'hcc06b50;
      121916: inst = 32'h20800011;
      121917: inst = 32'h10c00000;
      121918: inst = 32'hcc06b50;
      121919: inst = 32'h20800000;
      121920: inst = 32'h10c00000;
      121921: inst = 32'hcc06b50;
      121922: inst = 32'h20800001;
      121923: inst = 32'h10c00000;
      121924: inst = 32'hcc06b50;
      121925: inst = 32'h20800002;
      121926: inst = 32'h10c00000;
      121927: inst = 32'hcc06b50;
      121928: inst = 32'h20800003;
      121929: inst = 32'h10c00000;
      121930: inst = 32'hcc06b50;
      121931: inst = 32'h20800004;
      121932: inst = 32'h10c00000;
      121933: inst = 32'hcc06b50;
      121934: inst = 32'h20800005;
      121935: inst = 32'h10c00000;
      121936: inst = 32'hcc06b50;
      121937: inst = 32'h20800006;
      121938: inst = 32'h10c00000;
      121939: inst = 32'hcc0eeb6;
      121940: inst = 32'h20800007;
      121941: inst = 32'h10c00000;
      121942: inst = 32'hcc06b50;
      121943: inst = 32'h20800008;
      121944: inst = 32'h10c00000;
      121945: inst = 32'hcc0eeb6;
      121946: inst = 32'h20800009;
      121947: inst = 32'h10c00000;
      121948: inst = 32'hcc0eeb6;
      121949: inst = 32'h2080000a;
      121950: inst = 32'h10c00000;
      121951: inst = 32'hcc06b50;
      121952: inst = 32'h2080000b;
      121953: inst = 32'h10c00000;
      121954: inst = 32'hcc0eeb6;
      121955: inst = 32'h2080000c;
      121956: inst = 32'h10c00000;
      121957: inst = 32'hcc0eeb6;
      121958: inst = 32'h2080000d;
      121959: inst = 32'h10c00000;
      121960: inst = 32'hcc06b50;
      121961: inst = 32'h2080000e;
      121962: inst = 32'h10c00000;
      121963: inst = 32'hcc06b50;
      121964: inst = 32'h2080000f;
      121965: inst = 32'h10c00000;
      121966: inst = 32'hcc06b50;
      121967: inst = 32'h20800010;
      121968: inst = 32'h10c00000;
      121969: inst = 32'hcc06b50;
      121970: inst = 32'h20800011;
      121971: inst = 32'h10c00000;
      121972: inst = 32'hcc06b50;
      121973: inst = 32'h20800000;
      121974: inst = 32'h10c00000;
      121975: inst = 32'hcc06b50;
      121976: inst = 32'h20800001;
      121977: inst = 32'h10c00000;
      121978: inst = 32'hcc06b50;
      121979: inst = 32'h20800002;
      121980: inst = 32'h10c00000;
      121981: inst = 32'hcc06b50;
      121982: inst = 32'h20800003;
      121983: inst = 32'h10c00000;
      121984: inst = 32'hcc06b50;
      121985: inst = 32'h20800004;
      121986: inst = 32'h10c00000;
      121987: inst = 32'hcc06b50;
      121988: inst = 32'h20800005;
      121989: inst = 32'h10c00000;
      121990: inst = 32'hcc06b50;
      121991: inst = 32'h20800006;
      121992: inst = 32'h10c00000;
      121993: inst = 32'hcc0eeb6;
      121994: inst = 32'h20800007;
      121995: inst = 32'h10c00000;
      121996: inst = 32'hcc06b50;
      121997: inst = 32'h20800008;
      121998: inst = 32'h10c00000;
      121999: inst = 32'hcc0eeb6;
      122000: inst = 32'h20800009;
      122001: inst = 32'h10c00000;
      122002: inst = 32'hcc0eeb6;
      122003: inst = 32'h2080000a;
      122004: inst = 32'h10c00000;
      122005: inst = 32'hcc06b50;
      122006: inst = 32'h2080000b;
      122007: inst = 32'h10c00000;
      122008: inst = 32'hcc0eeb6;
      122009: inst = 32'h2080000c;
      122010: inst = 32'h10c00000;
      122011: inst = 32'hcc06b50;
      122012: inst = 32'h2080000d;
      122013: inst = 32'h10c00000;
      122014: inst = 32'hcc06b50;
      122015: inst = 32'h2080000e;
      122016: inst = 32'h10c00000;
      122017: inst = 32'hcc06b50;
      122018: inst = 32'h2080000f;
      122019: inst = 32'h10c00000;
      122020: inst = 32'hcc06b50;
      122021: inst = 32'h20800010;
      122022: inst = 32'h10c00000;
      122023: inst = 32'hcc06b50;
      122024: inst = 32'h20800011;
      122025: inst = 32'h10c00000;
      122026: inst = 32'hcc06b50;
      122027: inst = 32'h20800000;
      122028: inst = 32'h10c00000;
      122029: inst = 32'hcc06b50;
      122030: inst = 32'h20800001;
      122031: inst = 32'h10c00000;
      122032: inst = 32'hcc06b50;
      122033: inst = 32'h20800002;
      122034: inst = 32'h10c00000;
      122035: inst = 32'hcc06b50;
      122036: inst = 32'h20800003;
      122037: inst = 32'h10c00000;
      122038: inst = 32'hcc06b50;
      122039: inst = 32'h20800004;
      122040: inst = 32'h10c00000;
      122041: inst = 32'hcc06b50;
      122042: inst = 32'h20800005;
      122043: inst = 32'h10c00000;
      122044: inst = 32'hcc06b50;
      122045: inst = 32'h20800006;
      122046: inst = 32'h10c00000;
      122047: inst = 32'hcc0eeb6;
      122048: inst = 32'h20800007;
      122049: inst = 32'h10c00000;
      122050: inst = 32'hcc06b50;
      122051: inst = 32'h20800008;
      122052: inst = 32'h10c00000;
      122053: inst = 32'hcc0eeb6;
      122054: inst = 32'h20800009;
      122055: inst = 32'h10c00000;
      122056: inst = 32'hcc0eeb6;
      122057: inst = 32'h2080000a;
      122058: inst = 32'h10c00000;
      122059: inst = 32'hcc06b50;
      122060: inst = 32'h2080000b;
      122061: inst = 32'h10c00000;
      122062: inst = 32'hcc0eeb6;
      122063: inst = 32'h2080000c;
      122064: inst = 32'h10c00000;
      122065: inst = 32'hcc06b50;
      122066: inst = 32'h2080000d;
      122067: inst = 32'h10c00000;
      122068: inst = 32'hcc06b50;
      122069: inst = 32'h2080000e;
      122070: inst = 32'h10c00000;
      122071: inst = 32'hcc06b50;
      122072: inst = 32'h2080000f;
      122073: inst = 32'h10c00000;
      122074: inst = 32'hcc06b50;
      122075: inst = 32'h20800010;
      122076: inst = 32'h10c00000;
      122077: inst = 32'hcc06b50;
      122078: inst = 32'h20800011;
      122079: inst = 32'h10c00000;
      122080: inst = 32'hcc06b50;
      122081: inst = 32'h20800000;
      122082: inst = 32'h10c00000;
      122083: inst = 32'hcc06b50;
      122084: inst = 32'h20800001;
      122085: inst = 32'h10c00000;
      122086: inst = 32'hcc06b50;
      122087: inst = 32'h20800002;
      122088: inst = 32'h10c00000;
      122089: inst = 32'hcc06b50;
      122090: inst = 32'h20800003;
      122091: inst = 32'h10c00000;
      122092: inst = 32'hcc06b50;
      122093: inst = 32'h20800004;
      122094: inst = 32'h10c00000;
      122095: inst = 32'hcc06b50;
      122096: inst = 32'h20800005;
      122097: inst = 32'h10c00000;
      122098: inst = 32'hcc0eeb6;
      122099: inst = 32'h20800006;
      122100: inst = 32'h10c00000;
      122101: inst = 32'hcc0eeb6;
      122102: inst = 32'h20800007;
      122103: inst = 32'h10c00000;
      122104: inst = 32'hcc06b50;
      122105: inst = 32'h20800008;
      122106: inst = 32'h10c00000;
      122107: inst = 32'hcc0eeb6;
      122108: inst = 32'h20800009;
      122109: inst = 32'h10c00000;
      122110: inst = 32'hcc0eeb6;
      122111: inst = 32'h2080000a;
      122112: inst = 32'h10c00000;
      122113: inst = 32'hcc0eeb6;
      122114: inst = 32'h2080000b;
      122115: inst = 32'h10c00000;
      122116: inst = 32'hcc0eeb6;
      122117: inst = 32'h2080000c;
      122118: inst = 32'h10c00000;
      122119: inst = 32'hcc06b50;
      122120: inst = 32'h2080000d;
      122121: inst = 32'h10c00000;
      122122: inst = 32'hcc06b50;
      122123: inst = 32'h2080000e;
      122124: inst = 32'h10c00000;
      122125: inst = 32'hcc06b50;
      122126: inst = 32'h2080000f;
      122127: inst = 32'h10c00000;
      122128: inst = 32'hcc06b50;
      122129: inst = 32'h20800010;
      122130: inst = 32'h10c00000;
      122131: inst = 32'hcc06b50;
      122132: inst = 32'h20800011;
      122133: inst = 32'h10c00000;
      122134: inst = 32'hcc06b50;
      122135: inst = 32'h20800000;
      122136: inst = 32'h10c00000;
      122137: inst = 32'hcc06b50;
      122138: inst = 32'h20800001;
      122139: inst = 32'h10c00000;
      122140: inst = 32'hcc06b50;
      122141: inst = 32'h20800002;
      122142: inst = 32'h10c00000;
      122143: inst = 32'hcc06b50;
      122144: inst = 32'h20800003;
      122145: inst = 32'h10c00000;
      122146: inst = 32'hcc06b50;
      122147: inst = 32'h20800004;
      122148: inst = 32'h10c00000;
      122149: inst = 32'hcc06b50;
      122150: inst = 32'h20800005;
      122151: inst = 32'h10c00000;
      122152: inst = 32'hcc0eeb6;
      122153: inst = 32'h20800006;
      122154: inst = 32'h10c00000;
      122155: inst = 32'hcc0eeb6;
      122156: inst = 32'h20800007;
      122157: inst = 32'h10c00000;
      122158: inst = 32'hcc0eeb6;
      122159: inst = 32'h20800008;
      122160: inst = 32'h10c00000;
      122161: inst = 32'hcc0eeb6;
      122162: inst = 32'h20800009;
      122163: inst = 32'h10c00000;
      122164: inst = 32'hcc0eeb6;
      122165: inst = 32'h2080000a;
      122166: inst = 32'h10c00000;
      122167: inst = 32'hcc0eeb6;
      122168: inst = 32'h2080000b;
      122169: inst = 32'h10c00000;
      122170: inst = 32'hcc06b50;
      122171: inst = 32'h2080000c;
      122172: inst = 32'h10c00000;
      122173: inst = 32'hcc06b50;
      122174: inst = 32'h2080000d;
      122175: inst = 32'h10c00000;
      122176: inst = 32'hcc06b50;
      122177: inst = 32'h2080000e;
      122178: inst = 32'h10c00000;
      122179: inst = 32'hcc06b50;
      122180: inst = 32'h2080000f;
      122181: inst = 32'h10c00000;
      122182: inst = 32'hcc06b50;
      122183: inst = 32'h20800010;
      122184: inst = 32'h10c00000;
      122185: inst = 32'hcc06b50;
      122186: inst = 32'h20800011;
      122187: inst = 32'h10c00000;
      122188: inst = 32'hcc06b50;
      122189: inst = 32'h20800000;
      122190: inst = 32'h10c00000;
      122191: inst = 32'hcc06b50;
      122192: inst = 32'h20800001;
      122193: inst = 32'h10c00000;
      122194: inst = 32'hcc06b50;
      122195: inst = 32'h20800002;
      122196: inst = 32'h10c00000;
      122197: inst = 32'hcc06b50;
      122198: inst = 32'h20800003;
      122199: inst = 32'h10c00000;
      122200: inst = 32'hcc06b50;
      122201: inst = 32'h20800004;
      122202: inst = 32'h10c00000;
      122203: inst = 32'hcc06b50;
      122204: inst = 32'h20800005;
      122205: inst = 32'h10c00000;
      122206: inst = 32'hcc0eeb6;
      122207: inst = 32'h20800006;
      122208: inst = 32'h10c00000;
      122209: inst = 32'hcc0eeb6;
      122210: inst = 32'h20800007;
      122211: inst = 32'h10c00000;
      122212: inst = 32'hcc06b50;
      122213: inst = 32'h20800008;
      122214: inst = 32'h10c00000;
      122215: inst = 32'hcc0eeb6;
      122216: inst = 32'h20800009;
      122217: inst = 32'h10c00000;
      122218: inst = 32'hcc0eeb6;
      122219: inst = 32'h2080000a;
      122220: inst = 32'h10c00000;
      122221: inst = 32'hcc0eeb6;
      122222: inst = 32'h2080000b;
      122223: inst = 32'h10c00000;
      122224: inst = 32'hcc06b50;
      122225: inst = 32'h2080000c;
      122226: inst = 32'h10c00000;
      122227: inst = 32'hcc06b50;
      122228: inst = 32'h2080000d;
      122229: inst = 32'h10c00000;
      122230: inst = 32'hcc06b50;
      122231: inst = 32'h2080000e;
      122232: inst = 32'h10c00000;
      122233: inst = 32'hcc06b50;
      122234: inst = 32'h2080000f;
      122235: inst = 32'h10c00000;
      122236: inst = 32'hcc06b50;
      122237: inst = 32'h20800010;
      122238: inst = 32'h10c00000;
      122239: inst = 32'hcc06b50;
      122240: inst = 32'h20800011;
      122241: inst = 32'h10c00000;
      122242: inst = 32'hcc06b50;
      122243: inst = 32'h20800000;
      122244: inst = 32'h10c00000;
      122245: inst = 32'hcc06b50;
      122246: inst = 32'h20800001;
      122247: inst = 32'h10c00000;
      122248: inst = 32'hcc06b50;
      122249: inst = 32'h20800002;
      122250: inst = 32'h10c00000;
      122251: inst = 32'hcc06b50;
      122252: inst = 32'h20800003;
      122253: inst = 32'h10c00000;
      122254: inst = 32'hcc06b50;
      122255: inst = 32'h20800004;
      122256: inst = 32'h10c00000;
      122257: inst = 32'hcc06b50;
      122258: inst = 32'h20800005;
      122259: inst = 32'h10c00000;
      122260: inst = 32'hcc0eeb6;
      122261: inst = 32'h20800006;
      122262: inst = 32'h10c00000;
      122263: inst = 32'hcc0eeb6;
      122264: inst = 32'h20800007;
      122265: inst = 32'h10c00000;
      122266: inst = 32'hcc06b50;
      122267: inst = 32'h20800008;
      122268: inst = 32'h10c00000;
      122269: inst = 32'hcc0eeb6;
      122270: inst = 32'h20800009;
      122271: inst = 32'h10c00000;
      122272: inst = 32'hcc0eeb6;
      122273: inst = 32'h2080000a;
      122274: inst = 32'h10c00000;
      122275: inst = 32'hcc0eeb6;
      122276: inst = 32'h2080000b;
      122277: inst = 32'h10c00000;
      122278: inst = 32'hcc06b50;
      122279: inst = 32'h2080000c;
      122280: inst = 32'h10c00000;
      122281: inst = 32'hcc06b50;
      122282: inst = 32'h2080000d;
      122283: inst = 32'h10c00000;
      122284: inst = 32'hcc06b50;
      122285: inst = 32'h2080000e;
      122286: inst = 32'h10c00000;
      122287: inst = 32'hcc06b50;
      122288: inst = 32'h2080000f;
      122289: inst = 32'h10c00000;
      122290: inst = 32'hcc06b50;
      122291: inst = 32'h20800010;
      122292: inst = 32'h10c00000;
      122293: inst = 32'hcc06b50;
      122294: inst = 32'h20800011;
      122295: inst = 32'h10c00000;
      122296: inst = 32'hcc06b50;
      122297: inst = 32'h20800000;
      122298: inst = 32'h10c00000;
      122299: inst = 32'hcc06b50;
      122300: inst = 32'h20800001;
      122301: inst = 32'h10c00000;
      122302: inst = 32'hcc06b50;
      122303: inst = 32'h20800002;
      122304: inst = 32'h10c00000;
      122305: inst = 32'hcc06b50;
      122306: inst = 32'h20800003;
      122307: inst = 32'h10c00000;
      122308: inst = 32'hcc06b50;
      122309: inst = 32'h20800004;
      122310: inst = 32'h10c00000;
      122311: inst = 32'hcc06b50;
      122312: inst = 32'h20800005;
      122313: inst = 32'h10c00000;
      122314: inst = 32'hcc0eeb6;
      122315: inst = 32'h20800006;
      122316: inst = 32'h10c00000;
      122317: inst = 32'hcc0eeb6;
      122318: inst = 32'h20800007;
      122319: inst = 32'h10c00000;
      122320: inst = 32'hcc06b50;
      122321: inst = 32'h20800008;
      122322: inst = 32'h10c00000;
      122323: inst = 32'hcc0eeb6;
      122324: inst = 32'h20800009;
      122325: inst = 32'h10c00000;
      122326: inst = 32'hcc0eeb6;
      122327: inst = 32'h2080000a;
      122328: inst = 32'h10c00000;
      122329: inst = 32'hcc0eeb6;
      122330: inst = 32'h2080000b;
      122331: inst = 32'h10c00000;
      122332: inst = 32'hcc06b50;
      122333: inst = 32'h2080000c;
      122334: inst = 32'h10c00000;
      122335: inst = 32'hcc06b50;
      122336: inst = 32'h2080000d;
      122337: inst = 32'h10c00000;
      122338: inst = 32'hcc06b50;
      122339: inst = 32'h2080000e;
      122340: inst = 32'h10c00000;
      122341: inst = 32'hcc06b50;
      122342: inst = 32'h2080000f;
      122343: inst = 32'h10c00000;
      122344: inst = 32'hcc06b50;
      122345: inst = 32'h20800010;
      122346: inst = 32'h10c00000;
      122347: inst = 32'hcc06b50;
      122348: inst = 32'h20800011;
      122349: inst = 32'h10c00000;
      122350: inst = 32'hcc06b50;
      122351: inst = 32'h20800000;
      122352: inst = 32'h10c00000;
      122353: inst = 32'hcc06b50;
      122354: inst = 32'h20800001;
      122355: inst = 32'h10c00000;
      122356: inst = 32'hcc06b50;
      122357: inst = 32'h20800002;
      122358: inst = 32'h10c00000;
      122359: inst = 32'hcc06b50;
      122360: inst = 32'h20800003;
      122361: inst = 32'h10c00000;
      122362: inst = 32'hcc06b50;
      122363: inst = 32'h20800004;
      122364: inst = 32'h10c00000;
      122365: inst = 32'hcc06b50;
      122366: inst = 32'h20800005;
      122367: inst = 32'h10c00000;
      122368: inst = 32'hcc0eeb6;
      122369: inst = 32'h20800006;
      122370: inst = 32'h10c00000;
      122371: inst = 32'hcc0eeb6;
      122372: inst = 32'h20800007;
      122373: inst = 32'h10c00000;
      122374: inst = 32'hcc06b50;
      122375: inst = 32'h20800008;
      122376: inst = 32'h10c00000;
      122377: inst = 32'hcc0eeb6;
      122378: inst = 32'h20800009;
      122379: inst = 32'h10c00000;
      122380: inst = 32'hcc0eeb6;
      122381: inst = 32'h2080000a;
      122382: inst = 32'h10c00000;
      122383: inst = 32'hcc0eeb6;
      122384: inst = 32'h2080000b;
      122385: inst = 32'h10c00000;
      122386: inst = 32'hcc06b50;
      122387: inst = 32'h2080000c;
      122388: inst = 32'h10c00000;
      122389: inst = 32'hcc06b50;
      122390: inst = 32'h2080000d;
      122391: inst = 32'h10c00000;
      122392: inst = 32'hcc06b50;
      122393: inst = 32'h2080000e;
      122394: inst = 32'h10c00000;
      122395: inst = 32'hcc06b50;
      122396: inst = 32'h2080000f;
      122397: inst = 32'h10c00000;
      122398: inst = 32'hcc06b50;
      122399: inst = 32'h20800010;
      122400: inst = 32'h10c00000;
      122401: inst = 32'hcc06b50;
      122402: inst = 32'h20800011;
      122403: inst = 32'h10c00000;
      122404: inst = 32'hcc06b50;
      122405: inst = 32'h20800000;
      122406: inst = 32'h10c00000;
      122407: inst = 32'hcc06b50;
      122408: inst = 32'h20800001;
      122409: inst = 32'h10c00000;
      122410: inst = 32'hcc06b50;
      122411: inst = 32'h20800002;
      122412: inst = 32'h10c00000;
      122413: inst = 32'hcc06b50;
      122414: inst = 32'h20800003;
      122415: inst = 32'h10c00000;
      122416: inst = 32'hcc06b50;
      122417: inst = 32'h20800004;
      122418: inst = 32'h10c00000;
      122419: inst = 32'hcc06b50;
      122420: inst = 32'h20800005;
      122421: inst = 32'h10c00000;
      122422: inst = 32'hcc06b50;
      122423: inst = 32'h20800006;
      122424: inst = 32'h10c00000;
      122425: inst = 32'hcc06b50;
      122426: inst = 32'h20800007;
      122427: inst = 32'h10c00000;
      122428: inst = 32'hcc06b50;
      122429: inst = 32'h20800008;
      122430: inst = 32'h10c00000;
      122431: inst = 32'hcc06b50;
      122432: inst = 32'h20800009;
      122433: inst = 32'h10c00000;
      122434: inst = 32'hcc06b50;
      122435: inst = 32'h2080000a;
      122436: inst = 32'h10c00000;
      122437: inst = 32'hcc06b50;
      122438: inst = 32'h2080000b;
      122439: inst = 32'h10c00000;
      122440: inst = 32'hcc06b50;
      122441: inst = 32'h2080000c;
      122442: inst = 32'h10c00000;
      122443: inst = 32'hcc06b50;
      122444: inst = 32'h2080000d;
      122445: inst = 32'h10c00000;
      122446: inst = 32'hcc06b50;
      122447: inst = 32'h2080000e;
      122448: inst = 32'h10c00000;
      122449: inst = 32'hcc06b50;
      122450: inst = 32'h2080000f;
      122451: inst = 32'h10c00000;
      122452: inst = 32'hcc06b50;
      122453: inst = 32'h20800010;
      122454: inst = 32'h10c00000;
      122455: inst = 32'hcc06b50;
      122456: inst = 32'h20800011;
      122457: inst = 32'h10c00000;
      122458: inst = 32'hcc06b50;
      122459: inst = 32'h20800000;
      122460: inst = 32'h10c00000;
      122461: inst = 32'hcc06b50;
      122462: inst = 32'h20800001;
      122463: inst = 32'h10c00000;
      122464: inst = 32'hcc06b50;
      122465: inst = 32'h20800002;
      122466: inst = 32'h10c00000;
      122467: inst = 32'hcc06b50;
      122468: inst = 32'h20800003;
      122469: inst = 32'h10c00000;
      122470: inst = 32'hcc06b50;
      122471: inst = 32'h20800004;
      122472: inst = 32'h10c00000;
      122473: inst = 32'hcc06b50;
      122474: inst = 32'h20800005;
      122475: inst = 32'h10c00000;
      122476: inst = 32'hcc06b50;
      122477: inst = 32'h20800006;
      122478: inst = 32'h10c00000;
      122479: inst = 32'hcc06b50;
      122480: inst = 32'h20800007;
      122481: inst = 32'h10c00000;
      122482: inst = 32'hcc06b50;
      122483: inst = 32'h20800008;
      122484: inst = 32'h10c00000;
      122485: inst = 32'hcc06b50;
      122486: inst = 32'h20800009;
      122487: inst = 32'h10c00000;
      122488: inst = 32'hcc06b50;
      122489: inst = 32'h2080000a;
      122490: inst = 32'h10c00000;
      122491: inst = 32'hcc06b50;
      122492: inst = 32'h2080000b;
      122493: inst = 32'h10c00000;
      122494: inst = 32'hcc06b50;
      122495: inst = 32'h2080000c;
      122496: inst = 32'h10c00000;
      122497: inst = 32'hcc06b50;
      122498: inst = 32'h2080000d;
      122499: inst = 32'h10c00000;
      122500: inst = 32'hcc06b50;
      122501: inst = 32'h2080000e;
      122502: inst = 32'h10c00000;
      122503: inst = 32'hcc06b50;
      122504: inst = 32'h2080000f;
      122505: inst = 32'h10c00000;
      122506: inst = 32'hcc06b50;
      122507: inst = 32'h20800010;
      122508: inst = 32'h10c00000;
      122509: inst = 32'hcc06b50;
      122510: inst = 32'h20800011;
      122511: inst = 32'h10c00000;
      122512: inst = 32'hcc06b50;
      122513: inst = 32'h20800000;
      122514: inst = 32'h10c00000;
      122515: inst = 32'hcc06b50;
      122516: inst = 32'h20800001;
      122517: inst = 32'h10c00000;
      122518: inst = 32'hcc06b50;
      122519: inst = 32'h20800002;
      122520: inst = 32'h10c00000;
      122521: inst = 32'hcc06b50;
      122522: inst = 32'h20800003;
      122523: inst = 32'h10c00000;
      122524: inst = 32'hcc06b50;
      122525: inst = 32'h20800004;
      122526: inst = 32'h10c00000;
      122527: inst = 32'hcc06b50;
      122528: inst = 32'h20800005;
      122529: inst = 32'h10c00000;
      122530: inst = 32'hcc06b50;
      122531: inst = 32'h20800006;
      122532: inst = 32'h10c00000;
      122533: inst = 32'hcc06b50;
      122534: inst = 32'h20800007;
      122535: inst = 32'h10c00000;
      122536: inst = 32'hcc06b50;
      122537: inst = 32'h20800008;
      122538: inst = 32'h10c00000;
      122539: inst = 32'hcc06b50;
      122540: inst = 32'h20800009;
      122541: inst = 32'h10c00000;
      122542: inst = 32'hcc06b50;
      122543: inst = 32'h2080000a;
      122544: inst = 32'h10c00000;
      122545: inst = 32'hcc06b50;
      122546: inst = 32'h2080000b;
      122547: inst = 32'h10c00000;
      122548: inst = 32'hcc06b50;
      122549: inst = 32'h2080000c;
      122550: inst = 32'h10c00000;
      122551: inst = 32'hcc06b50;
      122552: inst = 32'h2080000d;
      122553: inst = 32'h10c00000;
      122554: inst = 32'hcc06b50;
      122555: inst = 32'h2080000e;
      122556: inst = 32'h10c00000;
      122557: inst = 32'hcc06b50;
      122558: inst = 32'h2080000f;
      122559: inst = 32'h10c00000;
      122560: inst = 32'hcc06b50;
      122561: inst = 32'h20800010;
      122562: inst = 32'h10c00000;
      122563: inst = 32'hcc06b50;
      122564: inst = 32'h20800011;
      122565: inst = 32'h10c00000;
      122566: inst = 32'hcc06b50;
      122567: inst = 32'h20800000;
      122568: inst = 32'h10c00000;
      122569: inst = 32'hcc06b50;
      122570: inst = 32'h20800001;
      122571: inst = 32'h10c00000;
      122572: inst = 32'hcc06b50;
      122573: inst = 32'h20800002;
      122574: inst = 32'h10c00000;
      122575: inst = 32'hcc06b50;
      122576: inst = 32'h20800003;
      122577: inst = 32'h10c00000;
      122578: inst = 32'hcc06b50;
      122579: inst = 32'h20800004;
      122580: inst = 32'h10c00000;
      122581: inst = 32'hcc06b50;
      122582: inst = 32'h20800005;
      122583: inst = 32'h10c00000;
      122584: inst = 32'hcc06b50;
      122585: inst = 32'h20800006;
      122586: inst = 32'h10c00000;
      122587: inst = 32'hcc06b50;
      122588: inst = 32'h20800007;
      122589: inst = 32'h10c00000;
      122590: inst = 32'hcc06b50;
      122591: inst = 32'h20800008;
      122592: inst = 32'h10c00000;
      122593: inst = 32'hcc06b50;
      122594: inst = 32'h20800009;
      122595: inst = 32'h10c00000;
      122596: inst = 32'hcc06b50;
      122597: inst = 32'h2080000a;
      122598: inst = 32'h10c00000;
      122599: inst = 32'hcc06b50;
      122600: inst = 32'h2080000b;
      122601: inst = 32'h10c00000;
      122602: inst = 32'hcc06b50;
      122603: inst = 32'h2080000c;
      122604: inst = 32'h10c00000;
      122605: inst = 32'hcc06b50;
      122606: inst = 32'h2080000d;
      122607: inst = 32'h10c00000;
      122608: inst = 32'hcc06b50;
      122609: inst = 32'h2080000e;
      122610: inst = 32'h10c00000;
      122611: inst = 32'hcc06b50;
      122612: inst = 32'h2080000f;
      122613: inst = 32'h10c00000;
      122614: inst = 32'hcc06b50;
      122615: inst = 32'h20800010;
      122616: inst = 32'h10c00000;
      122617: inst = 32'hcc06b50;
      122618: inst = 32'h20800011;
      122619: inst = 32'h10c00000;
      122620: inst = 32'hcc06b50;
      122621: inst = 32'h58a00000;
    endcase
  end
endmodule
