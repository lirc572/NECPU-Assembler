`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: lirc572
// Engineer: lirc572
// 
// Create Date: 
// Design Name: NECPU
// Module Name: InstMem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module instMem (
    input  [31:0]  address,
    output reg [31:0] inst
  );
  always @ (address) begin
    inst = 32'd0;
    case (address)
      0: inst = 32'h10000000;
      1: inst = 32'hc000005;
      2: inst = 32'h13e00000;
      3: inst = 32'hfe0004c;
      4: inst = 32'h5be00000;
      5: inst = 32'h13c0007f;
      6: inst = 32'hfc02815;
      7: inst = 32'h33de0001;
      8: inst = 32'h13e00000;
      9: inst = 32'hfe00007;
      10: inst = 32'h1fc00000;
      11: inst = 32'h5be00000;
      12: inst = 32'h10000000;
      13: inst = 32'hc000011;
      14: inst = 32'h13e00000;
      15: inst = 32'hfe048a4;
      16: inst = 32'h5be00000;
      17: inst = 32'h13c0007f;
      18: inst = 32'hfc02815;
      19: inst = 32'h33de0001;
      20: inst = 32'h13e00000;
      21: inst = 32'hfe00013;
      22: inst = 32'h1fc00000;
      23: inst = 32'h5be00000;
      24: inst = 32'h10000000;
      25: inst = 32'hc000000;
      26: inst = 32'h10200000;
      27: inst = 32'hc20001f;
      28: inst = 32'h13e00000;
      29: inst = 32'hfe065ff;
      30: inst = 32'h5be00000;
      31: inst = 32'h10000000;
      32: inst = 32'hc000024;
      33: inst = 32'h13e00000;
      34: inst = 32'hfe050f5;
      35: inst = 32'h5be00000;
      36: inst = 32'h13c001fc;
      37: inst = 32'hfc0a055;
      38: inst = 32'h33de0001;
      39: inst = 32'h13e00000;
      40: inst = 32'hfe00026;
      41: inst = 32'h1fc00000;
      42: inst = 32'h5be00000;
      43: inst = 32'h10000000;
      44: inst = 32'hc00002b;
      45: inst = 32'h10200000;
      46: inst = 32'hc200032;
      47: inst = 32'h13e00000;
      48: inst = 32'hfe065ff;
      49: inst = 32'h5be00000;
      50: inst = 32'h10200000;
      51: inst = 32'hc200000;
      52: inst = 32'h10000000;
      53: inst = 32'hc000039;
      54: inst = 32'h13e00000;
      55: inst = 32'hfe06369;
      56: inst = 32'h5be00000;
      57: inst = 32'h13e00000;
      58: inst = 32'hfe0003c;
      59: inst = 32'h5be00000;
      60: inst = 32'h10608000;
      61: inst = 32'hc600000;
      62: inst = 32'h10200000;
      63: inst = 32'hc20aaaa;
      64: inst = 32'h4c210000;
      65: inst = 32'h8230000;
      66: inst = 32'h104000fe;
      67: inst = 32'hc40502a;
      68: inst = 32'h30420001;
      69: inst = 32'h13e00000;
      70: inst = 32'hfe00044;
      71: inst = 32'h1c400000;
      72: inst = 32'h5be00000;
      73: inst = 32'h13e00000;
      74: inst = 32'hfe00040;
      75: inst = 32'h5be00000;
      76: inst = 32'hc20eeb6;
      77: inst = 32'h10408000;
      78: inst = 32'hc403fe0;
      79: inst = 32'h8220000;
      80: inst = 32'h10408000;
      81: inst = 32'hc403fe1;
      82: inst = 32'h8220000;
      83: inst = 32'h10408000;
      84: inst = 32'hc403fe2;
      85: inst = 32'h8220000;
      86: inst = 32'h10408000;
      87: inst = 32'hc403fe3;
      88: inst = 32'h8220000;
      89: inst = 32'h10408000;
      90: inst = 32'hc403fe4;
      91: inst = 32'h8220000;
      92: inst = 32'h10408000;
      93: inst = 32'hc403fe5;
      94: inst = 32'h8220000;
      95: inst = 32'h10408000;
      96: inst = 32'hc403fe6;
      97: inst = 32'h8220000;
      98: inst = 32'h10408000;
      99: inst = 32'hc403fe7;
      100: inst = 32'h8220000;
      101: inst = 32'h10408000;
      102: inst = 32'hc403fe8;
      103: inst = 32'h8220000;
      104: inst = 32'h10408000;
      105: inst = 32'hc403fe9;
      106: inst = 32'h8220000;
      107: inst = 32'h10408000;
      108: inst = 32'hc403fea;
      109: inst = 32'h8220000;
      110: inst = 32'h10408000;
      111: inst = 32'hc403fec;
      112: inst = 32'h8220000;
      113: inst = 32'h10408000;
      114: inst = 32'hc403fed;
      115: inst = 32'h8220000;
      116: inst = 32'h10408000;
      117: inst = 32'hc403fee;
      118: inst = 32'h8220000;
      119: inst = 32'h10408000;
      120: inst = 32'hc403fef;
      121: inst = 32'h8220000;
      122: inst = 32'h10408000;
      123: inst = 32'hc403ff0;
      124: inst = 32'h8220000;
      125: inst = 32'h10408000;
      126: inst = 32'hc403ff1;
      127: inst = 32'h8220000;
      128: inst = 32'h10408000;
      129: inst = 32'hc403ff2;
      130: inst = 32'h8220000;
      131: inst = 32'h10408000;
      132: inst = 32'hc403ff3;
      133: inst = 32'h8220000;
      134: inst = 32'h10408000;
      135: inst = 32'hc403ff4;
      136: inst = 32'h8220000;
      137: inst = 32'h10408000;
      138: inst = 32'hc403ff5;
      139: inst = 32'h8220000;
      140: inst = 32'h10408000;
      141: inst = 32'hc403ff6;
      142: inst = 32'h8220000;
      143: inst = 32'h10408000;
      144: inst = 32'hc403ff7;
      145: inst = 32'h8220000;
      146: inst = 32'h10408000;
      147: inst = 32'hc403ff8;
      148: inst = 32'h8220000;
      149: inst = 32'h10408000;
      150: inst = 32'hc403ff9;
      151: inst = 32'h8220000;
      152: inst = 32'h10408000;
      153: inst = 32'hc403ffa;
      154: inst = 32'h8220000;
      155: inst = 32'h10408000;
      156: inst = 32'hc403ffb;
      157: inst = 32'h8220000;
      158: inst = 32'h10408000;
      159: inst = 32'hc403ffc;
      160: inst = 32'h8220000;
      161: inst = 32'h10408000;
      162: inst = 32'hc403ffd;
      163: inst = 32'h8220000;
      164: inst = 32'h10408000;
      165: inst = 32'hc403ffe;
      166: inst = 32'h8220000;
      167: inst = 32'h10408000;
      168: inst = 32'hc403fff;
      169: inst = 32'h8220000;
      170: inst = 32'h10408000;
      171: inst = 32'hc404000;
      172: inst = 32'h8220000;
      173: inst = 32'h10408000;
      174: inst = 32'hc404001;
      175: inst = 32'h8220000;
      176: inst = 32'h10408000;
      177: inst = 32'hc404002;
      178: inst = 32'h8220000;
      179: inst = 32'h10408000;
      180: inst = 32'hc404003;
      181: inst = 32'h8220000;
      182: inst = 32'h10408000;
      183: inst = 32'hc404004;
      184: inst = 32'h8220000;
      185: inst = 32'h10408000;
      186: inst = 32'hc404005;
      187: inst = 32'h8220000;
      188: inst = 32'h10408000;
      189: inst = 32'hc404006;
      190: inst = 32'h8220000;
      191: inst = 32'h10408000;
      192: inst = 32'hc404007;
      193: inst = 32'h8220000;
      194: inst = 32'h10408000;
      195: inst = 32'hc404008;
      196: inst = 32'h8220000;
      197: inst = 32'h10408000;
      198: inst = 32'hc404009;
      199: inst = 32'h8220000;
      200: inst = 32'h10408000;
      201: inst = 32'hc40400a;
      202: inst = 32'h8220000;
      203: inst = 32'h10408000;
      204: inst = 32'hc40400b;
      205: inst = 32'h8220000;
      206: inst = 32'h10408000;
      207: inst = 32'hc40400c;
      208: inst = 32'h8220000;
      209: inst = 32'h10408000;
      210: inst = 32'hc40400d;
      211: inst = 32'h8220000;
      212: inst = 32'h10408000;
      213: inst = 32'hc40400e;
      214: inst = 32'h8220000;
      215: inst = 32'h10408000;
      216: inst = 32'hc40400f;
      217: inst = 32'h8220000;
      218: inst = 32'h10408000;
      219: inst = 32'hc404010;
      220: inst = 32'h8220000;
      221: inst = 32'h10408000;
      222: inst = 32'hc404011;
      223: inst = 32'h8220000;
      224: inst = 32'h10408000;
      225: inst = 32'hc404012;
      226: inst = 32'h8220000;
      227: inst = 32'h10408000;
      228: inst = 32'hc404013;
      229: inst = 32'h8220000;
      230: inst = 32'h10408000;
      231: inst = 32'hc404014;
      232: inst = 32'h8220000;
      233: inst = 32'h10408000;
      234: inst = 32'hc404015;
      235: inst = 32'h8220000;
      236: inst = 32'h10408000;
      237: inst = 32'hc404016;
      238: inst = 32'h8220000;
      239: inst = 32'h10408000;
      240: inst = 32'hc404017;
      241: inst = 32'h8220000;
      242: inst = 32'h10408000;
      243: inst = 32'hc404018;
      244: inst = 32'h8220000;
      245: inst = 32'h10408000;
      246: inst = 32'hc404019;
      247: inst = 32'h8220000;
      248: inst = 32'h10408000;
      249: inst = 32'hc40401a;
      250: inst = 32'h8220000;
      251: inst = 32'h10408000;
      252: inst = 32'hc40401b;
      253: inst = 32'h8220000;
      254: inst = 32'h10408000;
      255: inst = 32'hc40401c;
      256: inst = 32'h8220000;
      257: inst = 32'h10408000;
      258: inst = 32'hc40401d;
      259: inst = 32'h8220000;
      260: inst = 32'h10408000;
      261: inst = 32'hc40401e;
      262: inst = 32'h8220000;
      263: inst = 32'h10408000;
      264: inst = 32'hc40401f;
      265: inst = 32'h8220000;
      266: inst = 32'h10408000;
      267: inst = 32'hc404020;
      268: inst = 32'h8220000;
      269: inst = 32'h10408000;
      270: inst = 32'hc404021;
      271: inst = 32'h8220000;
      272: inst = 32'h10408000;
      273: inst = 32'hc404022;
      274: inst = 32'h8220000;
      275: inst = 32'h10408000;
      276: inst = 32'hc404023;
      277: inst = 32'h8220000;
      278: inst = 32'h10408000;
      279: inst = 32'hc404024;
      280: inst = 32'h8220000;
      281: inst = 32'h10408000;
      282: inst = 32'hc404025;
      283: inst = 32'h8220000;
      284: inst = 32'h10408000;
      285: inst = 32'hc404026;
      286: inst = 32'h8220000;
      287: inst = 32'h10408000;
      288: inst = 32'hc404027;
      289: inst = 32'h8220000;
      290: inst = 32'h10408000;
      291: inst = 32'hc404028;
      292: inst = 32'h8220000;
      293: inst = 32'h10408000;
      294: inst = 32'hc404029;
      295: inst = 32'h8220000;
      296: inst = 32'h10408000;
      297: inst = 32'hc40402a;
      298: inst = 32'h8220000;
      299: inst = 32'h10408000;
      300: inst = 32'hc40402b;
      301: inst = 32'h8220000;
      302: inst = 32'h10408000;
      303: inst = 32'hc40402c;
      304: inst = 32'h8220000;
      305: inst = 32'h10408000;
      306: inst = 32'hc40402d;
      307: inst = 32'h8220000;
      308: inst = 32'h10408000;
      309: inst = 32'hc40402e;
      310: inst = 32'h8220000;
      311: inst = 32'h10408000;
      312: inst = 32'hc40402f;
      313: inst = 32'h8220000;
      314: inst = 32'h10408000;
      315: inst = 32'hc404030;
      316: inst = 32'h8220000;
      317: inst = 32'h10408000;
      318: inst = 32'hc404031;
      319: inst = 32'h8220000;
      320: inst = 32'h10408000;
      321: inst = 32'hc404032;
      322: inst = 32'h8220000;
      323: inst = 32'h10408000;
      324: inst = 32'hc404033;
      325: inst = 32'h8220000;
      326: inst = 32'h10408000;
      327: inst = 32'hc404034;
      328: inst = 32'h8220000;
      329: inst = 32'h10408000;
      330: inst = 32'hc404035;
      331: inst = 32'h8220000;
      332: inst = 32'h10408000;
      333: inst = 32'hc404036;
      334: inst = 32'h8220000;
      335: inst = 32'h10408000;
      336: inst = 32'hc404037;
      337: inst = 32'h8220000;
      338: inst = 32'h10408000;
      339: inst = 32'hc404038;
      340: inst = 32'h8220000;
      341: inst = 32'h10408000;
      342: inst = 32'hc404039;
      343: inst = 32'h8220000;
      344: inst = 32'h10408000;
      345: inst = 32'hc40403a;
      346: inst = 32'h8220000;
      347: inst = 32'h10408000;
      348: inst = 32'hc40403b;
      349: inst = 32'h8220000;
      350: inst = 32'h10408000;
      351: inst = 32'hc40403c;
      352: inst = 32'h8220000;
      353: inst = 32'h10408000;
      354: inst = 32'hc40403d;
      355: inst = 32'h8220000;
      356: inst = 32'h10408000;
      357: inst = 32'hc40403e;
      358: inst = 32'h8220000;
      359: inst = 32'h10408000;
      360: inst = 32'hc40403f;
      361: inst = 32'h8220000;
      362: inst = 32'h10408000;
      363: inst = 32'hc404040;
      364: inst = 32'h8220000;
      365: inst = 32'h10408000;
      366: inst = 32'hc404041;
      367: inst = 32'h8220000;
      368: inst = 32'h10408000;
      369: inst = 32'hc404042;
      370: inst = 32'h8220000;
      371: inst = 32'h10408000;
      372: inst = 32'hc404043;
      373: inst = 32'h8220000;
      374: inst = 32'h10408000;
      375: inst = 32'hc404044;
      376: inst = 32'h8220000;
      377: inst = 32'h10408000;
      378: inst = 32'hc404045;
      379: inst = 32'h8220000;
      380: inst = 32'h10408000;
      381: inst = 32'hc404046;
      382: inst = 32'h8220000;
      383: inst = 32'h10408000;
      384: inst = 32'hc404047;
      385: inst = 32'h8220000;
      386: inst = 32'h10408000;
      387: inst = 32'hc404048;
      388: inst = 32'h8220000;
      389: inst = 32'h10408000;
      390: inst = 32'hc404049;
      391: inst = 32'h8220000;
      392: inst = 32'h10408000;
      393: inst = 32'hc40404a;
      394: inst = 32'h8220000;
      395: inst = 32'h10408000;
      396: inst = 32'hc40404c;
      397: inst = 32'h8220000;
      398: inst = 32'h10408000;
      399: inst = 32'hc40404d;
      400: inst = 32'h8220000;
      401: inst = 32'h10408000;
      402: inst = 32'hc40404e;
      403: inst = 32'h8220000;
      404: inst = 32'h10408000;
      405: inst = 32'hc40404f;
      406: inst = 32'h8220000;
      407: inst = 32'h10408000;
      408: inst = 32'hc404050;
      409: inst = 32'h8220000;
      410: inst = 32'h10408000;
      411: inst = 32'hc404051;
      412: inst = 32'h8220000;
      413: inst = 32'h10408000;
      414: inst = 32'hc404052;
      415: inst = 32'h8220000;
      416: inst = 32'h10408000;
      417: inst = 32'hc404053;
      418: inst = 32'h8220000;
      419: inst = 32'h10408000;
      420: inst = 32'hc404054;
      421: inst = 32'h8220000;
      422: inst = 32'h10408000;
      423: inst = 32'hc404055;
      424: inst = 32'h8220000;
      425: inst = 32'h10408000;
      426: inst = 32'hc404056;
      427: inst = 32'h8220000;
      428: inst = 32'h10408000;
      429: inst = 32'hc404057;
      430: inst = 32'h8220000;
      431: inst = 32'h10408000;
      432: inst = 32'hc404058;
      433: inst = 32'h8220000;
      434: inst = 32'h10408000;
      435: inst = 32'hc404059;
      436: inst = 32'h8220000;
      437: inst = 32'h10408000;
      438: inst = 32'hc40405a;
      439: inst = 32'h8220000;
      440: inst = 32'h10408000;
      441: inst = 32'hc40405b;
      442: inst = 32'h8220000;
      443: inst = 32'h10408000;
      444: inst = 32'hc40405c;
      445: inst = 32'h8220000;
      446: inst = 32'h10408000;
      447: inst = 32'hc40405d;
      448: inst = 32'h8220000;
      449: inst = 32'h10408000;
      450: inst = 32'hc40405e;
      451: inst = 32'h8220000;
      452: inst = 32'h10408000;
      453: inst = 32'hc40405f;
      454: inst = 32'h8220000;
      455: inst = 32'h10408000;
      456: inst = 32'hc404060;
      457: inst = 32'h8220000;
      458: inst = 32'h10408000;
      459: inst = 32'hc404061;
      460: inst = 32'h8220000;
      461: inst = 32'h10408000;
      462: inst = 32'hc404062;
      463: inst = 32'h8220000;
      464: inst = 32'h10408000;
      465: inst = 32'hc404063;
      466: inst = 32'h8220000;
      467: inst = 32'h10408000;
      468: inst = 32'hc404064;
      469: inst = 32'h8220000;
      470: inst = 32'h10408000;
      471: inst = 32'hc404065;
      472: inst = 32'h8220000;
      473: inst = 32'h10408000;
      474: inst = 32'hc404066;
      475: inst = 32'h8220000;
      476: inst = 32'h10408000;
      477: inst = 32'hc404067;
      478: inst = 32'h8220000;
      479: inst = 32'h10408000;
      480: inst = 32'hc404068;
      481: inst = 32'h8220000;
      482: inst = 32'h10408000;
      483: inst = 32'hc404069;
      484: inst = 32'h8220000;
      485: inst = 32'h10408000;
      486: inst = 32'hc40406a;
      487: inst = 32'h8220000;
      488: inst = 32'h10408000;
      489: inst = 32'hc40406b;
      490: inst = 32'h8220000;
      491: inst = 32'h10408000;
      492: inst = 32'hc40406c;
      493: inst = 32'h8220000;
      494: inst = 32'h10408000;
      495: inst = 32'hc40406d;
      496: inst = 32'h8220000;
      497: inst = 32'h10408000;
      498: inst = 32'hc40406e;
      499: inst = 32'h8220000;
      500: inst = 32'h10408000;
      501: inst = 32'hc40406f;
      502: inst = 32'h8220000;
      503: inst = 32'h10408000;
      504: inst = 32'hc404070;
      505: inst = 32'h8220000;
      506: inst = 32'h10408000;
      507: inst = 32'hc404071;
      508: inst = 32'h8220000;
      509: inst = 32'h10408000;
      510: inst = 32'hc404072;
      511: inst = 32'h8220000;
      512: inst = 32'h10408000;
      513: inst = 32'hc404073;
      514: inst = 32'h8220000;
      515: inst = 32'h10408000;
      516: inst = 32'hc404074;
      517: inst = 32'h8220000;
      518: inst = 32'h10408000;
      519: inst = 32'hc404075;
      520: inst = 32'h8220000;
      521: inst = 32'h10408000;
      522: inst = 32'hc404076;
      523: inst = 32'h8220000;
      524: inst = 32'h10408000;
      525: inst = 32'hc404077;
      526: inst = 32'h8220000;
      527: inst = 32'h10408000;
      528: inst = 32'hc404078;
      529: inst = 32'h8220000;
      530: inst = 32'h10408000;
      531: inst = 32'hc404079;
      532: inst = 32'h8220000;
      533: inst = 32'h10408000;
      534: inst = 32'hc40407a;
      535: inst = 32'h8220000;
      536: inst = 32'h10408000;
      537: inst = 32'hc40407b;
      538: inst = 32'h8220000;
      539: inst = 32'h10408000;
      540: inst = 32'hc40407c;
      541: inst = 32'h8220000;
      542: inst = 32'h10408000;
      543: inst = 32'hc40407d;
      544: inst = 32'h8220000;
      545: inst = 32'h10408000;
      546: inst = 32'hc40407e;
      547: inst = 32'h8220000;
      548: inst = 32'h10408000;
      549: inst = 32'hc40407f;
      550: inst = 32'h8220000;
      551: inst = 32'h10408000;
      552: inst = 32'hc404080;
      553: inst = 32'h8220000;
      554: inst = 32'h10408000;
      555: inst = 32'hc404081;
      556: inst = 32'h8220000;
      557: inst = 32'h10408000;
      558: inst = 32'hc404082;
      559: inst = 32'h8220000;
      560: inst = 32'h10408000;
      561: inst = 32'hc404083;
      562: inst = 32'h8220000;
      563: inst = 32'h10408000;
      564: inst = 32'hc404084;
      565: inst = 32'h8220000;
      566: inst = 32'h10408000;
      567: inst = 32'hc404085;
      568: inst = 32'h8220000;
      569: inst = 32'h10408000;
      570: inst = 32'hc404086;
      571: inst = 32'h8220000;
      572: inst = 32'h10408000;
      573: inst = 32'hc404087;
      574: inst = 32'h8220000;
      575: inst = 32'h10408000;
      576: inst = 32'hc404088;
      577: inst = 32'h8220000;
      578: inst = 32'h10408000;
      579: inst = 32'hc404089;
      580: inst = 32'h8220000;
      581: inst = 32'h10408000;
      582: inst = 32'hc40408a;
      583: inst = 32'h8220000;
      584: inst = 32'h10408000;
      585: inst = 32'hc40408b;
      586: inst = 32'h8220000;
      587: inst = 32'h10408000;
      588: inst = 32'hc40408c;
      589: inst = 32'h8220000;
      590: inst = 32'h10408000;
      591: inst = 32'hc40408d;
      592: inst = 32'h8220000;
      593: inst = 32'h10408000;
      594: inst = 32'hc40408e;
      595: inst = 32'h8220000;
      596: inst = 32'h10408000;
      597: inst = 32'hc40408f;
      598: inst = 32'h8220000;
      599: inst = 32'h10408000;
      600: inst = 32'hc404090;
      601: inst = 32'h8220000;
      602: inst = 32'h10408000;
      603: inst = 32'hc404091;
      604: inst = 32'h8220000;
      605: inst = 32'h10408000;
      606: inst = 32'hc404092;
      607: inst = 32'h8220000;
      608: inst = 32'h10408000;
      609: inst = 32'hc404093;
      610: inst = 32'h8220000;
      611: inst = 32'h10408000;
      612: inst = 32'hc404094;
      613: inst = 32'h8220000;
      614: inst = 32'h10408000;
      615: inst = 32'hc404095;
      616: inst = 32'h8220000;
      617: inst = 32'h10408000;
      618: inst = 32'hc404096;
      619: inst = 32'h8220000;
      620: inst = 32'h10408000;
      621: inst = 32'hc404097;
      622: inst = 32'h8220000;
      623: inst = 32'h10408000;
      624: inst = 32'hc404098;
      625: inst = 32'h8220000;
      626: inst = 32'h10408000;
      627: inst = 32'hc404099;
      628: inst = 32'h8220000;
      629: inst = 32'h10408000;
      630: inst = 32'hc40409a;
      631: inst = 32'h8220000;
      632: inst = 32'h10408000;
      633: inst = 32'hc40409b;
      634: inst = 32'h8220000;
      635: inst = 32'h10408000;
      636: inst = 32'hc40409c;
      637: inst = 32'h8220000;
      638: inst = 32'h10408000;
      639: inst = 32'hc40409d;
      640: inst = 32'h8220000;
      641: inst = 32'h10408000;
      642: inst = 32'hc40409e;
      643: inst = 32'h8220000;
      644: inst = 32'h10408000;
      645: inst = 32'hc40409f;
      646: inst = 32'h8220000;
      647: inst = 32'h10408000;
      648: inst = 32'hc4040a0;
      649: inst = 32'h8220000;
      650: inst = 32'h10408000;
      651: inst = 32'hc4040a1;
      652: inst = 32'h8220000;
      653: inst = 32'h10408000;
      654: inst = 32'hc4040a2;
      655: inst = 32'h8220000;
      656: inst = 32'h10408000;
      657: inst = 32'hc4040a3;
      658: inst = 32'h8220000;
      659: inst = 32'h10408000;
      660: inst = 32'hc4040a4;
      661: inst = 32'h8220000;
      662: inst = 32'h10408000;
      663: inst = 32'hc4040a5;
      664: inst = 32'h8220000;
      665: inst = 32'h10408000;
      666: inst = 32'hc4040a6;
      667: inst = 32'h8220000;
      668: inst = 32'h10408000;
      669: inst = 32'hc4040a7;
      670: inst = 32'h8220000;
      671: inst = 32'h10408000;
      672: inst = 32'hc4040a8;
      673: inst = 32'h8220000;
      674: inst = 32'h10408000;
      675: inst = 32'hc4040a9;
      676: inst = 32'h8220000;
      677: inst = 32'h10408000;
      678: inst = 32'hc4040aa;
      679: inst = 32'h8220000;
      680: inst = 32'h10408000;
      681: inst = 32'hc4040ac;
      682: inst = 32'h8220000;
      683: inst = 32'h10408000;
      684: inst = 32'hc4040ad;
      685: inst = 32'h8220000;
      686: inst = 32'h10408000;
      687: inst = 32'hc4040ae;
      688: inst = 32'h8220000;
      689: inst = 32'h10408000;
      690: inst = 32'hc4040af;
      691: inst = 32'h8220000;
      692: inst = 32'h10408000;
      693: inst = 32'hc4040b0;
      694: inst = 32'h8220000;
      695: inst = 32'h10408000;
      696: inst = 32'hc4040b1;
      697: inst = 32'h8220000;
      698: inst = 32'h10408000;
      699: inst = 32'hc4040b2;
      700: inst = 32'h8220000;
      701: inst = 32'h10408000;
      702: inst = 32'hc4040b3;
      703: inst = 32'h8220000;
      704: inst = 32'h10408000;
      705: inst = 32'hc4040b4;
      706: inst = 32'h8220000;
      707: inst = 32'h10408000;
      708: inst = 32'hc4040b5;
      709: inst = 32'h8220000;
      710: inst = 32'h10408000;
      711: inst = 32'hc4040b6;
      712: inst = 32'h8220000;
      713: inst = 32'h10408000;
      714: inst = 32'hc4040b7;
      715: inst = 32'h8220000;
      716: inst = 32'h10408000;
      717: inst = 32'hc4040b8;
      718: inst = 32'h8220000;
      719: inst = 32'h10408000;
      720: inst = 32'hc4040b9;
      721: inst = 32'h8220000;
      722: inst = 32'h10408000;
      723: inst = 32'hc4040ba;
      724: inst = 32'h8220000;
      725: inst = 32'h10408000;
      726: inst = 32'hc4040bb;
      727: inst = 32'h8220000;
      728: inst = 32'h10408000;
      729: inst = 32'hc4040bc;
      730: inst = 32'h8220000;
      731: inst = 32'h10408000;
      732: inst = 32'hc4040bd;
      733: inst = 32'h8220000;
      734: inst = 32'h10408000;
      735: inst = 32'hc4040be;
      736: inst = 32'h8220000;
      737: inst = 32'h10408000;
      738: inst = 32'hc4040bf;
      739: inst = 32'h8220000;
      740: inst = 32'h10408000;
      741: inst = 32'hc4040c0;
      742: inst = 32'h8220000;
      743: inst = 32'h10408000;
      744: inst = 32'hc4040c1;
      745: inst = 32'h8220000;
      746: inst = 32'h10408000;
      747: inst = 32'hc4040c2;
      748: inst = 32'h8220000;
      749: inst = 32'h10408000;
      750: inst = 32'hc4040c3;
      751: inst = 32'h8220000;
      752: inst = 32'h10408000;
      753: inst = 32'hc4040c4;
      754: inst = 32'h8220000;
      755: inst = 32'h10408000;
      756: inst = 32'hc4040c5;
      757: inst = 32'h8220000;
      758: inst = 32'h10408000;
      759: inst = 32'hc4040c6;
      760: inst = 32'h8220000;
      761: inst = 32'h10408000;
      762: inst = 32'hc4040c7;
      763: inst = 32'h8220000;
      764: inst = 32'h10408000;
      765: inst = 32'hc4040c8;
      766: inst = 32'h8220000;
      767: inst = 32'h10408000;
      768: inst = 32'hc4040c9;
      769: inst = 32'h8220000;
      770: inst = 32'h10408000;
      771: inst = 32'hc4040ca;
      772: inst = 32'h8220000;
      773: inst = 32'h10408000;
      774: inst = 32'hc4040cb;
      775: inst = 32'h8220000;
      776: inst = 32'h10408000;
      777: inst = 32'hc4040cc;
      778: inst = 32'h8220000;
      779: inst = 32'h10408000;
      780: inst = 32'hc4040cd;
      781: inst = 32'h8220000;
      782: inst = 32'h10408000;
      783: inst = 32'hc4040ce;
      784: inst = 32'h8220000;
      785: inst = 32'h10408000;
      786: inst = 32'hc4040cf;
      787: inst = 32'h8220000;
      788: inst = 32'h10408000;
      789: inst = 32'hc4040d0;
      790: inst = 32'h8220000;
      791: inst = 32'h10408000;
      792: inst = 32'hc4040d1;
      793: inst = 32'h8220000;
      794: inst = 32'h10408000;
      795: inst = 32'hc4040d2;
      796: inst = 32'h8220000;
      797: inst = 32'h10408000;
      798: inst = 32'hc4040d3;
      799: inst = 32'h8220000;
      800: inst = 32'h10408000;
      801: inst = 32'hc4040d4;
      802: inst = 32'h8220000;
      803: inst = 32'h10408000;
      804: inst = 32'hc4040d5;
      805: inst = 32'h8220000;
      806: inst = 32'h10408000;
      807: inst = 32'hc4040d6;
      808: inst = 32'h8220000;
      809: inst = 32'h10408000;
      810: inst = 32'hc4040d7;
      811: inst = 32'h8220000;
      812: inst = 32'h10408000;
      813: inst = 32'hc4040d8;
      814: inst = 32'h8220000;
      815: inst = 32'h10408000;
      816: inst = 32'hc4040d9;
      817: inst = 32'h8220000;
      818: inst = 32'h10408000;
      819: inst = 32'hc4040da;
      820: inst = 32'h8220000;
      821: inst = 32'h10408000;
      822: inst = 32'hc4040db;
      823: inst = 32'h8220000;
      824: inst = 32'h10408000;
      825: inst = 32'hc4040dc;
      826: inst = 32'h8220000;
      827: inst = 32'h10408000;
      828: inst = 32'hc4040dd;
      829: inst = 32'h8220000;
      830: inst = 32'h10408000;
      831: inst = 32'hc4040de;
      832: inst = 32'h8220000;
      833: inst = 32'h10408000;
      834: inst = 32'hc4040df;
      835: inst = 32'h8220000;
      836: inst = 32'h10408000;
      837: inst = 32'hc4040e0;
      838: inst = 32'h8220000;
      839: inst = 32'h10408000;
      840: inst = 32'hc4040e1;
      841: inst = 32'h8220000;
      842: inst = 32'h10408000;
      843: inst = 32'hc4040e2;
      844: inst = 32'h8220000;
      845: inst = 32'h10408000;
      846: inst = 32'hc4040e3;
      847: inst = 32'h8220000;
      848: inst = 32'h10408000;
      849: inst = 32'hc4040e4;
      850: inst = 32'h8220000;
      851: inst = 32'h10408000;
      852: inst = 32'hc4040e5;
      853: inst = 32'h8220000;
      854: inst = 32'h10408000;
      855: inst = 32'hc4040e6;
      856: inst = 32'h8220000;
      857: inst = 32'h10408000;
      858: inst = 32'hc4040e7;
      859: inst = 32'h8220000;
      860: inst = 32'h10408000;
      861: inst = 32'hc4040e8;
      862: inst = 32'h8220000;
      863: inst = 32'h10408000;
      864: inst = 32'hc4040e9;
      865: inst = 32'h8220000;
      866: inst = 32'h10408000;
      867: inst = 32'hc4040ea;
      868: inst = 32'h8220000;
      869: inst = 32'h10408000;
      870: inst = 32'hc4040eb;
      871: inst = 32'h8220000;
      872: inst = 32'h10408000;
      873: inst = 32'hc4040ec;
      874: inst = 32'h8220000;
      875: inst = 32'h10408000;
      876: inst = 32'hc4040ed;
      877: inst = 32'h8220000;
      878: inst = 32'h10408000;
      879: inst = 32'hc4040ee;
      880: inst = 32'h8220000;
      881: inst = 32'h10408000;
      882: inst = 32'hc4040ef;
      883: inst = 32'h8220000;
      884: inst = 32'h10408000;
      885: inst = 32'hc4040f0;
      886: inst = 32'h8220000;
      887: inst = 32'h10408000;
      888: inst = 32'hc4040f1;
      889: inst = 32'h8220000;
      890: inst = 32'h10408000;
      891: inst = 32'hc4040f2;
      892: inst = 32'h8220000;
      893: inst = 32'h10408000;
      894: inst = 32'hc4040f3;
      895: inst = 32'h8220000;
      896: inst = 32'h10408000;
      897: inst = 32'hc4040f4;
      898: inst = 32'h8220000;
      899: inst = 32'h10408000;
      900: inst = 32'hc4040f5;
      901: inst = 32'h8220000;
      902: inst = 32'h10408000;
      903: inst = 32'hc4040f6;
      904: inst = 32'h8220000;
      905: inst = 32'h10408000;
      906: inst = 32'hc4040f7;
      907: inst = 32'h8220000;
      908: inst = 32'h10408000;
      909: inst = 32'hc4040f8;
      910: inst = 32'h8220000;
      911: inst = 32'h10408000;
      912: inst = 32'hc4040f9;
      913: inst = 32'h8220000;
      914: inst = 32'h10408000;
      915: inst = 32'hc4040fa;
      916: inst = 32'h8220000;
      917: inst = 32'h10408000;
      918: inst = 32'hc4040fb;
      919: inst = 32'h8220000;
      920: inst = 32'h10408000;
      921: inst = 32'hc4040fc;
      922: inst = 32'h8220000;
      923: inst = 32'h10408000;
      924: inst = 32'hc4040fd;
      925: inst = 32'h8220000;
      926: inst = 32'h10408000;
      927: inst = 32'hc4040fe;
      928: inst = 32'h8220000;
      929: inst = 32'h10408000;
      930: inst = 32'hc4040ff;
      931: inst = 32'h8220000;
      932: inst = 32'h10408000;
      933: inst = 32'hc404100;
      934: inst = 32'h8220000;
      935: inst = 32'h10408000;
      936: inst = 32'hc404101;
      937: inst = 32'h8220000;
      938: inst = 32'h10408000;
      939: inst = 32'hc404102;
      940: inst = 32'h8220000;
      941: inst = 32'h10408000;
      942: inst = 32'hc404103;
      943: inst = 32'h8220000;
      944: inst = 32'h10408000;
      945: inst = 32'hc404104;
      946: inst = 32'h8220000;
      947: inst = 32'h10408000;
      948: inst = 32'hc404105;
      949: inst = 32'h8220000;
      950: inst = 32'h10408000;
      951: inst = 32'hc404106;
      952: inst = 32'h8220000;
      953: inst = 32'h10408000;
      954: inst = 32'hc404107;
      955: inst = 32'h8220000;
      956: inst = 32'h10408000;
      957: inst = 32'hc404108;
      958: inst = 32'h8220000;
      959: inst = 32'h10408000;
      960: inst = 32'hc404109;
      961: inst = 32'h8220000;
      962: inst = 32'h10408000;
      963: inst = 32'hc40410a;
      964: inst = 32'h8220000;
      965: inst = 32'h10408000;
      966: inst = 32'hc40410c;
      967: inst = 32'h8220000;
      968: inst = 32'h10408000;
      969: inst = 32'hc40410d;
      970: inst = 32'h8220000;
      971: inst = 32'h10408000;
      972: inst = 32'hc40410e;
      973: inst = 32'h8220000;
      974: inst = 32'h10408000;
      975: inst = 32'hc40410f;
      976: inst = 32'h8220000;
      977: inst = 32'h10408000;
      978: inst = 32'hc404110;
      979: inst = 32'h8220000;
      980: inst = 32'h10408000;
      981: inst = 32'hc404111;
      982: inst = 32'h8220000;
      983: inst = 32'h10408000;
      984: inst = 32'hc404112;
      985: inst = 32'h8220000;
      986: inst = 32'h10408000;
      987: inst = 32'hc404113;
      988: inst = 32'h8220000;
      989: inst = 32'h10408000;
      990: inst = 32'hc404114;
      991: inst = 32'h8220000;
      992: inst = 32'h10408000;
      993: inst = 32'hc404115;
      994: inst = 32'h8220000;
      995: inst = 32'h10408000;
      996: inst = 32'hc404116;
      997: inst = 32'h8220000;
      998: inst = 32'h10408000;
      999: inst = 32'hc404117;
      1000: inst = 32'h8220000;
      1001: inst = 32'h10408000;
      1002: inst = 32'hc404118;
      1003: inst = 32'h8220000;
      1004: inst = 32'h10408000;
      1005: inst = 32'hc404119;
      1006: inst = 32'h8220000;
      1007: inst = 32'h10408000;
      1008: inst = 32'hc40411a;
      1009: inst = 32'h8220000;
      1010: inst = 32'h10408000;
      1011: inst = 32'hc40411b;
      1012: inst = 32'h8220000;
      1013: inst = 32'h10408000;
      1014: inst = 32'hc40411c;
      1015: inst = 32'h8220000;
      1016: inst = 32'h10408000;
      1017: inst = 32'hc40411d;
      1018: inst = 32'h8220000;
      1019: inst = 32'h10408000;
      1020: inst = 32'hc40411e;
      1021: inst = 32'h8220000;
      1022: inst = 32'h10408000;
      1023: inst = 32'hc40411f;
      1024: inst = 32'h8220000;
      1025: inst = 32'h10408000;
      1026: inst = 32'hc404120;
      1027: inst = 32'h8220000;
      1028: inst = 32'h10408000;
      1029: inst = 32'hc404121;
      1030: inst = 32'h8220000;
      1031: inst = 32'h10408000;
      1032: inst = 32'hc404122;
      1033: inst = 32'h8220000;
      1034: inst = 32'h10408000;
      1035: inst = 32'hc404123;
      1036: inst = 32'h8220000;
      1037: inst = 32'h10408000;
      1038: inst = 32'hc404124;
      1039: inst = 32'h8220000;
      1040: inst = 32'h10408000;
      1041: inst = 32'hc404125;
      1042: inst = 32'h8220000;
      1043: inst = 32'h10408000;
      1044: inst = 32'hc404126;
      1045: inst = 32'h8220000;
      1046: inst = 32'h10408000;
      1047: inst = 32'hc404127;
      1048: inst = 32'h8220000;
      1049: inst = 32'h10408000;
      1050: inst = 32'hc404128;
      1051: inst = 32'h8220000;
      1052: inst = 32'h10408000;
      1053: inst = 32'hc404129;
      1054: inst = 32'h8220000;
      1055: inst = 32'h10408000;
      1056: inst = 32'hc40412a;
      1057: inst = 32'h8220000;
      1058: inst = 32'h10408000;
      1059: inst = 32'hc40412b;
      1060: inst = 32'h8220000;
      1061: inst = 32'h10408000;
      1062: inst = 32'hc40412c;
      1063: inst = 32'h8220000;
      1064: inst = 32'h10408000;
      1065: inst = 32'hc40412d;
      1066: inst = 32'h8220000;
      1067: inst = 32'h10408000;
      1068: inst = 32'hc40412e;
      1069: inst = 32'h8220000;
      1070: inst = 32'h10408000;
      1071: inst = 32'hc40412f;
      1072: inst = 32'h8220000;
      1073: inst = 32'h10408000;
      1074: inst = 32'hc404130;
      1075: inst = 32'h8220000;
      1076: inst = 32'h10408000;
      1077: inst = 32'hc404131;
      1078: inst = 32'h8220000;
      1079: inst = 32'h10408000;
      1080: inst = 32'hc404132;
      1081: inst = 32'h8220000;
      1082: inst = 32'h10408000;
      1083: inst = 32'hc404133;
      1084: inst = 32'h8220000;
      1085: inst = 32'h10408000;
      1086: inst = 32'hc404134;
      1087: inst = 32'h8220000;
      1088: inst = 32'h10408000;
      1089: inst = 32'hc404135;
      1090: inst = 32'h8220000;
      1091: inst = 32'h10408000;
      1092: inst = 32'hc404136;
      1093: inst = 32'h8220000;
      1094: inst = 32'h10408000;
      1095: inst = 32'hc404137;
      1096: inst = 32'h8220000;
      1097: inst = 32'h10408000;
      1098: inst = 32'hc404138;
      1099: inst = 32'h8220000;
      1100: inst = 32'h10408000;
      1101: inst = 32'hc404139;
      1102: inst = 32'h8220000;
      1103: inst = 32'h10408000;
      1104: inst = 32'hc40413a;
      1105: inst = 32'h8220000;
      1106: inst = 32'h10408000;
      1107: inst = 32'hc40413b;
      1108: inst = 32'h8220000;
      1109: inst = 32'h10408000;
      1110: inst = 32'hc40413c;
      1111: inst = 32'h8220000;
      1112: inst = 32'h10408000;
      1113: inst = 32'hc40413d;
      1114: inst = 32'h8220000;
      1115: inst = 32'h10408000;
      1116: inst = 32'hc40413e;
      1117: inst = 32'h8220000;
      1118: inst = 32'h10408000;
      1119: inst = 32'hc40413f;
      1120: inst = 32'h8220000;
      1121: inst = 32'h10408000;
      1122: inst = 32'hc404140;
      1123: inst = 32'h8220000;
      1124: inst = 32'h10408000;
      1125: inst = 32'hc404141;
      1126: inst = 32'h8220000;
      1127: inst = 32'h10408000;
      1128: inst = 32'hc404142;
      1129: inst = 32'h8220000;
      1130: inst = 32'h10408000;
      1131: inst = 32'hc404143;
      1132: inst = 32'h8220000;
      1133: inst = 32'h10408000;
      1134: inst = 32'hc404144;
      1135: inst = 32'h8220000;
      1136: inst = 32'h10408000;
      1137: inst = 32'hc404145;
      1138: inst = 32'h8220000;
      1139: inst = 32'h10408000;
      1140: inst = 32'hc404146;
      1141: inst = 32'h8220000;
      1142: inst = 32'h10408000;
      1143: inst = 32'hc404147;
      1144: inst = 32'h8220000;
      1145: inst = 32'h10408000;
      1146: inst = 32'hc404148;
      1147: inst = 32'h8220000;
      1148: inst = 32'h10408000;
      1149: inst = 32'hc404149;
      1150: inst = 32'h8220000;
      1151: inst = 32'h10408000;
      1152: inst = 32'hc40414a;
      1153: inst = 32'h8220000;
      1154: inst = 32'h10408000;
      1155: inst = 32'hc40414b;
      1156: inst = 32'h8220000;
      1157: inst = 32'h10408000;
      1158: inst = 32'hc40414c;
      1159: inst = 32'h8220000;
      1160: inst = 32'h10408000;
      1161: inst = 32'hc40414d;
      1162: inst = 32'h8220000;
      1163: inst = 32'h10408000;
      1164: inst = 32'hc40414e;
      1165: inst = 32'h8220000;
      1166: inst = 32'h10408000;
      1167: inst = 32'hc40414f;
      1168: inst = 32'h8220000;
      1169: inst = 32'h10408000;
      1170: inst = 32'hc404150;
      1171: inst = 32'h8220000;
      1172: inst = 32'h10408000;
      1173: inst = 32'hc404151;
      1174: inst = 32'h8220000;
      1175: inst = 32'h10408000;
      1176: inst = 32'hc404152;
      1177: inst = 32'h8220000;
      1178: inst = 32'h10408000;
      1179: inst = 32'hc404153;
      1180: inst = 32'h8220000;
      1181: inst = 32'h10408000;
      1182: inst = 32'hc404154;
      1183: inst = 32'h8220000;
      1184: inst = 32'h10408000;
      1185: inst = 32'hc404155;
      1186: inst = 32'h8220000;
      1187: inst = 32'h10408000;
      1188: inst = 32'hc404156;
      1189: inst = 32'h8220000;
      1190: inst = 32'h10408000;
      1191: inst = 32'hc404157;
      1192: inst = 32'h8220000;
      1193: inst = 32'h10408000;
      1194: inst = 32'hc404158;
      1195: inst = 32'h8220000;
      1196: inst = 32'h10408000;
      1197: inst = 32'hc404159;
      1198: inst = 32'h8220000;
      1199: inst = 32'h10408000;
      1200: inst = 32'hc40415a;
      1201: inst = 32'h8220000;
      1202: inst = 32'h10408000;
      1203: inst = 32'hc40415b;
      1204: inst = 32'h8220000;
      1205: inst = 32'h10408000;
      1206: inst = 32'hc40415c;
      1207: inst = 32'h8220000;
      1208: inst = 32'h10408000;
      1209: inst = 32'hc40415d;
      1210: inst = 32'h8220000;
      1211: inst = 32'h10408000;
      1212: inst = 32'hc40415e;
      1213: inst = 32'h8220000;
      1214: inst = 32'h10408000;
      1215: inst = 32'hc40415f;
      1216: inst = 32'h8220000;
      1217: inst = 32'h10408000;
      1218: inst = 32'hc404160;
      1219: inst = 32'h8220000;
      1220: inst = 32'h10408000;
      1221: inst = 32'hc404161;
      1222: inst = 32'h8220000;
      1223: inst = 32'h10408000;
      1224: inst = 32'hc404162;
      1225: inst = 32'h8220000;
      1226: inst = 32'h10408000;
      1227: inst = 32'hc404163;
      1228: inst = 32'h8220000;
      1229: inst = 32'h10408000;
      1230: inst = 32'hc404164;
      1231: inst = 32'h8220000;
      1232: inst = 32'h10408000;
      1233: inst = 32'hc404165;
      1234: inst = 32'h8220000;
      1235: inst = 32'h10408000;
      1236: inst = 32'hc404166;
      1237: inst = 32'h8220000;
      1238: inst = 32'h10408000;
      1239: inst = 32'hc404167;
      1240: inst = 32'h8220000;
      1241: inst = 32'h10408000;
      1242: inst = 32'hc404168;
      1243: inst = 32'h8220000;
      1244: inst = 32'h10408000;
      1245: inst = 32'hc404169;
      1246: inst = 32'h8220000;
      1247: inst = 32'h10408000;
      1248: inst = 32'hc40416a;
      1249: inst = 32'h8220000;
      1250: inst = 32'h10408000;
      1251: inst = 32'hc40416c;
      1252: inst = 32'h8220000;
      1253: inst = 32'h10408000;
      1254: inst = 32'hc40416d;
      1255: inst = 32'h8220000;
      1256: inst = 32'h10408000;
      1257: inst = 32'hc40416e;
      1258: inst = 32'h8220000;
      1259: inst = 32'h10408000;
      1260: inst = 32'hc40416f;
      1261: inst = 32'h8220000;
      1262: inst = 32'h10408000;
      1263: inst = 32'hc404170;
      1264: inst = 32'h8220000;
      1265: inst = 32'h10408000;
      1266: inst = 32'hc404171;
      1267: inst = 32'h8220000;
      1268: inst = 32'h10408000;
      1269: inst = 32'hc404172;
      1270: inst = 32'h8220000;
      1271: inst = 32'h10408000;
      1272: inst = 32'hc404173;
      1273: inst = 32'h8220000;
      1274: inst = 32'h10408000;
      1275: inst = 32'hc404174;
      1276: inst = 32'h8220000;
      1277: inst = 32'h10408000;
      1278: inst = 32'hc404175;
      1279: inst = 32'h8220000;
      1280: inst = 32'h10408000;
      1281: inst = 32'hc404176;
      1282: inst = 32'h8220000;
      1283: inst = 32'h10408000;
      1284: inst = 32'hc404177;
      1285: inst = 32'h8220000;
      1286: inst = 32'h10408000;
      1287: inst = 32'hc404178;
      1288: inst = 32'h8220000;
      1289: inst = 32'h10408000;
      1290: inst = 32'hc404179;
      1291: inst = 32'h8220000;
      1292: inst = 32'h10408000;
      1293: inst = 32'hc40417a;
      1294: inst = 32'h8220000;
      1295: inst = 32'h10408000;
      1296: inst = 32'hc40417b;
      1297: inst = 32'h8220000;
      1298: inst = 32'h10408000;
      1299: inst = 32'hc40417c;
      1300: inst = 32'h8220000;
      1301: inst = 32'h10408000;
      1302: inst = 32'hc40417d;
      1303: inst = 32'h8220000;
      1304: inst = 32'h10408000;
      1305: inst = 32'hc40417e;
      1306: inst = 32'h8220000;
      1307: inst = 32'h10408000;
      1308: inst = 32'hc40417f;
      1309: inst = 32'h8220000;
      1310: inst = 32'h10408000;
      1311: inst = 32'hc404180;
      1312: inst = 32'h8220000;
      1313: inst = 32'h10408000;
      1314: inst = 32'hc404181;
      1315: inst = 32'h8220000;
      1316: inst = 32'h10408000;
      1317: inst = 32'hc404182;
      1318: inst = 32'h8220000;
      1319: inst = 32'h10408000;
      1320: inst = 32'hc404183;
      1321: inst = 32'h8220000;
      1322: inst = 32'h10408000;
      1323: inst = 32'hc404184;
      1324: inst = 32'h8220000;
      1325: inst = 32'h10408000;
      1326: inst = 32'hc404185;
      1327: inst = 32'h8220000;
      1328: inst = 32'h10408000;
      1329: inst = 32'hc404186;
      1330: inst = 32'h8220000;
      1331: inst = 32'h10408000;
      1332: inst = 32'hc404187;
      1333: inst = 32'h8220000;
      1334: inst = 32'h10408000;
      1335: inst = 32'hc404188;
      1336: inst = 32'h8220000;
      1337: inst = 32'h10408000;
      1338: inst = 32'hc404189;
      1339: inst = 32'h8220000;
      1340: inst = 32'h10408000;
      1341: inst = 32'hc40418a;
      1342: inst = 32'h8220000;
      1343: inst = 32'h10408000;
      1344: inst = 32'hc40418b;
      1345: inst = 32'h8220000;
      1346: inst = 32'h10408000;
      1347: inst = 32'hc40418c;
      1348: inst = 32'h8220000;
      1349: inst = 32'h10408000;
      1350: inst = 32'hc40418d;
      1351: inst = 32'h8220000;
      1352: inst = 32'h10408000;
      1353: inst = 32'hc40418e;
      1354: inst = 32'h8220000;
      1355: inst = 32'h10408000;
      1356: inst = 32'hc40418f;
      1357: inst = 32'h8220000;
      1358: inst = 32'h10408000;
      1359: inst = 32'hc404190;
      1360: inst = 32'h8220000;
      1361: inst = 32'h10408000;
      1362: inst = 32'hc404191;
      1363: inst = 32'h8220000;
      1364: inst = 32'h10408000;
      1365: inst = 32'hc404192;
      1366: inst = 32'h8220000;
      1367: inst = 32'h10408000;
      1368: inst = 32'hc404193;
      1369: inst = 32'h8220000;
      1370: inst = 32'h10408000;
      1371: inst = 32'hc404194;
      1372: inst = 32'h8220000;
      1373: inst = 32'h10408000;
      1374: inst = 32'hc404195;
      1375: inst = 32'h8220000;
      1376: inst = 32'h10408000;
      1377: inst = 32'hc404196;
      1378: inst = 32'h8220000;
      1379: inst = 32'h10408000;
      1380: inst = 32'hc404197;
      1381: inst = 32'h8220000;
      1382: inst = 32'h10408000;
      1383: inst = 32'hc404198;
      1384: inst = 32'h8220000;
      1385: inst = 32'h10408000;
      1386: inst = 32'hc404199;
      1387: inst = 32'h8220000;
      1388: inst = 32'h10408000;
      1389: inst = 32'hc40419a;
      1390: inst = 32'h8220000;
      1391: inst = 32'h10408000;
      1392: inst = 32'hc40419b;
      1393: inst = 32'h8220000;
      1394: inst = 32'h10408000;
      1395: inst = 32'hc40419c;
      1396: inst = 32'h8220000;
      1397: inst = 32'h10408000;
      1398: inst = 32'hc40419d;
      1399: inst = 32'h8220000;
      1400: inst = 32'h10408000;
      1401: inst = 32'hc40419e;
      1402: inst = 32'h8220000;
      1403: inst = 32'h10408000;
      1404: inst = 32'hc40419f;
      1405: inst = 32'h8220000;
      1406: inst = 32'h10408000;
      1407: inst = 32'hc4041a0;
      1408: inst = 32'h8220000;
      1409: inst = 32'h10408000;
      1410: inst = 32'hc4041a1;
      1411: inst = 32'h8220000;
      1412: inst = 32'h10408000;
      1413: inst = 32'hc4041a2;
      1414: inst = 32'h8220000;
      1415: inst = 32'h10408000;
      1416: inst = 32'hc4041a3;
      1417: inst = 32'h8220000;
      1418: inst = 32'h10408000;
      1419: inst = 32'hc4041a4;
      1420: inst = 32'h8220000;
      1421: inst = 32'h10408000;
      1422: inst = 32'hc4041a5;
      1423: inst = 32'h8220000;
      1424: inst = 32'h10408000;
      1425: inst = 32'hc4041a6;
      1426: inst = 32'h8220000;
      1427: inst = 32'h10408000;
      1428: inst = 32'hc4041a7;
      1429: inst = 32'h8220000;
      1430: inst = 32'h10408000;
      1431: inst = 32'hc4041a8;
      1432: inst = 32'h8220000;
      1433: inst = 32'h10408000;
      1434: inst = 32'hc4041a9;
      1435: inst = 32'h8220000;
      1436: inst = 32'h10408000;
      1437: inst = 32'hc4041aa;
      1438: inst = 32'h8220000;
      1439: inst = 32'h10408000;
      1440: inst = 32'hc4041ab;
      1441: inst = 32'h8220000;
      1442: inst = 32'h10408000;
      1443: inst = 32'hc4041ac;
      1444: inst = 32'h8220000;
      1445: inst = 32'h10408000;
      1446: inst = 32'hc4041ad;
      1447: inst = 32'h8220000;
      1448: inst = 32'h10408000;
      1449: inst = 32'hc4041ae;
      1450: inst = 32'h8220000;
      1451: inst = 32'h10408000;
      1452: inst = 32'hc4041af;
      1453: inst = 32'h8220000;
      1454: inst = 32'h10408000;
      1455: inst = 32'hc4041b0;
      1456: inst = 32'h8220000;
      1457: inst = 32'h10408000;
      1458: inst = 32'hc4041b1;
      1459: inst = 32'h8220000;
      1460: inst = 32'h10408000;
      1461: inst = 32'hc4041b2;
      1462: inst = 32'h8220000;
      1463: inst = 32'h10408000;
      1464: inst = 32'hc4041b3;
      1465: inst = 32'h8220000;
      1466: inst = 32'h10408000;
      1467: inst = 32'hc4041b4;
      1468: inst = 32'h8220000;
      1469: inst = 32'h10408000;
      1470: inst = 32'hc4041b5;
      1471: inst = 32'h8220000;
      1472: inst = 32'h10408000;
      1473: inst = 32'hc4041b6;
      1474: inst = 32'h8220000;
      1475: inst = 32'h10408000;
      1476: inst = 32'hc4041b7;
      1477: inst = 32'h8220000;
      1478: inst = 32'h10408000;
      1479: inst = 32'hc4041b8;
      1480: inst = 32'h8220000;
      1481: inst = 32'h10408000;
      1482: inst = 32'hc4041b9;
      1483: inst = 32'h8220000;
      1484: inst = 32'h10408000;
      1485: inst = 32'hc4041ba;
      1486: inst = 32'h8220000;
      1487: inst = 32'h10408000;
      1488: inst = 32'hc4041bb;
      1489: inst = 32'h8220000;
      1490: inst = 32'h10408000;
      1491: inst = 32'hc4041bc;
      1492: inst = 32'h8220000;
      1493: inst = 32'h10408000;
      1494: inst = 32'hc4041bd;
      1495: inst = 32'h8220000;
      1496: inst = 32'h10408000;
      1497: inst = 32'hc4041be;
      1498: inst = 32'h8220000;
      1499: inst = 32'h10408000;
      1500: inst = 32'hc4041bf;
      1501: inst = 32'h8220000;
      1502: inst = 32'h10408000;
      1503: inst = 32'hc4041c0;
      1504: inst = 32'h8220000;
      1505: inst = 32'h10408000;
      1506: inst = 32'hc4041c1;
      1507: inst = 32'h8220000;
      1508: inst = 32'h10408000;
      1509: inst = 32'hc4041c2;
      1510: inst = 32'h8220000;
      1511: inst = 32'h10408000;
      1512: inst = 32'hc4041c3;
      1513: inst = 32'h8220000;
      1514: inst = 32'h10408000;
      1515: inst = 32'hc4041c4;
      1516: inst = 32'h8220000;
      1517: inst = 32'h10408000;
      1518: inst = 32'hc4041c5;
      1519: inst = 32'h8220000;
      1520: inst = 32'h10408000;
      1521: inst = 32'hc4041c6;
      1522: inst = 32'h8220000;
      1523: inst = 32'h10408000;
      1524: inst = 32'hc4041c7;
      1525: inst = 32'h8220000;
      1526: inst = 32'h10408000;
      1527: inst = 32'hc4041c8;
      1528: inst = 32'h8220000;
      1529: inst = 32'h10408000;
      1530: inst = 32'hc4041c9;
      1531: inst = 32'h8220000;
      1532: inst = 32'h10408000;
      1533: inst = 32'hc4041ca;
      1534: inst = 32'h8220000;
      1535: inst = 32'h10408000;
      1536: inst = 32'hc4041cc;
      1537: inst = 32'h8220000;
      1538: inst = 32'h10408000;
      1539: inst = 32'hc4041cd;
      1540: inst = 32'h8220000;
      1541: inst = 32'h10408000;
      1542: inst = 32'hc4041ce;
      1543: inst = 32'h8220000;
      1544: inst = 32'h10408000;
      1545: inst = 32'hc4041cf;
      1546: inst = 32'h8220000;
      1547: inst = 32'h10408000;
      1548: inst = 32'hc4041d0;
      1549: inst = 32'h8220000;
      1550: inst = 32'h10408000;
      1551: inst = 32'hc4041d1;
      1552: inst = 32'h8220000;
      1553: inst = 32'h10408000;
      1554: inst = 32'hc4041d2;
      1555: inst = 32'h8220000;
      1556: inst = 32'h10408000;
      1557: inst = 32'hc4041d3;
      1558: inst = 32'h8220000;
      1559: inst = 32'h10408000;
      1560: inst = 32'hc4041d4;
      1561: inst = 32'h8220000;
      1562: inst = 32'h10408000;
      1563: inst = 32'hc4041d5;
      1564: inst = 32'h8220000;
      1565: inst = 32'h10408000;
      1566: inst = 32'hc4041d6;
      1567: inst = 32'h8220000;
      1568: inst = 32'h10408000;
      1569: inst = 32'hc4041d7;
      1570: inst = 32'h8220000;
      1571: inst = 32'h10408000;
      1572: inst = 32'hc4041d8;
      1573: inst = 32'h8220000;
      1574: inst = 32'h10408000;
      1575: inst = 32'hc4041d9;
      1576: inst = 32'h8220000;
      1577: inst = 32'h10408000;
      1578: inst = 32'hc404206;
      1579: inst = 32'h8220000;
      1580: inst = 32'h10408000;
      1581: inst = 32'hc404207;
      1582: inst = 32'h8220000;
      1583: inst = 32'h10408000;
      1584: inst = 32'hc404208;
      1585: inst = 32'h8220000;
      1586: inst = 32'h10408000;
      1587: inst = 32'hc404209;
      1588: inst = 32'h8220000;
      1589: inst = 32'h10408000;
      1590: inst = 32'hc40420a;
      1591: inst = 32'h8220000;
      1592: inst = 32'h10408000;
      1593: inst = 32'hc40420b;
      1594: inst = 32'h8220000;
      1595: inst = 32'h10408000;
      1596: inst = 32'hc40420c;
      1597: inst = 32'h8220000;
      1598: inst = 32'h10408000;
      1599: inst = 32'hc40420d;
      1600: inst = 32'h8220000;
      1601: inst = 32'h10408000;
      1602: inst = 32'hc40420e;
      1603: inst = 32'h8220000;
      1604: inst = 32'h10408000;
      1605: inst = 32'hc40420f;
      1606: inst = 32'h8220000;
      1607: inst = 32'h10408000;
      1608: inst = 32'hc404210;
      1609: inst = 32'h8220000;
      1610: inst = 32'h10408000;
      1611: inst = 32'hc404211;
      1612: inst = 32'h8220000;
      1613: inst = 32'h10408000;
      1614: inst = 32'hc404212;
      1615: inst = 32'h8220000;
      1616: inst = 32'h10408000;
      1617: inst = 32'hc404213;
      1618: inst = 32'h8220000;
      1619: inst = 32'h10408000;
      1620: inst = 32'hc404214;
      1621: inst = 32'h8220000;
      1622: inst = 32'h10408000;
      1623: inst = 32'hc404215;
      1624: inst = 32'h8220000;
      1625: inst = 32'h10408000;
      1626: inst = 32'hc404216;
      1627: inst = 32'h8220000;
      1628: inst = 32'h10408000;
      1629: inst = 32'hc404217;
      1630: inst = 32'h8220000;
      1631: inst = 32'h10408000;
      1632: inst = 32'hc404218;
      1633: inst = 32'h8220000;
      1634: inst = 32'h10408000;
      1635: inst = 32'hc404219;
      1636: inst = 32'h8220000;
      1637: inst = 32'h10408000;
      1638: inst = 32'hc40421a;
      1639: inst = 32'h8220000;
      1640: inst = 32'h10408000;
      1641: inst = 32'hc40421b;
      1642: inst = 32'h8220000;
      1643: inst = 32'h10408000;
      1644: inst = 32'hc40421c;
      1645: inst = 32'h8220000;
      1646: inst = 32'h10408000;
      1647: inst = 32'hc40421d;
      1648: inst = 32'h8220000;
      1649: inst = 32'h10408000;
      1650: inst = 32'hc40421e;
      1651: inst = 32'h8220000;
      1652: inst = 32'h10408000;
      1653: inst = 32'hc40421f;
      1654: inst = 32'h8220000;
      1655: inst = 32'h10408000;
      1656: inst = 32'hc404220;
      1657: inst = 32'h8220000;
      1658: inst = 32'h10408000;
      1659: inst = 32'hc404221;
      1660: inst = 32'h8220000;
      1661: inst = 32'h10408000;
      1662: inst = 32'hc404222;
      1663: inst = 32'h8220000;
      1664: inst = 32'h10408000;
      1665: inst = 32'hc404223;
      1666: inst = 32'h8220000;
      1667: inst = 32'h10408000;
      1668: inst = 32'hc404224;
      1669: inst = 32'h8220000;
      1670: inst = 32'h10408000;
      1671: inst = 32'hc404225;
      1672: inst = 32'h8220000;
      1673: inst = 32'h10408000;
      1674: inst = 32'hc404226;
      1675: inst = 32'h8220000;
      1676: inst = 32'h10408000;
      1677: inst = 32'hc404227;
      1678: inst = 32'h8220000;
      1679: inst = 32'h10408000;
      1680: inst = 32'hc404228;
      1681: inst = 32'h8220000;
      1682: inst = 32'h10408000;
      1683: inst = 32'hc404229;
      1684: inst = 32'h8220000;
      1685: inst = 32'h10408000;
      1686: inst = 32'hc40422a;
      1687: inst = 32'h8220000;
      1688: inst = 32'h10408000;
      1689: inst = 32'hc40422c;
      1690: inst = 32'h8220000;
      1691: inst = 32'h10408000;
      1692: inst = 32'hc40422d;
      1693: inst = 32'h8220000;
      1694: inst = 32'h10408000;
      1695: inst = 32'hc40422e;
      1696: inst = 32'h8220000;
      1697: inst = 32'h10408000;
      1698: inst = 32'hc40422f;
      1699: inst = 32'h8220000;
      1700: inst = 32'h10408000;
      1701: inst = 32'hc404230;
      1702: inst = 32'h8220000;
      1703: inst = 32'h10408000;
      1704: inst = 32'hc404231;
      1705: inst = 32'h8220000;
      1706: inst = 32'h10408000;
      1707: inst = 32'hc404232;
      1708: inst = 32'h8220000;
      1709: inst = 32'h10408000;
      1710: inst = 32'hc404233;
      1711: inst = 32'h8220000;
      1712: inst = 32'h10408000;
      1713: inst = 32'hc404234;
      1714: inst = 32'h8220000;
      1715: inst = 32'h10408000;
      1716: inst = 32'hc404235;
      1717: inst = 32'h8220000;
      1718: inst = 32'h10408000;
      1719: inst = 32'hc404236;
      1720: inst = 32'h8220000;
      1721: inst = 32'h10408000;
      1722: inst = 32'hc404237;
      1723: inst = 32'h8220000;
      1724: inst = 32'h10408000;
      1725: inst = 32'hc404238;
      1726: inst = 32'h8220000;
      1727: inst = 32'h10408000;
      1728: inst = 32'hc404239;
      1729: inst = 32'h8220000;
      1730: inst = 32'h10408000;
      1731: inst = 32'hc40423a;
      1732: inst = 32'h8220000;
      1733: inst = 32'h10408000;
      1734: inst = 32'hc40423b;
      1735: inst = 32'h8220000;
      1736: inst = 32'h10408000;
      1737: inst = 32'hc404264;
      1738: inst = 32'h8220000;
      1739: inst = 32'h10408000;
      1740: inst = 32'hc404265;
      1741: inst = 32'h8220000;
      1742: inst = 32'h10408000;
      1743: inst = 32'hc404266;
      1744: inst = 32'h8220000;
      1745: inst = 32'h10408000;
      1746: inst = 32'hc404267;
      1747: inst = 32'h8220000;
      1748: inst = 32'h10408000;
      1749: inst = 32'hc404268;
      1750: inst = 32'h8220000;
      1751: inst = 32'h10408000;
      1752: inst = 32'hc404269;
      1753: inst = 32'h8220000;
      1754: inst = 32'h10408000;
      1755: inst = 32'hc40426a;
      1756: inst = 32'h8220000;
      1757: inst = 32'h10408000;
      1758: inst = 32'hc40426b;
      1759: inst = 32'h8220000;
      1760: inst = 32'h10408000;
      1761: inst = 32'hc40426c;
      1762: inst = 32'h8220000;
      1763: inst = 32'h10408000;
      1764: inst = 32'hc40426d;
      1765: inst = 32'h8220000;
      1766: inst = 32'h10408000;
      1767: inst = 32'hc40426e;
      1768: inst = 32'h8220000;
      1769: inst = 32'h10408000;
      1770: inst = 32'hc40426f;
      1771: inst = 32'h8220000;
      1772: inst = 32'h10408000;
      1773: inst = 32'hc404270;
      1774: inst = 32'h8220000;
      1775: inst = 32'h10408000;
      1776: inst = 32'hc404271;
      1777: inst = 32'h8220000;
      1778: inst = 32'h10408000;
      1779: inst = 32'hc404272;
      1780: inst = 32'h8220000;
      1781: inst = 32'h10408000;
      1782: inst = 32'hc404273;
      1783: inst = 32'h8220000;
      1784: inst = 32'h10408000;
      1785: inst = 32'hc404274;
      1786: inst = 32'h8220000;
      1787: inst = 32'h10408000;
      1788: inst = 32'hc404275;
      1789: inst = 32'h8220000;
      1790: inst = 32'h10408000;
      1791: inst = 32'hc404276;
      1792: inst = 32'h8220000;
      1793: inst = 32'h10408000;
      1794: inst = 32'hc404277;
      1795: inst = 32'h8220000;
      1796: inst = 32'h10408000;
      1797: inst = 32'hc404278;
      1798: inst = 32'h8220000;
      1799: inst = 32'h10408000;
      1800: inst = 32'hc404279;
      1801: inst = 32'h8220000;
      1802: inst = 32'h10408000;
      1803: inst = 32'hc40427a;
      1804: inst = 32'h8220000;
      1805: inst = 32'h10408000;
      1806: inst = 32'hc40427b;
      1807: inst = 32'h8220000;
      1808: inst = 32'h10408000;
      1809: inst = 32'hc40427c;
      1810: inst = 32'h8220000;
      1811: inst = 32'h10408000;
      1812: inst = 32'hc40427d;
      1813: inst = 32'h8220000;
      1814: inst = 32'h10408000;
      1815: inst = 32'hc40427e;
      1816: inst = 32'h8220000;
      1817: inst = 32'h10408000;
      1818: inst = 32'hc40427f;
      1819: inst = 32'h8220000;
      1820: inst = 32'h10408000;
      1821: inst = 32'hc404280;
      1822: inst = 32'h8220000;
      1823: inst = 32'h10408000;
      1824: inst = 32'hc404281;
      1825: inst = 32'h8220000;
      1826: inst = 32'h10408000;
      1827: inst = 32'hc404282;
      1828: inst = 32'h8220000;
      1829: inst = 32'h10408000;
      1830: inst = 32'hc404283;
      1831: inst = 32'h8220000;
      1832: inst = 32'h10408000;
      1833: inst = 32'hc404284;
      1834: inst = 32'h8220000;
      1835: inst = 32'h10408000;
      1836: inst = 32'hc404285;
      1837: inst = 32'h8220000;
      1838: inst = 32'h10408000;
      1839: inst = 32'hc404286;
      1840: inst = 32'h8220000;
      1841: inst = 32'h10408000;
      1842: inst = 32'hc404287;
      1843: inst = 32'h8220000;
      1844: inst = 32'h10408000;
      1845: inst = 32'hc404288;
      1846: inst = 32'h8220000;
      1847: inst = 32'h10408000;
      1848: inst = 32'hc404289;
      1849: inst = 32'h8220000;
      1850: inst = 32'h10408000;
      1851: inst = 32'hc40428a;
      1852: inst = 32'h8220000;
      1853: inst = 32'h10408000;
      1854: inst = 32'hc40428c;
      1855: inst = 32'h8220000;
      1856: inst = 32'h10408000;
      1857: inst = 32'hc40428d;
      1858: inst = 32'h8220000;
      1859: inst = 32'h10408000;
      1860: inst = 32'hc40428e;
      1861: inst = 32'h8220000;
      1862: inst = 32'h10408000;
      1863: inst = 32'hc40428f;
      1864: inst = 32'h8220000;
      1865: inst = 32'h10408000;
      1866: inst = 32'hc404290;
      1867: inst = 32'h8220000;
      1868: inst = 32'h10408000;
      1869: inst = 32'hc404291;
      1870: inst = 32'h8220000;
      1871: inst = 32'h10408000;
      1872: inst = 32'hc404292;
      1873: inst = 32'h8220000;
      1874: inst = 32'h10408000;
      1875: inst = 32'hc404293;
      1876: inst = 32'h8220000;
      1877: inst = 32'h10408000;
      1878: inst = 32'hc404294;
      1879: inst = 32'h8220000;
      1880: inst = 32'h10408000;
      1881: inst = 32'hc404295;
      1882: inst = 32'h8220000;
      1883: inst = 32'h10408000;
      1884: inst = 32'hc404296;
      1885: inst = 32'h8220000;
      1886: inst = 32'h10408000;
      1887: inst = 32'hc404297;
      1888: inst = 32'h8220000;
      1889: inst = 32'h10408000;
      1890: inst = 32'hc404298;
      1891: inst = 32'h8220000;
      1892: inst = 32'h10408000;
      1893: inst = 32'hc404299;
      1894: inst = 32'h8220000;
      1895: inst = 32'h10408000;
      1896: inst = 32'hc40429a;
      1897: inst = 32'h8220000;
      1898: inst = 32'h10408000;
      1899: inst = 32'hc40429b;
      1900: inst = 32'h8220000;
      1901: inst = 32'h10408000;
      1902: inst = 32'hc4042c4;
      1903: inst = 32'h8220000;
      1904: inst = 32'h10408000;
      1905: inst = 32'hc4042c5;
      1906: inst = 32'h8220000;
      1907: inst = 32'h10408000;
      1908: inst = 32'hc4042c6;
      1909: inst = 32'h8220000;
      1910: inst = 32'h10408000;
      1911: inst = 32'hc4042c7;
      1912: inst = 32'h8220000;
      1913: inst = 32'h10408000;
      1914: inst = 32'hc4042c8;
      1915: inst = 32'h8220000;
      1916: inst = 32'h10408000;
      1917: inst = 32'hc4042c9;
      1918: inst = 32'h8220000;
      1919: inst = 32'h10408000;
      1920: inst = 32'hc4042ca;
      1921: inst = 32'h8220000;
      1922: inst = 32'h10408000;
      1923: inst = 32'hc4042cb;
      1924: inst = 32'h8220000;
      1925: inst = 32'h10408000;
      1926: inst = 32'hc4042cc;
      1927: inst = 32'h8220000;
      1928: inst = 32'h10408000;
      1929: inst = 32'hc4042cd;
      1930: inst = 32'h8220000;
      1931: inst = 32'h10408000;
      1932: inst = 32'hc4042ce;
      1933: inst = 32'h8220000;
      1934: inst = 32'h10408000;
      1935: inst = 32'hc4042cf;
      1936: inst = 32'h8220000;
      1937: inst = 32'h10408000;
      1938: inst = 32'hc4042d0;
      1939: inst = 32'h8220000;
      1940: inst = 32'h10408000;
      1941: inst = 32'hc4042d1;
      1942: inst = 32'h8220000;
      1943: inst = 32'h10408000;
      1944: inst = 32'hc4042d2;
      1945: inst = 32'h8220000;
      1946: inst = 32'h10408000;
      1947: inst = 32'hc4042d3;
      1948: inst = 32'h8220000;
      1949: inst = 32'h10408000;
      1950: inst = 32'hc4042d4;
      1951: inst = 32'h8220000;
      1952: inst = 32'h10408000;
      1953: inst = 32'hc4042d5;
      1954: inst = 32'h8220000;
      1955: inst = 32'h10408000;
      1956: inst = 32'hc4042d6;
      1957: inst = 32'h8220000;
      1958: inst = 32'h10408000;
      1959: inst = 32'hc4042d7;
      1960: inst = 32'h8220000;
      1961: inst = 32'h10408000;
      1962: inst = 32'hc4042d8;
      1963: inst = 32'h8220000;
      1964: inst = 32'h10408000;
      1965: inst = 32'hc4042d9;
      1966: inst = 32'h8220000;
      1967: inst = 32'h10408000;
      1968: inst = 32'hc4042da;
      1969: inst = 32'h8220000;
      1970: inst = 32'h10408000;
      1971: inst = 32'hc4042db;
      1972: inst = 32'h8220000;
      1973: inst = 32'h10408000;
      1974: inst = 32'hc4042dc;
      1975: inst = 32'h8220000;
      1976: inst = 32'h10408000;
      1977: inst = 32'hc4042dd;
      1978: inst = 32'h8220000;
      1979: inst = 32'h10408000;
      1980: inst = 32'hc4042de;
      1981: inst = 32'h8220000;
      1982: inst = 32'h10408000;
      1983: inst = 32'hc4042df;
      1984: inst = 32'h8220000;
      1985: inst = 32'h10408000;
      1986: inst = 32'hc4042e0;
      1987: inst = 32'h8220000;
      1988: inst = 32'h10408000;
      1989: inst = 32'hc4042e1;
      1990: inst = 32'h8220000;
      1991: inst = 32'h10408000;
      1992: inst = 32'hc4042e2;
      1993: inst = 32'h8220000;
      1994: inst = 32'h10408000;
      1995: inst = 32'hc4042e3;
      1996: inst = 32'h8220000;
      1997: inst = 32'h10408000;
      1998: inst = 32'hc4042e4;
      1999: inst = 32'h8220000;
      2000: inst = 32'h10408000;
      2001: inst = 32'hc4042e5;
      2002: inst = 32'h8220000;
      2003: inst = 32'h10408000;
      2004: inst = 32'hc4042e6;
      2005: inst = 32'h8220000;
      2006: inst = 32'h10408000;
      2007: inst = 32'hc4042e7;
      2008: inst = 32'h8220000;
      2009: inst = 32'h10408000;
      2010: inst = 32'hc4042e8;
      2011: inst = 32'h8220000;
      2012: inst = 32'h10408000;
      2013: inst = 32'hc4042e9;
      2014: inst = 32'h8220000;
      2015: inst = 32'h10408000;
      2016: inst = 32'hc4042ee;
      2017: inst = 32'h8220000;
      2018: inst = 32'h10408000;
      2019: inst = 32'hc4042ef;
      2020: inst = 32'h8220000;
      2021: inst = 32'h10408000;
      2022: inst = 32'hc4042f0;
      2023: inst = 32'h8220000;
      2024: inst = 32'h10408000;
      2025: inst = 32'hc4042f1;
      2026: inst = 32'h8220000;
      2027: inst = 32'h10408000;
      2028: inst = 32'hc4042f2;
      2029: inst = 32'h8220000;
      2030: inst = 32'h10408000;
      2031: inst = 32'hc4042f3;
      2032: inst = 32'h8220000;
      2033: inst = 32'h10408000;
      2034: inst = 32'hc4042f4;
      2035: inst = 32'h8220000;
      2036: inst = 32'h10408000;
      2037: inst = 32'hc4042f5;
      2038: inst = 32'h8220000;
      2039: inst = 32'h10408000;
      2040: inst = 32'hc4042f6;
      2041: inst = 32'h8220000;
      2042: inst = 32'h10408000;
      2043: inst = 32'hc4042f7;
      2044: inst = 32'h8220000;
      2045: inst = 32'h10408000;
      2046: inst = 32'hc4042f8;
      2047: inst = 32'h8220000;
      2048: inst = 32'h10408000;
      2049: inst = 32'hc4042f9;
      2050: inst = 32'h8220000;
      2051: inst = 32'h10408000;
      2052: inst = 32'hc4042fa;
      2053: inst = 32'h8220000;
      2054: inst = 32'h10408000;
      2055: inst = 32'hc4042fb;
      2056: inst = 32'h8220000;
      2057: inst = 32'h10408000;
      2058: inst = 32'hc404324;
      2059: inst = 32'h8220000;
      2060: inst = 32'h10408000;
      2061: inst = 32'hc404325;
      2062: inst = 32'h8220000;
      2063: inst = 32'h10408000;
      2064: inst = 32'hc404326;
      2065: inst = 32'h8220000;
      2066: inst = 32'h10408000;
      2067: inst = 32'hc404327;
      2068: inst = 32'h8220000;
      2069: inst = 32'h10408000;
      2070: inst = 32'hc404328;
      2071: inst = 32'h8220000;
      2072: inst = 32'h10408000;
      2073: inst = 32'hc404329;
      2074: inst = 32'h8220000;
      2075: inst = 32'h10408000;
      2076: inst = 32'hc40432a;
      2077: inst = 32'h8220000;
      2078: inst = 32'h10408000;
      2079: inst = 32'hc40432b;
      2080: inst = 32'h8220000;
      2081: inst = 32'h10408000;
      2082: inst = 32'hc40432c;
      2083: inst = 32'h8220000;
      2084: inst = 32'h10408000;
      2085: inst = 32'hc40432d;
      2086: inst = 32'h8220000;
      2087: inst = 32'h10408000;
      2088: inst = 32'hc40432e;
      2089: inst = 32'h8220000;
      2090: inst = 32'h10408000;
      2091: inst = 32'hc40432f;
      2092: inst = 32'h8220000;
      2093: inst = 32'h10408000;
      2094: inst = 32'hc404330;
      2095: inst = 32'h8220000;
      2096: inst = 32'h10408000;
      2097: inst = 32'hc404331;
      2098: inst = 32'h8220000;
      2099: inst = 32'h10408000;
      2100: inst = 32'hc404332;
      2101: inst = 32'h8220000;
      2102: inst = 32'h10408000;
      2103: inst = 32'hc404333;
      2104: inst = 32'h8220000;
      2105: inst = 32'h10408000;
      2106: inst = 32'hc404334;
      2107: inst = 32'h8220000;
      2108: inst = 32'h10408000;
      2109: inst = 32'hc404335;
      2110: inst = 32'h8220000;
      2111: inst = 32'h10408000;
      2112: inst = 32'hc404336;
      2113: inst = 32'h8220000;
      2114: inst = 32'h10408000;
      2115: inst = 32'hc404337;
      2116: inst = 32'h8220000;
      2117: inst = 32'h10408000;
      2118: inst = 32'hc404338;
      2119: inst = 32'h8220000;
      2120: inst = 32'h10408000;
      2121: inst = 32'hc404339;
      2122: inst = 32'h8220000;
      2123: inst = 32'h10408000;
      2124: inst = 32'hc40433a;
      2125: inst = 32'h8220000;
      2126: inst = 32'h10408000;
      2127: inst = 32'hc40433b;
      2128: inst = 32'h8220000;
      2129: inst = 32'h10408000;
      2130: inst = 32'hc40433c;
      2131: inst = 32'h8220000;
      2132: inst = 32'h10408000;
      2133: inst = 32'hc40433d;
      2134: inst = 32'h8220000;
      2135: inst = 32'h10408000;
      2136: inst = 32'hc40433e;
      2137: inst = 32'h8220000;
      2138: inst = 32'h10408000;
      2139: inst = 32'hc40433f;
      2140: inst = 32'h8220000;
      2141: inst = 32'h10408000;
      2142: inst = 32'hc404340;
      2143: inst = 32'h8220000;
      2144: inst = 32'h10408000;
      2145: inst = 32'hc404341;
      2146: inst = 32'h8220000;
      2147: inst = 32'h10408000;
      2148: inst = 32'hc404342;
      2149: inst = 32'h8220000;
      2150: inst = 32'h10408000;
      2151: inst = 32'hc404343;
      2152: inst = 32'h8220000;
      2153: inst = 32'h10408000;
      2154: inst = 32'hc404344;
      2155: inst = 32'h8220000;
      2156: inst = 32'h10408000;
      2157: inst = 32'hc404345;
      2158: inst = 32'h8220000;
      2159: inst = 32'h10408000;
      2160: inst = 32'hc404346;
      2161: inst = 32'h8220000;
      2162: inst = 32'h10408000;
      2163: inst = 32'hc404347;
      2164: inst = 32'h8220000;
      2165: inst = 32'h10408000;
      2166: inst = 32'hc404348;
      2167: inst = 32'h8220000;
      2168: inst = 32'h10408000;
      2169: inst = 32'hc40434f;
      2170: inst = 32'h8220000;
      2171: inst = 32'h10408000;
      2172: inst = 32'hc404350;
      2173: inst = 32'h8220000;
      2174: inst = 32'h10408000;
      2175: inst = 32'hc404351;
      2176: inst = 32'h8220000;
      2177: inst = 32'h10408000;
      2178: inst = 32'hc404352;
      2179: inst = 32'h8220000;
      2180: inst = 32'h10408000;
      2181: inst = 32'hc404353;
      2182: inst = 32'h8220000;
      2183: inst = 32'h10408000;
      2184: inst = 32'hc404354;
      2185: inst = 32'h8220000;
      2186: inst = 32'h10408000;
      2187: inst = 32'hc404355;
      2188: inst = 32'h8220000;
      2189: inst = 32'h10408000;
      2190: inst = 32'hc404356;
      2191: inst = 32'h8220000;
      2192: inst = 32'h10408000;
      2193: inst = 32'hc404357;
      2194: inst = 32'h8220000;
      2195: inst = 32'h10408000;
      2196: inst = 32'hc404358;
      2197: inst = 32'h8220000;
      2198: inst = 32'h10408000;
      2199: inst = 32'hc404359;
      2200: inst = 32'h8220000;
      2201: inst = 32'h10408000;
      2202: inst = 32'hc40435a;
      2203: inst = 32'h8220000;
      2204: inst = 32'h10408000;
      2205: inst = 32'hc40435b;
      2206: inst = 32'h8220000;
      2207: inst = 32'h10408000;
      2208: inst = 32'hc404384;
      2209: inst = 32'h8220000;
      2210: inst = 32'h10408000;
      2211: inst = 32'hc404385;
      2212: inst = 32'h8220000;
      2213: inst = 32'h10408000;
      2214: inst = 32'hc404386;
      2215: inst = 32'h8220000;
      2216: inst = 32'h10408000;
      2217: inst = 32'hc404387;
      2218: inst = 32'h8220000;
      2219: inst = 32'h10408000;
      2220: inst = 32'hc404388;
      2221: inst = 32'h8220000;
      2222: inst = 32'h10408000;
      2223: inst = 32'hc404389;
      2224: inst = 32'h8220000;
      2225: inst = 32'h10408000;
      2226: inst = 32'hc40438a;
      2227: inst = 32'h8220000;
      2228: inst = 32'h10408000;
      2229: inst = 32'hc40438b;
      2230: inst = 32'h8220000;
      2231: inst = 32'h10408000;
      2232: inst = 32'hc40438c;
      2233: inst = 32'h8220000;
      2234: inst = 32'h10408000;
      2235: inst = 32'hc40438d;
      2236: inst = 32'h8220000;
      2237: inst = 32'h10408000;
      2238: inst = 32'hc40438e;
      2239: inst = 32'h8220000;
      2240: inst = 32'h10408000;
      2241: inst = 32'hc40438f;
      2242: inst = 32'h8220000;
      2243: inst = 32'h10408000;
      2244: inst = 32'hc404390;
      2245: inst = 32'h8220000;
      2246: inst = 32'h10408000;
      2247: inst = 32'hc404391;
      2248: inst = 32'h8220000;
      2249: inst = 32'h10408000;
      2250: inst = 32'hc404392;
      2251: inst = 32'h8220000;
      2252: inst = 32'h10408000;
      2253: inst = 32'hc404393;
      2254: inst = 32'h8220000;
      2255: inst = 32'h10408000;
      2256: inst = 32'hc404394;
      2257: inst = 32'h8220000;
      2258: inst = 32'h10408000;
      2259: inst = 32'hc404395;
      2260: inst = 32'h8220000;
      2261: inst = 32'h10408000;
      2262: inst = 32'hc404396;
      2263: inst = 32'h8220000;
      2264: inst = 32'h10408000;
      2265: inst = 32'hc404397;
      2266: inst = 32'h8220000;
      2267: inst = 32'h10408000;
      2268: inst = 32'hc404398;
      2269: inst = 32'h8220000;
      2270: inst = 32'h10408000;
      2271: inst = 32'hc404399;
      2272: inst = 32'h8220000;
      2273: inst = 32'h10408000;
      2274: inst = 32'hc40439a;
      2275: inst = 32'h8220000;
      2276: inst = 32'h10408000;
      2277: inst = 32'hc40439b;
      2278: inst = 32'h8220000;
      2279: inst = 32'h10408000;
      2280: inst = 32'hc40439c;
      2281: inst = 32'h8220000;
      2282: inst = 32'h10408000;
      2283: inst = 32'hc40439d;
      2284: inst = 32'h8220000;
      2285: inst = 32'h10408000;
      2286: inst = 32'hc40439e;
      2287: inst = 32'h8220000;
      2288: inst = 32'h10408000;
      2289: inst = 32'hc40439f;
      2290: inst = 32'h8220000;
      2291: inst = 32'h10408000;
      2292: inst = 32'hc4043a0;
      2293: inst = 32'h8220000;
      2294: inst = 32'h10408000;
      2295: inst = 32'hc4043a1;
      2296: inst = 32'h8220000;
      2297: inst = 32'h10408000;
      2298: inst = 32'hc4043a2;
      2299: inst = 32'h8220000;
      2300: inst = 32'h10408000;
      2301: inst = 32'hc4043a3;
      2302: inst = 32'h8220000;
      2303: inst = 32'h10408000;
      2304: inst = 32'hc4043a4;
      2305: inst = 32'h8220000;
      2306: inst = 32'h10408000;
      2307: inst = 32'hc4043a5;
      2308: inst = 32'h8220000;
      2309: inst = 32'h10408000;
      2310: inst = 32'hc4043a6;
      2311: inst = 32'h8220000;
      2312: inst = 32'h10408000;
      2313: inst = 32'hc4043b1;
      2314: inst = 32'h8220000;
      2315: inst = 32'h10408000;
      2316: inst = 32'hc4043b2;
      2317: inst = 32'h8220000;
      2318: inst = 32'h10408000;
      2319: inst = 32'hc4043b3;
      2320: inst = 32'h8220000;
      2321: inst = 32'h10408000;
      2322: inst = 32'hc4043b4;
      2323: inst = 32'h8220000;
      2324: inst = 32'h10408000;
      2325: inst = 32'hc4043b5;
      2326: inst = 32'h8220000;
      2327: inst = 32'h10408000;
      2328: inst = 32'hc4043b6;
      2329: inst = 32'h8220000;
      2330: inst = 32'h10408000;
      2331: inst = 32'hc4043b7;
      2332: inst = 32'h8220000;
      2333: inst = 32'h10408000;
      2334: inst = 32'hc4043b8;
      2335: inst = 32'h8220000;
      2336: inst = 32'h10408000;
      2337: inst = 32'hc4043b9;
      2338: inst = 32'h8220000;
      2339: inst = 32'h10408000;
      2340: inst = 32'hc4043ba;
      2341: inst = 32'h8220000;
      2342: inst = 32'h10408000;
      2343: inst = 32'hc4043bb;
      2344: inst = 32'h8220000;
      2345: inst = 32'h10408000;
      2346: inst = 32'hc4043e4;
      2347: inst = 32'h8220000;
      2348: inst = 32'h10408000;
      2349: inst = 32'hc4043e5;
      2350: inst = 32'h8220000;
      2351: inst = 32'h10408000;
      2352: inst = 32'hc4043e6;
      2353: inst = 32'h8220000;
      2354: inst = 32'h10408000;
      2355: inst = 32'hc4043e7;
      2356: inst = 32'h8220000;
      2357: inst = 32'h10408000;
      2358: inst = 32'hc4043e8;
      2359: inst = 32'h8220000;
      2360: inst = 32'h10408000;
      2361: inst = 32'hc4043e9;
      2362: inst = 32'h8220000;
      2363: inst = 32'h10408000;
      2364: inst = 32'hc4043ea;
      2365: inst = 32'h8220000;
      2366: inst = 32'h10408000;
      2367: inst = 32'hc4043eb;
      2368: inst = 32'h8220000;
      2369: inst = 32'h10408000;
      2370: inst = 32'hc4043ec;
      2371: inst = 32'h8220000;
      2372: inst = 32'h10408000;
      2373: inst = 32'hc4043ed;
      2374: inst = 32'h8220000;
      2375: inst = 32'h10408000;
      2376: inst = 32'hc4043ee;
      2377: inst = 32'h8220000;
      2378: inst = 32'h10408000;
      2379: inst = 32'hc4043ef;
      2380: inst = 32'h8220000;
      2381: inst = 32'h10408000;
      2382: inst = 32'hc4043f0;
      2383: inst = 32'h8220000;
      2384: inst = 32'h10408000;
      2385: inst = 32'hc4043f1;
      2386: inst = 32'h8220000;
      2387: inst = 32'h10408000;
      2388: inst = 32'hc4043f2;
      2389: inst = 32'h8220000;
      2390: inst = 32'h10408000;
      2391: inst = 32'hc4043f3;
      2392: inst = 32'h8220000;
      2393: inst = 32'h10408000;
      2394: inst = 32'hc4043f4;
      2395: inst = 32'h8220000;
      2396: inst = 32'h10408000;
      2397: inst = 32'hc4043f5;
      2398: inst = 32'h8220000;
      2399: inst = 32'h10408000;
      2400: inst = 32'hc4043f6;
      2401: inst = 32'h8220000;
      2402: inst = 32'h10408000;
      2403: inst = 32'hc4043f7;
      2404: inst = 32'h8220000;
      2405: inst = 32'h10408000;
      2406: inst = 32'hc4043f8;
      2407: inst = 32'h8220000;
      2408: inst = 32'h10408000;
      2409: inst = 32'hc4043f9;
      2410: inst = 32'h8220000;
      2411: inst = 32'h10408000;
      2412: inst = 32'hc4043fa;
      2413: inst = 32'h8220000;
      2414: inst = 32'h10408000;
      2415: inst = 32'hc4043fb;
      2416: inst = 32'h8220000;
      2417: inst = 32'h10408000;
      2418: inst = 32'hc4043fc;
      2419: inst = 32'h8220000;
      2420: inst = 32'h10408000;
      2421: inst = 32'hc4043fd;
      2422: inst = 32'h8220000;
      2423: inst = 32'h10408000;
      2424: inst = 32'hc4043fe;
      2425: inst = 32'h8220000;
      2426: inst = 32'h10408000;
      2427: inst = 32'hc4043ff;
      2428: inst = 32'h8220000;
      2429: inst = 32'h10408000;
      2430: inst = 32'hc404400;
      2431: inst = 32'h8220000;
      2432: inst = 32'h10408000;
      2433: inst = 32'hc404401;
      2434: inst = 32'h8220000;
      2435: inst = 32'h10408000;
      2436: inst = 32'hc404402;
      2437: inst = 32'h8220000;
      2438: inst = 32'h10408000;
      2439: inst = 32'hc404403;
      2440: inst = 32'h8220000;
      2441: inst = 32'h10408000;
      2442: inst = 32'hc404404;
      2443: inst = 32'h8220000;
      2444: inst = 32'h10408000;
      2445: inst = 32'hc404405;
      2446: inst = 32'h8220000;
      2447: inst = 32'h10408000;
      2448: inst = 32'hc404412;
      2449: inst = 32'h8220000;
      2450: inst = 32'h10408000;
      2451: inst = 32'hc404413;
      2452: inst = 32'h8220000;
      2453: inst = 32'h10408000;
      2454: inst = 32'hc404414;
      2455: inst = 32'h8220000;
      2456: inst = 32'h10408000;
      2457: inst = 32'hc404415;
      2458: inst = 32'h8220000;
      2459: inst = 32'h10408000;
      2460: inst = 32'hc404416;
      2461: inst = 32'h8220000;
      2462: inst = 32'h10408000;
      2463: inst = 32'hc404417;
      2464: inst = 32'h8220000;
      2465: inst = 32'h10408000;
      2466: inst = 32'hc404418;
      2467: inst = 32'h8220000;
      2468: inst = 32'h10408000;
      2469: inst = 32'hc404419;
      2470: inst = 32'h8220000;
      2471: inst = 32'h10408000;
      2472: inst = 32'hc40441a;
      2473: inst = 32'h8220000;
      2474: inst = 32'h10408000;
      2475: inst = 32'hc40441b;
      2476: inst = 32'h8220000;
      2477: inst = 32'h10408000;
      2478: inst = 32'hc404444;
      2479: inst = 32'h8220000;
      2480: inst = 32'h10408000;
      2481: inst = 32'hc404445;
      2482: inst = 32'h8220000;
      2483: inst = 32'h10408000;
      2484: inst = 32'hc404446;
      2485: inst = 32'h8220000;
      2486: inst = 32'h10408000;
      2487: inst = 32'hc404447;
      2488: inst = 32'h8220000;
      2489: inst = 32'h10408000;
      2490: inst = 32'hc404448;
      2491: inst = 32'h8220000;
      2492: inst = 32'h10408000;
      2493: inst = 32'hc404449;
      2494: inst = 32'h8220000;
      2495: inst = 32'h10408000;
      2496: inst = 32'hc40444a;
      2497: inst = 32'h8220000;
      2498: inst = 32'h10408000;
      2499: inst = 32'hc40444b;
      2500: inst = 32'h8220000;
      2501: inst = 32'h10408000;
      2502: inst = 32'hc40444c;
      2503: inst = 32'h8220000;
      2504: inst = 32'h10408000;
      2505: inst = 32'hc40444d;
      2506: inst = 32'h8220000;
      2507: inst = 32'h10408000;
      2508: inst = 32'hc40444e;
      2509: inst = 32'h8220000;
      2510: inst = 32'h10408000;
      2511: inst = 32'hc40444f;
      2512: inst = 32'h8220000;
      2513: inst = 32'h10408000;
      2514: inst = 32'hc404450;
      2515: inst = 32'h8220000;
      2516: inst = 32'h10408000;
      2517: inst = 32'hc404451;
      2518: inst = 32'h8220000;
      2519: inst = 32'h10408000;
      2520: inst = 32'hc404452;
      2521: inst = 32'h8220000;
      2522: inst = 32'h10408000;
      2523: inst = 32'hc404453;
      2524: inst = 32'h8220000;
      2525: inst = 32'h10408000;
      2526: inst = 32'hc404454;
      2527: inst = 32'h8220000;
      2528: inst = 32'h10408000;
      2529: inst = 32'hc404455;
      2530: inst = 32'h8220000;
      2531: inst = 32'h10408000;
      2532: inst = 32'hc404456;
      2533: inst = 32'h8220000;
      2534: inst = 32'h10408000;
      2535: inst = 32'hc404457;
      2536: inst = 32'h8220000;
      2537: inst = 32'h10408000;
      2538: inst = 32'hc404458;
      2539: inst = 32'h8220000;
      2540: inst = 32'h10408000;
      2541: inst = 32'hc404459;
      2542: inst = 32'h8220000;
      2543: inst = 32'h10408000;
      2544: inst = 32'hc40445a;
      2545: inst = 32'h8220000;
      2546: inst = 32'h10408000;
      2547: inst = 32'hc40445b;
      2548: inst = 32'h8220000;
      2549: inst = 32'h10408000;
      2550: inst = 32'hc40445c;
      2551: inst = 32'h8220000;
      2552: inst = 32'h10408000;
      2553: inst = 32'hc40445d;
      2554: inst = 32'h8220000;
      2555: inst = 32'h10408000;
      2556: inst = 32'hc40445e;
      2557: inst = 32'h8220000;
      2558: inst = 32'h10408000;
      2559: inst = 32'hc40445f;
      2560: inst = 32'h8220000;
      2561: inst = 32'h10408000;
      2562: inst = 32'hc404460;
      2563: inst = 32'h8220000;
      2564: inst = 32'h10408000;
      2565: inst = 32'hc404461;
      2566: inst = 32'h8220000;
      2567: inst = 32'h10408000;
      2568: inst = 32'hc404462;
      2569: inst = 32'h8220000;
      2570: inst = 32'h10408000;
      2571: inst = 32'hc404463;
      2572: inst = 32'h8220000;
      2573: inst = 32'h10408000;
      2574: inst = 32'hc404464;
      2575: inst = 32'h8220000;
      2576: inst = 32'h10408000;
      2577: inst = 32'hc404465;
      2578: inst = 32'h8220000;
      2579: inst = 32'h10408000;
      2580: inst = 32'hc404466;
      2581: inst = 32'h8220000;
      2582: inst = 32'h10408000;
      2583: inst = 32'hc404467;
      2584: inst = 32'h8220000;
      2585: inst = 32'h10408000;
      2586: inst = 32'hc404468;
      2587: inst = 32'h8220000;
      2588: inst = 32'h10408000;
      2589: inst = 32'hc404469;
      2590: inst = 32'h8220000;
      2591: inst = 32'h10408000;
      2592: inst = 32'hc40446e;
      2593: inst = 32'h8220000;
      2594: inst = 32'h10408000;
      2595: inst = 32'hc40446f;
      2596: inst = 32'h8220000;
      2597: inst = 32'h10408000;
      2598: inst = 32'hc404470;
      2599: inst = 32'h8220000;
      2600: inst = 32'h10408000;
      2601: inst = 32'hc404471;
      2602: inst = 32'h8220000;
      2603: inst = 32'h10408000;
      2604: inst = 32'hc404472;
      2605: inst = 32'h8220000;
      2606: inst = 32'h10408000;
      2607: inst = 32'hc404473;
      2608: inst = 32'h8220000;
      2609: inst = 32'h10408000;
      2610: inst = 32'hc404474;
      2611: inst = 32'h8220000;
      2612: inst = 32'h10408000;
      2613: inst = 32'hc404475;
      2614: inst = 32'h8220000;
      2615: inst = 32'h10408000;
      2616: inst = 32'hc404476;
      2617: inst = 32'h8220000;
      2618: inst = 32'h10408000;
      2619: inst = 32'hc404477;
      2620: inst = 32'h8220000;
      2621: inst = 32'h10408000;
      2622: inst = 32'hc404478;
      2623: inst = 32'h8220000;
      2624: inst = 32'h10408000;
      2625: inst = 32'hc404479;
      2626: inst = 32'h8220000;
      2627: inst = 32'h10408000;
      2628: inst = 32'hc40447a;
      2629: inst = 32'h8220000;
      2630: inst = 32'h10408000;
      2631: inst = 32'hc40447b;
      2632: inst = 32'h8220000;
      2633: inst = 32'h10408000;
      2634: inst = 32'hc4044a4;
      2635: inst = 32'h8220000;
      2636: inst = 32'h10408000;
      2637: inst = 32'hc4044a5;
      2638: inst = 32'h8220000;
      2639: inst = 32'h10408000;
      2640: inst = 32'hc4044a6;
      2641: inst = 32'h8220000;
      2642: inst = 32'h10408000;
      2643: inst = 32'hc4044a7;
      2644: inst = 32'h8220000;
      2645: inst = 32'h10408000;
      2646: inst = 32'hc4044a8;
      2647: inst = 32'h8220000;
      2648: inst = 32'h10408000;
      2649: inst = 32'hc4044a9;
      2650: inst = 32'h8220000;
      2651: inst = 32'h10408000;
      2652: inst = 32'hc4044aa;
      2653: inst = 32'h8220000;
      2654: inst = 32'h10408000;
      2655: inst = 32'hc4044ab;
      2656: inst = 32'h8220000;
      2657: inst = 32'h10408000;
      2658: inst = 32'hc4044ac;
      2659: inst = 32'h8220000;
      2660: inst = 32'h10408000;
      2661: inst = 32'hc4044ad;
      2662: inst = 32'h8220000;
      2663: inst = 32'h10408000;
      2664: inst = 32'hc4044ae;
      2665: inst = 32'h8220000;
      2666: inst = 32'h10408000;
      2667: inst = 32'hc4044af;
      2668: inst = 32'h8220000;
      2669: inst = 32'h10408000;
      2670: inst = 32'hc4044b0;
      2671: inst = 32'h8220000;
      2672: inst = 32'h10408000;
      2673: inst = 32'hc4044b1;
      2674: inst = 32'h8220000;
      2675: inst = 32'h10408000;
      2676: inst = 32'hc4044b6;
      2677: inst = 32'h8220000;
      2678: inst = 32'h10408000;
      2679: inst = 32'hc4044b7;
      2680: inst = 32'h8220000;
      2681: inst = 32'h10408000;
      2682: inst = 32'hc4044b8;
      2683: inst = 32'h8220000;
      2684: inst = 32'h10408000;
      2685: inst = 32'hc4044b9;
      2686: inst = 32'h8220000;
      2687: inst = 32'h10408000;
      2688: inst = 32'hc4044ba;
      2689: inst = 32'h8220000;
      2690: inst = 32'h10408000;
      2691: inst = 32'hc4044bb;
      2692: inst = 32'h8220000;
      2693: inst = 32'h10408000;
      2694: inst = 32'hc4044bc;
      2695: inst = 32'h8220000;
      2696: inst = 32'h10408000;
      2697: inst = 32'hc4044bd;
      2698: inst = 32'h8220000;
      2699: inst = 32'h10408000;
      2700: inst = 32'hc4044be;
      2701: inst = 32'h8220000;
      2702: inst = 32'h10408000;
      2703: inst = 32'hc4044bf;
      2704: inst = 32'h8220000;
      2705: inst = 32'h10408000;
      2706: inst = 32'hc4044c0;
      2707: inst = 32'h8220000;
      2708: inst = 32'h10408000;
      2709: inst = 32'hc4044c1;
      2710: inst = 32'h8220000;
      2711: inst = 32'h10408000;
      2712: inst = 32'hc4044c2;
      2713: inst = 32'h8220000;
      2714: inst = 32'h10408000;
      2715: inst = 32'hc4044c3;
      2716: inst = 32'h8220000;
      2717: inst = 32'h10408000;
      2718: inst = 32'hc4044c4;
      2719: inst = 32'h8220000;
      2720: inst = 32'h10408000;
      2721: inst = 32'hc4044c5;
      2722: inst = 32'h8220000;
      2723: inst = 32'h10408000;
      2724: inst = 32'hc4044c6;
      2725: inst = 32'h8220000;
      2726: inst = 32'h10408000;
      2727: inst = 32'hc4044c7;
      2728: inst = 32'h8220000;
      2729: inst = 32'h10408000;
      2730: inst = 32'hc4044c8;
      2731: inst = 32'h8220000;
      2732: inst = 32'h10408000;
      2733: inst = 32'hc4044c9;
      2734: inst = 32'h8220000;
      2735: inst = 32'h10408000;
      2736: inst = 32'hc4044ca;
      2737: inst = 32'h8220000;
      2738: inst = 32'h10408000;
      2739: inst = 32'hc4044cd;
      2740: inst = 32'h8220000;
      2741: inst = 32'h10408000;
      2742: inst = 32'hc4044ce;
      2743: inst = 32'h8220000;
      2744: inst = 32'h10408000;
      2745: inst = 32'hc4044cf;
      2746: inst = 32'h8220000;
      2747: inst = 32'h10408000;
      2748: inst = 32'hc4044d0;
      2749: inst = 32'h8220000;
      2750: inst = 32'h10408000;
      2751: inst = 32'hc4044d1;
      2752: inst = 32'h8220000;
      2753: inst = 32'h10408000;
      2754: inst = 32'hc4044d2;
      2755: inst = 32'h8220000;
      2756: inst = 32'h10408000;
      2757: inst = 32'hc4044d3;
      2758: inst = 32'h8220000;
      2759: inst = 32'h10408000;
      2760: inst = 32'hc4044d4;
      2761: inst = 32'h8220000;
      2762: inst = 32'h10408000;
      2763: inst = 32'hc4044d5;
      2764: inst = 32'h8220000;
      2765: inst = 32'h10408000;
      2766: inst = 32'hc4044d6;
      2767: inst = 32'h8220000;
      2768: inst = 32'h10408000;
      2769: inst = 32'hc4044d7;
      2770: inst = 32'h8220000;
      2771: inst = 32'h10408000;
      2772: inst = 32'hc4044d8;
      2773: inst = 32'h8220000;
      2774: inst = 32'h10408000;
      2775: inst = 32'hc4044d9;
      2776: inst = 32'h8220000;
      2777: inst = 32'h10408000;
      2778: inst = 32'hc4044da;
      2779: inst = 32'h8220000;
      2780: inst = 32'h10408000;
      2781: inst = 32'hc4044db;
      2782: inst = 32'h8220000;
      2783: inst = 32'h10408000;
      2784: inst = 32'hc404504;
      2785: inst = 32'h8220000;
      2786: inst = 32'h10408000;
      2787: inst = 32'hc404505;
      2788: inst = 32'h8220000;
      2789: inst = 32'h10408000;
      2790: inst = 32'hc404506;
      2791: inst = 32'h8220000;
      2792: inst = 32'h10408000;
      2793: inst = 32'hc404507;
      2794: inst = 32'h8220000;
      2795: inst = 32'h10408000;
      2796: inst = 32'hc404508;
      2797: inst = 32'h8220000;
      2798: inst = 32'h10408000;
      2799: inst = 32'hc404509;
      2800: inst = 32'h8220000;
      2801: inst = 32'h10408000;
      2802: inst = 32'hc40450a;
      2803: inst = 32'h8220000;
      2804: inst = 32'h10408000;
      2805: inst = 32'hc40450b;
      2806: inst = 32'h8220000;
      2807: inst = 32'h10408000;
      2808: inst = 32'hc40450c;
      2809: inst = 32'h8220000;
      2810: inst = 32'h10408000;
      2811: inst = 32'hc40450d;
      2812: inst = 32'h8220000;
      2813: inst = 32'h10408000;
      2814: inst = 32'hc40450e;
      2815: inst = 32'h8220000;
      2816: inst = 32'h10408000;
      2817: inst = 32'hc40450f;
      2818: inst = 32'h8220000;
      2819: inst = 32'h10408000;
      2820: inst = 32'hc404510;
      2821: inst = 32'h8220000;
      2822: inst = 32'h10408000;
      2823: inst = 32'hc404511;
      2824: inst = 32'h8220000;
      2825: inst = 32'h10408000;
      2826: inst = 32'hc404512;
      2827: inst = 32'h8220000;
      2828: inst = 32'h10408000;
      2829: inst = 32'hc404515;
      2830: inst = 32'h8220000;
      2831: inst = 32'h10408000;
      2832: inst = 32'hc404516;
      2833: inst = 32'h8220000;
      2834: inst = 32'h10408000;
      2835: inst = 32'hc404517;
      2836: inst = 32'h8220000;
      2837: inst = 32'h10408000;
      2838: inst = 32'hc404518;
      2839: inst = 32'h8220000;
      2840: inst = 32'h10408000;
      2841: inst = 32'hc404519;
      2842: inst = 32'h8220000;
      2843: inst = 32'h10408000;
      2844: inst = 32'hc40451a;
      2845: inst = 32'h8220000;
      2846: inst = 32'h10408000;
      2847: inst = 32'hc40451b;
      2848: inst = 32'h8220000;
      2849: inst = 32'h10408000;
      2850: inst = 32'hc40451c;
      2851: inst = 32'h8220000;
      2852: inst = 32'h10408000;
      2853: inst = 32'hc40451d;
      2854: inst = 32'h8220000;
      2855: inst = 32'h10408000;
      2856: inst = 32'hc40451e;
      2857: inst = 32'h8220000;
      2858: inst = 32'h10408000;
      2859: inst = 32'hc40451f;
      2860: inst = 32'h8220000;
      2861: inst = 32'h10408000;
      2862: inst = 32'hc404520;
      2863: inst = 32'h8220000;
      2864: inst = 32'h10408000;
      2865: inst = 32'hc404521;
      2866: inst = 32'h8220000;
      2867: inst = 32'h10408000;
      2868: inst = 32'hc404522;
      2869: inst = 32'h8220000;
      2870: inst = 32'h10408000;
      2871: inst = 32'hc404523;
      2872: inst = 32'h8220000;
      2873: inst = 32'h10408000;
      2874: inst = 32'hc404524;
      2875: inst = 32'h8220000;
      2876: inst = 32'h10408000;
      2877: inst = 32'hc404525;
      2878: inst = 32'h8220000;
      2879: inst = 32'h10408000;
      2880: inst = 32'hc404526;
      2881: inst = 32'h8220000;
      2882: inst = 32'h10408000;
      2883: inst = 32'hc404527;
      2884: inst = 32'h8220000;
      2885: inst = 32'h10408000;
      2886: inst = 32'hc404528;
      2887: inst = 32'h8220000;
      2888: inst = 32'h10408000;
      2889: inst = 32'hc404529;
      2890: inst = 32'h8220000;
      2891: inst = 32'h10408000;
      2892: inst = 32'hc40452a;
      2893: inst = 32'h8220000;
      2894: inst = 32'h10408000;
      2895: inst = 32'hc40452b;
      2896: inst = 32'h8220000;
      2897: inst = 32'h10408000;
      2898: inst = 32'hc40452c;
      2899: inst = 32'h8220000;
      2900: inst = 32'h10408000;
      2901: inst = 32'hc40452d;
      2902: inst = 32'h8220000;
      2903: inst = 32'h10408000;
      2904: inst = 32'hc40452e;
      2905: inst = 32'h8220000;
      2906: inst = 32'h10408000;
      2907: inst = 32'hc40452f;
      2908: inst = 32'h8220000;
      2909: inst = 32'h10408000;
      2910: inst = 32'hc404530;
      2911: inst = 32'h8220000;
      2912: inst = 32'h10408000;
      2913: inst = 32'hc404531;
      2914: inst = 32'h8220000;
      2915: inst = 32'h10408000;
      2916: inst = 32'hc404532;
      2917: inst = 32'h8220000;
      2918: inst = 32'h10408000;
      2919: inst = 32'hc404533;
      2920: inst = 32'h8220000;
      2921: inst = 32'h10408000;
      2922: inst = 32'hc404534;
      2923: inst = 32'h8220000;
      2924: inst = 32'h10408000;
      2925: inst = 32'hc404535;
      2926: inst = 32'h8220000;
      2927: inst = 32'h10408000;
      2928: inst = 32'hc404536;
      2929: inst = 32'h8220000;
      2930: inst = 32'h10408000;
      2931: inst = 32'hc404537;
      2932: inst = 32'h8220000;
      2933: inst = 32'h10408000;
      2934: inst = 32'hc404538;
      2935: inst = 32'h8220000;
      2936: inst = 32'h10408000;
      2937: inst = 32'hc404539;
      2938: inst = 32'h8220000;
      2939: inst = 32'h10408000;
      2940: inst = 32'hc40453a;
      2941: inst = 32'h8220000;
      2942: inst = 32'h10408000;
      2943: inst = 32'hc40453b;
      2944: inst = 32'h8220000;
      2945: inst = 32'h10408000;
      2946: inst = 32'hc404564;
      2947: inst = 32'h8220000;
      2948: inst = 32'h10408000;
      2949: inst = 32'hc404565;
      2950: inst = 32'h8220000;
      2951: inst = 32'h10408000;
      2952: inst = 32'hc404566;
      2953: inst = 32'h8220000;
      2954: inst = 32'h10408000;
      2955: inst = 32'hc404567;
      2956: inst = 32'h8220000;
      2957: inst = 32'h10408000;
      2958: inst = 32'hc404568;
      2959: inst = 32'h8220000;
      2960: inst = 32'h10408000;
      2961: inst = 32'hc404569;
      2962: inst = 32'h8220000;
      2963: inst = 32'h10408000;
      2964: inst = 32'hc40456a;
      2965: inst = 32'h8220000;
      2966: inst = 32'h10408000;
      2967: inst = 32'hc40456b;
      2968: inst = 32'h8220000;
      2969: inst = 32'h10408000;
      2970: inst = 32'hc40456c;
      2971: inst = 32'h8220000;
      2972: inst = 32'h10408000;
      2973: inst = 32'hc40456d;
      2974: inst = 32'h8220000;
      2975: inst = 32'h10408000;
      2976: inst = 32'hc40456e;
      2977: inst = 32'h8220000;
      2978: inst = 32'h10408000;
      2979: inst = 32'hc40456f;
      2980: inst = 32'h8220000;
      2981: inst = 32'h10408000;
      2982: inst = 32'hc404570;
      2983: inst = 32'h8220000;
      2984: inst = 32'h10408000;
      2985: inst = 32'hc404571;
      2986: inst = 32'h8220000;
      2987: inst = 32'h10408000;
      2988: inst = 32'hc404572;
      2989: inst = 32'h8220000;
      2990: inst = 32'h10408000;
      2991: inst = 32'hc404573;
      2992: inst = 32'h8220000;
      2993: inst = 32'h10408000;
      2994: inst = 32'hc404574;
      2995: inst = 32'h8220000;
      2996: inst = 32'h10408000;
      2997: inst = 32'hc404575;
      2998: inst = 32'h8220000;
      2999: inst = 32'h10408000;
      3000: inst = 32'hc404576;
      3001: inst = 32'h8220000;
      3002: inst = 32'h10408000;
      3003: inst = 32'hc404577;
      3004: inst = 32'h8220000;
      3005: inst = 32'h10408000;
      3006: inst = 32'hc404578;
      3007: inst = 32'h8220000;
      3008: inst = 32'h10408000;
      3009: inst = 32'hc404579;
      3010: inst = 32'h8220000;
      3011: inst = 32'h10408000;
      3012: inst = 32'hc40457a;
      3013: inst = 32'h8220000;
      3014: inst = 32'h10408000;
      3015: inst = 32'hc40457b;
      3016: inst = 32'h8220000;
      3017: inst = 32'h10408000;
      3018: inst = 32'hc40457c;
      3019: inst = 32'h8220000;
      3020: inst = 32'h10408000;
      3021: inst = 32'hc40457d;
      3022: inst = 32'h8220000;
      3023: inst = 32'h10408000;
      3024: inst = 32'hc40457e;
      3025: inst = 32'h8220000;
      3026: inst = 32'h10408000;
      3027: inst = 32'hc40457f;
      3028: inst = 32'h8220000;
      3029: inst = 32'h10408000;
      3030: inst = 32'hc404580;
      3031: inst = 32'h8220000;
      3032: inst = 32'h10408000;
      3033: inst = 32'hc404581;
      3034: inst = 32'h8220000;
      3035: inst = 32'h10408000;
      3036: inst = 32'hc404582;
      3037: inst = 32'h8220000;
      3038: inst = 32'h10408000;
      3039: inst = 32'hc404583;
      3040: inst = 32'h8220000;
      3041: inst = 32'h10408000;
      3042: inst = 32'hc404584;
      3043: inst = 32'h8220000;
      3044: inst = 32'h10408000;
      3045: inst = 32'hc404585;
      3046: inst = 32'h8220000;
      3047: inst = 32'h10408000;
      3048: inst = 32'hc404586;
      3049: inst = 32'h8220000;
      3050: inst = 32'h10408000;
      3051: inst = 32'hc404587;
      3052: inst = 32'h8220000;
      3053: inst = 32'h10408000;
      3054: inst = 32'hc404588;
      3055: inst = 32'h8220000;
      3056: inst = 32'h10408000;
      3057: inst = 32'hc404589;
      3058: inst = 32'h8220000;
      3059: inst = 32'h10408000;
      3060: inst = 32'hc40458a;
      3061: inst = 32'h8220000;
      3062: inst = 32'h10408000;
      3063: inst = 32'hc40458b;
      3064: inst = 32'h8220000;
      3065: inst = 32'h10408000;
      3066: inst = 32'hc40458c;
      3067: inst = 32'h8220000;
      3068: inst = 32'h10408000;
      3069: inst = 32'hc40458d;
      3070: inst = 32'h8220000;
      3071: inst = 32'h10408000;
      3072: inst = 32'hc40458e;
      3073: inst = 32'h8220000;
      3074: inst = 32'h10408000;
      3075: inst = 32'hc40458f;
      3076: inst = 32'h8220000;
      3077: inst = 32'h10408000;
      3078: inst = 32'hc404590;
      3079: inst = 32'h8220000;
      3080: inst = 32'h10408000;
      3081: inst = 32'hc404591;
      3082: inst = 32'h8220000;
      3083: inst = 32'h10408000;
      3084: inst = 32'hc404592;
      3085: inst = 32'h8220000;
      3086: inst = 32'h10408000;
      3087: inst = 32'hc404593;
      3088: inst = 32'h8220000;
      3089: inst = 32'h10408000;
      3090: inst = 32'hc404594;
      3091: inst = 32'h8220000;
      3092: inst = 32'h10408000;
      3093: inst = 32'hc404595;
      3094: inst = 32'h8220000;
      3095: inst = 32'h10408000;
      3096: inst = 32'hc404596;
      3097: inst = 32'h8220000;
      3098: inst = 32'h10408000;
      3099: inst = 32'hc404597;
      3100: inst = 32'h8220000;
      3101: inst = 32'h10408000;
      3102: inst = 32'hc404598;
      3103: inst = 32'h8220000;
      3104: inst = 32'h10408000;
      3105: inst = 32'hc404599;
      3106: inst = 32'h8220000;
      3107: inst = 32'h10408000;
      3108: inst = 32'hc40459a;
      3109: inst = 32'h8220000;
      3110: inst = 32'h10408000;
      3111: inst = 32'hc40459b;
      3112: inst = 32'h8220000;
      3113: inst = 32'h10408000;
      3114: inst = 32'hc4045c4;
      3115: inst = 32'h8220000;
      3116: inst = 32'h10408000;
      3117: inst = 32'hc4045c5;
      3118: inst = 32'h8220000;
      3119: inst = 32'h10408000;
      3120: inst = 32'hc4045c6;
      3121: inst = 32'h8220000;
      3122: inst = 32'h10408000;
      3123: inst = 32'hc4045c7;
      3124: inst = 32'h8220000;
      3125: inst = 32'h10408000;
      3126: inst = 32'hc4045c8;
      3127: inst = 32'h8220000;
      3128: inst = 32'h10408000;
      3129: inst = 32'hc4045c9;
      3130: inst = 32'h8220000;
      3131: inst = 32'h10408000;
      3132: inst = 32'hc4045ca;
      3133: inst = 32'h8220000;
      3134: inst = 32'h10408000;
      3135: inst = 32'hc4045cb;
      3136: inst = 32'h8220000;
      3137: inst = 32'h10408000;
      3138: inst = 32'hc4045cc;
      3139: inst = 32'h8220000;
      3140: inst = 32'h10408000;
      3141: inst = 32'hc4045cd;
      3142: inst = 32'h8220000;
      3143: inst = 32'h10408000;
      3144: inst = 32'hc4045ce;
      3145: inst = 32'h8220000;
      3146: inst = 32'h10408000;
      3147: inst = 32'hc4045cf;
      3148: inst = 32'h8220000;
      3149: inst = 32'h10408000;
      3150: inst = 32'hc4045d0;
      3151: inst = 32'h8220000;
      3152: inst = 32'h10408000;
      3153: inst = 32'hc4045d1;
      3154: inst = 32'h8220000;
      3155: inst = 32'h10408000;
      3156: inst = 32'hc4045d2;
      3157: inst = 32'h8220000;
      3158: inst = 32'h10408000;
      3159: inst = 32'hc4045d3;
      3160: inst = 32'h8220000;
      3161: inst = 32'h10408000;
      3162: inst = 32'hc4045d4;
      3163: inst = 32'h8220000;
      3164: inst = 32'h10408000;
      3165: inst = 32'hc4045d5;
      3166: inst = 32'h8220000;
      3167: inst = 32'h10408000;
      3168: inst = 32'hc4045d6;
      3169: inst = 32'h8220000;
      3170: inst = 32'h10408000;
      3171: inst = 32'hc4045d7;
      3172: inst = 32'h8220000;
      3173: inst = 32'h10408000;
      3174: inst = 32'hc4045d8;
      3175: inst = 32'h8220000;
      3176: inst = 32'h10408000;
      3177: inst = 32'hc4045d9;
      3178: inst = 32'h8220000;
      3179: inst = 32'h10408000;
      3180: inst = 32'hc4045da;
      3181: inst = 32'h8220000;
      3182: inst = 32'h10408000;
      3183: inst = 32'hc4045db;
      3184: inst = 32'h8220000;
      3185: inst = 32'h10408000;
      3186: inst = 32'hc4045dc;
      3187: inst = 32'h8220000;
      3188: inst = 32'h10408000;
      3189: inst = 32'hc4045dd;
      3190: inst = 32'h8220000;
      3191: inst = 32'h10408000;
      3192: inst = 32'hc4045de;
      3193: inst = 32'h8220000;
      3194: inst = 32'h10408000;
      3195: inst = 32'hc4045df;
      3196: inst = 32'h8220000;
      3197: inst = 32'h10408000;
      3198: inst = 32'hc4045e0;
      3199: inst = 32'h8220000;
      3200: inst = 32'h10408000;
      3201: inst = 32'hc4045e1;
      3202: inst = 32'h8220000;
      3203: inst = 32'h10408000;
      3204: inst = 32'hc4045e2;
      3205: inst = 32'h8220000;
      3206: inst = 32'h10408000;
      3207: inst = 32'hc4045e3;
      3208: inst = 32'h8220000;
      3209: inst = 32'h10408000;
      3210: inst = 32'hc4045e4;
      3211: inst = 32'h8220000;
      3212: inst = 32'h10408000;
      3213: inst = 32'hc4045e5;
      3214: inst = 32'h8220000;
      3215: inst = 32'h10408000;
      3216: inst = 32'hc4045e6;
      3217: inst = 32'h8220000;
      3218: inst = 32'h10408000;
      3219: inst = 32'hc4045e7;
      3220: inst = 32'h8220000;
      3221: inst = 32'h10408000;
      3222: inst = 32'hc4045e8;
      3223: inst = 32'h8220000;
      3224: inst = 32'h10408000;
      3225: inst = 32'hc4045e9;
      3226: inst = 32'h8220000;
      3227: inst = 32'h10408000;
      3228: inst = 32'hc4045ea;
      3229: inst = 32'h8220000;
      3230: inst = 32'h10408000;
      3231: inst = 32'hc4045eb;
      3232: inst = 32'h8220000;
      3233: inst = 32'h10408000;
      3234: inst = 32'hc4045ec;
      3235: inst = 32'h8220000;
      3236: inst = 32'h10408000;
      3237: inst = 32'hc4045ed;
      3238: inst = 32'h8220000;
      3239: inst = 32'h10408000;
      3240: inst = 32'hc4045ee;
      3241: inst = 32'h8220000;
      3242: inst = 32'h10408000;
      3243: inst = 32'hc4045ef;
      3244: inst = 32'h8220000;
      3245: inst = 32'h10408000;
      3246: inst = 32'hc4045f0;
      3247: inst = 32'h8220000;
      3248: inst = 32'h10408000;
      3249: inst = 32'hc4045f1;
      3250: inst = 32'h8220000;
      3251: inst = 32'h10408000;
      3252: inst = 32'hc4045f2;
      3253: inst = 32'h8220000;
      3254: inst = 32'h10408000;
      3255: inst = 32'hc4045f3;
      3256: inst = 32'h8220000;
      3257: inst = 32'h10408000;
      3258: inst = 32'hc4045f4;
      3259: inst = 32'h8220000;
      3260: inst = 32'h10408000;
      3261: inst = 32'hc4045f5;
      3262: inst = 32'h8220000;
      3263: inst = 32'h10408000;
      3264: inst = 32'hc4045f6;
      3265: inst = 32'h8220000;
      3266: inst = 32'h10408000;
      3267: inst = 32'hc4045f7;
      3268: inst = 32'h8220000;
      3269: inst = 32'h10408000;
      3270: inst = 32'hc4045f8;
      3271: inst = 32'h8220000;
      3272: inst = 32'h10408000;
      3273: inst = 32'hc4045f9;
      3274: inst = 32'h8220000;
      3275: inst = 32'h10408000;
      3276: inst = 32'hc4045fa;
      3277: inst = 32'h8220000;
      3278: inst = 32'h10408000;
      3279: inst = 32'hc4045fb;
      3280: inst = 32'h8220000;
      3281: inst = 32'h10408000;
      3282: inst = 32'hc404624;
      3283: inst = 32'h8220000;
      3284: inst = 32'h10408000;
      3285: inst = 32'hc404625;
      3286: inst = 32'h8220000;
      3287: inst = 32'h10408000;
      3288: inst = 32'hc404626;
      3289: inst = 32'h8220000;
      3290: inst = 32'h10408000;
      3291: inst = 32'hc404627;
      3292: inst = 32'h8220000;
      3293: inst = 32'h10408000;
      3294: inst = 32'hc404628;
      3295: inst = 32'h8220000;
      3296: inst = 32'h10408000;
      3297: inst = 32'hc404629;
      3298: inst = 32'h8220000;
      3299: inst = 32'h10408000;
      3300: inst = 32'hc40462a;
      3301: inst = 32'h8220000;
      3302: inst = 32'h10408000;
      3303: inst = 32'hc40462b;
      3304: inst = 32'h8220000;
      3305: inst = 32'h10408000;
      3306: inst = 32'hc40462c;
      3307: inst = 32'h8220000;
      3308: inst = 32'h10408000;
      3309: inst = 32'hc40462d;
      3310: inst = 32'h8220000;
      3311: inst = 32'h10408000;
      3312: inst = 32'hc40462e;
      3313: inst = 32'h8220000;
      3314: inst = 32'h10408000;
      3315: inst = 32'hc40462f;
      3316: inst = 32'h8220000;
      3317: inst = 32'h10408000;
      3318: inst = 32'hc404630;
      3319: inst = 32'h8220000;
      3320: inst = 32'h10408000;
      3321: inst = 32'hc404631;
      3322: inst = 32'h8220000;
      3323: inst = 32'h10408000;
      3324: inst = 32'hc404632;
      3325: inst = 32'h8220000;
      3326: inst = 32'h10408000;
      3327: inst = 32'hc404633;
      3328: inst = 32'h8220000;
      3329: inst = 32'h10408000;
      3330: inst = 32'hc404634;
      3331: inst = 32'h8220000;
      3332: inst = 32'h10408000;
      3333: inst = 32'hc404635;
      3334: inst = 32'h8220000;
      3335: inst = 32'h10408000;
      3336: inst = 32'hc404636;
      3337: inst = 32'h8220000;
      3338: inst = 32'h10408000;
      3339: inst = 32'hc404637;
      3340: inst = 32'h8220000;
      3341: inst = 32'h10408000;
      3342: inst = 32'hc404638;
      3343: inst = 32'h8220000;
      3344: inst = 32'h10408000;
      3345: inst = 32'hc404639;
      3346: inst = 32'h8220000;
      3347: inst = 32'h10408000;
      3348: inst = 32'hc40463a;
      3349: inst = 32'h8220000;
      3350: inst = 32'h10408000;
      3351: inst = 32'hc40463b;
      3352: inst = 32'h8220000;
      3353: inst = 32'h10408000;
      3354: inst = 32'hc40463c;
      3355: inst = 32'h8220000;
      3356: inst = 32'h10408000;
      3357: inst = 32'hc40463d;
      3358: inst = 32'h8220000;
      3359: inst = 32'h10408000;
      3360: inst = 32'hc40463e;
      3361: inst = 32'h8220000;
      3362: inst = 32'h10408000;
      3363: inst = 32'hc40463f;
      3364: inst = 32'h8220000;
      3365: inst = 32'h10408000;
      3366: inst = 32'hc404640;
      3367: inst = 32'h8220000;
      3368: inst = 32'h10408000;
      3369: inst = 32'hc404641;
      3370: inst = 32'h8220000;
      3371: inst = 32'h10408000;
      3372: inst = 32'hc404642;
      3373: inst = 32'h8220000;
      3374: inst = 32'h10408000;
      3375: inst = 32'hc404643;
      3376: inst = 32'h8220000;
      3377: inst = 32'h10408000;
      3378: inst = 32'hc404644;
      3379: inst = 32'h8220000;
      3380: inst = 32'h10408000;
      3381: inst = 32'hc404645;
      3382: inst = 32'h8220000;
      3383: inst = 32'h10408000;
      3384: inst = 32'hc404646;
      3385: inst = 32'h8220000;
      3386: inst = 32'h10408000;
      3387: inst = 32'hc404647;
      3388: inst = 32'h8220000;
      3389: inst = 32'h10408000;
      3390: inst = 32'hc404648;
      3391: inst = 32'h8220000;
      3392: inst = 32'h10408000;
      3393: inst = 32'hc404649;
      3394: inst = 32'h8220000;
      3395: inst = 32'h10408000;
      3396: inst = 32'hc40464a;
      3397: inst = 32'h8220000;
      3398: inst = 32'h10408000;
      3399: inst = 32'hc40464b;
      3400: inst = 32'h8220000;
      3401: inst = 32'h10408000;
      3402: inst = 32'hc40464c;
      3403: inst = 32'h8220000;
      3404: inst = 32'h10408000;
      3405: inst = 32'hc40464d;
      3406: inst = 32'h8220000;
      3407: inst = 32'h10408000;
      3408: inst = 32'hc40464e;
      3409: inst = 32'h8220000;
      3410: inst = 32'h10408000;
      3411: inst = 32'hc40464f;
      3412: inst = 32'h8220000;
      3413: inst = 32'h10408000;
      3414: inst = 32'hc404650;
      3415: inst = 32'h8220000;
      3416: inst = 32'h10408000;
      3417: inst = 32'hc404651;
      3418: inst = 32'h8220000;
      3419: inst = 32'h10408000;
      3420: inst = 32'hc404652;
      3421: inst = 32'h8220000;
      3422: inst = 32'h10408000;
      3423: inst = 32'hc404653;
      3424: inst = 32'h8220000;
      3425: inst = 32'h10408000;
      3426: inst = 32'hc404654;
      3427: inst = 32'h8220000;
      3428: inst = 32'h10408000;
      3429: inst = 32'hc404655;
      3430: inst = 32'h8220000;
      3431: inst = 32'h10408000;
      3432: inst = 32'hc404656;
      3433: inst = 32'h8220000;
      3434: inst = 32'h10408000;
      3435: inst = 32'hc404657;
      3436: inst = 32'h8220000;
      3437: inst = 32'h10408000;
      3438: inst = 32'hc404658;
      3439: inst = 32'h8220000;
      3440: inst = 32'h10408000;
      3441: inst = 32'hc404659;
      3442: inst = 32'h8220000;
      3443: inst = 32'h10408000;
      3444: inst = 32'hc40465a;
      3445: inst = 32'h8220000;
      3446: inst = 32'h10408000;
      3447: inst = 32'hc40465b;
      3448: inst = 32'h8220000;
      3449: inst = 32'h10408000;
      3450: inst = 32'hc404684;
      3451: inst = 32'h8220000;
      3452: inst = 32'h10408000;
      3453: inst = 32'hc404685;
      3454: inst = 32'h8220000;
      3455: inst = 32'h10408000;
      3456: inst = 32'hc404686;
      3457: inst = 32'h8220000;
      3458: inst = 32'h10408000;
      3459: inst = 32'hc404687;
      3460: inst = 32'h8220000;
      3461: inst = 32'h10408000;
      3462: inst = 32'hc404688;
      3463: inst = 32'h8220000;
      3464: inst = 32'h10408000;
      3465: inst = 32'hc404689;
      3466: inst = 32'h8220000;
      3467: inst = 32'h10408000;
      3468: inst = 32'hc40468a;
      3469: inst = 32'h8220000;
      3470: inst = 32'h10408000;
      3471: inst = 32'hc40468b;
      3472: inst = 32'h8220000;
      3473: inst = 32'h10408000;
      3474: inst = 32'hc40468c;
      3475: inst = 32'h8220000;
      3476: inst = 32'h10408000;
      3477: inst = 32'hc40468d;
      3478: inst = 32'h8220000;
      3479: inst = 32'h10408000;
      3480: inst = 32'hc40468e;
      3481: inst = 32'h8220000;
      3482: inst = 32'h10408000;
      3483: inst = 32'hc40468f;
      3484: inst = 32'h8220000;
      3485: inst = 32'h10408000;
      3486: inst = 32'hc404690;
      3487: inst = 32'h8220000;
      3488: inst = 32'h10408000;
      3489: inst = 32'hc404691;
      3490: inst = 32'h8220000;
      3491: inst = 32'h10408000;
      3492: inst = 32'hc404692;
      3493: inst = 32'h8220000;
      3494: inst = 32'h10408000;
      3495: inst = 32'hc404693;
      3496: inst = 32'h8220000;
      3497: inst = 32'h10408000;
      3498: inst = 32'hc404694;
      3499: inst = 32'h8220000;
      3500: inst = 32'h10408000;
      3501: inst = 32'hc404695;
      3502: inst = 32'h8220000;
      3503: inst = 32'h10408000;
      3504: inst = 32'hc404696;
      3505: inst = 32'h8220000;
      3506: inst = 32'h10408000;
      3507: inst = 32'hc404697;
      3508: inst = 32'h8220000;
      3509: inst = 32'h10408000;
      3510: inst = 32'hc404698;
      3511: inst = 32'h8220000;
      3512: inst = 32'h10408000;
      3513: inst = 32'hc404699;
      3514: inst = 32'h8220000;
      3515: inst = 32'h10408000;
      3516: inst = 32'hc40469a;
      3517: inst = 32'h8220000;
      3518: inst = 32'h10408000;
      3519: inst = 32'hc40469b;
      3520: inst = 32'h8220000;
      3521: inst = 32'h10408000;
      3522: inst = 32'hc40469c;
      3523: inst = 32'h8220000;
      3524: inst = 32'h10408000;
      3525: inst = 32'hc40469d;
      3526: inst = 32'h8220000;
      3527: inst = 32'h10408000;
      3528: inst = 32'hc40469e;
      3529: inst = 32'h8220000;
      3530: inst = 32'h10408000;
      3531: inst = 32'hc40469f;
      3532: inst = 32'h8220000;
      3533: inst = 32'h10408000;
      3534: inst = 32'hc4046a0;
      3535: inst = 32'h8220000;
      3536: inst = 32'h10408000;
      3537: inst = 32'hc4046a1;
      3538: inst = 32'h8220000;
      3539: inst = 32'h10408000;
      3540: inst = 32'hc4046a2;
      3541: inst = 32'h8220000;
      3542: inst = 32'h10408000;
      3543: inst = 32'hc4046a3;
      3544: inst = 32'h8220000;
      3545: inst = 32'h10408000;
      3546: inst = 32'hc4046a4;
      3547: inst = 32'h8220000;
      3548: inst = 32'h10408000;
      3549: inst = 32'hc4046a5;
      3550: inst = 32'h8220000;
      3551: inst = 32'h10408000;
      3552: inst = 32'hc4046a6;
      3553: inst = 32'h8220000;
      3554: inst = 32'h10408000;
      3555: inst = 32'hc4046a7;
      3556: inst = 32'h8220000;
      3557: inst = 32'h10408000;
      3558: inst = 32'hc4046a8;
      3559: inst = 32'h8220000;
      3560: inst = 32'h10408000;
      3561: inst = 32'hc4046a9;
      3562: inst = 32'h8220000;
      3563: inst = 32'h10408000;
      3564: inst = 32'hc4046aa;
      3565: inst = 32'h8220000;
      3566: inst = 32'h10408000;
      3567: inst = 32'hc4046ab;
      3568: inst = 32'h8220000;
      3569: inst = 32'h10408000;
      3570: inst = 32'hc4046ac;
      3571: inst = 32'h8220000;
      3572: inst = 32'h10408000;
      3573: inst = 32'hc4046ad;
      3574: inst = 32'h8220000;
      3575: inst = 32'h10408000;
      3576: inst = 32'hc4046ae;
      3577: inst = 32'h8220000;
      3578: inst = 32'h10408000;
      3579: inst = 32'hc4046af;
      3580: inst = 32'h8220000;
      3581: inst = 32'h10408000;
      3582: inst = 32'hc4046b0;
      3583: inst = 32'h8220000;
      3584: inst = 32'h10408000;
      3585: inst = 32'hc4046b1;
      3586: inst = 32'h8220000;
      3587: inst = 32'h10408000;
      3588: inst = 32'hc4046b2;
      3589: inst = 32'h8220000;
      3590: inst = 32'h10408000;
      3591: inst = 32'hc4046b3;
      3592: inst = 32'h8220000;
      3593: inst = 32'h10408000;
      3594: inst = 32'hc4046b4;
      3595: inst = 32'h8220000;
      3596: inst = 32'h10408000;
      3597: inst = 32'hc4046b5;
      3598: inst = 32'h8220000;
      3599: inst = 32'h10408000;
      3600: inst = 32'hc4046b6;
      3601: inst = 32'h8220000;
      3602: inst = 32'h10408000;
      3603: inst = 32'hc4046b7;
      3604: inst = 32'h8220000;
      3605: inst = 32'h10408000;
      3606: inst = 32'hc4046b8;
      3607: inst = 32'h8220000;
      3608: inst = 32'h10408000;
      3609: inst = 32'hc4046b9;
      3610: inst = 32'h8220000;
      3611: inst = 32'h10408000;
      3612: inst = 32'hc4046ba;
      3613: inst = 32'h8220000;
      3614: inst = 32'h10408000;
      3615: inst = 32'hc4046bb;
      3616: inst = 32'h8220000;
      3617: inst = 32'h10408000;
      3618: inst = 32'hc4046e4;
      3619: inst = 32'h8220000;
      3620: inst = 32'h10408000;
      3621: inst = 32'hc4046e5;
      3622: inst = 32'h8220000;
      3623: inst = 32'h10408000;
      3624: inst = 32'hc4046e6;
      3625: inst = 32'h8220000;
      3626: inst = 32'h10408000;
      3627: inst = 32'hc4046e7;
      3628: inst = 32'h8220000;
      3629: inst = 32'h10408000;
      3630: inst = 32'hc4046e8;
      3631: inst = 32'h8220000;
      3632: inst = 32'h10408000;
      3633: inst = 32'hc4046e9;
      3634: inst = 32'h8220000;
      3635: inst = 32'h10408000;
      3636: inst = 32'hc4046ea;
      3637: inst = 32'h8220000;
      3638: inst = 32'h10408000;
      3639: inst = 32'hc4046eb;
      3640: inst = 32'h8220000;
      3641: inst = 32'h10408000;
      3642: inst = 32'hc4046ec;
      3643: inst = 32'h8220000;
      3644: inst = 32'h10408000;
      3645: inst = 32'hc4046ed;
      3646: inst = 32'h8220000;
      3647: inst = 32'h10408000;
      3648: inst = 32'hc4046ee;
      3649: inst = 32'h8220000;
      3650: inst = 32'h10408000;
      3651: inst = 32'hc404700;
      3652: inst = 32'h8220000;
      3653: inst = 32'h10408000;
      3654: inst = 32'hc404701;
      3655: inst = 32'h8220000;
      3656: inst = 32'h10408000;
      3657: inst = 32'hc404702;
      3658: inst = 32'h8220000;
      3659: inst = 32'h10408000;
      3660: inst = 32'hc404703;
      3661: inst = 32'h8220000;
      3662: inst = 32'h10408000;
      3663: inst = 32'hc404704;
      3664: inst = 32'h8220000;
      3665: inst = 32'h10408000;
      3666: inst = 32'hc404705;
      3667: inst = 32'h8220000;
      3668: inst = 32'h10408000;
      3669: inst = 32'hc404706;
      3670: inst = 32'h8220000;
      3671: inst = 32'h10408000;
      3672: inst = 32'hc404707;
      3673: inst = 32'h8220000;
      3674: inst = 32'h10408000;
      3675: inst = 32'hc404708;
      3676: inst = 32'h8220000;
      3677: inst = 32'h10408000;
      3678: inst = 32'hc404709;
      3679: inst = 32'h8220000;
      3680: inst = 32'h10408000;
      3681: inst = 32'hc40470a;
      3682: inst = 32'h8220000;
      3683: inst = 32'h10408000;
      3684: inst = 32'hc40470b;
      3685: inst = 32'h8220000;
      3686: inst = 32'h10408000;
      3687: inst = 32'hc40470c;
      3688: inst = 32'h8220000;
      3689: inst = 32'h10408000;
      3690: inst = 32'hc40470d;
      3691: inst = 32'h8220000;
      3692: inst = 32'h10408000;
      3693: inst = 32'hc40470e;
      3694: inst = 32'h8220000;
      3695: inst = 32'h10408000;
      3696: inst = 32'hc40470f;
      3697: inst = 32'h8220000;
      3698: inst = 32'h10408000;
      3699: inst = 32'hc404710;
      3700: inst = 32'h8220000;
      3701: inst = 32'h10408000;
      3702: inst = 32'hc404711;
      3703: inst = 32'h8220000;
      3704: inst = 32'h10408000;
      3705: inst = 32'hc404712;
      3706: inst = 32'h8220000;
      3707: inst = 32'h10408000;
      3708: inst = 32'hc404713;
      3709: inst = 32'h8220000;
      3710: inst = 32'h10408000;
      3711: inst = 32'hc404714;
      3712: inst = 32'h8220000;
      3713: inst = 32'h10408000;
      3714: inst = 32'hc404715;
      3715: inst = 32'h8220000;
      3716: inst = 32'h10408000;
      3717: inst = 32'hc404716;
      3718: inst = 32'h8220000;
      3719: inst = 32'h10408000;
      3720: inst = 32'hc404717;
      3721: inst = 32'h8220000;
      3722: inst = 32'h10408000;
      3723: inst = 32'hc404718;
      3724: inst = 32'h8220000;
      3725: inst = 32'h10408000;
      3726: inst = 32'hc404719;
      3727: inst = 32'h8220000;
      3728: inst = 32'h10408000;
      3729: inst = 32'hc40471a;
      3730: inst = 32'h8220000;
      3731: inst = 32'h10408000;
      3732: inst = 32'hc40471b;
      3733: inst = 32'h8220000;
      3734: inst = 32'h10408000;
      3735: inst = 32'hc404744;
      3736: inst = 32'h8220000;
      3737: inst = 32'h10408000;
      3738: inst = 32'hc404745;
      3739: inst = 32'h8220000;
      3740: inst = 32'h10408000;
      3741: inst = 32'hc404746;
      3742: inst = 32'h8220000;
      3743: inst = 32'h10408000;
      3744: inst = 32'hc404747;
      3745: inst = 32'h8220000;
      3746: inst = 32'h10408000;
      3747: inst = 32'hc404748;
      3748: inst = 32'h8220000;
      3749: inst = 32'h10408000;
      3750: inst = 32'hc404749;
      3751: inst = 32'h8220000;
      3752: inst = 32'h10408000;
      3753: inst = 32'hc40474a;
      3754: inst = 32'h8220000;
      3755: inst = 32'h10408000;
      3756: inst = 32'hc40474b;
      3757: inst = 32'h8220000;
      3758: inst = 32'h10408000;
      3759: inst = 32'hc40474c;
      3760: inst = 32'h8220000;
      3761: inst = 32'h10408000;
      3762: inst = 32'hc40474d;
      3763: inst = 32'h8220000;
      3764: inst = 32'h10408000;
      3765: inst = 32'hc40474e;
      3766: inst = 32'h8220000;
      3767: inst = 32'h10408000;
      3768: inst = 32'hc404760;
      3769: inst = 32'h8220000;
      3770: inst = 32'h10408000;
      3771: inst = 32'hc404761;
      3772: inst = 32'h8220000;
      3773: inst = 32'h10408000;
      3774: inst = 32'hc404762;
      3775: inst = 32'h8220000;
      3776: inst = 32'h10408000;
      3777: inst = 32'hc404763;
      3778: inst = 32'h8220000;
      3779: inst = 32'h10408000;
      3780: inst = 32'hc404764;
      3781: inst = 32'h8220000;
      3782: inst = 32'h10408000;
      3783: inst = 32'hc404765;
      3784: inst = 32'h8220000;
      3785: inst = 32'h10408000;
      3786: inst = 32'hc404766;
      3787: inst = 32'h8220000;
      3788: inst = 32'h10408000;
      3789: inst = 32'hc404767;
      3790: inst = 32'h8220000;
      3791: inst = 32'h10408000;
      3792: inst = 32'hc404768;
      3793: inst = 32'h8220000;
      3794: inst = 32'h10408000;
      3795: inst = 32'hc404769;
      3796: inst = 32'h8220000;
      3797: inst = 32'h10408000;
      3798: inst = 32'hc40476a;
      3799: inst = 32'h8220000;
      3800: inst = 32'h10408000;
      3801: inst = 32'hc40476b;
      3802: inst = 32'h8220000;
      3803: inst = 32'h10408000;
      3804: inst = 32'hc40476c;
      3805: inst = 32'h8220000;
      3806: inst = 32'h10408000;
      3807: inst = 32'hc40476d;
      3808: inst = 32'h8220000;
      3809: inst = 32'h10408000;
      3810: inst = 32'hc40476e;
      3811: inst = 32'h8220000;
      3812: inst = 32'h10408000;
      3813: inst = 32'hc40476f;
      3814: inst = 32'h8220000;
      3815: inst = 32'h10408000;
      3816: inst = 32'hc404770;
      3817: inst = 32'h8220000;
      3818: inst = 32'h10408000;
      3819: inst = 32'hc404771;
      3820: inst = 32'h8220000;
      3821: inst = 32'h10408000;
      3822: inst = 32'hc404772;
      3823: inst = 32'h8220000;
      3824: inst = 32'h10408000;
      3825: inst = 32'hc404773;
      3826: inst = 32'h8220000;
      3827: inst = 32'h10408000;
      3828: inst = 32'hc404774;
      3829: inst = 32'h8220000;
      3830: inst = 32'h10408000;
      3831: inst = 32'hc404775;
      3832: inst = 32'h8220000;
      3833: inst = 32'h10408000;
      3834: inst = 32'hc404776;
      3835: inst = 32'h8220000;
      3836: inst = 32'h10408000;
      3837: inst = 32'hc404777;
      3838: inst = 32'h8220000;
      3839: inst = 32'h10408000;
      3840: inst = 32'hc404778;
      3841: inst = 32'h8220000;
      3842: inst = 32'h10408000;
      3843: inst = 32'hc404779;
      3844: inst = 32'h8220000;
      3845: inst = 32'h10408000;
      3846: inst = 32'hc40477a;
      3847: inst = 32'h8220000;
      3848: inst = 32'h10408000;
      3849: inst = 32'hc40477b;
      3850: inst = 32'h8220000;
      3851: inst = 32'h10408000;
      3852: inst = 32'hc4047a4;
      3853: inst = 32'h8220000;
      3854: inst = 32'h10408000;
      3855: inst = 32'hc4047a5;
      3856: inst = 32'h8220000;
      3857: inst = 32'h10408000;
      3858: inst = 32'hc4047a6;
      3859: inst = 32'h8220000;
      3860: inst = 32'h10408000;
      3861: inst = 32'hc4047a7;
      3862: inst = 32'h8220000;
      3863: inst = 32'h10408000;
      3864: inst = 32'hc4047a8;
      3865: inst = 32'h8220000;
      3866: inst = 32'h10408000;
      3867: inst = 32'hc4047a9;
      3868: inst = 32'h8220000;
      3869: inst = 32'h10408000;
      3870: inst = 32'hc4047aa;
      3871: inst = 32'h8220000;
      3872: inst = 32'h10408000;
      3873: inst = 32'hc4047ab;
      3874: inst = 32'h8220000;
      3875: inst = 32'h10408000;
      3876: inst = 32'hc4047ac;
      3877: inst = 32'h8220000;
      3878: inst = 32'h10408000;
      3879: inst = 32'hc4047ad;
      3880: inst = 32'h8220000;
      3881: inst = 32'h10408000;
      3882: inst = 32'hc4047ae;
      3883: inst = 32'h8220000;
      3884: inst = 32'h10408000;
      3885: inst = 32'hc4047c0;
      3886: inst = 32'h8220000;
      3887: inst = 32'h10408000;
      3888: inst = 32'hc4047c1;
      3889: inst = 32'h8220000;
      3890: inst = 32'h10408000;
      3891: inst = 32'hc4047c2;
      3892: inst = 32'h8220000;
      3893: inst = 32'h10408000;
      3894: inst = 32'hc4047c3;
      3895: inst = 32'h8220000;
      3896: inst = 32'h10408000;
      3897: inst = 32'hc4047c4;
      3898: inst = 32'h8220000;
      3899: inst = 32'h10408000;
      3900: inst = 32'hc4047c5;
      3901: inst = 32'h8220000;
      3902: inst = 32'h10408000;
      3903: inst = 32'hc4047c6;
      3904: inst = 32'h8220000;
      3905: inst = 32'h10408000;
      3906: inst = 32'hc4047c7;
      3907: inst = 32'h8220000;
      3908: inst = 32'h10408000;
      3909: inst = 32'hc4047c8;
      3910: inst = 32'h8220000;
      3911: inst = 32'h10408000;
      3912: inst = 32'hc4047c9;
      3913: inst = 32'h8220000;
      3914: inst = 32'h10408000;
      3915: inst = 32'hc4047ca;
      3916: inst = 32'h8220000;
      3917: inst = 32'h10408000;
      3918: inst = 32'hc4047cb;
      3919: inst = 32'h8220000;
      3920: inst = 32'h10408000;
      3921: inst = 32'hc4047cc;
      3922: inst = 32'h8220000;
      3923: inst = 32'h10408000;
      3924: inst = 32'hc4047cd;
      3925: inst = 32'h8220000;
      3926: inst = 32'h10408000;
      3927: inst = 32'hc4047ce;
      3928: inst = 32'h8220000;
      3929: inst = 32'h10408000;
      3930: inst = 32'hc4047cf;
      3931: inst = 32'h8220000;
      3932: inst = 32'h10408000;
      3933: inst = 32'hc4047d0;
      3934: inst = 32'h8220000;
      3935: inst = 32'h10408000;
      3936: inst = 32'hc4047d1;
      3937: inst = 32'h8220000;
      3938: inst = 32'h10408000;
      3939: inst = 32'hc4047d2;
      3940: inst = 32'h8220000;
      3941: inst = 32'h10408000;
      3942: inst = 32'hc4047d3;
      3943: inst = 32'h8220000;
      3944: inst = 32'h10408000;
      3945: inst = 32'hc4047d4;
      3946: inst = 32'h8220000;
      3947: inst = 32'h10408000;
      3948: inst = 32'hc4047d5;
      3949: inst = 32'h8220000;
      3950: inst = 32'h10408000;
      3951: inst = 32'hc4047d6;
      3952: inst = 32'h8220000;
      3953: inst = 32'h10408000;
      3954: inst = 32'hc4047d7;
      3955: inst = 32'h8220000;
      3956: inst = 32'h10408000;
      3957: inst = 32'hc4047d8;
      3958: inst = 32'h8220000;
      3959: inst = 32'h10408000;
      3960: inst = 32'hc4047d9;
      3961: inst = 32'h8220000;
      3962: inst = 32'h10408000;
      3963: inst = 32'hc4047da;
      3964: inst = 32'h8220000;
      3965: inst = 32'h10408000;
      3966: inst = 32'hc4047db;
      3967: inst = 32'h8220000;
      3968: inst = 32'h10408000;
      3969: inst = 32'hc404804;
      3970: inst = 32'h8220000;
      3971: inst = 32'h10408000;
      3972: inst = 32'hc404805;
      3973: inst = 32'h8220000;
      3974: inst = 32'h10408000;
      3975: inst = 32'hc404806;
      3976: inst = 32'h8220000;
      3977: inst = 32'h10408000;
      3978: inst = 32'hc404807;
      3979: inst = 32'h8220000;
      3980: inst = 32'h10408000;
      3981: inst = 32'hc404808;
      3982: inst = 32'h8220000;
      3983: inst = 32'h10408000;
      3984: inst = 32'hc404809;
      3985: inst = 32'h8220000;
      3986: inst = 32'h10408000;
      3987: inst = 32'hc40480a;
      3988: inst = 32'h8220000;
      3989: inst = 32'h10408000;
      3990: inst = 32'hc40480b;
      3991: inst = 32'h8220000;
      3992: inst = 32'h10408000;
      3993: inst = 32'hc40480c;
      3994: inst = 32'h8220000;
      3995: inst = 32'h10408000;
      3996: inst = 32'hc40480d;
      3997: inst = 32'h8220000;
      3998: inst = 32'h10408000;
      3999: inst = 32'hc40480e;
      4000: inst = 32'h8220000;
      4001: inst = 32'h10408000;
      4002: inst = 32'hc404820;
      4003: inst = 32'h8220000;
      4004: inst = 32'h10408000;
      4005: inst = 32'hc404821;
      4006: inst = 32'h8220000;
      4007: inst = 32'h10408000;
      4008: inst = 32'hc404822;
      4009: inst = 32'h8220000;
      4010: inst = 32'h10408000;
      4011: inst = 32'hc404823;
      4012: inst = 32'h8220000;
      4013: inst = 32'h10408000;
      4014: inst = 32'hc404824;
      4015: inst = 32'h8220000;
      4016: inst = 32'h10408000;
      4017: inst = 32'hc404825;
      4018: inst = 32'h8220000;
      4019: inst = 32'h10408000;
      4020: inst = 32'hc404826;
      4021: inst = 32'h8220000;
      4022: inst = 32'h10408000;
      4023: inst = 32'hc404827;
      4024: inst = 32'h8220000;
      4025: inst = 32'h10408000;
      4026: inst = 32'hc404828;
      4027: inst = 32'h8220000;
      4028: inst = 32'h10408000;
      4029: inst = 32'hc404829;
      4030: inst = 32'h8220000;
      4031: inst = 32'h10408000;
      4032: inst = 32'hc40482a;
      4033: inst = 32'h8220000;
      4034: inst = 32'h10408000;
      4035: inst = 32'hc40482b;
      4036: inst = 32'h8220000;
      4037: inst = 32'h10408000;
      4038: inst = 32'hc40482c;
      4039: inst = 32'h8220000;
      4040: inst = 32'h10408000;
      4041: inst = 32'hc40482d;
      4042: inst = 32'h8220000;
      4043: inst = 32'h10408000;
      4044: inst = 32'hc40482e;
      4045: inst = 32'h8220000;
      4046: inst = 32'h10408000;
      4047: inst = 32'hc40482f;
      4048: inst = 32'h8220000;
      4049: inst = 32'h10408000;
      4050: inst = 32'hc404830;
      4051: inst = 32'h8220000;
      4052: inst = 32'h10408000;
      4053: inst = 32'hc404831;
      4054: inst = 32'h8220000;
      4055: inst = 32'h10408000;
      4056: inst = 32'hc404832;
      4057: inst = 32'h8220000;
      4058: inst = 32'h10408000;
      4059: inst = 32'hc404833;
      4060: inst = 32'h8220000;
      4061: inst = 32'h10408000;
      4062: inst = 32'hc404834;
      4063: inst = 32'h8220000;
      4064: inst = 32'h10408000;
      4065: inst = 32'hc404835;
      4066: inst = 32'h8220000;
      4067: inst = 32'h10408000;
      4068: inst = 32'hc404836;
      4069: inst = 32'h8220000;
      4070: inst = 32'h10408000;
      4071: inst = 32'hc404837;
      4072: inst = 32'h8220000;
      4073: inst = 32'h10408000;
      4074: inst = 32'hc404838;
      4075: inst = 32'h8220000;
      4076: inst = 32'h10408000;
      4077: inst = 32'hc404839;
      4078: inst = 32'h8220000;
      4079: inst = 32'h10408000;
      4080: inst = 32'hc40483a;
      4081: inst = 32'h8220000;
      4082: inst = 32'h10408000;
      4083: inst = 32'hc40483b;
      4084: inst = 32'h8220000;
      4085: inst = 32'h10408000;
      4086: inst = 32'hc404864;
      4087: inst = 32'h8220000;
      4088: inst = 32'h10408000;
      4089: inst = 32'hc404865;
      4090: inst = 32'h8220000;
      4091: inst = 32'h10408000;
      4092: inst = 32'hc404866;
      4093: inst = 32'h8220000;
      4094: inst = 32'h10408000;
      4095: inst = 32'hc404867;
      4096: inst = 32'h8220000;
      4097: inst = 32'h10408000;
      4098: inst = 32'hc404868;
      4099: inst = 32'h8220000;
      4100: inst = 32'h10408000;
      4101: inst = 32'hc404869;
      4102: inst = 32'h8220000;
      4103: inst = 32'h10408000;
      4104: inst = 32'hc40486a;
      4105: inst = 32'h8220000;
      4106: inst = 32'h10408000;
      4107: inst = 32'hc40486b;
      4108: inst = 32'h8220000;
      4109: inst = 32'h10408000;
      4110: inst = 32'hc40486c;
      4111: inst = 32'h8220000;
      4112: inst = 32'h10408000;
      4113: inst = 32'hc40486d;
      4114: inst = 32'h8220000;
      4115: inst = 32'h10408000;
      4116: inst = 32'hc40486e;
      4117: inst = 32'h8220000;
      4118: inst = 32'h10408000;
      4119: inst = 32'hc404880;
      4120: inst = 32'h8220000;
      4121: inst = 32'h10408000;
      4122: inst = 32'hc404881;
      4123: inst = 32'h8220000;
      4124: inst = 32'h10408000;
      4125: inst = 32'hc404882;
      4126: inst = 32'h8220000;
      4127: inst = 32'h10408000;
      4128: inst = 32'hc404883;
      4129: inst = 32'h8220000;
      4130: inst = 32'h10408000;
      4131: inst = 32'hc404884;
      4132: inst = 32'h8220000;
      4133: inst = 32'h10408000;
      4134: inst = 32'hc404885;
      4135: inst = 32'h8220000;
      4136: inst = 32'h10408000;
      4137: inst = 32'hc404886;
      4138: inst = 32'h8220000;
      4139: inst = 32'h10408000;
      4140: inst = 32'hc404887;
      4141: inst = 32'h8220000;
      4142: inst = 32'h10408000;
      4143: inst = 32'hc404888;
      4144: inst = 32'h8220000;
      4145: inst = 32'h10408000;
      4146: inst = 32'hc404889;
      4147: inst = 32'h8220000;
      4148: inst = 32'h10408000;
      4149: inst = 32'hc40488a;
      4150: inst = 32'h8220000;
      4151: inst = 32'h10408000;
      4152: inst = 32'hc40488b;
      4153: inst = 32'h8220000;
      4154: inst = 32'h10408000;
      4155: inst = 32'hc40488c;
      4156: inst = 32'h8220000;
      4157: inst = 32'h10408000;
      4158: inst = 32'hc40488d;
      4159: inst = 32'h8220000;
      4160: inst = 32'h10408000;
      4161: inst = 32'hc40488e;
      4162: inst = 32'h8220000;
      4163: inst = 32'h10408000;
      4164: inst = 32'hc40488f;
      4165: inst = 32'h8220000;
      4166: inst = 32'h10408000;
      4167: inst = 32'hc404890;
      4168: inst = 32'h8220000;
      4169: inst = 32'h10408000;
      4170: inst = 32'hc404891;
      4171: inst = 32'h8220000;
      4172: inst = 32'h10408000;
      4173: inst = 32'hc404892;
      4174: inst = 32'h8220000;
      4175: inst = 32'h10408000;
      4176: inst = 32'hc404893;
      4177: inst = 32'h8220000;
      4178: inst = 32'h10408000;
      4179: inst = 32'hc404894;
      4180: inst = 32'h8220000;
      4181: inst = 32'h10408000;
      4182: inst = 32'hc404895;
      4183: inst = 32'h8220000;
      4184: inst = 32'h10408000;
      4185: inst = 32'hc404896;
      4186: inst = 32'h8220000;
      4187: inst = 32'h10408000;
      4188: inst = 32'hc404897;
      4189: inst = 32'h8220000;
      4190: inst = 32'h10408000;
      4191: inst = 32'hc404898;
      4192: inst = 32'h8220000;
      4193: inst = 32'h10408000;
      4194: inst = 32'hc404899;
      4195: inst = 32'h8220000;
      4196: inst = 32'h10408000;
      4197: inst = 32'hc40489a;
      4198: inst = 32'h8220000;
      4199: inst = 32'h10408000;
      4200: inst = 32'hc40489b;
      4201: inst = 32'h8220000;
      4202: inst = 32'h10408000;
      4203: inst = 32'hc4048c4;
      4204: inst = 32'h8220000;
      4205: inst = 32'h10408000;
      4206: inst = 32'hc4048c5;
      4207: inst = 32'h8220000;
      4208: inst = 32'h10408000;
      4209: inst = 32'hc4048c6;
      4210: inst = 32'h8220000;
      4211: inst = 32'h10408000;
      4212: inst = 32'hc4048c7;
      4213: inst = 32'h8220000;
      4214: inst = 32'h10408000;
      4215: inst = 32'hc4048c8;
      4216: inst = 32'h8220000;
      4217: inst = 32'h10408000;
      4218: inst = 32'hc4048c9;
      4219: inst = 32'h8220000;
      4220: inst = 32'h10408000;
      4221: inst = 32'hc4048ca;
      4222: inst = 32'h8220000;
      4223: inst = 32'h10408000;
      4224: inst = 32'hc4048cb;
      4225: inst = 32'h8220000;
      4226: inst = 32'h10408000;
      4227: inst = 32'hc4048cc;
      4228: inst = 32'h8220000;
      4229: inst = 32'h10408000;
      4230: inst = 32'hc4048cd;
      4231: inst = 32'h8220000;
      4232: inst = 32'h10408000;
      4233: inst = 32'hc4048ce;
      4234: inst = 32'h8220000;
      4235: inst = 32'h10408000;
      4236: inst = 32'hc4048e0;
      4237: inst = 32'h8220000;
      4238: inst = 32'h10408000;
      4239: inst = 32'hc4048e1;
      4240: inst = 32'h8220000;
      4241: inst = 32'h10408000;
      4242: inst = 32'hc4048e2;
      4243: inst = 32'h8220000;
      4244: inst = 32'h10408000;
      4245: inst = 32'hc4048e3;
      4246: inst = 32'h8220000;
      4247: inst = 32'h10408000;
      4248: inst = 32'hc4048e4;
      4249: inst = 32'h8220000;
      4250: inst = 32'h10408000;
      4251: inst = 32'hc4048e5;
      4252: inst = 32'h8220000;
      4253: inst = 32'h10408000;
      4254: inst = 32'hc4048e6;
      4255: inst = 32'h8220000;
      4256: inst = 32'h10408000;
      4257: inst = 32'hc4048e7;
      4258: inst = 32'h8220000;
      4259: inst = 32'h10408000;
      4260: inst = 32'hc4048e8;
      4261: inst = 32'h8220000;
      4262: inst = 32'h10408000;
      4263: inst = 32'hc4048e9;
      4264: inst = 32'h8220000;
      4265: inst = 32'h10408000;
      4266: inst = 32'hc4048ea;
      4267: inst = 32'h8220000;
      4268: inst = 32'h10408000;
      4269: inst = 32'hc4048eb;
      4270: inst = 32'h8220000;
      4271: inst = 32'h10408000;
      4272: inst = 32'hc4048ec;
      4273: inst = 32'h8220000;
      4274: inst = 32'h10408000;
      4275: inst = 32'hc4048ed;
      4276: inst = 32'h8220000;
      4277: inst = 32'h10408000;
      4278: inst = 32'hc4048ee;
      4279: inst = 32'h8220000;
      4280: inst = 32'h10408000;
      4281: inst = 32'hc4048ef;
      4282: inst = 32'h8220000;
      4283: inst = 32'h10408000;
      4284: inst = 32'hc4048f0;
      4285: inst = 32'h8220000;
      4286: inst = 32'h10408000;
      4287: inst = 32'hc4048f1;
      4288: inst = 32'h8220000;
      4289: inst = 32'h10408000;
      4290: inst = 32'hc4048f2;
      4291: inst = 32'h8220000;
      4292: inst = 32'h10408000;
      4293: inst = 32'hc4048f3;
      4294: inst = 32'h8220000;
      4295: inst = 32'h10408000;
      4296: inst = 32'hc4048f4;
      4297: inst = 32'h8220000;
      4298: inst = 32'h10408000;
      4299: inst = 32'hc4048f5;
      4300: inst = 32'h8220000;
      4301: inst = 32'h10408000;
      4302: inst = 32'hc4048f6;
      4303: inst = 32'h8220000;
      4304: inst = 32'h10408000;
      4305: inst = 32'hc4048f7;
      4306: inst = 32'h8220000;
      4307: inst = 32'h10408000;
      4308: inst = 32'hc4048f8;
      4309: inst = 32'h8220000;
      4310: inst = 32'h10408000;
      4311: inst = 32'hc4048f9;
      4312: inst = 32'h8220000;
      4313: inst = 32'h10408000;
      4314: inst = 32'hc4048fa;
      4315: inst = 32'h8220000;
      4316: inst = 32'h10408000;
      4317: inst = 32'hc4048fb;
      4318: inst = 32'h8220000;
      4319: inst = 32'h10408000;
      4320: inst = 32'hc404924;
      4321: inst = 32'h8220000;
      4322: inst = 32'h10408000;
      4323: inst = 32'hc404925;
      4324: inst = 32'h8220000;
      4325: inst = 32'h10408000;
      4326: inst = 32'hc404926;
      4327: inst = 32'h8220000;
      4328: inst = 32'h10408000;
      4329: inst = 32'hc404927;
      4330: inst = 32'h8220000;
      4331: inst = 32'h10408000;
      4332: inst = 32'hc404928;
      4333: inst = 32'h8220000;
      4334: inst = 32'h10408000;
      4335: inst = 32'hc404929;
      4336: inst = 32'h8220000;
      4337: inst = 32'h10408000;
      4338: inst = 32'hc40492a;
      4339: inst = 32'h8220000;
      4340: inst = 32'h10408000;
      4341: inst = 32'hc40492b;
      4342: inst = 32'h8220000;
      4343: inst = 32'h10408000;
      4344: inst = 32'hc40492c;
      4345: inst = 32'h8220000;
      4346: inst = 32'h10408000;
      4347: inst = 32'hc40492d;
      4348: inst = 32'h8220000;
      4349: inst = 32'h10408000;
      4350: inst = 32'hc40492e;
      4351: inst = 32'h8220000;
      4352: inst = 32'h10408000;
      4353: inst = 32'hc404940;
      4354: inst = 32'h8220000;
      4355: inst = 32'h10408000;
      4356: inst = 32'hc404941;
      4357: inst = 32'h8220000;
      4358: inst = 32'h10408000;
      4359: inst = 32'hc404942;
      4360: inst = 32'h8220000;
      4361: inst = 32'h10408000;
      4362: inst = 32'hc404943;
      4363: inst = 32'h8220000;
      4364: inst = 32'h10408000;
      4365: inst = 32'hc404944;
      4366: inst = 32'h8220000;
      4367: inst = 32'h10408000;
      4368: inst = 32'hc404945;
      4369: inst = 32'h8220000;
      4370: inst = 32'h10408000;
      4371: inst = 32'hc404946;
      4372: inst = 32'h8220000;
      4373: inst = 32'h10408000;
      4374: inst = 32'hc404947;
      4375: inst = 32'h8220000;
      4376: inst = 32'h10408000;
      4377: inst = 32'hc404948;
      4378: inst = 32'h8220000;
      4379: inst = 32'h10408000;
      4380: inst = 32'hc404949;
      4381: inst = 32'h8220000;
      4382: inst = 32'h10408000;
      4383: inst = 32'hc40494a;
      4384: inst = 32'h8220000;
      4385: inst = 32'h10408000;
      4386: inst = 32'hc40494b;
      4387: inst = 32'h8220000;
      4388: inst = 32'h10408000;
      4389: inst = 32'hc40494c;
      4390: inst = 32'h8220000;
      4391: inst = 32'h10408000;
      4392: inst = 32'hc40494d;
      4393: inst = 32'h8220000;
      4394: inst = 32'h10408000;
      4395: inst = 32'hc40494e;
      4396: inst = 32'h8220000;
      4397: inst = 32'h10408000;
      4398: inst = 32'hc40494f;
      4399: inst = 32'h8220000;
      4400: inst = 32'h10408000;
      4401: inst = 32'hc404950;
      4402: inst = 32'h8220000;
      4403: inst = 32'h10408000;
      4404: inst = 32'hc404951;
      4405: inst = 32'h8220000;
      4406: inst = 32'h10408000;
      4407: inst = 32'hc404952;
      4408: inst = 32'h8220000;
      4409: inst = 32'h10408000;
      4410: inst = 32'hc404953;
      4411: inst = 32'h8220000;
      4412: inst = 32'h10408000;
      4413: inst = 32'hc404954;
      4414: inst = 32'h8220000;
      4415: inst = 32'h10408000;
      4416: inst = 32'hc404955;
      4417: inst = 32'h8220000;
      4418: inst = 32'h10408000;
      4419: inst = 32'hc404956;
      4420: inst = 32'h8220000;
      4421: inst = 32'h10408000;
      4422: inst = 32'hc404957;
      4423: inst = 32'h8220000;
      4424: inst = 32'h10408000;
      4425: inst = 32'hc404958;
      4426: inst = 32'h8220000;
      4427: inst = 32'h10408000;
      4428: inst = 32'hc404959;
      4429: inst = 32'h8220000;
      4430: inst = 32'h10408000;
      4431: inst = 32'hc40495a;
      4432: inst = 32'h8220000;
      4433: inst = 32'h10408000;
      4434: inst = 32'hc40495b;
      4435: inst = 32'h8220000;
      4436: inst = 32'h10408000;
      4437: inst = 32'hc404984;
      4438: inst = 32'h8220000;
      4439: inst = 32'h10408000;
      4440: inst = 32'hc404985;
      4441: inst = 32'h8220000;
      4442: inst = 32'h10408000;
      4443: inst = 32'hc404986;
      4444: inst = 32'h8220000;
      4445: inst = 32'h10408000;
      4446: inst = 32'hc404987;
      4447: inst = 32'h8220000;
      4448: inst = 32'h10408000;
      4449: inst = 32'hc404988;
      4450: inst = 32'h8220000;
      4451: inst = 32'h10408000;
      4452: inst = 32'hc404989;
      4453: inst = 32'h8220000;
      4454: inst = 32'h10408000;
      4455: inst = 32'hc40498a;
      4456: inst = 32'h8220000;
      4457: inst = 32'h10408000;
      4458: inst = 32'hc40498b;
      4459: inst = 32'h8220000;
      4460: inst = 32'h10408000;
      4461: inst = 32'hc40498c;
      4462: inst = 32'h8220000;
      4463: inst = 32'h10408000;
      4464: inst = 32'hc40498d;
      4465: inst = 32'h8220000;
      4466: inst = 32'h10408000;
      4467: inst = 32'hc40498e;
      4468: inst = 32'h8220000;
      4469: inst = 32'h10408000;
      4470: inst = 32'hc4049a0;
      4471: inst = 32'h8220000;
      4472: inst = 32'h10408000;
      4473: inst = 32'hc4049a1;
      4474: inst = 32'h8220000;
      4475: inst = 32'h10408000;
      4476: inst = 32'hc4049a2;
      4477: inst = 32'h8220000;
      4478: inst = 32'h10408000;
      4479: inst = 32'hc4049a3;
      4480: inst = 32'h8220000;
      4481: inst = 32'h10408000;
      4482: inst = 32'hc4049a4;
      4483: inst = 32'h8220000;
      4484: inst = 32'h10408000;
      4485: inst = 32'hc4049a5;
      4486: inst = 32'h8220000;
      4487: inst = 32'h10408000;
      4488: inst = 32'hc4049a6;
      4489: inst = 32'h8220000;
      4490: inst = 32'h10408000;
      4491: inst = 32'hc4049a7;
      4492: inst = 32'h8220000;
      4493: inst = 32'h10408000;
      4494: inst = 32'hc4049a8;
      4495: inst = 32'h8220000;
      4496: inst = 32'h10408000;
      4497: inst = 32'hc4049a9;
      4498: inst = 32'h8220000;
      4499: inst = 32'h10408000;
      4500: inst = 32'hc4049aa;
      4501: inst = 32'h8220000;
      4502: inst = 32'h10408000;
      4503: inst = 32'hc4049ab;
      4504: inst = 32'h8220000;
      4505: inst = 32'h10408000;
      4506: inst = 32'hc4049ac;
      4507: inst = 32'h8220000;
      4508: inst = 32'h10408000;
      4509: inst = 32'hc4049ad;
      4510: inst = 32'h8220000;
      4511: inst = 32'h10408000;
      4512: inst = 32'hc4049ae;
      4513: inst = 32'h8220000;
      4514: inst = 32'h10408000;
      4515: inst = 32'hc4049af;
      4516: inst = 32'h8220000;
      4517: inst = 32'h10408000;
      4518: inst = 32'hc4049b0;
      4519: inst = 32'h8220000;
      4520: inst = 32'h10408000;
      4521: inst = 32'hc4049b1;
      4522: inst = 32'h8220000;
      4523: inst = 32'h10408000;
      4524: inst = 32'hc4049b2;
      4525: inst = 32'h8220000;
      4526: inst = 32'h10408000;
      4527: inst = 32'hc4049b3;
      4528: inst = 32'h8220000;
      4529: inst = 32'h10408000;
      4530: inst = 32'hc4049b4;
      4531: inst = 32'h8220000;
      4532: inst = 32'h10408000;
      4533: inst = 32'hc4049b5;
      4534: inst = 32'h8220000;
      4535: inst = 32'h10408000;
      4536: inst = 32'hc4049b6;
      4537: inst = 32'h8220000;
      4538: inst = 32'h10408000;
      4539: inst = 32'hc4049b7;
      4540: inst = 32'h8220000;
      4541: inst = 32'h10408000;
      4542: inst = 32'hc4049b8;
      4543: inst = 32'h8220000;
      4544: inst = 32'h10408000;
      4545: inst = 32'hc4049b9;
      4546: inst = 32'h8220000;
      4547: inst = 32'h10408000;
      4548: inst = 32'hc4049ba;
      4549: inst = 32'h8220000;
      4550: inst = 32'h10408000;
      4551: inst = 32'hc4049bb;
      4552: inst = 32'h8220000;
      4553: inst = 32'h10408000;
      4554: inst = 32'hc4049e4;
      4555: inst = 32'h8220000;
      4556: inst = 32'h10408000;
      4557: inst = 32'hc4049e5;
      4558: inst = 32'h8220000;
      4559: inst = 32'h10408000;
      4560: inst = 32'hc4049e6;
      4561: inst = 32'h8220000;
      4562: inst = 32'h10408000;
      4563: inst = 32'hc4049e7;
      4564: inst = 32'h8220000;
      4565: inst = 32'h10408000;
      4566: inst = 32'hc4049e8;
      4567: inst = 32'h8220000;
      4568: inst = 32'h10408000;
      4569: inst = 32'hc4049e9;
      4570: inst = 32'h8220000;
      4571: inst = 32'h10408000;
      4572: inst = 32'hc4049ea;
      4573: inst = 32'h8220000;
      4574: inst = 32'h10408000;
      4575: inst = 32'hc4049eb;
      4576: inst = 32'h8220000;
      4577: inst = 32'h10408000;
      4578: inst = 32'hc4049ec;
      4579: inst = 32'h8220000;
      4580: inst = 32'h10408000;
      4581: inst = 32'hc4049ed;
      4582: inst = 32'h8220000;
      4583: inst = 32'h10408000;
      4584: inst = 32'hc4049ee;
      4585: inst = 32'h8220000;
      4586: inst = 32'h10408000;
      4587: inst = 32'hc404a00;
      4588: inst = 32'h8220000;
      4589: inst = 32'h10408000;
      4590: inst = 32'hc404a01;
      4591: inst = 32'h8220000;
      4592: inst = 32'h10408000;
      4593: inst = 32'hc404a02;
      4594: inst = 32'h8220000;
      4595: inst = 32'h10408000;
      4596: inst = 32'hc404a03;
      4597: inst = 32'h8220000;
      4598: inst = 32'h10408000;
      4599: inst = 32'hc404a04;
      4600: inst = 32'h8220000;
      4601: inst = 32'h10408000;
      4602: inst = 32'hc404a05;
      4603: inst = 32'h8220000;
      4604: inst = 32'h10408000;
      4605: inst = 32'hc404a06;
      4606: inst = 32'h8220000;
      4607: inst = 32'h10408000;
      4608: inst = 32'hc404a07;
      4609: inst = 32'h8220000;
      4610: inst = 32'h10408000;
      4611: inst = 32'hc404a0f;
      4612: inst = 32'h8220000;
      4613: inst = 32'h10408000;
      4614: inst = 32'hc404a10;
      4615: inst = 32'h8220000;
      4616: inst = 32'h10408000;
      4617: inst = 32'hc404a11;
      4618: inst = 32'h8220000;
      4619: inst = 32'h10408000;
      4620: inst = 32'hc404a12;
      4621: inst = 32'h8220000;
      4622: inst = 32'h10408000;
      4623: inst = 32'hc404a13;
      4624: inst = 32'h8220000;
      4625: inst = 32'h10408000;
      4626: inst = 32'hc404a14;
      4627: inst = 32'h8220000;
      4628: inst = 32'h10408000;
      4629: inst = 32'hc404a15;
      4630: inst = 32'h8220000;
      4631: inst = 32'h10408000;
      4632: inst = 32'hc404a16;
      4633: inst = 32'h8220000;
      4634: inst = 32'h10408000;
      4635: inst = 32'hc404a17;
      4636: inst = 32'h8220000;
      4637: inst = 32'h10408000;
      4638: inst = 32'hc404a18;
      4639: inst = 32'h8220000;
      4640: inst = 32'h10408000;
      4641: inst = 32'hc404a19;
      4642: inst = 32'h8220000;
      4643: inst = 32'h10408000;
      4644: inst = 32'hc404a1a;
      4645: inst = 32'h8220000;
      4646: inst = 32'h10408000;
      4647: inst = 32'hc404a1b;
      4648: inst = 32'h8220000;
      4649: inst = 32'h10408000;
      4650: inst = 32'hc404a44;
      4651: inst = 32'h8220000;
      4652: inst = 32'h10408000;
      4653: inst = 32'hc404a45;
      4654: inst = 32'h8220000;
      4655: inst = 32'h10408000;
      4656: inst = 32'hc404a46;
      4657: inst = 32'h8220000;
      4658: inst = 32'h10408000;
      4659: inst = 32'hc404a47;
      4660: inst = 32'h8220000;
      4661: inst = 32'h10408000;
      4662: inst = 32'hc404a48;
      4663: inst = 32'h8220000;
      4664: inst = 32'h10408000;
      4665: inst = 32'hc404a49;
      4666: inst = 32'h8220000;
      4667: inst = 32'h10408000;
      4668: inst = 32'hc404a4a;
      4669: inst = 32'h8220000;
      4670: inst = 32'h10408000;
      4671: inst = 32'hc404a4b;
      4672: inst = 32'h8220000;
      4673: inst = 32'h10408000;
      4674: inst = 32'hc404a4c;
      4675: inst = 32'h8220000;
      4676: inst = 32'h10408000;
      4677: inst = 32'hc404a4d;
      4678: inst = 32'h8220000;
      4679: inst = 32'h10408000;
      4680: inst = 32'hc404a4e;
      4681: inst = 32'h8220000;
      4682: inst = 32'h10408000;
      4683: inst = 32'hc404a60;
      4684: inst = 32'h8220000;
      4685: inst = 32'h10408000;
      4686: inst = 32'hc404a61;
      4687: inst = 32'h8220000;
      4688: inst = 32'h10408000;
      4689: inst = 32'hc404a62;
      4690: inst = 32'h8220000;
      4691: inst = 32'h10408000;
      4692: inst = 32'hc404a63;
      4693: inst = 32'h8220000;
      4694: inst = 32'h10408000;
      4695: inst = 32'hc404a64;
      4696: inst = 32'h8220000;
      4697: inst = 32'h10408000;
      4698: inst = 32'hc404a65;
      4699: inst = 32'h8220000;
      4700: inst = 32'h10408000;
      4701: inst = 32'hc404a66;
      4702: inst = 32'h8220000;
      4703: inst = 32'h10408000;
      4704: inst = 32'hc404a70;
      4705: inst = 32'h8220000;
      4706: inst = 32'h10408000;
      4707: inst = 32'hc404a71;
      4708: inst = 32'h8220000;
      4709: inst = 32'h10408000;
      4710: inst = 32'hc404a72;
      4711: inst = 32'h8220000;
      4712: inst = 32'h10408000;
      4713: inst = 32'hc404a73;
      4714: inst = 32'h8220000;
      4715: inst = 32'h10408000;
      4716: inst = 32'hc404a74;
      4717: inst = 32'h8220000;
      4718: inst = 32'h10408000;
      4719: inst = 32'hc404a75;
      4720: inst = 32'h8220000;
      4721: inst = 32'h10408000;
      4722: inst = 32'hc404a76;
      4723: inst = 32'h8220000;
      4724: inst = 32'h10408000;
      4725: inst = 32'hc404a77;
      4726: inst = 32'h8220000;
      4727: inst = 32'h10408000;
      4728: inst = 32'hc404a78;
      4729: inst = 32'h8220000;
      4730: inst = 32'h10408000;
      4731: inst = 32'hc404a79;
      4732: inst = 32'h8220000;
      4733: inst = 32'h10408000;
      4734: inst = 32'hc404a7a;
      4735: inst = 32'h8220000;
      4736: inst = 32'h10408000;
      4737: inst = 32'hc404a7b;
      4738: inst = 32'h8220000;
      4739: inst = 32'h10408000;
      4740: inst = 32'hc404aa4;
      4741: inst = 32'h8220000;
      4742: inst = 32'h10408000;
      4743: inst = 32'hc404aa5;
      4744: inst = 32'h8220000;
      4745: inst = 32'h10408000;
      4746: inst = 32'hc404aa6;
      4747: inst = 32'h8220000;
      4748: inst = 32'h10408000;
      4749: inst = 32'hc404aa7;
      4750: inst = 32'h8220000;
      4751: inst = 32'h10408000;
      4752: inst = 32'hc404aa8;
      4753: inst = 32'h8220000;
      4754: inst = 32'h10408000;
      4755: inst = 32'hc404aa9;
      4756: inst = 32'h8220000;
      4757: inst = 32'h10408000;
      4758: inst = 32'hc404aaa;
      4759: inst = 32'h8220000;
      4760: inst = 32'h10408000;
      4761: inst = 32'hc404aab;
      4762: inst = 32'h8220000;
      4763: inst = 32'h10408000;
      4764: inst = 32'hc404aac;
      4765: inst = 32'h8220000;
      4766: inst = 32'h10408000;
      4767: inst = 32'hc404aad;
      4768: inst = 32'h8220000;
      4769: inst = 32'h10408000;
      4770: inst = 32'hc404aae;
      4771: inst = 32'h8220000;
      4772: inst = 32'h10408000;
      4773: inst = 32'hc404ac0;
      4774: inst = 32'h8220000;
      4775: inst = 32'h10408000;
      4776: inst = 32'hc404ac1;
      4777: inst = 32'h8220000;
      4778: inst = 32'h10408000;
      4779: inst = 32'hc404ac2;
      4780: inst = 32'h8220000;
      4781: inst = 32'h10408000;
      4782: inst = 32'hc404ac3;
      4783: inst = 32'h8220000;
      4784: inst = 32'h10408000;
      4785: inst = 32'hc404ac4;
      4786: inst = 32'h8220000;
      4787: inst = 32'h10408000;
      4788: inst = 32'hc404ac5;
      4789: inst = 32'h8220000;
      4790: inst = 32'h10408000;
      4791: inst = 32'hc404ac6;
      4792: inst = 32'h8220000;
      4793: inst = 32'h10408000;
      4794: inst = 32'hc404ad0;
      4795: inst = 32'h8220000;
      4796: inst = 32'h10408000;
      4797: inst = 32'hc404ad1;
      4798: inst = 32'h8220000;
      4799: inst = 32'h10408000;
      4800: inst = 32'hc404ad2;
      4801: inst = 32'h8220000;
      4802: inst = 32'h10408000;
      4803: inst = 32'hc404ad3;
      4804: inst = 32'h8220000;
      4805: inst = 32'h10408000;
      4806: inst = 32'hc404ad4;
      4807: inst = 32'h8220000;
      4808: inst = 32'h10408000;
      4809: inst = 32'hc404ad5;
      4810: inst = 32'h8220000;
      4811: inst = 32'h10408000;
      4812: inst = 32'hc404ad6;
      4813: inst = 32'h8220000;
      4814: inst = 32'h10408000;
      4815: inst = 32'hc404ad7;
      4816: inst = 32'h8220000;
      4817: inst = 32'h10408000;
      4818: inst = 32'hc404ad8;
      4819: inst = 32'h8220000;
      4820: inst = 32'h10408000;
      4821: inst = 32'hc404ad9;
      4822: inst = 32'h8220000;
      4823: inst = 32'h10408000;
      4824: inst = 32'hc404ada;
      4825: inst = 32'h8220000;
      4826: inst = 32'h10408000;
      4827: inst = 32'hc404adb;
      4828: inst = 32'h8220000;
      4829: inst = 32'h10408000;
      4830: inst = 32'hc404b04;
      4831: inst = 32'h8220000;
      4832: inst = 32'h10408000;
      4833: inst = 32'hc404b05;
      4834: inst = 32'h8220000;
      4835: inst = 32'h10408000;
      4836: inst = 32'hc404b06;
      4837: inst = 32'h8220000;
      4838: inst = 32'h10408000;
      4839: inst = 32'hc404b07;
      4840: inst = 32'h8220000;
      4841: inst = 32'h10408000;
      4842: inst = 32'hc404b08;
      4843: inst = 32'h8220000;
      4844: inst = 32'h10408000;
      4845: inst = 32'hc404b09;
      4846: inst = 32'h8220000;
      4847: inst = 32'h10408000;
      4848: inst = 32'hc404b0a;
      4849: inst = 32'h8220000;
      4850: inst = 32'h10408000;
      4851: inst = 32'hc404b0b;
      4852: inst = 32'h8220000;
      4853: inst = 32'h10408000;
      4854: inst = 32'hc404b0c;
      4855: inst = 32'h8220000;
      4856: inst = 32'h10408000;
      4857: inst = 32'hc404b0d;
      4858: inst = 32'h8220000;
      4859: inst = 32'h10408000;
      4860: inst = 32'hc404b0e;
      4861: inst = 32'h8220000;
      4862: inst = 32'h10408000;
      4863: inst = 32'hc404b20;
      4864: inst = 32'h8220000;
      4865: inst = 32'h10408000;
      4866: inst = 32'hc404b21;
      4867: inst = 32'h8220000;
      4868: inst = 32'h10408000;
      4869: inst = 32'hc404b22;
      4870: inst = 32'h8220000;
      4871: inst = 32'h10408000;
      4872: inst = 32'hc404b23;
      4873: inst = 32'h8220000;
      4874: inst = 32'h10408000;
      4875: inst = 32'hc404b24;
      4876: inst = 32'h8220000;
      4877: inst = 32'h10408000;
      4878: inst = 32'hc404b25;
      4879: inst = 32'h8220000;
      4880: inst = 32'h10408000;
      4881: inst = 32'hc404b26;
      4882: inst = 32'h8220000;
      4883: inst = 32'h10408000;
      4884: inst = 32'hc404b30;
      4885: inst = 32'h8220000;
      4886: inst = 32'h10408000;
      4887: inst = 32'hc404b31;
      4888: inst = 32'h8220000;
      4889: inst = 32'h10408000;
      4890: inst = 32'hc404b32;
      4891: inst = 32'h8220000;
      4892: inst = 32'h10408000;
      4893: inst = 32'hc404b33;
      4894: inst = 32'h8220000;
      4895: inst = 32'h10408000;
      4896: inst = 32'hc404b34;
      4897: inst = 32'h8220000;
      4898: inst = 32'h10408000;
      4899: inst = 32'hc404b35;
      4900: inst = 32'h8220000;
      4901: inst = 32'h10408000;
      4902: inst = 32'hc404b36;
      4903: inst = 32'h8220000;
      4904: inst = 32'h10408000;
      4905: inst = 32'hc404b37;
      4906: inst = 32'h8220000;
      4907: inst = 32'h10408000;
      4908: inst = 32'hc404b38;
      4909: inst = 32'h8220000;
      4910: inst = 32'h10408000;
      4911: inst = 32'hc404b39;
      4912: inst = 32'h8220000;
      4913: inst = 32'h10408000;
      4914: inst = 32'hc404b3a;
      4915: inst = 32'h8220000;
      4916: inst = 32'h10408000;
      4917: inst = 32'hc404b3b;
      4918: inst = 32'h8220000;
      4919: inst = 32'h10408000;
      4920: inst = 32'hc404b64;
      4921: inst = 32'h8220000;
      4922: inst = 32'h10408000;
      4923: inst = 32'hc404b65;
      4924: inst = 32'h8220000;
      4925: inst = 32'h10408000;
      4926: inst = 32'hc404b66;
      4927: inst = 32'h8220000;
      4928: inst = 32'h10408000;
      4929: inst = 32'hc404b67;
      4930: inst = 32'h8220000;
      4931: inst = 32'h10408000;
      4932: inst = 32'hc404b68;
      4933: inst = 32'h8220000;
      4934: inst = 32'h10408000;
      4935: inst = 32'hc404b69;
      4936: inst = 32'h8220000;
      4937: inst = 32'h10408000;
      4938: inst = 32'hc404b6a;
      4939: inst = 32'h8220000;
      4940: inst = 32'h10408000;
      4941: inst = 32'hc404b6b;
      4942: inst = 32'h8220000;
      4943: inst = 32'h10408000;
      4944: inst = 32'hc404b6c;
      4945: inst = 32'h8220000;
      4946: inst = 32'h10408000;
      4947: inst = 32'hc404b6d;
      4948: inst = 32'h8220000;
      4949: inst = 32'h10408000;
      4950: inst = 32'hc404b6e;
      4951: inst = 32'h8220000;
      4952: inst = 32'h10408000;
      4953: inst = 32'hc404b80;
      4954: inst = 32'h8220000;
      4955: inst = 32'h10408000;
      4956: inst = 32'hc404b81;
      4957: inst = 32'h8220000;
      4958: inst = 32'h10408000;
      4959: inst = 32'hc404b82;
      4960: inst = 32'h8220000;
      4961: inst = 32'h10408000;
      4962: inst = 32'hc404b83;
      4963: inst = 32'h8220000;
      4964: inst = 32'h10408000;
      4965: inst = 32'hc404b84;
      4966: inst = 32'h8220000;
      4967: inst = 32'h10408000;
      4968: inst = 32'hc404b85;
      4969: inst = 32'h8220000;
      4970: inst = 32'h10408000;
      4971: inst = 32'hc404b86;
      4972: inst = 32'h8220000;
      4973: inst = 32'h10408000;
      4974: inst = 32'hc404b90;
      4975: inst = 32'h8220000;
      4976: inst = 32'h10408000;
      4977: inst = 32'hc404b91;
      4978: inst = 32'h8220000;
      4979: inst = 32'h10408000;
      4980: inst = 32'hc404b92;
      4981: inst = 32'h8220000;
      4982: inst = 32'h10408000;
      4983: inst = 32'hc404b93;
      4984: inst = 32'h8220000;
      4985: inst = 32'h10408000;
      4986: inst = 32'hc404b94;
      4987: inst = 32'h8220000;
      4988: inst = 32'h10408000;
      4989: inst = 32'hc404b95;
      4990: inst = 32'h8220000;
      4991: inst = 32'h10408000;
      4992: inst = 32'hc404b96;
      4993: inst = 32'h8220000;
      4994: inst = 32'h10408000;
      4995: inst = 32'hc404b97;
      4996: inst = 32'h8220000;
      4997: inst = 32'h10408000;
      4998: inst = 32'hc404b98;
      4999: inst = 32'h8220000;
      5000: inst = 32'h10408000;
      5001: inst = 32'hc404b99;
      5002: inst = 32'h8220000;
      5003: inst = 32'h10408000;
      5004: inst = 32'hc404b9a;
      5005: inst = 32'h8220000;
      5006: inst = 32'h10408000;
      5007: inst = 32'hc404b9b;
      5008: inst = 32'h8220000;
      5009: inst = 32'h10408000;
      5010: inst = 32'hc404bc4;
      5011: inst = 32'h8220000;
      5012: inst = 32'h10408000;
      5013: inst = 32'hc404bc5;
      5014: inst = 32'h8220000;
      5015: inst = 32'h10408000;
      5016: inst = 32'hc404bc6;
      5017: inst = 32'h8220000;
      5018: inst = 32'h10408000;
      5019: inst = 32'hc404bc7;
      5020: inst = 32'h8220000;
      5021: inst = 32'h10408000;
      5022: inst = 32'hc404bc8;
      5023: inst = 32'h8220000;
      5024: inst = 32'h10408000;
      5025: inst = 32'hc404bc9;
      5026: inst = 32'h8220000;
      5027: inst = 32'h10408000;
      5028: inst = 32'hc404bca;
      5029: inst = 32'h8220000;
      5030: inst = 32'h10408000;
      5031: inst = 32'hc404bcb;
      5032: inst = 32'h8220000;
      5033: inst = 32'h10408000;
      5034: inst = 32'hc404bcc;
      5035: inst = 32'h8220000;
      5036: inst = 32'h10408000;
      5037: inst = 32'hc404bcd;
      5038: inst = 32'h8220000;
      5039: inst = 32'h10408000;
      5040: inst = 32'hc404bce;
      5041: inst = 32'h8220000;
      5042: inst = 32'h10408000;
      5043: inst = 32'hc404be0;
      5044: inst = 32'h8220000;
      5045: inst = 32'h10408000;
      5046: inst = 32'hc404be1;
      5047: inst = 32'h8220000;
      5048: inst = 32'h10408000;
      5049: inst = 32'hc404be2;
      5050: inst = 32'h8220000;
      5051: inst = 32'h10408000;
      5052: inst = 32'hc404be3;
      5053: inst = 32'h8220000;
      5054: inst = 32'h10408000;
      5055: inst = 32'hc404be4;
      5056: inst = 32'h8220000;
      5057: inst = 32'h10408000;
      5058: inst = 32'hc404be5;
      5059: inst = 32'h8220000;
      5060: inst = 32'h10408000;
      5061: inst = 32'hc404be6;
      5062: inst = 32'h8220000;
      5063: inst = 32'h10408000;
      5064: inst = 32'hc404bf0;
      5065: inst = 32'h8220000;
      5066: inst = 32'h10408000;
      5067: inst = 32'hc404bf1;
      5068: inst = 32'h8220000;
      5069: inst = 32'h10408000;
      5070: inst = 32'hc404bf2;
      5071: inst = 32'h8220000;
      5072: inst = 32'h10408000;
      5073: inst = 32'hc404bf3;
      5074: inst = 32'h8220000;
      5075: inst = 32'h10408000;
      5076: inst = 32'hc404bf4;
      5077: inst = 32'h8220000;
      5078: inst = 32'h10408000;
      5079: inst = 32'hc404bf5;
      5080: inst = 32'h8220000;
      5081: inst = 32'h10408000;
      5082: inst = 32'hc404bf6;
      5083: inst = 32'h8220000;
      5084: inst = 32'h10408000;
      5085: inst = 32'hc404bf7;
      5086: inst = 32'h8220000;
      5087: inst = 32'h10408000;
      5088: inst = 32'hc404bf8;
      5089: inst = 32'h8220000;
      5090: inst = 32'h10408000;
      5091: inst = 32'hc404bf9;
      5092: inst = 32'h8220000;
      5093: inst = 32'h10408000;
      5094: inst = 32'hc404c26;
      5095: inst = 32'h8220000;
      5096: inst = 32'h10408000;
      5097: inst = 32'hc404c27;
      5098: inst = 32'h8220000;
      5099: inst = 32'h10408000;
      5100: inst = 32'hc404c28;
      5101: inst = 32'h8220000;
      5102: inst = 32'h10408000;
      5103: inst = 32'hc404c29;
      5104: inst = 32'h8220000;
      5105: inst = 32'h10408000;
      5106: inst = 32'hc404c2a;
      5107: inst = 32'h8220000;
      5108: inst = 32'h10408000;
      5109: inst = 32'hc404c2b;
      5110: inst = 32'h8220000;
      5111: inst = 32'h10408000;
      5112: inst = 32'hc404c2c;
      5113: inst = 32'h8220000;
      5114: inst = 32'h10408000;
      5115: inst = 32'hc404c2d;
      5116: inst = 32'h8220000;
      5117: inst = 32'h10408000;
      5118: inst = 32'hc404c2e;
      5119: inst = 32'h8220000;
      5120: inst = 32'h10408000;
      5121: inst = 32'hc404c40;
      5122: inst = 32'h8220000;
      5123: inst = 32'h10408000;
      5124: inst = 32'hc404c41;
      5125: inst = 32'h8220000;
      5126: inst = 32'h10408000;
      5127: inst = 32'hc404c42;
      5128: inst = 32'h8220000;
      5129: inst = 32'h10408000;
      5130: inst = 32'hc404c43;
      5131: inst = 32'h8220000;
      5132: inst = 32'h10408000;
      5133: inst = 32'hc404c44;
      5134: inst = 32'h8220000;
      5135: inst = 32'h10408000;
      5136: inst = 32'hc404c45;
      5137: inst = 32'h8220000;
      5138: inst = 32'h10408000;
      5139: inst = 32'hc404c46;
      5140: inst = 32'h8220000;
      5141: inst = 32'h10408000;
      5142: inst = 32'hc404c4f;
      5143: inst = 32'h8220000;
      5144: inst = 32'h10408000;
      5145: inst = 32'hc404c50;
      5146: inst = 32'h8220000;
      5147: inst = 32'h10408000;
      5148: inst = 32'hc404c51;
      5149: inst = 32'h8220000;
      5150: inst = 32'h10408000;
      5151: inst = 32'hc404c52;
      5152: inst = 32'h8220000;
      5153: inst = 32'h10408000;
      5154: inst = 32'hc404c53;
      5155: inst = 32'h8220000;
      5156: inst = 32'h10408000;
      5157: inst = 32'hc404c54;
      5158: inst = 32'h8220000;
      5159: inst = 32'h10408000;
      5160: inst = 32'hc404c55;
      5161: inst = 32'h8220000;
      5162: inst = 32'h10408000;
      5163: inst = 32'hc404c56;
      5164: inst = 32'h8220000;
      5165: inst = 32'h10408000;
      5166: inst = 32'hc404c57;
      5167: inst = 32'h8220000;
      5168: inst = 32'h10408000;
      5169: inst = 32'hc404c58;
      5170: inst = 32'h8220000;
      5171: inst = 32'h10408000;
      5172: inst = 32'hc404c59;
      5173: inst = 32'h8220000;
      5174: inst = 32'h10408000;
      5175: inst = 32'hc404c5a;
      5176: inst = 32'h8220000;
      5177: inst = 32'h10408000;
      5178: inst = 32'hc404c5b;
      5179: inst = 32'h8220000;
      5180: inst = 32'h10408000;
      5181: inst = 32'hc404c5c;
      5182: inst = 32'h8220000;
      5183: inst = 32'h10408000;
      5184: inst = 32'hc404c5d;
      5185: inst = 32'h8220000;
      5186: inst = 32'h10408000;
      5187: inst = 32'hc404c5e;
      5188: inst = 32'h8220000;
      5189: inst = 32'h10408000;
      5190: inst = 32'hc404c5f;
      5191: inst = 32'h8220000;
      5192: inst = 32'h10408000;
      5193: inst = 32'hc404c60;
      5194: inst = 32'h8220000;
      5195: inst = 32'h10408000;
      5196: inst = 32'hc404c61;
      5197: inst = 32'h8220000;
      5198: inst = 32'h10408000;
      5199: inst = 32'hc404c62;
      5200: inst = 32'h8220000;
      5201: inst = 32'h10408000;
      5202: inst = 32'hc404c63;
      5203: inst = 32'h8220000;
      5204: inst = 32'h10408000;
      5205: inst = 32'hc404c64;
      5206: inst = 32'h8220000;
      5207: inst = 32'h10408000;
      5208: inst = 32'hc404c65;
      5209: inst = 32'h8220000;
      5210: inst = 32'h10408000;
      5211: inst = 32'hc404c66;
      5212: inst = 32'h8220000;
      5213: inst = 32'h10408000;
      5214: inst = 32'hc404c67;
      5215: inst = 32'h8220000;
      5216: inst = 32'h10408000;
      5217: inst = 32'hc404c68;
      5218: inst = 32'h8220000;
      5219: inst = 32'h10408000;
      5220: inst = 32'hc404c69;
      5221: inst = 32'h8220000;
      5222: inst = 32'h10408000;
      5223: inst = 32'hc404c6a;
      5224: inst = 32'h8220000;
      5225: inst = 32'h10408000;
      5226: inst = 32'hc404c6b;
      5227: inst = 32'h8220000;
      5228: inst = 32'h10408000;
      5229: inst = 32'hc404c6c;
      5230: inst = 32'h8220000;
      5231: inst = 32'h10408000;
      5232: inst = 32'hc404c6d;
      5233: inst = 32'h8220000;
      5234: inst = 32'h10408000;
      5235: inst = 32'hc404c6e;
      5236: inst = 32'h8220000;
      5237: inst = 32'h10408000;
      5238: inst = 32'hc404c6f;
      5239: inst = 32'h8220000;
      5240: inst = 32'h10408000;
      5241: inst = 32'hc404c70;
      5242: inst = 32'h8220000;
      5243: inst = 32'h10408000;
      5244: inst = 32'hc404c71;
      5245: inst = 32'h8220000;
      5246: inst = 32'h10408000;
      5247: inst = 32'hc404c72;
      5248: inst = 32'h8220000;
      5249: inst = 32'h10408000;
      5250: inst = 32'hc404c73;
      5251: inst = 32'h8220000;
      5252: inst = 32'h10408000;
      5253: inst = 32'hc404c74;
      5254: inst = 32'h8220000;
      5255: inst = 32'h10408000;
      5256: inst = 32'hc404c75;
      5257: inst = 32'h8220000;
      5258: inst = 32'h10408000;
      5259: inst = 32'hc404c76;
      5260: inst = 32'h8220000;
      5261: inst = 32'h10408000;
      5262: inst = 32'hc404c77;
      5263: inst = 32'h8220000;
      5264: inst = 32'h10408000;
      5265: inst = 32'hc404c78;
      5266: inst = 32'h8220000;
      5267: inst = 32'h10408000;
      5268: inst = 32'hc404c79;
      5269: inst = 32'h8220000;
      5270: inst = 32'h10408000;
      5271: inst = 32'hc404c7a;
      5272: inst = 32'h8220000;
      5273: inst = 32'h10408000;
      5274: inst = 32'hc404c7b;
      5275: inst = 32'h8220000;
      5276: inst = 32'h10408000;
      5277: inst = 32'hc404c7c;
      5278: inst = 32'h8220000;
      5279: inst = 32'h10408000;
      5280: inst = 32'hc404c7d;
      5281: inst = 32'h8220000;
      5282: inst = 32'h10408000;
      5283: inst = 32'hc404c7e;
      5284: inst = 32'h8220000;
      5285: inst = 32'h10408000;
      5286: inst = 32'hc404c7f;
      5287: inst = 32'h8220000;
      5288: inst = 32'h10408000;
      5289: inst = 32'hc404c80;
      5290: inst = 32'h8220000;
      5291: inst = 32'h10408000;
      5292: inst = 32'hc404c81;
      5293: inst = 32'h8220000;
      5294: inst = 32'h10408000;
      5295: inst = 32'hc404c82;
      5296: inst = 32'h8220000;
      5297: inst = 32'h10408000;
      5298: inst = 32'hc404c83;
      5299: inst = 32'h8220000;
      5300: inst = 32'h10408000;
      5301: inst = 32'hc404c84;
      5302: inst = 32'h8220000;
      5303: inst = 32'h10408000;
      5304: inst = 32'hc404c85;
      5305: inst = 32'h8220000;
      5306: inst = 32'h10408000;
      5307: inst = 32'hc404c86;
      5308: inst = 32'h8220000;
      5309: inst = 32'h10408000;
      5310: inst = 32'hc404c87;
      5311: inst = 32'h8220000;
      5312: inst = 32'h10408000;
      5313: inst = 32'hc404c88;
      5314: inst = 32'h8220000;
      5315: inst = 32'h10408000;
      5316: inst = 32'hc404c89;
      5317: inst = 32'h8220000;
      5318: inst = 32'h10408000;
      5319: inst = 32'hc404c8a;
      5320: inst = 32'h8220000;
      5321: inst = 32'h10408000;
      5322: inst = 32'hc404c8b;
      5323: inst = 32'h8220000;
      5324: inst = 32'h10408000;
      5325: inst = 32'hc404c8c;
      5326: inst = 32'h8220000;
      5327: inst = 32'h10408000;
      5328: inst = 32'hc404c8d;
      5329: inst = 32'h8220000;
      5330: inst = 32'h10408000;
      5331: inst = 32'hc404c8e;
      5332: inst = 32'h8220000;
      5333: inst = 32'h10408000;
      5334: inst = 32'hc404ca0;
      5335: inst = 32'h8220000;
      5336: inst = 32'h10408000;
      5337: inst = 32'hc404ca1;
      5338: inst = 32'h8220000;
      5339: inst = 32'h10408000;
      5340: inst = 32'hc404cb7;
      5341: inst = 32'h8220000;
      5342: inst = 32'h10408000;
      5343: inst = 32'hc404cb8;
      5344: inst = 32'h8220000;
      5345: inst = 32'h10408000;
      5346: inst = 32'hc404cb9;
      5347: inst = 32'h8220000;
      5348: inst = 32'h10408000;
      5349: inst = 32'hc404cba;
      5350: inst = 32'h8220000;
      5351: inst = 32'h10408000;
      5352: inst = 32'hc404cbb;
      5353: inst = 32'h8220000;
      5354: inst = 32'h10408000;
      5355: inst = 32'hc404cbc;
      5356: inst = 32'h8220000;
      5357: inst = 32'h10408000;
      5358: inst = 32'hc404cbd;
      5359: inst = 32'h8220000;
      5360: inst = 32'h10408000;
      5361: inst = 32'hc404cbe;
      5362: inst = 32'h8220000;
      5363: inst = 32'h10408000;
      5364: inst = 32'hc404cbf;
      5365: inst = 32'h8220000;
      5366: inst = 32'h10408000;
      5367: inst = 32'hc404cc0;
      5368: inst = 32'h8220000;
      5369: inst = 32'h10408000;
      5370: inst = 32'hc404cc1;
      5371: inst = 32'h8220000;
      5372: inst = 32'h10408000;
      5373: inst = 32'hc404cc2;
      5374: inst = 32'h8220000;
      5375: inst = 32'h10408000;
      5376: inst = 32'hc404cc3;
      5377: inst = 32'h8220000;
      5378: inst = 32'h10408000;
      5379: inst = 32'hc404cc4;
      5380: inst = 32'h8220000;
      5381: inst = 32'h10408000;
      5382: inst = 32'hc404cc5;
      5383: inst = 32'h8220000;
      5384: inst = 32'h10408000;
      5385: inst = 32'hc404cc6;
      5386: inst = 32'h8220000;
      5387: inst = 32'h10408000;
      5388: inst = 32'hc404cc7;
      5389: inst = 32'h8220000;
      5390: inst = 32'h10408000;
      5391: inst = 32'hc404cc8;
      5392: inst = 32'h8220000;
      5393: inst = 32'h10408000;
      5394: inst = 32'hc404cc9;
      5395: inst = 32'h8220000;
      5396: inst = 32'h10408000;
      5397: inst = 32'hc404cca;
      5398: inst = 32'h8220000;
      5399: inst = 32'h10408000;
      5400: inst = 32'hc404ccb;
      5401: inst = 32'h8220000;
      5402: inst = 32'h10408000;
      5403: inst = 32'hc404ccc;
      5404: inst = 32'h8220000;
      5405: inst = 32'h10408000;
      5406: inst = 32'hc404ccd;
      5407: inst = 32'h8220000;
      5408: inst = 32'h10408000;
      5409: inst = 32'hc404cce;
      5410: inst = 32'h8220000;
      5411: inst = 32'h10408000;
      5412: inst = 32'hc404ccf;
      5413: inst = 32'h8220000;
      5414: inst = 32'h10408000;
      5415: inst = 32'hc404cd0;
      5416: inst = 32'h8220000;
      5417: inst = 32'h10408000;
      5418: inst = 32'hc404cd1;
      5419: inst = 32'h8220000;
      5420: inst = 32'h10408000;
      5421: inst = 32'hc404cd2;
      5422: inst = 32'h8220000;
      5423: inst = 32'h10408000;
      5424: inst = 32'hc404cd3;
      5425: inst = 32'h8220000;
      5426: inst = 32'h10408000;
      5427: inst = 32'hc404cd4;
      5428: inst = 32'h8220000;
      5429: inst = 32'h10408000;
      5430: inst = 32'hc404cd5;
      5431: inst = 32'h8220000;
      5432: inst = 32'h10408000;
      5433: inst = 32'hc404cd6;
      5434: inst = 32'h8220000;
      5435: inst = 32'h10408000;
      5436: inst = 32'hc404cd7;
      5437: inst = 32'h8220000;
      5438: inst = 32'h10408000;
      5439: inst = 32'hc404cd8;
      5440: inst = 32'h8220000;
      5441: inst = 32'h10408000;
      5442: inst = 32'hc404cd9;
      5443: inst = 32'h8220000;
      5444: inst = 32'h10408000;
      5445: inst = 32'hc404cda;
      5446: inst = 32'h8220000;
      5447: inst = 32'h10408000;
      5448: inst = 32'hc404cdb;
      5449: inst = 32'h8220000;
      5450: inst = 32'h10408000;
      5451: inst = 32'hc404cdc;
      5452: inst = 32'h8220000;
      5453: inst = 32'h10408000;
      5454: inst = 32'hc404cdd;
      5455: inst = 32'h8220000;
      5456: inst = 32'h10408000;
      5457: inst = 32'hc404cde;
      5458: inst = 32'h8220000;
      5459: inst = 32'h10408000;
      5460: inst = 32'hc404cdf;
      5461: inst = 32'h8220000;
      5462: inst = 32'h10408000;
      5463: inst = 32'hc404ce0;
      5464: inst = 32'h8220000;
      5465: inst = 32'h10408000;
      5466: inst = 32'hc404ce1;
      5467: inst = 32'h8220000;
      5468: inst = 32'h10408000;
      5469: inst = 32'hc404ce2;
      5470: inst = 32'h8220000;
      5471: inst = 32'h10408000;
      5472: inst = 32'hc404ce3;
      5473: inst = 32'h8220000;
      5474: inst = 32'h10408000;
      5475: inst = 32'hc404ce4;
      5476: inst = 32'h8220000;
      5477: inst = 32'h10408000;
      5478: inst = 32'hc404ce5;
      5479: inst = 32'h8220000;
      5480: inst = 32'h10408000;
      5481: inst = 32'hc404ce6;
      5482: inst = 32'h8220000;
      5483: inst = 32'h10408000;
      5484: inst = 32'hc404ce7;
      5485: inst = 32'h8220000;
      5486: inst = 32'h10408000;
      5487: inst = 32'hc404ce8;
      5488: inst = 32'h8220000;
      5489: inst = 32'h10408000;
      5490: inst = 32'hc404ce9;
      5491: inst = 32'h8220000;
      5492: inst = 32'h10408000;
      5493: inst = 32'hc404cea;
      5494: inst = 32'h8220000;
      5495: inst = 32'h10408000;
      5496: inst = 32'hc404ceb;
      5497: inst = 32'h8220000;
      5498: inst = 32'h10408000;
      5499: inst = 32'hc404cec;
      5500: inst = 32'h8220000;
      5501: inst = 32'h10408000;
      5502: inst = 32'hc404ced;
      5503: inst = 32'h8220000;
      5504: inst = 32'h10408000;
      5505: inst = 32'hc404cee;
      5506: inst = 32'h8220000;
      5507: inst = 32'h10408000;
      5508: inst = 32'hc404d17;
      5509: inst = 32'h8220000;
      5510: inst = 32'h10408000;
      5511: inst = 32'hc404d18;
      5512: inst = 32'h8220000;
      5513: inst = 32'h10408000;
      5514: inst = 32'hc404d19;
      5515: inst = 32'h8220000;
      5516: inst = 32'h10408000;
      5517: inst = 32'hc404d1a;
      5518: inst = 32'h8220000;
      5519: inst = 32'h10408000;
      5520: inst = 32'hc404d1b;
      5521: inst = 32'h8220000;
      5522: inst = 32'h10408000;
      5523: inst = 32'hc404d1c;
      5524: inst = 32'h8220000;
      5525: inst = 32'h10408000;
      5526: inst = 32'hc404d1d;
      5527: inst = 32'h8220000;
      5528: inst = 32'h10408000;
      5529: inst = 32'hc404d1e;
      5530: inst = 32'h8220000;
      5531: inst = 32'h10408000;
      5532: inst = 32'hc404d1f;
      5533: inst = 32'h8220000;
      5534: inst = 32'h10408000;
      5535: inst = 32'hc404d20;
      5536: inst = 32'h8220000;
      5537: inst = 32'h10408000;
      5538: inst = 32'hc404d21;
      5539: inst = 32'h8220000;
      5540: inst = 32'h10408000;
      5541: inst = 32'hc404d22;
      5542: inst = 32'h8220000;
      5543: inst = 32'h10408000;
      5544: inst = 32'hc404d23;
      5545: inst = 32'h8220000;
      5546: inst = 32'h10408000;
      5547: inst = 32'hc404d24;
      5548: inst = 32'h8220000;
      5549: inst = 32'h10408000;
      5550: inst = 32'hc404d25;
      5551: inst = 32'h8220000;
      5552: inst = 32'h10408000;
      5553: inst = 32'hc404d26;
      5554: inst = 32'h8220000;
      5555: inst = 32'h10408000;
      5556: inst = 32'hc404d27;
      5557: inst = 32'h8220000;
      5558: inst = 32'h10408000;
      5559: inst = 32'hc404d28;
      5560: inst = 32'h8220000;
      5561: inst = 32'h10408000;
      5562: inst = 32'hc404d29;
      5563: inst = 32'h8220000;
      5564: inst = 32'h10408000;
      5565: inst = 32'hc404d2a;
      5566: inst = 32'h8220000;
      5567: inst = 32'h10408000;
      5568: inst = 32'hc404d2b;
      5569: inst = 32'h8220000;
      5570: inst = 32'h10408000;
      5571: inst = 32'hc404d2c;
      5572: inst = 32'h8220000;
      5573: inst = 32'h10408000;
      5574: inst = 32'hc404d2d;
      5575: inst = 32'h8220000;
      5576: inst = 32'h10408000;
      5577: inst = 32'hc404d2e;
      5578: inst = 32'h8220000;
      5579: inst = 32'h10408000;
      5580: inst = 32'hc404d2f;
      5581: inst = 32'h8220000;
      5582: inst = 32'h10408000;
      5583: inst = 32'hc404d30;
      5584: inst = 32'h8220000;
      5585: inst = 32'h10408000;
      5586: inst = 32'hc404d31;
      5587: inst = 32'h8220000;
      5588: inst = 32'h10408000;
      5589: inst = 32'hc404d32;
      5590: inst = 32'h8220000;
      5591: inst = 32'h10408000;
      5592: inst = 32'hc404d33;
      5593: inst = 32'h8220000;
      5594: inst = 32'h10408000;
      5595: inst = 32'hc404d34;
      5596: inst = 32'h8220000;
      5597: inst = 32'h10408000;
      5598: inst = 32'hc404d35;
      5599: inst = 32'h8220000;
      5600: inst = 32'h10408000;
      5601: inst = 32'hc404d36;
      5602: inst = 32'h8220000;
      5603: inst = 32'h10408000;
      5604: inst = 32'hc404d37;
      5605: inst = 32'h8220000;
      5606: inst = 32'h10408000;
      5607: inst = 32'hc404d38;
      5608: inst = 32'h8220000;
      5609: inst = 32'h10408000;
      5610: inst = 32'hc404d39;
      5611: inst = 32'h8220000;
      5612: inst = 32'h10408000;
      5613: inst = 32'hc404d3a;
      5614: inst = 32'h8220000;
      5615: inst = 32'h10408000;
      5616: inst = 32'hc404d3b;
      5617: inst = 32'h8220000;
      5618: inst = 32'h10408000;
      5619: inst = 32'hc404d3c;
      5620: inst = 32'h8220000;
      5621: inst = 32'h10408000;
      5622: inst = 32'hc404d3d;
      5623: inst = 32'h8220000;
      5624: inst = 32'h10408000;
      5625: inst = 32'hc404d3e;
      5626: inst = 32'h8220000;
      5627: inst = 32'h10408000;
      5628: inst = 32'hc404d3f;
      5629: inst = 32'h8220000;
      5630: inst = 32'h10408000;
      5631: inst = 32'hc404d40;
      5632: inst = 32'h8220000;
      5633: inst = 32'h10408000;
      5634: inst = 32'hc404d41;
      5635: inst = 32'h8220000;
      5636: inst = 32'h10408000;
      5637: inst = 32'hc404d42;
      5638: inst = 32'h8220000;
      5639: inst = 32'h10408000;
      5640: inst = 32'hc404d43;
      5641: inst = 32'h8220000;
      5642: inst = 32'h10408000;
      5643: inst = 32'hc404d44;
      5644: inst = 32'h8220000;
      5645: inst = 32'h10408000;
      5646: inst = 32'hc404d45;
      5647: inst = 32'h8220000;
      5648: inst = 32'h10408000;
      5649: inst = 32'hc404d46;
      5650: inst = 32'h8220000;
      5651: inst = 32'h10408000;
      5652: inst = 32'hc404d47;
      5653: inst = 32'h8220000;
      5654: inst = 32'h10408000;
      5655: inst = 32'hc404d48;
      5656: inst = 32'h8220000;
      5657: inst = 32'h10408000;
      5658: inst = 32'hc404d49;
      5659: inst = 32'h8220000;
      5660: inst = 32'h10408000;
      5661: inst = 32'hc404d4a;
      5662: inst = 32'h8220000;
      5663: inst = 32'h10408000;
      5664: inst = 32'hc404d4b;
      5665: inst = 32'h8220000;
      5666: inst = 32'h10408000;
      5667: inst = 32'hc404d4c;
      5668: inst = 32'h8220000;
      5669: inst = 32'h10408000;
      5670: inst = 32'hc404d4d;
      5671: inst = 32'h8220000;
      5672: inst = 32'h10408000;
      5673: inst = 32'hc404d4e;
      5674: inst = 32'h8220000;
      5675: inst = 32'h10408000;
      5676: inst = 32'hc404d77;
      5677: inst = 32'h8220000;
      5678: inst = 32'h10408000;
      5679: inst = 32'hc404d78;
      5680: inst = 32'h8220000;
      5681: inst = 32'h10408000;
      5682: inst = 32'hc404d79;
      5683: inst = 32'h8220000;
      5684: inst = 32'h10408000;
      5685: inst = 32'hc404d7a;
      5686: inst = 32'h8220000;
      5687: inst = 32'h10408000;
      5688: inst = 32'hc404d7b;
      5689: inst = 32'h8220000;
      5690: inst = 32'h10408000;
      5691: inst = 32'hc404d7c;
      5692: inst = 32'h8220000;
      5693: inst = 32'h10408000;
      5694: inst = 32'hc404d7d;
      5695: inst = 32'h8220000;
      5696: inst = 32'h10408000;
      5697: inst = 32'hc404d7e;
      5698: inst = 32'h8220000;
      5699: inst = 32'h10408000;
      5700: inst = 32'hc404d7f;
      5701: inst = 32'h8220000;
      5702: inst = 32'h10408000;
      5703: inst = 32'hc404d80;
      5704: inst = 32'h8220000;
      5705: inst = 32'h10408000;
      5706: inst = 32'hc404d81;
      5707: inst = 32'h8220000;
      5708: inst = 32'h10408000;
      5709: inst = 32'hc404d82;
      5710: inst = 32'h8220000;
      5711: inst = 32'h10408000;
      5712: inst = 32'hc404d83;
      5713: inst = 32'h8220000;
      5714: inst = 32'h10408000;
      5715: inst = 32'hc404d84;
      5716: inst = 32'h8220000;
      5717: inst = 32'h10408000;
      5718: inst = 32'hc404d85;
      5719: inst = 32'h8220000;
      5720: inst = 32'h10408000;
      5721: inst = 32'hc404d86;
      5722: inst = 32'h8220000;
      5723: inst = 32'h10408000;
      5724: inst = 32'hc404d87;
      5725: inst = 32'h8220000;
      5726: inst = 32'h10408000;
      5727: inst = 32'hc404d88;
      5728: inst = 32'h8220000;
      5729: inst = 32'h10408000;
      5730: inst = 32'hc404d89;
      5731: inst = 32'h8220000;
      5732: inst = 32'h10408000;
      5733: inst = 32'hc404d8a;
      5734: inst = 32'h8220000;
      5735: inst = 32'h10408000;
      5736: inst = 32'hc404d8b;
      5737: inst = 32'h8220000;
      5738: inst = 32'h10408000;
      5739: inst = 32'hc404d8c;
      5740: inst = 32'h8220000;
      5741: inst = 32'h10408000;
      5742: inst = 32'hc404d8d;
      5743: inst = 32'h8220000;
      5744: inst = 32'h10408000;
      5745: inst = 32'hc404d8e;
      5746: inst = 32'h8220000;
      5747: inst = 32'h10408000;
      5748: inst = 32'hc404d8f;
      5749: inst = 32'h8220000;
      5750: inst = 32'h10408000;
      5751: inst = 32'hc404d90;
      5752: inst = 32'h8220000;
      5753: inst = 32'h10408000;
      5754: inst = 32'hc404d91;
      5755: inst = 32'h8220000;
      5756: inst = 32'h10408000;
      5757: inst = 32'hc404d92;
      5758: inst = 32'h8220000;
      5759: inst = 32'h10408000;
      5760: inst = 32'hc404d93;
      5761: inst = 32'h8220000;
      5762: inst = 32'h10408000;
      5763: inst = 32'hc404d94;
      5764: inst = 32'h8220000;
      5765: inst = 32'h10408000;
      5766: inst = 32'hc404d95;
      5767: inst = 32'h8220000;
      5768: inst = 32'h10408000;
      5769: inst = 32'hc404d96;
      5770: inst = 32'h8220000;
      5771: inst = 32'h10408000;
      5772: inst = 32'hc404d97;
      5773: inst = 32'h8220000;
      5774: inst = 32'h10408000;
      5775: inst = 32'hc404d98;
      5776: inst = 32'h8220000;
      5777: inst = 32'h10408000;
      5778: inst = 32'hc404d99;
      5779: inst = 32'h8220000;
      5780: inst = 32'h10408000;
      5781: inst = 32'hc404d9a;
      5782: inst = 32'h8220000;
      5783: inst = 32'h10408000;
      5784: inst = 32'hc404d9b;
      5785: inst = 32'h8220000;
      5786: inst = 32'h10408000;
      5787: inst = 32'hc404d9c;
      5788: inst = 32'h8220000;
      5789: inst = 32'h10408000;
      5790: inst = 32'hc404d9d;
      5791: inst = 32'h8220000;
      5792: inst = 32'h10408000;
      5793: inst = 32'hc404d9e;
      5794: inst = 32'h8220000;
      5795: inst = 32'h10408000;
      5796: inst = 32'hc404d9f;
      5797: inst = 32'h8220000;
      5798: inst = 32'h10408000;
      5799: inst = 32'hc404da0;
      5800: inst = 32'h8220000;
      5801: inst = 32'h10408000;
      5802: inst = 32'hc404da1;
      5803: inst = 32'h8220000;
      5804: inst = 32'h10408000;
      5805: inst = 32'hc404da2;
      5806: inst = 32'h8220000;
      5807: inst = 32'h10408000;
      5808: inst = 32'hc404da3;
      5809: inst = 32'h8220000;
      5810: inst = 32'h10408000;
      5811: inst = 32'hc404da4;
      5812: inst = 32'h8220000;
      5813: inst = 32'h10408000;
      5814: inst = 32'hc404da5;
      5815: inst = 32'h8220000;
      5816: inst = 32'h10408000;
      5817: inst = 32'hc404da6;
      5818: inst = 32'h8220000;
      5819: inst = 32'h10408000;
      5820: inst = 32'hc404da7;
      5821: inst = 32'h8220000;
      5822: inst = 32'h10408000;
      5823: inst = 32'hc404da8;
      5824: inst = 32'h8220000;
      5825: inst = 32'h10408000;
      5826: inst = 32'hc404da9;
      5827: inst = 32'h8220000;
      5828: inst = 32'h10408000;
      5829: inst = 32'hc404daa;
      5830: inst = 32'h8220000;
      5831: inst = 32'h10408000;
      5832: inst = 32'hc404dab;
      5833: inst = 32'h8220000;
      5834: inst = 32'h10408000;
      5835: inst = 32'hc404dac;
      5836: inst = 32'h8220000;
      5837: inst = 32'h10408000;
      5838: inst = 32'hc404dad;
      5839: inst = 32'h8220000;
      5840: inst = 32'h10408000;
      5841: inst = 32'hc404dae;
      5842: inst = 32'h8220000;
      5843: inst = 32'h10408000;
      5844: inst = 32'hc404dd7;
      5845: inst = 32'h8220000;
      5846: inst = 32'h10408000;
      5847: inst = 32'hc404dd8;
      5848: inst = 32'h8220000;
      5849: inst = 32'h10408000;
      5850: inst = 32'hc404dd9;
      5851: inst = 32'h8220000;
      5852: inst = 32'h10408000;
      5853: inst = 32'hc404dda;
      5854: inst = 32'h8220000;
      5855: inst = 32'h10408000;
      5856: inst = 32'hc404ddb;
      5857: inst = 32'h8220000;
      5858: inst = 32'h10408000;
      5859: inst = 32'hc404ddc;
      5860: inst = 32'h8220000;
      5861: inst = 32'h10408000;
      5862: inst = 32'hc404ddd;
      5863: inst = 32'h8220000;
      5864: inst = 32'h10408000;
      5865: inst = 32'hc404dde;
      5866: inst = 32'h8220000;
      5867: inst = 32'h10408000;
      5868: inst = 32'hc404ddf;
      5869: inst = 32'h8220000;
      5870: inst = 32'h10408000;
      5871: inst = 32'hc404de0;
      5872: inst = 32'h8220000;
      5873: inst = 32'h10408000;
      5874: inst = 32'hc404de1;
      5875: inst = 32'h8220000;
      5876: inst = 32'h10408000;
      5877: inst = 32'hc404de2;
      5878: inst = 32'h8220000;
      5879: inst = 32'h10408000;
      5880: inst = 32'hc404de3;
      5881: inst = 32'h8220000;
      5882: inst = 32'h10408000;
      5883: inst = 32'hc404de4;
      5884: inst = 32'h8220000;
      5885: inst = 32'h10408000;
      5886: inst = 32'hc404de5;
      5887: inst = 32'h8220000;
      5888: inst = 32'h10408000;
      5889: inst = 32'hc404de6;
      5890: inst = 32'h8220000;
      5891: inst = 32'h10408000;
      5892: inst = 32'hc404de7;
      5893: inst = 32'h8220000;
      5894: inst = 32'h10408000;
      5895: inst = 32'hc404de8;
      5896: inst = 32'h8220000;
      5897: inst = 32'h10408000;
      5898: inst = 32'hc404de9;
      5899: inst = 32'h8220000;
      5900: inst = 32'h10408000;
      5901: inst = 32'hc404dea;
      5902: inst = 32'h8220000;
      5903: inst = 32'h10408000;
      5904: inst = 32'hc404deb;
      5905: inst = 32'h8220000;
      5906: inst = 32'h10408000;
      5907: inst = 32'hc404dec;
      5908: inst = 32'h8220000;
      5909: inst = 32'h10408000;
      5910: inst = 32'hc404ded;
      5911: inst = 32'h8220000;
      5912: inst = 32'h10408000;
      5913: inst = 32'hc404dee;
      5914: inst = 32'h8220000;
      5915: inst = 32'h10408000;
      5916: inst = 32'hc404def;
      5917: inst = 32'h8220000;
      5918: inst = 32'h10408000;
      5919: inst = 32'hc404df0;
      5920: inst = 32'h8220000;
      5921: inst = 32'h10408000;
      5922: inst = 32'hc404df1;
      5923: inst = 32'h8220000;
      5924: inst = 32'h10408000;
      5925: inst = 32'hc404df2;
      5926: inst = 32'h8220000;
      5927: inst = 32'h10408000;
      5928: inst = 32'hc404df3;
      5929: inst = 32'h8220000;
      5930: inst = 32'h10408000;
      5931: inst = 32'hc404df4;
      5932: inst = 32'h8220000;
      5933: inst = 32'h10408000;
      5934: inst = 32'hc404df5;
      5935: inst = 32'h8220000;
      5936: inst = 32'h10408000;
      5937: inst = 32'hc404df6;
      5938: inst = 32'h8220000;
      5939: inst = 32'h10408000;
      5940: inst = 32'hc404df7;
      5941: inst = 32'h8220000;
      5942: inst = 32'h10408000;
      5943: inst = 32'hc404df8;
      5944: inst = 32'h8220000;
      5945: inst = 32'h10408000;
      5946: inst = 32'hc404df9;
      5947: inst = 32'h8220000;
      5948: inst = 32'h10408000;
      5949: inst = 32'hc404dfa;
      5950: inst = 32'h8220000;
      5951: inst = 32'h10408000;
      5952: inst = 32'hc404dfb;
      5953: inst = 32'h8220000;
      5954: inst = 32'h10408000;
      5955: inst = 32'hc404dfc;
      5956: inst = 32'h8220000;
      5957: inst = 32'h10408000;
      5958: inst = 32'hc404dfd;
      5959: inst = 32'h8220000;
      5960: inst = 32'h10408000;
      5961: inst = 32'hc404dfe;
      5962: inst = 32'h8220000;
      5963: inst = 32'h10408000;
      5964: inst = 32'hc404dff;
      5965: inst = 32'h8220000;
      5966: inst = 32'h10408000;
      5967: inst = 32'hc404e00;
      5968: inst = 32'h8220000;
      5969: inst = 32'h10408000;
      5970: inst = 32'hc404e01;
      5971: inst = 32'h8220000;
      5972: inst = 32'h10408000;
      5973: inst = 32'hc404e02;
      5974: inst = 32'h8220000;
      5975: inst = 32'h10408000;
      5976: inst = 32'hc404e03;
      5977: inst = 32'h8220000;
      5978: inst = 32'h10408000;
      5979: inst = 32'hc404e04;
      5980: inst = 32'h8220000;
      5981: inst = 32'h10408000;
      5982: inst = 32'hc404e05;
      5983: inst = 32'h8220000;
      5984: inst = 32'h10408000;
      5985: inst = 32'hc404e06;
      5986: inst = 32'h8220000;
      5987: inst = 32'h10408000;
      5988: inst = 32'hc404e07;
      5989: inst = 32'h8220000;
      5990: inst = 32'h10408000;
      5991: inst = 32'hc404e08;
      5992: inst = 32'h8220000;
      5993: inst = 32'h10408000;
      5994: inst = 32'hc404e09;
      5995: inst = 32'h8220000;
      5996: inst = 32'h10408000;
      5997: inst = 32'hc404e0a;
      5998: inst = 32'h8220000;
      5999: inst = 32'h10408000;
      6000: inst = 32'hc404e0b;
      6001: inst = 32'h8220000;
      6002: inst = 32'h10408000;
      6003: inst = 32'hc404e0c;
      6004: inst = 32'h8220000;
      6005: inst = 32'h10408000;
      6006: inst = 32'hc404e0d;
      6007: inst = 32'h8220000;
      6008: inst = 32'h10408000;
      6009: inst = 32'hc404e0e;
      6010: inst = 32'h8220000;
      6011: inst = 32'h10408000;
      6012: inst = 32'hc404e37;
      6013: inst = 32'h8220000;
      6014: inst = 32'h10408000;
      6015: inst = 32'hc404e38;
      6016: inst = 32'h8220000;
      6017: inst = 32'h10408000;
      6018: inst = 32'hc404e39;
      6019: inst = 32'h8220000;
      6020: inst = 32'h10408000;
      6021: inst = 32'hc404e3a;
      6022: inst = 32'h8220000;
      6023: inst = 32'h10408000;
      6024: inst = 32'hc404e3b;
      6025: inst = 32'h8220000;
      6026: inst = 32'h10408000;
      6027: inst = 32'hc404e3c;
      6028: inst = 32'h8220000;
      6029: inst = 32'h10408000;
      6030: inst = 32'hc404e3d;
      6031: inst = 32'h8220000;
      6032: inst = 32'h10408000;
      6033: inst = 32'hc404e3e;
      6034: inst = 32'h8220000;
      6035: inst = 32'h10408000;
      6036: inst = 32'hc404e3f;
      6037: inst = 32'h8220000;
      6038: inst = 32'h10408000;
      6039: inst = 32'hc404e40;
      6040: inst = 32'h8220000;
      6041: inst = 32'h10408000;
      6042: inst = 32'hc404e41;
      6043: inst = 32'h8220000;
      6044: inst = 32'h10408000;
      6045: inst = 32'hc404e42;
      6046: inst = 32'h8220000;
      6047: inst = 32'h10408000;
      6048: inst = 32'hc404e43;
      6049: inst = 32'h8220000;
      6050: inst = 32'h10408000;
      6051: inst = 32'hc404e44;
      6052: inst = 32'h8220000;
      6053: inst = 32'h10408000;
      6054: inst = 32'hc404e45;
      6055: inst = 32'h8220000;
      6056: inst = 32'h10408000;
      6057: inst = 32'hc404e46;
      6058: inst = 32'h8220000;
      6059: inst = 32'h10408000;
      6060: inst = 32'hc404e47;
      6061: inst = 32'h8220000;
      6062: inst = 32'h10408000;
      6063: inst = 32'hc404e48;
      6064: inst = 32'h8220000;
      6065: inst = 32'h10408000;
      6066: inst = 32'hc404e49;
      6067: inst = 32'h8220000;
      6068: inst = 32'h10408000;
      6069: inst = 32'hc404e4a;
      6070: inst = 32'h8220000;
      6071: inst = 32'h10408000;
      6072: inst = 32'hc404e4b;
      6073: inst = 32'h8220000;
      6074: inst = 32'h10408000;
      6075: inst = 32'hc404e4c;
      6076: inst = 32'h8220000;
      6077: inst = 32'h10408000;
      6078: inst = 32'hc404e4d;
      6079: inst = 32'h8220000;
      6080: inst = 32'h10408000;
      6081: inst = 32'hc404e4e;
      6082: inst = 32'h8220000;
      6083: inst = 32'h10408000;
      6084: inst = 32'hc404e4f;
      6085: inst = 32'h8220000;
      6086: inst = 32'h10408000;
      6087: inst = 32'hc404e50;
      6088: inst = 32'h8220000;
      6089: inst = 32'h10408000;
      6090: inst = 32'hc404e51;
      6091: inst = 32'h8220000;
      6092: inst = 32'h10408000;
      6093: inst = 32'hc404e52;
      6094: inst = 32'h8220000;
      6095: inst = 32'h10408000;
      6096: inst = 32'hc404e53;
      6097: inst = 32'h8220000;
      6098: inst = 32'h10408000;
      6099: inst = 32'hc404e54;
      6100: inst = 32'h8220000;
      6101: inst = 32'h10408000;
      6102: inst = 32'hc404e55;
      6103: inst = 32'h8220000;
      6104: inst = 32'h10408000;
      6105: inst = 32'hc404e56;
      6106: inst = 32'h8220000;
      6107: inst = 32'h10408000;
      6108: inst = 32'hc404e57;
      6109: inst = 32'h8220000;
      6110: inst = 32'h10408000;
      6111: inst = 32'hc404e58;
      6112: inst = 32'h8220000;
      6113: inst = 32'h10408000;
      6114: inst = 32'hc404e59;
      6115: inst = 32'h8220000;
      6116: inst = 32'h10408000;
      6117: inst = 32'hc404e5a;
      6118: inst = 32'h8220000;
      6119: inst = 32'h10408000;
      6120: inst = 32'hc404e5b;
      6121: inst = 32'h8220000;
      6122: inst = 32'h10408000;
      6123: inst = 32'hc404e5c;
      6124: inst = 32'h8220000;
      6125: inst = 32'h10408000;
      6126: inst = 32'hc404e5d;
      6127: inst = 32'h8220000;
      6128: inst = 32'h10408000;
      6129: inst = 32'hc404e5e;
      6130: inst = 32'h8220000;
      6131: inst = 32'h10408000;
      6132: inst = 32'hc404e5f;
      6133: inst = 32'h8220000;
      6134: inst = 32'h10408000;
      6135: inst = 32'hc404e60;
      6136: inst = 32'h8220000;
      6137: inst = 32'h10408000;
      6138: inst = 32'hc404e61;
      6139: inst = 32'h8220000;
      6140: inst = 32'h10408000;
      6141: inst = 32'hc404e62;
      6142: inst = 32'h8220000;
      6143: inst = 32'h10408000;
      6144: inst = 32'hc404e63;
      6145: inst = 32'h8220000;
      6146: inst = 32'h10408000;
      6147: inst = 32'hc404e64;
      6148: inst = 32'h8220000;
      6149: inst = 32'h10408000;
      6150: inst = 32'hc404e65;
      6151: inst = 32'h8220000;
      6152: inst = 32'h10408000;
      6153: inst = 32'hc404e66;
      6154: inst = 32'h8220000;
      6155: inst = 32'h10408000;
      6156: inst = 32'hc404e67;
      6157: inst = 32'h8220000;
      6158: inst = 32'h10408000;
      6159: inst = 32'hc404e68;
      6160: inst = 32'h8220000;
      6161: inst = 32'h10408000;
      6162: inst = 32'hc404e69;
      6163: inst = 32'h8220000;
      6164: inst = 32'h10408000;
      6165: inst = 32'hc404e6a;
      6166: inst = 32'h8220000;
      6167: inst = 32'h10408000;
      6168: inst = 32'hc404e6b;
      6169: inst = 32'h8220000;
      6170: inst = 32'h10408000;
      6171: inst = 32'hc404e6c;
      6172: inst = 32'h8220000;
      6173: inst = 32'h10408000;
      6174: inst = 32'hc404e6d;
      6175: inst = 32'h8220000;
      6176: inst = 32'h10408000;
      6177: inst = 32'hc404e6e;
      6178: inst = 32'h8220000;
      6179: inst = 32'h10408000;
      6180: inst = 32'hc404e97;
      6181: inst = 32'h8220000;
      6182: inst = 32'h10408000;
      6183: inst = 32'hc404e98;
      6184: inst = 32'h8220000;
      6185: inst = 32'h10408000;
      6186: inst = 32'hc404e99;
      6187: inst = 32'h8220000;
      6188: inst = 32'h10408000;
      6189: inst = 32'hc404e9a;
      6190: inst = 32'h8220000;
      6191: inst = 32'h10408000;
      6192: inst = 32'hc404e9b;
      6193: inst = 32'h8220000;
      6194: inst = 32'h10408000;
      6195: inst = 32'hc404e9c;
      6196: inst = 32'h8220000;
      6197: inst = 32'h10408000;
      6198: inst = 32'hc404e9d;
      6199: inst = 32'h8220000;
      6200: inst = 32'h10408000;
      6201: inst = 32'hc404e9e;
      6202: inst = 32'h8220000;
      6203: inst = 32'h10408000;
      6204: inst = 32'hc404ea8;
      6205: inst = 32'h8220000;
      6206: inst = 32'h10408000;
      6207: inst = 32'hc404ea9;
      6208: inst = 32'h8220000;
      6209: inst = 32'h10408000;
      6210: inst = 32'hc404eaa;
      6211: inst = 32'h8220000;
      6212: inst = 32'h10408000;
      6213: inst = 32'hc404eab;
      6214: inst = 32'h8220000;
      6215: inst = 32'h10408000;
      6216: inst = 32'hc404eac;
      6217: inst = 32'h8220000;
      6218: inst = 32'h10408000;
      6219: inst = 32'hc404ead;
      6220: inst = 32'h8220000;
      6221: inst = 32'h10408000;
      6222: inst = 32'hc404eae;
      6223: inst = 32'h8220000;
      6224: inst = 32'h10408000;
      6225: inst = 32'hc404eaf;
      6226: inst = 32'h8220000;
      6227: inst = 32'h10408000;
      6228: inst = 32'hc404eb0;
      6229: inst = 32'h8220000;
      6230: inst = 32'h10408000;
      6231: inst = 32'hc404eb1;
      6232: inst = 32'h8220000;
      6233: inst = 32'h10408000;
      6234: inst = 32'hc404eb2;
      6235: inst = 32'h8220000;
      6236: inst = 32'h10408000;
      6237: inst = 32'hc404eb3;
      6238: inst = 32'h8220000;
      6239: inst = 32'h10408000;
      6240: inst = 32'hc404eb4;
      6241: inst = 32'h8220000;
      6242: inst = 32'h10408000;
      6243: inst = 32'hc404eb5;
      6244: inst = 32'h8220000;
      6245: inst = 32'h10408000;
      6246: inst = 32'hc404eb6;
      6247: inst = 32'h8220000;
      6248: inst = 32'h10408000;
      6249: inst = 32'hc404eb7;
      6250: inst = 32'h8220000;
      6251: inst = 32'h10408000;
      6252: inst = 32'hc404ec1;
      6253: inst = 32'h8220000;
      6254: inst = 32'h10408000;
      6255: inst = 32'hc404ec2;
      6256: inst = 32'h8220000;
      6257: inst = 32'h10408000;
      6258: inst = 32'hc404ec3;
      6259: inst = 32'h8220000;
      6260: inst = 32'h10408000;
      6261: inst = 32'hc404ec4;
      6262: inst = 32'h8220000;
      6263: inst = 32'h10408000;
      6264: inst = 32'hc404ec5;
      6265: inst = 32'h8220000;
      6266: inst = 32'h10408000;
      6267: inst = 32'hc404ec6;
      6268: inst = 32'h8220000;
      6269: inst = 32'h10408000;
      6270: inst = 32'hc404ec7;
      6271: inst = 32'h8220000;
      6272: inst = 32'h10408000;
      6273: inst = 32'hc404ec8;
      6274: inst = 32'h8220000;
      6275: inst = 32'h10408000;
      6276: inst = 32'hc404ec9;
      6277: inst = 32'h8220000;
      6278: inst = 32'h10408000;
      6279: inst = 32'hc404eca;
      6280: inst = 32'h8220000;
      6281: inst = 32'h10408000;
      6282: inst = 32'hc404ecb;
      6283: inst = 32'h8220000;
      6284: inst = 32'h10408000;
      6285: inst = 32'hc404ecc;
      6286: inst = 32'h8220000;
      6287: inst = 32'h10408000;
      6288: inst = 32'hc404ecd;
      6289: inst = 32'h8220000;
      6290: inst = 32'h10408000;
      6291: inst = 32'hc404ece;
      6292: inst = 32'h8220000;
      6293: inst = 32'h10408000;
      6294: inst = 32'hc404ef7;
      6295: inst = 32'h8220000;
      6296: inst = 32'h10408000;
      6297: inst = 32'hc404ef8;
      6298: inst = 32'h8220000;
      6299: inst = 32'h10408000;
      6300: inst = 32'hc404ef9;
      6301: inst = 32'h8220000;
      6302: inst = 32'h10408000;
      6303: inst = 32'hc404efa;
      6304: inst = 32'h8220000;
      6305: inst = 32'h10408000;
      6306: inst = 32'hc404efb;
      6307: inst = 32'h8220000;
      6308: inst = 32'h10408000;
      6309: inst = 32'hc404efc;
      6310: inst = 32'h8220000;
      6311: inst = 32'h10408000;
      6312: inst = 32'hc404efd;
      6313: inst = 32'h8220000;
      6314: inst = 32'h10408000;
      6315: inst = 32'hc404efe;
      6316: inst = 32'h8220000;
      6317: inst = 32'h10408000;
      6318: inst = 32'hc404f08;
      6319: inst = 32'h8220000;
      6320: inst = 32'h10408000;
      6321: inst = 32'hc404f09;
      6322: inst = 32'h8220000;
      6323: inst = 32'h10408000;
      6324: inst = 32'hc404f0a;
      6325: inst = 32'h8220000;
      6326: inst = 32'h10408000;
      6327: inst = 32'hc404f0b;
      6328: inst = 32'h8220000;
      6329: inst = 32'h10408000;
      6330: inst = 32'hc404f0c;
      6331: inst = 32'h8220000;
      6332: inst = 32'h10408000;
      6333: inst = 32'hc404f0d;
      6334: inst = 32'h8220000;
      6335: inst = 32'h10408000;
      6336: inst = 32'hc404f0e;
      6337: inst = 32'h8220000;
      6338: inst = 32'h10408000;
      6339: inst = 32'hc404f0f;
      6340: inst = 32'h8220000;
      6341: inst = 32'h10408000;
      6342: inst = 32'hc404f10;
      6343: inst = 32'h8220000;
      6344: inst = 32'h10408000;
      6345: inst = 32'hc404f11;
      6346: inst = 32'h8220000;
      6347: inst = 32'h10408000;
      6348: inst = 32'hc404f12;
      6349: inst = 32'h8220000;
      6350: inst = 32'h10408000;
      6351: inst = 32'hc404f13;
      6352: inst = 32'h8220000;
      6353: inst = 32'h10408000;
      6354: inst = 32'hc404f14;
      6355: inst = 32'h8220000;
      6356: inst = 32'h10408000;
      6357: inst = 32'hc404f15;
      6358: inst = 32'h8220000;
      6359: inst = 32'h10408000;
      6360: inst = 32'hc404f16;
      6361: inst = 32'h8220000;
      6362: inst = 32'h10408000;
      6363: inst = 32'hc404f17;
      6364: inst = 32'h8220000;
      6365: inst = 32'h10408000;
      6366: inst = 32'hc404f21;
      6367: inst = 32'h8220000;
      6368: inst = 32'h10408000;
      6369: inst = 32'hc404f22;
      6370: inst = 32'h8220000;
      6371: inst = 32'h10408000;
      6372: inst = 32'hc404f23;
      6373: inst = 32'h8220000;
      6374: inst = 32'h10408000;
      6375: inst = 32'hc404f24;
      6376: inst = 32'h8220000;
      6377: inst = 32'h10408000;
      6378: inst = 32'hc404f25;
      6379: inst = 32'h8220000;
      6380: inst = 32'h10408000;
      6381: inst = 32'hc404f26;
      6382: inst = 32'h8220000;
      6383: inst = 32'h10408000;
      6384: inst = 32'hc404f27;
      6385: inst = 32'h8220000;
      6386: inst = 32'h10408000;
      6387: inst = 32'hc404f28;
      6388: inst = 32'h8220000;
      6389: inst = 32'h10408000;
      6390: inst = 32'hc404f29;
      6391: inst = 32'h8220000;
      6392: inst = 32'h10408000;
      6393: inst = 32'hc404f2a;
      6394: inst = 32'h8220000;
      6395: inst = 32'h10408000;
      6396: inst = 32'hc404f2b;
      6397: inst = 32'h8220000;
      6398: inst = 32'h10408000;
      6399: inst = 32'hc404f2c;
      6400: inst = 32'h8220000;
      6401: inst = 32'h10408000;
      6402: inst = 32'hc404f2d;
      6403: inst = 32'h8220000;
      6404: inst = 32'h10408000;
      6405: inst = 32'hc404f2e;
      6406: inst = 32'h8220000;
      6407: inst = 32'h10408000;
      6408: inst = 32'hc404f57;
      6409: inst = 32'h8220000;
      6410: inst = 32'h10408000;
      6411: inst = 32'hc404f58;
      6412: inst = 32'h8220000;
      6413: inst = 32'h10408000;
      6414: inst = 32'hc404f59;
      6415: inst = 32'h8220000;
      6416: inst = 32'h10408000;
      6417: inst = 32'hc404f5a;
      6418: inst = 32'h8220000;
      6419: inst = 32'h10408000;
      6420: inst = 32'hc404f5b;
      6421: inst = 32'h8220000;
      6422: inst = 32'h10408000;
      6423: inst = 32'hc404f5c;
      6424: inst = 32'h8220000;
      6425: inst = 32'h10408000;
      6426: inst = 32'hc404f5d;
      6427: inst = 32'h8220000;
      6428: inst = 32'h10408000;
      6429: inst = 32'hc404f5e;
      6430: inst = 32'h8220000;
      6431: inst = 32'h10408000;
      6432: inst = 32'hc404f68;
      6433: inst = 32'h8220000;
      6434: inst = 32'h10408000;
      6435: inst = 32'hc404f69;
      6436: inst = 32'h8220000;
      6437: inst = 32'h10408000;
      6438: inst = 32'hc404f6a;
      6439: inst = 32'h8220000;
      6440: inst = 32'h10408000;
      6441: inst = 32'hc404f6b;
      6442: inst = 32'h8220000;
      6443: inst = 32'h10408000;
      6444: inst = 32'hc404f6c;
      6445: inst = 32'h8220000;
      6446: inst = 32'h10408000;
      6447: inst = 32'hc404f6d;
      6448: inst = 32'h8220000;
      6449: inst = 32'h10408000;
      6450: inst = 32'hc404f6e;
      6451: inst = 32'h8220000;
      6452: inst = 32'h10408000;
      6453: inst = 32'hc404f6f;
      6454: inst = 32'h8220000;
      6455: inst = 32'h10408000;
      6456: inst = 32'hc404f70;
      6457: inst = 32'h8220000;
      6458: inst = 32'h10408000;
      6459: inst = 32'hc404f71;
      6460: inst = 32'h8220000;
      6461: inst = 32'h10408000;
      6462: inst = 32'hc404f72;
      6463: inst = 32'h8220000;
      6464: inst = 32'h10408000;
      6465: inst = 32'hc404f73;
      6466: inst = 32'h8220000;
      6467: inst = 32'h10408000;
      6468: inst = 32'hc404f74;
      6469: inst = 32'h8220000;
      6470: inst = 32'h10408000;
      6471: inst = 32'hc404f75;
      6472: inst = 32'h8220000;
      6473: inst = 32'h10408000;
      6474: inst = 32'hc404f76;
      6475: inst = 32'h8220000;
      6476: inst = 32'h10408000;
      6477: inst = 32'hc404f77;
      6478: inst = 32'h8220000;
      6479: inst = 32'h10408000;
      6480: inst = 32'hc404f81;
      6481: inst = 32'h8220000;
      6482: inst = 32'h10408000;
      6483: inst = 32'hc404f82;
      6484: inst = 32'h8220000;
      6485: inst = 32'h10408000;
      6486: inst = 32'hc404f83;
      6487: inst = 32'h8220000;
      6488: inst = 32'h10408000;
      6489: inst = 32'hc404f84;
      6490: inst = 32'h8220000;
      6491: inst = 32'h10408000;
      6492: inst = 32'hc404f85;
      6493: inst = 32'h8220000;
      6494: inst = 32'h10408000;
      6495: inst = 32'hc404f86;
      6496: inst = 32'h8220000;
      6497: inst = 32'h10408000;
      6498: inst = 32'hc404f87;
      6499: inst = 32'h8220000;
      6500: inst = 32'h10408000;
      6501: inst = 32'hc404f88;
      6502: inst = 32'h8220000;
      6503: inst = 32'h10408000;
      6504: inst = 32'hc404f89;
      6505: inst = 32'h8220000;
      6506: inst = 32'h10408000;
      6507: inst = 32'hc404f8a;
      6508: inst = 32'h8220000;
      6509: inst = 32'h10408000;
      6510: inst = 32'hc404f8b;
      6511: inst = 32'h8220000;
      6512: inst = 32'h10408000;
      6513: inst = 32'hc404f8c;
      6514: inst = 32'h8220000;
      6515: inst = 32'h10408000;
      6516: inst = 32'hc404f8d;
      6517: inst = 32'h8220000;
      6518: inst = 32'h10408000;
      6519: inst = 32'hc404f8e;
      6520: inst = 32'h8220000;
      6521: inst = 32'h10408000;
      6522: inst = 32'hc404fb7;
      6523: inst = 32'h8220000;
      6524: inst = 32'h10408000;
      6525: inst = 32'hc404fb8;
      6526: inst = 32'h8220000;
      6527: inst = 32'h10408000;
      6528: inst = 32'hc404fb9;
      6529: inst = 32'h8220000;
      6530: inst = 32'h10408000;
      6531: inst = 32'hc404fba;
      6532: inst = 32'h8220000;
      6533: inst = 32'h10408000;
      6534: inst = 32'hc404fbb;
      6535: inst = 32'h8220000;
      6536: inst = 32'h10408000;
      6537: inst = 32'hc404fbc;
      6538: inst = 32'h8220000;
      6539: inst = 32'h10408000;
      6540: inst = 32'hc404fbd;
      6541: inst = 32'h8220000;
      6542: inst = 32'h10408000;
      6543: inst = 32'hc404fbe;
      6544: inst = 32'h8220000;
      6545: inst = 32'h10408000;
      6546: inst = 32'hc404fc8;
      6547: inst = 32'h8220000;
      6548: inst = 32'h10408000;
      6549: inst = 32'hc404fc9;
      6550: inst = 32'h8220000;
      6551: inst = 32'h10408000;
      6552: inst = 32'hc404fca;
      6553: inst = 32'h8220000;
      6554: inst = 32'h10408000;
      6555: inst = 32'hc404fcb;
      6556: inst = 32'h8220000;
      6557: inst = 32'h10408000;
      6558: inst = 32'hc404fcc;
      6559: inst = 32'h8220000;
      6560: inst = 32'h10408000;
      6561: inst = 32'hc404fcd;
      6562: inst = 32'h8220000;
      6563: inst = 32'h10408000;
      6564: inst = 32'hc404fce;
      6565: inst = 32'h8220000;
      6566: inst = 32'h10408000;
      6567: inst = 32'hc404fcf;
      6568: inst = 32'h8220000;
      6569: inst = 32'h10408000;
      6570: inst = 32'hc404fd0;
      6571: inst = 32'h8220000;
      6572: inst = 32'h10408000;
      6573: inst = 32'hc404fd1;
      6574: inst = 32'h8220000;
      6575: inst = 32'h10408000;
      6576: inst = 32'hc404fd2;
      6577: inst = 32'h8220000;
      6578: inst = 32'h10408000;
      6579: inst = 32'hc404fd3;
      6580: inst = 32'h8220000;
      6581: inst = 32'h10408000;
      6582: inst = 32'hc404fd4;
      6583: inst = 32'h8220000;
      6584: inst = 32'h10408000;
      6585: inst = 32'hc404fd5;
      6586: inst = 32'h8220000;
      6587: inst = 32'h10408000;
      6588: inst = 32'hc404fd6;
      6589: inst = 32'h8220000;
      6590: inst = 32'h10408000;
      6591: inst = 32'hc404fd7;
      6592: inst = 32'h8220000;
      6593: inst = 32'h10408000;
      6594: inst = 32'hc404fe1;
      6595: inst = 32'h8220000;
      6596: inst = 32'h10408000;
      6597: inst = 32'hc404fe2;
      6598: inst = 32'h8220000;
      6599: inst = 32'h10408000;
      6600: inst = 32'hc404fe3;
      6601: inst = 32'h8220000;
      6602: inst = 32'h10408000;
      6603: inst = 32'hc404fe4;
      6604: inst = 32'h8220000;
      6605: inst = 32'h10408000;
      6606: inst = 32'hc404fe5;
      6607: inst = 32'h8220000;
      6608: inst = 32'h10408000;
      6609: inst = 32'hc404fe6;
      6610: inst = 32'h8220000;
      6611: inst = 32'h10408000;
      6612: inst = 32'hc404fe7;
      6613: inst = 32'h8220000;
      6614: inst = 32'h10408000;
      6615: inst = 32'hc404fe8;
      6616: inst = 32'h8220000;
      6617: inst = 32'h10408000;
      6618: inst = 32'hc404fe9;
      6619: inst = 32'h8220000;
      6620: inst = 32'h10408000;
      6621: inst = 32'hc404fea;
      6622: inst = 32'h8220000;
      6623: inst = 32'h10408000;
      6624: inst = 32'hc404feb;
      6625: inst = 32'h8220000;
      6626: inst = 32'h10408000;
      6627: inst = 32'hc404fec;
      6628: inst = 32'h8220000;
      6629: inst = 32'h10408000;
      6630: inst = 32'hc404fed;
      6631: inst = 32'h8220000;
      6632: inst = 32'h10408000;
      6633: inst = 32'hc404fee;
      6634: inst = 32'h8220000;
      6635: inst = 32'h10408000;
      6636: inst = 32'hc405017;
      6637: inst = 32'h8220000;
      6638: inst = 32'h10408000;
      6639: inst = 32'hc405018;
      6640: inst = 32'h8220000;
      6641: inst = 32'h10408000;
      6642: inst = 32'hc405019;
      6643: inst = 32'h8220000;
      6644: inst = 32'h10408000;
      6645: inst = 32'hc40501a;
      6646: inst = 32'h8220000;
      6647: inst = 32'h10408000;
      6648: inst = 32'hc40501b;
      6649: inst = 32'h8220000;
      6650: inst = 32'h10408000;
      6651: inst = 32'hc40501c;
      6652: inst = 32'h8220000;
      6653: inst = 32'h10408000;
      6654: inst = 32'hc40501d;
      6655: inst = 32'h8220000;
      6656: inst = 32'h10408000;
      6657: inst = 32'hc40501e;
      6658: inst = 32'h8220000;
      6659: inst = 32'h10408000;
      6660: inst = 32'hc405028;
      6661: inst = 32'h8220000;
      6662: inst = 32'h10408000;
      6663: inst = 32'hc405029;
      6664: inst = 32'h8220000;
      6665: inst = 32'h10408000;
      6666: inst = 32'hc40502a;
      6667: inst = 32'h8220000;
      6668: inst = 32'h10408000;
      6669: inst = 32'hc40502b;
      6670: inst = 32'h8220000;
      6671: inst = 32'h10408000;
      6672: inst = 32'hc40502c;
      6673: inst = 32'h8220000;
      6674: inst = 32'h10408000;
      6675: inst = 32'hc40502d;
      6676: inst = 32'h8220000;
      6677: inst = 32'h10408000;
      6678: inst = 32'hc40502e;
      6679: inst = 32'h8220000;
      6680: inst = 32'h10408000;
      6681: inst = 32'hc40502f;
      6682: inst = 32'h8220000;
      6683: inst = 32'h10408000;
      6684: inst = 32'hc405030;
      6685: inst = 32'h8220000;
      6686: inst = 32'h10408000;
      6687: inst = 32'hc405031;
      6688: inst = 32'h8220000;
      6689: inst = 32'h10408000;
      6690: inst = 32'hc405032;
      6691: inst = 32'h8220000;
      6692: inst = 32'h10408000;
      6693: inst = 32'hc405033;
      6694: inst = 32'h8220000;
      6695: inst = 32'h10408000;
      6696: inst = 32'hc405034;
      6697: inst = 32'h8220000;
      6698: inst = 32'h10408000;
      6699: inst = 32'hc405035;
      6700: inst = 32'h8220000;
      6701: inst = 32'h10408000;
      6702: inst = 32'hc405036;
      6703: inst = 32'h8220000;
      6704: inst = 32'h10408000;
      6705: inst = 32'hc405037;
      6706: inst = 32'h8220000;
      6707: inst = 32'h10408000;
      6708: inst = 32'hc405041;
      6709: inst = 32'h8220000;
      6710: inst = 32'h10408000;
      6711: inst = 32'hc405042;
      6712: inst = 32'h8220000;
      6713: inst = 32'h10408000;
      6714: inst = 32'hc405043;
      6715: inst = 32'h8220000;
      6716: inst = 32'h10408000;
      6717: inst = 32'hc405044;
      6718: inst = 32'h8220000;
      6719: inst = 32'h10408000;
      6720: inst = 32'hc405045;
      6721: inst = 32'h8220000;
      6722: inst = 32'h10408000;
      6723: inst = 32'hc405046;
      6724: inst = 32'h8220000;
      6725: inst = 32'h10408000;
      6726: inst = 32'hc405047;
      6727: inst = 32'h8220000;
      6728: inst = 32'h10408000;
      6729: inst = 32'hc405048;
      6730: inst = 32'h8220000;
      6731: inst = 32'h10408000;
      6732: inst = 32'hc405049;
      6733: inst = 32'h8220000;
      6734: inst = 32'h10408000;
      6735: inst = 32'hc40504a;
      6736: inst = 32'h8220000;
      6737: inst = 32'h10408000;
      6738: inst = 32'hc40504b;
      6739: inst = 32'h8220000;
      6740: inst = 32'h10408000;
      6741: inst = 32'hc40504c;
      6742: inst = 32'h8220000;
      6743: inst = 32'h10408000;
      6744: inst = 32'hc40504d;
      6745: inst = 32'h8220000;
      6746: inst = 32'h10408000;
      6747: inst = 32'hc40504e;
      6748: inst = 32'h8220000;
      6749: inst = 32'h10408000;
      6750: inst = 32'hc405077;
      6751: inst = 32'h8220000;
      6752: inst = 32'h10408000;
      6753: inst = 32'hc405078;
      6754: inst = 32'h8220000;
      6755: inst = 32'h10408000;
      6756: inst = 32'hc405079;
      6757: inst = 32'h8220000;
      6758: inst = 32'h10408000;
      6759: inst = 32'hc40507a;
      6760: inst = 32'h8220000;
      6761: inst = 32'h10408000;
      6762: inst = 32'hc40507b;
      6763: inst = 32'h8220000;
      6764: inst = 32'h10408000;
      6765: inst = 32'hc40507c;
      6766: inst = 32'h8220000;
      6767: inst = 32'h10408000;
      6768: inst = 32'hc40507d;
      6769: inst = 32'h8220000;
      6770: inst = 32'h10408000;
      6771: inst = 32'hc40507e;
      6772: inst = 32'h8220000;
      6773: inst = 32'h10408000;
      6774: inst = 32'hc405088;
      6775: inst = 32'h8220000;
      6776: inst = 32'h10408000;
      6777: inst = 32'hc405089;
      6778: inst = 32'h8220000;
      6779: inst = 32'h10408000;
      6780: inst = 32'hc40508a;
      6781: inst = 32'h8220000;
      6782: inst = 32'h10408000;
      6783: inst = 32'hc40508b;
      6784: inst = 32'h8220000;
      6785: inst = 32'h10408000;
      6786: inst = 32'hc40508c;
      6787: inst = 32'h8220000;
      6788: inst = 32'h10408000;
      6789: inst = 32'hc40508d;
      6790: inst = 32'h8220000;
      6791: inst = 32'h10408000;
      6792: inst = 32'hc40508e;
      6793: inst = 32'h8220000;
      6794: inst = 32'h10408000;
      6795: inst = 32'hc40508f;
      6796: inst = 32'h8220000;
      6797: inst = 32'h10408000;
      6798: inst = 32'hc405090;
      6799: inst = 32'h8220000;
      6800: inst = 32'h10408000;
      6801: inst = 32'hc405091;
      6802: inst = 32'h8220000;
      6803: inst = 32'h10408000;
      6804: inst = 32'hc405092;
      6805: inst = 32'h8220000;
      6806: inst = 32'h10408000;
      6807: inst = 32'hc405093;
      6808: inst = 32'h8220000;
      6809: inst = 32'h10408000;
      6810: inst = 32'hc405094;
      6811: inst = 32'h8220000;
      6812: inst = 32'h10408000;
      6813: inst = 32'hc405095;
      6814: inst = 32'h8220000;
      6815: inst = 32'h10408000;
      6816: inst = 32'hc405096;
      6817: inst = 32'h8220000;
      6818: inst = 32'h10408000;
      6819: inst = 32'hc405097;
      6820: inst = 32'h8220000;
      6821: inst = 32'h10408000;
      6822: inst = 32'hc4050a1;
      6823: inst = 32'h8220000;
      6824: inst = 32'h10408000;
      6825: inst = 32'hc4050a2;
      6826: inst = 32'h8220000;
      6827: inst = 32'h10408000;
      6828: inst = 32'hc4050a3;
      6829: inst = 32'h8220000;
      6830: inst = 32'h10408000;
      6831: inst = 32'hc4050a4;
      6832: inst = 32'h8220000;
      6833: inst = 32'h10408000;
      6834: inst = 32'hc4050a5;
      6835: inst = 32'h8220000;
      6836: inst = 32'h10408000;
      6837: inst = 32'hc4050a6;
      6838: inst = 32'h8220000;
      6839: inst = 32'h10408000;
      6840: inst = 32'hc4050a7;
      6841: inst = 32'h8220000;
      6842: inst = 32'h10408000;
      6843: inst = 32'hc4050a8;
      6844: inst = 32'h8220000;
      6845: inst = 32'h10408000;
      6846: inst = 32'hc4050a9;
      6847: inst = 32'h8220000;
      6848: inst = 32'h10408000;
      6849: inst = 32'hc4050aa;
      6850: inst = 32'h8220000;
      6851: inst = 32'h10408000;
      6852: inst = 32'hc4050ab;
      6853: inst = 32'h8220000;
      6854: inst = 32'h10408000;
      6855: inst = 32'hc4050ac;
      6856: inst = 32'h8220000;
      6857: inst = 32'h10408000;
      6858: inst = 32'hc4050ad;
      6859: inst = 32'h8220000;
      6860: inst = 32'h10408000;
      6861: inst = 32'hc4050ae;
      6862: inst = 32'h8220000;
      6863: inst = 32'h10408000;
      6864: inst = 32'hc4050d7;
      6865: inst = 32'h8220000;
      6866: inst = 32'h10408000;
      6867: inst = 32'hc4050d8;
      6868: inst = 32'h8220000;
      6869: inst = 32'h10408000;
      6870: inst = 32'hc4050d9;
      6871: inst = 32'h8220000;
      6872: inst = 32'h10408000;
      6873: inst = 32'hc4050da;
      6874: inst = 32'h8220000;
      6875: inst = 32'h10408000;
      6876: inst = 32'hc4050db;
      6877: inst = 32'h8220000;
      6878: inst = 32'h10408000;
      6879: inst = 32'hc4050dc;
      6880: inst = 32'h8220000;
      6881: inst = 32'h10408000;
      6882: inst = 32'hc4050dd;
      6883: inst = 32'h8220000;
      6884: inst = 32'h10408000;
      6885: inst = 32'hc4050de;
      6886: inst = 32'h8220000;
      6887: inst = 32'h10408000;
      6888: inst = 32'hc4050e8;
      6889: inst = 32'h8220000;
      6890: inst = 32'h10408000;
      6891: inst = 32'hc4050e9;
      6892: inst = 32'h8220000;
      6893: inst = 32'h10408000;
      6894: inst = 32'hc4050ea;
      6895: inst = 32'h8220000;
      6896: inst = 32'h10408000;
      6897: inst = 32'hc4050eb;
      6898: inst = 32'h8220000;
      6899: inst = 32'h10408000;
      6900: inst = 32'hc4050ec;
      6901: inst = 32'h8220000;
      6902: inst = 32'h10408000;
      6903: inst = 32'hc4050ed;
      6904: inst = 32'h8220000;
      6905: inst = 32'h10408000;
      6906: inst = 32'hc4050ee;
      6907: inst = 32'h8220000;
      6908: inst = 32'h10408000;
      6909: inst = 32'hc4050ef;
      6910: inst = 32'h8220000;
      6911: inst = 32'h10408000;
      6912: inst = 32'hc4050f0;
      6913: inst = 32'h8220000;
      6914: inst = 32'h10408000;
      6915: inst = 32'hc4050f1;
      6916: inst = 32'h8220000;
      6917: inst = 32'h10408000;
      6918: inst = 32'hc4050f2;
      6919: inst = 32'h8220000;
      6920: inst = 32'h10408000;
      6921: inst = 32'hc4050f3;
      6922: inst = 32'h8220000;
      6923: inst = 32'h10408000;
      6924: inst = 32'hc4050f4;
      6925: inst = 32'h8220000;
      6926: inst = 32'h10408000;
      6927: inst = 32'hc4050f5;
      6928: inst = 32'h8220000;
      6929: inst = 32'h10408000;
      6930: inst = 32'hc4050f6;
      6931: inst = 32'h8220000;
      6932: inst = 32'h10408000;
      6933: inst = 32'hc4050f7;
      6934: inst = 32'h8220000;
      6935: inst = 32'h10408000;
      6936: inst = 32'hc405101;
      6937: inst = 32'h8220000;
      6938: inst = 32'h10408000;
      6939: inst = 32'hc405102;
      6940: inst = 32'h8220000;
      6941: inst = 32'h10408000;
      6942: inst = 32'hc405103;
      6943: inst = 32'h8220000;
      6944: inst = 32'h10408000;
      6945: inst = 32'hc405104;
      6946: inst = 32'h8220000;
      6947: inst = 32'h10408000;
      6948: inst = 32'hc405105;
      6949: inst = 32'h8220000;
      6950: inst = 32'h10408000;
      6951: inst = 32'hc405106;
      6952: inst = 32'h8220000;
      6953: inst = 32'h10408000;
      6954: inst = 32'hc405107;
      6955: inst = 32'h8220000;
      6956: inst = 32'h10408000;
      6957: inst = 32'hc405108;
      6958: inst = 32'h8220000;
      6959: inst = 32'h10408000;
      6960: inst = 32'hc405109;
      6961: inst = 32'h8220000;
      6962: inst = 32'h10408000;
      6963: inst = 32'hc40510a;
      6964: inst = 32'h8220000;
      6965: inst = 32'h10408000;
      6966: inst = 32'hc40510b;
      6967: inst = 32'h8220000;
      6968: inst = 32'h10408000;
      6969: inst = 32'hc40510c;
      6970: inst = 32'h8220000;
      6971: inst = 32'h10408000;
      6972: inst = 32'hc40510d;
      6973: inst = 32'h8220000;
      6974: inst = 32'h10408000;
      6975: inst = 32'hc40510e;
      6976: inst = 32'h8220000;
      6977: inst = 32'h10408000;
      6978: inst = 32'hc405137;
      6979: inst = 32'h8220000;
      6980: inst = 32'h10408000;
      6981: inst = 32'hc405138;
      6982: inst = 32'h8220000;
      6983: inst = 32'h10408000;
      6984: inst = 32'hc405139;
      6985: inst = 32'h8220000;
      6986: inst = 32'h10408000;
      6987: inst = 32'hc40513a;
      6988: inst = 32'h8220000;
      6989: inst = 32'h10408000;
      6990: inst = 32'hc40513b;
      6991: inst = 32'h8220000;
      6992: inst = 32'h10408000;
      6993: inst = 32'hc40513c;
      6994: inst = 32'h8220000;
      6995: inst = 32'h10408000;
      6996: inst = 32'hc40513d;
      6997: inst = 32'h8220000;
      6998: inst = 32'h10408000;
      6999: inst = 32'hc40513e;
      7000: inst = 32'h8220000;
      7001: inst = 32'h10408000;
      7002: inst = 32'hc405148;
      7003: inst = 32'h8220000;
      7004: inst = 32'h10408000;
      7005: inst = 32'hc405149;
      7006: inst = 32'h8220000;
      7007: inst = 32'h10408000;
      7008: inst = 32'hc40514a;
      7009: inst = 32'h8220000;
      7010: inst = 32'h10408000;
      7011: inst = 32'hc40514b;
      7012: inst = 32'h8220000;
      7013: inst = 32'h10408000;
      7014: inst = 32'hc40514c;
      7015: inst = 32'h8220000;
      7016: inst = 32'h10408000;
      7017: inst = 32'hc40514d;
      7018: inst = 32'h8220000;
      7019: inst = 32'h10408000;
      7020: inst = 32'hc40514e;
      7021: inst = 32'h8220000;
      7022: inst = 32'h10408000;
      7023: inst = 32'hc40514f;
      7024: inst = 32'h8220000;
      7025: inst = 32'h10408000;
      7026: inst = 32'hc405150;
      7027: inst = 32'h8220000;
      7028: inst = 32'h10408000;
      7029: inst = 32'hc405151;
      7030: inst = 32'h8220000;
      7031: inst = 32'h10408000;
      7032: inst = 32'hc405152;
      7033: inst = 32'h8220000;
      7034: inst = 32'h10408000;
      7035: inst = 32'hc405153;
      7036: inst = 32'h8220000;
      7037: inst = 32'h10408000;
      7038: inst = 32'hc405154;
      7039: inst = 32'h8220000;
      7040: inst = 32'h10408000;
      7041: inst = 32'hc405155;
      7042: inst = 32'h8220000;
      7043: inst = 32'h10408000;
      7044: inst = 32'hc405156;
      7045: inst = 32'h8220000;
      7046: inst = 32'h10408000;
      7047: inst = 32'hc405157;
      7048: inst = 32'h8220000;
      7049: inst = 32'h10408000;
      7050: inst = 32'hc405161;
      7051: inst = 32'h8220000;
      7052: inst = 32'h10408000;
      7053: inst = 32'hc405162;
      7054: inst = 32'h8220000;
      7055: inst = 32'h10408000;
      7056: inst = 32'hc405163;
      7057: inst = 32'h8220000;
      7058: inst = 32'h10408000;
      7059: inst = 32'hc405164;
      7060: inst = 32'h8220000;
      7061: inst = 32'h10408000;
      7062: inst = 32'hc405165;
      7063: inst = 32'h8220000;
      7064: inst = 32'h10408000;
      7065: inst = 32'hc405166;
      7066: inst = 32'h8220000;
      7067: inst = 32'h10408000;
      7068: inst = 32'hc405167;
      7069: inst = 32'h8220000;
      7070: inst = 32'h10408000;
      7071: inst = 32'hc405168;
      7072: inst = 32'h8220000;
      7073: inst = 32'h10408000;
      7074: inst = 32'hc405169;
      7075: inst = 32'h8220000;
      7076: inst = 32'h10408000;
      7077: inst = 32'hc40516a;
      7078: inst = 32'h8220000;
      7079: inst = 32'h10408000;
      7080: inst = 32'hc40516b;
      7081: inst = 32'h8220000;
      7082: inst = 32'h10408000;
      7083: inst = 32'hc40516c;
      7084: inst = 32'h8220000;
      7085: inst = 32'h10408000;
      7086: inst = 32'hc40516d;
      7087: inst = 32'h8220000;
      7088: inst = 32'h10408000;
      7089: inst = 32'hc40516e;
      7090: inst = 32'h8220000;
      7091: inst = 32'h10408000;
      7092: inst = 32'hc405197;
      7093: inst = 32'h8220000;
      7094: inst = 32'h10408000;
      7095: inst = 32'hc405198;
      7096: inst = 32'h8220000;
      7097: inst = 32'h10408000;
      7098: inst = 32'hc405199;
      7099: inst = 32'h8220000;
      7100: inst = 32'h10408000;
      7101: inst = 32'hc40519a;
      7102: inst = 32'h8220000;
      7103: inst = 32'h10408000;
      7104: inst = 32'hc40519b;
      7105: inst = 32'h8220000;
      7106: inst = 32'h10408000;
      7107: inst = 32'hc40519c;
      7108: inst = 32'h8220000;
      7109: inst = 32'h10408000;
      7110: inst = 32'hc40519d;
      7111: inst = 32'h8220000;
      7112: inst = 32'h10408000;
      7113: inst = 32'hc4051aa;
      7114: inst = 32'h8220000;
      7115: inst = 32'h10408000;
      7116: inst = 32'hc4051ab;
      7117: inst = 32'h8220000;
      7118: inst = 32'h10408000;
      7119: inst = 32'hc4051ac;
      7120: inst = 32'h8220000;
      7121: inst = 32'h10408000;
      7122: inst = 32'hc4051ad;
      7123: inst = 32'h8220000;
      7124: inst = 32'h10408000;
      7125: inst = 32'hc4051ae;
      7126: inst = 32'h8220000;
      7127: inst = 32'h10408000;
      7128: inst = 32'hc4051af;
      7129: inst = 32'h8220000;
      7130: inst = 32'h10408000;
      7131: inst = 32'hc4051b0;
      7132: inst = 32'h8220000;
      7133: inst = 32'h10408000;
      7134: inst = 32'hc4051b1;
      7135: inst = 32'h8220000;
      7136: inst = 32'h10408000;
      7137: inst = 32'hc4051b2;
      7138: inst = 32'h8220000;
      7139: inst = 32'h10408000;
      7140: inst = 32'hc4051b3;
      7141: inst = 32'h8220000;
      7142: inst = 32'h10408000;
      7143: inst = 32'hc4051b4;
      7144: inst = 32'h8220000;
      7145: inst = 32'h10408000;
      7146: inst = 32'hc4051b5;
      7147: inst = 32'h8220000;
      7148: inst = 32'h10408000;
      7149: inst = 32'hc4051c2;
      7150: inst = 32'h8220000;
      7151: inst = 32'h10408000;
      7152: inst = 32'hc4051c3;
      7153: inst = 32'h8220000;
      7154: inst = 32'h10408000;
      7155: inst = 32'hc4051c4;
      7156: inst = 32'h8220000;
      7157: inst = 32'h10408000;
      7158: inst = 32'hc4051c5;
      7159: inst = 32'h8220000;
      7160: inst = 32'h10408000;
      7161: inst = 32'hc4051c6;
      7162: inst = 32'h8220000;
      7163: inst = 32'h10408000;
      7164: inst = 32'hc4051c7;
      7165: inst = 32'h8220000;
      7166: inst = 32'h10408000;
      7167: inst = 32'hc4051c8;
      7168: inst = 32'h8220000;
      7169: inst = 32'h10408000;
      7170: inst = 32'hc4051c9;
      7171: inst = 32'h8220000;
      7172: inst = 32'h10408000;
      7173: inst = 32'hc4051ca;
      7174: inst = 32'h8220000;
      7175: inst = 32'h10408000;
      7176: inst = 32'hc4051cb;
      7177: inst = 32'h8220000;
      7178: inst = 32'h10408000;
      7179: inst = 32'hc4051cc;
      7180: inst = 32'h8220000;
      7181: inst = 32'h10408000;
      7182: inst = 32'hc4051cd;
      7183: inst = 32'h8220000;
      7184: inst = 32'h10408000;
      7185: inst = 32'hc4051ce;
      7186: inst = 32'h8220000;
      7187: inst = 32'h10408000;
      7188: inst = 32'hc4051f7;
      7189: inst = 32'h8220000;
      7190: inst = 32'h10408000;
      7191: inst = 32'hc4051f8;
      7192: inst = 32'h8220000;
      7193: inst = 32'h10408000;
      7194: inst = 32'hc4051f9;
      7195: inst = 32'h8220000;
      7196: inst = 32'h10408000;
      7197: inst = 32'hc4051fa;
      7198: inst = 32'h8220000;
      7199: inst = 32'h10408000;
      7200: inst = 32'hc4051fb;
      7201: inst = 32'h8220000;
      7202: inst = 32'h10408000;
      7203: inst = 32'hc4051fc;
      7204: inst = 32'h8220000;
      7205: inst = 32'h10408000;
      7206: inst = 32'hc40520a;
      7207: inst = 32'h8220000;
      7208: inst = 32'h10408000;
      7209: inst = 32'hc40520b;
      7210: inst = 32'h8220000;
      7211: inst = 32'h10408000;
      7212: inst = 32'hc40520c;
      7213: inst = 32'h8220000;
      7214: inst = 32'h10408000;
      7215: inst = 32'hc40520d;
      7216: inst = 32'h8220000;
      7217: inst = 32'h10408000;
      7218: inst = 32'hc40520e;
      7219: inst = 32'h8220000;
      7220: inst = 32'h10408000;
      7221: inst = 32'hc40520f;
      7222: inst = 32'h8220000;
      7223: inst = 32'h10408000;
      7224: inst = 32'hc405210;
      7225: inst = 32'h8220000;
      7226: inst = 32'h10408000;
      7227: inst = 32'hc405211;
      7228: inst = 32'h8220000;
      7229: inst = 32'h10408000;
      7230: inst = 32'hc405212;
      7231: inst = 32'h8220000;
      7232: inst = 32'h10408000;
      7233: inst = 32'hc405213;
      7234: inst = 32'h8220000;
      7235: inst = 32'h10408000;
      7236: inst = 32'hc405214;
      7237: inst = 32'h8220000;
      7238: inst = 32'h10408000;
      7239: inst = 32'hc405215;
      7240: inst = 32'h8220000;
      7241: inst = 32'h10408000;
      7242: inst = 32'hc405223;
      7243: inst = 32'h8220000;
      7244: inst = 32'h10408000;
      7245: inst = 32'hc405224;
      7246: inst = 32'h8220000;
      7247: inst = 32'h10408000;
      7248: inst = 32'hc405225;
      7249: inst = 32'h8220000;
      7250: inst = 32'h10408000;
      7251: inst = 32'hc405226;
      7252: inst = 32'h8220000;
      7253: inst = 32'h10408000;
      7254: inst = 32'hc405227;
      7255: inst = 32'h8220000;
      7256: inst = 32'h10408000;
      7257: inst = 32'hc405228;
      7258: inst = 32'h8220000;
      7259: inst = 32'h10408000;
      7260: inst = 32'hc405229;
      7261: inst = 32'h8220000;
      7262: inst = 32'h10408000;
      7263: inst = 32'hc40522a;
      7264: inst = 32'h8220000;
      7265: inst = 32'h10408000;
      7266: inst = 32'hc40522b;
      7267: inst = 32'h8220000;
      7268: inst = 32'h10408000;
      7269: inst = 32'hc40522c;
      7270: inst = 32'h8220000;
      7271: inst = 32'h10408000;
      7272: inst = 32'hc40522d;
      7273: inst = 32'h8220000;
      7274: inst = 32'h10408000;
      7275: inst = 32'hc40522e;
      7276: inst = 32'h8220000;
      7277: inst = 32'h10408000;
      7278: inst = 32'hc405257;
      7279: inst = 32'h8220000;
      7280: inst = 32'h10408000;
      7281: inst = 32'hc405258;
      7282: inst = 32'h8220000;
      7283: inst = 32'h10408000;
      7284: inst = 32'hc405259;
      7285: inst = 32'h8220000;
      7286: inst = 32'h10408000;
      7287: inst = 32'hc40525a;
      7288: inst = 32'h8220000;
      7289: inst = 32'h10408000;
      7290: inst = 32'hc40525b;
      7291: inst = 32'h8220000;
      7292: inst = 32'h10408000;
      7293: inst = 32'hc40526a;
      7294: inst = 32'h8220000;
      7295: inst = 32'h10408000;
      7296: inst = 32'hc40526b;
      7297: inst = 32'h8220000;
      7298: inst = 32'h10408000;
      7299: inst = 32'hc40526c;
      7300: inst = 32'h8220000;
      7301: inst = 32'h10408000;
      7302: inst = 32'hc40526d;
      7303: inst = 32'h8220000;
      7304: inst = 32'h10408000;
      7305: inst = 32'hc40526e;
      7306: inst = 32'h8220000;
      7307: inst = 32'h10408000;
      7308: inst = 32'hc40526f;
      7309: inst = 32'h8220000;
      7310: inst = 32'h10408000;
      7311: inst = 32'hc405270;
      7312: inst = 32'h8220000;
      7313: inst = 32'h10408000;
      7314: inst = 32'hc405271;
      7315: inst = 32'h8220000;
      7316: inst = 32'h10408000;
      7317: inst = 32'hc405272;
      7318: inst = 32'h8220000;
      7319: inst = 32'h10408000;
      7320: inst = 32'hc405273;
      7321: inst = 32'h8220000;
      7322: inst = 32'h10408000;
      7323: inst = 32'hc405274;
      7324: inst = 32'h8220000;
      7325: inst = 32'h10408000;
      7326: inst = 32'hc405275;
      7327: inst = 32'h8220000;
      7328: inst = 32'h10408000;
      7329: inst = 32'hc405284;
      7330: inst = 32'h8220000;
      7331: inst = 32'h10408000;
      7332: inst = 32'hc405285;
      7333: inst = 32'h8220000;
      7334: inst = 32'h10408000;
      7335: inst = 32'hc405286;
      7336: inst = 32'h8220000;
      7337: inst = 32'h10408000;
      7338: inst = 32'hc405287;
      7339: inst = 32'h8220000;
      7340: inst = 32'h10408000;
      7341: inst = 32'hc405288;
      7342: inst = 32'h8220000;
      7343: inst = 32'h10408000;
      7344: inst = 32'hc405289;
      7345: inst = 32'h8220000;
      7346: inst = 32'h10408000;
      7347: inst = 32'hc40528a;
      7348: inst = 32'h8220000;
      7349: inst = 32'h10408000;
      7350: inst = 32'hc40528b;
      7351: inst = 32'h8220000;
      7352: inst = 32'h10408000;
      7353: inst = 32'hc40528c;
      7354: inst = 32'h8220000;
      7355: inst = 32'h10408000;
      7356: inst = 32'hc40528d;
      7357: inst = 32'h8220000;
      7358: inst = 32'h10408000;
      7359: inst = 32'hc40528e;
      7360: inst = 32'h8220000;
      7361: inst = 32'h10408000;
      7362: inst = 32'hc4052b7;
      7363: inst = 32'h8220000;
      7364: inst = 32'h10408000;
      7365: inst = 32'hc4052b8;
      7366: inst = 32'h8220000;
      7367: inst = 32'h10408000;
      7368: inst = 32'hc4052b9;
      7369: inst = 32'h8220000;
      7370: inst = 32'h10408000;
      7371: inst = 32'hc4052ba;
      7372: inst = 32'h8220000;
      7373: inst = 32'h10408000;
      7374: inst = 32'hc4052bb;
      7375: inst = 32'h8220000;
      7376: inst = 32'h10408000;
      7377: inst = 32'hc4052ca;
      7378: inst = 32'h8220000;
      7379: inst = 32'h10408000;
      7380: inst = 32'hc4052cb;
      7381: inst = 32'h8220000;
      7382: inst = 32'h10408000;
      7383: inst = 32'hc4052cc;
      7384: inst = 32'h8220000;
      7385: inst = 32'h10408000;
      7386: inst = 32'hc4052cd;
      7387: inst = 32'h8220000;
      7388: inst = 32'h10408000;
      7389: inst = 32'hc4052ce;
      7390: inst = 32'h8220000;
      7391: inst = 32'h10408000;
      7392: inst = 32'hc4052cf;
      7393: inst = 32'h8220000;
      7394: inst = 32'h10408000;
      7395: inst = 32'hc4052d0;
      7396: inst = 32'h8220000;
      7397: inst = 32'h10408000;
      7398: inst = 32'hc4052d1;
      7399: inst = 32'h8220000;
      7400: inst = 32'h10408000;
      7401: inst = 32'hc4052d2;
      7402: inst = 32'h8220000;
      7403: inst = 32'h10408000;
      7404: inst = 32'hc4052d3;
      7405: inst = 32'h8220000;
      7406: inst = 32'h10408000;
      7407: inst = 32'hc4052d4;
      7408: inst = 32'h8220000;
      7409: inst = 32'h10408000;
      7410: inst = 32'hc4052d5;
      7411: inst = 32'h8220000;
      7412: inst = 32'h10408000;
      7413: inst = 32'hc4052e4;
      7414: inst = 32'h8220000;
      7415: inst = 32'h10408000;
      7416: inst = 32'hc4052e5;
      7417: inst = 32'h8220000;
      7418: inst = 32'h10408000;
      7419: inst = 32'hc4052e6;
      7420: inst = 32'h8220000;
      7421: inst = 32'h10408000;
      7422: inst = 32'hc4052e7;
      7423: inst = 32'h8220000;
      7424: inst = 32'h10408000;
      7425: inst = 32'hc4052e8;
      7426: inst = 32'h8220000;
      7427: inst = 32'h10408000;
      7428: inst = 32'hc4052e9;
      7429: inst = 32'h8220000;
      7430: inst = 32'h10408000;
      7431: inst = 32'hc4052ea;
      7432: inst = 32'h8220000;
      7433: inst = 32'h10408000;
      7434: inst = 32'hc4052eb;
      7435: inst = 32'h8220000;
      7436: inst = 32'h10408000;
      7437: inst = 32'hc4052ec;
      7438: inst = 32'h8220000;
      7439: inst = 32'h10408000;
      7440: inst = 32'hc4052ed;
      7441: inst = 32'h8220000;
      7442: inst = 32'h10408000;
      7443: inst = 32'hc4052ee;
      7444: inst = 32'h8220000;
      7445: inst = 32'hc2094b2;
      7446: inst = 32'h10408000;
      7447: inst = 32'hc403feb;
      7448: inst = 32'h8220000;
      7449: inst = 32'h10408000;
      7450: inst = 32'hc40404b;
      7451: inst = 32'h8220000;
      7452: inst = 32'h10408000;
      7453: inst = 32'hc4040ab;
      7454: inst = 32'h8220000;
      7455: inst = 32'h10408000;
      7456: inst = 32'hc40410b;
      7457: inst = 32'h8220000;
      7458: inst = 32'h10408000;
      7459: inst = 32'hc40416b;
      7460: inst = 32'h8220000;
      7461: inst = 32'h10408000;
      7462: inst = 32'hc4041cb;
      7463: inst = 32'h8220000;
      7464: inst = 32'h10408000;
      7465: inst = 32'hc40422b;
      7466: inst = 32'h8220000;
      7467: inst = 32'h10408000;
      7468: inst = 32'hc40428b;
      7469: inst = 32'h8220000;
      7470: inst = 32'hc20b596;
      7471: inst = 32'h10408000;
      7472: inst = 32'hc4041da;
      7473: inst = 32'h8220000;
      7474: inst = 32'h10408000;
      7475: inst = 32'hc4041db;
      7476: inst = 32'h8220000;
      7477: inst = 32'h10408000;
      7478: inst = 32'hc4041dc;
      7479: inst = 32'h8220000;
      7480: inst = 32'h10408000;
      7481: inst = 32'hc4041dd;
      7482: inst = 32'h8220000;
      7483: inst = 32'h10408000;
      7484: inst = 32'hc4041de;
      7485: inst = 32'h8220000;
      7486: inst = 32'h10408000;
      7487: inst = 32'hc4041df;
      7488: inst = 32'h8220000;
      7489: inst = 32'h10408000;
      7490: inst = 32'hc4041e0;
      7491: inst = 32'h8220000;
      7492: inst = 32'h10408000;
      7493: inst = 32'hc4041e1;
      7494: inst = 32'h8220000;
      7495: inst = 32'h10408000;
      7496: inst = 32'hc4041e2;
      7497: inst = 32'h8220000;
      7498: inst = 32'h10408000;
      7499: inst = 32'hc4041e3;
      7500: inst = 32'h8220000;
      7501: inst = 32'h10408000;
      7502: inst = 32'hc4041e4;
      7503: inst = 32'h8220000;
      7504: inst = 32'h10408000;
      7505: inst = 32'hc4041e5;
      7506: inst = 32'h8220000;
      7507: inst = 32'h10408000;
      7508: inst = 32'hc4041e6;
      7509: inst = 32'h8220000;
      7510: inst = 32'h10408000;
      7511: inst = 32'hc4041e7;
      7512: inst = 32'h8220000;
      7513: inst = 32'h10408000;
      7514: inst = 32'hc4041e8;
      7515: inst = 32'h8220000;
      7516: inst = 32'h10408000;
      7517: inst = 32'hc4041e9;
      7518: inst = 32'h8220000;
      7519: inst = 32'h10408000;
      7520: inst = 32'hc4041ea;
      7521: inst = 32'h8220000;
      7522: inst = 32'h10408000;
      7523: inst = 32'hc4041eb;
      7524: inst = 32'h8220000;
      7525: inst = 32'h10408000;
      7526: inst = 32'hc4041ec;
      7527: inst = 32'h8220000;
      7528: inst = 32'h10408000;
      7529: inst = 32'hc4041ed;
      7530: inst = 32'h8220000;
      7531: inst = 32'h10408000;
      7532: inst = 32'hc4041ee;
      7533: inst = 32'h8220000;
      7534: inst = 32'h10408000;
      7535: inst = 32'hc4041ef;
      7536: inst = 32'h8220000;
      7537: inst = 32'h10408000;
      7538: inst = 32'hc4041f0;
      7539: inst = 32'h8220000;
      7540: inst = 32'h10408000;
      7541: inst = 32'hc4041f1;
      7542: inst = 32'h8220000;
      7543: inst = 32'h10408000;
      7544: inst = 32'hc4041f2;
      7545: inst = 32'h8220000;
      7546: inst = 32'h10408000;
      7547: inst = 32'hc4041f3;
      7548: inst = 32'h8220000;
      7549: inst = 32'h10408000;
      7550: inst = 32'hc4041f4;
      7551: inst = 32'h8220000;
      7552: inst = 32'h10408000;
      7553: inst = 32'hc4041f5;
      7554: inst = 32'h8220000;
      7555: inst = 32'h10408000;
      7556: inst = 32'hc4041f6;
      7557: inst = 32'h8220000;
      7558: inst = 32'h10408000;
      7559: inst = 32'hc4041f7;
      7560: inst = 32'h8220000;
      7561: inst = 32'h10408000;
      7562: inst = 32'hc4041f8;
      7563: inst = 32'h8220000;
      7564: inst = 32'h10408000;
      7565: inst = 32'hc4041f9;
      7566: inst = 32'h8220000;
      7567: inst = 32'h10408000;
      7568: inst = 32'hc4041fa;
      7569: inst = 32'h8220000;
      7570: inst = 32'h10408000;
      7571: inst = 32'hc4041fb;
      7572: inst = 32'h8220000;
      7573: inst = 32'h10408000;
      7574: inst = 32'hc4041fc;
      7575: inst = 32'h8220000;
      7576: inst = 32'h10408000;
      7577: inst = 32'hc4041fd;
      7578: inst = 32'h8220000;
      7579: inst = 32'h10408000;
      7580: inst = 32'hc4041fe;
      7581: inst = 32'h8220000;
      7582: inst = 32'h10408000;
      7583: inst = 32'hc4041ff;
      7584: inst = 32'h8220000;
      7585: inst = 32'h10408000;
      7586: inst = 32'hc404200;
      7587: inst = 32'h8220000;
      7588: inst = 32'h10408000;
      7589: inst = 32'hc404201;
      7590: inst = 32'h8220000;
      7591: inst = 32'h10408000;
      7592: inst = 32'hc404202;
      7593: inst = 32'h8220000;
      7594: inst = 32'h10408000;
      7595: inst = 32'hc404203;
      7596: inst = 32'h8220000;
      7597: inst = 32'h10408000;
      7598: inst = 32'hc404204;
      7599: inst = 32'h8220000;
      7600: inst = 32'h10408000;
      7601: inst = 32'hc404205;
      7602: inst = 32'h8220000;
      7603: inst = 32'h10408000;
      7604: inst = 32'hc404bfa;
      7605: inst = 32'h8220000;
      7606: inst = 32'h10408000;
      7607: inst = 32'hc404bfb;
      7608: inst = 32'h8220000;
      7609: inst = 32'h10408000;
      7610: inst = 32'hc404bfc;
      7611: inst = 32'h8220000;
      7612: inst = 32'h10408000;
      7613: inst = 32'hc404bfd;
      7614: inst = 32'h8220000;
      7615: inst = 32'h10408000;
      7616: inst = 32'hc404bfe;
      7617: inst = 32'h8220000;
      7618: inst = 32'h10408000;
      7619: inst = 32'hc404bff;
      7620: inst = 32'h8220000;
      7621: inst = 32'h10408000;
      7622: inst = 32'hc404c00;
      7623: inst = 32'h8220000;
      7624: inst = 32'h10408000;
      7625: inst = 32'hc404c01;
      7626: inst = 32'h8220000;
      7627: inst = 32'h10408000;
      7628: inst = 32'hc404c02;
      7629: inst = 32'h8220000;
      7630: inst = 32'h10408000;
      7631: inst = 32'hc404c03;
      7632: inst = 32'h8220000;
      7633: inst = 32'h10408000;
      7634: inst = 32'hc404c04;
      7635: inst = 32'h8220000;
      7636: inst = 32'h10408000;
      7637: inst = 32'hc404c05;
      7638: inst = 32'h8220000;
      7639: inst = 32'h10408000;
      7640: inst = 32'hc404c06;
      7641: inst = 32'h8220000;
      7642: inst = 32'h10408000;
      7643: inst = 32'hc404c07;
      7644: inst = 32'h8220000;
      7645: inst = 32'h10408000;
      7646: inst = 32'hc404c08;
      7647: inst = 32'h8220000;
      7648: inst = 32'h10408000;
      7649: inst = 32'hc404c09;
      7650: inst = 32'h8220000;
      7651: inst = 32'h10408000;
      7652: inst = 32'hc404c0a;
      7653: inst = 32'h8220000;
      7654: inst = 32'h10408000;
      7655: inst = 32'hc404c0b;
      7656: inst = 32'h8220000;
      7657: inst = 32'h10408000;
      7658: inst = 32'hc404c0c;
      7659: inst = 32'h8220000;
      7660: inst = 32'h10408000;
      7661: inst = 32'hc404c0d;
      7662: inst = 32'h8220000;
      7663: inst = 32'h10408000;
      7664: inst = 32'hc404c0e;
      7665: inst = 32'h8220000;
      7666: inst = 32'h10408000;
      7667: inst = 32'hc404c0f;
      7668: inst = 32'h8220000;
      7669: inst = 32'h10408000;
      7670: inst = 32'hc404c10;
      7671: inst = 32'h8220000;
      7672: inst = 32'h10408000;
      7673: inst = 32'hc404c11;
      7674: inst = 32'h8220000;
      7675: inst = 32'h10408000;
      7676: inst = 32'hc404c12;
      7677: inst = 32'h8220000;
      7678: inst = 32'h10408000;
      7679: inst = 32'hc404c13;
      7680: inst = 32'h8220000;
      7681: inst = 32'h10408000;
      7682: inst = 32'hc404c14;
      7683: inst = 32'h8220000;
      7684: inst = 32'h10408000;
      7685: inst = 32'hc404c15;
      7686: inst = 32'h8220000;
      7687: inst = 32'h10408000;
      7688: inst = 32'hc404c16;
      7689: inst = 32'h8220000;
      7690: inst = 32'h10408000;
      7691: inst = 32'hc404c17;
      7692: inst = 32'h8220000;
      7693: inst = 32'h10408000;
      7694: inst = 32'hc404c18;
      7695: inst = 32'h8220000;
      7696: inst = 32'h10408000;
      7697: inst = 32'hc404c19;
      7698: inst = 32'h8220000;
      7699: inst = 32'h10408000;
      7700: inst = 32'hc404c1a;
      7701: inst = 32'h8220000;
      7702: inst = 32'h10408000;
      7703: inst = 32'hc404c1b;
      7704: inst = 32'h8220000;
      7705: inst = 32'h10408000;
      7706: inst = 32'hc404c1c;
      7707: inst = 32'h8220000;
      7708: inst = 32'h10408000;
      7709: inst = 32'hc404c1d;
      7710: inst = 32'h8220000;
      7711: inst = 32'h10408000;
      7712: inst = 32'hc404c1e;
      7713: inst = 32'h8220000;
      7714: inst = 32'h10408000;
      7715: inst = 32'hc404c1f;
      7716: inst = 32'h8220000;
      7717: inst = 32'h10408000;
      7718: inst = 32'hc404c20;
      7719: inst = 32'h8220000;
      7720: inst = 32'h10408000;
      7721: inst = 32'hc404c21;
      7722: inst = 32'h8220000;
      7723: inst = 32'h10408000;
      7724: inst = 32'hc404c22;
      7725: inst = 32'h8220000;
      7726: inst = 32'h10408000;
      7727: inst = 32'hc404c23;
      7728: inst = 32'h8220000;
      7729: inst = 32'h10408000;
      7730: inst = 32'hc404c24;
      7731: inst = 32'h8220000;
      7732: inst = 32'h10408000;
      7733: inst = 32'hc404c25;
      7734: inst = 32'h8220000;
      7735: inst = 32'hc20ffff;
      7736: inst = 32'h10408000;
      7737: inst = 32'hc40423c;
      7738: inst = 32'h8220000;
      7739: inst = 32'h10408000;
      7740: inst = 32'hc40423d;
      7741: inst = 32'h8220000;
      7742: inst = 32'h10408000;
      7743: inst = 32'hc40423e;
      7744: inst = 32'h8220000;
      7745: inst = 32'h10408000;
      7746: inst = 32'hc40423f;
      7747: inst = 32'h8220000;
      7748: inst = 32'h10408000;
      7749: inst = 32'hc404240;
      7750: inst = 32'h8220000;
      7751: inst = 32'h10408000;
      7752: inst = 32'hc404241;
      7753: inst = 32'h8220000;
      7754: inst = 32'h10408000;
      7755: inst = 32'hc404242;
      7756: inst = 32'h8220000;
      7757: inst = 32'h10408000;
      7758: inst = 32'hc404243;
      7759: inst = 32'h8220000;
      7760: inst = 32'h10408000;
      7761: inst = 32'hc404244;
      7762: inst = 32'h8220000;
      7763: inst = 32'h10408000;
      7764: inst = 32'hc404245;
      7765: inst = 32'h8220000;
      7766: inst = 32'h10408000;
      7767: inst = 32'hc404246;
      7768: inst = 32'h8220000;
      7769: inst = 32'h10408000;
      7770: inst = 32'hc404247;
      7771: inst = 32'h8220000;
      7772: inst = 32'h10408000;
      7773: inst = 32'hc404248;
      7774: inst = 32'h8220000;
      7775: inst = 32'h10408000;
      7776: inst = 32'hc404249;
      7777: inst = 32'h8220000;
      7778: inst = 32'h10408000;
      7779: inst = 32'hc40424a;
      7780: inst = 32'h8220000;
      7781: inst = 32'h10408000;
      7782: inst = 32'hc40424b;
      7783: inst = 32'h8220000;
      7784: inst = 32'h10408000;
      7785: inst = 32'hc40424c;
      7786: inst = 32'h8220000;
      7787: inst = 32'h10408000;
      7788: inst = 32'hc40424d;
      7789: inst = 32'h8220000;
      7790: inst = 32'h10408000;
      7791: inst = 32'hc40424e;
      7792: inst = 32'h8220000;
      7793: inst = 32'h10408000;
      7794: inst = 32'hc40424f;
      7795: inst = 32'h8220000;
      7796: inst = 32'h10408000;
      7797: inst = 32'hc404250;
      7798: inst = 32'h8220000;
      7799: inst = 32'h10408000;
      7800: inst = 32'hc404251;
      7801: inst = 32'h8220000;
      7802: inst = 32'h10408000;
      7803: inst = 32'hc404252;
      7804: inst = 32'h8220000;
      7805: inst = 32'h10408000;
      7806: inst = 32'hc404253;
      7807: inst = 32'h8220000;
      7808: inst = 32'h10408000;
      7809: inst = 32'hc404254;
      7810: inst = 32'h8220000;
      7811: inst = 32'h10408000;
      7812: inst = 32'hc404255;
      7813: inst = 32'h8220000;
      7814: inst = 32'h10408000;
      7815: inst = 32'hc404256;
      7816: inst = 32'h8220000;
      7817: inst = 32'h10408000;
      7818: inst = 32'hc404257;
      7819: inst = 32'h8220000;
      7820: inst = 32'h10408000;
      7821: inst = 32'hc404258;
      7822: inst = 32'h8220000;
      7823: inst = 32'h10408000;
      7824: inst = 32'hc404259;
      7825: inst = 32'h8220000;
      7826: inst = 32'h10408000;
      7827: inst = 32'hc40425a;
      7828: inst = 32'h8220000;
      7829: inst = 32'h10408000;
      7830: inst = 32'hc40425b;
      7831: inst = 32'h8220000;
      7832: inst = 32'h10408000;
      7833: inst = 32'hc40425c;
      7834: inst = 32'h8220000;
      7835: inst = 32'h10408000;
      7836: inst = 32'hc40425d;
      7837: inst = 32'h8220000;
      7838: inst = 32'h10408000;
      7839: inst = 32'hc40425e;
      7840: inst = 32'h8220000;
      7841: inst = 32'h10408000;
      7842: inst = 32'hc40425f;
      7843: inst = 32'h8220000;
      7844: inst = 32'h10408000;
      7845: inst = 32'hc404260;
      7846: inst = 32'h8220000;
      7847: inst = 32'h10408000;
      7848: inst = 32'hc404261;
      7849: inst = 32'h8220000;
      7850: inst = 32'h10408000;
      7851: inst = 32'hc404262;
      7852: inst = 32'h8220000;
      7853: inst = 32'h10408000;
      7854: inst = 32'hc404263;
      7855: inst = 32'h8220000;
      7856: inst = 32'h10408000;
      7857: inst = 32'hc40429c;
      7858: inst = 32'h8220000;
      7859: inst = 32'h10408000;
      7860: inst = 32'hc40429d;
      7861: inst = 32'h8220000;
      7862: inst = 32'h10408000;
      7863: inst = 32'hc40429e;
      7864: inst = 32'h8220000;
      7865: inst = 32'h10408000;
      7866: inst = 32'hc40429f;
      7867: inst = 32'h8220000;
      7868: inst = 32'h10408000;
      7869: inst = 32'hc4042a0;
      7870: inst = 32'h8220000;
      7871: inst = 32'h10408000;
      7872: inst = 32'hc4042a1;
      7873: inst = 32'h8220000;
      7874: inst = 32'h10408000;
      7875: inst = 32'hc4042a2;
      7876: inst = 32'h8220000;
      7877: inst = 32'h10408000;
      7878: inst = 32'hc4042a3;
      7879: inst = 32'h8220000;
      7880: inst = 32'h10408000;
      7881: inst = 32'hc4042a4;
      7882: inst = 32'h8220000;
      7883: inst = 32'h10408000;
      7884: inst = 32'hc4042a5;
      7885: inst = 32'h8220000;
      7886: inst = 32'h10408000;
      7887: inst = 32'hc4042a6;
      7888: inst = 32'h8220000;
      7889: inst = 32'h10408000;
      7890: inst = 32'hc4042a7;
      7891: inst = 32'h8220000;
      7892: inst = 32'h10408000;
      7893: inst = 32'hc4042a8;
      7894: inst = 32'h8220000;
      7895: inst = 32'h10408000;
      7896: inst = 32'hc4042a9;
      7897: inst = 32'h8220000;
      7898: inst = 32'h10408000;
      7899: inst = 32'hc4042aa;
      7900: inst = 32'h8220000;
      7901: inst = 32'h10408000;
      7902: inst = 32'hc4042ab;
      7903: inst = 32'h8220000;
      7904: inst = 32'h10408000;
      7905: inst = 32'hc4042ac;
      7906: inst = 32'h8220000;
      7907: inst = 32'h10408000;
      7908: inst = 32'hc4042ad;
      7909: inst = 32'h8220000;
      7910: inst = 32'h10408000;
      7911: inst = 32'hc4042ae;
      7912: inst = 32'h8220000;
      7913: inst = 32'h10408000;
      7914: inst = 32'hc4042af;
      7915: inst = 32'h8220000;
      7916: inst = 32'h10408000;
      7917: inst = 32'hc4042b0;
      7918: inst = 32'h8220000;
      7919: inst = 32'h10408000;
      7920: inst = 32'hc4042b1;
      7921: inst = 32'h8220000;
      7922: inst = 32'h10408000;
      7923: inst = 32'hc4042b2;
      7924: inst = 32'h8220000;
      7925: inst = 32'h10408000;
      7926: inst = 32'hc4042b3;
      7927: inst = 32'h8220000;
      7928: inst = 32'h10408000;
      7929: inst = 32'hc4042b4;
      7930: inst = 32'h8220000;
      7931: inst = 32'h10408000;
      7932: inst = 32'hc4042b5;
      7933: inst = 32'h8220000;
      7934: inst = 32'h10408000;
      7935: inst = 32'hc4042b6;
      7936: inst = 32'h8220000;
      7937: inst = 32'h10408000;
      7938: inst = 32'hc4042b7;
      7939: inst = 32'h8220000;
      7940: inst = 32'h10408000;
      7941: inst = 32'hc4042b8;
      7942: inst = 32'h8220000;
      7943: inst = 32'h10408000;
      7944: inst = 32'hc4042b9;
      7945: inst = 32'h8220000;
      7946: inst = 32'h10408000;
      7947: inst = 32'hc4042ba;
      7948: inst = 32'h8220000;
      7949: inst = 32'h10408000;
      7950: inst = 32'hc4042bb;
      7951: inst = 32'h8220000;
      7952: inst = 32'h10408000;
      7953: inst = 32'hc4042bc;
      7954: inst = 32'h8220000;
      7955: inst = 32'h10408000;
      7956: inst = 32'hc4042bd;
      7957: inst = 32'h8220000;
      7958: inst = 32'h10408000;
      7959: inst = 32'hc4042be;
      7960: inst = 32'h8220000;
      7961: inst = 32'h10408000;
      7962: inst = 32'hc4042bf;
      7963: inst = 32'h8220000;
      7964: inst = 32'h10408000;
      7965: inst = 32'hc4042c0;
      7966: inst = 32'h8220000;
      7967: inst = 32'h10408000;
      7968: inst = 32'hc4042c1;
      7969: inst = 32'h8220000;
      7970: inst = 32'h10408000;
      7971: inst = 32'hc4042c2;
      7972: inst = 32'h8220000;
      7973: inst = 32'h10408000;
      7974: inst = 32'hc4042c3;
      7975: inst = 32'h8220000;
      7976: inst = 32'h10408000;
      7977: inst = 32'hc4042fc;
      7978: inst = 32'h8220000;
      7979: inst = 32'h10408000;
      7980: inst = 32'hc4042fd;
      7981: inst = 32'h8220000;
      7982: inst = 32'h10408000;
      7983: inst = 32'hc4042fe;
      7984: inst = 32'h8220000;
      7985: inst = 32'h10408000;
      7986: inst = 32'hc4042ff;
      7987: inst = 32'h8220000;
      7988: inst = 32'h10408000;
      7989: inst = 32'hc404300;
      7990: inst = 32'h8220000;
      7991: inst = 32'h10408000;
      7992: inst = 32'hc404301;
      7993: inst = 32'h8220000;
      7994: inst = 32'h10408000;
      7995: inst = 32'hc404302;
      7996: inst = 32'h8220000;
      7997: inst = 32'h10408000;
      7998: inst = 32'hc404303;
      7999: inst = 32'h8220000;
      8000: inst = 32'h10408000;
      8001: inst = 32'hc404304;
      8002: inst = 32'h8220000;
      8003: inst = 32'h10408000;
      8004: inst = 32'hc404305;
      8005: inst = 32'h8220000;
      8006: inst = 32'h10408000;
      8007: inst = 32'hc404306;
      8008: inst = 32'h8220000;
      8009: inst = 32'h10408000;
      8010: inst = 32'hc404307;
      8011: inst = 32'h8220000;
      8012: inst = 32'h10408000;
      8013: inst = 32'hc404308;
      8014: inst = 32'h8220000;
      8015: inst = 32'h10408000;
      8016: inst = 32'hc404309;
      8017: inst = 32'h8220000;
      8018: inst = 32'h10408000;
      8019: inst = 32'hc40430a;
      8020: inst = 32'h8220000;
      8021: inst = 32'h10408000;
      8022: inst = 32'hc40430b;
      8023: inst = 32'h8220000;
      8024: inst = 32'h10408000;
      8025: inst = 32'hc40430c;
      8026: inst = 32'h8220000;
      8027: inst = 32'h10408000;
      8028: inst = 32'hc40430d;
      8029: inst = 32'h8220000;
      8030: inst = 32'h10408000;
      8031: inst = 32'hc40430e;
      8032: inst = 32'h8220000;
      8033: inst = 32'h10408000;
      8034: inst = 32'hc40430f;
      8035: inst = 32'h8220000;
      8036: inst = 32'h10408000;
      8037: inst = 32'hc404310;
      8038: inst = 32'h8220000;
      8039: inst = 32'h10408000;
      8040: inst = 32'hc404311;
      8041: inst = 32'h8220000;
      8042: inst = 32'h10408000;
      8043: inst = 32'hc404312;
      8044: inst = 32'h8220000;
      8045: inst = 32'h10408000;
      8046: inst = 32'hc404313;
      8047: inst = 32'h8220000;
      8048: inst = 32'h10408000;
      8049: inst = 32'hc404314;
      8050: inst = 32'h8220000;
      8051: inst = 32'h10408000;
      8052: inst = 32'hc404315;
      8053: inst = 32'h8220000;
      8054: inst = 32'h10408000;
      8055: inst = 32'hc404316;
      8056: inst = 32'h8220000;
      8057: inst = 32'h10408000;
      8058: inst = 32'hc404317;
      8059: inst = 32'h8220000;
      8060: inst = 32'h10408000;
      8061: inst = 32'hc404318;
      8062: inst = 32'h8220000;
      8063: inst = 32'h10408000;
      8064: inst = 32'hc404319;
      8065: inst = 32'h8220000;
      8066: inst = 32'h10408000;
      8067: inst = 32'hc40431a;
      8068: inst = 32'h8220000;
      8069: inst = 32'h10408000;
      8070: inst = 32'hc40431b;
      8071: inst = 32'h8220000;
      8072: inst = 32'h10408000;
      8073: inst = 32'hc40431c;
      8074: inst = 32'h8220000;
      8075: inst = 32'h10408000;
      8076: inst = 32'hc40431d;
      8077: inst = 32'h8220000;
      8078: inst = 32'h10408000;
      8079: inst = 32'hc40431e;
      8080: inst = 32'h8220000;
      8081: inst = 32'h10408000;
      8082: inst = 32'hc40431f;
      8083: inst = 32'h8220000;
      8084: inst = 32'h10408000;
      8085: inst = 32'hc404320;
      8086: inst = 32'h8220000;
      8087: inst = 32'h10408000;
      8088: inst = 32'hc404321;
      8089: inst = 32'h8220000;
      8090: inst = 32'h10408000;
      8091: inst = 32'hc404322;
      8092: inst = 32'h8220000;
      8093: inst = 32'h10408000;
      8094: inst = 32'hc404323;
      8095: inst = 32'h8220000;
      8096: inst = 32'h10408000;
      8097: inst = 32'hc40435c;
      8098: inst = 32'h8220000;
      8099: inst = 32'h10408000;
      8100: inst = 32'hc40435d;
      8101: inst = 32'h8220000;
      8102: inst = 32'h10408000;
      8103: inst = 32'hc40435e;
      8104: inst = 32'h8220000;
      8105: inst = 32'h10408000;
      8106: inst = 32'hc40435f;
      8107: inst = 32'h8220000;
      8108: inst = 32'h10408000;
      8109: inst = 32'hc404360;
      8110: inst = 32'h8220000;
      8111: inst = 32'h10408000;
      8112: inst = 32'hc404361;
      8113: inst = 32'h8220000;
      8114: inst = 32'h10408000;
      8115: inst = 32'hc404362;
      8116: inst = 32'h8220000;
      8117: inst = 32'h10408000;
      8118: inst = 32'hc404363;
      8119: inst = 32'h8220000;
      8120: inst = 32'h10408000;
      8121: inst = 32'hc404364;
      8122: inst = 32'h8220000;
      8123: inst = 32'h10408000;
      8124: inst = 32'hc404365;
      8125: inst = 32'h8220000;
      8126: inst = 32'h10408000;
      8127: inst = 32'hc404366;
      8128: inst = 32'h8220000;
      8129: inst = 32'h10408000;
      8130: inst = 32'hc404367;
      8131: inst = 32'h8220000;
      8132: inst = 32'h10408000;
      8133: inst = 32'hc404368;
      8134: inst = 32'h8220000;
      8135: inst = 32'h10408000;
      8136: inst = 32'hc404369;
      8137: inst = 32'h8220000;
      8138: inst = 32'h10408000;
      8139: inst = 32'hc40436a;
      8140: inst = 32'h8220000;
      8141: inst = 32'h10408000;
      8142: inst = 32'hc40436b;
      8143: inst = 32'h8220000;
      8144: inst = 32'h10408000;
      8145: inst = 32'hc40436c;
      8146: inst = 32'h8220000;
      8147: inst = 32'h10408000;
      8148: inst = 32'hc40436d;
      8149: inst = 32'h8220000;
      8150: inst = 32'h10408000;
      8151: inst = 32'hc40436e;
      8152: inst = 32'h8220000;
      8153: inst = 32'h10408000;
      8154: inst = 32'hc40436f;
      8155: inst = 32'h8220000;
      8156: inst = 32'h10408000;
      8157: inst = 32'hc404370;
      8158: inst = 32'h8220000;
      8159: inst = 32'h10408000;
      8160: inst = 32'hc404371;
      8161: inst = 32'h8220000;
      8162: inst = 32'h10408000;
      8163: inst = 32'hc404372;
      8164: inst = 32'h8220000;
      8165: inst = 32'h10408000;
      8166: inst = 32'hc404373;
      8167: inst = 32'h8220000;
      8168: inst = 32'h10408000;
      8169: inst = 32'hc404374;
      8170: inst = 32'h8220000;
      8171: inst = 32'h10408000;
      8172: inst = 32'hc404375;
      8173: inst = 32'h8220000;
      8174: inst = 32'h10408000;
      8175: inst = 32'hc404376;
      8176: inst = 32'h8220000;
      8177: inst = 32'h10408000;
      8178: inst = 32'hc404377;
      8179: inst = 32'h8220000;
      8180: inst = 32'h10408000;
      8181: inst = 32'hc404378;
      8182: inst = 32'h8220000;
      8183: inst = 32'h10408000;
      8184: inst = 32'hc404379;
      8185: inst = 32'h8220000;
      8186: inst = 32'h10408000;
      8187: inst = 32'hc40437a;
      8188: inst = 32'h8220000;
      8189: inst = 32'h10408000;
      8190: inst = 32'hc40437b;
      8191: inst = 32'h8220000;
      8192: inst = 32'h10408000;
      8193: inst = 32'hc40437c;
      8194: inst = 32'h8220000;
      8195: inst = 32'h10408000;
      8196: inst = 32'hc40437d;
      8197: inst = 32'h8220000;
      8198: inst = 32'h10408000;
      8199: inst = 32'hc40437e;
      8200: inst = 32'h8220000;
      8201: inst = 32'h10408000;
      8202: inst = 32'hc40437f;
      8203: inst = 32'h8220000;
      8204: inst = 32'h10408000;
      8205: inst = 32'hc404380;
      8206: inst = 32'h8220000;
      8207: inst = 32'h10408000;
      8208: inst = 32'hc404381;
      8209: inst = 32'h8220000;
      8210: inst = 32'h10408000;
      8211: inst = 32'hc404382;
      8212: inst = 32'h8220000;
      8213: inst = 32'h10408000;
      8214: inst = 32'hc404383;
      8215: inst = 32'h8220000;
      8216: inst = 32'h10408000;
      8217: inst = 32'hc4043bc;
      8218: inst = 32'h8220000;
      8219: inst = 32'h10408000;
      8220: inst = 32'hc4043bd;
      8221: inst = 32'h8220000;
      8222: inst = 32'h10408000;
      8223: inst = 32'hc4043be;
      8224: inst = 32'h8220000;
      8225: inst = 32'h10408000;
      8226: inst = 32'hc4043bf;
      8227: inst = 32'h8220000;
      8228: inst = 32'h10408000;
      8229: inst = 32'hc4043c0;
      8230: inst = 32'h8220000;
      8231: inst = 32'h10408000;
      8232: inst = 32'hc4043c1;
      8233: inst = 32'h8220000;
      8234: inst = 32'h10408000;
      8235: inst = 32'hc4043c2;
      8236: inst = 32'h8220000;
      8237: inst = 32'h10408000;
      8238: inst = 32'hc4043c3;
      8239: inst = 32'h8220000;
      8240: inst = 32'h10408000;
      8241: inst = 32'hc4043c4;
      8242: inst = 32'h8220000;
      8243: inst = 32'h10408000;
      8244: inst = 32'hc4043c5;
      8245: inst = 32'h8220000;
      8246: inst = 32'h10408000;
      8247: inst = 32'hc4043c6;
      8248: inst = 32'h8220000;
      8249: inst = 32'h10408000;
      8250: inst = 32'hc4043c7;
      8251: inst = 32'h8220000;
      8252: inst = 32'h10408000;
      8253: inst = 32'hc4043c8;
      8254: inst = 32'h8220000;
      8255: inst = 32'h10408000;
      8256: inst = 32'hc4043c9;
      8257: inst = 32'h8220000;
      8258: inst = 32'h10408000;
      8259: inst = 32'hc4043ca;
      8260: inst = 32'h8220000;
      8261: inst = 32'h10408000;
      8262: inst = 32'hc4043cb;
      8263: inst = 32'h8220000;
      8264: inst = 32'h10408000;
      8265: inst = 32'hc4043cc;
      8266: inst = 32'h8220000;
      8267: inst = 32'h10408000;
      8268: inst = 32'hc4043cd;
      8269: inst = 32'h8220000;
      8270: inst = 32'h10408000;
      8271: inst = 32'hc4043ce;
      8272: inst = 32'h8220000;
      8273: inst = 32'h10408000;
      8274: inst = 32'hc4043cf;
      8275: inst = 32'h8220000;
      8276: inst = 32'h10408000;
      8277: inst = 32'hc4043d0;
      8278: inst = 32'h8220000;
      8279: inst = 32'h10408000;
      8280: inst = 32'hc4043d1;
      8281: inst = 32'h8220000;
      8282: inst = 32'h10408000;
      8283: inst = 32'hc4043d2;
      8284: inst = 32'h8220000;
      8285: inst = 32'h10408000;
      8286: inst = 32'hc4043d3;
      8287: inst = 32'h8220000;
      8288: inst = 32'h10408000;
      8289: inst = 32'hc4043d4;
      8290: inst = 32'h8220000;
      8291: inst = 32'h10408000;
      8292: inst = 32'hc4043d5;
      8293: inst = 32'h8220000;
      8294: inst = 32'h10408000;
      8295: inst = 32'hc4043d6;
      8296: inst = 32'h8220000;
      8297: inst = 32'h10408000;
      8298: inst = 32'hc4043d7;
      8299: inst = 32'h8220000;
      8300: inst = 32'h10408000;
      8301: inst = 32'hc4043d8;
      8302: inst = 32'h8220000;
      8303: inst = 32'h10408000;
      8304: inst = 32'hc4043d9;
      8305: inst = 32'h8220000;
      8306: inst = 32'h10408000;
      8307: inst = 32'hc4043da;
      8308: inst = 32'h8220000;
      8309: inst = 32'h10408000;
      8310: inst = 32'hc4043db;
      8311: inst = 32'h8220000;
      8312: inst = 32'h10408000;
      8313: inst = 32'hc4043dc;
      8314: inst = 32'h8220000;
      8315: inst = 32'h10408000;
      8316: inst = 32'hc4043dd;
      8317: inst = 32'h8220000;
      8318: inst = 32'h10408000;
      8319: inst = 32'hc4043de;
      8320: inst = 32'h8220000;
      8321: inst = 32'h10408000;
      8322: inst = 32'hc4043df;
      8323: inst = 32'h8220000;
      8324: inst = 32'h10408000;
      8325: inst = 32'hc4043e0;
      8326: inst = 32'h8220000;
      8327: inst = 32'h10408000;
      8328: inst = 32'hc4043e1;
      8329: inst = 32'h8220000;
      8330: inst = 32'h10408000;
      8331: inst = 32'hc4043e2;
      8332: inst = 32'h8220000;
      8333: inst = 32'h10408000;
      8334: inst = 32'hc4043e3;
      8335: inst = 32'h8220000;
      8336: inst = 32'h10408000;
      8337: inst = 32'hc40441c;
      8338: inst = 32'h8220000;
      8339: inst = 32'h10408000;
      8340: inst = 32'hc40441d;
      8341: inst = 32'h8220000;
      8342: inst = 32'h10408000;
      8343: inst = 32'hc40441e;
      8344: inst = 32'h8220000;
      8345: inst = 32'h10408000;
      8346: inst = 32'hc40441f;
      8347: inst = 32'h8220000;
      8348: inst = 32'h10408000;
      8349: inst = 32'hc404420;
      8350: inst = 32'h8220000;
      8351: inst = 32'h10408000;
      8352: inst = 32'hc404421;
      8353: inst = 32'h8220000;
      8354: inst = 32'h10408000;
      8355: inst = 32'hc404422;
      8356: inst = 32'h8220000;
      8357: inst = 32'h10408000;
      8358: inst = 32'hc404423;
      8359: inst = 32'h8220000;
      8360: inst = 32'h10408000;
      8361: inst = 32'hc404424;
      8362: inst = 32'h8220000;
      8363: inst = 32'h10408000;
      8364: inst = 32'hc404425;
      8365: inst = 32'h8220000;
      8366: inst = 32'h10408000;
      8367: inst = 32'hc404426;
      8368: inst = 32'h8220000;
      8369: inst = 32'h10408000;
      8370: inst = 32'hc404427;
      8371: inst = 32'h8220000;
      8372: inst = 32'h10408000;
      8373: inst = 32'hc404428;
      8374: inst = 32'h8220000;
      8375: inst = 32'h10408000;
      8376: inst = 32'hc404429;
      8377: inst = 32'h8220000;
      8378: inst = 32'h10408000;
      8379: inst = 32'hc40442a;
      8380: inst = 32'h8220000;
      8381: inst = 32'h10408000;
      8382: inst = 32'hc40442b;
      8383: inst = 32'h8220000;
      8384: inst = 32'h10408000;
      8385: inst = 32'hc40442c;
      8386: inst = 32'h8220000;
      8387: inst = 32'h10408000;
      8388: inst = 32'hc40442d;
      8389: inst = 32'h8220000;
      8390: inst = 32'h10408000;
      8391: inst = 32'hc40442e;
      8392: inst = 32'h8220000;
      8393: inst = 32'h10408000;
      8394: inst = 32'hc40442f;
      8395: inst = 32'h8220000;
      8396: inst = 32'h10408000;
      8397: inst = 32'hc404430;
      8398: inst = 32'h8220000;
      8399: inst = 32'h10408000;
      8400: inst = 32'hc404431;
      8401: inst = 32'h8220000;
      8402: inst = 32'h10408000;
      8403: inst = 32'hc404432;
      8404: inst = 32'h8220000;
      8405: inst = 32'h10408000;
      8406: inst = 32'hc404433;
      8407: inst = 32'h8220000;
      8408: inst = 32'h10408000;
      8409: inst = 32'hc404434;
      8410: inst = 32'h8220000;
      8411: inst = 32'h10408000;
      8412: inst = 32'hc404435;
      8413: inst = 32'h8220000;
      8414: inst = 32'h10408000;
      8415: inst = 32'hc404436;
      8416: inst = 32'h8220000;
      8417: inst = 32'h10408000;
      8418: inst = 32'hc404437;
      8419: inst = 32'h8220000;
      8420: inst = 32'h10408000;
      8421: inst = 32'hc404438;
      8422: inst = 32'h8220000;
      8423: inst = 32'h10408000;
      8424: inst = 32'hc404439;
      8425: inst = 32'h8220000;
      8426: inst = 32'h10408000;
      8427: inst = 32'hc40443a;
      8428: inst = 32'h8220000;
      8429: inst = 32'h10408000;
      8430: inst = 32'hc40443b;
      8431: inst = 32'h8220000;
      8432: inst = 32'h10408000;
      8433: inst = 32'hc40443c;
      8434: inst = 32'h8220000;
      8435: inst = 32'h10408000;
      8436: inst = 32'hc40443d;
      8437: inst = 32'h8220000;
      8438: inst = 32'h10408000;
      8439: inst = 32'hc40443e;
      8440: inst = 32'h8220000;
      8441: inst = 32'h10408000;
      8442: inst = 32'hc40443f;
      8443: inst = 32'h8220000;
      8444: inst = 32'h10408000;
      8445: inst = 32'hc404440;
      8446: inst = 32'h8220000;
      8447: inst = 32'h10408000;
      8448: inst = 32'hc404441;
      8449: inst = 32'h8220000;
      8450: inst = 32'h10408000;
      8451: inst = 32'hc404442;
      8452: inst = 32'h8220000;
      8453: inst = 32'h10408000;
      8454: inst = 32'hc404443;
      8455: inst = 32'h8220000;
      8456: inst = 32'h10408000;
      8457: inst = 32'hc40447c;
      8458: inst = 32'h8220000;
      8459: inst = 32'h10408000;
      8460: inst = 32'hc40447d;
      8461: inst = 32'h8220000;
      8462: inst = 32'h10408000;
      8463: inst = 32'hc40447e;
      8464: inst = 32'h8220000;
      8465: inst = 32'h10408000;
      8466: inst = 32'hc40447f;
      8467: inst = 32'h8220000;
      8468: inst = 32'h10408000;
      8469: inst = 32'hc404480;
      8470: inst = 32'h8220000;
      8471: inst = 32'h10408000;
      8472: inst = 32'hc404481;
      8473: inst = 32'h8220000;
      8474: inst = 32'h10408000;
      8475: inst = 32'hc404482;
      8476: inst = 32'h8220000;
      8477: inst = 32'h10408000;
      8478: inst = 32'hc404483;
      8479: inst = 32'h8220000;
      8480: inst = 32'h10408000;
      8481: inst = 32'hc404484;
      8482: inst = 32'h8220000;
      8483: inst = 32'h10408000;
      8484: inst = 32'hc404485;
      8485: inst = 32'h8220000;
      8486: inst = 32'h10408000;
      8487: inst = 32'hc404486;
      8488: inst = 32'h8220000;
      8489: inst = 32'h10408000;
      8490: inst = 32'hc404487;
      8491: inst = 32'h8220000;
      8492: inst = 32'h10408000;
      8493: inst = 32'hc404488;
      8494: inst = 32'h8220000;
      8495: inst = 32'h10408000;
      8496: inst = 32'hc404489;
      8497: inst = 32'h8220000;
      8498: inst = 32'h10408000;
      8499: inst = 32'hc40448a;
      8500: inst = 32'h8220000;
      8501: inst = 32'h10408000;
      8502: inst = 32'hc40448b;
      8503: inst = 32'h8220000;
      8504: inst = 32'h10408000;
      8505: inst = 32'hc40448c;
      8506: inst = 32'h8220000;
      8507: inst = 32'h10408000;
      8508: inst = 32'hc40448d;
      8509: inst = 32'h8220000;
      8510: inst = 32'h10408000;
      8511: inst = 32'hc40448e;
      8512: inst = 32'h8220000;
      8513: inst = 32'h10408000;
      8514: inst = 32'hc40448f;
      8515: inst = 32'h8220000;
      8516: inst = 32'h10408000;
      8517: inst = 32'hc404490;
      8518: inst = 32'h8220000;
      8519: inst = 32'h10408000;
      8520: inst = 32'hc404491;
      8521: inst = 32'h8220000;
      8522: inst = 32'h10408000;
      8523: inst = 32'hc404492;
      8524: inst = 32'h8220000;
      8525: inst = 32'h10408000;
      8526: inst = 32'hc404493;
      8527: inst = 32'h8220000;
      8528: inst = 32'h10408000;
      8529: inst = 32'hc404494;
      8530: inst = 32'h8220000;
      8531: inst = 32'h10408000;
      8532: inst = 32'hc404495;
      8533: inst = 32'h8220000;
      8534: inst = 32'h10408000;
      8535: inst = 32'hc404496;
      8536: inst = 32'h8220000;
      8537: inst = 32'h10408000;
      8538: inst = 32'hc404497;
      8539: inst = 32'h8220000;
      8540: inst = 32'h10408000;
      8541: inst = 32'hc404498;
      8542: inst = 32'h8220000;
      8543: inst = 32'h10408000;
      8544: inst = 32'hc404499;
      8545: inst = 32'h8220000;
      8546: inst = 32'h10408000;
      8547: inst = 32'hc40449a;
      8548: inst = 32'h8220000;
      8549: inst = 32'h10408000;
      8550: inst = 32'hc40449b;
      8551: inst = 32'h8220000;
      8552: inst = 32'h10408000;
      8553: inst = 32'hc40449c;
      8554: inst = 32'h8220000;
      8555: inst = 32'h10408000;
      8556: inst = 32'hc40449d;
      8557: inst = 32'h8220000;
      8558: inst = 32'h10408000;
      8559: inst = 32'hc40449e;
      8560: inst = 32'h8220000;
      8561: inst = 32'h10408000;
      8562: inst = 32'hc40449f;
      8563: inst = 32'h8220000;
      8564: inst = 32'h10408000;
      8565: inst = 32'hc4044a0;
      8566: inst = 32'h8220000;
      8567: inst = 32'h10408000;
      8568: inst = 32'hc4044a1;
      8569: inst = 32'h8220000;
      8570: inst = 32'h10408000;
      8571: inst = 32'hc4044a2;
      8572: inst = 32'h8220000;
      8573: inst = 32'h10408000;
      8574: inst = 32'hc4044a3;
      8575: inst = 32'h8220000;
      8576: inst = 32'h10408000;
      8577: inst = 32'hc4044dc;
      8578: inst = 32'h8220000;
      8579: inst = 32'h10408000;
      8580: inst = 32'hc4044dd;
      8581: inst = 32'h8220000;
      8582: inst = 32'h10408000;
      8583: inst = 32'hc4044de;
      8584: inst = 32'h8220000;
      8585: inst = 32'h10408000;
      8586: inst = 32'hc4044df;
      8587: inst = 32'h8220000;
      8588: inst = 32'h10408000;
      8589: inst = 32'hc4044e0;
      8590: inst = 32'h8220000;
      8591: inst = 32'h10408000;
      8592: inst = 32'hc4044e1;
      8593: inst = 32'h8220000;
      8594: inst = 32'h10408000;
      8595: inst = 32'hc4044e2;
      8596: inst = 32'h8220000;
      8597: inst = 32'h10408000;
      8598: inst = 32'hc4044e3;
      8599: inst = 32'h8220000;
      8600: inst = 32'h10408000;
      8601: inst = 32'hc4044e4;
      8602: inst = 32'h8220000;
      8603: inst = 32'h10408000;
      8604: inst = 32'hc4044e5;
      8605: inst = 32'h8220000;
      8606: inst = 32'h10408000;
      8607: inst = 32'hc4044e6;
      8608: inst = 32'h8220000;
      8609: inst = 32'h10408000;
      8610: inst = 32'hc4044e7;
      8611: inst = 32'h8220000;
      8612: inst = 32'h10408000;
      8613: inst = 32'hc4044e8;
      8614: inst = 32'h8220000;
      8615: inst = 32'h10408000;
      8616: inst = 32'hc4044e9;
      8617: inst = 32'h8220000;
      8618: inst = 32'h10408000;
      8619: inst = 32'hc4044ea;
      8620: inst = 32'h8220000;
      8621: inst = 32'h10408000;
      8622: inst = 32'hc4044eb;
      8623: inst = 32'h8220000;
      8624: inst = 32'h10408000;
      8625: inst = 32'hc4044ec;
      8626: inst = 32'h8220000;
      8627: inst = 32'h10408000;
      8628: inst = 32'hc4044ed;
      8629: inst = 32'h8220000;
      8630: inst = 32'h10408000;
      8631: inst = 32'hc4044ee;
      8632: inst = 32'h8220000;
      8633: inst = 32'h10408000;
      8634: inst = 32'hc4044ef;
      8635: inst = 32'h8220000;
      8636: inst = 32'h10408000;
      8637: inst = 32'hc4044f0;
      8638: inst = 32'h8220000;
      8639: inst = 32'h10408000;
      8640: inst = 32'hc4044f1;
      8641: inst = 32'h8220000;
      8642: inst = 32'h10408000;
      8643: inst = 32'hc4044f2;
      8644: inst = 32'h8220000;
      8645: inst = 32'h10408000;
      8646: inst = 32'hc4044f3;
      8647: inst = 32'h8220000;
      8648: inst = 32'h10408000;
      8649: inst = 32'hc4044f4;
      8650: inst = 32'h8220000;
      8651: inst = 32'h10408000;
      8652: inst = 32'hc4044f5;
      8653: inst = 32'h8220000;
      8654: inst = 32'h10408000;
      8655: inst = 32'hc4044f6;
      8656: inst = 32'h8220000;
      8657: inst = 32'h10408000;
      8658: inst = 32'hc4044f7;
      8659: inst = 32'h8220000;
      8660: inst = 32'h10408000;
      8661: inst = 32'hc4044f8;
      8662: inst = 32'h8220000;
      8663: inst = 32'h10408000;
      8664: inst = 32'hc4044f9;
      8665: inst = 32'h8220000;
      8666: inst = 32'h10408000;
      8667: inst = 32'hc4044fa;
      8668: inst = 32'h8220000;
      8669: inst = 32'h10408000;
      8670: inst = 32'hc4044fb;
      8671: inst = 32'h8220000;
      8672: inst = 32'h10408000;
      8673: inst = 32'hc4044fc;
      8674: inst = 32'h8220000;
      8675: inst = 32'h10408000;
      8676: inst = 32'hc4044fd;
      8677: inst = 32'h8220000;
      8678: inst = 32'h10408000;
      8679: inst = 32'hc4044fe;
      8680: inst = 32'h8220000;
      8681: inst = 32'h10408000;
      8682: inst = 32'hc4044ff;
      8683: inst = 32'h8220000;
      8684: inst = 32'h10408000;
      8685: inst = 32'hc404500;
      8686: inst = 32'h8220000;
      8687: inst = 32'h10408000;
      8688: inst = 32'hc404501;
      8689: inst = 32'h8220000;
      8690: inst = 32'h10408000;
      8691: inst = 32'hc404502;
      8692: inst = 32'h8220000;
      8693: inst = 32'h10408000;
      8694: inst = 32'hc404503;
      8695: inst = 32'h8220000;
      8696: inst = 32'h10408000;
      8697: inst = 32'hc40453c;
      8698: inst = 32'h8220000;
      8699: inst = 32'h10408000;
      8700: inst = 32'hc40453d;
      8701: inst = 32'h8220000;
      8702: inst = 32'h10408000;
      8703: inst = 32'hc40453e;
      8704: inst = 32'h8220000;
      8705: inst = 32'h10408000;
      8706: inst = 32'hc40453f;
      8707: inst = 32'h8220000;
      8708: inst = 32'h10408000;
      8709: inst = 32'hc404540;
      8710: inst = 32'h8220000;
      8711: inst = 32'h10408000;
      8712: inst = 32'hc404541;
      8713: inst = 32'h8220000;
      8714: inst = 32'h10408000;
      8715: inst = 32'hc404542;
      8716: inst = 32'h8220000;
      8717: inst = 32'h10408000;
      8718: inst = 32'hc404543;
      8719: inst = 32'h8220000;
      8720: inst = 32'h10408000;
      8721: inst = 32'hc404544;
      8722: inst = 32'h8220000;
      8723: inst = 32'h10408000;
      8724: inst = 32'hc404545;
      8725: inst = 32'h8220000;
      8726: inst = 32'h10408000;
      8727: inst = 32'hc404546;
      8728: inst = 32'h8220000;
      8729: inst = 32'h10408000;
      8730: inst = 32'hc404547;
      8731: inst = 32'h8220000;
      8732: inst = 32'h10408000;
      8733: inst = 32'hc404548;
      8734: inst = 32'h8220000;
      8735: inst = 32'h10408000;
      8736: inst = 32'hc404549;
      8737: inst = 32'h8220000;
      8738: inst = 32'h10408000;
      8739: inst = 32'hc40454a;
      8740: inst = 32'h8220000;
      8741: inst = 32'h10408000;
      8742: inst = 32'hc40454b;
      8743: inst = 32'h8220000;
      8744: inst = 32'h10408000;
      8745: inst = 32'hc40454c;
      8746: inst = 32'h8220000;
      8747: inst = 32'h10408000;
      8748: inst = 32'hc40454d;
      8749: inst = 32'h8220000;
      8750: inst = 32'h10408000;
      8751: inst = 32'hc40454e;
      8752: inst = 32'h8220000;
      8753: inst = 32'h10408000;
      8754: inst = 32'hc40454f;
      8755: inst = 32'h8220000;
      8756: inst = 32'h10408000;
      8757: inst = 32'hc404550;
      8758: inst = 32'h8220000;
      8759: inst = 32'h10408000;
      8760: inst = 32'hc404551;
      8761: inst = 32'h8220000;
      8762: inst = 32'h10408000;
      8763: inst = 32'hc404552;
      8764: inst = 32'h8220000;
      8765: inst = 32'h10408000;
      8766: inst = 32'hc404553;
      8767: inst = 32'h8220000;
      8768: inst = 32'h10408000;
      8769: inst = 32'hc404554;
      8770: inst = 32'h8220000;
      8771: inst = 32'h10408000;
      8772: inst = 32'hc404555;
      8773: inst = 32'h8220000;
      8774: inst = 32'h10408000;
      8775: inst = 32'hc404556;
      8776: inst = 32'h8220000;
      8777: inst = 32'h10408000;
      8778: inst = 32'hc404557;
      8779: inst = 32'h8220000;
      8780: inst = 32'h10408000;
      8781: inst = 32'hc404558;
      8782: inst = 32'h8220000;
      8783: inst = 32'h10408000;
      8784: inst = 32'hc404559;
      8785: inst = 32'h8220000;
      8786: inst = 32'h10408000;
      8787: inst = 32'hc40455a;
      8788: inst = 32'h8220000;
      8789: inst = 32'h10408000;
      8790: inst = 32'hc40455b;
      8791: inst = 32'h8220000;
      8792: inst = 32'h10408000;
      8793: inst = 32'hc40455c;
      8794: inst = 32'h8220000;
      8795: inst = 32'h10408000;
      8796: inst = 32'hc40455d;
      8797: inst = 32'h8220000;
      8798: inst = 32'h10408000;
      8799: inst = 32'hc40455e;
      8800: inst = 32'h8220000;
      8801: inst = 32'h10408000;
      8802: inst = 32'hc40455f;
      8803: inst = 32'h8220000;
      8804: inst = 32'h10408000;
      8805: inst = 32'hc404560;
      8806: inst = 32'h8220000;
      8807: inst = 32'h10408000;
      8808: inst = 32'hc404561;
      8809: inst = 32'h8220000;
      8810: inst = 32'h10408000;
      8811: inst = 32'hc404562;
      8812: inst = 32'h8220000;
      8813: inst = 32'h10408000;
      8814: inst = 32'hc404563;
      8815: inst = 32'h8220000;
      8816: inst = 32'h10408000;
      8817: inst = 32'hc40459c;
      8818: inst = 32'h8220000;
      8819: inst = 32'h10408000;
      8820: inst = 32'hc40459d;
      8821: inst = 32'h8220000;
      8822: inst = 32'h10408000;
      8823: inst = 32'hc40459e;
      8824: inst = 32'h8220000;
      8825: inst = 32'h10408000;
      8826: inst = 32'hc40459f;
      8827: inst = 32'h8220000;
      8828: inst = 32'h10408000;
      8829: inst = 32'hc4045a0;
      8830: inst = 32'h8220000;
      8831: inst = 32'h10408000;
      8832: inst = 32'hc4045a1;
      8833: inst = 32'h8220000;
      8834: inst = 32'h10408000;
      8835: inst = 32'hc4045a2;
      8836: inst = 32'h8220000;
      8837: inst = 32'h10408000;
      8838: inst = 32'hc4045a3;
      8839: inst = 32'h8220000;
      8840: inst = 32'h10408000;
      8841: inst = 32'hc4045a4;
      8842: inst = 32'h8220000;
      8843: inst = 32'h10408000;
      8844: inst = 32'hc4045a5;
      8845: inst = 32'h8220000;
      8846: inst = 32'h10408000;
      8847: inst = 32'hc4045a6;
      8848: inst = 32'h8220000;
      8849: inst = 32'h10408000;
      8850: inst = 32'hc4045a7;
      8851: inst = 32'h8220000;
      8852: inst = 32'h10408000;
      8853: inst = 32'hc4045a8;
      8854: inst = 32'h8220000;
      8855: inst = 32'h10408000;
      8856: inst = 32'hc4045a9;
      8857: inst = 32'h8220000;
      8858: inst = 32'h10408000;
      8859: inst = 32'hc4045aa;
      8860: inst = 32'h8220000;
      8861: inst = 32'h10408000;
      8862: inst = 32'hc4045ab;
      8863: inst = 32'h8220000;
      8864: inst = 32'h10408000;
      8865: inst = 32'hc4045ac;
      8866: inst = 32'h8220000;
      8867: inst = 32'h10408000;
      8868: inst = 32'hc4045ad;
      8869: inst = 32'h8220000;
      8870: inst = 32'h10408000;
      8871: inst = 32'hc4045ae;
      8872: inst = 32'h8220000;
      8873: inst = 32'h10408000;
      8874: inst = 32'hc4045af;
      8875: inst = 32'h8220000;
      8876: inst = 32'h10408000;
      8877: inst = 32'hc4045b0;
      8878: inst = 32'h8220000;
      8879: inst = 32'h10408000;
      8880: inst = 32'hc4045b1;
      8881: inst = 32'h8220000;
      8882: inst = 32'h10408000;
      8883: inst = 32'hc4045b2;
      8884: inst = 32'h8220000;
      8885: inst = 32'h10408000;
      8886: inst = 32'hc4045b3;
      8887: inst = 32'h8220000;
      8888: inst = 32'h10408000;
      8889: inst = 32'hc4045b4;
      8890: inst = 32'h8220000;
      8891: inst = 32'h10408000;
      8892: inst = 32'hc4045b5;
      8893: inst = 32'h8220000;
      8894: inst = 32'h10408000;
      8895: inst = 32'hc4045b6;
      8896: inst = 32'h8220000;
      8897: inst = 32'h10408000;
      8898: inst = 32'hc4045b7;
      8899: inst = 32'h8220000;
      8900: inst = 32'h10408000;
      8901: inst = 32'hc4045b8;
      8902: inst = 32'h8220000;
      8903: inst = 32'h10408000;
      8904: inst = 32'hc4045b9;
      8905: inst = 32'h8220000;
      8906: inst = 32'h10408000;
      8907: inst = 32'hc4045ba;
      8908: inst = 32'h8220000;
      8909: inst = 32'h10408000;
      8910: inst = 32'hc4045bb;
      8911: inst = 32'h8220000;
      8912: inst = 32'h10408000;
      8913: inst = 32'hc4045bc;
      8914: inst = 32'h8220000;
      8915: inst = 32'h10408000;
      8916: inst = 32'hc4045bd;
      8917: inst = 32'h8220000;
      8918: inst = 32'h10408000;
      8919: inst = 32'hc4045be;
      8920: inst = 32'h8220000;
      8921: inst = 32'h10408000;
      8922: inst = 32'hc4045bf;
      8923: inst = 32'h8220000;
      8924: inst = 32'h10408000;
      8925: inst = 32'hc4045c0;
      8926: inst = 32'h8220000;
      8927: inst = 32'h10408000;
      8928: inst = 32'hc4045c1;
      8929: inst = 32'h8220000;
      8930: inst = 32'h10408000;
      8931: inst = 32'hc4045c2;
      8932: inst = 32'h8220000;
      8933: inst = 32'h10408000;
      8934: inst = 32'hc4045c3;
      8935: inst = 32'h8220000;
      8936: inst = 32'h10408000;
      8937: inst = 32'hc4045fc;
      8938: inst = 32'h8220000;
      8939: inst = 32'h10408000;
      8940: inst = 32'hc4045fd;
      8941: inst = 32'h8220000;
      8942: inst = 32'h10408000;
      8943: inst = 32'hc4045fe;
      8944: inst = 32'h8220000;
      8945: inst = 32'h10408000;
      8946: inst = 32'hc4045ff;
      8947: inst = 32'h8220000;
      8948: inst = 32'h10408000;
      8949: inst = 32'hc404600;
      8950: inst = 32'h8220000;
      8951: inst = 32'h10408000;
      8952: inst = 32'hc404601;
      8953: inst = 32'h8220000;
      8954: inst = 32'h10408000;
      8955: inst = 32'hc404602;
      8956: inst = 32'h8220000;
      8957: inst = 32'h10408000;
      8958: inst = 32'hc404603;
      8959: inst = 32'h8220000;
      8960: inst = 32'h10408000;
      8961: inst = 32'hc404604;
      8962: inst = 32'h8220000;
      8963: inst = 32'h10408000;
      8964: inst = 32'hc404605;
      8965: inst = 32'h8220000;
      8966: inst = 32'h10408000;
      8967: inst = 32'hc404606;
      8968: inst = 32'h8220000;
      8969: inst = 32'h10408000;
      8970: inst = 32'hc404607;
      8971: inst = 32'h8220000;
      8972: inst = 32'h10408000;
      8973: inst = 32'hc404608;
      8974: inst = 32'h8220000;
      8975: inst = 32'h10408000;
      8976: inst = 32'hc404609;
      8977: inst = 32'h8220000;
      8978: inst = 32'h10408000;
      8979: inst = 32'hc40460a;
      8980: inst = 32'h8220000;
      8981: inst = 32'h10408000;
      8982: inst = 32'hc40460b;
      8983: inst = 32'h8220000;
      8984: inst = 32'h10408000;
      8985: inst = 32'hc40460c;
      8986: inst = 32'h8220000;
      8987: inst = 32'h10408000;
      8988: inst = 32'hc40460d;
      8989: inst = 32'h8220000;
      8990: inst = 32'h10408000;
      8991: inst = 32'hc40460e;
      8992: inst = 32'h8220000;
      8993: inst = 32'h10408000;
      8994: inst = 32'hc40460f;
      8995: inst = 32'h8220000;
      8996: inst = 32'h10408000;
      8997: inst = 32'hc404610;
      8998: inst = 32'h8220000;
      8999: inst = 32'h10408000;
      9000: inst = 32'hc404611;
      9001: inst = 32'h8220000;
      9002: inst = 32'h10408000;
      9003: inst = 32'hc404612;
      9004: inst = 32'h8220000;
      9005: inst = 32'h10408000;
      9006: inst = 32'hc404613;
      9007: inst = 32'h8220000;
      9008: inst = 32'h10408000;
      9009: inst = 32'hc404614;
      9010: inst = 32'h8220000;
      9011: inst = 32'h10408000;
      9012: inst = 32'hc404615;
      9013: inst = 32'h8220000;
      9014: inst = 32'h10408000;
      9015: inst = 32'hc404616;
      9016: inst = 32'h8220000;
      9017: inst = 32'h10408000;
      9018: inst = 32'hc404617;
      9019: inst = 32'h8220000;
      9020: inst = 32'h10408000;
      9021: inst = 32'hc404618;
      9022: inst = 32'h8220000;
      9023: inst = 32'h10408000;
      9024: inst = 32'hc404619;
      9025: inst = 32'h8220000;
      9026: inst = 32'h10408000;
      9027: inst = 32'hc40461a;
      9028: inst = 32'h8220000;
      9029: inst = 32'h10408000;
      9030: inst = 32'hc40461b;
      9031: inst = 32'h8220000;
      9032: inst = 32'h10408000;
      9033: inst = 32'hc40461c;
      9034: inst = 32'h8220000;
      9035: inst = 32'h10408000;
      9036: inst = 32'hc40461d;
      9037: inst = 32'h8220000;
      9038: inst = 32'h10408000;
      9039: inst = 32'hc40461e;
      9040: inst = 32'h8220000;
      9041: inst = 32'h10408000;
      9042: inst = 32'hc40461f;
      9043: inst = 32'h8220000;
      9044: inst = 32'h10408000;
      9045: inst = 32'hc404620;
      9046: inst = 32'h8220000;
      9047: inst = 32'h10408000;
      9048: inst = 32'hc404621;
      9049: inst = 32'h8220000;
      9050: inst = 32'h10408000;
      9051: inst = 32'hc404622;
      9052: inst = 32'h8220000;
      9053: inst = 32'h10408000;
      9054: inst = 32'hc404623;
      9055: inst = 32'h8220000;
      9056: inst = 32'h10408000;
      9057: inst = 32'hc40465c;
      9058: inst = 32'h8220000;
      9059: inst = 32'h10408000;
      9060: inst = 32'hc40465d;
      9061: inst = 32'h8220000;
      9062: inst = 32'h10408000;
      9063: inst = 32'hc40465e;
      9064: inst = 32'h8220000;
      9065: inst = 32'h10408000;
      9066: inst = 32'hc40465f;
      9067: inst = 32'h8220000;
      9068: inst = 32'h10408000;
      9069: inst = 32'hc404660;
      9070: inst = 32'h8220000;
      9071: inst = 32'h10408000;
      9072: inst = 32'hc404661;
      9073: inst = 32'h8220000;
      9074: inst = 32'h10408000;
      9075: inst = 32'hc404662;
      9076: inst = 32'h8220000;
      9077: inst = 32'h10408000;
      9078: inst = 32'hc404663;
      9079: inst = 32'h8220000;
      9080: inst = 32'h10408000;
      9081: inst = 32'hc404664;
      9082: inst = 32'h8220000;
      9083: inst = 32'h10408000;
      9084: inst = 32'hc404665;
      9085: inst = 32'h8220000;
      9086: inst = 32'h10408000;
      9087: inst = 32'hc404666;
      9088: inst = 32'h8220000;
      9089: inst = 32'h10408000;
      9090: inst = 32'hc404667;
      9091: inst = 32'h8220000;
      9092: inst = 32'h10408000;
      9093: inst = 32'hc404668;
      9094: inst = 32'h8220000;
      9095: inst = 32'h10408000;
      9096: inst = 32'hc404669;
      9097: inst = 32'h8220000;
      9098: inst = 32'h10408000;
      9099: inst = 32'hc40466a;
      9100: inst = 32'h8220000;
      9101: inst = 32'h10408000;
      9102: inst = 32'hc40466b;
      9103: inst = 32'h8220000;
      9104: inst = 32'h10408000;
      9105: inst = 32'hc40466c;
      9106: inst = 32'h8220000;
      9107: inst = 32'h10408000;
      9108: inst = 32'hc40466d;
      9109: inst = 32'h8220000;
      9110: inst = 32'h10408000;
      9111: inst = 32'hc40466e;
      9112: inst = 32'h8220000;
      9113: inst = 32'h10408000;
      9114: inst = 32'hc40466f;
      9115: inst = 32'h8220000;
      9116: inst = 32'h10408000;
      9117: inst = 32'hc404670;
      9118: inst = 32'h8220000;
      9119: inst = 32'h10408000;
      9120: inst = 32'hc404671;
      9121: inst = 32'h8220000;
      9122: inst = 32'h10408000;
      9123: inst = 32'hc404672;
      9124: inst = 32'h8220000;
      9125: inst = 32'h10408000;
      9126: inst = 32'hc404673;
      9127: inst = 32'h8220000;
      9128: inst = 32'h10408000;
      9129: inst = 32'hc404674;
      9130: inst = 32'h8220000;
      9131: inst = 32'h10408000;
      9132: inst = 32'hc404675;
      9133: inst = 32'h8220000;
      9134: inst = 32'h10408000;
      9135: inst = 32'hc404676;
      9136: inst = 32'h8220000;
      9137: inst = 32'h10408000;
      9138: inst = 32'hc404677;
      9139: inst = 32'h8220000;
      9140: inst = 32'h10408000;
      9141: inst = 32'hc404678;
      9142: inst = 32'h8220000;
      9143: inst = 32'h10408000;
      9144: inst = 32'hc404679;
      9145: inst = 32'h8220000;
      9146: inst = 32'h10408000;
      9147: inst = 32'hc40467a;
      9148: inst = 32'h8220000;
      9149: inst = 32'h10408000;
      9150: inst = 32'hc40467b;
      9151: inst = 32'h8220000;
      9152: inst = 32'h10408000;
      9153: inst = 32'hc40467c;
      9154: inst = 32'h8220000;
      9155: inst = 32'h10408000;
      9156: inst = 32'hc40467d;
      9157: inst = 32'h8220000;
      9158: inst = 32'h10408000;
      9159: inst = 32'hc40467e;
      9160: inst = 32'h8220000;
      9161: inst = 32'h10408000;
      9162: inst = 32'hc40467f;
      9163: inst = 32'h8220000;
      9164: inst = 32'h10408000;
      9165: inst = 32'hc404680;
      9166: inst = 32'h8220000;
      9167: inst = 32'h10408000;
      9168: inst = 32'hc404681;
      9169: inst = 32'h8220000;
      9170: inst = 32'h10408000;
      9171: inst = 32'hc404682;
      9172: inst = 32'h8220000;
      9173: inst = 32'h10408000;
      9174: inst = 32'hc404683;
      9175: inst = 32'h8220000;
      9176: inst = 32'h10408000;
      9177: inst = 32'hc4046bc;
      9178: inst = 32'h8220000;
      9179: inst = 32'h10408000;
      9180: inst = 32'hc4046bd;
      9181: inst = 32'h8220000;
      9182: inst = 32'h10408000;
      9183: inst = 32'hc4046be;
      9184: inst = 32'h8220000;
      9185: inst = 32'h10408000;
      9186: inst = 32'hc4046bf;
      9187: inst = 32'h8220000;
      9188: inst = 32'h10408000;
      9189: inst = 32'hc4046c0;
      9190: inst = 32'h8220000;
      9191: inst = 32'h10408000;
      9192: inst = 32'hc4046c1;
      9193: inst = 32'h8220000;
      9194: inst = 32'h10408000;
      9195: inst = 32'hc4046c2;
      9196: inst = 32'h8220000;
      9197: inst = 32'h10408000;
      9198: inst = 32'hc4046c3;
      9199: inst = 32'h8220000;
      9200: inst = 32'h10408000;
      9201: inst = 32'hc4046c4;
      9202: inst = 32'h8220000;
      9203: inst = 32'h10408000;
      9204: inst = 32'hc4046c5;
      9205: inst = 32'h8220000;
      9206: inst = 32'h10408000;
      9207: inst = 32'hc4046c6;
      9208: inst = 32'h8220000;
      9209: inst = 32'h10408000;
      9210: inst = 32'hc4046c7;
      9211: inst = 32'h8220000;
      9212: inst = 32'h10408000;
      9213: inst = 32'hc4046c8;
      9214: inst = 32'h8220000;
      9215: inst = 32'h10408000;
      9216: inst = 32'hc4046c9;
      9217: inst = 32'h8220000;
      9218: inst = 32'h10408000;
      9219: inst = 32'hc4046ca;
      9220: inst = 32'h8220000;
      9221: inst = 32'h10408000;
      9222: inst = 32'hc4046cb;
      9223: inst = 32'h8220000;
      9224: inst = 32'h10408000;
      9225: inst = 32'hc4046cc;
      9226: inst = 32'h8220000;
      9227: inst = 32'h10408000;
      9228: inst = 32'hc4046cd;
      9229: inst = 32'h8220000;
      9230: inst = 32'h10408000;
      9231: inst = 32'hc4046ce;
      9232: inst = 32'h8220000;
      9233: inst = 32'h10408000;
      9234: inst = 32'hc4046cf;
      9235: inst = 32'h8220000;
      9236: inst = 32'h10408000;
      9237: inst = 32'hc4046d0;
      9238: inst = 32'h8220000;
      9239: inst = 32'h10408000;
      9240: inst = 32'hc4046d1;
      9241: inst = 32'h8220000;
      9242: inst = 32'h10408000;
      9243: inst = 32'hc4046d2;
      9244: inst = 32'h8220000;
      9245: inst = 32'h10408000;
      9246: inst = 32'hc4046d3;
      9247: inst = 32'h8220000;
      9248: inst = 32'h10408000;
      9249: inst = 32'hc4046d4;
      9250: inst = 32'h8220000;
      9251: inst = 32'h10408000;
      9252: inst = 32'hc4046d5;
      9253: inst = 32'h8220000;
      9254: inst = 32'h10408000;
      9255: inst = 32'hc4046d6;
      9256: inst = 32'h8220000;
      9257: inst = 32'h10408000;
      9258: inst = 32'hc4046d7;
      9259: inst = 32'h8220000;
      9260: inst = 32'h10408000;
      9261: inst = 32'hc4046d8;
      9262: inst = 32'h8220000;
      9263: inst = 32'h10408000;
      9264: inst = 32'hc4046d9;
      9265: inst = 32'h8220000;
      9266: inst = 32'h10408000;
      9267: inst = 32'hc4046da;
      9268: inst = 32'h8220000;
      9269: inst = 32'h10408000;
      9270: inst = 32'hc4046db;
      9271: inst = 32'h8220000;
      9272: inst = 32'h10408000;
      9273: inst = 32'hc4046dc;
      9274: inst = 32'h8220000;
      9275: inst = 32'h10408000;
      9276: inst = 32'hc4046dd;
      9277: inst = 32'h8220000;
      9278: inst = 32'h10408000;
      9279: inst = 32'hc4046de;
      9280: inst = 32'h8220000;
      9281: inst = 32'h10408000;
      9282: inst = 32'hc4046df;
      9283: inst = 32'h8220000;
      9284: inst = 32'h10408000;
      9285: inst = 32'hc4046e0;
      9286: inst = 32'h8220000;
      9287: inst = 32'h10408000;
      9288: inst = 32'hc4046e1;
      9289: inst = 32'h8220000;
      9290: inst = 32'h10408000;
      9291: inst = 32'hc4046e2;
      9292: inst = 32'h8220000;
      9293: inst = 32'h10408000;
      9294: inst = 32'hc4046e3;
      9295: inst = 32'h8220000;
      9296: inst = 32'h10408000;
      9297: inst = 32'hc40471c;
      9298: inst = 32'h8220000;
      9299: inst = 32'h10408000;
      9300: inst = 32'hc40471d;
      9301: inst = 32'h8220000;
      9302: inst = 32'h10408000;
      9303: inst = 32'hc40471e;
      9304: inst = 32'h8220000;
      9305: inst = 32'h10408000;
      9306: inst = 32'hc40471f;
      9307: inst = 32'h8220000;
      9308: inst = 32'h10408000;
      9309: inst = 32'hc404720;
      9310: inst = 32'h8220000;
      9311: inst = 32'h10408000;
      9312: inst = 32'hc404721;
      9313: inst = 32'h8220000;
      9314: inst = 32'h10408000;
      9315: inst = 32'hc404722;
      9316: inst = 32'h8220000;
      9317: inst = 32'h10408000;
      9318: inst = 32'hc404723;
      9319: inst = 32'h8220000;
      9320: inst = 32'h10408000;
      9321: inst = 32'hc404724;
      9322: inst = 32'h8220000;
      9323: inst = 32'h10408000;
      9324: inst = 32'hc404725;
      9325: inst = 32'h8220000;
      9326: inst = 32'h10408000;
      9327: inst = 32'hc404726;
      9328: inst = 32'h8220000;
      9329: inst = 32'h10408000;
      9330: inst = 32'hc404727;
      9331: inst = 32'h8220000;
      9332: inst = 32'h10408000;
      9333: inst = 32'hc404728;
      9334: inst = 32'h8220000;
      9335: inst = 32'h10408000;
      9336: inst = 32'hc404729;
      9337: inst = 32'h8220000;
      9338: inst = 32'h10408000;
      9339: inst = 32'hc40472a;
      9340: inst = 32'h8220000;
      9341: inst = 32'h10408000;
      9342: inst = 32'hc40472b;
      9343: inst = 32'h8220000;
      9344: inst = 32'h10408000;
      9345: inst = 32'hc40472c;
      9346: inst = 32'h8220000;
      9347: inst = 32'h10408000;
      9348: inst = 32'hc40472d;
      9349: inst = 32'h8220000;
      9350: inst = 32'h10408000;
      9351: inst = 32'hc40472e;
      9352: inst = 32'h8220000;
      9353: inst = 32'h10408000;
      9354: inst = 32'hc40472f;
      9355: inst = 32'h8220000;
      9356: inst = 32'h10408000;
      9357: inst = 32'hc404730;
      9358: inst = 32'h8220000;
      9359: inst = 32'h10408000;
      9360: inst = 32'hc404731;
      9361: inst = 32'h8220000;
      9362: inst = 32'h10408000;
      9363: inst = 32'hc404732;
      9364: inst = 32'h8220000;
      9365: inst = 32'h10408000;
      9366: inst = 32'hc404733;
      9367: inst = 32'h8220000;
      9368: inst = 32'h10408000;
      9369: inst = 32'hc404734;
      9370: inst = 32'h8220000;
      9371: inst = 32'h10408000;
      9372: inst = 32'hc404735;
      9373: inst = 32'h8220000;
      9374: inst = 32'h10408000;
      9375: inst = 32'hc404736;
      9376: inst = 32'h8220000;
      9377: inst = 32'h10408000;
      9378: inst = 32'hc404737;
      9379: inst = 32'h8220000;
      9380: inst = 32'h10408000;
      9381: inst = 32'hc404738;
      9382: inst = 32'h8220000;
      9383: inst = 32'h10408000;
      9384: inst = 32'hc404739;
      9385: inst = 32'h8220000;
      9386: inst = 32'h10408000;
      9387: inst = 32'hc40473a;
      9388: inst = 32'h8220000;
      9389: inst = 32'h10408000;
      9390: inst = 32'hc40473b;
      9391: inst = 32'h8220000;
      9392: inst = 32'h10408000;
      9393: inst = 32'hc40473c;
      9394: inst = 32'h8220000;
      9395: inst = 32'h10408000;
      9396: inst = 32'hc40473d;
      9397: inst = 32'h8220000;
      9398: inst = 32'h10408000;
      9399: inst = 32'hc40473e;
      9400: inst = 32'h8220000;
      9401: inst = 32'h10408000;
      9402: inst = 32'hc40473f;
      9403: inst = 32'h8220000;
      9404: inst = 32'h10408000;
      9405: inst = 32'hc404740;
      9406: inst = 32'h8220000;
      9407: inst = 32'h10408000;
      9408: inst = 32'hc404741;
      9409: inst = 32'h8220000;
      9410: inst = 32'h10408000;
      9411: inst = 32'hc404742;
      9412: inst = 32'h8220000;
      9413: inst = 32'h10408000;
      9414: inst = 32'hc404743;
      9415: inst = 32'h8220000;
      9416: inst = 32'h10408000;
      9417: inst = 32'hc40477c;
      9418: inst = 32'h8220000;
      9419: inst = 32'h10408000;
      9420: inst = 32'hc40477d;
      9421: inst = 32'h8220000;
      9422: inst = 32'h10408000;
      9423: inst = 32'hc40477e;
      9424: inst = 32'h8220000;
      9425: inst = 32'h10408000;
      9426: inst = 32'hc40477f;
      9427: inst = 32'h8220000;
      9428: inst = 32'h10408000;
      9429: inst = 32'hc404780;
      9430: inst = 32'h8220000;
      9431: inst = 32'h10408000;
      9432: inst = 32'hc404781;
      9433: inst = 32'h8220000;
      9434: inst = 32'h10408000;
      9435: inst = 32'hc404782;
      9436: inst = 32'h8220000;
      9437: inst = 32'h10408000;
      9438: inst = 32'hc404783;
      9439: inst = 32'h8220000;
      9440: inst = 32'h10408000;
      9441: inst = 32'hc404784;
      9442: inst = 32'h8220000;
      9443: inst = 32'h10408000;
      9444: inst = 32'hc404785;
      9445: inst = 32'h8220000;
      9446: inst = 32'h10408000;
      9447: inst = 32'hc404786;
      9448: inst = 32'h8220000;
      9449: inst = 32'h10408000;
      9450: inst = 32'hc404787;
      9451: inst = 32'h8220000;
      9452: inst = 32'h10408000;
      9453: inst = 32'hc404788;
      9454: inst = 32'h8220000;
      9455: inst = 32'h10408000;
      9456: inst = 32'hc404789;
      9457: inst = 32'h8220000;
      9458: inst = 32'h10408000;
      9459: inst = 32'hc40478a;
      9460: inst = 32'h8220000;
      9461: inst = 32'h10408000;
      9462: inst = 32'hc40478b;
      9463: inst = 32'h8220000;
      9464: inst = 32'h10408000;
      9465: inst = 32'hc40478c;
      9466: inst = 32'h8220000;
      9467: inst = 32'h10408000;
      9468: inst = 32'hc40478d;
      9469: inst = 32'h8220000;
      9470: inst = 32'h10408000;
      9471: inst = 32'hc40478e;
      9472: inst = 32'h8220000;
      9473: inst = 32'h10408000;
      9474: inst = 32'hc40478f;
      9475: inst = 32'h8220000;
      9476: inst = 32'h10408000;
      9477: inst = 32'hc404790;
      9478: inst = 32'h8220000;
      9479: inst = 32'h10408000;
      9480: inst = 32'hc404791;
      9481: inst = 32'h8220000;
      9482: inst = 32'h10408000;
      9483: inst = 32'hc404792;
      9484: inst = 32'h8220000;
      9485: inst = 32'h10408000;
      9486: inst = 32'hc404793;
      9487: inst = 32'h8220000;
      9488: inst = 32'h10408000;
      9489: inst = 32'hc404794;
      9490: inst = 32'h8220000;
      9491: inst = 32'h10408000;
      9492: inst = 32'hc404795;
      9493: inst = 32'h8220000;
      9494: inst = 32'h10408000;
      9495: inst = 32'hc404796;
      9496: inst = 32'h8220000;
      9497: inst = 32'h10408000;
      9498: inst = 32'hc404797;
      9499: inst = 32'h8220000;
      9500: inst = 32'h10408000;
      9501: inst = 32'hc404798;
      9502: inst = 32'h8220000;
      9503: inst = 32'h10408000;
      9504: inst = 32'hc404799;
      9505: inst = 32'h8220000;
      9506: inst = 32'h10408000;
      9507: inst = 32'hc40479a;
      9508: inst = 32'h8220000;
      9509: inst = 32'h10408000;
      9510: inst = 32'hc40479b;
      9511: inst = 32'h8220000;
      9512: inst = 32'h10408000;
      9513: inst = 32'hc40479c;
      9514: inst = 32'h8220000;
      9515: inst = 32'h10408000;
      9516: inst = 32'hc40479d;
      9517: inst = 32'h8220000;
      9518: inst = 32'h10408000;
      9519: inst = 32'hc40479e;
      9520: inst = 32'h8220000;
      9521: inst = 32'h10408000;
      9522: inst = 32'hc40479f;
      9523: inst = 32'h8220000;
      9524: inst = 32'h10408000;
      9525: inst = 32'hc4047a0;
      9526: inst = 32'h8220000;
      9527: inst = 32'h10408000;
      9528: inst = 32'hc4047a1;
      9529: inst = 32'h8220000;
      9530: inst = 32'h10408000;
      9531: inst = 32'hc4047a2;
      9532: inst = 32'h8220000;
      9533: inst = 32'h10408000;
      9534: inst = 32'hc4047a3;
      9535: inst = 32'h8220000;
      9536: inst = 32'h10408000;
      9537: inst = 32'hc4047dc;
      9538: inst = 32'h8220000;
      9539: inst = 32'h10408000;
      9540: inst = 32'hc4047dd;
      9541: inst = 32'h8220000;
      9542: inst = 32'h10408000;
      9543: inst = 32'hc4047de;
      9544: inst = 32'h8220000;
      9545: inst = 32'h10408000;
      9546: inst = 32'hc4047df;
      9547: inst = 32'h8220000;
      9548: inst = 32'h10408000;
      9549: inst = 32'hc4047e0;
      9550: inst = 32'h8220000;
      9551: inst = 32'h10408000;
      9552: inst = 32'hc4047e1;
      9553: inst = 32'h8220000;
      9554: inst = 32'h10408000;
      9555: inst = 32'hc4047e2;
      9556: inst = 32'h8220000;
      9557: inst = 32'h10408000;
      9558: inst = 32'hc4047e3;
      9559: inst = 32'h8220000;
      9560: inst = 32'h10408000;
      9561: inst = 32'hc4047e4;
      9562: inst = 32'h8220000;
      9563: inst = 32'h10408000;
      9564: inst = 32'hc4047e5;
      9565: inst = 32'h8220000;
      9566: inst = 32'h10408000;
      9567: inst = 32'hc4047e6;
      9568: inst = 32'h8220000;
      9569: inst = 32'h10408000;
      9570: inst = 32'hc4047e7;
      9571: inst = 32'h8220000;
      9572: inst = 32'h10408000;
      9573: inst = 32'hc4047e8;
      9574: inst = 32'h8220000;
      9575: inst = 32'h10408000;
      9576: inst = 32'hc4047e9;
      9577: inst = 32'h8220000;
      9578: inst = 32'h10408000;
      9579: inst = 32'hc4047ea;
      9580: inst = 32'h8220000;
      9581: inst = 32'h10408000;
      9582: inst = 32'hc4047eb;
      9583: inst = 32'h8220000;
      9584: inst = 32'h10408000;
      9585: inst = 32'hc4047ec;
      9586: inst = 32'h8220000;
      9587: inst = 32'h10408000;
      9588: inst = 32'hc4047ed;
      9589: inst = 32'h8220000;
      9590: inst = 32'h10408000;
      9591: inst = 32'hc4047ee;
      9592: inst = 32'h8220000;
      9593: inst = 32'h10408000;
      9594: inst = 32'hc4047ef;
      9595: inst = 32'h8220000;
      9596: inst = 32'h10408000;
      9597: inst = 32'hc4047f0;
      9598: inst = 32'h8220000;
      9599: inst = 32'h10408000;
      9600: inst = 32'hc4047f1;
      9601: inst = 32'h8220000;
      9602: inst = 32'h10408000;
      9603: inst = 32'hc4047f2;
      9604: inst = 32'h8220000;
      9605: inst = 32'h10408000;
      9606: inst = 32'hc4047f3;
      9607: inst = 32'h8220000;
      9608: inst = 32'h10408000;
      9609: inst = 32'hc4047f4;
      9610: inst = 32'h8220000;
      9611: inst = 32'h10408000;
      9612: inst = 32'hc4047f5;
      9613: inst = 32'h8220000;
      9614: inst = 32'h10408000;
      9615: inst = 32'hc4047f6;
      9616: inst = 32'h8220000;
      9617: inst = 32'h10408000;
      9618: inst = 32'hc4047f7;
      9619: inst = 32'h8220000;
      9620: inst = 32'h10408000;
      9621: inst = 32'hc4047f8;
      9622: inst = 32'h8220000;
      9623: inst = 32'h10408000;
      9624: inst = 32'hc4047f9;
      9625: inst = 32'h8220000;
      9626: inst = 32'h10408000;
      9627: inst = 32'hc4047fa;
      9628: inst = 32'h8220000;
      9629: inst = 32'h10408000;
      9630: inst = 32'hc4047fb;
      9631: inst = 32'h8220000;
      9632: inst = 32'h10408000;
      9633: inst = 32'hc4047fc;
      9634: inst = 32'h8220000;
      9635: inst = 32'h10408000;
      9636: inst = 32'hc4047fd;
      9637: inst = 32'h8220000;
      9638: inst = 32'h10408000;
      9639: inst = 32'hc4047fe;
      9640: inst = 32'h8220000;
      9641: inst = 32'h10408000;
      9642: inst = 32'hc4047ff;
      9643: inst = 32'h8220000;
      9644: inst = 32'h10408000;
      9645: inst = 32'hc404800;
      9646: inst = 32'h8220000;
      9647: inst = 32'h10408000;
      9648: inst = 32'hc404801;
      9649: inst = 32'h8220000;
      9650: inst = 32'h10408000;
      9651: inst = 32'hc404802;
      9652: inst = 32'h8220000;
      9653: inst = 32'h10408000;
      9654: inst = 32'hc404803;
      9655: inst = 32'h8220000;
      9656: inst = 32'h10408000;
      9657: inst = 32'hc40483c;
      9658: inst = 32'h8220000;
      9659: inst = 32'h10408000;
      9660: inst = 32'hc40483d;
      9661: inst = 32'h8220000;
      9662: inst = 32'h10408000;
      9663: inst = 32'hc40483e;
      9664: inst = 32'h8220000;
      9665: inst = 32'h10408000;
      9666: inst = 32'hc40483f;
      9667: inst = 32'h8220000;
      9668: inst = 32'h10408000;
      9669: inst = 32'hc404840;
      9670: inst = 32'h8220000;
      9671: inst = 32'h10408000;
      9672: inst = 32'hc404841;
      9673: inst = 32'h8220000;
      9674: inst = 32'h10408000;
      9675: inst = 32'hc404842;
      9676: inst = 32'h8220000;
      9677: inst = 32'h10408000;
      9678: inst = 32'hc404843;
      9679: inst = 32'h8220000;
      9680: inst = 32'h10408000;
      9681: inst = 32'hc404844;
      9682: inst = 32'h8220000;
      9683: inst = 32'h10408000;
      9684: inst = 32'hc404845;
      9685: inst = 32'h8220000;
      9686: inst = 32'h10408000;
      9687: inst = 32'hc404846;
      9688: inst = 32'h8220000;
      9689: inst = 32'h10408000;
      9690: inst = 32'hc404847;
      9691: inst = 32'h8220000;
      9692: inst = 32'h10408000;
      9693: inst = 32'hc404848;
      9694: inst = 32'h8220000;
      9695: inst = 32'h10408000;
      9696: inst = 32'hc404849;
      9697: inst = 32'h8220000;
      9698: inst = 32'h10408000;
      9699: inst = 32'hc40484a;
      9700: inst = 32'h8220000;
      9701: inst = 32'h10408000;
      9702: inst = 32'hc40484b;
      9703: inst = 32'h8220000;
      9704: inst = 32'h10408000;
      9705: inst = 32'hc40484c;
      9706: inst = 32'h8220000;
      9707: inst = 32'h10408000;
      9708: inst = 32'hc40484d;
      9709: inst = 32'h8220000;
      9710: inst = 32'h10408000;
      9711: inst = 32'hc40484e;
      9712: inst = 32'h8220000;
      9713: inst = 32'h10408000;
      9714: inst = 32'hc40484f;
      9715: inst = 32'h8220000;
      9716: inst = 32'h10408000;
      9717: inst = 32'hc404850;
      9718: inst = 32'h8220000;
      9719: inst = 32'h10408000;
      9720: inst = 32'hc404851;
      9721: inst = 32'h8220000;
      9722: inst = 32'h10408000;
      9723: inst = 32'hc404852;
      9724: inst = 32'h8220000;
      9725: inst = 32'h10408000;
      9726: inst = 32'hc404853;
      9727: inst = 32'h8220000;
      9728: inst = 32'h10408000;
      9729: inst = 32'hc404854;
      9730: inst = 32'h8220000;
      9731: inst = 32'h10408000;
      9732: inst = 32'hc404855;
      9733: inst = 32'h8220000;
      9734: inst = 32'h10408000;
      9735: inst = 32'hc404856;
      9736: inst = 32'h8220000;
      9737: inst = 32'h10408000;
      9738: inst = 32'hc404857;
      9739: inst = 32'h8220000;
      9740: inst = 32'h10408000;
      9741: inst = 32'hc404858;
      9742: inst = 32'h8220000;
      9743: inst = 32'h10408000;
      9744: inst = 32'hc404859;
      9745: inst = 32'h8220000;
      9746: inst = 32'h10408000;
      9747: inst = 32'hc40485a;
      9748: inst = 32'h8220000;
      9749: inst = 32'h10408000;
      9750: inst = 32'hc40485b;
      9751: inst = 32'h8220000;
      9752: inst = 32'h10408000;
      9753: inst = 32'hc40485c;
      9754: inst = 32'h8220000;
      9755: inst = 32'h10408000;
      9756: inst = 32'hc40485d;
      9757: inst = 32'h8220000;
      9758: inst = 32'h10408000;
      9759: inst = 32'hc40485e;
      9760: inst = 32'h8220000;
      9761: inst = 32'h10408000;
      9762: inst = 32'hc40485f;
      9763: inst = 32'h8220000;
      9764: inst = 32'h10408000;
      9765: inst = 32'hc404860;
      9766: inst = 32'h8220000;
      9767: inst = 32'h10408000;
      9768: inst = 32'hc404861;
      9769: inst = 32'h8220000;
      9770: inst = 32'h10408000;
      9771: inst = 32'hc404862;
      9772: inst = 32'h8220000;
      9773: inst = 32'h10408000;
      9774: inst = 32'hc404863;
      9775: inst = 32'h8220000;
      9776: inst = 32'h10408000;
      9777: inst = 32'hc40489c;
      9778: inst = 32'h8220000;
      9779: inst = 32'h10408000;
      9780: inst = 32'hc40489d;
      9781: inst = 32'h8220000;
      9782: inst = 32'h10408000;
      9783: inst = 32'hc40489e;
      9784: inst = 32'h8220000;
      9785: inst = 32'h10408000;
      9786: inst = 32'hc40489f;
      9787: inst = 32'h8220000;
      9788: inst = 32'h10408000;
      9789: inst = 32'hc4048a0;
      9790: inst = 32'h8220000;
      9791: inst = 32'h10408000;
      9792: inst = 32'hc4048a1;
      9793: inst = 32'h8220000;
      9794: inst = 32'h10408000;
      9795: inst = 32'hc4048a2;
      9796: inst = 32'h8220000;
      9797: inst = 32'h10408000;
      9798: inst = 32'hc4048a3;
      9799: inst = 32'h8220000;
      9800: inst = 32'h10408000;
      9801: inst = 32'hc4048a4;
      9802: inst = 32'h8220000;
      9803: inst = 32'h10408000;
      9804: inst = 32'hc4048a5;
      9805: inst = 32'h8220000;
      9806: inst = 32'h10408000;
      9807: inst = 32'hc4048a6;
      9808: inst = 32'h8220000;
      9809: inst = 32'h10408000;
      9810: inst = 32'hc4048a7;
      9811: inst = 32'h8220000;
      9812: inst = 32'h10408000;
      9813: inst = 32'hc4048a8;
      9814: inst = 32'h8220000;
      9815: inst = 32'h10408000;
      9816: inst = 32'hc4048a9;
      9817: inst = 32'h8220000;
      9818: inst = 32'h10408000;
      9819: inst = 32'hc4048aa;
      9820: inst = 32'h8220000;
      9821: inst = 32'h10408000;
      9822: inst = 32'hc4048ab;
      9823: inst = 32'h8220000;
      9824: inst = 32'h10408000;
      9825: inst = 32'hc4048ac;
      9826: inst = 32'h8220000;
      9827: inst = 32'h10408000;
      9828: inst = 32'hc4048ad;
      9829: inst = 32'h8220000;
      9830: inst = 32'h10408000;
      9831: inst = 32'hc4048ae;
      9832: inst = 32'h8220000;
      9833: inst = 32'h10408000;
      9834: inst = 32'hc4048af;
      9835: inst = 32'h8220000;
      9836: inst = 32'h10408000;
      9837: inst = 32'hc4048b0;
      9838: inst = 32'h8220000;
      9839: inst = 32'h10408000;
      9840: inst = 32'hc4048b1;
      9841: inst = 32'h8220000;
      9842: inst = 32'h10408000;
      9843: inst = 32'hc4048b2;
      9844: inst = 32'h8220000;
      9845: inst = 32'h10408000;
      9846: inst = 32'hc4048b3;
      9847: inst = 32'h8220000;
      9848: inst = 32'h10408000;
      9849: inst = 32'hc4048b4;
      9850: inst = 32'h8220000;
      9851: inst = 32'h10408000;
      9852: inst = 32'hc4048b5;
      9853: inst = 32'h8220000;
      9854: inst = 32'h10408000;
      9855: inst = 32'hc4048b6;
      9856: inst = 32'h8220000;
      9857: inst = 32'h10408000;
      9858: inst = 32'hc4048b7;
      9859: inst = 32'h8220000;
      9860: inst = 32'h10408000;
      9861: inst = 32'hc4048b8;
      9862: inst = 32'h8220000;
      9863: inst = 32'h10408000;
      9864: inst = 32'hc4048b9;
      9865: inst = 32'h8220000;
      9866: inst = 32'h10408000;
      9867: inst = 32'hc4048ba;
      9868: inst = 32'h8220000;
      9869: inst = 32'h10408000;
      9870: inst = 32'hc4048bb;
      9871: inst = 32'h8220000;
      9872: inst = 32'h10408000;
      9873: inst = 32'hc4048bc;
      9874: inst = 32'h8220000;
      9875: inst = 32'h10408000;
      9876: inst = 32'hc4048bd;
      9877: inst = 32'h8220000;
      9878: inst = 32'h10408000;
      9879: inst = 32'hc4048be;
      9880: inst = 32'h8220000;
      9881: inst = 32'h10408000;
      9882: inst = 32'hc4048bf;
      9883: inst = 32'h8220000;
      9884: inst = 32'h10408000;
      9885: inst = 32'hc4048c0;
      9886: inst = 32'h8220000;
      9887: inst = 32'h10408000;
      9888: inst = 32'hc4048c1;
      9889: inst = 32'h8220000;
      9890: inst = 32'h10408000;
      9891: inst = 32'hc4048c2;
      9892: inst = 32'h8220000;
      9893: inst = 32'h10408000;
      9894: inst = 32'hc4048c3;
      9895: inst = 32'h8220000;
      9896: inst = 32'h10408000;
      9897: inst = 32'hc4048fc;
      9898: inst = 32'h8220000;
      9899: inst = 32'h10408000;
      9900: inst = 32'hc4048fd;
      9901: inst = 32'h8220000;
      9902: inst = 32'h10408000;
      9903: inst = 32'hc4048fe;
      9904: inst = 32'h8220000;
      9905: inst = 32'h10408000;
      9906: inst = 32'hc4048ff;
      9907: inst = 32'h8220000;
      9908: inst = 32'h10408000;
      9909: inst = 32'hc404900;
      9910: inst = 32'h8220000;
      9911: inst = 32'h10408000;
      9912: inst = 32'hc404901;
      9913: inst = 32'h8220000;
      9914: inst = 32'h10408000;
      9915: inst = 32'hc404902;
      9916: inst = 32'h8220000;
      9917: inst = 32'h10408000;
      9918: inst = 32'hc404903;
      9919: inst = 32'h8220000;
      9920: inst = 32'h10408000;
      9921: inst = 32'hc404904;
      9922: inst = 32'h8220000;
      9923: inst = 32'h10408000;
      9924: inst = 32'hc404905;
      9925: inst = 32'h8220000;
      9926: inst = 32'h10408000;
      9927: inst = 32'hc404906;
      9928: inst = 32'h8220000;
      9929: inst = 32'h10408000;
      9930: inst = 32'hc404907;
      9931: inst = 32'h8220000;
      9932: inst = 32'h10408000;
      9933: inst = 32'hc404908;
      9934: inst = 32'h8220000;
      9935: inst = 32'h10408000;
      9936: inst = 32'hc404909;
      9937: inst = 32'h8220000;
      9938: inst = 32'h10408000;
      9939: inst = 32'hc40490a;
      9940: inst = 32'h8220000;
      9941: inst = 32'h10408000;
      9942: inst = 32'hc40490b;
      9943: inst = 32'h8220000;
      9944: inst = 32'h10408000;
      9945: inst = 32'hc40490c;
      9946: inst = 32'h8220000;
      9947: inst = 32'h10408000;
      9948: inst = 32'hc40490d;
      9949: inst = 32'h8220000;
      9950: inst = 32'h10408000;
      9951: inst = 32'hc40490e;
      9952: inst = 32'h8220000;
      9953: inst = 32'h10408000;
      9954: inst = 32'hc40490f;
      9955: inst = 32'h8220000;
      9956: inst = 32'h10408000;
      9957: inst = 32'hc404910;
      9958: inst = 32'h8220000;
      9959: inst = 32'h10408000;
      9960: inst = 32'hc404911;
      9961: inst = 32'h8220000;
      9962: inst = 32'h10408000;
      9963: inst = 32'hc404912;
      9964: inst = 32'h8220000;
      9965: inst = 32'h10408000;
      9966: inst = 32'hc404913;
      9967: inst = 32'h8220000;
      9968: inst = 32'h10408000;
      9969: inst = 32'hc404914;
      9970: inst = 32'h8220000;
      9971: inst = 32'h10408000;
      9972: inst = 32'hc404915;
      9973: inst = 32'h8220000;
      9974: inst = 32'h10408000;
      9975: inst = 32'hc404916;
      9976: inst = 32'h8220000;
      9977: inst = 32'h10408000;
      9978: inst = 32'hc404917;
      9979: inst = 32'h8220000;
      9980: inst = 32'h10408000;
      9981: inst = 32'hc404918;
      9982: inst = 32'h8220000;
      9983: inst = 32'h10408000;
      9984: inst = 32'hc404919;
      9985: inst = 32'h8220000;
      9986: inst = 32'h10408000;
      9987: inst = 32'hc40491a;
      9988: inst = 32'h8220000;
      9989: inst = 32'h10408000;
      9990: inst = 32'hc40491b;
      9991: inst = 32'h8220000;
      9992: inst = 32'h10408000;
      9993: inst = 32'hc40491c;
      9994: inst = 32'h8220000;
      9995: inst = 32'h10408000;
      9996: inst = 32'hc40491d;
      9997: inst = 32'h8220000;
      9998: inst = 32'h10408000;
      9999: inst = 32'hc40491e;
      10000: inst = 32'h8220000;
      10001: inst = 32'h10408000;
      10002: inst = 32'hc40491f;
      10003: inst = 32'h8220000;
      10004: inst = 32'h10408000;
      10005: inst = 32'hc404920;
      10006: inst = 32'h8220000;
      10007: inst = 32'h10408000;
      10008: inst = 32'hc404921;
      10009: inst = 32'h8220000;
      10010: inst = 32'h10408000;
      10011: inst = 32'hc404922;
      10012: inst = 32'h8220000;
      10013: inst = 32'h10408000;
      10014: inst = 32'hc404923;
      10015: inst = 32'h8220000;
      10016: inst = 32'h10408000;
      10017: inst = 32'hc40495c;
      10018: inst = 32'h8220000;
      10019: inst = 32'h10408000;
      10020: inst = 32'hc40495d;
      10021: inst = 32'h8220000;
      10022: inst = 32'h10408000;
      10023: inst = 32'hc40495e;
      10024: inst = 32'h8220000;
      10025: inst = 32'h10408000;
      10026: inst = 32'hc40495f;
      10027: inst = 32'h8220000;
      10028: inst = 32'h10408000;
      10029: inst = 32'hc404960;
      10030: inst = 32'h8220000;
      10031: inst = 32'h10408000;
      10032: inst = 32'hc404961;
      10033: inst = 32'h8220000;
      10034: inst = 32'h10408000;
      10035: inst = 32'hc404962;
      10036: inst = 32'h8220000;
      10037: inst = 32'h10408000;
      10038: inst = 32'hc404963;
      10039: inst = 32'h8220000;
      10040: inst = 32'h10408000;
      10041: inst = 32'hc404964;
      10042: inst = 32'h8220000;
      10043: inst = 32'h10408000;
      10044: inst = 32'hc404965;
      10045: inst = 32'h8220000;
      10046: inst = 32'h10408000;
      10047: inst = 32'hc404966;
      10048: inst = 32'h8220000;
      10049: inst = 32'h10408000;
      10050: inst = 32'hc404967;
      10051: inst = 32'h8220000;
      10052: inst = 32'h10408000;
      10053: inst = 32'hc404968;
      10054: inst = 32'h8220000;
      10055: inst = 32'h10408000;
      10056: inst = 32'hc404969;
      10057: inst = 32'h8220000;
      10058: inst = 32'h10408000;
      10059: inst = 32'hc40496a;
      10060: inst = 32'h8220000;
      10061: inst = 32'h10408000;
      10062: inst = 32'hc40496b;
      10063: inst = 32'h8220000;
      10064: inst = 32'h10408000;
      10065: inst = 32'hc40496c;
      10066: inst = 32'h8220000;
      10067: inst = 32'h10408000;
      10068: inst = 32'hc40496d;
      10069: inst = 32'h8220000;
      10070: inst = 32'h10408000;
      10071: inst = 32'hc40496e;
      10072: inst = 32'h8220000;
      10073: inst = 32'h10408000;
      10074: inst = 32'hc40496f;
      10075: inst = 32'h8220000;
      10076: inst = 32'h10408000;
      10077: inst = 32'hc404970;
      10078: inst = 32'h8220000;
      10079: inst = 32'h10408000;
      10080: inst = 32'hc404971;
      10081: inst = 32'h8220000;
      10082: inst = 32'h10408000;
      10083: inst = 32'hc404972;
      10084: inst = 32'h8220000;
      10085: inst = 32'h10408000;
      10086: inst = 32'hc404973;
      10087: inst = 32'h8220000;
      10088: inst = 32'h10408000;
      10089: inst = 32'hc404974;
      10090: inst = 32'h8220000;
      10091: inst = 32'h10408000;
      10092: inst = 32'hc404975;
      10093: inst = 32'h8220000;
      10094: inst = 32'h10408000;
      10095: inst = 32'hc404976;
      10096: inst = 32'h8220000;
      10097: inst = 32'h10408000;
      10098: inst = 32'hc404977;
      10099: inst = 32'h8220000;
      10100: inst = 32'h10408000;
      10101: inst = 32'hc404978;
      10102: inst = 32'h8220000;
      10103: inst = 32'h10408000;
      10104: inst = 32'hc404979;
      10105: inst = 32'h8220000;
      10106: inst = 32'h10408000;
      10107: inst = 32'hc40497a;
      10108: inst = 32'h8220000;
      10109: inst = 32'h10408000;
      10110: inst = 32'hc40497b;
      10111: inst = 32'h8220000;
      10112: inst = 32'h10408000;
      10113: inst = 32'hc40497c;
      10114: inst = 32'h8220000;
      10115: inst = 32'h10408000;
      10116: inst = 32'hc40497d;
      10117: inst = 32'h8220000;
      10118: inst = 32'h10408000;
      10119: inst = 32'hc40497e;
      10120: inst = 32'h8220000;
      10121: inst = 32'h10408000;
      10122: inst = 32'hc40497f;
      10123: inst = 32'h8220000;
      10124: inst = 32'h10408000;
      10125: inst = 32'hc404980;
      10126: inst = 32'h8220000;
      10127: inst = 32'h10408000;
      10128: inst = 32'hc404981;
      10129: inst = 32'h8220000;
      10130: inst = 32'h10408000;
      10131: inst = 32'hc404982;
      10132: inst = 32'h8220000;
      10133: inst = 32'h10408000;
      10134: inst = 32'hc404983;
      10135: inst = 32'h8220000;
      10136: inst = 32'h10408000;
      10137: inst = 32'hc404992;
      10138: inst = 32'h8220000;
      10139: inst = 32'h10408000;
      10140: inst = 32'hc4049bc;
      10141: inst = 32'h8220000;
      10142: inst = 32'h10408000;
      10143: inst = 32'hc4049bd;
      10144: inst = 32'h8220000;
      10145: inst = 32'h10408000;
      10146: inst = 32'hc4049be;
      10147: inst = 32'h8220000;
      10148: inst = 32'h10408000;
      10149: inst = 32'hc4049bf;
      10150: inst = 32'h8220000;
      10151: inst = 32'h10408000;
      10152: inst = 32'hc4049c0;
      10153: inst = 32'h8220000;
      10154: inst = 32'h10408000;
      10155: inst = 32'hc4049c1;
      10156: inst = 32'h8220000;
      10157: inst = 32'h10408000;
      10158: inst = 32'hc4049c2;
      10159: inst = 32'h8220000;
      10160: inst = 32'h10408000;
      10161: inst = 32'hc4049c3;
      10162: inst = 32'h8220000;
      10163: inst = 32'h10408000;
      10164: inst = 32'hc4049c4;
      10165: inst = 32'h8220000;
      10166: inst = 32'h10408000;
      10167: inst = 32'hc4049c5;
      10168: inst = 32'h8220000;
      10169: inst = 32'h10408000;
      10170: inst = 32'hc4049c6;
      10171: inst = 32'h8220000;
      10172: inst = 32'h10408000;
      10173: inst = 32'hc4049c7;
      10174: inst = 32'h8220000;
      10175: inst = 32'h10408000;
      10176: inst = 32'hc4049c8;
      10177: inst = 32'h8220000;
      10178: inst = 32'h10408000;
      10179: inst = 32'hc4049c9;
      10180: inst = 32'h8220000;
      10181: inst = 32'h10408000;
      10182: inst = 32'hc4049ca;
      10183: inst = 32'h8220000;
      10184: inst = 32'h10408000;
      10185: inst = 32'hc4049cb;
      10186: inst = 32'h8220000;
      10187: inst = 32'h10408000;
      10188: inst = 32'hc4049cc;
      10189: inst = 32'h8220000;
      10190: inst = 32'h10408000;
      10191: inst = 32'hc4049cd;
      10192: inst = 32'h8220000;
      10193: inst = 32'h10408000;
      10194: inst = 32'hc4049ce;
      10195: inst = 32'h8220000;
      10196: inst = 32'h10408000;
      10197: inst = 32'hc4049cf;
      10198: inst = 32'h8220000;
      10199: inst = 32'h10408000;
      10200: inst = 32'hc4049d0;
      10201: inst = 32'h8220000;
      10202: inst = 32'h10408000;
      10203: inst = 32'hc4049d1;
      10204: inst = 32'h8220000;
      10205: inst = 32'h10408000;
      10206: inst = 32'hc4049d2;
      10207: inst = 32'h8220000;
      10208: inst = 32'h10408000;
      10209: inst = 32'hc4049d3;
      10210: inst = 32'h8220000;
      10211: inst = 32'h10408000;
      10212: inst = 32'hc4049d4;
      10213: inst = 32'h8220000;
      10214: inst = 32'h10408000;
      10215: inst = 32'hc4049d5;
      10216: inst = 32'h8220000;
      10217: inst = 32'h10408000;
      10218: inst = 32'hc4049d6;
      10219: inst = 32'h8220000;
      10220: inst = 32'h10408000;
      10221: inst = 32'hc4049d7;
      10222: inst = 32'h8220000;
      10223: inst = 32'h10408000;
      10224: inst = 32'hc4049d8;
      10225: inst = 32'h8220000;
      10226: inst = 32'h10408000;
      10227: inst = 32'hc4049d9;
      10228: inst = 32'h8220000;
      10229: inst = 32'h10408000;
      10230: inst = 32'hc4049da;
      10231: inst = 32'h8220000;
      10232: inst = 32'h10408000;
      10233: inst = 32'hc4049db;
      10234: inst = 32'h8220000;
      10235: inst = 32'h10408000;
      10236: inst = 32'hc4049dc;
      10237: inst = 32'h8220000;
      10238: inst = 32'h10408000;
      10239: inst = 32'hc4049dd;
      10240: inst = 32'h8220000;
      10241: inst = 32'h10408000;
      10242: inst = 32'hc4049de;
      10243: inst = 32'h8220000;
      10244: inst = 32'h10408000;
      10245: inst = 32'hc4049df;
      10246: inst = 32'h8220000;
      10247: inst = 32'h10408000;
      10248: inst = 32'hc4049e0;
      10249: inst = 32'h8220000;
      10250: inst = 32'h10408000;
      10251: inst = 32'hc4049e1;
      10252: inst = 32'h8220000;
      10253: inst = 32'h10408000;
      10254: inst = 32'hc4049e2;
      10255: inst = 32'h8220000;
      10256: inst = 32'h10408000;
      10257: inst = 32'hc4049e3;
      10258: inst = 32'h8220000;
      10259: inst = 32'h10408000;
      10260: inst = 32'hc4049f2;
      10261: inst = 32'h8220000;
      10262: inst = 32'h10408000;
      10263: inst = 32'hc404a1c;
      10264: inst = 32'h8220000;
      10265: inst = 32'h10408000;
      10266: inst = 32'hc404a1d;
      10267: inst = 32'h8220000;
      10268: inst = 32'h10408000;
      10269: inst = 32'hc404a1e;
      10270: inst = 32'h8220000;
      10271: inst = 32'h10408000;
      10272: inst = 32'hc404a1f;
      10273: inst = 32'h8220000;
      10274: inst = 32'h10408000;
      10275: inst = 32'hc404a20;
      10276: inst = 32'h8220000;
      10277: inst = 32'h10408000;
      10278: inst = 32'hc404a21;
      10279: inst = 32'h8220000;
      10280: inst = 32'h10408000;
      10281: inst = 32'hc404a22;
      10282: inst = 32'h8220000;
      10283: inst = 32'h10408000;
      10284: inst = 32'hc404a23;
      10285: inst = 32'h8220000;
      10286: inst = 32'h10408000;
      10287: inst = 32'hc404a24;
      10288: inst = 32'h8220000;
      10289: inst = 32'h10408000;
      10290: inst = 32'hc404a25;
      10291: inst = 32'h8220000;
      10292: inst = 32'h10408000;
      10293: inst = 32'hc404a26;
      10294: inst = 32'h8220000;
      10295: inst = 32'h10408000;
      10296: inst = 32'hc404a27;
      10297: inst = 32'h8220000;
      10298: inst = 32'h10408000;
      10299: inst = 32'hc404a28;
      10300: inst = 32'h8220000;
      10301: inst = 32'h10408000;
      10302: inst = 32'hc404a29;
      10303: inst = 32'h8220000;
      10304: inst = 32'h10408000;
      10305: inst = 32'hc404a2a;
      10306: inst = 32'h8220000;
      10307: inst = 32'h10408000;
      10308: inst = 32'hc404a2b;
      10309: inst = 32'h8220000;
      10310: inst = 32'h10408000;
      10311: inst = 32'hc404a2c;
      10312: inst = 32'h8220000;
      10313: inst = 32'h10408000;
      10314: inst = 32'hc404a2d;
      10315: inst = 32'h8220000;
      10316: inst = 32'h10408000;
      10317: inst = 32'hc404a2e;
      10318: inst = 32'h8220000;
      10319: inst = 32'h10408000;
      10320: inst = 32'hc404a2f;
      10321: inst = 32'h8220000;
      10322: inst = 32'h10408000;
      10323: inst = 32'hc404a30;
      10324: inst = 32'h8220000;
      10325: inst = 32'h10408000;
      10326: inst = 32'hc404a31;
      10327: inst = 32'h8220000;
      10328: inst = 32'h10408000;
      10329: inst = 32'hc404a32;
      10330: inst = 32'h8220000;
      10331: inst = 32'h10408000;
      10332: inst = 32'hc404a33;
      10333: inst = 32'h8220000;
      10334: inst = 32'h10408000;
      10335: inst = 32'hc404a34;
      10336: inst = 32'h8220000;
      10337: inst = 32'h10408000;
      10338: inst = 32'hc404a35;
      10339: inst = 32'h8220000;
      10340: inst = 32'h10408000;
      10341: inst = 32'hc404a36;
      10342: inst = 32'h8220000;
      10343: inst = 32'h10408000;
      10344: inst = 32'hc404a37;
      10345: inst = 32'h8220000;
      10346: inst = 32'h10408000;
      10347: inst = 32'hc404a38;
      10348: inst = 32'h8220000;
      10349: inst = 32'h10408000;
      10350: inst = 32'hc404a39;
      10351: inst = 32'h8220000;
      10352: inst = 32'h10408000;
      10353: inst = 32'hc404a3a;
      10354: inst = 32'h8220000;
      10355: inst = 32'h10408000;
      10356: inst = 32'hc404a3b;
      10357: inst = 32'h8220000;
      10358: inst = 32'h10408000;
      10359: inst = 32'hc404a3c;
      10360: inst = 32'h8220000;
      10361: inst = 32'h10408000;
      10362: inst = 32'hc404a3d;
      10363: inst = 32'h8220000;
      10364: inst = 32'h10408000;
      10365: inst = 32'hc404a3e;
      10366: inst = 32'h8220000;
      10367: inst = 32'h10408000;
      10368: inst = 32'hc404a3f;
      10369: inst = 32'h8220000;
      10370: inst = 32'h10408000;
      10371: inst = 32'hc404a40;
      10372: inst = 32'h8220000;
      10373: inst = 32'h10408000;
      10374: inst = 32'hc404a41;
      10375: inst = 32'h8220000;
      10376: inst = 32'h10408000;
      10377: inst = 32'hc404a42;
      10378: inst = 32'h8220000;
      10379: inst = 32'h10408000;
      10380: inst = 32'hc404a43;
      10381: inst = 32'h8220000;
      10382: inst = 32'h10408000;
      10383: inst = 32'hc404a52;
      10384: inst = 32'h8220000;
      10385: inst = 32'h10408000;
      10386: inst = 32'hc404a7c;
      10387: inst = 32'h8220000;
      10388: inst = 32'h10408000;
      10389: inst = 32'hc404a7d;
      10390: inst = 32'h8220000;
      10391: inst = 32'h10408000;
      10392: inst = 32'hc404a7e;
      10393: inst = 32'h8220000;
      10394: inst = 32'h10408000;
      10395: inst = 32'hc404a7f;
      10396: inst = 32'h8220000;
      10397: inst = 32'h10408000;
      10398: inst = 32'hc404a80;
      10399: inst = 32'h8220000;
      10400: inst = 32'h10408000;
      10401: inst = 32'hc404a81;
      10402: inst = 32'h8220000;
      10403: inst = 32'h10408000;
      10404: inst = 32'hc404a82;
      10405: inst = 32'h8220000;
      10406: inst = 32'h10408000;
      10407: inst = 32'hc404a83;
      10408: inst = 32'h8220000;
      10409: inst = 32'h10408000;
      10410: inst = 32'hc404a84;
      10411: inst = 32'h8220000;
      10412: inst = 32'h10408000;
      10413: inst = 32'hc404a85;
      10414: inst = 32'h8220000;
      10415: inst = 32'h10408000;
      10416: inst = 32'hc404a86;
      10417: inst = 32'h8220000;
      10418: inst = 32'h10408000;
      10419: inst = 32'hc404a87;
      10420: inst = 32'h8220000;
      10421: inst = 32'h10408000;
      10422: inst = 32'hc404a88;
      10423: inst = 32'h8220000;
      10424: inst = 32'h10408000;
      10425: inst = 32'hc404a89;
      10426: inst = 32'h8220000;
      10427: inst = 32'h10408000;
      10428: inst = 32'hc404a8a;
      10429: inst = 32'h8220000;
      10430: inst = 32'h10408000;
      10431: inst = 32'hc404a8b;
      10432: inst = 32'h8220000;
      10433: inst = 32'h10408000;
      10434: inst = 32'hc404a8c;
      10435: inst = 32'h8220000;
      10436: inst = 32'h10408000;
      10437: inst = 32'hc404a8d;
      10438: inst = 32'h8220000;
      10439: inst = 32'h10408000;
      10440: inst = 32'hc404a8e;
      10441: inst = 32'h8220000;
      10442: inst = 32'h10408000;
      10443: inst = 32'hc404a8f;
      10444: inst = 32'h8220000;
      10445: inst = 32'h10408000;
      10446: inst = 32'hc404a90;
      10447: inst = 32'h8220000;
      10448: inst = 32'h10408000;
      10449: inst = 32'hc404a91;
      10450: inst = 32'h8220000;
      10451: inst = 32'h10408000;
      10452: inst = 32'hc404a92;
      10453: inst = 32'h8220000;
      10454: inst = 32'h10408000;
      10455: inst = 32'hc404a93;
      10456: inst = 32'h8220000;
      10457: inst = 32'h10408000;
      10458: inst = 32'hc404a94;
      10459: inst = 32'h8220000;
      10460: inst = 32'h10408000;
      10461: inst = 32'hc404a95;
      10462: inst = 32'h8220000;
      10463: inst = 32'h10408000;
      10464: inst = 32'hc404a96;
      10465: inst = 32'h8220000;
      10466: inst = 32'h10408000;
      10467: inst = 32'hc404a97;
      10468: inst = 32'h8220000;
      10469: inst = 32'h10408000;
      10470: inst = 32'hc404a98;
      10471: inst = 32'h8220000;
      10472: inst = 32'h10408000;
      10473: inst = 32'hc404a99;
      10474: inst = 32'h8220000;
      10475: inst = 32'h10408000;
      10476: inst = 32'hc404a9a;
      10477: inst = 32'h8220000;
      10478: inst = 32'h10408000;
      10479: inst = 32'hc404a9b;
      10480: inst = 32'h8220000;
      10481: inst = 32'h10408000;
      10482: inst = 32'hc404a9c;
      10483: inst = 32'h8220000;
      10484: inst = 32'h10408000;
      10485: inst = 32'hc404a9d;
      10486: inst = 32'h8220000;
      10487: inst = 32'h10408000;
      10488: inst = 32'hc404a9e;
      10489: inst = 32'h8220000;
      10490: inst = 32'h10408000;
      10491: inst = 32'hc404a9f;
      10492: inst = 32'h8220000;
      10493: inst = 32'h10408000;
      10494: inst = 32'hc404aa0;
      10495: inst = 32'h8220000;
      10496: inst = 32'h10408000;
      10497: inst = 32'hc404aa1;
      10498: inst = 32'h8220000;
      10499: inst = 32'h10408000;
      10500: inst = 32'hc404aa2;
      10501: inst = 32'h8220000;
      10502: inst = 32'h10408000;
      10503: inst = 32'hc404aa3;
      10504: inst = 32'h8220000;
      10505: inst = 32'h10408000;
      10506: inst = 32'hc404ab4;
      10507: inst = 32'h8220000;
      10508: inst = 32'h10408000;
      10509: inst = 32'hc404adc;
      10510: inst = 32'h8220000;
      10511: inst = 32'h10408000;
      10512: inst = 32'hc404add;
      10513: inst = 32'h8220000;
      10514: inst = 32'h10408000;
      10515: inst = 32'hc404ade;
      10516: inst = 32'h8220000;
      10517: inst = 32'h10408000;
      10518: inst = 32'hc404adf;
      10519: inst = 32'h8220000;
      10520: inst = 32'h10408000;
      10521: inst = 32'hc404ae0;
      10522: inst = 32'h8220000;
      10523: inst = 32'h10408000;
      10524: inst = 32'hc404ae1;
      10525: inst = 32'h8220000;
      10526: inst = 32'h10408000;
      10527: inst = 32'hc404ae2;
      10528: inst = 32'h8220000;
      10529: inst = 32'h10408000;
      10530: inst = 32'hc404ae3;
      10531: inst = 32'h8220000;
      10532: inst = 32'h10408000;
      10533: inst = 32'hc404ae4;
      10534: inst = 32'h8220000;
      10535: inst = 32'h10408000;
      10536: inst = 32'hc404ae5;
      10537: inst = 32'h8220000;
      10538: inst = 32'h10408000;
      10539: inst = 32'hc404ae6;
      10540: inst = 32'h8220000;
      10541: inst = 32'h10408000;
      10542: inst = 32'hc404ae7;
      10543: inst = 32'h8220000;
      10544: inst = 32'h10408000;
      10545: inst = 32'hc404ae8;
      10546: inst = 32'h8220000;
      10547: inst = 32'h10408000;
      10548: inst = 32'hc404ae9;
      10549: inst = 32'h8220000;
      10550: inst = 32'h10408000;
      10551: inst = 32'hc404aea;
      10552: inst = 32'h8220000;
      10553: inst = 32'h10408000;
      10554: inst = 32'hc404aeb;
      10555: inst = 32'h8220000;
      10556: inst = 32'h10408000;
      10557: inst = 32'hc404aec;
      10558: inst = 32'h8220000;
      10559: inst = 32'h10408000;
      10560: inst = 32'hc404aed;
      10561: inst = 32'h8220000;
      10562: inst = 32'h10408000;
      10563: inst = 32'hc404aee;
      10564: inst = 32'h8220000;
      10565: inst = 32'h10408000;
      10566: inst = 32'hc404aef;
      10567: inst = 32'h8220000;
      10568: inst = 32'h10408000;
      10569: inst = 32'hc404af0;
      10570: inst = 32'h8220000;
      10571: inst = 32'h10408000;
      10572: inst = 32'hc404af1;
      10573: inst = 32'h8220000;
      10574: inst = 32'h10408000;
      10575: inst = 32'hc404af2;
      10576: inst = 32'h8220000;
      10577: inst = 32'h10408000;
      10578: inst = 32'hc404af3;
      10579: inst = 32'h8220000;
      10580: inst = 32'h10408000;
      10581: inst = 32'hc404af4;
      10582: inst = 32'h8220000;
      10583: inst = 32'h10408000;
      10584: inst = 32'hc404af5;
      10585: inst = 32'h8220000;
      10586: inst = 32'h10408000;
      10587: inst = 32'hc404af6;
      10588: inst = 32'h8220000;
      10589: inst = 32'h10408000;
      10590: inst = 32'hc404af7;
      10591: inst = 32'h8220000;
      10592: inst = 32'h10408000;
      10593: inst = 32'hc404af8;
      10594: inst = 32'h8220000;
      10595: inst = 32'h10408000;
      10596: inst = 32'hc404af9;
      10597: inst = 32'h8220000;
      10598: inst = 32'h10408000;
      10599: inst = 32'hc404afa;
      10600: inst = 32'h8220000;
      10601: inst = 32'h10408000;
      10602: inst = 32'hc404afb;
      10603: inst = 32'h8220000;
      10604: inst = 32'h10408000;
      10605: inst = 32'hc404afc;
      10606: inst = 32'h8220000;
      10607: inst = 32'h10408000;
      10608: inst = 32'hc404afd;
      10609: inst = 32'h8220000;
      10610: inst = 32'h10408000;
      10611: inst = 32'hc404afe;
      10612: inst = 32'h8220000;
      10613: inst = 32'h10408000;
      10614: inst = 32'hc404aff;
      10615: inst = 32'h8220000;
      10616: inst = 32'h10408000;
      10617: inst = 32'hc404b00;
      10618: inst = 32'h8220000;
      10619: inst = 32'h10408000;
      10620: inst = 32'hc404b01;
      10621: inst = 32'h8220000;
      10622: inst = 32'h10408000;
      10623: inst = 32'hc404b02;
      10624: inst = 32'h8220000;
      10625: inst = 32'h10408000;
      10626: inst = 32'hc404b03;
      10627: inst = 32'h8220000;
      10628: inst = 32'h10408000;
      10629: inst = 32'hc404b14;
      10630: inst = 32'h8220000;
      10631: inst = 32'h10408000;
      10632: inst = 32'hc404b3c;
      10633: inst = 32'h8220000;
      10634: inst = 32'h10408000;
      10635: inst = 32'hc404b3d;
      10636: inst = 32'h8220000;
      10637: inst = 32'h10408000;
      10638: inst = 32'hc404b3e;
      10639: inst = 32'h8220000;
      10640: inst = 32'h10408000;
      10641: inst = 32'hc404b3f;
      10642: inst = 32'h8220000;
      10643: inst = 32'h10408000;
      10644: inst = 32'hc404b40;
      10645: inst = 32'h8220000;
      10646: inst = 32'h10408000;
      10647: inst = 32'hc404b41;
      10648: inst = 32'h8220000;
      10649: inst = 32'h10408000;
      10650: inst = 32'hc404b42;
      10651: inst = 32'h8220000;
      10652: inst = 32'h10408000;
      10653: inst = 32'hc404b43;
      10654: inst = 32'h8220000;
      10655: inst = 32'h10408000;
      10656: inst = 32'hc404b44;
      10657: inst = 32'h8220000;
      10658: inst = 32'h10408000;
      10659: inst = 32'hc404b45;
      10660: inst = 32'h8220000;
      10661: inst = 32'h10408000;
      10662: inst = 32'hc404b46;
      10663: inst = 32'h8220000;
      10664: inst = 32'h10408000;
      10665: inst = 32'hc404b47;
      10666: inst = 32'h8220000;
      10667: inst = 32'h10408000;
      10668: inst = 32'hc404b48;
      10669: inst = 32'h8220000;
      10670: inst = 32'h10408000;
      10671: inst = 32'hc404b49;
      10672: inst = 32'h8220000;
      10673: inst = 32'h10408000;
      10674: inst = 32'hc404b4a;
      10675: inst = 32'h8220000;
      10676: inst = 32'h10408000;
      10677: inst = 32'hc404b4b;
      10678: inst = 32'h8220000;
      10679: inst = 32'h10408000;
      10680: inst = 32'hc404b4c;
      10681: inst = 32'h8220000;
      10682: inst = 32'h10408000;
      10683: inst = 32'hc404b4d;
      10684: inst = 32'h8220000;
      10685: inst = 32'h10408000;
      10686: inst = 32'hc404b4e;
      10687: inst = 32'h8220000;
      10688: inst = 32'h10408000;
      10689: inst = 32'hc404b4f;
      10690: inst = 32'h8220000;
      10691: inst = 32'h10408000;
      10692: inst = 32'hc404b50;
      10693: inst = 32'h8220000;
      10694: inst = 32'h10408000;
      10695: inst = 32'hc404b51;
      10696: inst = 32'h8220000;
      10697: inst = 32'h10408000;
      10698: inst = 32'hc404b52;
      10699: inst = 32'h8220000;
      10700: inst = 32'h10408000;
      10701: inst = 32'hc404b53;
      10702: inst = 32'h8220000;
      10703: inst = 32'h10408000;
      10704: inst = 32'hc404b54;
      10705: inst = 32'h8220000;
      10706: inst = 32'h10408000;
      10707: inst = 32'hc404b55;
      10708: inst = 32'h8220000;
      10709: inst = 32'h10408000;
      10710: inst = 32'hc404b56;
      10711: inst = 32'h8220000;
      10712: inst = 32'h10408000;
      10713: inst = 32'hc404b57;
      10714: inst = 32'h8220000;
      10715: inst = 32'h10408000;
      10716: inst = 32'hc404b58;
      10717: inst = 32'h8220000;
      10718: inst = 32'h10408000;
      10719: inst = 32'hc404b59;
      10720: inst = 32'h8220000;
      10721: inst = 32'h10408000;
      10722: inst = 32'hc404b5a;
      10723: inst = 32'h8220000;
      10724: inst = 32'h10408000;
      10725: inst = 32'hc404b5b;
      10726: inst = 32'h8220000;
      10727: inst = 32'h10408000;
      10728: inst = 32'hc404b5c;
      10729: inst = 32'h8220000;
      10730: inst = 32'h10408000;
      10731: inst = 32'hc404b5d;
      10732: inst = 32'h8220000;
      10733: inst = 32'h10408000;
      10734: inst = 32'hc404b5e;
      10735: inst = 32'h8220000;
      10736: inst = 32'h10408000;
      10737: inst = 32'hc404b5f;
      10738: inst = 32'h8220000;
      10739: inst = 32'h10408000;
      10740: inst = 32'hc404b60;
      10741: inst = 32'h8220000;
      10742: inst = 32'h10408000;
      10743: inst = 32'hc404b61;
      10744: inst = 32'h8220000;
      10745: inst = 32'h10408000;
      10746: inst = 32'hc404b62;
      10747: inst = 32'h8220000;
      10748: inst = 32'h10408000;
      10749: inst = 32'hc404b63;
      10750: inst = 32'h8220000;
      10751: inst = 32'h10408000;
      10752: inst = 32'hc404b9c;
      10753: inst = 32'h8220000;
      10754: inst = 32'h10408000;
      10755: inst = 32'hc404b9d;
      10756: inst = 32'h8220000;
      10757: inst = 32'h10408000;
      10758: inst = 32'hc404b9e;
      10759: inst = 32'h8220000;
      10760: inst = 32'h10408000;
      10761: inst = 32'hc404b9f;
      10762: inst = 32'h8220000;
      10763: inst = 32'h10408000;
      10764: inst = 32'hc404ba0;
      10765: inst = 32'h8220000;
      10766: inst = 32'h10408000;
      10767: inst = 32'hc404ba1;
      10768: inst = 32'h8220000;
      10769: inst = 32'h10408000;
      10770: inst = 32'hc404ba2;
      10771: inst = 32'h8220000;
      10772: inst = 32'h10408000;
      10773: inst = 32'hc404ba3;
      10774: inst = 32'h8220000;
      10775: inst = 32'h10408000;
      10776: inst = 32'hc404ba4;
      10777: inst = 32'h8220000;
      10778: inst = 32'h10408000;
      10779: inst = 32'hc404ba5;
      10780: inst = 32'h8220000;
      10781: inst = 32'h10408000;
      10782: inst = 32'hc404ba6;
      10783: inst = 32'h8220000;
      10784: inst = 32'h10408000;
      10785: inst = 32'hc404ba7;
      10786: inst = 32'h8220000;
      10787: inst = 32'h10408000;
      10788: inst = 32'hc404ba8;
      10789: inst = 32'h8220000;
      10790: inst = 32'h10408000;
      10791: inst = 32'hc404ba9;
      10792: inst = 32'h8220000;
      10793: inst = 32'h10408000;
      10794: inst = 32'hc404baa;
      10795: inst = 32'h8220000;
      10796: inst = 32'h10408000;
      10797: inst = 32'hc404bab;
      10798: inst = 32'h8220000;
      10799: inst = 32'h10408000;
      10800: inst = 32'hc404bac;
      10801: inst = 32'h8220000;
      10802: inst = 32'h10408000;
      10803: inst = 32'hc404bad;
      10804: inst = 32'h8220000;
      10805: inst = 32'h10408000;
      10806: inst = 32'hc404bae;
      10807: inst = 32'h8220000;
      10808: inst = 32'h10408000;
      10809: inst = 32'hc404baf;
      10810: inst = 32'h8220000;
      10811: inst = 32'h10408000;
      10812: inst = 32'hc404bb0;
      10813: inst = 32'h8220000;
      10814: inst = 32'h10408000;
      10815: inst = 32'hc404bb1;
      10816: inst = 32'h8220000;
      10817: inst = 32'h10408000;
      10818: inst = 32'hc404bb2;
      10819: inst = 32'h8220000;
      10820: inst = 32'h10408000;
      10821: inst = 32'hc404bb3;
      10822: inst = 32'h8220000;
      10823: inst = 32'h10408000;
      10824: inst = 32'hc404bb4;
      10825: inst = 32'h8220000;
      10826: inst = 32'h10408000;
      10827: inst = 32'hc404bb5;
      10828: inst = 32'h8220000;
      10829: inst = 32'h10408000;
      10830: inst = 32'hc404bb6;
      10831: inst = 32'h8220000;
      10832: inst = 32'h10408000;
      10833: inst = 32'hc404bb7;
      10834: inst = 32'h8220000;
      10835: inst = 32'h10408000;
      10836: inst = 32'hc404bb8;
      10837: inst = 32'h8220000;
      10838: inst = 32'h10408000;
      10839: inst = 32'hc404bb9;
      10840: inst = 32'h8220000;
      10841: inst = 32'h10408000;
      10842: inst = 32'hc404bba;
      10843: inst = 32'h8220000;
      10844: inst = 32'h10408000;
      10845: inst = 32'hc404bbb;
      10846: inst = 32'h8220000;
      10847: inst = 32'h10408000;
      10848: inst = 32'hc404bbc;
      10849: inst = 32'h8220000;
      10850: inst = 32'h10408000;
      10851: inst = 32'hc404bbd;
      10852: inst = 32'h8220000;
      10853: inst = 32'h10408000;
      10854: inst = 32'hc404bbe;
      10855: inst = 32'h8220000;
      10856: inst = 32'h10408000;
      10857: inst = 32'hc404bbf;
      10858: inst = 32'h8220000;
      10859: inst = 32'h10408000;
      10860: inst = 32'hc404bc0;
      10861: inst = 32'h8220000;
      10862: inst = 32'h10408000;
      10863: inst = 32'hc404bc1;
      10864: inst = 32'h8220000;
      10865: inst = 32'h10408000;
      10866: inst = 32'hc404bc2;
      10867: inst = 32'h8220000;
      10868: inst = 32'h10408000;
      10869: inst = 32'hc404bc3;
      10870: inst = 32'h8220000;
      10871: inst = 32'hc20ee75;
      10872: inst = 32'h10408000;
      10873: inst = 32'hc4042ea;
      10874: inst = 32'h8220000;
      10875: inst = 32'h10408000;
      10876: inst = 32'hc4043a7;
      10877: inst = 32'h8220000;
      10878: inst = 32'hc20d42c;
      10879: inst = 32'h10408000;
      10880: inst = 32'hc4042eb;
      10881: inst = 32'h8220000;
      10882: inst = 32'h10408000;
      10883: inst = 32'hc4042ec;
      10884: inst = 32'h8220000;
      10885: inst = 32'h10408000;
      10886: inst = 32'hc4043a8;
      10887: inst = 32'h8220000;
      10888: inst = 32'hc20ee55;
      10889: inst = 32'h10408000;
      10890: inst = 32'hc4042ed;
      10891: inst = 32'h8220000;
      10892: inst = 32'h10408000;
      10893: inst = 32'hc4043b0;
      10894: inst = 32'h8220000;
      10895: inst = 32'hc20e571;
      10896: inst = 32'h10408000;
      10897: inst = 32'hc404349;
      10898: inst = 32'h8220000;
      10899: inst = 32'h10408000;
      10900: inst = 32'hc40434e;
      10901: inst = 32'h8220000;
      10902: inst = 32'h10408000;
      10903: inst = 32'hc404406;
      10904: inst = 32'h8220000;
      10905: inst = 32'h10408000;
      10906: inst = 32'hc404411;
      10907: inst = 32'h8220000;
      10908: inst = 32'hc20cb28;
      10909: inst = 32'h10408000;
      10910: inst = 32'hc40434a;
      10911: inst = 32'h8220000;
      10912: inst = 32'h10408000;
      10913: inst = 32'hc40434d;
      10914: inst = 32'h8220000;
      10915: inst = 32'h10408000;
      10916: inst = 32'hc404407;
      10917: inst = 32'h8220000;
      10918: inst = 32'h10408000;
      10919: inst = 32'hc404410;
      10920: inst = 32'h8220000;
      10921: inst = 32'hc20cac7;
      10922: inst = 32'h10408000;
      10923: inst = 32'hc40434b;
      10924: inst = 32'h8220000;
      10925: inst = 32'h10408000;
      10926: inst = 32'hc40434c;
      10927: inst = 32'h8220000;
      10928: inst = 32'h10408000;
      10929: inst = 32'hc4043a9;
      10930: inst = 32'h8220000;
      10931: inst = 32'h10408000;
      10932: inst = 32'hc4043aa;
      10933: inst = 32'h8220000;
      10934: inst = 32'h10408000;
      10935: inst = 32'hc4043ab;
      10936: inst = 32'h8220000;
      10937: inst = 32'h10408000;
      10938: inst = 32'hc4043ac;
      10939: inst = 32'h8220000;
      10940: inst = 32'h10408000;
      10941: inst = 32'hc4043ad;
      10942: inst = 32'h8220000;
      10943: inst = 32'h10408000;
      10944: inst = 32'hc4043ae;
      10945: inst = 32'h8220000;
      10946: inst = 32'h10408000;
      10947: inst = 32'hc404408;
      10948: inst = 32'h8220000;
      10949: inst = 32'h10408000;
      10950: inst = 32'hc404409;
      10951: inst = 32'h8220000;
      10952: inst = 32'h10408000;
      10953: inst = 32'hc40440a;
      10954: inst = 32'h8220000;
      10955: inst = 32'h10408000;
      10956: inst = 32'hc40440b;
      10957: inst = 32'h8220000;
      10958: inst = 32'h10408000;
      10959: inst = 32'hc40440c;
      10960: inst = 32'h8220000;
      10961: inst = 32'h10408000;
      10962: inst = 32'hc40440d;
      10963: inst = 32'h8220000;
      10964: inst = 32'h10408000;
      10965: inst = 32'hc40440e;
      10966: inst = 32'h8220000;
      10967: inst = 32'h10408000;
      10968: inst = 32'hc40440f;
      10969: inst = 32'h8220000;
      10970: inst = 32'hc20d40c;
      10971: inst = 32'h10408000;
      10972: inst = 32'hc4043af;
      10973: inst = 32'h8220000;
      10974: inst = 32'hc20ee8e;
      10975: inst = 32'h10408000;
      10976: inst = 32'hc40446a;
      10977: inst = 32'h8220000;
      10978: inst = 32'h10408000;
      10979: inst = 32'hc4044b5;
      10980: inst = 32'h8220000;
      10981: inst = 32'hc20ee48;
      10982: inst = 32'h10408000;
      10983: inst = 32'hc40446b;
      10984: inst = 32'h8220000;
      10985: inst = 32'h10408000;
      10986: inst = 32'hc40446c;
      10987: inst = 32'h8220000;
      10988: inst = 32'h10408000;
      10989: inst = 32'hc4044b3;
      10990: inst = 32'h8220000;
      10991: inst = 32'h10408000;
      10992: inst = 32'hc4044b4;
      10993: inst = 32'h8220000;
      10994: inst = 32'hc20ee90;
      10995: inst = 32'h10408000;
      10996: inst = 32'hc40446d;
      10997: inst = 32'h8220000;
      10998: inst = 32'h10408000;
      10999: inst = 32'hc4044b2;
      11000: inst = 32'h8220000;
      11001: inst = 32'hc20eeb5;
      11002: inst = 32'h10408000;
      11003: inst = 32'hc4044cb;
      11004: inst = 32'h8220000;
      11005: inst = 32'h10408000;
      11006: inst = 32'hc4044cc;
      11007: inst = 32'h8220000;
      11008: inst = 32'h10408000;
      11009: inst = 32'hc404513;
      11010: inst = 32'h8220000;
      11011: inst = 32'h10408000;
      11012: inst = 32'hc404514;
      11013: inst = 32'h8220000;
      11014: inst = 32'hc20c2e2;
      11015: inst = 32'h10408000;
      11016: inst = 32'hc4046ef;
      11017: inst = 32'h8220000;
      11018: inst = 32'h10408000;
      11019: inst = 32'hc4046f0;
      11020: inst = 32'h8220000;
      11021: inst = 32'h10408000;
      11022: inst = 32'hc4046f1;
      11023: inst = 32'h8220000;
      11024: inst = 32'h10408000;
      11025: inst = 32'hc4046f2;
      11026: inst = 32'h8220000;
      11027: inst = 32'h10408000;
      11028: inst = 32'hc4046f3;
      11029: inst = 32'h8220000;
      11030: inst = 32'h10408000;
      11031: inst = 32'hc4046f4;
      11032: inst = 32'h8220000;
      11033: inst = 32'h10408000;
      11034: inst = 32'hc4046f5;
      11035: inst = 32'h8220000;
      11036: inst = 32'h10408000;
      11037: inst = 32'hc4046f6;
      11038: inst = 32'h8220000;
      11039: inst = 32'h10408000;
      11040: inst = 32'hc4046f7;
      11041: inst = 32'h8220000;
      11042: inst = 32'h10408000;
      11043: inst = 32'hc4046f8;
      11044: inst = 32'h8220000;
      11045: inst = 32'h10408000;
      11046: inst = 32'hc4046f9;
      11047: inst = 32'h8220000;
      11048: inst = 32'h10408000;
      11049: inst = 32'hc4046fa;
      11050: inst = 32'h8220000;
      11051: inst = 32'h10408000;
      11052: inst = 32'hc4046fb;
      11053: inst = 32'h8220000;
      11054: inst = 32'h10408000;
      11055: inst = 32'hc4046fc;
      11056: inst = 32'h8220000;
      11057: inst = 32'h10408000;
      11058: inst = 32'hc4046fd;
      11059: inst = 32'h8220000;
      11060: inst = 32'h10408000;
      11061: inst = 32'hc4046fe;
      11062: inst = 32'h8220000;
      11063: inst = 32'h10408000;
      11064: inst = 32'hc4046ff;
      11065: inst = 32'h8220000;
      11066: inst = 32'h10408000;
      11067: inst = 32'hc40474f;
      11068: inst = 32'h8220000;
      11069: inst = 32'h10408000;
      11070: inst = 32'hc40475f;
      11071: inst = 32'h8220000;
      11072: inst = 32'h10408000;
      11073: inst = 32'hc4047af;
      11074: inst = 32'h8220000;
      11075: inst = 32'h10408000;
      11076: inst = 32'hc4047bf;
      11077: inst = 32'h8220000;
      11078: inst = 32'h10408000;
      11079: inst = 32'hc40480f;
      11080: inst = 32'h8220000;
      11081: inst = 32'h10408000;
      11082: inst = 32'hc40481f;
      11083: inst = 32'h8220000;
      11084: inst = 32'h10408000;
      11085: inst = 32'hc40486f;
      11086: inst = 32'h8220000;
      11087: inst = 32'h10408000;
      11088: inst = 32'hc40487f;
      11089: inst = 32'h8220000;
      11090: inst = 32'h10408000;
      11091: inst = 32'hc4048cf;
      11092: inst = 32'h8220000;
      11093: inst = 32'h10408000;
      11094: inst = 32'hc4048df;
      11095: inst = 32'h8220000;
      11096: inst = 32'h10408000;
      11097: inst = 32'hc40492f;
      11098: inst = 32'h8220000;
      11099: inst = 32'h10408000;
      11100: inst = 32'hc40493f;
      11101: inst = 32'h8220000;
      11102: inst = 32'h10408000;
      11103: inst = 32'hc40498f;
      11104: inst = 32'h8220000;
      11105: inst = 32'h10408000;
      11106: inst = 32'hc40499f;
      11107: inst = 32'h8220000;
      11108: inst = 32'h10408000;
      11109: inst = 32'hc4049ef;
      11110: inst = 32'h8220000;
      11111: inst = 32'h10408000;
      11112: inst = 32'hc4049ff;
      11113: inst = 32'h8220000;
      11114: inst = 32'h10408000;
      11115: inst = 32'hc404a4f;
      11116: inst = 32'h8220000;
      11117: inst = 32'h10408000;
      11118: inst = 32'hc404a5f;
      11119: inst = 32'h8220000;
      11120: inst = 32'h10408000;
      11121: inst = 32'hc404aaf;
      11122: inst = 32'h8220000;
      11123: inst = 32'h10408000;
      11124: inst = 32'hc404abf;
      11125: inst = 32'h8220000;
      11126: inst = 32'h10408000;
      11127: inst = 32'hc404b0f;
      11128: inst = 32'h8220000;
      11129: inst = 32'h10408000;
      11130: inst = 32'hc404b1f;
      11131: inst = 32'h8220000;
      11132: inst = 32'h10408000;
      11133: inst = 32'hc404b6f;
      11134: inst = 32'h8220000;
      11135: inst = 32'h10408000;
      11136: inst = 32'hc404b7f;
      11137: inst = 32'h8220000;
      11138: inst = 32'h10408000;
      11139: inst = 32'hc404bcf;
      11140: inst = 32'h8220000;
      11141: inst = 32'h10408000;
      11142: inst = 32'hc404bdf;
      11143: inst = 32'h8220000;
      11144: inst = 32'h10408000;
      11145: inst = 32'hc404c2f;
      11146: inst = 32'h8220000;
      11147: inst = 32'h10408000;
      11148: inst = 32'hc404c3f;
      11149: inst = 32'h8220000;
      11150: inst = 32'h10408000;
      11151: inst = 32'hc404c8f;
      11152: inst = 32'h8220000;
      11153: inst = 32'h10408000;
      11154: inst = 32'hc404c9f;
      11155: inst = 32'h8220000;
      11156: inst = 32'h10408000;
      11157: inst = 32'hc404cef;
      11158: inst = 32'h8220000;
      11159: inst = 32'h10408000;
      11160: inst = 32'hc404cff;
      11161: inst = 32'h8220000;
      11162: inst = 32'h10408000;
      11163: inst = 32'hc404d4f;
      11164: inst = 32'h8220000;
      11165: inst = 32'h10408000;
      11166: inst = 32'hc404d5f;
      11167: inst = 32'h8220000;
      11168: inst = 32'h10408000;
      11169: inst = 32'hc404daf;
      11170: inst = 32'h8220000;
      11171: inst = 32'h10408000;
      11172: inst = 32'hc404dbf;
      11173: inst = 32'h8220000;
      11174: inst = 32'h10408000;
      11175: inst = 32'hc404e0f;
      11176: inst = 32'h8220000;
      11177: inst = 32'h10408000;
      11178: inst = 32'hc404e1f;
      11179: inst = 32'h8220000;
      11180: inst = 32'h10408000;
      11181: inst = 32'hc404e6f;
      11182: inst = 32'h8220000;
      11183: inst = 32'h10408000;
      11184: inst = 32'hc404e7f;
      11185: inst = 32'h8220000;
      11186: inst = 32'h10408000;
      11187: inst = 32'hc404ecf;
      11188: inst = 32'h8220000;
      11189: inst = 32'h10408000;
      11190: inst = 32'hc404edf;
      11191: inst = 32'h8220000;
      11192: inst = 32'h10408000;
      11193: inst = 32'hc404f2f;
      11194: inst = 32'h8220000;
      11195: inst = 32'h10408000;
      11196: inst = 32'hc404f3f;
      11197: inst = 32'h8220000;
      11198: inst = 32'h10408000;
      11199: inst = 32'hc404f8f;
      11200: inst = 32'h8220000;
      11201: inst = 32'h10408000;
      11202: inst = 32'hc404f9f;
      11203: inst = 32'h8220000;
      11204: inst = 32'h10408000;
      11205: inst = 32'hc404fef;
      11206: inst = 32'h8220000;
      11207: inst = 32'h10408000;
      11208: inst = 32'hc404fff;
      11209: inst = 32'h8220000;
      11210: inst = 32'h10408000;
      11211: inst = 32'hc40504f;
      11212: inst = 32'h8220000;
      11213: inst = 32'h10408000;
      11214: inst = 32'hc40505f;
      11215: inst = 32'h8220000;
      11216: inst = 32'h10408000;
      11217: inst = 32'hc4050af;
      11218: inst = 32'h8220000;
      11219: inst = 32'h10408000;
      11220: inst = 32'hc4050bf;
      11221: inst = 32'h8220000;
      11222: inst = 32'h10408000;
      11223: inst = 32'hc40510f;
      11224: inst = 32'h8220000;
      11225: inst = 32'h10408000;
      11226: inst = 32'hc40511f;
      11227: inst = 32'h8220000;
      11228: inst = 32'h10408000;
      11229: inst = 32'hc40516f;
      11230: inst = 32'h8220000;
      11231: inst = 32'h10408000;
      11232: inst = 32'hc40517f;
      11233: inst = 32'h8220000;
      11234: inst = 32'h10408000;
      11235: inst = 32'hc4051cf;
      11236: inst = 32'h8220000;
      11237: inst = 32'h10408000;
      11238: inst = 32'hc4051df;
      11239: inst = 32'h8220000;
      11240: inst = 32'h10408000;
      11241: inst = 32'hc40522f;
      11242: inst = 32'h8220000;
      11243: inst = 32'h10408000;
      11244: inst = 32'hc40523f;
      11245: inst = 32'h8220000;
      11246: inst = 32'h10408000;
      11247: inst = 32'hc40528f;
      11248: inst = 32'h8220000;
      11249: inst = 32'h10408000;
      11250: inst = 32'hc40529f;
      11251: inst = 32'h8220000;
      11252: inst = 32'h10408000;
      11253: inst = 32'hc4052ef;
      11254: inst = 32'h8220000;
      11255: inst = 32'h10408000;
      11256: inst = 32'hc4052f0;
      11257: inst = 32'h8220000;
      11258: inst = 32'h10408000;
      11259: inst = 32'hc4052f1;
      11260: inst = 32'h8220000;
      11261: inst = 32'h10408000;
      11262: inst = 32'hc4052f2;
      11263: inst = 32'h8220000;
      11264: inst = 32'h10408000;
      11265: inst = 32'hc4052f3;
      11266: inst = 32'h8220000;
      11267: inst = 32'h10408000;
      11268: inst = 32'hc4052f4;
      11269: inst = 32'h8220000;
      11270: inst = 32'h10408000;
      11271: inst = 32'hc4052f5;
      11272: inst = 32'h8220000;
      11273: inst = 32'h10408000;
      11274: inst = 32'hc4052f6;
      11275: inst = 32'h8220000;
      11276: inst = 32'h10408000;
      11277: inst = 32'hc4052f7;
      11278: inst = 32'h8220000;
      11279: inst = 32'h10408000;
      11280: inst = 32'hc4052f8;
      11281: inst = 32'h8220000;
      11282: inst = 32'h10408000;
      11283: inst = 32'hc4052f9;
      11284: inst = 32'h8220000;
      11285: inst = 32'h10408000;
      11286: inst = 32'hc4052fa;
      11287: inst = 32'h8220000;
      11288: inst = 32'h10408000;
      11289: inst = 32'hc4052fb;
      11290: inst = 32'h8220000;
      11291: inst = 32'h10408000;
      11292: inst = 32'hc4052fc;
      11293: inst = 32'h8220000;
      11294: inst = 32'h10408000;
      11295: inst = 32'hc4052fd;
      11296: inst = 32'h8220000;
      11297: inst = 32'h10408000;
      11298: inst = 32'hc4052fe;
      11299: inst = 32'h8220000;
      11300: inst = 32'h10408000;
      11301: inst = 32'hc4052ff;
      11302: inst = 32'h8220000;
      11303: inst = 32'hc20dbc5;
      11304: inst = 32'h10408000;
      11305: inst = 32'hc404750;
      11306: inst = 32'h8220000;
      11307: inst = 32'h10408000;
      11308: inst = 32'hc404751;
      11309: inst = 32'h8220000;
      11310: inst = 32'h10408000;
      11311: inst = 32'hc404752;
      11312: inst = 32'h8220000;
      11313: inst = 32'h10408000;
      11314: inst = 32'hc404753;
      11315: inst = 32'h8220000;
      11316: inst = 32'h10408000;
      11317: inst = 32'hc404754;
      11318: inst = 32'h8220000;
      11319: inst = 32'h10408000;
      11320: inst = 32'hc404755;
      11321: inst = 32'h8220000;
      11322: inst = 32'h10408000;
      11323: inst = 32'hc404756;
      11324: inst = 32'h8220000;
      11325: inst = 32'h10408000;
      11326: inst = 32'hc404757;
      11327: inst = 32'h8220000;
      11328: inst = 32'h10408000;
      11329: inst = 32'hc404758;
      11330: inst = 32'h8220000;
      11331: inst = 32'h10408000;
      11332: inst = 32'hc404759;
      11333: inst = 32'h8220000;
      11334: inst = 32'h10408000;
      11335: inst = 32'hc40475a;
      11336: inst = 32'h8220000;
      11337: inst = 32'h10408000;
      11338: inst = 32'hc40475b;
      11339: inst = 32'h8220000;
      11340: inst = 32'h10408000;
      11341: inst = 32'hc40475c;
      11342: inst = 32'h8220000;
      11343: inst = 32'h10408000;
      11344: inst = 32'hc40475d;
      11345: inst = 32'h8220000;
      11346: inst = 32'h10408000;
      11347: inst = 32'hc40475e;
      11348: inst = 32'h8220000;
      11349: inst = 32'h10408000;
      11350: inst = 32'hc4047b0;
      11351: inst = 32'h8220000;
      11352: inst = 32'h10408000;
      11353: inst = 32'hc4047b1;
      11354: inst = 32'h8220000;
      11355: inst = 32'h10408000;
      11356: inst = 32'hc4047b2;
      11357: inst = 32'h8220000;
      11358: inst = 32'h10408000;
      11359: inst = 32'hc4047b3;
      11360: inst = 32'h8220000;
      11361: inst = 32'h10408000;
      11362: inst = 32'hc4047b4;
      11363: inst = 32'h8220000;
      11364: inst = 32'h10408000;
      11365: inst = 32'hc4047b5;
      11366: inst = 32'h8220000;
      11367: inst = 32'h10408000;
      11368: inst = 32'hc4047b6;
      11369: inst = 32'h8220000;
      11370: inst = 32'h10408000;
      11371: inst = 32'hc4047b7;
      11372: inst = 32'h8220000;
      11373: inst = 32'h10408000;
      11374: inst = 32'hc4047b8;
      11375: inst = 32'h8220000;
      11376: inst = 32'h10408000;
      11377: inst = 32'hc4047b9;
      11378: inst = 32'h8220000;
      11379: inst = 32'h10408000;
      11380: inst = 32'hc4047ba;
      11381: inst = 32'h8220000;
      11382: inst = 32'h10408000;
      11383: inst = 32'hc4047bb;
      11384: inst = 32'h8220000;
      11385: inst = 32'h10408000;
      11386: inst = 32'hc4047bc;
      11387: inst = 32'h8220000;
      11388: inst = 32'h10408000;
      11389: inst = 32'hc4047bd;
      11390: inst = 32'h8220000;
      11391: inst = 32'h10408000;
      11392: inst = 32'hc4047be;
      11393: inst = 32'h8220000;
      11394: inst = 32'h10408000;
      11395: inst = 32'hc404810;
      11396: inst = 32'h8220000;
      11397: inst = 32'h10408000;
      11398: inst = 32'hc404811;
      11399: inst = 32'h8220000;
      11400: inst = 32'h10408000;
      11401: inst = 32'hc404812;
      11402: inst = 32'h8220000;
      11403: inst = 32'h10408000;
      11404: inst = 32'hc404813;
      11405: inst = 32'h8220000;
      11406: inst = 32'h10408000;
      11407: inst = 32'hc404814;
      11408: inst = 32'h8220000;
      11409: inst = 32'h10408000;
      11410: inst = 32'hc404815;
      11411: inst = 32'h8220000;
      11412: inst = 32'h10408000;
      11413: inst = 32'hc404816;
      11414: inst = 32'h8220000;
      11415: inst = 32'h10408000;
      11416: inst = 32'hc404817;
      11417: inst = 32'h8220000;
      11418: inst = 32'h10408000;
      11419: inst = 32'hc404818;
      11420: inst = 32'h8220000;
      11421: inst = 32'h10408000;
      11422: inst = 32'hc404819;
      11423: inst = 32'h8220000;
      11424: inst = 32'h10408000;
      11425: inst = 32'hc40481a;
      11426: inst = 32'h8220000;
      11427: inst = 32'h10408000;
      11428: inst = 32'hc40481b;
      11429: inst = 32'h8220000;
      11430: inst = 32'h10408000;
      11431: inst = 32'hc40481c;
      11432: inst = 32'h8220000;
      11433: inst = 32'h10408000;
      11434: inst = 32'hc40481d;
      11435: inst = 32'h8220000;
      11436: inst = 32'h10408000;
      11437: inst = 32'hc40481e;
      11438: inst = 32'h8220000;
      11439: inst = 32'h10408000;
      11440: inst = 32'hc404870;
      11441: inst = 32'h8220000;
      11442: inst = 32'h10408000;
      11443: inst = 32'hc404871;
      11444: inst = 32'h8220000;
      11445: inst = 32'h10408000;
      11446: inst = 32'hc404872;
      11447: inst = 32'h8220000;
      11448: inst = 32'h10408000;
      11449: inst = 32'hc404873;
      11450: inst = 32'h8220000;
      11451: inst = 32'h10408000;
      11452: inst = 32'hc404874;
      11453: inst = 32'h8220000;
      11454: inst = 32'h10408000;
      11455: inst = 32'hc404875;
      11456: inst = 32'h8220000;
      11457: inst = 32'h10408000;
      11458: inst = 32'hc404876;
      11459: inst = 32'h8220000;
      11460: inst = 32'h10408000;
      11461: inst = 32'hc404877;
      11462: inst = 32'h8220000;
      11463: inst = 32'h10408000;
      11464: inst = 32'hc404878;
      11465: inst = 32'h8220000;
      11466: inst = 32'h10408000;
      11467: inst = 32'hc404879;
      11468: inst = 32'h8220000;
      11469: inst = 32'h10408000;
      11470: inst = 32'hc40487a;
      11471: inst = 32'h8220000;
      11472: inst = 32'h10408000;
      11473: inst = 32'hc40487b;
      11474: inst = 32'h8220000;
      11475: inst = 32'h10408000;
      11476: inst = 32'hc40487c;
      11477: inst = 32'h8220000;
      11478: inst = 32'h10408000;
      11479: inst = 32'hc40487d;
      11480: inst = 32'h8220000;
      11481: inst = 32'h10408000;
      11482: inst = 32'hc40487e;
      11483: inst = 32'h8220000;
      11484: inst = 32'h10408000;
      11485: inst = 32'hc4048d0;
      11486: inst = 32'h8220000;
      11487: inst = 32'h10408000;
      11488: inst = 32'hc4048d1;
      11489: inst = 32'h8220000;
      11490: inst = 32'h10408000;
      11491: inst = 32'hc4048d2;
      11492: inst = 32'h8220000;
      11493: inst = 32'h10408000;
      11494: inst = 32'hc4048d3;
      11495: inst = 32'h8220000;
      11496: inst = 32'h10408000;
      11497: inst = 32'hc4048d4;
      11498: inst = 32'h8220000;
      11499: inst = 32'h10408000;
      11500: inst = 32'hc4048d5;
      11501: inst = 32'h8220000;
      11502: inst = 32'h10408000;
      11503: inst = 32'hc4048d6;
      11504: inst = 32'h8220000;
      11505: inst = 32'h10408000;
      11506: inst = 32'hc4048d7;
      11507: inst = 32'h8220000;
      11508: inst = 32'h10408000;
      11509: inst = 32'hc4048d8;
      11510: inst = 32'h8220000;
      11511: inst = 32'h10408000;
      11512: inst = 32'hc4048d9;
      11513: inst = 32'h8220000;
      11514: inst = 32'h10408000;
      11515: inst = 32'hc4048da;
      11516: inst = 32'h8220000;
      11517: inst = 32'h10408000;
      11518: inst = 32'hc4048db;
      11519: inst = 32'h8220000;
      11520: inst = 32'h10408000;
      11521: inst = 32'hc4048dc;
      11522: inst = 32'h8220000;
      11523: inst = 32'h10408000;
      11524: inst = 32'hc4048dd;
      11525: inst = 32'h8220000;
      11526: inst = 32'h10408000;
      11527: inst = 32'hc4048de;
      11528: inst = 32'h8220000;
      11529: inst = 32'h10408000;
      11530: inst = 32'hc404930;
      11531: inst = 32'h8220000;
      11532: inst = 32'h10408000;
      11533: inst = 32'hc404931;
      11534: inst = 32'h8220000;
      11535: inst = 32'h10408000;
      11536: inst = 32'hc404936;
      11537: inst = 32'h8220000;
      11538: inst = 32'h10408000;
      11539: inst = 32'hc404937;
      11540: inst = 32'h8220000;
      11541: inst = 32'h10408000;
      11542: inst = 32'hc404938;
      11543: inst = 32'h8220000;
      11544: inst = 32'h10408000;
      11545: inst = 32'hc404939;
      11546: inst = 32'h8220000;
      11547: inst = 32'h10408000;
      11548: inst = 32'hc40493a;
      11549: inst = 32'h8220000;
      11550: inst = 32'h10408000;
      11551: inst = 32'hc40493b;
      11552: inst = 32'h8220000;
      11553: inst = 32'h10408000;
      11554: inst = 32'hc40493c;
      11555: inst = 32'h8220000;
      11556: inst = 32'h10408000;
      11557: inst = 32'hc40493d;
      11558: inst = 32'h8220000;
      11559: inst = 32'h10408000;
      11560: inst = 32'hc40493e;
      11561: inst = 32'h8220000;
      11562: inst = 32'h10408000;
      11563: inst = 32'hc404990;
      11564: inst = 32'h8220000;
      11565: inst = 32'h10408000;
      11566: inst = 32'hc404991;
      11567: inst = 32'h8220000;
      11568: inst = 32'h10408000;
      11569: inst = 32'hc404996;
      11570: inst = 32'h8220000;
      11571: inst = 32'h10408000;
      11572: inst = 32'hc404997;
      11573: inst = 32'h8220000;
      11574: inst = 32'h10408000;
      11575: inst = 32'hc404998;
      11576: inst = 32'h8220000;
      11577: inst = 32'h10408000;
      11578: inst = 32'hc404999;
      11579: inst = 32'h8220000;
      11580: inst = 32'h10408000;
      11581: inst = 32'hc40499a;
      11582: inst = 32'h8220000;
      11583: inst = 32'h10408000;
      11584: inst = 32'hc40499b;
      11585: inst = 32'h8220000;
      11586: inst = 32'h10408000;
      11587: inst = 32'hc40499c;
      11588: inst = 32'h8220000;
      11589: inst = 32'h10408000;
      11590: inst = 32'hc40499d;
      11591: inst = 32'h8220000;
      11592: inst = 32'h10408000;
      11593: inst = 32'hc40499e;
      11594: inst = 32'h8220000;
      11595: inst = 32'h10408000;
      11596: inst = 32'hc4049f0;
      11597: inst = 32'h8220000;
      11598: inst = 32'h10408000;
      11599: inst = 32'hc4049f1;
      11600: inst = 32'h8220000;
      11601: inst = 32'h10408000;
      11602: inst = 32'hc4049f6;
      11603: inst = 32'h8220000;
      11604: inst = 32'h10408000;
      11605: inst = 32'hc4049f7;
      11606: inst = 32'h8220000;
      11607: inst = 32'h10408000;
      11608: inst = 32'hc4049f8;
      11609: inst = 32'h8220000;
      11610: inst = 32'h10408000;
      11611: inst = 32'hc4049f9;
      11612: inst = 32'h8220000;
      11613: inst = 32'h10408000;
      11614: inst = 32'hc4049fa;
      11615: inst = 32'h8220000;
      11616: inst = 32'h10408000;
      11617: inst = 32'hc4049fb;
      11618: inst = 32'h8220000;
      11619: inst = 32'h10408000;
      11620: inst = 32'hc4049fc;
      11621: inst = 32'h8220000;
      11622: inst = 32'h10408000;
      11623: inst = 32'hc4049fd;
      11624: inst = 32'h8220000;
      11625: inst = 32'h10408000;
      11626: inst = 32'hc4049fe;
      11627: inst = 32'h8220000;
      11628: inst = 32'h10408000;
      11629: inst = 32'hc404a50;
      11630: inst = 32'h8220000;
      11631: inst = 32'h10408000;
      11632: inst = 32'hc404a51;
      11633: inst = 32'h8220000;
      11634: inst = 32'h10408000;
      11635: inst = 32'hc404a56;
      11636: inst = 32'h8220000;
      11637: inst = 32'h10408000;
      11638: inst = 32'hc404a57;
      11639: inst = 32'h8220000;
      11640: inst = 32'h10408000;
      11641: inst = 32'hc404a58;
      11642: inst = 32'h8220000;
      11643: inst = 32'h10408000;
      11644: inst = 32'hc404a59;
      11645: inst = 32'h8220000;
      11646: inst = 32'h10408000;
      11647: inst = 32'hc404a5a;
      11648: inst = 32'h8220000;
      11649: inst = 32'h10408000;
      11650: inst = 32'hc404a5b;
      11651: inst = 32'h8220000;
      11652: inst = 32'h10408000;
      11653: inst = 32'hc404a5c;
      11654: inst = 32'h8220000;
      11655: inst = 32'h10408000;
      11656: inst = 32'hc404a5d;
      11657: inst = 32'h8220000;
      11658: inst = 32'h10408000;
      11659: inst = 32'hc404a5e;
      11660: inst = 32'h8220000;
      11661: inst = 32'h10408000;
      11662: inst = 32'hc404ab0;
      11663: inst = 32'h8220000;
      11664: inst = 32'h10408000;
      11665: inst = 32'hc404ab1;
      11666: inst = 32'h8220000;
      11667: inst = 32'h10408000;
      11668: inst = 32'hc404ab6;
      11669: inst = 32'h8220000;
      11670: inst = 32'h10408000;
      11671: inst = 32'hc404ab7;
      11672: inst = 32'h8220000;
      11673: inst = 32'h10408000;
      11674: inst = 32'hc404ab8;
      11675: inst = 32'h8220000;
      11676: inst = 32'h10408000;
      11677: inst = 32'hc404ab9;
      11678: inst = 32'h8220000;
      11679: inst = 32'h10408000;
      11680: inst = 32'hc404aba;
      11681: inst = 32'h8220000;
      11682: inst = 32'h10408000;
      11683: inst = 32'hc404abb;
      11684: inst = 32'h8220000;
      11685: inst = 32'h10408000;
      11686: inst = 32'hc404abc;
      11687: inst = 32'h8220000;
      11688: inst = 32'h10408000;
      11689: inst = 32'hc404abd;
      11690: inst = 32'h8220000;
      11691: inst = 32'h10408000;
      11692: inst = 32'hc404abe;
      11693: inst = 32'h8220000;
      11694: inst = 32'h10408000;
      11695: inst = 32'hc404b10;
      11696: inst = 32'h8220000;
      11697: inst = 32'h10408000;
      11698: inst = 32'hc404b11;
      11699: inst = 32'h8220000;
      11700: inst = 32'h10408000;
      11701: inst = 32'hc404b16;
      11702: inst = 32'h8220000;
      11703: inst = 32'h10408000;
      11704: inst = 32'hc404b17;
      11705: inst = 32'h8220000;
      11706: inst = 32'h10408000;
      11707: inst = 32'hc404b18;
      11708: inst = 32'h8220000;
      11709: inst = 32'h10408000;
      11710: inst = 32'hc404b19;
      11711: inst = 32'h8220000;
      11712: inst = 32'h10408000;
      11713: inst = 32'hc404b1a;
      11714: inst = 32'h8220000;
      11715: inst = 32'h10408000;
      11716: inst = 32'hc404b1b;
      11717: inst = 32'h8220000;
      11718: inst = 32'h10408000;
      11719: inst = 32'hc404b1c;
      11720: inst = 32'h8220000;
      11721: inst = 32'h10408000;
      11722: inst = 32'hc404b1d;
      11723: inst = 32'h8220000;
      11724: inst = 32'h10408000;
      11725: inst = 32'hc404b1e;
      11726: inst = 32'h8220000;
      11727: inst = 32'h10408000;
      11728: inst = 32'hc404b70;
      11729: inst = 32'h8220000;
      11730: inst = 32'h10408000;
      11731: inst = 32'hc404b71;
      11732: inst = 32'h8220000;
      11733: inst = 32'h10408000;
      11734: inst = 32'hc404b76;
      11735: inst = 32'h8220000;
      11736: inst = 32'h10408000;
      11737: inst = 32'hc404b77;
      11738: inst = 32'h8220000;
      11739: inst = 32'h10408000;
      11740: inst = 32'hc404b78;
      11741: inst = 32'h8220000;
      11742: inst = 32'h10408000;
      11743: inst = 32'hc404b79;
      11744: inst = 32'h8220000;
      11745: inst = 32'h10408000;
      11746: inst = 32'hc404b7a;
      11747: inst = 32'h8220000;
      11748: inst = 32'h10408000;
      11749: inst = 32'hc404b7b;
      11750: inst = 32'h8220000;
      11751: inst = 32'h10408000;
      11752: inst = 32'hc404b7c;
      11753: inst = 32'h8220000;
      11754: inst = 32'h10408000;
      11755: inst = 32'hc404b7d;
      11756: inst = 32'h8220000;
      11757: inst = 32'h10408000;
      11758: inst = 32'hc404b7e;
      11759: inst = 32'h8220000;
      11760: inst = 32'h10408000;
      11761: inst = 32'hc404bd0;
      11762: inst = 32'h8220000;
      11763: inst = 32'h10408000;
      11764: inst = 32'hc404bd1;
      11765: inst = 32'h8220000;
      11766: inst = 32'h10408000;
      11767: inst = 32'hc404bd2;
      11768: inst = 32'h8220000;
      11769: inst = 32'h10408000;
      11770: inst = 32'hc404bd3;
      11771: inst = 32'h8220000;
      11772: inst = 32'h10408000;
      11773: inst = 32'hc404bd4;
      11774: inst = 32'h8220000;
      11775: inst = 32'h10408000;
      11776: inst = 32'hc404bd5;
      11777: inst = 32'h8220000;
      11778: inst = 32'h10408000;
      11779: inst = 32'hc404bd6;
      11780: inst = 32'h8220000;
      11781: inst = 32'h10408000;
      11782: inst = 32'hc404bd7;
      11783: inst = 32'h8220000;
      11784: inst = 32'h10408000;
      11785: inst = 32'hc404bd8;
      11786: inst = 32'h8220000;
      11787: inst = 32'h10408000;
      11788: inst = 32'hc404bd9;
      11789: inst = 32'h8220000;
      11790: inst = 32'h10408000;
      11791: inst = 32'hc404bda;
      11792: inst = 32'h8220000;
      11793: inst = 32'h10408000;
      11794: inst = 32'hc404bdb;
      11795: inst = 32'h8220000;
      11796: inst = 32'h10408000;
      11797: inst = 32'hc404bdc;
      11798: inst = 32'h8220000;
      11799: inst = 32'h10408000;
      11800: inst = 32'hc404bdd;
      11801: inst = 32'h8220000;
      11802: inst = 32'h10408000;
      11803: inst = 32'hc404bde;
      11804: inst = 32'h8220000;
      11805: inst = 32'h10408000;
      11806: inst = 32'hc404c30;
      11807: inst = 32'h8220000;
      11808: inst = 32'h10408000;
      11809: inst = 32'hc404c31;
      11810: inst = 32'h8220000;
      11811: inst = 32'h10408000;
      11812: inst = 32'hc404c32;
      11813: inst = 32'h8220000;
      11814: inst = 32'h10408000;
      11815: inst = 32'hc404c33;
      11816: inst = 32'h8220000;
      11817: inst = 32'h10408000;
      11818: inst = 32'hc404c34;
      11819: inst = 32'h8220000;
      11820: inst = 32'h10408000;
      11821: inst = 32'hc404c35;
      11822: inst = 32'h8220000;
      11823: inst = 32'h10408000;
      11824: inst = 32'hc404c36;
      11825: inst = 32'h8220000;
      11826: inst = 32'h10408000;
      11827: inst = 32'hc404c37;
      11828: inst = 32'h8220000;
      11829: inst = 32'h10408000;
      11830: inst = 32'hc404c38;
      11831: inst = 32'h8220000;
      11832: inst = 32'h10408000;
      11833: inst = 32'hc404c39;
      11834: inst = 32'h8220000;
      11835: inst = 32'h10408000;
      11836: inst = 32'hc404c3a;
      11837: inst = 32'h8220000;
      11838: inst = 32'h10408000;
      11839: inst = 32'hc404c3b;
      11840: inst = 32'h8220000;
      11841: inst = 32'h10408000;
      11842: inst = 32'hc404c3c;
      11843: inst = 32'h8220000;
      11844: inst = 32'h10408000;
      11845: inst = 32'hc404c3d;
      11846: inst = 32'h8220000;
      11847: inst = 32'h10408000;
      11848: inst = 32'hc404c3e;
      11849: inst = 32'h8220000;
      11850: inst = 32'h10408000;
      11851: inst = 32'hc404c90;
      11852: inst = 32'h8220000;
      11853: inst = 32'h10408000;
      11854: inst = 32'hc404c91;
      11855: inst = 32'h8220000;
      11856: inst = 32'h10408000;
      11857: inst = 32'hc404c92;
      11858: inst = 32'h8220000;
      11859: inst = 32'h10408000;
      11860: inst = 32'hc404c93;
      11861: inst = 32'h8220000;
      11862: inst = 32'h10408000;
      11863: inst = 32'hc404c94;
      11864: inst = 32'h8220000;
      11865: inst = 32'h10408000;
      11866: inst = 32'hc404c95;
      11867: inst = 32'h8220000;
      11868: inst = 32'h10408000;
      11869: inst = 32'hc404c96;
      11870: inst = 32'h8220000;
      11871: inst = 32'h10408000;
      11872: inst = 32'hc404c97;
      11873: inst = 32'h8220000;
      11874: inst = 32'h10408000;
      11875: inst = 32'hc404c98;
      11876: inst = 32'h8220000;
      11877: inst = 32'h10408000;
      11878: inst = 32'hc404c99;
      11879: inst = 32'h8220000;
      11880: inst = 32'h10408000;
      11881: inst = 32'hc404c9a;
      11882: inst = 32'h8220000;
      11883: inst = 32'h10408000;
      11884: inst = 32'hc404c9b;
      11885: inst = 32'h8220000;
      11886: inst = 32'h10408000;
      11887: inst = 32'hc404c9c;
      11888: inst = 32'h8220000;
      11889: inst = 32'h10408000;
      11890: inst = 32'hc404c9d;
      11891: inst = 32'h8220000;
      11892: inst = 32'h10408000;
      11893: inst = 32'hc404c9e;
      11894: inst = 32'h8220000;
      11895: inst = 32'h10408000;
      11896: inst = 32'hc404cf0;
      11897: inst = 32'h8220000;
      11898: inst = 32'h10408000;
      11899: inst = 32'hc404cf1;
      11900: inst = 32'h8220000;
      11901: inst = 32'h10408000;
      11902: inst = 32'hc404cf2;
      11903: inst = 32'h8220000;
      11904: inst = 32'h10408000;
      11905: inst = 32'hc404cf3;
      11906: inst = 32'h8220000;
      11907: inst = 32'h10408000;
      11908: inst = 32'hc404cf4;
      11909: inst = 32'h8220000;
      11910: inst = 32'h10408000;
      11911: inst = 32'hc404cf5;
      11912: inst = 32'h8220000;
      11913: inst = 32'h10408000;
      11914: inst = 32'hc404cf6;
      11915: inst = 32'h8220000;
      11916: inst = 32'h10408000;
      11917: inst = 32'hc404cf7;
      11918: inst = 32'h8220000;
      11919: inst = 32'h10408000;
      11920: inst = 32'hc404cf8;
      11921: inst = 32'h8220000;
      11922: inst = 32'h10408000;
      11923: inst = 32'hc404cf9;
      11924: inst = 32'h8220000;
      11925: inst = 32'h10408000;
      11926: inst = 32'hc404cfa;
      11927: inst = 32'h8220000;
      11928: inst = 32'h10408000;
      11929: inst = 32'hc404cfe;
      11930: inst = 32'h8220000;
      11931: inst = 32'h10408000;
      11932: inst = 32'hc404d50;
      11933: inst = 32'h8220000;
      11934: inst = 32'h10408000;
      11935: inst = 32'hc404d51;
      11936: inst = 32'h8220000;
      11937: inst = 32'h10408000;
      11938: inst = 32'hc404d52;
      11939: inst = 32'h8220000;
      11940: inst = 32'h10408000;
      11941: inst = 32'hc404d53;
      11942: inst = 32'h8220000;
      11943: inst = 32'h10408000;
      11944: inst = 32'hc404d54;
      11945: inst = 32'h8220000;
      11946: inst = 32'h10408000;
      11947: inst = 32'hc404d55;
      11948: inst = 32'h8220000;
      11949: inst = 32'h10408000;
      11950: inst = 32'hc404d56;
      11951: inst = 32'h8220000;
      11952: inst = 32'h10408000;
      11953: inst = 32'hc404d57;
      11954: inst = 32'h8220000;
      11955: inst = 32'h10408000;
      11956: inst = 32'hc404d58;
      11957: inst = 32'h8220000;
      11958: inst = 32'h10408000;
      11959: inst = 32'hc404d59;
      11960: inst = 32'h8220000;
      11961: inst = 32'h10408000;
      11962: inst = 32'hc404d5a;
      11963: inst = 32'h8220000;
      11964: inst = 32'h10408000;
      11965: inst = 32'hc404d5c;
      11966: inst = 32'h8220000;
      11967: inst = 32'h10408000;
      11968: inst = 32'hc404d5d;
      11969: inst = 32'h8220000;
      11970: inst = 32'h10408000;
      11971: inst = 32'hc404d5e;
      11972: inst = 32'h8220000;
      11973: inst = 32'h10408000;
      11974: inst = 32'hc404db0;
      11975: inst = 32'h8220000;
      11976: inst = 32'h10408000;
      11977: inst = 32'hc404db1;
      11978: inst = 32'h8220000;
      11979: inst = 32'h10408000;
      11980: inst = 32'hc404db2;
      11981: inst = 32'h8220000;
      11982: inst = 32'h10408000;
      11983: inst = 32'hc404db3;
      11984: inst = 32'h8220000;
      11985: inst = 32'h10408000;
      11986: inst = 32'hc404db4;
      11987: inst = 32'h8220000;
      11988: inst = 32'h10408000;
      11989: inst = 32'hc404db5;
      11990: inst = 32'h8220000;
      11991: inst = 32'h10408000;
      11992: inst = 32'hc404db6;
      11993: inst = 32'h8220000;
      11994: inst = 32'h10408000;
      11995: inst = 32'hc404db7;
      11996: inst = 32'h8220000;
      11997: inst = 32'h10408000;
      11998: inst = 32'hc404db8;
      11999: inst = 32'h8220000;
      12000: inst = 32'h10408000;
      12001: inst = 32'hc404db9;
      12002: inst = 32'h8220000;
      12003: inst = 32'h10408000;
      12004: inst = 32'hc404dba;
      12005: inst = 32'h8220000;
      12006: inst = 32'h10408000;
      12007: inst = 32'hc404dbb;
      12008: inst = 32'h8220000;
      12009: inst = 32'h10408000;
      12010: inst = 32'hc404dbc;
      12011: inst = 32'h8220000;
      12012: inst = 32'h10408000;
      12013: inst = 32'hc404dbd;
      12014: inst = 32'h8220000;
      12015: inst = 32'h10408000;
      12016: inst = 32'hc404dbe;
      12017: inst = 32'h8220000;
      12018: inst = 32'h10408000;
      12019: inst = 32'hc404e10;
      12020: inst = 32'h8220000;
      12021: inst = 32'h10408000;
      12022: inst = 32'hc404e11;
      12023: inst = 32'h8220000;
      12024: inst = 32'h10408000;
      12025: inst = 32'hc404e12;
      12026: inst = 32'h8220000;
      12027: inst = 32'h10408000;
      12028: inst = 32'hc404e13;
      12029: inst = 32'h8220000;
      12030: inst = 32'h10408000;
      12031: inst = 32'hc404e14;
      12032: inst = 32'h8220000;
      12033: inst = 32'h10408000;
      12034: inst = 32'hc404e15;
      12035: inst = 32'h8220000;
      12036: inst = 32'h10408000;
      12037: inst = 32'hc404e16;
      12038: inst = 32'h8220000;
      12039: inst = 32'h10408000;
      12040: inst = 32'hc404e17;
      12041: inst = 32'h8220000;
      12042: inst = 32'h10408000;
      12043: inst = 32'hc404e18;
      12044: inst = 32'h8220000;
      12045: inst = 32'h10408000;
      12046: inst = 32'hc404e19;
      12047: inst = 32'h8220000;
      12048: inst = 32'h10408000;
      12049: inst = 32'hc404e1a;
      12050: inst = 32'h8220000;
      12051: inst = 32'h10408000;
      12052: inst = 32'hc404e1b;
      12053: inst = 32'h8220000;
      12054: inst = 32'h10408000;
      12055: inst = 32'hc404e1c;
      12056: inst = 32'h8220000;
      12057: inst = 32'h10408000;
      12058: inst = 32'hc404e1d;
      12059: inst = 32'h8220000;
      12060: inst = 32'h10408000;
      12061: inst = 32'hc404e1e;
      12062: inst = 32'h8220000;
      12063: inst = 32'h10408000;
      12064: inst = 32'hc404e70;
      12065: inst = 32'h8220000;
      12066: inst = 32'h10408000;
      12067: inst = 32'hc404e71;
      12068: inst = 32'h8220000;
      12069: inst = 32'h10408000;
      12070: inst = 32'hc404e72;
      12071: inst = 32'h8220000;
      12072: inst = 32'h10408000;
      12073: inst = 32'hc404e73;
      12074: inst = 32'h8220000;
      12075: inst = 32'h10408000;
      12076: inst = 32'hc404e74;
      12077: inst = 32'h8220000;
      12078: inst = 32'h10408000;
      12079: inst = 32'hc404e75;
      12080: inst = 32'h8220000;
      12081: inst = 32'h10408000;
      12082: inst = 32'hc404e76;
      12083: inst = 32'h8220000;
      12084: inst = 32'h10408000;
      12085: inst = 32'hc404e77;
      12086: inst = 32'h8220000;
      12087: inst = 32'h10408000;
      12088: inst = 32'hc404e78;
      12089: inst = 32'h8220000;
      12090: inst = 32'h10408000;
      12091: inst = 32'hc404e79;
      12092: inst = 32'h8220000;
      12093: inst = 32'h10408000;
      12094: inst = 32'hc404e7a;
      12095: inst = 32'h8220000;
      12096: inst = 32'h10408000;
      12097: inst = 32'hc404e7b;
      12098: inst = 32'h8220000;
      12099: inst = 32'h10408000;
      12100: inst = 32'hc404e7c;
      12101: inst = 32'h8220000;
      12102: inst = 32'h10408000;
      12103: inst = 32'hc404e7d;
      12104: inst = 32'h8220000;
      12105: inst = 32'h10408000;
      12106: inst = 32'hc404e7e;
      12107: inst = 32'h8220000;
      12108: inst = 32'h10408000;
      12109: inst = 32'hc404ed0;
      12110: inst = 32'h8220000;
      12111: inst = 32'h10408000;
      12112: inst = 32'hc404ed1;
      12113: inst = 32'h8220000;
      12114: inst = 32'h10408000;
      12115: inst = 32'hc404ed2;
      12116: inst = 32'h8220000;
      12117: inst = 32'h10408000;
      12118: inst = 32'hc404ed3;
      12119: inst = 32'h8220000;
      12120: inst = 32'h10408000;
      12121: inst = 32'hc404ed4;
      12122: inst = 32'h8220000;
      12123: inst = 32'h10408000;
      12124: inst = 32'hc404ed5;
      12125: inst = 32'h8220000;
      12126: inst = 32'h10408000;
      12127: inst = 32'hc404ed6;
      12128: inst = 32'h8220000;
      12129: inst = 32'h10408000;
      12130: inst = 32'hc404ed7;
      12131: inst = 32'h8220000;
      12132: inst = 32'h10408000;
      12133: inst = 32'hc404ed8;
      12134: inst = 32'h8220000;
      12135: inst = 32'h10408000;
      12136: inst = 32'hc404ed9;
      12137: inst = 32'h8220000;
      12138: inst = 32'h10408000;
      12139: inst = 32'hc404eda;
      12140: inst = 32'h8220000;
      12141: inst = 32'h10408000;
      12142: inst = 32'hc404edb;
      12143: inst = 32'h8220000;
      12144: inst = 32'h10408000;
      12145: inst = 32'hc404edc;
      12146: inst = 32'h8220000;
      12147: inst = 32'h10408000;
      12148: inst = 32'hc404edd;
      12149: inst = 32'h8220000;
      12150: inst = 32'h10408000;
      12151: inst = 32'hc404ede;
      12152: inst = 32'h8220000;
      12153: inst = 32'h10408000;
      12154: inst = 32'hc404f30;
      12155: inst = 32'h8220000;
      12156: inst = 32'h10408000;
      12157: inst = 32'hc404f31;
      12158: inst = 32'h8220000;
      12159: inst = 32'h10408000;
      12160: inst = 32'hc404f32;
      12161: inst = 32'h8220000;
      12162: inst = 32'h10408000;
      12163: inst = 32'hc404f33;
      12164: inst = 32'h8220000;
      12165: inst = 32'h10408000;
      12166: inst = 32'hc404f34;
      12167: inst = 32'h8220000;
      12168: inst = 32'h10408000;
      12169: inst = 32'hc404f35;
      12170: inst = 32'h8220000;
      12171: inst = 32'h10408000;
      12172: inst = 32'hc404f36;
      12173: inst = 32'h8220000;
      12174: inst = 32'h10408000;
      12175: inst = 32'hc404f37;
      12176: inst = 32'h8220000;
      12177: inst = 32'h10408000;
      12178: inst = 32'hc404f38;
      12179: inst = 32'h8220000;
      12180: inst = 32'h10408000;
      12181: inst = 32'hc404f39;
      12182: inst = 32'h8220000;
      12183: inst = 32'h10408000;
      12184: inst = 32'hc404f3a;
      12185: inst = 32'h8220000;
      12186: inst = 32'h10408000;
      12187: inst = 32'hc404f3b;
      12188: inst = 32'h8220000;
      12189: inst = 32'h10408000;
      12190: inst = 32'hc404f3c;
      12191: inst = 32'h8220000;
      12192: inst = 32'h10408000;
      12193: inst = 32'hc404f3d;
      12194: inst = 32'h8220000;
      12195: inst = 32'h10408000;
      12196: inst = 32'hc404f3e;
      12197: inst = 32'h8220000;
      12198: inst = 32'h10408000;
      12199: inst = 32'hc404f90;
      12200: inst = 32'h8220000;
      12201: inst = 32'h10408000;
      12202: inst = 32'hc404f91;
      12203: inst = 32'h8220000;
      12204: inst = 32'h10408000;
      12205: inst = 32'hc404f92;
      12206: inst = 32'h8220000;
      12207: inst = 32'h10408000;
      12208: inst = 32'hc404f93;
      12209: inst = 32'h8220000;
      12210: inst = 32'h10408000;
      12211: inst = 32'hc404f94;
      12212: inst = 32'h8220000;
      12213: inst = 32'h10408000;
      12214: inst = 32'hc404f95;
      12215: inst = 32'h8220000;
      12216: inst = 32'h10408000;
      12217: inst = 32'hc404f96;
      12218: inst = 32'h8220000;
      12219: inst = 32'h10408000;
      12220: inst = 32'hc404f97;
      12221: inst = 32'h8220000;
      12222: inst = 32'h10408000;
      12223: inst = 32'hc404f98;
      12224: inst = 32'h8220000;
      12225: inst = 32'h10408000;
      12226: inst = 32'hc404f99;
      12227: inst = 32'h8220000;
      12228: inst = 32'h10408000;
      12229: inst = 32'hc404f9a;
      12230: inst = 32'h8220000;
      12231: inst = 32'h10408000;
      12232: inst = 32'hc404f9b;
      12233: inst = 32'h8220000;
      12234: inst = 32'h10408000;
      12235: inst = 32'hc404f9c;
      12236: inst = 32'h8220000;
      12237: inst = 32'h10408000;
      12238: inst = 32'hc404f9d;
      12239: inst = 32'h8220000;
      12240: inst = 32'h10408000;
      12241: inst = 32'hc404f9e;
      12242: inst = 32'h8220000;
      12243: inst = 32'h10408000;
      12244: inst = 32'hc404ff0;
      12245: inst = 32'h8220000;
      12246: inst = 32'h10408000;
      12247: inst = 32'hc404ff1;
      12248: inst = 32'h8220000;
      12249: inst = 32'h10408000;
      12250: inst = 32'hc404ff2;
      12251: inst = 32'h8220000;
      12252: inst = 32'h10408000;
      12253: inst = 32'hc404ff3;
      12254: inst = 32'h8220000;
      12255: inst = 32'h10408000;
      12256: inst = 32'hc404ff4;
      12257: inst = 32'h8220000;
      12258: inst = 32'h10408000;
      12259: inst = 32'hc404ff5;
      12260: inst = 32'h8220000;
      12261: inst = 32'h10408000;
      12262: inst = 32'hc404ff6;
      12263: inst = 32'h8220000;
      12264: inst = 32'h10408000;
      12265: inst = 32'hc404ff7;
      12266: inst = 32'h8220000;
      12267: inst = 32'h10408000;
      12268: inst = 32'hc404ff8;
      12269: inst = 32'h8220000;
      12270: inst = 32'h10408000;
      12271: inst = 32'hc404ff9;
      12272: inst = 32'h8220000;
      12273: inst = 32'h10408000;
      12274: inst = 32'hc404ffa;
      12275: inst = 32'h8220000;
      12276: inst = 32'h10408000;
      12277: inst = 32'hc404ffb;
      12278: inst = 32'h8220000;
      12279: inst = 32'h10408000;
      12280: inst = 32'hc404ffc;
      12281: inst = 32'h8220000;
      12282: inst = 32'h10408000;
      12283: inst = 32'hc404ffd;
      12284: inst = 32'h8220000;
      12285: inst = 32'h10408000;
      12286: inst = 32'hc404ffe;
      12287: inst = 32'h8220000;
      12288: inst = 32'h10408000;
      12289: inst = 32'hc405050;
      12290: inst = 32'h8220000;
      12291: inst = 32'h10408000;
      12292: inst = 32'hc405051;
      12293: inst = 32'h8220000;
      12294: inst = 32'h10408000;
      12295: inst = 32'hc405052;
      12296: inst = 32'h8220000;
      12297: inst = 32'h10408000;
      12298: inst = 32'hc405053;
      12299: inst = 32'h8220000;
      12300: inst = 32'h10408000;
      12301: inst = 32'hc405054;
      12302: inst = 32'h8220000;
      12303: inst = 32'h10408000;
      12304: inst = 32'hc405055;
      12305: inst = 32'h8220000;
      12306: inst = 32'h10408000;
      12307: inst = 32'hc405056;
      12308: inst = 32'h8220000;
      12309: inst = 32'h10408000;
      12310: inst = 32'hc405057;
      12311: inst = 32'h8220000;
      12312: inst = 32'h10408000;
      12313: inst = 32'hc405058;
      12314: inst = 32'h8220000;
      12315: inst = 32'h10408000;
      12316: inst = 32'hc405059;
      12317: inst = 32'h8220000;
      12318: inst = 32'h10408000;
      12319: inst = 32'hc40505a;
      12320: inst = 32'h8220000;
      12321: inst = 32'h10408000;
      12322: inst = 32'hc40505b;
      12323: inst = 32'h8220000;
      12324: inst = 32'h10408000;
      12325: inst = 32'hc40505c;
      12326: inst = 32'h8220000;
      12327: inst = 32'h10408000;
      12328: inst = 32'hc40505d;
      12329: inst = 32'h8220000;
      12330: inst = 32'h10408000;
      12331: inst = 32'hc40505e;
      12332: inst = 32'h8220000;
      12333: inst = 32'h10408000;
      12334: inst = 32'hc4050b0;
      12335: inst = 32'h8220000;
      12336: inst = 32'h10408000;
      12337: inst = 32'hc4050b1;
      12338: inst = 32'h8220000;
      12339: inst = 32'h10408000;
      12340: inst = 32'hc4050b2;
      12341: inst = 32'h8220000;
      12342: inst = 32'h10408000;
      12343: inst = 32'hc4050b3;
      12344: inst = 32'h8220000;
      12345: inst = 32'h10408000;
      12346: inst = 32'hc4050b4;
      12347: inst = 32'h8220000;
      12348: inst = 32'h10408000;
      12349: inst = 32'hc4050b5;
      12350: inst = 32'h8220000;
      12351: inst = 32'h10408000;
      12352: inst = 32'hc4050b6;
      12353: inst = 32'h8220000;
      12354: inst = 32'h10408000;
      12355: inst = 32'hc4050b7;
      12356: inst = 32'h8220000;
      12357: inst = 32'h10408000;
      12358: inst = 32'hc4050b8;
      12359: inst = 32'h8220000;
      12360: inst = 32'h10408000;
      12361: inst = 32'hc4050b9;
      12362: inst = 32'h8220000;
      12363: inst = 32'h10408000;
      12364: inst = 32'hc4050ba;
      12365: inst = 32'h8220000;
      12366: inst = 32'h10408000;
      12367: inst = 32'hc4050bb;
      12368: inst = 32'h8220000;
      12369: inst = 32'h10408000;
      12370: inst = 32'hc4050bc;
      12371: inst = 32'h8220000;
      12372: inst = 32'h10408000;
      12373: inst = 32'hc4050bd;
      12374: inst = 32'h8220000;
      12375: inst = 32'h10408000;
      12376: inst = 32'hc4050be;
      12377: inst = 32'h8220000;
      12378: inst = 32'h10408000;
      12379: inst = 32'hc405110;
      12380: inst = 32'h8220000;
      12381: inst = 32'h10408000;
      12382: inst = 32'hc405111;
      12383: inst = 32'h8220000;
      12384: inst = 32'h10408000;
      12385: inst = 32'hc405112;
      12386: inst = 32'h8220000;
      12387: inst = 32'h10408000;
      12388: inst = 32'hc405113;
      12389: inst = 32'h8220000;
      12390: inst = 32'h10408000;
      12391: inst = 32'hc405114;
      12392: inst = 32'h8220000;
      12393: inst = 32'h10408000;
      12394: inst = 32'hc405115;
      12395: inst = 32'h8220000;
      12396: inst = 32'h10408000;
      12397: inst = 32'hc405116;
      12398: inst = 32'h8220000;
      12399: inst = 32'h10408000;
      12400: inst = 32'hc405117;
      12401: inst = 32'h8220000;
      12402: inst = 32'h10408000;
      12403: inst = 32'hc405118;
      12404: inst = 32'h8220000;
      12405: inst = 32'h10408000;
      12406: inst = 32'hc405119;
      12407: inst = 32'h8220000;
      12408: inst = 32'h10408000;
      12409: inst = 32'hc40511a;
      12410: inst = 32'h8220000;
      12411: inst = 32'h10408000;
      12412: inst = 32'hc40511b;
      12413: inst = 32'h8220000;
      12414: inst = 32'h10408000;
      12415: inst = 32'hc40511c;
      12416: inst = 32'h8220000;
      12417: inst = 32'h10408000;
      12418: inst = 32'hc40511d;
      12419: inst = 32'h8220000;
      12420: inst = 32'h10408000;
      12421: inst = 32'hc40511e;
      12422: inst = 32'h8220000;
      12423: inst = 32'h10408000;
      12424: inst = 32'hc405170;
      12425: inst = 32'h8220000;
      12426: inst = 32'h10408000;
      12427: inst = 32'hc405171;
      12428: inst = 32'h8220000;
      12429: inst = 32'h10408000;
      12430: inst = 32'hc405172;
      12431: inst = 32'h8220000;
      12432: inst = 32'h10408000;
      12433: inst = 32'hc405173;
      12434: inst = 32'h8220000;
      12435: inst = 32'h10408000;
      12436: inst = 32'hc405174;
      12437: inst = 32'h8220000;
      12438: inst = 32'h10408000;
      12439: inst = 32'hc405175;
      12440: inst = 32'h8220000;
      12441: inst = 32'h10408000;
      12442: inst = 32'hc405176;
      12443: inst = 32'h8220000;
      12444: inst = 32'h10408000;
      12445: inst = 32'hc405177;
      12446: inst = 32'h8220000;
      12447: inst = 32'h10408000;
      12448: inst = 32'hc405178;
      12449: inst = 32'h8220000;
      12450: inst = 32'h10408000;
      12451: inst = 32'hc405179;
      12452: inst = 32'h8220000;
      12453: inst = 32'h10408000;
      12454: inst = 32'hc40517a;
      12455: inst = 32'h8220000;
      12456: inst = 32'h10408000;
      12457: inst = 32'hc40517b;
      12458: inst = 32'h8220000;
      12459: inst = 32'h10408000;
      12460: inst = 32'hc40517c;
      12461: inst = 32'h8220000;
      12462: inst = 32'h10408000;
      12463: inst = 32'hc40517d;
      12464: inst = 32'h8220000;
      12465: inst = 32'h10408000;
      12466: inst = 32'hc40517e;
      12467: inst = 32'h8220000;
      12468: inst = 32'h10408000;
      12469: inst = 32'hc4051d0;
      12470: inst = 32'h8220000;
      12471: inst = 32'h10408000;
      12472: inst = 32'hc4051d1;
      12473: inst = 32'h8220000;
      12474: inst = 32'h10408000;
      12475: inst = 32'hc4051d2;
      12476: inst = 32'h8220000;
      12477: inst = 32'h10408000;
      12478: inst = 32'hc4051d3;
      12479: inst = 32'h8220000;
      12480: inst = 32'h10408000;
      12481: inst = 32'hc4051d4;
      12482: inst = 32'h8220000;
      12483: inst = 32'h10408000;
      12484: inst = 32'hc4051d5;
      12485: inst = 32'h8220000;
      12486: inst = 32'h10408000;
      12487: inst = 32'hc4051d6;
      12488: inst = 32'h8220000;
      12489: inst = 32'h10408000;
      12490: inst = 32'hc4051d7;
      12491: inst = 32'h8220000;
      12492: inst = 32'h10408000;
      12493: inst = 32'hc4051d8;
      12494: inst = 32'h8220000;
      12495: inst = 32'h10408000;
      12496: inst = 32'hc4051d9;
      12497: inst = 32'h8220000;
      12498: inst = 32'h10408000;
      12499: inst = 32'hc4051da;
      12500: inst = 32'h8220000;
      12501: inst = 32'h10408000;
      12502: inst = 32'hc4051db;
      12503: inst = 32'h8220000;
      12504: inst = 32'h10408000;
      12505: inst = 32'hc4051dc;
      12506: inst = 32'h8220000;
      12507: inst = 32'h10408000;
      12508: inst = 32'hc4051dd;
      12509: inst = 32'h8220000;
      12510: inst = 32'h10408000;
      12511: inst = 32'hc4051de;
      12512: inst = 32'h8220000;
      12513: inst = 32'h10408000;
      12514: inst = 32'hc405230;
      12515: inst = 32'h8220000;
      12516: inst = 32'h10408000;
      12517: inst = 32'hc405231;
      12518: inst = 32'h8220000;
      12519: inst = 32'h10408000;
      12520: inst = 32'hc405232;
      12521: inst = 32'h8220000;
      12522: inst = 32'h10408000;
      12523: inst = 32'hc405233;
      12524: inst = 32'h8220000;
      12525: inst = 32'h10408000;
      12526: inst = 32'hc405234;
      12527: inst = 32'h8220000;
      12528: inst = 32'h10408000;
      12529: inst = 32'hc405235;
      12530: inst = 32'h8220000;
      12531: inst = 32'h10408000;
      12532: inst = 32'hc405236;
      12533: inst = 32'h8220000;
      12534: inst = 32'h10408000;
      12535: inst = 32'hc405237;
      12536: inst = 32'h8220000;
      12537: inst = 32'h10408000;
      12538: inst = 32'hc405238;
      12539: inst = 32'h8220000;
      12540: inst = 32'h10408000;
      12541: inst = 32'hc405239;
      12542: inst = 32'h8220000;
      12543: inst = 32'h10408000;
      12544: inst = 32'hc40523a;
      12545: inst = 32'h8220000;
      12546: inst = 32'h10408000;
      12547: inst = 32'hc40523b;
      12548: inst = 32'h8220000;
      12549: inst = 32'h10408000;
      12550: inst = 32'hc40523c;
      12551: inst = 32'h8220000;
      12552: inst = 32'h10408000;
      12553: inst = 32'hc40523d;
      12554: inst = 32'h8220000;
      12555: inst = 32'h10408000;
      12556: inst = 32'hc40523e;
      12557: inst = 32'h8220000;
      12558: inst = 32'h10408000;
      12559: inst = 32'hc405290;
      12560: inst = 32'h8220000;
      12561: inst = 32'h10408000;
      12562: inst = 32'hc405291;
      12563: inst = 32'h8220000;
      12564: inst = 32'h10408000;
      12565: inst = 32'hc405292;
      12566: inst = 32'h8220000;
      12567: inst = 32'h10408000;
      12568: inst = 32'hc405293;
      12569: inst = 32'h8220000;
      12570: inst = 32'h10408000;
      12571: inst = 32'hc405294;
      12572: inst = 32'h8220000;
      12573: inst = 32'h10408000;
      12574: inst = 32'hc405295;
      12575: inst = 32'h8220000;
      12576: inst = 32'h10408000;
      12577: inst = 32'hc405296;
      12578: inst = 32'h8220000;
      12579: inst = 32'h10408000;
      12580: inst = 32'hc405297;
      12581: inst = 32'h8220000;
      12582: inst = 32'h10408000;
      12583: inst = 32'hc405298;
      12584: inst = 32'h8220000;
      12585: inst = 32'h10408000;
      12586: inst = 32'hc405299;
      12587: inst = 32'h8220000;
      12588: inst = 32'h10408000;
      12589: inst = 32'hc40529a;
      12590: inst = 32'h8220000;
      12591: inst = 32'h10408000;
      12592: inst = 32'hc40529b;
      12593: inst = 32'h8220000;
      12594: inst = 32'h10408000;
      12595: inst = 32'hc40529c;
      12596: inst = 32'h8220000;
      12597: inst = 32'h10408000;
      12598: inst = 32'hc40529d;
      12599: inst = 32'h8220000;
      12600: inst = 32'h10408000;
      12601: inst = 32'hc40529e;
      12602: inst = 32'h8220000;
      12603: inst = 32'hc20ef7c;
      12604: inst = 32'h10408000;
      12605: inst = 32'hc404932;
      12606: inst = 32'h8220000;
      12607: inst = 32'h10408000;
      12608: inst = 32'hc404933;
      12609: inst = 32'h8220000;
      12610: inst = 32'h10408000;
      12611: inst = 32'hc404934;
      12612: inst = 32'h8220000;
      12613: inst = 32'h10408000;
      12614: inst = 32'hc404935;
      12615: inst = 32'h8220000;
      12616: inst = 32'h10408000;
      12617: inst = 32'hc404993;
      12618: inst = 32'h8220000;
      12619: inst = 32'h10408000;
      12620: inst = 32'hc404994;
      12621: inst = 32'h8220000;
      12622: inst = 32'h10408000;
      12623: inst = 32'hc404995;
      12624: inst = 32'h8220000;
      12625: inst = 32'h10408000;
      12626: inst = 32'hc4049f3;
      12627: inst = 32'h8220000;
      12628: inst = 32'h10408000;
      12629: inst = 32'hc4049f4;
      12630: inst = 32'h8220000;
      12631: inst = 32'h10408000;
      12632: inst = 32'hc4049f5;
      12633: inst = 32'h8220000;
      12634: inst = 32'h10408000;
      12635: inst = 32'hc404a53;
      12636: inst = 32'h8220000;
      12637: inst = 32'h10408000;
      12638: inst = 32'hc404a54;
      12639: inst = 32'h8220000;
      12640: inst = 32'h10408000;
      12641: inst = 32'hc404a55;
      12642: inst = 32'h8220000;
      12643: inst = 32'h10408000;
      12644: inst = 32'hc404ab2;
      12645: inst = 32'h8220000;
      12646: inst = 32'h10408000;
      12647: inst = 32'hc404ab3;
      12648: inst = 32'h8220000;
      12649: inst = 32'h10408000;
      12650: inst = 32'hc404ab5;
      12651: inst = 32'h8220000;
      12652: inst = 32'h10408000;
      12653: inst = 32'hc404b12;
      12654: inst = 32'h8220000;
      12655: inst = 32'h10408000;
      12656: inst = 32'hc404b13;
      12657: inst = 32'h8220000;
      12658: inst = 32'h10408000;
      12659: inst = 32'hc404b15;
      12660: inst = 32'h8220000;
      12661: inst = 32'h10408000;
      12662: inst = 32'hc404b72;
      12663: inst = 32'h8220000;
      12664: inst = 32'h10408000;
      12665: inst = 32'hc404b73;
      12666: inst = 32'h8220000;
      12667: inst = 32'h10408000;
      12668: inst = 32'hc404b74;
      12669: inst = 32'h8220000;
      12670: inst = 32'h10408000;
      12671: inst = 32'hc404b75;
      12672: inst = 32'h8220000;
      12673: inst = 32'hc20eed7;
      12674: inst = 32'h10408000;
      12675: inst = 32'hc404a08;
      12676: inst = 32'h8220000;
      12677: inst = 32'h10408000;
      12678: inst = 32'hc404a0e;
      12679: inst = 32'h8220000;
      12680: inst = 32'hc20e6fa;
      12681: inst = 32'h10408000;
      12682: inst = 32'hc404a09;
      12683: inst = 32'h8220000;
      12684: inst = 32'h10408000;
      12685: inst = 32'hc404a0d;
      12686: inst = 32'h8220000;
      12687: inst = 32'h10408000;
      12688: inst = 32'hc404be7;
      12689: inst = 32'h8220000;
      12690: inst = 32'hc20e6fb;
      12691: inst = 32'h10408000;
      12692: inst = 32'hc404a0a;
      12693: inst = 32'h8220000;
      12694: inst = 32'h10408000;
      12695: inst = 32'hc404a0c;
      12696: inst = 32'h8220000;
      12697: inst = 32'h10408000;
      12698: inst = 32'hc404ac7;
      12699: inst = 32'h8220000;
      12700: inst = 32'h10408000;
      12701: inst = 32'hc404acf;
      12702: inst = 32'h8220000;
      12703: inst = 32'h10408000;
      12704: inst = 32'hc404b87;
      12705: inst = 32'h8220000;
      12706: inst = 32'h10408000;
      12707: inst = 32'hc404b8f;
      12708: inst = 32'h8220000;
      12709: inst = 32'h10408000;
      12710: inst = 32'hc404c4d;
      12711: inst = 32'h8220000;
      12712: inst = 32'hc20defb;
      12713: inst = 32'h10408000;
      12714: inst = 32'hc404a0b;
      12715: inst = 32'h8220000;
      12716: inst = 32'h10408000;
      12717: inst = 32'hc404a68;
      12718: inst = 32'h8220000;
      12719: inst = 32'h10408000;
      12720: inst = 32'hc404a69;
      12721: inst = 32'h8220000;
      12722: inst = 32'h10408000;
      12723: inst = 32'hc404a6a;
      12724: inst = 32'h8220000;
      12725: inst = 32'h10408000;
      12726: inst = 32'hc404a6b;
      12727: inst = 32'h8220000;
      12728: inst = 32'h10408000;
      12729: inst = 32'hc404a6c;
      12730: inst = 32'h8220000;
      12731: inst = 32'h10408000;
      12732: inst = 32'hc404a6d;
      12733: inst = 32'h8220000;
      12734: inst = 32'h10408000;
      12735: inst = 32'hc404a6e;
      12736: inst = 32'h8220000;
      12737: inst = 32'h10408000;
      12738: inst = 32'hc404ac8;
      12739: inst = 32'h8220000;
      12740: inst = 32'h10408000;
      12741: inst = 32'hc404ac9;
      12742: inst = 32'h8220000;
      12743: inst = 32'h10408000;
      12744: inst = 32'hc404aca;
      12745: inst = 32'h8220000;
      12746: inst = 32'h10408000;
      12747: inst = 32'hc404acb;
      12748: inst = 32'h8220000;
      12749: inst = 32'h10408000;
      12750: inst = 32'hc404acc;
      12751: inst = 32'h8220000;
      12752: inst = 32'h10408000;
      12753: inst = 32'hc404acd;
      12754: inst = 32'h8220000;
      12755: inst = 32'h10408000;
      12756: inst = 32'hc404ace;
      12757: inst = 32'h8220000;
      12758: inst = 32'h10408000;
      12759: inst = 32'hc404b27;
      12760: inst = 32'h8220000;
      12761: inst = 32'h10408000;
      12762: inst = 32'hc404b2a;
      12763: inst = 32'h8220000;
      12764: inst = 32'h10408000;
      12765: inst = 32'hc404b2d;
      12766: inst = 32'h8220000;
      12767: inst = 32'h10408000;
      12768: inst = 32'hc404b2e;
      12769: inst = 32'h8220000;
      12770: inst = 32'h10408000;
      12771: inst = 32'hc404b2f;
      12772: inst = 32'h8220000;
      12773: inst = 32'h10408000;
      12774: inst = 32'hc404b8a;
      12775: inst = 32'h8220000;
      12776: inst = 32'h10408000;
      12777: inst = 32'hc404b8d;
      12778: inst = 32'h8220000;
      12779: inst = 32'h10408000;
      12780: inst = 32'hc404b8e;
      12781: inst = 32'h8220000;
      12782: inst = 32'h10408000;
      12783: inst = 32'hc404be8;
      12784: inst = 32'h8220000;
      12785: inst = 32'h10408000;
      12786: inst = 32'hc404be9;
      12787: inst = 32'h8220000;
      12788: inst = 32'h10408000;
      12789: inst = 32'hc404bea;
      12790: inst = 32'h8220000;
      12791: inst = 32'h10408000;
      12792: inst = 32'hc404beb;
      12793: inst = 32'h8220000;
      12794: inst = 32'h10408000;
      12795: inst = 32'hc404bec;
      12796: inst = 32'h8220000;
      12797: inst = 32'h10408000;
      12798: inst = 32'hc404bed;
      12799: inst = 32'h8220000;
      12800: inst = 32'h10408000;
      12801: inst = 32'hc404bee;
      12802: inst = 32'h8220000;
      12803: inst = 32'h10408000;
      12804: inst = 32'hc404c49;
      12805: inst = 32'h8220000;
      12806: inst = 32'h10408000;
      12807: inst = 32'hc404c4b;
      12808: inst = 32'h8220000;
      12809: inst = 32'h10408000;
      12810: inst = 32'hc404ca9;
      12811: inst = 32'h8220000;
      12812: inst = 32'h10408000;
      12813: inst = 32'hc404cab;
      12814: inst = 32'h8220000;
      12815: inst = 32'hc20eed8;
      12816: inst = 32'h10408000;
      12817: inst = 32'hc404a67;
      12818: inst = 32'h8220000;
      12819: inst = 32'h10408000;
      12820: inst = 32'hc404a6f;
      12821: inst = 32'h8220000;
      12822: inst = 32'hc204a69;
      12823: inst = 32'h10408000;
      12824: inst = 32'hc404b28;
      12825: inst = 32'h8220000;
      12826: inst = 32'h10408000;
      12827: inst = 32'hc404b29;
      12828: inst = 32'h8220000;
      12829: inst = 32'h10408000;
      12830: inst = 32'hc404b2b;
      12831: inst = 32'h8220000;
      12832: inst = 32'h10408000;
      12833: inst = 32'hc404b2c;
      12834: inst = 32'h8220000;
      12835: inst = 32'h10408000;
      12836: inst = 32'hc404b88;
      12837: inst = 32'h8220000;
      12838: inst = 32'h10408000;
      12839: inst = 32'hc404b89;
      12840: inst = 32'h8220000;
      12841: inst = 32'h10408000;
      12842: inst = 32'hc404b8b;
      12843: inst = 32'h8220000;
      12844: inst = 32'h10408000;
      12845: inst = 32'hc404b8c;
      12846: inst = 32'h8220000;
      12847: inst = 32'h10408000;
      12848: inst = 32'hc404c48;
      12849: inst = 32'h8220000;
      12850: inst = 32'h10408000;
      12851: inst = 32'hc404c4a;
      12852: inst = 32'h8220000;
      12853: inst = 32'h10408000;
      12854: inst = 32'hc404c4c;
      12855: inst = 32'h8220000;
      12856: inst = 32'h10408000;
      12857: inst = 32'hc404ca8;
      12858: inst = 32'h8220000;
      12859: inst = 32'h10408000;
      12860: inst = 32'hc404caa;
      12861: inst = 32'h8220000;
      12862: inst = 32'h10408000;
      12863: inst = 32'hc404cac;
      12864: inst = 32'h8220000;
      12865: inst = 32'h10408000;
      12866: inst = 32'hc405085;
      12867: inst = 32'h8220000;
      12868: inst = 32'h10408000;
      12869: inst = 32'hc40509a;
      12870: inst = 32'h8220000;
      12871: inst = 32'h10408000;
      12872: inst = 32'hc4050e4;
      12873: inst = 32'h8220000;
      12874: inst = 32'h10408000;
      12875: inst = 32'hc4050e5;
      12876: inst = 32'h8220000;
      12877: inst = 32'h10408000;
      12878: inst = 32'hc4050fa;
      12879: inst = 32'h8220000;
      12880: inst = 32'h10408000;
      12881: inst = 32'hc4050fb;
      12882: inst = 32'h8220000;
      12883: inst = 32'h10408000;
      12884: inst = 32'hc405143;
      12885: inst = 32'h8220000;
      12886: inst = 32'h10408000;
      12887: inst = 32'hc405144;
      12888: inst = 32'h8220000;
      12889: inst = 32'h10408000;
      12890: inst = 32'hc405145;
      12891: inst = 32'h8220000;
      12892: inst = 32'h10408000;
      12893: inst = 32'hc40515a;
      12894: inst = 32'h8220000;
      12895: inst = 32'h10408000;
      12896: inst = 32'hc40515b;
      12897: inst = 32'h8220000;
      12898: inst = 32'h10408000;
      12899: inst = 32'hc40515c;
      12900: inst = 32'h8220000;
      12901: inst = 32'h10408000;
      12902: inst = 32'hc4051a2;
      12903: inst = 32'h8220000;
      12904: inst = 32'h10408000;
      12905: inst = 32'hc4051a3;
      12906: inst = 32'h8220000;
      12907: inst = 32'h10408000;
      12908: inst = 32'hc4051a4;
      12909: inst = 32'h8220000;
      12910: inst = 32'h10408000;
      12911: inst = 32'hc4051a5;
      12912: inst = 32'h8220000;
      12913: inst = 32'h10408000;
      12914: inst = 32'hc4051ba;
      12915: inst = 32'h8220000;
      12916: inst = 32'h10408000;
      12917: inst = 32'hc4051bb;
      12918: inst = 32'h8220000;
      12919: inst = 32'h10408000;
      12920: inst = 32'hc4051bc;
      12921: inst = 32'h8220000;
      12922: inst = 32'h10408000;
      12923: inst = 32'hc4051bd;
      12924: inst = 32'h8220000;
      12925: inst = 32'h10408000;
      12926: inst = 32'hc405202;
      12927: inst = 32'h8220000;
      12928: inst = 32'h10408000;
      12929: inst = 32'hc405203;
      12930: inst = 32'h8220000;
      12931: inst = 32'h10408000;
      12932: inst = 32'hc405204;
      12933: inst = 32'h8220000;
      12934: inst = 32'h10408000;
      12935: inst = 32'hc405205;
      12936: inst = 32'h8220000;
      12937: inst = 32'h10408000;
      12938: inst = 32'hc40521a;
      12939: inst = 32'h8220000;
      12940: inst = 32'h10408000;
      12941: inst = 32'hc40521b;
      12942: inst = 32'h8220000;
      12943: inst = 32'h10408000;
      12944: inst = 32'hc40521c;
      12945: inst = 32'h8220000;
      12946: inst = 32'h10408000;
      12947: inst = 32'hc40521d;
      12948: inst = 32'h8220000;
      12949: inst = 32'h10408000;
      12950: inst = 32'hc405262;
      12951: inst = 32'h8220000;
      12952: inst = 32'h10408000;
      12953: inst = 32'hc405263;
      12954: inst = 32'h8220000;
      12955: inst = 32'h10408000;
      12956: inst = 32'hc405264;
      12957: inst = 32'h8220000;
      12958: inst = 32'h10408000;
      12959: inst = 32'hc405265;
      12960: inst = 32'h8220000;
      12961: inst = 32'h10408000;
      12962: inst = 32'hc40527a;
      12963: inst = 32'h8220000;
      12964: inst = 32'h10408000;
      12965: inst = 32'hc40527b;
      12966: inst = 32'h8220000;
      12967: inst = 32'h10408000;
      12968: inst = 32'hc40527c;
      12969: inst = 32'h8220000;
      12970: inst = 32'h10408000;
      12971: inst = 32'hc40527d;
      12972: inst = 32'h8220000;
      12973: inst = 32'h10408000;
      12974: inst = 32'hc4052c2;
      12975: inst = 32'h8220000;
      12976: inst = 32'h10408000;
      12977: inst = 32'hc4052c3;
      12978: inst = 32'h8220000;
      12979: inst = 32'h10408000;
      12980: inst = 32'hc4052c4;
      12981: inst = 32'h8220000;
      12982: inst = 32'h10408000;
      12983: inst = 32'hc4052db;
      12984: inst = 32'h8220000;
      12985: inst = 32'h10408000;
      12986: inst = 32'hc4052dc;
      12987: inst = 32'h8220000;
      12988: inst = 32'h10408000;
      12989: inst = 32'hc4052dd;
      12990: inst = 32'h8220000;
      12991: inst = 32'h10408000;
      12992: inst = 32'hc405322;
      12993: inst = 32'h8220000;
      12994: inst = 32'h10408000;
      12995: inst = 32'hc405323;
      12996: inst = 32'h8220000;
      12997: inst = 32'h10408000;
      12998: inst = 32'hc405324;
      12999: inst = 32'h8220000;
      13000: inst = 32'h10408000;
      13001: inst = 32'hc40533b;
      13002: inst = 32'h8220000;
      13003: inst = 32'h10408000;
      13004: inst = 32'hc40533c;
      13005: inst = 32'h8220000;
      13006: inst = 32'h10408000;
      13007: inst = 32'hc40533d;
      13008: inst = 32'h8220000;
      13009: inst = 32'h10408000;
      13010: inst = 32'hc40537f;
      13011: inst = 32'h8220000;
      13012: inst = 32'h10408000;
      13013: inst = 32'hc405382;
      13014: inst = 32'h8220000;
      13015: inst = 32'h10408000;
      13016: inst = 32'hc405383;
      13017: inst = 32'h8220000;
      13018: inst = 32'h10408000;
      13019: inst = 32'hc405384;
      13020: inst = 32'h8220000;
      13021: inst = 32'h10408000;
      13022: inst = 32'hc40539b;
      13023: inst = 32'h8220000;
      13024: inst = 32'h10408000;
      13025: inst = 32'hc40539c;
      13026: inst = 32'h8220000;
      13027: inst = 32'h10408000;
      13028: inst = 32'hc40539d;
      13029: inst = 32'h8220000;
      13030: inst = 32'h10408000;
      13031: inst = 32'hc4053a0;
      13032: inst = 32'h8220000;
      13033: inst = 32'h10408000;
      13034: inst = 32'hc4053de;
      13035: inst = 32'h8220000;
      13036: inst = 32'h10408000;
      13037: inst = 32'hc4053df;
      13038: inst = 32'h8220000;
      13039: inst = 32'h10408000;
      13040: inst = 32'hc4053e2;
      13041: inst = 32'h8220000;
      13042: inst = 32'h10408000;
      13043: inst = 32'hc4053e3;
      13044: inst = 32'h8220000;
      13045: inst = 32'h10408000;
      13046: inst = 32'hc4053fc;
      13047: inst = 32'h8220000;
      13048: inst = 32'h10408000;
      13049: inst = 32'hc4053fd;
      13050: inst = 32'h8220000;
      13051: inst = 32'h10408000;
      13052: inst = 32'hc405400;
      13053: inst = 32'h8220000;
      13054: inst = 32'h10408000;
      13055: inst = 32'hc405401;
      13056: inst = 32'h8220000;
      13057: inst = 32'h10408000;
      13058: inst = 32'hc40543d;
      13059: inst = 32'h8220000;
      13060: inst = 32'h10408000;
      13061: inst = 32'hc40543e;
      13062: inst = 32'h8220000;
      13063: inst = 32'h10408000;
      13064: inst = 32'hc40543f;
      13065: inst = 32'h8220000;
      13066: inst = 32'h10408000;
      13067: inst = 32'hc405442;
      13068: inst = 32'h8220000;
      13069: inst = 32'h10408000;
      13070: inst = 32'hc405443;
      13071: inst = 32'h8220000;
      13072: inst = 32'h10408000;
      13073: inst = 32'hc40545c;
      13074: inst = 32'h8220000;
      13075: inst = 32'h10408000;
      13076: inst = 32'hc40545d;
      13077: inst = 32'h8220000;
      13078: inst = 32'h10408000;
      13079: inst = 32'hc405460;
      13080: inst = 32'h8220000;
      13081: inst = 32'h10408000;
      13082: inst = 32'hc405461;
      13083: inst = 32'h8220000;
      13084: inst = 32'h10408000;
      13085: inst = 32'hc405462;
      13086: inst = 32'h8220000;
      13087: inst = 32'h10408000;
      13088: inst = 32'hc40549d;
      13089: inst = 32'h8220000;
      13090: inst = 32'h10408000;
      13091: inst = 32'hc40549e;
      13092: inst = 32'h8220000;
      13093: inst = 32'h10408000;
      13094: inst = 32'hc4054a0;
      13095: inst = 32'h8220000;
      13096: inst = 32'h10408000;
      13097: inst = 32'hc4054a1;
      13098: inst = 32'h8220000;
      13099: inst = 32'h10408000;
      13100: inst = 32'hc4054a2;
      13101: inst = 32'h8220000;
      13102: inst = 32'h10408000;
      13103: inst = 32'hc4054a3;
      13104: inst = 32'h8220000;
      13105: inst = 32'h10408000;
      13106: inst = 32'hc4054bc;
      13107: inst = 32'h8220000;
      13108: inst = 32'h10408000;
      13109: inst = 32'hc4054bd;
      13110: inst = 32'h8220000;
      13111: inst = 32'h10408000;
      13112: inst = 32'hc4054be;
      13113: inst = 32'h8220000;
      13114: inst = 32'h10408000;
      13115: inst = 32'hc4054bf;
      13116: inst = 32'h8220000;
      13117: inst = 32'h10408000;
      13118: inst = 32'hc4054c1;
      13119: inst = 32'h8220000;
      13120: inst = 32'h10408000;
      13121: inst = 32'hc4054c2;
      13122: inst = 32'h8220000;
      13123: inst = 32'h10408000;
      13124: inst = 32'hc4054fc;
      13125: inst = 32'h8220000;
      13126: inst = 32'h10408000;
      13127: inst = 32'hc4054fd;
      13128: inst = 32'h8220000;
      13129: inst = 32'h10408000;
      13130: inst = 32'hc4054fe;
      13131: inst = 32'h8220000;
      13132: inst = 32'h10408000;
      13133: inst = 32'hc405502;
      13134: inst = 32'h8220000;
      13135: inst = 32'h10408000;
      13136: inst = 32'hc40551d;
      13137: inst = 32'h8220000;
      13138: inst = 32'h10408000;
      13139: inst = 32'hc405521;
      13140: inst = 32'h8220000;
      13141: inst = 32'h10408000;
      13142: inst = 32'hc405522;
      13143: inst = 32'h8220000;
      13144: inst = 32'h10408000;
      13145: inst = 32'hc405523;
      13146: inst = 32'h8220000;
      13147: inst = 32'h10408000;
      13148: inst = 32'hc40555b;
      13149: inst = 32'h8220000;
      13150: inst = 32'h10408000;
      13151: inst = 32'hc40555c;
      13152: inst = 32'h8220000;
      13153: inst = 32'h10408000;
      13154: inst = 32'hc40555d;
      13155: inst = 32'h8220000;
      13156: inst = 32'h10408000;
      13157: inst = 32'hc405562;
      13158: inst = 32'h8220000;
      13159: inst = 32'h10408000;
      13160: inst = 32'hc40557d;
      13161: inst = 32'h8220000;
      13162: inst = 32'h10408000;
      13163: inst = 32'hc405582;
      13164: inst = 32'h8220000;
      13165: inst = 32'h10408000;
      13166: inst = 32'hc405583;
      13167: inst = 32'h8220000;
      13168: inst = 32'h10408000;
      13169: inst = 32'hc405584;
      13170: inst = 32'h8220000;
      13171: inst = 32'h10408000;
      13172: inst = 32'hc4055ba;
      13173: inst = 32'h8220000;
      13174: inst = 32'h10408000;
      13175: inst = 32'hc4055bb;
      13176: inst = 32'h8220000;
      13177: inst = 32'h10408000;
      13178: inst = 32'hc4055bc;
      13179: inst = 32'h8220000;
      13180: inst = 32'h10408000;
      13181: inst = 32'hc4055bd;
      13182: inst = 32'h8220000;
      13183: inst = 32'h10408000;
      13184: inst = 32'hc4055c2;
      13185: inst = 32'h8220000;
      13186: inst = 32'h10408000;
      13187: inst = 32'hc4055dd;
      13188: inst = 32'h8220000;
      13189: inst = 32'h10408000;
      13190: inst = 32'hc4055e2;
      13191: inst = 32'h8220000;
      13192: inst = 32'h10408000;
      13193: inst = 32'hc4055e3;
      13194: inst = 32'h8220000;
      13195: inst = 32'h10408000;
      13196: inst = 32'hc4055e4;
      13197: inst = 32'h8220000;
      13198: inst = 32'h10408000;
      13199: inst = 32'hc4055e5;
      13200: inst = 32'h8220000;
      13201: inst = 32'h10408000;
      13202: inst = 32'hc40561a;
      13203: inst = 32'h8220000;
      13204: inst = 32'h10408000;
      13205: inst = 32'hc40561b;
      13206: inst = 32'h8220000;
      13207: inst = 32'h10408000;
      13208: inst = 32'hc40561c;
      13209: inst = 32'h8220000;
      13210: inst = 32'h10408000;
      13211: inst = 32'hc40561d;
      13212: inst = 32'h8220000;
      13213: inst = 32'h10408000;
      13214: inst = 32'hc405642;
      13215: inst = 32'h8220000;
      13216: inst = 32'h10408000;
      13217: inst = 32'hc405643;
      13218: inst = 32'h8220000;
      13219: inst = 32'h10408000;
      13220: inst = 32'hc405644;
      13221: inst = 32'h8220000;
      13222: inst = 32'h10408000;
      13223: inst = 32'hc405645;
      13224: inst = 32'h8220000;
      13225: inst = 32'h10408000;
      13226: inst = 32'hc405679;
      13227: inst = 32'h8220000;
      13228: inst = 32'h10408000;
      13229: inst = 32'hc40567a;
      13230: inst = 32'h8220000;
      13231: inst = 32'h10408000;
      13232: inst = 32'hc40567b;
      13233: inst = 32'h8220000;
      13234: inst = 32'h10408000;
      13235: inst = 32'hc40567c;
      13236: inst = 32'h8220000;
      13237: inst = 32'h10408000;
      13238: inst = 32'hc4056a3;
      13239: inst = 32'h8220000;
      13240: inst = 32'h10408000;
      13241: inst = 32'hc4056a4;
      13242: inst = 32'h8220000;
      13243: inst = 32'h10408000;
      13244: inst = 32'hc4056a5;
      13245: inst = 32'h8220000;
      13246: inst = 32'h10408000;
      13247: inst = 32'hc4056a6;
      13248: inst = 32'h8220000;
      13249: inst = 32'hc20e6d9;
      13250: inst = 32'h10408000;
      13251: inst = 32'hc404bef;
      13252: inst = 32'h8220000;
      13253: inst = 32'h10408000;
      13254: inst = 32'hc404c4e;
      13255: inst = 32'h8220000;
      13256: inst = 32'hc20eeb7;
      13257: inst = 32'h10408000;
      13258: inst = 32'hc404c47;
      13259: inst = 32'h8220000;
      13260: inst = 32'hc20d615;
      13261: inst = 32'h10408000;
      13262: inst = 32'hc404ca2;
      13263: inst = 32'h8220000;
      13264: inst = 32'h10408000;
      13265: inst = 32'hc404d00;
      13266: inst = 32'h8220000;
      13267: inst = 32'hc209c91;
      13268: inst = 32'h10408000;
      13269: inst = 32'hc404ca3;
      13270: inst = 32'h8220000;
      13271: inst = 32'h10408000;
      13272: inst = 32'hc404d01;
      13273: inst = 32'h8220000;
      13274: inst = 32'hc207bf0;
      13275: inst = 32'h10408000;
      13276: inst = 32'hc404ca4;
      13277: inst = 32'h8220000;
      13278: inst = 32'h10408000;
      13279: inst = 32'hc404ca5;
      13280: inst = 32'h8220000;
      13281: inst = 32'h10408000;
      13282: inst = 32'hc404ca6;
      13283: inst = 32'h8220000;
      13284: inst = 32'h10408000;
      13285: inst = 32'hc404ca7;
      13286: inst = 32'h8220000;
      13287: inst = 32'h10408000;
      13288: inst = 32'hc404d02;
      13289: inst = 32'h8220000;
      13290: inst = 32'h10408000;
      13291: inst = 32'hc404d03;
      13292: inst = 32'h8220000;
      13293: inst = 32'h10408000;
      13294: inst = 32'hc404d04;
      13295: inst = 32'h8220000;
      13296: inst = 32'h10408000;
      13297: inst = 32'hc404d05;
      13298: inst = 32'h8220000;
      13299: inst = 32'h10408000;
      13300: inst = 32'hc404d06;
      13301: inst = 32'h8220000;
      13302: inst = 32'h10408000;
      13303: inst = 32'hc404d07;
      13304: inst = 32'h8220000;
      13305: inst = 32'h10408000;
      13306: inst = 32'hc404d08;
      13307: inst = 32'h8220000;
      13308: inst = 32'h10408000;
      13309: inst = 32'hc404d09;
      13310: inst = 32'h8220000;
      13311: inst = 32'h10408000;
      13312: inst = 32'hc404d0a;
      13313: inst = 32'h8220000;
      13314: inst = 32'h10408000;
      13315: inst = 32'hc404d0b;
      13316: inst = 32'h8220000;
      13317: inst = 32'h10408000;
      13318: inst = 32'hc404d0c;
      13319: inst = 32'h8220000;
      13320: inst = 32'h10408000;
      13321: inst = 32'hc404d0d;
      13322: inst = 32'h8220000;
      13323: inst = 32'h10408000;
      13324: inst = 32'hc404d0e;
      13325: inst = 32'h8220000;
      13326: inst = 32'h10408000;
      13327: inst = 32'hc404d0f;
      13328: inst = 32'h8220000;
      13329: inst = 32'h10408000;
      13330: inst = 32'hc404d10;
      13331: inst = 32'h8220000;
      13332: inst = 32'h10408000;
      13333: inst = 32'hc404d11;
      13334: inst = 32'h8220000;
      13335: inst = 32'h10408000;
      13336: inst = 32'hc404d12;
      13337: inst = 32'h8220000;
      13338: inst = 32'h10408000;
      13339: inst = 32'hc404d13;
      13340: inst = 32'h8220000;
      13341: inst = 32'h10408000;
      13342: inst = 32'hc404d14;
      13343: inst = 32'h8220000;
      13344: inst = 32'h10408000;
      13345: inst = 32'hc4055c3;
      13346: inst = 32'h8220000;
      13347: inst = 32'h10408000;
      13348: inst = 32'hc4055dc;
      13349: inst = 32'h8220000;
      13350: inst = 32'hc20ad55;
      13351: inst = 32'h10408000;
      13352: inst = 32'hc404cad;
      13353: inst = 32'h8220000;
      13354: inst = 32'hc208410;
      13355: inst = 32'h10408000;
      13356: inst = 32'hc404cae;
      13357: inst = 32'h8220000;
      13358: inst = 32'h10408000;
      13359: inst = 32'hc404caf;
      13360: inst = 32'h8220000;
      13361: inst = 32'h10408000;
      13362: inst = 32'hc404cb0;
      13363: inst = 32'h8220000;
      13364: inst = 32'h10408000;
      13365: inst = 32'hc404cb1;
      13366: inst = 32'h8220000;
      13367: inst = 32'h10408000;
      13368: inst = 32'hc404cb2;
      13369: inst = 32'h8220000;
      13370: inst = 32'h10408000;
      13371: inst = 32'hc404cb3;
      13372: inst = 32'h8220000;
      13373: inst = 32'h10408000;
      13374: inst = 32'hc404cb4;
      13375: inst = 32'h8220000;
      13376: inst = 32'h10408000;
      13377: inst = 32'hc404cb5;
      13378: inst = 32'h8220000;
      13379: inst = 32'h10408000;
      13380: inst = 32'hc40537d;
      13381: inst = 32'h8220000;
      13382: inst = 32'h10408000;
      13383: inst = 32'hc405385;
      13384: inst = 32'h8220000;
      13385: inst = 32'h10408000;
      13386: inst = 32'hc40539a;
      13387: inst = 32'h8220000;
      13388: inst = 32'h10408000;
      13389: inst = 32'hc4053a2;
      13390: inst = 32'h8220000;
      13391: inst = 32'h10408000;
      13392: inst = 32'hc4054a4;
      13393: inst = 32'h8220000;
      13394: inst = 32'h10408000;
      13395: inst = 32'hc4054bb;
      13396: inst = 32'h8220000;
      13397: inst = 32'h10408000;
      13398: inst = 32'hc405741;
      13399: inst = 32'h8220000;
      13400: inst = 32'h10408000;
      13401: inst = 32'hc40575e;
      13402: inst = 32'h8220000;
      13403: inst = 32'hc209470;
      13404: inst = 32'h10408000;
      13405: inst = 32'hc404cb6;
      13406: inst = 32'h8220000;
      13407: inst = 32'h10408000;
      13408: inst = 32'hc404d15;
      13409: inst = 32'h8220000;
      13410: inst = 32'hc20a534;
      13411: inst = 32'h10408000;
      13412: inst = 32'hc404cfb;
      13413: inst = 32'h8220000;
      13414: inst = 32'hc208c51;
      13415: inst = 32'h10408000;
      13416: inst = 32'hc404cfc;
      13417: inst = 32'h8220000;
      13418: inst = 32'h10408000;
      13419: inst = 32'hc404cfd;
      13420: inst = 32'h8220000;
      13421: inst = 32'h10408000;
      13422: inst = 32'hc4053da;
      13423: inst = 32'h8220000;
      13424: inst = 32'h10408000;
      13425: inst = 32'hc4053dc;
      13426: inst = 32'h8220000;
      13427: inst = 32'h10408000;
      13428: inst = 32'hc405403;
      13429: inst = 32'h8220000;
      13430: inst = 32'h10408000;
      13431: inst = 32'hc405405;
      13432: inst = 32'h8220000;
      13433: inst = 32'h10408000;
      13434: inst = 32'hc4054fa;
      13435: inst = 32'h8220000;
      13436: inst = 32'h10408000;
      13437: inst = 32'hc405525;
      13438: inst = 32'h8220000;
      13439: inst = 32'h10408000;
      13440: inst = 32'hc405557;
      13441: inst = 32'h8220000;
      13442: inst = 32'h10408000;
      13443: inst = 32'hc40555f;
      13444: inst = 32'h8220000;
      13445: inst = 32'h10408000;
      13446: inst = 32'hc405580;
      13447: inst = 32'h8220000;
      13448: inst = 32'h10408000;
      13449: inst = 32'hc405588;
      13450: inst = 32'h8220000;
      13451: inst = 32'h10408000;
      13452: inst = 32'hc405618;
      13453: inst = 32'h8220000;
      13454: inst = 32'h10408000;
      13455: inst = 32'hc405627;
      13456: inst = 32'h8220000;
      13457: inst = 32'h10408000;
      13458: inst = 32'hc405638;
      13459: inst = 32'h8220000;
      13460: inst = 32'h10408000;
      13461: inst = 32'hc405647;
      13462: inst = 32'h8220000;
      13463: inst = 32'h10408000;
      13464: inst = 32'hc40570b;
      13465: inst = 32'h8220000;
      13466: inst = 32'hc206b6d;
      13467: inst = 32'h10408000;
      13468: inst = 32'hc404d16;
      13469: inst = 32'h8220000;
      13470: inst = 32'h10408000;
      13471: inst = 32'hc404d75;
      13472: inst = 32'h8220000;
      13473: inst = 32'h10408000;
      13474: inst = 32'hc404d76;
      13475: inst = 32'h8220000;
      13476: inst = 32'h10408000;
      13477: inst = 32'hc404dd5;
      13478: inst = 32'h8220000;
      13479: inst = 32'h10408000;
      13480: inst = 32'hc404dd6;
      13481: inst = 32'h8220000;
      13482: inst = 32'h10408000;
      13483: inst = 32'hc404e35;
      13484: inst = 32'h8220000;
      13485: inst = 32'h10408000;
      13486: inst = 32'hc404e36;
      13487: inst = 32'h8220000;
      13488: inst = 32'h10408000;
      13489: inst = 32'hc404e95;
      13490: inst = 32'h8220000;
      13491: inst = 32'h10408000;
      13492: inst = 32'hc404e96;
      13493: inst = 32'h8220000;
      13494: inst = 32'h10408000;
      13495: inst = 32'hc404ef5;
      13496: inst = 32'h8220000;
      13497: inst = 32'h10408000;
      13498: inst = 32'hc404ef6;
      13499: inst = 32'h8220000;
      13500: inst = 32'h10408000;
      13501: inst = 32'hc404f55;
      13502: inst = 32'h8220000;
      13503: inst = 32'h10408000;
      13504: inst = 32'hc404f56;
      13505: inst = 32'h8220000;
      13506: inst = 32'h10408000;
      13507: inst = 32'hc404fb5;
      13508: inst = 32'h8220000;
      13509: inst = 32'h10408000;
      13510: inst = 32'hc404fb6;
      13511: inst = 32'h8220000;
      13512: inst = 32'h10408000;
      13513: inst = 32'hc405015;
      13514: inst = 32'h8220000;
      13515: inst = 32'h10408000;
      13516: inst = 32'hc405016;
      13517: inst = 32'h8220000;
      13518: inst = 32'h10408000;
      13519: inst = 32'hc405075;
      13520: inst = 32'h8220000;
      13521: inst = 32'h10408000;
      13522: inst = 32'hc405076;
      13523: inst = 32'h8220000;
      13524: inst = 32'h10408000;
      13525: inst = 32'hc4050d5;
      13526: inst = 32'h8220000;
      13527: inst = 32'h10408000;
      13528: inst = 32'hc4050d6;
      13529: inst = 32'h8220000;
      13530: inst = 32'h10408000;
      13531: inst = 32'hc405135;
      13532: inst = 32'h8220000;
      13533: inst = 32'h10408000;
      13534: inst = 32'hc405136;
      13535: inst = 32'h8220000;
      13536: inst = 32'h10408000;
      13537: inst = 32'hc405195;
      13538: inst = 32'h8220000;
      13539: inst = 32'h10408000;
      13540: inst = 32'hc405196;
      13541: inst = 32'h8220000;
      13542: inst = 32'h10408000;
      13543: inst = 32'hc4051f5;
      13544: inst = 32'h8220000;
      13545: inst = 32'h10408000;
      13546: inst = 32'hc4051f6;
      13547: inst = 32'h8220000;
      13548: inst = 32'h10408000;
      13549: inst = 32'hc405255;
      13550: inst = 32'h8220000;
      13551: inst = 32'h10408000;
      13552: inst = 32'hc405256;
      13553: inst = 32'h8220000;
      13554: inst = 32'h10408000;
      13555: inst = 32'hc4052b5;
      13556: inst = 32'h8220000;
      13557: inst = 32'h10408000;
      13558: inst = 32'hc4052b6;
      13559: inst = 32'h8220000;
      13560: inst = 32'h10408000;
      13561: inst = 32'hc405325;
      13562: inst = 32'h8220000;
      13563: inst = 32'h10408000;
      13564: inst = 32'hc40533a;
      13565: inst = 32'h8220000;
      13566: inst = 32'hc20c638;
      13567: inst = 32'h10408000;
      13568: inst = 32'hc404d5b;
      13569: inst = 32'h8220000;
      13570: inst = 32'hc208c71;
      13571: inst = 32'h10408000;
      13572: inst = 32'hc404d60;
      13573: inst = 32'h8220000;
      13574: inst = 32'h10408000;
      13575: inst = 32'hc404d61;
      13576: inst = 32'h8220000;
      13577: inst = 32'h10408000;
      13578: inst = 32'hc404d62;
      13579: inst = 32'h8220000;
      13580: inst = 32'h10408000;
      13581: inst = 32'hc404d63;
      13582: inst = 32'h8220000;
      13583: inst = 32'h10408000;
      13584: inst = 32'hc404d64;
      13585: inst = 32'h8220000;
      13586: inst = 32'h10408000;
      13587: inst = 32'hc404d65;
      13588: inst = 32'h8220000;
      13589: inst = 32'h10408000;
      13590: inst = 32'hc404d66;
      13591: inst = 32'h8220000;
      13592: inst = 32'h10408000;
      13593: inst = 32'hc404d67;
      13594: inst = 32'h8220000;
      13595: inst = 32'h10408000;
      13596: inst = 32'hc404d68;
      13597: inst = 32'h8220000;
      13598: inst = 32'h10408000;
      13599: inst = 32'hc404d69;
      13600: inst = 32'h8220000;
      13601: inst = 32'h10408000;
      13602: inst = 32'hc404d6a;
      13603: inst = 32'h8220000;
      13604: inst = 32'h10408000;
      13605: inst = 32'hc404d6b;
      13606: inst = 32'h8220000;
      13607: inst = 32'h10408000;
      13608: inst = 32'hc404d6c;
      13609: inst = 32'h8220000;
      13610: inst = 32'h10408000;
      13611: inst = 32'hc404d6d;
      13612: inst = 32'h8220000;
      13613: inst = 32'h10408000;
      13614: inst = 32'hc404d6e;
      13615: inst = 32'h8220000;
      13616: inst = 32'h10408000;
      13617: inst = 32'hc404d6f;
      13618: inst = 32'h8220000;
      13619: inst = 32'h10408000;
      13620: inst = 32'hc404d70;
      13621: inst = 32'h8220000;
      13622: inst = 32'h10408000;
      13623: inst = 32'hc404d71;
      13624: inst = 32'h8220000;
      13625: inst = 32'h10408000;
      13626: inst = 32'hc404d72;
      13627: inst = 32'h8220000;
      13628: inst = 32'h10408000;
      13629: inst = 32'hc404d73;
      13630: inst = 32'h8220000;
      13631: inst = 32'h10408000;
      13632: inst = 32'hc404d74;
      13633: inst = 32'h8220000;
      13634: inst = 32'h10408000;
      13635: inst = 32'hc404dc0;
      13636: inst = 32'h8220000;
      13637: inst = 32'h10408000;
      13638: inst = 32'hc404dca;
      13639: inst = 32'h8220000;
      13640: inst = 32'h10408000;
      13641: inst = 32'hc404dd4;
      13642: inst = 32'h8220000;
      13643: inst = 32'h10408000;
      13644: inst = 32'hc404e20;
      13645: inst = 32'h8220000;
      13646: inst = 32'h10408000;
      13647: inst = 32'hc404e2a;
      13648: inst = 32'h8220000;
      13649: inst = 32'h10408000;
      13650: inst = 32'hc404e34;
      13651: inst = 32'h8220000;
      13652: inst = 32'h10408000;
      13653: inst = 32'hc404e80;
      13654: inst = 32'h8220000;
      13655: inst = 32'h10408000;
      13656: inst = 32'hc404e8a;
      13657: inst = 32'h8220000;
      13658: inst = 32'h10408000;
      13659: inst = 32'hc404e94;
      13660: inst = 32'h8220000;
      13661: inst = 32'h10408000;
      13662: inst = 32'hc404ee0;
      13663: inst = 32'h8220000;
      13664: inst = 32'h10408000;
      13665: inst = 32'hc404eea;
      13666: inst = 32'h8220000;
      13667: inst = 32'h10408000;
      13668: inst = 32'hc404ef4;
      13669: inst = 32'h8220000;
      13670: inst = 32'h10408000;
      13671: inst = 32'hc404f40;
      13672: inst = 32'h8220000;
      13673: inst = 32'h10408000;
      13674: inst = 32'hc404f4a;
      13675: inst = 32'h8220000;
      13676: inst = 32'h10408000;
      13677: inst = 32'hc404f54;
      13678: inst = 32'h8220000;
      13679: inst = 32'h10408000;
      13680: inst = 32'hc404fa0;
      13681: inst = 32'h8220000;
      13682: inst = 32'h10408000;
      13683: inst = 32'hc404faa;
      13684: inst = 32'h8220000;
      13685: inst = 32'h10408000;
      13686: inst = 32'hc404fb4;
      13687: inst = 32'h8220000;
      13688: inst = 32'h10408000;
      13689: inst = 32'hc405000;
      13690: inst = 32'h8220000;
      13691: inst = 32'h10408000;
      13692: inst = 32'hc40500a;
      13693: inst = 32'h8220000;
      13694: inst = 32'h10408000;
      13695: inst = 32'hc405014;
      13696: inst = 32'h8220000;
      13697: inst = 32'h10408000;
      13698: inst = 32'hc405060;
      13699: inst = 32'h8220000;
      13700: inst = 32'h10408000;
      13701: inst = 32'hc40506a;
      13702: inst = 32'h8220000;
      13703: inst = 32'h10408000;
      13704: inst = 32'hc405074;
      13705: inst = 32'h8220000;
      13706: inst = 32'h10408000;
      13707: inst = 32'hc4050c0;
      13708: inst = 32'h8220000;
      13709: inst = 32'h10408000;
      13710: inst = 32'hc4050ca;
      13711: inst = 32'h8220000;
      13712: inst = 32'h10408000;
      13713: inst = 32'hc4050d4;
      13714: inst = 32'h8220000;
      13715: inst = 32'h10408000;
      13716: inst = 32'hc405120;
      13717: inst = 32'h8220000;
      13718: inst = 32'h10408000;
      13719: inst = 32'hc40512a;
      13720: inst = 32'h8220000;
      13721: inst = 32'h10408000;
      13722: inst = 32'hc405134;
      13723: inst = 32'h8220000;
      13724: inst = 32'h10408000;
      13725: inst = 32'hc405180;
      13726: inst = 32'h8220000;
      13727: inst = 32'h10408000;
      13728: inst = 32'hc40518a;
      13729: inst = 32'h8220000;
      13730: inst = 32'h10408000;
      13731: inst = 32'hc405194;
      13732: inst = 32'h8220000;
      13733: inst = 32'h10408000;
      13734: inst = 32'hc4051a8;
      13735: inst = 32'h8220000;
      13736: inst = 32'h10408000;
      13737: inst = 32'hc4051a9;
      13738: inst = 32'h8220000;
      13739: inst = 32'h10408000;
      13740: inst = 32'hc4051b7;
      13741: inst = 32'h8220000;
      13742: inst = 32'h10408000;
      13743: inst = 32'hc4051e0;
      13744: inst = 32'h8220000;
      13745: inst = 32'h10408000;
      13746: inst = 32'hc4051ea;
      13747: inst = 32'h8220000;
      13748: inst = 32'h10408000;
      13749: inst = 32'hc4051f4;
      13750: inst = 32'h8220000;
      13751: inst = 32'h10408000;
      13752: inst = 32'hc405208;
      13753: inst = 32'h8220000;
      13754: inst = 32'h10408000;
      13755: inst = 32'hc405217;
      13756: inst = 32'h8220000;
      13757: inst = 32'h10408000;
      13758: inst = 32'hc405240;
      13759: inst = 32'h8220000;
      13760: inst = 32'h10408000;
      13761: inst = 32'hc40524a;
      13762: inst = 32'h8220000;
      13763: inst = 32'h10408000;
      13764: inst = 32'hc405254;
      13765: inst = 32'h8220000;
      13766: inst = 32'h10408000;
      13767: inst = 32'hc40525e;
      13768: inst = 32'h8220000;
      13769: inst = 32'h10408000;
      13770: inst = 32'hc405268;
      13771: inst = 32'h8220000;
      13772: inst = 32'h10408000;
      13773: inst = 32'hc405277;
      13774: inst = 32'h8220000;
      13775: inst = 32'h10408000;
      13776: inst = 32'hc405281;
      13777: inst = 32'h8220000;
      13778: inst = 32'h10408000;
      13779: inst = 32'hc4052a0;
      13780: inst = 32'h8220000;
      13781: inst = 32'h10408000;
      13782: inst = 32'hc4052a1;
      13783: inst = 32'h8220000;
      13784: inst = 32'h10408000;
      13785: inst = 32'hc4052a2;
      13786: inst = 32'h8220000;
      13787: inst = 32'h10408000;
      13788: inst = 32'hc4052a3;
      13789: inst = 32'h8220000;
      13790: inst = 32'h10408000;
      13791: inst = 32'hc4052a4;
      13792: inst = 32'h8220000;
      13793: inst = 32'h10408000;
      13794: inst = 32'hc4052a5;
      13795: inst = 32'h8220000;
      13796: inst = 32'h10408000;
      13797: inst = 32'hc4052a6;
      13798: inst = 32'h8220000;
      13799: inst = 32'h10408000;
      13800: inst = 32'hc4052a7;
      13801: inst = 32'h8220000;
      13802: inst = 32'h10408000;
      13803: inst = 32'hc4052a8;
      13804: inst = 32'h8220000;
      13805: inst = 32'h10408000;
      13806: inst = 32'hc4052a9;
      13807: inst = 32'h8220000;
      13808: inst = 32'h10408000;
      13809: inst = 32'hc4052aa;
      13810: inst = 32'h8220000;
      13811: inst = 32'h10408000;
      13812: inst = 32'hc4052ab;
      13813: inst = 32'h8220000;
      13814: inst = 32'h10408000;
      13815: inst = 32'hc4052ac;
      13816: inst = 32'h8220000;
      13817: inst = 32'h10408000;
      13818: inst = 32'hc4052ad;
      13819: inst = 32'h8220000;
      13820: inst = 32'h10408000;
      13821: inst = 32'hc4052ae;
      13822: inst = 32'h8220000;
      13823: inst = 32'h10408000;
      13824: inst = 32'hc4052af;
      13825: inst = 32'h8220000;
      13826: inst = 32'h10408000;
      13827: inst = 32'hc4052b0;
      13828: inst = 32'h8220000;
      13829: inst = 32'h10408000;
      13830: inst = 32'hc4052b1;
      13831: inst = 32'h8220000;
      13832: inst = 32'h10408000;
      13833: inst = 32'hc4052b2;
      13834: inst = 32'h8220000;
      13835: inst = 32'h10408000;
      13836: inst = 32'hc4052b3;
      13837: inst = 32'h8220000;
      13838: inst = 32'h10408000;
      13839: inst = 32'hc4052b4;
      13840: inst = 32'h8220000;
      13841: inst = 32'h10408000;
      13842: inst = 32'hc4052bd;
      13843: inst = 32'h8220000;
      13844: inst = 32'h10408000;
      13845: inst = 32'hc4052be;
      13846: inst = 32'h8220000;
      13847: inst = 32'h10408000;
      13848: inst = 32'hc4052c8;
      13849: inst = 32'h8220000;
      13850: inst = 32'h10408000;
      13851: inst = 32'hc4052d7;
      13852: inst = 32'h8220000;
      13853: inst = 32'h10408000;
      13854: inst = 32'hc4052e1;
      13855: inst = 32'h8220000;
      13856: inst = 32'h10408000;
      13857: inst = 32'hc4052e2;
      13858: inst = 32'h8220000;
      13859: inst = 32'h10408000;
      13860: inst = 32'hc40531c;
      13861: inst = 32'h8220000;
      13862: inst = 32'h10408000;
      13863: inst = 32'hc40531d;
      13864: inst = 32'h8220000;
      13865: inst = 32'h10408000;
      13866: inst = 32'hc40531e;
      13867: inst = 32'h8220000;
      13868: inst = 32'h10408000;
      13869: inst = 32'hc40531f;
      13870: inst = 32'h8220000;
      13871: inst = 32'h10408000;
      13872: inst = 32'hc405320;
      13873: inst = 32'h8220000;
      13874: inst = 32'h10408000;
      13875: inst = 32'hc405326;
      13876: inst = 32'h8220000;
      13877: inst = 32'h10408000;
      13878: inst = 32'hc405327;
      13879: inst = 32'h8220000;
      13880: inst = 32'h10408000;
      13881: inst = 32'hc405328;
      13882: inst = 32'h8220000;
      13883: inst = 32'h10408000;
      13884: inst = 32'hc405337;
      13885: inst = 32'h8220000;
      13886: inst = 32'h10408000;
      13887: inst = 32'hc405338;
      13888: inst = 32'h8220000;
      13889: inst = 32'h10408000;
      13890: inst = 32'hc405339;
      13891: inst = 32'h8220000;
      13892: inst = 32'h10408000;
      13893: inst = 32'hc40533f;
      13894: inst = 32'h8220000;
      13895: inst = 32'h10408000;
      13896: inst = 32'hc405340;
      13897: inst = 32'h8220000;
      13898: inst = 32'h10408000;
      13899: inst = 32'hc405341;
      13900: inst = 32'h8220000;
      13901: inst = 32'h10408000;
      13902: inst = 32'hc405342;
      13903: inst = 32'h8220000;
      13904: inst = 32'h10408000;
      13905: inst = 32'hc405343;
      13906: inst = 32'h8220000;
      13907: inst = 32'h10408000;
      13908: inst = 32'hc40537b;
      13909: inst = 32'h8220000;
      13910: inst = 32'h10408000;
      13911: inst = 32'hc40537c;
      13912: inst = 32'h8220000;
      13913: inst = 32'h10408000;
      13914: inst = 32'hc405386;
      13915: inst = 32'h8220000;
      13916: inst = 32'h10408000;
      13917: inst = 32'hc405387;
      13918: inst = 32'h8220000;
      13919: inst = 32'h10408000;
      13920: inst = 32'hc405388;
      13921: inst = 32'h8220000;
      13922: inst = 32'h10408000;
      13923: inst = 32'hc405397;
      13924: inst = 32'h8220000;
      13925: inst = 32'h10408000;
      13926: inst = 32'hc405398;
      13927: inst = 32'h8220000;
      13928: inst = 32'h10408000;
      13929: inst = 32'hc405399;
      13930: inst = 32'h8220000;
      13931: inst = 32'h10408000;
      13932: inst = 32'hc4053a3;
      13933: inst = 32'h8220000;
      13934: inst = 32'h10408000;
      13935: inst = 32'hc4053a4;
      13936: inst = 32'h8220000;
      13937: inst = 32'h10408000;
      13938: inst = 32'hc4053db;
      13939: inst = 32'h8220000;
      13940: inst = 32'h10408000;
      13941: inst = 32'hc4053e5;
      13942: inst = 32'h8220000;
      13943: inst = 32'h10408000;
      13944: inst = 32'hc4053e6;
      13945: inst = 32'h8220000;
      13946: inst = 32'h10408000;
      13947: inst = 32'hc4053e7;
      13948: inst = 32'h8220000;
      13949: inst = 32'h10408000;
      13950: inst = 32'hc4053f8;
      13951: inst = 32'h8220000;
      13952: inst = 32'h10408000;
      13953: inst = 32'hc4053f9;
      13954: inst = 32'h8220000;
      13955: inst = 32'h10408000;
      13956: inst = 32'hc4053fa;
      13957: inst = 32'h8220000;
      13958: inst = 32'h10408000;
      13959: inst = 32'hc405404;
      13960: inst = 32'h8220000;
      13961: inst = 32'h10408000;
      13962: inst = 32'hc40543a;
      13963: inst = 32'h8220000;
      13964: inst = 32'h10408000;
      13965: inst = 32'hc40543b;
      13966: inst = 32'h8220000;
      13967: inst = 32'h10408000;
      13968: inst = 32'hc405445;
      13969: inst = 32'h8220000;
      13970: inst = 32'h10408000;
      13971: inst = 32'hc405446;
      13972: inst = 32'h8220000;
      13973: inst = 32'h10408000;
      13974: inst = 32'hc405447;
      13975: inst = 32'h8220000;
      13976: inst = 32'h10408000;
      13977: inst = 32'hc405458;
      13978: inst = 32'h8220000;
      13979: inst = 32'h10408000;
      13980: inst = 32'hc405459;
      13981: inst = 32'h8220000;
      13982: inst = 32'h10408000;
      13983: inst = 32'hc40545a;
      13984: inst = 32'h8220000;
      13985: inst = 32'h10408000;
      13986: inst = 32'hc405464;
      13987: inst = 32'h8220000;
      13988: inst = 32'h10408000;
      13989: inst = 32'hc405465;
      13990: inst = 32'h8220000;
      13991: inst = 32'h10408000;
      13992: inst = 32'hc405499;
      13993: inst = 32'h8220000;
      13994: inst = 32'h10408000;
      13995: inst = 32'hc40549a;
      13996: inst = 32'h8220000;
      13997: inst = 32'h10408000;
      13998: inst = 32'hc4054a5;
      13999: inst = 32'h8220000;
      14000: inst = 32'h10408000;
      14001: inst = 32'hc4054a6;
      14002: inst = 32'h8220000;
      14003: inst = 32'h10408000;
      14004: inst = 32'hc4054a7;
      14005: inst = 32'h8220000;
      14006: inst = 32'h10408000;
      14007: inst = 32'hc4054b8;
      14008: inst = 32'h8220000;
      14009: inst = 32'h10408000;
      14010: inst = 32'hc4054b9;
      14011: inst = 32'h8220000;
      14012: inst = 32'h10408000;
      14013: inst = 32'hc4054ba;
      14014: inst = 32'h8220000;
      14015: inst = 32'h10408000;
      14016: inst = 32'hc4054c5;
      14017: inst = 32'h8220000;
      14018: inst = 32'h10408000;
      14019: inst = 32'hc4054c6;
      14020: inst = 32'h8220000;
      14021: inst = 32'h10408000;
      14022: inst = 32'hc4054f8;
      14023: inst = 32'h8220000;
      14024: inst = 32'h10408000;
      14025: inst = 32'hc4054f9;
      14026: inst = 32'h8220000;
      14027: inst = 32'h10408000;
      14028: inst = 32'hc405500;
      14029: inst = 32'h8220000;
      14030: inst = 32'h10408000;
      14031: inst = 32'hc405504;
      14032: inst = 32'h8220000;
      14033: inst = 32'h10408000;
      14034: inst = 32'hc405505;
      14035: inst = 32'h8220000;
      14036: inst = 32'h10408000;
      14037: inst = 32'hc405506;
      14038: inst = 32'h8220000;
      14039: inst = 32'h10408000;
      14040: inst = 32'hc405507;
      14041: inst = 32'h8220000;
      14042: inst = 32'h10408000;
      14043: inst = 32'hc405518;
      14044: inst = 32'h8220000;
      14045: inst = 32'h10408000;
      14046: inst = 32'hc405519;
      14047: inst = 32'h8220000;
      14048: inst = 32'h10408000;
      14049: inst = 32'hc40551a;
      14050: inst = 32'h8220000;
      14051: inst = 32'h10408000;
      14052: inst = 32'hc40551b;
      14053: inst = 32'h8220000;
      14054: inst = 32'h10408000;
      14055: inst = 32'hc40551f;
      14056: inst = 32'h8220000;
      14057: inst = 32'h10408000;
      14058: inst = 32'hc405526;
      14059: inst = 32'h8220000;
      14060: inst = 32'h10408000;
      14061: inst = 32'hc405527;
      14062: inst = 32'h8220000;
      14063: inst = 32'h10408000;
      14064: inst = 32'hc405558;
      14065: inst = 32'h8220000;
      14066: inst = 32'h10408000;
      14067: inst = 32'hc405559;
      14068: inst = 32'h8220000;
      14069: inst = 32'h10408000;
      14070: inst = 32'hc405560;
      14071: inst = 32'h8220000;
      14072: inst = 32'h10408000;
      14073: inst = 32'hc405564;
      14074: inst = 32'h8220000;
      14075: inst = 32'h10408000;
      14076: inst = 32'hc405565;
      14077: inst = 32'h8220000;
      14078: inst = 32'h10408000;
      14079: inst = 32'hc405566;
      14080: inst = 32'h8220000;
      14081: inst = 32'h10408000;
      14082: inst = 32'hc405567;
      14083: inst = 32'h8220000;
      14084: inst = 32'h10408000;
      14085: inst = 32'hc405578;
      14086: inst = 32'h8220000;
      14087: inst = 32'h10408000;
      14088: inst = 32'hc405579;
      14089: inst = 32'h8220000;
      14090: inst = 32'h10408000;
      14091: inst = 32'hc40557a;
      14092: inst = 32'h8220000;
      14093: inst = 32'h10408000;
      14094: inst = 32'hc40557b;
      14095: inst = 32'h8220000;
      14096: inst = 32'h10408000;
      14097: inst = 32'hc40557f;
      14098: inst = 32'h8220000;
      14099: inst = 32'h10408000;
      14100: inst = 32'hc405586;
      14101: inst = 32'h8220000;
      14102: inst = 32'h10408000;
      14103: inst = 32'hc405587;
      14104: inst = 32'h8220000;
      14105: inst = 32'h10408000;
      14106: inst = 32'hc4055b7;
      14107: inst = 32'h8220000;
      14108: inst = 32'h10408000;
      14109: inst = 32'hc4055b8;
      14110: inst = 32'h8220000;
      14111: inst = 32'h10408000;
      14112: inst = 32'hc4055bf;
      14113: inst = 32'h8220000;
      14114: inst = 32'h10408000;
      14115: inst = 32'hc4055c0;
      14116: inst = 32'h8220000;
      14117: inst = 32'h10408000;
      14118: inst = 32'hc4055c4;
      14119: inst = 32'h8220000;
      14120: inst = 32'h10408000;
      14121: inst = 32'hc4055c5;
      14122: inst = 32'h8220000;
      14123: inst = 32'h10408000;
      14124: inst = 32'hc4055c6;
      14125: inst = 32'h8220000;
      14126: inst = 32'h10408000;
      14127: inst = 32'hc4055c7;
      14128: inst = 32'h8220000;
      14129: inst = 32'h10408000;
      14130: inst = 32'hc4055d8;
      14131: inst = 32'h8220000;
      14132: inst = 32'h10408000;
      14133: inst = 32'hc4055d9;
      14134: inst = 32'h8220000;
      14135: inst = 32'h10408000;
      14136: inst = 32'hc4055da;
      14137: inst = 32'h8220000;
      14138: inst = 32'h10408000;
      14139: inst = 32'hc4055db;
      14140: inst = 32'h8220000;
      14141: inst = 32'h10408000;
      14142: inst = 32'hc4055df;
      14143: inst = 32'h8220000;
      14144: inst = 32'h10408000;
      14145: inst = 32'hc4055e0;
      14146: inst = 32'h8220000;
      14147: inst = 32'h10408000;
      14148: inst = 32'hc4055e7;
      14149: inst = 32'h8220000;
      14150: inst = 32'h10408000;
      14151: inst = 32'hc4055e8;
      14152: inst = 32'h8220000;
      14153: inst = 32'h10408000;
      14154: inst = 32'hc405616;
      14155: inst = 32'h8220000;
      14156: inst = 32'h10408000;
      14157: inst = 32'hc405617;
      14158: inst = 32'h8220000;
      14159: inst = 32'h10408000;
      14160: inst = 32'hc40561f;
      14161: inst = 32'h8220000;
      14162: inst = 32'h10408000;
      14163: inst = 32'hc405620;
      14164: inst = 32'h8220000;
      14165: inst = 32'h10408000;
      14166: inst = 32'hc405623;
      14167: inst = 32'h8220000;
      14168: inst = 32'h10408000;
      14169: inst = 32'hc405624;
      14170: inst = 32'h8220000;
      14171: inst = 32'h10408000;
      14172: inst = 32'hc405625;
      14173: inst = 32'h8220000;
      14174: inst = 32'h10408000;
      14175: inst = 32'hc405626;
      14176: inst = 32'h8220000;
      14177: inst = 32'h10408000;
      14178: inst = 32'hc405639;
      14179: inst = 32'h8220000;
      14180: inst = 32'h10408000;
      14181: inst = 32'hc40563a;
      14182: inst = 32'h8220000;
      14183: inst = 32'h10408000;
      14184: inst = 32'hc40563b;
      14185: inst = 32'h8220000;
      14186: inst = 32'h10408000;
      14187: inst = 32'hc40563c;
      14188: inst = 32'h8220000;
      14189: inst = 32'h10408000;
      14190: inst = 32'hc40563f;
      14191: inst = 32'h8220000;
      14192: inst = 32'h10408000;
      14193: inst = 32'hc405640;
      14194: inst = 32'h8220000;
      14195: inst = 32'h10408000;
      14196: inst = 32'hc405648;
      14197: inst = 32'h8220000;
      14198: inst = 32'h10408000;
      14199: inst = 32'hc405649;
      14200: inst = 32'h8220000;
      14201: inst = 32'h10408000;
      14202: inst = 32'hc405675;
      14203: inst = 32'h8220000;
      14204: inst = 32'h10408000;
      14205: inst = 32'hc405676;
      14206: inst = 32'h8220000;
      14207: inst = 32'h10408000;
      14208: inst = 32'hc405677;
      14209: inst = 32'h8220000;
      14210: inst = 32'h10408000;
      14211: inst = 32'hc40567e;
      14212: inst = 32'h8220000;
      14213: inst = 32'h10408000;
      14214: inst = 32'hc40567f;
      14215: inst = 32'h8220000;
      14216: inst = 32'h10408000;
      14217: inst = 32'hc405680;
      14218: inst = 32'h8220000;
      14219: inst = 32'h10408000;
      14220: inst = 32'hc405683;
      14221: inst = 32'h8220000;
      14222: inst = 32'h10408000;
      14223: inst = 32'hc405684;
      14224: inst = 32'h8220000;
      14225: inst = 32'h10408000;
      14226: inst = 32'hc405685;
      14227: inst = 32'h8220000;
      14228: inst = 32'h10408000;
      14229: inst = 32'hc405686;
      14230: inst = 32'h8220000;
      14231: inst = 32'h10408000;
      14232: inst = 32'hc405699;
      14233: inst = 32'h8220000;
      14234: inst = 32'h10408000;
      14235: inst = 32'hc40569a;
      14236: inst = 32'h8220000;
      14237: inst = 32'h10408000;
      14238: inst = 32'hc40569b;
      14239: inst = 32'h8220000;
      14240: inst = 32'h10408000;
      14241: inst = 32'hc40569c;
      14242: inst = 32'h8220000;
      14243: inst = 32'h10408000;
      14244: inst = 32'hc40569f;
      14245: inst = 32'h8220000;
      14246: inst = 32'h10408000;
      14247: inst = 32'hc4056a0;
      14248: inst = 32'h8220000;
      14249: inst = 32'h10408000;
      14250: inst = 32'hc4056a1;
      14251: inst = 32'h8220000;
      14252: inst = 32'h10408000;
      14253: inst = 32'hc4056a8;
      14254: inst = 32'h8220000;
      14255: inst = 32'h10408000;
      14256: inst = 32'hc4056a9;
      14257: inst = 32'h8220000;
      14258: inst = 32'h10408000;
      14259: inst = 32'hc4056aa;
      14260: inst = 32'h8220000;
      14261: inst = 32'h10408000;
      14262: inst = 32'hc4056d4;
      14263: inst = 32'h8220000;
      14264: inst = 32'h10408000;
      14265: inst = 32'hc4056d5;
      14266: inst = 32'h8220000;
      14267: inst = 32'h10408000;
      14268: inst = 32'hc4056d6;
      14269: inst = 32'h8220000;
      14270: inst = 32'h10408000;
      14271: inst = 32'hc4056d7;
      14272: inst = 32'h8220000;
      14273: inst = 32'h10408000;
      14274: inst = 32'hc4056d8;
      14275: inst = 32'h8220000;
      14276: inst = 32'h10408000;
      14277: inst = 32'hc4056d9;
      14278: inst = 32'h8220000;
      14279: inst = 32'h10408000;
      14280: inst = 32'hc4056da;
      14281: inst = 32'h8220000;
      14282: inst = 32'h10408000;
      14283: inst = 32'hc4056db;
      14284: inst = 32'h8220000;
      14285: inst = 32'h10408000;
      14286: inst = 32'hc4056dc;
      14287: inst = 32'h8220000;
      14288: inst = 32'h10408000;
      14289: inst = 32'hc4056dd;
      14290: inst = 32'h8220000;
      14291: inst = 32'h10408000;
      14292: inst = 32'hc4056de;
      14293: inst = 32'h8220000;
      14294: inst = 32'h10408000;
      14295: inst = 32'hc4056df;
      14296: inst = 32'h8220000;
      14297: inst = 32'h10408000;
      14298: inst = 32'hc4056e0;
      14299: inst = 32'h8220000;
      14300: inst = 32'h10408000;
      14301: inst = 32'hc4056e3;
      14302: inst = 32'h8220000;
      14303: inst = 32'h10408000;
      14304: inst = 32'hc4056e4;
      14305: inst = 32'h8220000;
      14306: inst = 32'h10408000;
      14307: inst = 32'hc4056e5;
      14308: inst = 32'h8220000;
      14309: inst = 32'h10408000;
      14310: inst = 32'hc4056e6;
      14311: inst = 32'h8220000;
      14312: inst = 32'h10408000;
      14313: inst = 32'hc4056f9;
      14314: inst = 32'h8220000;
      14315: inst = 32'h10408000;
      14316: inst = 32'hc4056fa;
      14317: inst = 32'h8220000;
      14318: inst = 32'h10408000;
      14319: inst = 32'hc4056fb;
      14320: inst = 32'h8220000;
      14321: inst = 32'h10408000;
      14322: inst = 32'hc4056fc;
      14323: inst = 32'h8220000;
      14324: inst = 32'h10408000;
      14325: inst = 32'hc4056ff;
      14326: inst = 32'h8220000;
      14327: inst = 32'h10408000;
      14328: inst = 32'hc405700;
      14329: inst = 32'h8220000;
      14330: inst = 32'h10408000;
      14331: inst = 32'hc405701;
      14332: inst = 32'h8220000;
      14333: inst = 32'h10408000;
      14334: inst = 32'hc405702;
      14335: inst = 32'h8220000;
      14336: inst = 32'h10408000;
      14337: inst = 32'hc405703;
      14338: inst = 32'h8220000;
      14339: inst = 32'h10408000;
      14340: inst = 32'hc405704;
      14341: inst = 32'h8220000;
      14342: inst = 32'h10408000;
      14343: inst = 32'hc405705;
      14344: inst = 32'h8220000;
      14345: inst = 32'h10408000;
      14346: inst = 32'hc405706;
      14347: inst = 32'h8220000;
      14348: inst = 32'h10408000;
      14349: inst = 32'hc405707;
      14350: inst = 32'h8220000;
      14351: inst = 32'h10408000;
      14352: inst = 32'hc405708;
      14353: inst = 32'h8220000;
      14354: inst = 32'h10408000;
      14355: inst = 32'hc405709;
      14356: inst = 32'h8220000;
      14357: inst = 32'h10408000;
      14358: inst = 32'hc40570a;
      14359: inst = 32'h8220000;
      14360: inst = 32'h10408000;
      14361: inst = 32'hc405734;
      14362: inst = 32'h8220000;
      14363: inst = 32'h10408000;
      14364: inst = 32'hc405735;
      14365: inst = 32'h8220000;
      14366: inst = 32'h10408000;
      14367: inst = 32'hc405736;
      14368: inst = 32'h8220000;
      14369: inst = 32'h10408000;
      14370: inst = 32'hc405737;
      14371: inst = 32'h8220000;
      14372: inst = 32'h10408000;
      14373: inst = 32'hc405738;
      14374: inst = 32'h8220000;
      14375: inst = 32'h10408000;
      14376: inst = 32'hc405739;
      14377: inst = 32'h8220000;
      14378: inst = 32'h10408000;
      14379: inst = 32'hc40573a;
      14380: inst = 32'h8220000;
      14381: inst = 32'h10408000;
      14382: inst = 32'hc40573b;
      14383: inst = 32'h8220000;
      14384: inst = 32'h10408000;
      14385: inst = 32'hc40573c;
      14386: inst = 32'h8220000;
      14387: inst = 32'h10408000;
      14388: inst = 32'hc40573d;
      14389: inst = 32'h8220000;
      14390: inst = 32'h10408000;
      14391: inst = 32'hc40573e;
      14392: inst = 32'h8220000;
      14393: inst = 32'h10408000;
      14394: inst = 32'hc40573f;
      14395: inst = 32'h8220000;
      14396: inst = 32'h10408000;
      14397: inst = 32'hc405740;
      14398: inst = 32'h8220000;
      14399: inst = 32'h10408000;
      14400: inst = 32'hc405742;
      14401: inst = 32'h8220000;
      14402: inst = 32'h10408000;
      14403: inst = 32'hc405743;
      14404: inst = 32'h8220000;
      14405: inst = 32'h10408000;
      14406: inst = 32'hc405744;
      14407: inst = 32'h8220000;
      14408: inst = 32'h10408000;
      14409: inst = 32'hc405745;
      14410: inst = 32'h8220000;
      14411: inst = 32'h10408000;
      14412: inst = 32'hc405746;
      14413: inst = 32'h8220000;
      14414: inst = 32'h10408000;
      14415: inst = 32'hc405759;
      14416: inst = 32'h8220000;
      14417: inst = 32'h10408000;
      14418: inst = 32'hc40575a;
      14419: inst = 32'h8220000;
      14420: inst = 32'h10408000;
      14421: inst = 32'hc40575b;
      14422: inst = 32'h8220000;
      14423: inst = 32'h10408000;
      14424: inst = 32'hc40575c;
      14425: inst = 32'h8220000;
      14426: inst = 32'h10408000;
      14427: inst = 32'hc40575d;
      14428: inst = 32'h8220000;
      14429: inst = 32'h10408000;
      14430: inst = 32'hc40575f;
      14431: inst = 32'h8220000;
      14432: inst = 32'h10408000;
      14433: inst = 32'hc405760;
      14434: inst = 32'h8220000;
      14435: inst = 32'h10408000;
      14436: inst = 32'hc405761;
      14437: inst = 32'h8220000;
      14438: inst = 32'h10408000;
      14439: inst = 32'hc405762;
      14440: inst = 32'h8220000;
      14441: inst = 32'h10408000;
      14442: inst = 32'hc405763;
      14443: inst = 32'h8220000;
      14444: inst = 32'h10408000;
      14445: inst = 32'hc405764;
      14446: inst = 32'h8220000;
      14447: inst = 32'h10408000;
      14448: inst = 32'hc405765;
      14449: inst = 32'h8220000;
      14450: inst = 32'h10408000;
      14451: inst = 32'hc405766;
      14452: inst = 32'h8220000;
      14453: inst = 32'h10408000;
      14454: inst = 32'hc405767;
      14455: inst = 32'h8220000;
      14456: inst = 32'h10408000;
      14457: inst = 32'hc405768;
      14458: inst = 32'h8220000;
      14459: inst = 32'h10408000;
      14460: inst = 32'hc405769;
      14461: inst = 32'h8220000;
      14462: inst = 32'h10408000;
      14463: inst = 32'hc40576a;
      14464: inst = 32'h8220000;
      14465: inst = 32'h10408000;
      14466: inst = 32'hc40576b;
      14467: inst = 32'h8220000;
      14468: inst = 32'h10408000;
      14469: inst = 32'hc405793;
      14470: inst = 32'h8220000;
      14471: inst = 32'h10408000;
      14472: inst = 32'hc405794;
      14473: inst = 32'h8220000;
      14474: inst = 32'h10408000;
      14475: inst = 32'hc405795;
      14476: inst = 32'h8220000;
      14477: inst = 32'h10408000;
      14478: inst = 32'hc405796;
      14479: inst = 32'h8220000;
      14480: inst = 32'h10408000;
      14481: inst = 32'hc405797;
      14482: inst = 32'h8220000;
      14483: inst = 32'h10408000;
      14484: inst = 32'hc405798;
      14485: inst = 32'h8220000;
      14486: inst = 32'h10408000;
      14487: inst = 32'hc405799;
      14488: inst = 32'h8220000;
      14489: inst = 32'h10408000;
      14490: inst = 32'hc40579a;
      14491: inst = 32'h8220000;
      14492: inst = 32'h10408000;
      14493: inst = 32'hc40579b;
      14494: inst = 32'h8220000;
      14495: inst = 32'h10408000;
      14496: inst = 32'hc40579c;
      14497: inst = 32'h8220000;
      14498: inst = 32'h10408000;
      14499: inst = 32'hc40579d;
      14500: inst = 32'h8220000;
      14501: inst = 32'h10408000;
      14502: inst = 32'hc40579e;
      14503: inst = 32'h8220000;
      14504: inst = 32'h10408000;
      14505: inst = 32'hc40579f;
      14506: inst = 32'h8220000;
      14507: inst = 32'h10408000;
      14508: inst = 32'hc4057a0;
      14509: inst = 32'h8220000;
      14510: inst = 32'h10408000;
      14511: inst = 32'hc4057a1;
      14512: inst = 32'h8220000;
      14513: inst = 32'h10408000;
      14514: inst = 32'hc4057a2;
      14515: inst = 32'h8220000;
      14516: inst = 32'h10408000;
      14517: inst = 32'hc4057a3;
      14518: inst = 32'h8220000;
      14519: inst = 32'h10408000;
      14520: inst = 32'hc4057a4;
      14521: inst = 32'h8220000;
      14522: inst = 32'h10408000;
      14523: inst = 32'hc4057a5;
      14524: inst = 32'h8220000;
      14525: inst = 32'h10408000;
      14526: inst = 32'hc4057a6;
      14527: inst = 32'h8220000;
      14528: inst = 32'h10408000;
      14529: inst = 32'hc4057b9;
      14530: inst = 32'h8220000;
      14531: inst = 32'h10408000;
      14532: inst = 32'hc4057ba;
      14533: inst = 32'h8220000;
      14534: inst = 32'h10408000;
      14535: inst = 32'hc4057bb;
      14536: inst = 32'h8220000;
      14537: inst = 32'h10408000;
      14538: inst = 32'hc4057bc;
      14539: inst = 32'h8220000;
      14540: inst = 32'h10408000;
      14541: inst = 32'hc4057bd;
      14542: inst = 32'h8220000;
      14543: inst = 32'h10408000;
      14544: inst = 32'hc4057be;
      14545: inst = 32'h8220000;
      14546: inst = 32'h10408000;
      14547: inst = 32'hc4057bf;
      14548: inst = 32'h8220000;
      14549: inst = 32'h10408000;
      14550: inst = 32'hc4057c0;
      14551: inst = 32'h8220000;
      14552: inst = 32'h10408000;
      14553: inst = 32'hc4057c1;
      14554: inst = 32'h8220000;
      14555: inst = 32'h10408000;
      14556: inst = 32'hc4057c2;
      14557: inst = 32'h8220000;
      14558: inst = 32'h10408000;
      14559: inst = 32'hc4057c3;
      14560: inst = 32'h8220000;
      14561: inst = 32'h10408000;
      14562: inst = 32'hc4057c4;
      14563: inst = 32'h8220000;
      14564: inst = 32'h10408000;
      14565: inst = 32'hc4057c5;
      14566: inst = 32'h8220000;
      14567: inst = 32'h10408000;
      14568: inst = 32'hc4057c6;
      14569: inst = 32'h8220000;
      14570: inst = 32'h10408000;
      14571: inst = 32'hc4057c7;
      14572: inst = 32'h8220000;
      14573: inst = 32'h10408000;
      14574: inst = 32'hc4057c8;
      14575: inst = 32'h8220000;
      14576: inst = 32'h10408000;
      14577: inst = 32'hc4057c9;
      14578: inst = 32'h8220000;
      14579: inst = 32'h10408000;
      14580: inst = 32'hc4057ca;
      14581: inst = 32'h8220000;
      14582: inst = 32'h10408000;
      14583: inst = 32'hc4057cb;
      14584: inst = 32'h8220000;
      14585: inst = 32'h10408000;
      14586: inst = 32'hc4057cc;
      14587: inst = 32'h8220000;
      14588: inst = 32'hc20bdd7;
      14589: inst = 32'h10408000;
      14590: inst = 32'hc404dc1;
      14591: inst = 32'h8220000;
      14592: inst = 32'h10408000;
      14593: inst = 32'hc404dc2;
      14594: inst = 32'h8220000;
      14595: inst = 32'h10408000;
      14596: inst = 32'hc404dc3;
      14597: inst = 32'h8220000;
      14598: inst = 32'h10408000;
      14599: inst = 32'hc404dc4;
      14600: inst = 32'h8220000;
      14601: inst = 32'h10408000;
      14602: inst = 32'hc404dc5;
      14603: inst = 32'h8220000;
      14604: inst = 32'h10408000;
      14605: inst = 32'hc404dc6;
      14606: inst = 32'h8220000;
      14607: inst = 32'h10408000;
      14608: inst = 32'hc404dc7;
      14609: inst = 32'h8220000;
      14610: inst = 32'h10408000;
      14611: inst = 32'hc404dc8;
      14612: inst = 32'h8220000;
      14613: inst = 32'h10408000;
      14614: inst = 32'hc404dc9;
      14615: inst = 32'h8220000;
      14616: inst = 32'h10408000;
      14617: inst = 32'hc404dcb;
      14618: inst = 32'h8220000;
      14619: inst = 32'h10408000;
      14620: inst = 32'hc404dcc;
      14621: inst = 32'h8220000;
      14622: inst = 32'h10408000;
      14623: inst = 32'hc404dcd;
      14624: inst = 32'h8220000;
      14625: inst = 32'h10408000;
      14626: inst = 32'hc404dce;
      14627: inst = 32'h8220000;
      14628: inst = 32'h10408000;
      14629: inst = 32'hc404dcf;
      14630: inst = 32'h8220000;
      14631: inst = 32'h10408000;
      14632: inst = 32'hc404dd0;
      14633: inst = 32'h8220000;
      14634: inst = 32'h10408000;
      14635: inst = 32'hc404dd1;
      14636: inst = 32'h8220000;
      14637: inst = 32'h10408000;
      14638: inst = 32'hc404dd2;
      14639: inst = 32'h8220000;
      14640: inst = 32'h10408000;
      14641: inst = 32'hc404dd3;
      14642: inst = 32'h8220000;
      14643: inst = 32'h10408000;
      14644: inst = 32'hc404e21;
      14645: inst = 32'h8220000;
      14646: inst = 32'h10408000;
      14647: inst = 32'hc404e22;
      14648: inst = 32'h8220000;
      14649: inst = 32'h10408000;
      14650: inst = 32'hc404e23;
      14651: inst = 32'h8220000;
      14652: inst = 32'h10408000;
      14653: inst = 32'hc404e24;
      14654: inst = 32'h8220000;
      14655: inst = 32'h10408000;
      14656: inst = 32'hc404e25;
      14657: inst = 32'h8220000;
      14658: inst = 32'h10408000;
      14659: inst = 32'hc404e26;
      14660: inst = 32'h8220000;
      14661: inst = 32'h10408000;
      14662: inst = 32'hc404e27;
      14663: inst = 32'h8220000;
      14664: inst = 32'h10408000;
      14665: inst = 32'hc404e28;
      14666: inst = 32'h8220000;
      14667: inst = 32'h10408000;
      14668: inst = 32'hc404e29;
      14669: inst = 32'h8220000;
      14670: inst = 32'h10408000;
      14671: inst = 32'hc404e2b;
      14672: inst = 32'h8220000;
      14673: inst = 32'h10408000;
      14674: inst = 32'hc404e2c;
      14675: inst = 32'h8220000;
      14676: inst = 32'h10408000;
      14677: inst = 32'hc404e2d;
      14678: inst = 32'h8220000;
      14679: inst = 32'h10408000;
      14680: inst = 32'hc404e2e;
      14681: inst = 32'h8220000;
      14682: inst = 32'h10408000;
      14683: inst = 32'hc404e2f;
      14684: inst = 32'h8220000;
      14685: inst = 32'h10408000;
      14686: inst = 32'hc404e30;
      14687: inst = 32'h8220000;
      14688: inst = 32'h10408000;
      14689: inst = 32'hc404e31;
      14690: inst = 32'h8220000;
      14691: inst = 32'h10408000;
      14692: inst = 32'hc404e32;
      14693: inst = 32'h8220000;
      14694: inst = 32'h10408000;
      14695: inst = 32'hc404e33;
      14696: inst = 32'h8220000;
      14697: inst = 32'h10408000;
      14698: inst = 32'hc404e81;
      14699: inst = 32'h8220000;
      14700: inst = 32'h10408000;
      14701: inst = 32'hc404e82;
      14702: inst = 32'h8220000;
      14703: inst = 32'h10408000;
      14704: inst = 32'hc404e83;
      14705: inst = 32'h8220000;
      14706: inst = 32'h10408000;
      14707: inst = 32'hc404e84;
      14708: inst = 32'h8220000;
      14709: inst = 32'h10408000;
      14710: inst = 32'hc404e85;
      14711: inst = 32'h8220000;
      14712: inst = 32'h10408000;
      14713: inst = 32'hc404e86;
      14714: inst = 32'h8220000;
      14715: inst = 32'h10408000;
      14716: inst = 32'hc404e87;
      14717: inst = 32'h8220000;
      14718: inst = 32'h10408000;
      14719: inst = 32'hc404e88;
      14720: inst = 32'h8220000;
      14721: inst = 32'h10408000;
      14722: inst = 32'hc404e89;
      14723: inst = 32'h8220000;
      14724: inst = 32'h10408000;
      14725: inst = 32'hc404e8b;
      14726: inst = 32'h8220000;
      14727: inst = 32'h10408000;
      14728: inst = 32'hc404e8c;
      14729: inst = 32'h8220000;
      14730: inst = 32'h10408000;
      14731: inst = 32'hc404e8d;
      14732: inst = 32'h8220000;
      14733: inst = 32'h10408000;
      14734: inst = 32'hc404e8e;
      14735: inst = 32'h8220000;
      14736: inst = 32'h10408000;
      14737: inst = 32'hc404e8f;
      14738: inst = 32'h8220000;
      14739: inst = 32'h10408000;
      14740: inst = 32'hc404e90;
      14741: inst = 32'h8220000;
      14742: inst = 32'h10408000;
      14743: inst = 32'hc404e91;
      14744: inst = 32'h8220000;
      14745: inst = 32'h10408000;
      14746: inst = 32'hc404e92;
      14747: inst = 32'h8220000;
      14748: inst = 32'h10408000;
      14749: inst = 32'hc404e93;
      14750: inst = 32'h8220000;
      14751: inst = 32'h10408000;
      14752: inst = 32'hc404ee1;
      14753: inst = 32'h8220000;
      14754: inst = 32'h10408000;
      14755: inst = 32'hc404ee2;
      14756: inst = 32'h8220000;
      14757: inst = 32'h10408000;
      14758: inst = 32'hc404ee3;
      14759: inst = 32'h8220000;
      14760: inst = 32'h10408000;
      14761: inst = 32'hc404ee4;
      14762: inst = 32'h8220000;
      14763: inst = 32'h10408000;
      14764: inst = 32'hc404ee5;
      14765: inst = 32'h8220000;
      14766: inst = 32'h10408000;
      14767: inst = 32'hc404ee6;
      14768: inst = 32'h8220000;
      14769: inst = 32'h10408000;
      14770: inst = 32'hc404ee7;
      14771: inst = 32'h8220000;
      14772: inst = 32'h10408000;
      14773: inst = 32'hc404ee8;
      14774: inst = 32'h8220000;
      14775: inst = 32'h10408000;
      14776: inst = 32'hc404ee9;
      14777: inst = 32'h8220000;
      14778: inst = 32'h10408000;
      14779: inst = 32'hc404eeb;
      14780: inst = 32'h8220000;
      14781: inst = 32'h10408000;
      14782: inst = 32'hc404eec;
      14783: inst = 32'h8220000;
      14784: inst = 32'h10408000;
      14785: inst = 32'hc404eed;
      14786: inst = 32'h8220000;
      14787: inst = 32'h10408000;
      14788: inst = 32'hc404eee;
      14789: inst = 32'h8220000;
      14790: inst = 32'h10408000;
      14791: inst = 32'hc404eef;
      14792: inst = 32'h8220000;
      14793: inst = 32'h10408000;
      14794: inst = 32'hc404ef0;
      14795: inst = 32'h8220000;
      14796: inst = 32'h10408000;
      14797: inst = 32'hc404ef1;
      14798: inst = 32'h8220000;
      14799: inst = 32'h10408000;
      14800: inst = 32'hc404ef2;
      14801: inst = 32'h8220000;
      14802: inst = 32'h10408000;
      14803: inst = 32'hc404ef3;
      14804: inst = 32'h8220000;
      14805: inst = 32'h10408000;
      14806: inst = 32'hc404f41;
      14807: inst = 32'h8220000;
      14808: inst = 32'h10408000;
      14809: inst = 32'hc404f42;
      14810: inst = 32'h8220000;
      14811: inst = 32'h10408000;
      14812: inst = 32'hc404f43;
      14813: inst = 32'h8220000;
      14814: inst = 32'h10408000;
      14815: inst = 32'hc404f44;
      14816: inst = 32'h8220000;
      14817: inst = 32'h10408000;
      14818: inst = 32'hc404f45;
      14819: inst = 32'h8220000;
      14820: inst = 32'h10408000;
      14821: inst = 32'hc404f46;
      14822: inst = 32'h8220000;
      14823: inst = 32'h10408000;
      14824: inst = 32'hc404f47;
      14825: inst = 32'h8220000;
      14826: inst = 32'h10408000;
      14827: inst = 32'hc404f48;
      14828: inst = 32'h8220000;
      14829: inst = 32'h10408000;
      14830: inst = 32'hc404f49;
      14831: inst = 32'h8220000;
      14832: inst = 32'h10408000;
      14833: inst = 32'hc404f4b;
      14834: inst = 32'h8220000;
      14835: inst = 32'h10408000;
      14836: inst = 32'hc404f4c;
      14837: inst = 32'h8220000;
      14838: inst = 32'h10408000;
      14839: inst = 32'hc404f4d;
      14840: inst = 32'h8220000;
      14841: inst = 32'h10408000;
      14842: inst = 32'hc404f4e;
      14843: inst = 32'h8220000;
      14844: inst = 32'h10408000;
      14845: inst = 32'hc404f4f;
      14846: inst = 32'h8220000;
      14847: inst = 32'h10408000;
      14848: inst = 32'hc404f50;
      14849: inst = 32'h8220000;
      14850: inst = 32'h10408000;
      14851: inst = 32'hc404f51;
      14852: inst = 32'h8220000;
      14853: inst = 32'h10408000;
      14854: inst = 32'hc404f52;
      14855: inst = 32'h8220000;
      14856: inst = 32'h10408000;
      14857: inst = 32'hc404f53;
      14858: inst = 32'h8220000;
      14859: inst = 32'h10408000;
      14860: inst = 32'hc404fa1;
      14861: inst = 32'h8220000;
      14862: inst = 32'h10408000;
      14863: inst = 32'hc404fa2;
      14864: inst = 32'h8220000;
      14865: inst = 32'h10408000;
      14866: inst = 32'hc404fa3;
      14867: inst = 32'h8220000;
      14868: inst = 32'h10408000;
      14869: inst = 32'hc404fa4;
      14870: inst = 32'h8220000;
      14871: inst = 32'h10408000;
      14872: inst = 32'hc404fa5;
      14873: inst = 32'h8220000;
      14874: inst = 32'h10408000;
      14875: inst = 32'hc404fa6;
      14876: inst = 32'h8220000;
      14877: inst = 32'h10408000;
      14878: inst = 32'hc404fa7;
      14879: inst = 32'h8220000;
      14880: inst = 32'h10408000;
      14881: inst = 32'hc404fa9;
      14882: inst = 32'h8220000;
      14883: inst = 32'h10408000;
      14884: inst = 32'hc404fab;
      14885: inst = 32'h8220000;
      14886: inst = 32'h10408000;
      14887: inst = 32'hc404fad;
      14888: inst = 32'h8220000;
      14889: inst = 32'h10408000;
      14890: inst = 32'hc404fae;
      14891: inst = 32'h8220000;
      14892: inst = 32'h10408000;
      14893: inst = 32'hc404faf;
      14894: inst = 32'h8220000;
      14895: inst = 32'h10408000;
      14896: inst = 32'hc404fb0;
      14897: inst = 32'h8220000;
      14898: inst = 32'h10408000;
      14899: inst = 32'hc404fb1;
      14900: inst = 32'h8220000;
      14901: inst = 32'h10408000;
      14902: inst = 32'hc404fb2;
      14903: inst = 32'h8220000;
      14904: inst = 32'h10408000;
      14905: inst = 32'hc404fb3;
      14906: inst = 32'h8220000;
      14907: inst = 32'h10408000;
      14908: inst = 32'hc405001;
      14909: inst = 32'h8220000;
      14910: inst = 32'h10408000;
      14911: inst = 32'hc405002;
      14912: inst = 32'h8220000;
      14913: inst = 32'h10408000;
      14914: inst = 32'hc405003;
      14915: inst = 32'h8220000;
      14916: inst = 32'h10408000;
      14917: inst = 32'hc405004;
      14918: inst = 32'h8220000;
      14919: inst = 32'h10408000;
      14920: inst = 32'hc405005;
      14921: inst = 32'h8220000;
      14922: inst = 32'h10408000;
      14923: inst = 32'hc405006;
      14924: inst = 32'h8220000;
      14925: inst = 32'h10408000;
      14926: inst = 32'hc405007;
      14927: inst = 32'h8220000;
      14928: inst = 32'h10408000;
      14929: inst = 32'hc405009;
      14930: inst = 32'h8220000;
      14931: inst = 32'h10408000;
      14932: inst = 32'hc40500b;
      14933: inst = 32'h8220000;
      14934: inst = 32'h10408000;
      14935: inst = 32'hc40500d;
      14936: inst = 32'h8220000;
      14937: inst = 32'h10408000;
      14938: inst = 32'hc40500e;
      14939: inst = 32'h8220000;
      14940: inst = 32'h10408000;
      14941: inst = 32'hc40500f;
      14942: inst = 32'h8220000;
      14943: inst = 32'h10408000;
      14944: inst = 32'hc405010;
      14945: inst = 32'h8220000;
      14946: inst = 32'h10408000;
      14947: inst = 32'hc405011;
      14948: inst = 32'h8220000;
      14949: inst = 32'h10408000;
      14950: inst = 32'hc405012;
      14951: inst = 32'h8220000;
      14952: inst = 32'h10408000;
      14953: inst = 32'hc405013;
      14954: inst = 32'h8220000;
      14955: inst = 32'h10408000;
      14956: inst = 32'hc405061;
      14957: inst = 32'h8220000;
      14958: inst = 32'h10408000;
      14959: inst = 32'hc405062;
      14960: inst = 32'h8220000;
      14961: inst = 32'h10408000;
      14962: inst = 32'hc405063;
      14963: inst = 32'h8220000;
      14964: inst = 32'h10408000;
      14965: inst = 32'hc405064;
      14966: inst = 32'h8220000;
      14967: inst = 32'h10408000;
      14968: inst = 32'hc405065;
      14969: inst = 32'h8220000;
      14970: inst = 32'h10408000;
      14971: inst = 32'hc405066;
      14972: inst = 32'h8220000;
      14973: inst = 32'h10408000;
      14974: inst = 32'hc405067;
      14975: inst = 32'h8220000;
      14976: inst = 32'h10408000;
      14977: inst = 32'hc405068;
      14978: inst = 32'h8220000;
      14979: inst = 32'h10408000;
      14980: inst = 32'hc405069;
      14981: inst = 32'h8220000;
      14982: inst = 32'h10408000;
      14983: inst = 32'hc40506b;
      14984: inst = 32'h8220000;
      14985: inst = 32'h10408000;
      14986: inst = 32'hc40506c;
      14987: inst = 32'h8220000;
      14988: inst = 32'h10408000;
      14989: inst = 32'hc40506d;
      14990: inst = 32'h8220000;
      14991: inst = 32'h10408000;
      14992: inst = 32'hc40506e;
      14993: inst = 32'h8220000;
      14994: inst = 32'h10408000;
      14995: inst = 32'hc40506f;
      14996: inst = 32'h8220000;
      14997: inst = 32'h10408000;
      14998: inst = 32'hc405070;
      14999: inst = 32'h8220000;
      15000: inst = 32'h10408000;
      15001: inst = 32'hc405071;
      15002: inst = 32'h8220000;
      15003: inst = 32'h10408000;
      15004: inst = 32'hc405072;
      15005: inst = 32'h8220000;
      15006: inst = 32'h10408000;
      15007: inst = 32'hc405073;
      15008: inst = 32'h8220000;
      15009: inst = 32'h10408000;
      15010: inst = 32'hc4050c1;
      15011: inst = 32'h8220000;
      15012: inst = 32'h10408000;
      15013: inst = 32'hc4050c2;
      15014: inst = 32'h8220000;
      15015: inst = 32'h10408000;
      15016: inst = 32'hc4050c3;
      15017: inst = 32'h8220000;
      15018: inst = 32'h10408000;
      15019: inst = 32'hc4050c4;
      15020: inst = 32'h8220000;
      15021: inst = 32'h10408000;
      15022: inst = 32'hc4050c5;
      15023: inst = 32'h8220000;
      15024: inst = 32'h10408000;
      15025: inst = 32'hc4050c6;
      15026: inst = 32'h8220000;
      15027: inst = 32'h10408000;
      15028: inst = 32'hc4050c7;
      15029: inst = 32'h8220000;
      15030: inst = 32'h10408000;
      15031: inst = 32'hc4050c8;
      15032: inst = 32'h8220000;
      15033: inst = 32'h10408000;
      15034: inst = 32'hc4050c9;
      15035: inst = 32'h8220000;
      15036: inst = 32'h10408000;
      15037: inst = 32'hc4050cb;
      15038: inst = 32'h8220000;
      15039: inst = 32'h10408000;
      15040: inst = 32'hc4050cc;
      15041: inst = 32'h8220000;
      15042: inst = 32'h10408000;
      15043: inst = 32'hc4050cd;
      15044: inst = 32'h8220000;
      15045: inst = 32'h10408000;
      15046: inst = 32'hc4050ce;
      15047: inst = 32'h8220000;
      15048: inst = 32'h10408000;
      15049: inst = 32'hc4050cf;
      15050: inst = 32'h8220000;
      15051: inst = 32'h10408000;
      15052: inst = 32'hc4050d0;
      15053: inst = 32'h8220000;
      15054: inst = 32'h10408000;
      15055: inst = 32'hc4050d1;
      15056: inst = 32'h8220000;
      15057: inst = 32'h10408000;
      15058: inst = 32'hc4050d2;
      15059: inst = 32'h8220000;
      15060: inst = 32'h10408000;
      15061: inst = 32'hc4050d3;
      15062: inst = 32'h8220000;
      15063: inst = 32'h10408000;
      15064: inst = 32'hc405121;
      15065: inst = 32'h8220000;
      15066: inst = 32'h10408000;
      15067: inst = 32'hc405122;
      15068: inst = 32'h8220000;
      15069: inst = 32'h10408000;
      15070: inst = 32'hc405123;
      15071: inst = 32'h8220000;
      15072: inst = 32'h10408000;
      15073: inst = 32'hc405124;
      15074: inst = 32'h8220000;
      15075: inst = 32'h10408000;
      15076: inst = 32'hc405125;
      15077: inst = 32'h8220000;
      15078: inst = 32'h10408000;
      15079: inst = 32'hc405126;
      15080: inst = 32'h8220000;
      15081: inst = 32'h10408000;
      15082: inst = 32'hc405127;
      15083: inst = 32'h8220000;
      15084: inst = 32'h10408000;
      15085: inst = 32'hc405128;
      15086: inst = 32'h8220000;
      15087: inst = 32'h10408000;
      15088: inst = 32'hc405129;
      15089: inst = 32'h8220000;
      15090: inst = 32'h10408000;
      15091: inst = 32'hc40512b;
      15092: inst = 32'h8220000;
      15093: inst = 32'h10408000;
      15094: inst = 32'hc40512c;
      15095: inst = 32'h8220000;
      15096: inst = 32'h10408000;
      15097: inst = 32'hc40512d;
      15098: inst = 32'h8220000;
      15099: inst = 32'h10408000;
      15100: inst = 32'hc40512e;
      15101: inst = 32'h8220000;
      15102: inst = 32'h10408000;
      15103: inst = 32'hc40512f;
      15104: inst = 32'h8220000;
      15105: inst = 32'h10408000;
      15106: inst = 32'hc405130;
      15107: inst = 32'h8220000;
      15108: inst = 32'h10408000;
      15109: inst = 32'hc405131;
      15110: inst = 32'h8220000;
      15111: inst = 32'h10408000;
      15112: inst = 32'hc405132;
      15113: inst = 32'h8220000;
      15114: inst = 32'h10408000;
      15115: inst = 32'hc405133;
      15116: inst = 32'h8220000;
      15117: inst = 32'h10408000;
      15118: inst = 32'hc405181;
      15119: inst = 32'h8220000;
      15120: inst = 32'h10408000;
      15121: inst = 32'hc405182;
      15122: inst = 32'h8220000;
      15123: inst = 32'h10408000;
      15124: inst = 32'hc405183;
      15125: inst = 32'h8220000;
      15126: inst = 32'h10408000;
      15127: inst = 32'hc405184;
      15128: inst = 32'h8220000;
      15129: inst = 32'h10408000;
      15130: inst = 32'hc405185;
      15131: inst = 32'h8220000;
      15132: inst = 32'h10408000;
      15133: inst = 32'hc405186;
      15134: inst = 32'h8220000;
      15135: inst = 32'h10408000;
      15136: inst = 32'hc405187;
      15137: inst = 32'h8220000;
      15138: inst = 32'h10408000;
      15139: inst = 32'hc405188;
      15140: inst = 32'h8220000;
      15141: inst = 32'h10408000;
      15142: inst = 32'hc405189;
      15143: inst = 32'h8220000;
      15144: inst = 32'h10408000;
      15145: inst = 32'hc40518b;
      15146: inst = 32'h8220000;
      15147: inst = 32'h10408000;
      15148: inst = 32'hc40518c;
      15149: inst = 32'h8220000;
      15150: inst = 32'h10408000;
      15151: inst = 32'hc40518d;
      15152: inst = 32'h8220000;
      15153: inst = 32'h10408000;
      15154: inst = 32'hc40518e;
      15155: inst = 32'h8220000;
      15156: inst = 32'h10408000;
      15157: inst = 32'hc40518f;
      15158: inst = 32'h8220000;
      15159: inst = 32'h10408000;
      15160: inst = 32'hc405190;
      15161: inst = 32'h8220000;
      15162: inst = 32'h10408000;
      15163: inst = 32'hc405191;
      15164: inst = 32'h8220000;
      15165: inst = 32'h10408000;
      15166: inst = 32'hc405192;
      15167: inst = 32'h8220000;
      15168: inst = 32'h10408000;
      15169: inst = 32'hc405193;
      15170: inst = 32'h8220000;
      15171: inst = 32'h10408000;
      15172: inst = 32'hc4051e1;
      15173: inst = 32'h8220000;
      15174: inst = 32'h10408000;
      15175: inst = 32'hc4051e2;
      15176: inst = 32'h8220000;
      15177: inst = 32'h10408000;
      15178: inst = 32'hc4051e3;
      15179: inst = 32'h8220000;
      15180: inst = 32'h10408000;
      15181: inst = 32'hc4051e4;
      15182: inst = 32'h8220000;
      15183: inst = 32'h10408000;
      15184: inst = 32'hc4051e5;
      15185: inst = 32'h8220000;
      15186: inst = 32'h10408000;
      15187: inst = 32'hc4051e6;
      15188: inst = 32'h8220000;
      15189: inst = 32'h10408000;
      15190: inst = 32'hc4051e7;
      15191: inst = 32'h8220000;
      15192: inst = 32'h10408000;
      15193: inst = 32'hc4051e8;
      15194: inst = 32'h8220000;
      15195: inst = 32'h10408000;
      15196: inst = 32'hc4051e9;
      15197: inst = 32'h8220000;
      15198: inst = 32'h10408000;
      15199: inst = 32'hc4051eb;
      15200: inst = 32'h8220000;
      15201: inst = 32'h10408000;
      15202: inst = 32'hc4051ec;
      15203: inst = 32'h8220000;
      15204: inst = 32'h10408000;
      15205: inst = 32'hc4051ed;
      15206: inst = 32'h8220000;
      15207: inst = 32'h10408000;
      15208: inst = 32'hc4051ee;
      15209: inst = 32'h8220000;
      15210: inst = 32'h10408000;
      15211: inst = 32'hc4051ef;
      15212: inst = 32'h8220000;
      15213: inst = 32'h10408000;
      15214: inst = 32'hc4051f0;
      15215: inst = 32'h8220000;
      15216: inst = 32'h10408000;
      15217: inst = 32'hc4051f1;
      15218: inst = 32'h8220000;
      15219: inst = 32'h10408000;
      15220: inst = 32'hc4051f2;
      15221: inst = 32'h8220000;
      15222: inst = 32'h10408000;
      15223: inst = 32'hc4051f3;
      15224: inst = 32'h8220000;
      15225: inst = 32'h10408000;
      15226: inst = 32'hc405241;
      15227: inst = 32'h8220000;
      15228: inst = 32'h10408000;
      15229: inst = 32'hc405242;
      15230: inst = 32'h8220000;
      15231: inst = 32'h10408000;
      15232: inst = 32'hc405243;
      15233: inst = 32'h8220000;
      15234: inst = 32'h10408000;
      15235: inst = 32'hc405244;
      15236: inst = 32'h8220000;
      15237: inst = 32'h10408000;
      15238: inst = 32'hc405245;
      15239: inst = 32'h8220000;
      15240: inst = 32'h10408000;
      15241: inst = 32'hc405246;
      15242: inst = 32'h8220000;
      15243: inst = 32'h10408000;
      15244: inst = 32'hc405247;
      15245: inst = 32'h8220000;
      15246: inst = 32'h10408000;
      15247: inst = 32'hc405248;
      15248: inst = 32'h8220000;
      15249: inst = 32'h10408000;
      15250: inst = 32'hc405249;
      15251: inst = 32'h8220000;
      15252: inst = 32'h10408000;
      15253: inst = 32'hc40524b;
      15254: inst = 32'h8220000;
      15255: inst = 32'h10408000;
      15256: inst = 32'hc40524c;
      15257: inst = 32'h8220000;
      15258: inst = 32'h10408000;
      15259: inst = 32'hc40524d;
      15260: inst = 32'h8220000;
      15261: inst = 32'h10408000;
      15262: inst = 32'hc40524e;
      15263: inst = 32'h8220000;
      15264: inst = 32'h10408000;
      15265: inst = 32'hc40524f;
      15266: inst = 32'h8220000;
      15267: inst = 32'h10408000;
      15268: inst = 32'hc405250;
      15269: inst = 32'h8220000;
      15270: inst = 32'h10408000;
      15271: inst = 32'hc405251;
      15272: inst = 32'h8220000;
      15273: inst = 32'h10408000;
      15274: inst = 32'hc405252;
      15275: inst = 32'h8220000;
      15276: inst = 32'h10408000;
      15277: inst = 32'hc405253;
      15278: inst = 32'h8220000;
      15279: inst = 32'hc20bd73;
      15280: inst = 32'h10408000;
      15281: inst = 32'hc404e9f;
      15282: inst = 32'h8220000;
      15283: inst = 32'h10408000;
      15284: inst = 32'hc404ec0;
      15285: inst = 32'h8220000;
      15286: inst = 32'hc205aed;
      15287: inst = 32'h10408000;
      15288: inst = 32'hc404ea0;
      15289: inst = 32'h8220000;
      15290: inst = 32'h10408000;
      15291: inst = 32'hc404ea1;
      15292: inst = 32'h8220000;
      15293: inst = 32'h10408000;
      15294: inst = 32'hc404ea2;
      15295: inst = 32'h8220000;
      15296: inst = 32'h10408000;
      15297: inst = 32'hc404ea3;
      15298: inst = 32'h8220000;
      15299: inst = 32'h10408000;
      15300: inst = 32'hc404ea4;
      15301: inst = 32'h8220000;
      15302: inst = 32'h10408000;
      15303: inst = 32'hc404ebb;
      15304: inst = 32'h8220000;
      15305: inst = 32'h10408000;
      15306: inst = 32'hc404ebc;
      15307: inst = 32'h8220000;
      15308: inst = 32'h10408000;
      15309: inst = 32'hc404ebd;
      15310: inst = 32'h8220000;
      15311: inst = 32'h10408000;
      15312: inst = 32'hc404ebe;
      15313: inst = 32'h8220000;
      15314: inst = 32'h10408000;
      15315: inst = 32'hc404ebf;
      15316: inst = 32'h8220000;
      15317: inst = 32'h10408000;
      15318: inst = 32'hc404f00;
      15319: inst = 32'h8220000;
      15320: inst = 32'h10408000;
      15321: inst = 32'hc404f01;
      15322: inst = 32'h8220000;
      15323: inst = 32'h10408000;
      15324: inst = 32'hc404f02;
      15325: inst = 32'h8220000;
      15326: inst = 32'h10408000;
      15327: inst = 32'hc404f03;
      15328: inst = 32'h8220000;
      15329: inst = 32'h10408000;
      15330: inst = 32'hc404f04;
      15331: inst = 32'h8220000;
      15332: inst = 32'h10408000;
      15333: inst = 32'hc404f05;
      15334: inst = 32'h8220000;
      15335: inst = 32'h10408000;
      15336: inst = 32'hc404f1a;
      15337: inst = 32'h8220000;
      15338: inst = 32'h10408000;
      15339: inst = 32'hc404f1b;
      15340: inst = 32'h8220000;
      15341: inst = 32'h10408000;
      15342: inst = 32'hc404f1c;
      15343: inst = 32'h8220000;
      15344: inst = 32'h10408000;
      15345: inst = 32'hc404f1d;
      15346: inst = 32'h8220000;
      15347: inst = 32'h10408000;
      15348: inst = 32'hc404f1e;
      15349: inst = 32'h8220000;
      15350: inst = 32'h10408000;
      15351: inst = 32'hc404f1f;
      15352: inst = 32'h8220000;
      15353: inst = 32'h10408000;
      15354: inst = 32'hc404f60;
      15355: inst = 32'h8220000;
      15356: inst = 32'h10408000;
      15357: inst = 32'hc404f61;
      15358: inst = 32'h8220000;
      15359: inst = 32'h10408000;
      15360: inst = 32'hc404f62;
      15361: inst = 32'h8220000;
      15362: inst = 32'h10408000;
      15363: inst = 32'hc404f63;
      15364: inst = 32'h8220000;
      15365: inst = 32'h10408000;
      15366: inst = 32'hc404f64;
      15367: inst = 32'h8220000;
      15368: inst = 32'h10408000;
      15369: inst = 32'hc404f65;
      15370: inst = 32'h8220000;
      15371: inst = 32'h10408000;
      15372: inst = 32'hc404f66;
      15373: inst = 32'h8220000;
      15374: inst = 32'h10408000;
      15375: inst = 32'hc404f67;
      15376: inst = 32'h8220000;
      15377: inst = 32'h10408000;
      15378: inst = 32'hc404f78;
      15379: inst = 32'h8220000;
      15380: inst = 32'h10408000;
      15381: inst = 32'hc404f79;
      15382: inst = 32'h8220000;
      15383: inst = 32'h10408000;
      15384: inst = 32'hc404f7a;
      15385: inst = 32'h8220000;
      15386: inst = 32'h10408000;
      15387: inst = 32'hc404f7b;
      15388: inst = 32'h8220000;
      15389: inst = 32'h10408000;
      15390: inst = 32'hc404f7c;
      15391: inst = 32'h8220000;
      15392: inst = 32'h10408000;
      15393: inst = 32'hc404f7d;
      15394: inst = 32'h8220000;
      15395: inst = 32'h10408000;
      15396: inst = 32'hc404f7e;
      15397: inst = 32'h8220000;
      15398: inst = 32'h10408000;
      15399: inst = 32'hc404f7f;
      15400: inst = 32'h8220000;
      15401: inst = 32'h10408000;
      15402: inst = 32'hc404fc0;
      15403: inst = 32'h8220000;
      15404: inst = 32'h10408000;
      15405: inst = 32'hc404fc1;
      15406: inst = 32'h8220000;
      15407: inst = 32'h10408000;
      15408: inst = 32'hc404fc2;
      15409: inst = 32'h8220000;
      15410: inst = 32'h10408000;
      15411: inst = 32'hc404fc3;
      15412: inst = 32'h8220000;
      15413: inst = 32'h10408000;
      15414: inst = 32'hc404fc4;
      15415: inst = 32'h8220000;
      15416: inst = 32'h10408000;
      15417: inst = 32'hc404fc6;
      15418: inst = 32'h8220000;
      15419: inst = 32'h10408000;
      15420: inst = 32'hc404fc7;
      15421: inst = 32'h8220000;
      15422: inst = 32'h10408000;
      15423: inst = 32'hc404fd8;
      15424: inst = 32'h8220000;
      15425: inst = 32'h10408000;
      15426: inst = 32'hc404fd9;
      15427: inst = 32'h8220000;
      15428: inst = 32'h10408000;
      15429: inst = 32'hc404fdb;
      15430: inst = 32'h8220000;
      15431: inst = 32'h10408000;
      15432: inst = 32'hc404fdc;
      15433: inst = 32'h8220000;
      15434: inst = 32'h10408000;
      15435: inst = 32'hc404fdd;
      15436: inst = 32'h8220000;
      15437: inst = 32'h10408000;
      15438: inst = 32'hc404fde;
      15439: inst = 32'h8220000;
      15440: inst = 32'h10408000;
      15441: inst = 32'hc404fdf;
      15442: inst = 32'h8220000;
      15443: inst = 32'h10408000;
      15444: inst = 32'hc405020;
      15445: inst = 32'h8220000;
      15446: inst = 32'h10408000;
      15447: inst = 32'hc405021;
      15448: inst = 32'h8220000;
      15449: inst = 32'h10408000;
      15450: inst = 32'hc405022;
      15451: inst = 32'h8220000;
      15452: inst = 32'h10408000;
      15453: inst = 32'hc405023;
      15454: inst = 32'h8220000;
      15455: inst = 32'h10408000;
      15456: inst = 32'hc405026;
      15457: inst = 32'h8220000;
      15458: inst = 32'h10408000;
      15459: inst = 32'hc405027;
      15460: inst = 32'h8220000;
      15461: inst = 32'h10408000;
      15462: inst = 32'hc405038;
      15463: inst = 32'h8220000;
      15464: inst = 32'h10408000;
      15465: inst = 32'hc405039;
      15466: inst = 32'h8220000;
      15467: inst = 32'h10408000;
      15468: inst = 32'hc40503c;
      15469: inst = 32'h8220000;
      15470: inst = 32'h10408000;
      15471: inst = 32'hc40503d;
      15472: inst = 32'h8220000;
      15473: inst = 32'h10408000;
      15474: inst = 32'hc40503e;
      15475: inst = 32'h8220000;
      15476: inst = 32'h10408000;
      15477: inst = 32'hc40503f;
      15478: inst = 32'h8220000;
      15479: inst = 32'h10408000;
      15480: inst = 32'hc40507f;
      15481: inst = 32'h8220000;
      15482: inst = 32'h10408000;
      15483: inst = 32'hc405080;
      15484: inst = 32'h8220000;
      15485: inst = 32'h10408000;
      15486: inst = 32'hc405081;
      15487: inst = 32'h8220000;
      15488: inst = 32'h10408000;
      15489: inst = 32'hc405082;
      15490: inst = 32'h8220000;
      15491: inst = 32'h10408000;
      15492: inst = 32'hc405086;
      15493: inst = 32'h8220000;
      15494: inst = 32'h10408000;
      15495: inst = 32'hc405087;
      15496: inst = 32'h8220000;
      15497: inst = 32'h10408000;
      15498: inst = 32'hc405098;
      15499: inst = 32'h8220000;
      15500: inst = 32'h10408000;
      15501: inst = 32'hc405099;
      15502: inst = 32'h8220000;
      15503: inst = 32'h10408000;
      15504: inst = 32'hc40509d;
      15505: inst = 32'h8220000;
      15506: inst = 32'h10408000;
      15507: inst = 32'hc40509e;
      15508: inst = 32'h8220000;
      15509: inst = 32'h10408000;
      15510: inst = 32'hc40509f;
      15511: inst = 32'h8220000;
      15512: inst = 32'h10408000;
      15513: inst = 32'hc4050a0;
      15514: inst = 32'h8220000;
      15515: inst = 32'h10408000;
      15516: inst = 32'hc4050df;
      15517: inst = 32'h8220000;
      15518: inst = 32'h10408000;
      15519: inst = 32'hc4050e0;
      15520: inst = 32'h8220000;
      15521: inst = 32'h10408000;
      15522: inst = 32'hc4050e1;
      15523: inst = 32'h8220000;
      15524: inst = 32'h10408000;
      15525: inst = 32'hc4050e2;
      15526: inst = 32'h8220000;
      15527: inst = 32'h10408000;
      15528: inst = 32'hc4050e6;
      15529: inst = 32'h8220000;
      15530: inst = 32'h10408000;
      15531: inst = 32'hc4050e7;
      15532: inst = 32'h8220000;
      15533: inst = 32'h10408000;
      15534: inst = 32'hc4050f8;
      15535: inst = 32'h8220000;
      15536: inst = 32'h10408000;
      15537: inst = 32'hc4050f9;
      15538: inst = 32'h8220000;
      15539: inst = 32'h10408000;
      15540: inst = 32'hc4050fd;
      15541: inst = 32'h8220000;
      15542: inst = 32'h10408000;
      15543: inst = 32'hc4050fe;
      15544: inst = 32'h8220000;
      15545: inst = 32'h10408000;
      15546: inst = 32'hc4050ff;
      15547: inst = 32'h8220000;
      15548: inst = 32'h10408000;
      15549: inst = 32'hc405100;
      15550: inst = 32'h8220000;
      15551: inst = 32'h10408000;
      15552: inst = 32'hc40513f;
      15553: inst = 32'h8220000;
      15554: inst = 32'h10408000;
      15555: inst = 32'hc405140;
      15556: inst = 32'h8220000;
      15557: inst = 32'h10408000;
      15558: inst = 32'hc405141;
      15559: inst = 32'h8220000;
      15560: inst = 32'h10408000;
      15561: inst = 32'hc405146;
      15562: inst = 32'h8220000;
      15563: inst = 32'h10408000;
      15564: inst = 32'hc405147;
      15565: inst = 32'h8220000;
      15566: inst = 32'h10408000;
      15567: inst = 32'hc405158;
      15568: inst = 32'h8220000;
      15569: inst = 32'h10408000;
      15570: inst = 32'hc405159;
      15571: inst = 32'h8220000;
      15572: inst = 32'h10408000;
      15573: inst = 32'hc40515e;
      15574: inst = 32'h8220000;
      15575: inst = 32'h10408000;
      15576: inst = 32'hc40515f;
      15577: inst = 32'h8220000;
      15578: inst = 32'h10408000;
      15579: inst = 32'hc405160;
      15580: inst = 32'h8220000;
      15581: inst = 32'h10408000;
      15582: inst = 32'hc40519f;
      15583: inst = 32'h8220000;
      15584: inst = 32'h10408000;
      15585: inst = 32'hc4051a0;
      15586: inst = 32'h8220000;
      15587: inst = 32'h10408000;
      15588: inst = 32'hc4051a6;
      15589: inst = 32'h8220000;
      15590: inst = 32'h10408000;
      15591: inst = 32'hc4051a7;
      15592: inst = 32'h8220000;
      15593: inst = 32'h10408000;
      15594: inst = 32'hc4051b8;
      15595: inst = 32'h8220000;
      15596: inst = 32'h10408000;
      15597: inst = 32'hc4051b9;
      15598: inst = 32'h8220000;
      15599: inst = 32'h10408000;
      15600: inst = 32'hc4051bf;
      15601: inst = 32'h8220000;
      15602: inst = 32'h10408000;
      15603: inst = 32'hc4051c0;
      15604: inst = 32'h8220000;
      15605: inst = 32'h10408000;
      15606: inst = 32'hc4051ff;
      15607: inst = 32'h8220000;
      15608: inst = 32'h10408000;
      15609: inst = 32'hc405200;
      15610: inst = 32'h8220000;
      15611: inst = 32'h10408000;
      15612: inst = 32'hc405206;
      15613: inst = 32'h8220000;
      15614: inst = 32'h10408000;
      15615: inst = 32'hc405207;
      15616: inst = 32'h8220000;
      15617: inst = 32'h10408000;
      15618: inst = 32'hc405218;
      15619: inst = 32'h8220000;
      15620: inst = 32'h10408000;
      15621: inst = 32'hc405219;
      15622: inst = 32'h8220000;
      15623: inst = 32'h10408000;
      15624: inst = 32'hc40521f;
      15625: inst = 32'h8220000;
      15626: inst = 32'h10408000;
      15627: inst = 32'hc405220;
      15628: inst = 32'h8220000;
      15629: inst = 32'h10408000;
      15630: inst = 32'hc40525f;
      15631: inst = 32'h8220000;
      15632: inst = 32'h10408000;
      15633: inst = 32'hc405260;
      15634: inst = 32'h8220000;
      15635: inst = 32'h10408000;
      15636: inst = 32'hc405266;
      15637: inst = 32'h8220000;
      15638: inst = 32'h10408000;
      15639: inst = 32'hc405267;
      15640: inst = 32'h8220000;
      15641: inst = 32'h10408000;
      15642: inst = 32'hc405278;
      15643: inst = 32'h8220000;
      15644: inst = 32'h10408000;
      15645: inst = 32'hc405279;
      15646: inst = 32'h8220000;
      15647: inst = 32'h10408000;
      15648: inst = 32'hc40527f;
      15649: inst = 32'h8220000;
      15650: inst = 32'h10408000;
      15651: inst = 32'hc405280;
      15652: inst = 32'h8220000;
      15653: inst = 32'h10408000;
      15654: inst = 32'hc4052bf;
      15655: inst = 32'h8220000;
      15656: inst = 32'h10408000;
      15657: inst = 32'hc4052c0;
      15658: inst = 32'h8220000;
      15659: inst = 32'h10408000;
      15660: inst = 32'hc4052c6;
      15661: inst = 32'h8220000;
      15662: inst = 32'h10408000;
      15663: inst = 32'hc4052c7;
      15664: inst = 32'h8220000;
      15665: inst = 32'h10408000;
      15666: inst = 32'hc4052d8;
      15667: inst = 32'h8220000;
      15668: inst = 32'h10408000;
      15669: inst = 32'hc4052d9;
      15670: inst = 32'h8220000;
      15671: inst = 32'h10408000;
      15672: inst = 32'hc4052df;
      15673: inst = 32'h8220000;
      15674: inst = 32'h10408000;
      15675: inst = 32'hc4052e0;
      15676: inst = 32'h8220000;
      15677: inst = 32'hc207bae;
      15678: inst = 32'h10408000;
      15679: inst = 32'hc404ea5;
      15680: inst = 32'h8220000;
      15681: inst = 32'h10408000;
      15682: inst = 32'hc404eba;
      15683: inst = 32'h8220000;
      15684: inst = 32'hc20c5b4;
      15685: inst = 32'h10408000;
      15686: inst = 32'hc404ea6;
      15687: inst = 32'h8220000;
      15688: inst = 32'h10408000;
      15689: inst = 32'hc404eb9;
      15690: inst = 32'h8220000;
      15691: inst = 32'hc20d5f4;
      15692: inst = 32'h10408000;
      15693: inst = 32'hc404ea7;
      15694: inst = 32'h8220000;
      15695: inst = 32'h10408000;
      15696: inst = 32'hc404eb8;
      15697: inst = 32'h8220000;
      15698: inst = 32'hc20a4b1;
      15699: inst = 32'h10408000;
      15700: inst = 32'hc404eff;
      15701: inst = 32'h8220000;
      15702: inst = 32'h10408000;
      15703: inst = 32'hc404f20;
      15704: inst = 32'h8220000;
      15705: inst = 32'h10408000;
      15706: inst = 32'hc404fbf;
      15707: inst = 32'h8220000;
      15708: inst = 32'h10408000;
      15709: inst = 32'hc404fe0;
      15710: inst = 32'h8220000;
      15711: inst = 32'hc2062ed;
      15712: inst = 32'h10408000;
      15713: inst = 32'hc404f06;
      15714: inst = 32'h8220000;
      15715: inst = 32'h10408000;
      15716: inst = 32'hc404f19;
      15717: inst = 32'h8220000;
      15718: inst = 32'hc209450;
      15719: inst = 32'h10408000;
      15720: inst = 32'hc404f07;
      15721: inst = 32'h8220000;
      15722: inst = 32'h10408000;
      15723: inst = 32'hc404f18;
      15724: inst = 32'h8220000;
      15725: inst = 32'h10408000;
      15726: inst = 32'hc405209;
      15727: inst = 32'h8220000;
      15728: inst = 32'h10408000;
      15729: inst = 32'hc405216;
      15730: inst = 32'h8220000;
      15731: inst = 32'hc20a4d1;
      15732: inst = 32'h10408000;
      15733: inst = 32'hc404f5f;
      15734: inst = 32'h8220000;
      15735: inst = 32'h10408000;
      15736: inst = 32'hc404f80;
      15737: inst = 32'h8220000;
      15738: inst = 32'hc204a49;
      15739: inst = 32'h10408000;
      15740: inst = 32'hc404fa8;
      15741: inst = 32'h8220000;
      15742: inst = 32'h10408000;
      15743: inst = 32'hc404fac;
      15744: inst = 32'h8220000;
      15745: inst = 32'h10408000;
      15746: inst = 32'hc405008;
      15747: inst = 32'h8220000;
      15748: inst = 32'h10408000;
      15749: inst = 32'hc40500c;
      15750: inst = 32'h8220000;
      15751: inst = 32'hc205acb;
      15752: inst = 32'h10408000;
      15753: inst = 32'hc404fc5;
      15754: inst = 32'h8220000;
      15755: inst = 32'h10408000;
      15756: inst = 32'hc404fda;
      15757: inst = 32'h8220000;
      15758: inst = 32'h10408000;
      15759: inst = 32'hc405336;
      15760: inst = 32'h8220000;
      15761: inst = 32'h10408000;
      15762: inst = 32'hc405380;
      15763: inst = 32'h8220000;
      15764: inst = 32'h10408000;
      15765: inst = 32'hc40539f;
      15766: inst = 32'h8220000;
      15767: inst = 32'h10408000;
      15768: inst = 32'hc4053dd;
      15769: inst = 32'h8220000;
      15770: inst = 32'h10408000;
      15771: inst = 32'hc405402;
      15772: inst = 32'h8220000;
      15773: inst = 32'hc20630d;
      15774: inst = 32'h10408000;
      15775: inst = 32'hc40501f;
      15776: inst = 32'h8220000;
      15777: inst = 32'h10408000;
      15778: inst = 32'hc405040;
      15779: inst = 32'h8220000;
      15780: inst = 32'hc205aec;
      15781: inst = 32'h10408000;
      15782: inst = 32'hc405024;
      15783: inst = 32'h8220000;
      15784: inst = 32'h10408000;
      15785: inst = 32'hc40503b;
      15786: inst = 32'h8220000;
      15787: inst = 32'h10408000;
      15788: inst = 32'hc405083;
      15789: inst = 32'h8220000;
      15790: inst = 32'h10408000;
      15791: inst = 32'hc40509c;
      15792: inst = 32'h8220000;
      15793: inst = 32'h10408000;
      15794: inst = 32'hc4051a1;
      15795: inst = 32'h8220000;
      15796: inst = 32'h10408000;
      15797: inst = 32'hc4051be;
      15798: inst = 32'h8220000;
      15799: inst = 32'h10408000;
      15800: inst = 32'hc405329;
      15801: inst = 32'h8220000;
      15802: inst = 32'h10408000;
      15803: inst = 32'hc405568;
      15804: inst = 32'h8220000;
      15805: inst = 32'h10408000;
      15806: inst = 32'hc405577;
      15807: inst = 32'h8220000;
      15808: inst = 32'h10408000;
      15809: inst = 32'hc4057a7;
      15810: inst = 32'h8220000;
      15811: inst = 32'h10408000;
      15812: inst = 32'hc4057b8;
      15813: inst = 32'h8220000;
      15814: inst = 32'hc205269;
      15815: inst = 32'h10408000;
      15816: inst = 32'hc405025;
      15817: inst = 32'h8220000;
      15818: inst = 32'h10408000;
      15819: inst = 32'hc40503a;
      15820: inst = 32'h8220000;
      15821: inst = 32'h10408000;
      15822: inst = 32'hc40537e;
      15823: inst = 32'h8220000;
      15824: inst = 32'h10408000;
      15825: inst = 32'hc4053a1;
      15826: inst = 32'h8220000;
      15827: inst = 32'h10408000;
      15828: inst = 32'hc40549c;
      15829: inst = 32'h8220000;
      15830: inst = 32'h10408000;
      15831: inst = 32'hc4054c3;
      15832: inst = 32'h8220000;
      15833: inst = 32'hc20528a;
      15834: inst = 32'h10408000;
      15835: inst = 32'hc405084;
      15836: inst = 32'h8220000;
      15837: inst = 32'h10408000;
      15838: inst = 32'hc40509b;
      15839: inst = 32'h8220000;
      15840: inst = 32'h10408000;
      15841: inst = 32'hc4050e3;
      15842: inst = 32'h8220000;
      15843: inst = 32'h10408000;
      15844: inst = 32'hc4050fc;
      15845: inst = 32'h8220000;
      15846: inst = 32'h10408000;
      15847: inst = 32'hc4052c5;
      15848: inst = 32'h8220000;
      15849: inst = 32'h10408000;
      15850: inst = 32'hc4052da;
      15851: inst = 32'h8220000;
      15852: inst = 32'h10408000;
      15853: inst = 32'hc4053e9;
      15854: inst = 32'h8220000;
      15855: inst = 32'h10408000;
      15856: inst = 32'hc4053f6;
      15857: inst = 32'h8220000;
      15858: inst = 32'h10408000;
      15859: inst = 32'hc405449;
      15860: inst = 32'h8220000;
      15861: inst = 32'h10408000;
      15862: inst = 32'hc405456;
      15863: inst = 32'h8220000;
      15864: inst = 32'h10408000;
      15865: inst = 32'hc4054a9;
      15866: inst = 32'h8220000;
      15867: inst = 32'h10408000;
      15868: inst = 32'hc4054b6;
      15869: inst = 32'h8220000;
      15870: inst = 32'h10408000;
      15871: inst = 32'hc405509;
      15872: inst = 32'h8220000;
      15873: inst = 32'h10408000;
      15874: inst = 32'hc405516;
      15875: inst = 32'h8220000;
      15876: inst = 32'h10408000;
      15877: inst = 32'hc40555e;
      15878: inst = 32'h8220000;
      15879: inst = 32'h10408000;
      15880: inst = 32'hc405569;
      15881: inst = 32'h8220000;
      15882: inst = 32'h10408000;
      15883: inst = 32'hc405576;
      15884: inst = 32'h8220000;
      15885: inst = 32'h10408000;
      15886: inst = 32'hc405581;
      15887: inst = 32'h8220000;
      15888: inst = 32'h10408000;
      15889: inst = 32'hc4055c9;
      15890: inst = 32'h8220000;
      15891: inst = 32'h10408000;
      15892: inst = 32'hc4055d6;
      15893: inst = 32'h8220000;
      15894: inst = 32'h10408000;
      15895: inst = 32'hc405628;
      15896: inst = 32'h8220000;
      15897: inst = 32'h10408000;
      15898: inst = 32'hc405629;
      15899: inst = 32'h8220000;
      15900: inst = 32'h10408000;
      15901: inst = 32'hc405636;
      15902: inst = 32'h8220000;
      15903: inst = 32'h10408000;
      15904: inst = 32'hc405637;
      15905: inst = 32'h8220000;
      15906: inst = 32'h10408000;
      15907: inst = 32'hc40567d;
      15908: inst = 32'h8220000;
      15909: inst = 32'h10408000;
      15910: inst = 32'hc405688;
      15911: inst = 32'h8220000;
      15912: inst = 32'h10408000;
      15913: inst = 32'hc405689;
      15914: inst = 32'h8220000;
      15915: inst = 32'h10408000;
      15916: inst = 32'hc405696;
      15917: inst = 32'h8220000;
      15918: inst = 32'h10408000;
      15919: inst = 32'hc405697;
      15920: inst = 32'h8220000;
      15921: inst = 32'h10408000;
      15922: inst = 32'hc4056a2;
      15923: inst = 32'h8220000;
      15924: inst = 32'h10408000;
      15925: inst = 32'hc4056e8;
      15926: inst = 32'h8220000;
      15927: inst = 32'h10408000;
      15928: inst = 32'hc4056e9;
      15929: inst = 32'h8220000;
      15930: inst = 32'h10408000;
      15931: inst = 32'hc4056f6;
      15932: inst = 32'h8220000;
      15933: inst = 32'h10408000;
      15934: inst = 32'hc4056f7;
      15935: inst = 32'h8220000;
      15936: inst = 32'h10408000;
      15937: inst = 32'hc405748;
      15938: inst = 32'h8220000;
      15939: inst = 32'h10408000;
      15940: inst = 32'hc405749;
      15941: inst = 32'h8220000;
      15942: inst = 32'h10408000;
      15943: inst = 32'hc405756;
      15944: inst = 32'h8220000;
      15945: inst = 32'h10408000;
      15946: inst = 32'hc405757;
      15947: inst = 32'h8220000;
      15948: inst = 32'h10408000;
      15949: inst = 32'hc4057a8;
      15950: inst = 32'h8220000;
      15951: inst = 32'h10408000;
      15952: inst = 32'hc4057a9;
      15953: inst = 32'h8220000;
      15954: inst = 32'h10408000;
      15955: inst = 32'hc4057b6;
      15956: inst = 32'h8220000;
      15957: inst = 32'h10408000;
      15958: inst = 32'hc4057b7;
      15959: inst = 32'h8220000;
      15960: inst = 32'hc205aab;
      15961: inst = 32'h10408000;
      15962: inst = 32'hc405142;
      15963: inst = 32'h8220000;
      15964: inst = 32'h10408000;
      15965: inst = 32'hc40515d;
      15966: inst = 32'h8220000;
      15967: inst = 32'hc20cdd4;
      15968: inst = 32'h10408000;
      15969: inst = 32'hc40519e;
      15970: inst = 32'h8220000;
      15971: inst = 32'h10408000;
      15972: inst = 32'hc4051c1;
      15973: inst = 32'h8220000;
      15974: inst = 32'hc209471;
      15975: inst = 32'h10408000;
      15976: inst = 32'hc4051b6;
      15977: inst = 32'h8220000;
      15978: inst = 32'hc20de55;
      15979: inst = 32'h10408000;
      15980: inst = 32'hc4051fd;
      15981: inst = 32'h8220000;
      15982: inst = 32'h10408000;
      15983: inst = 32'hc405222;
      15984: inst = 32'h8220000;
      15985: inst = 32'hc209492;
      15986: inst = 32'h10408000;
      15987: inst = 32'hc4051fe;
      15988: inst = 32'h8220000;
      15989: inst = 32'h10408000;
      15990: inst = 32'hc405221;
      15991: inst = 32'h8220000;
      15992: inst = 32'hc205acc;
      15993: inst = 32'h10408000;
      15994: inst = 32'hc405201;
      15995: inst = 32'h8220000;
      15996: inst = 32'h10408000;
      15997: inst = 32'hc40521e;
      15998: inst = 32'h8220000;
      15999: inst = 32'h10408000;
      16000: inst = 32'hc405261;
      16001: inst = 32'h8220000;
      16002: inst = 32'h10408000;
      16003: inst = 32'hc40527e;
      16004: inst = 32'h8220000;
      16005: inst = 32'h10408000;
      16006: inst = 32'hc4052c1;
      16007: inst = 32'h8220000;
      16008: inst = 32'h10408000;
      16009: inst = 32'hc4052de;
      16010: inst = 32'h8220000;
      16011: inst = 32'hc20e696;
      16012: inst = 32'h10408000;
      16013: inst = 32'hc40525c;
      16014: inst = 32'h8220000;
      16015: inst = 32'h10408000;
      16016: inst = 32'hc405283;
      16017: inst = 32'h8220000;
      16018: inst = 32'hc209cb2;
      16019: inst = 32'h10408000;
      16020: inst = 32'hc40525d;
      16021: inst = 32'h8220000;
      16022: inst = 32'h10408000;
      16023: inst = 32'hc405282;
      16024: inst = 32'h8220000;
      16025: inst = 32'hc208c2f;
      16026: inst = 32'h10408000;
      16027: inst = 32'hc405269;
      16028: inst = 32'h8220000;
      16029: inst = 32'h10408000;
      16030: inst = 32'hc405276;
      16031: inst = 32'h8220000;
      16032: inst = 32'hc20ad33;
      16033: inst = 32'h10408000;
      16034: inst = 32'hc4052bc;
      16035: inst = 32'h8220000;
      16036: inst = 32'h10408000;
      16037: inst = 32'hc4052e3;
      16038: inst = 32'h8220000;
      16039: inst = 32'hc2083ee;
      16040: inst = 32'h10408000;
      16041: inst = 32'hc4052c9;
      16042: inst = 32'h8220000;
      16043: inst = 32'h10408000;
      16044: inst = 32'hc4052d6;
      16045: inst = 32'h8220000;
      16046: inst = 32'hc206b50;
      16047: inst = 32'h10408000;
      16048: inst = 32'hc405300;
      16049: inst = 32'h8220000;
      16050: inst = 32'h10408000;
      16051: inst = 32'hc405301;
      16052: inst = 32'h8220000;
      16053: inst = 32'h10408000;
      16054: inst = 32'hc405302;
      16055: inst = 32'h8220000;
      16056: inst = 32'h10408000;
      16057: inst = 32'hc405303;
      16058: inst = 32'h8220000;
      16059: inst = 32'h10408000;
      16060: inst = 32'hc405304;
      16061: inst = 32'h8220000;
      16062: inst = 32'h10408000;
      16063: inst = 32'hc405305;
      16064: inst = 32'h8220000;
      16065: inst = 32'h10408000;
      16066: inst = 32'hc405306;
      16067: inst = 32'h8220000;
      16068: inst = 32'h10408000;
      16069: inst = 32'hc405307;
      16070: inst = 32'h8220000;
      16071: inst = 32'h10408000;
      16072: inst = 32'hc405308;
      16073: inst = 32'h8220000;
      16074: inst = 32'h10408000;
      16075: inst = 32'hc405309;
      16076: inst = 32'h8220000;
      16077: inst = 32'h10408000;
      16078: inst = 32'hc40530a;
      16079: inst = 32'h8220000;
      16080: inst = 32'h10408000;
      16081: inst = 32'hc40530b;
      16082: inst = 32'h8220000;
      16083: inst = 32'h10408000;
      16084: inst = 32'hc40530c;
      16085: inst = 32'h8220000;
      16086: inst = 32'h10408000;
      16087: inst = 32'hc40530d;
      16088: inst = 32'h8220000;
      16089: inst = 32'h10408000;
      16090: inst = 32'hc40530e;
      16091: inst = 32'h8220000;
      16092: inst = 32'h10408000;
      16093: inst = 32'hc40530f;
      16094: inst = 32'h8220000;
      16095: inst = 32'h10408000;
      16096: inst = 32'hc405310;
      16097: inst = 32'h8220000;
      16098: inst = 32'h10408000;
      16099: inst = 32'hc405311;
      16100: inst = 32'h8220000;
      16101: inst = 32'h10408000;
      16102: inst = 32'hc405312;
      16103: inst = 32'h8220000;
      16104: inst = 32'h10408000;
      16105: inst = 32'hc405313;
      16106: inst = 32'h8220000;
      16107: inst = 32'h10408000;
      16108: inst = 32'hc405314;
      16109: inst = 32'h8220000;
      16110: inst = 32'h10408000;
      16111: inst = 32'hc405315;
      16112: inst = 32'h8220000;
      16113: inst = 32'h10408000;
      16114: inst = 32'hc405316;
      16115: inst = 32'h8220000;
      16116: inst = 32'h10408000;
      16117: inst = 32'hc405317;
      16118: inst = 32'h8220000;
      16119: inst = 32'h10408000;
      16120: inst = 32'hc405318;
      16121: inst = 32'h8220000;
      16122: inst = 32'h10408000;
      16123: inst = 32'hc405319;
      16124: inst = 32'h8220000;
      16125: inst = 32'h10408000;
      16126: inst = 32'hc40531a;
      16127: inst = 32'h8220000;
      16128: inst = 32'h10408000;
      16129: inst = 32'hc40532a;
      16130: inst = 32'h8220000;
      16131: inst = 32'h10408000;
      16132: inst = 32'hc40532b;
      16133: inst = 32'h8220000;
      16134: inst = 32'h10408000;
      16135: inst = 32'hc40532c;
      16136: inst = 32'h8220000;
      16137: inst = 32'h10408000;
      16138: inst = 32'hc40532d;
      16139: inst = 32'h8220000;
      16140: inst = 32'h10408000;
      16141: inst = 32'hc40532e;
      16142: inst = 32'h8220000;
      16143: inst = 32'h10408000;
      16144: inst = 32'hc40532f;
      16145: inst = 32'h8220000;
      16146: inst = 32'h10408000;
      16147: inst = 32'hc405330;
      16148: inst = 32'h8220000;
      16149: inst = 32'h10408000;
      16150: inst = 32'hc405331;
      16151: inst = 32'h8220000;
      16152: inst = 32'h10408000;
      16153: inst = 32'hc405332;
      16154: inst = 32'h8220000;
      16155: inst = 32'h10408000;
      16156: inst = 32'hc405333;
      16157: inst = 32'h8220000;
      16158: inst = 32'h10408000;
      16159: inst = 32'hc405334;
      16160: inst = 32'h8220000;
      16161: inst = 32'h10408000;
      16162: inst = 32'hc405335;
      16163: inst = 32'h8220000;
      16164: inst = 32'h10408000;
      16165: inst = 32'hc405345;
      16166: inst = 32'h8220000;
      16167: inst = 32'h10408000;
      16168: inst = 32'hc405346;
      16169: inst = 32'h8220000;
      16170: inst = 32'h10408000;
      16171: inst = 32'hc405347;
      16172: inst = 32'h8220000;
      16173: inst = 32'h10408000;
      16174: inst = 32'hc405348;
      16175: inst = 32'h8220000;
      16176: inst = 32'h10408000;
      16177: inst = 32'hc405349;
      16178: inst = 32'h8220000;
      16179: inst = 32'h10408000;
      16180: inst = 32'hc40534a;
      16181: inst = 32'h8220000;
      16182: inst = 32'h10408000;
      16183: inst = 32'hc40534b;
      16184: inst = 32'h8220000;
      16185: inst = 32'h10408000;
      16186: inst = 32'hc40534c;
      16187: inst = 32'h8220000;
      16188: inst = 32'h10408000;
      16189: inst = 32'hc40534d;
      16190: inst = 32'h8220000;
      16191: inst = 32'h10408000;
      16192: inst = 32'hc40534e;
      16193: inst = 32'h8220000;
      16194: inst = 32'h10408000;
      16195: inst = 32'hc40534f;
      16196: inst = 32'h8220000;
      16197: inst = 32'h10408000;
      16198: inst = 32'hc405350;
      16199: inst = 32'h8220000;
      16200: inst = 32'h10408000;
      16201: inst = 32'hc405351;
      16202: inst = 32'h8220000;
      16203: inst = 32'h10408000;
      16204: inst = 32'hc405352;
      16205: inst = 32'h8220000;
      16206: inst = 32'h10408000;
      16207: inst = 32'hc405353;
      16208: inst = 32'h8220000;
      16209: inst = 32'h10408000;
      16210: inst = 32'hc405354;
      16211: inst = 32'h8220000;
      16212: inst = 32'h10408000;
      16213: inst = 32'hc405355;
      16214: inst = 32'h8220000;
      16215: inst = 32'h10408000;
      16216: inst = 32'hc405356;
      16217: inst = 32'h8220000;
      16218: inst = 32'h10408000;
      16219: inst = 32'hc405357;
      16220: inst = 32'h8220000;
      16221: inst = 32'h10408000;
      16222: inst = 32'hc405358;
      16223: inst = 32'h8220000;
      16224: inst = 32'h10408000;
      16225: inst = 32'hc405359;
      16226: inst = 32'h8220000;
      16227: inst = 32'h10408000;
      16228: inst = 32'hc40535a;
      16229: inst = 32'h8220000;
      16230: inst = 32'h10408000;
      16231: inst = 32'hc40535b;
      16232: inst = 32'h8220000;
      16233: inst = 32'h10408000;
      16234: inst = 32'hc40535c;
      16235: inst = 32'h8220000;
      16236: inst = 32'h10408000;
      16237: inst = 32'hc40535d;
      16238: inst = 32'h8220000;
      16239: inst = 32'h10408000;
      16240: inst = 32'hc40535e;
      16241: inst = 32'h8220000;
      16242: inst = 32'h10408000;
      16243: inst = 32'hc40535f;
      16244: inst = 32'h8220000;
      16245: inst = 32'h10408000;
      16246: inst = 32'hc405360;
      16247: inst = 32'h8220000;
      16248: inst = 32'h10408000;
      16249: inst = 32'hc405361;
      16250: inst = 32'h8220000;
      16251: inst = 32'h10408000;
      16252: inst = 32'hc405362;
      16253: inst = 32'h8220000;
      16254: inst = 32'h10408000;
      16255: inst = 32'hc405363;
      16256: inst = 32'h8220000;
      16257: inst = 32'h10408000;
      16258: inst = 32'hc405364;
      16259: inst = 32'h8220000;
      16260: inst = 32'h10408000;
      16261: inst = 32'hc405365;
      16262: inst = 32'h8220000;
      16263: inst = 32'h10408000;
      16264: inst = 32'hc405366;
      16265: inst = 32'h8220000;
      16266: inst = 32'h10408000;
      16267: inst = 32'hc405367;
      16268: inst = 32'h8220000;
      16269: inst = 32'h10408000;
      16270: inst = 32'hc405368;
      16271: inst = 32'h8220000;
      16272: inst = 32'h10408000;
      16273: inst = 32'hc405369;
      16274: inst = 32'h8220000;
      16275: inst = 32'h10408000;
      16276: inst = 32'hc40536a;
      16277: inst = 32'h8220000;
      16278: inst = 32'h10408000;
      16279: inst = 32'hc40536b;
      16280: inst = 32'h8220000;
      16281: inst = 32'h10408000;
      16282: inst = 32'hc40536c;
      16283: inst = 32'h8220000;
      16284: inst = 32'h10408000;
      16285: inst = 32'hc40536d;
      16286: inst = 32'h8220000;
      16287: inst = 32'h10408000;
      16288: inst = 32'hc40536e;
      16289: inst = 32'h8220000;
      16290: inst = 32'h10408000;
      16291: inst = 32'hc40536f;
      16292: inst = 32'h8220000;
      16293: inst = 32'h10408000;
      16294: inst = 32'hc405370;
      16295: inst = 32'h8220000;
      16296: inst = 32'h10408000;
      16297: inst = 32'hc405371;
      16298: inst = 32'h8220000;
      16299: inst = 32'h10408000;
      16300: inst = 32'hc405372;
      16301: inst = 32'h8220000;
      16302: inst = 32'h10408000;
      16303: inst = 32'hc405373;
      16304: inst = 32'h8220000;
      16305: inst = 32'h10408000;
      16306: inst = 32'hc405374;
      16307: inst = 32'h8220000;
      16308: inst = 32'h10408000;
      16309: inst = 32'hc405375;
      16310: inst = 32'h8220000;
      16311: inst = 32'h10408000;
      16312: inst = 32'hc405376;
      16313: inst = 32'h8220000;
      16314: inst = 32'h10408000;
      16315: inst = 32'hc405377;
      16316: inst = 32'h8220000;
      16317: inst = 32'h10408000;
      16318: inst = 32'hc405378;
      16319: inst = 32'h8220000;
      16320: inst = 32'h10408000;
      16321: inst = 32'hc405379;
      16322: inst = 32'h8220000;
      16323: inst = 32'h10408000;
      16324: inst = 32'hc40538a;
      16325: inst = 32'h8220000;
      16326: inst = 32'h10408000;
      16327: inst = 32'hc40538b;
      16328: inst = 32'h8220000;
      16329: inst = 32'h10408000;
      16330: inst = 32'hc40538c;
      16331: inst = 32'h8220000;
      16332: inst = 32'h10408000;
      16333: inst = 32'hc40538d;
      16334: inst = 32'h8220000;
      16335: inst = 32'h10408000;
      16336: inst = 32'hc40538e;
      16337: inst = 32'h8220000;
      16338: inst = 32'h10408000;
      16339: inst = 32'hc40538f;
      16340: inst = 32'h8220000;
      16341: inst = 32'h10408000;
      16342: inst = 32'hc405390;
      16343: inst = 32'h8220000;
      16344: inst = 32'h10408000;
      16345: inst = 32'hc405391;
      16346: inst = 32'h8220000;
      16347: inst = 32'h10408000;
      16348: inst = 32'hc405392;
      16349: inst = 32'h8220000;
      16350: inst = 32'h10408000;
      16351: inst = 32'hc405393;
      16352: inst = 32'h8220000;
      16353: inst = 32'h10408000;
      16354: inst = 32'hc405394;
      16355: inst = 32'h8220000;
      16356: inst = 32'h10408000;
      16357: inst = 32'hc405395;
      16358: inst = 32'h8220000;
      16359: inst = 32'h10408000;
      16360: inst = 32'hc4053a6;
      16361: inst = 32'h8220000;
      16362: inst = 32'h10408000;
      16363: inst = 32'hc4053a7;
      16364: inst = 32'h8220000;
      16365: inst = 32'h10408000;
      16366: inst = 32'hc4053a8;
      16367: inst = 32'h8220000;
      16368: inst = 32'h10408000;
      16369: inst = 32'hc4053a9;
      16370: inst = 32'h8220000;
      16371: inst = 32'h10408000;
      16372: inst = 32'hc4053aa;
      16373: inst = 32'h8220000;
      16374: inst = 32'h10408000;
      16375: inst = 32'hc4053ab;
      16376: inst = 32'h8220000;
      16377: inst = 32'h10408000;
      16378: inst = 32'hc4053ac;
      16379: inst = 32'h8220000;
      16380: inst = 32'h10408000;
      16381: inst = 32'hc4053ad;
      16382: inst = 32'h8220000;
      16383: inst = 32'h10408000;
      16384: inst = 32'hc4053ae;
      16385: inst = 32'h8220000;
      16386: inst = 32'h10408000;
      16387: inst = 32'hc4053af;
      16388: inst = 32'h8220000;
      16389: inst = 32'h10408000;
      16390: inst = 32'hc4053b0;
      16391: inst = 32'h8220000;
      16392: inst = 32'h10408000;
      16393: inst = 32'hc4053b1;
      16394: inst = 32'h8220000;
      16395: inst = 32'h10408000;
      16396: inst = 32'hc4053b2;
      16397: inst = 32'h8220000;
      16398: inst = 32'h10408000;
      16399: inst = 32'hc4053b3;
      16400: inst = 32'h8220000;
      16401: inst = 32'h10408000;
      16402: inst = 32'hc4053b4;
      16403: inst = 32'h8220000;
      16404: inst = 32'h10408000;
      16405: inst = 32'hc4053b5;
      16406: inst = 32'h8220000;
      16407: inst = 32'h10408000;
      16408: inst = 32'hc4053b6;
      16409: inst = 32'h8220000;
      16410: inst = 32'h10408000;
      16411: inst = 32'hc4053b7;
      16412: inst = 32'h8220000;
      16413: inst = 32'h10408000;
      16414: inst = 32'hc4053b8;
      16415: inst = 32'h8220000;
      16416: inst = 32'h10408000;
      16417: inst = 32'hc4053b9;
      16418: inst = 32'h8220000;
      16419: inst = 32'h10408000;
      16420: inst = 32'hc4053ba;
      16421: inst = 32'h8220000;
      16422: inst = 32'h10408000;
      16423: inst = 32'hc4053bb;
      16424: inst = 32'h8220000;
      16425: inst = 32'h10408000;
      16426: inst = 32'hc4053bc;
      16427: inst = 32'h8220000;
      16428: inst = 32'h10408000;
      16429: inst = 32'hc4053bd;
      16430: inst = 32'h8220000;
      16431: inst = 32'h10408000;
      16432: inst = 32'hc4053be;
      16433: inst = 32'h8220000;
      16434: inst = 32'h10408000;
      16435: inst = 32'hc4053bf;
      16436: inst = 32'h8220000;
      16437: inst = 32'h10408000;
      16438: inst = 32'hc4053c0;
      16439: inst = 32'h8220000;
      16440: inst = 32'h10408000;
      16441: inst = 32'hc4053c1;
      16442: inst = 32'h8220000;
      16443: inst = 32'h10408000;
      16444: inst = 32'hc4053c2;
      16445: inst = 32'h8220000;
      16446: inst = 32'h10408000;
      16447: inst = 32'hc4053c3;
      16448: inst = 32'h8220000;
      16449: inst = 32'h10408000;
      16450: inst = 32'hc4053c4;
      16451: inst = 32'h8220000;
      16452: inst = 32'h10408000;
      16453: inst = 32'hc4053c5;
      16454: inst = 32'h8220000;
      16455: inst = 32'h10408000;
      16456: inst = 32'hc4053c6;
      16457: inst = 32'h8220000;
      16458: inst = 32'h10408000;
      16459: inst = 32'hc4053c7;
      16460: inst = 32'h8220000;
      16461: inst = 32'h10408000;
      16462: inst = 32'hc4053c8;
      16463: inst = 32'h8220000;
      16464: inst = 32'h10408000;
      16465: inst = 32'hc4053c9;
      16466: inst = 32'h8220000;
      16467: inst = 32'h10408000;
      16468: inst = 32'hc4053ca;
      16469: inst = 32'h8220000;
      16470: inst = 32'h10408000;
      16471: inst = 32'hc4053cb;
      16472: inst = 32'h8220000;
      16473: inst = 32'h10408000;
      16474: inst = 32'hc4053cc;
      16475: inst = 32'h8220000;
      16476: inst = 32'h10408000;
      16477: inst = 32'hc4053cd;
      16478: inst = 32'h8220000;
      16479: inst = 32'h10408000;
      16480: inst = 32'hc4053ce;
      16481: inst = 32'h8220000;
      16482: inst = 32'h10408000;
      16483: inst = 32'hc4053cf;
      16484: inst = 32'h8220000;
      16485: inst = 32'h10408000;
      16486: inst = 32'hc4053d0;
      16487: inst = 32'h8220000;
      16488: inst = 32'h10408000;
      16489: inst = 32'hc4053d1;
      16490: inst = 32'h8220000;
      16491: inst = 32'h10408000;
      16492: inst = 32'hc4053d2;
      16493: inst = 32'h8220000;
      16494: inst = 32'h10408000;
      16495: inst = 32'hc4053d3;
      16496: inst = 32'h8220000;
      16497: inst = 32'h10408000;
      16498: inst = 32'hc4053d4;
      16499: inst = 32'h8220000;
      16500: inst = 32'h10408000;
      16501: inst = 32'hc4053d5;
      16502: inst = 32'h8220000;
      16503: inst = 32'h10408000;
      16504: inst = 32'hc4053d6;
      16505: inst = 32'h8220000;
      16506: inst = 32'h10408000;
      16507: inst = 32'hc4053d7;
      16508: inst = 32'h8220000;
      16509: inst = 32'h10408000;
      16510: inst = 32'hc4053d8;
      16511: inst = 32'h8220000;
      16512: inst = 32'h10408000;
      16513: inst = 32'hc4053ea;
      16514: inst = 32'h8220000;
      16515: inst = 32'h10408000;
      16516: inst = 32'hc4053eb;
      16517: inst = 32'h8220000;
      16518: inst = 32'h10408000;
      16519: inst = 32'hc4053ec;
      16520: inst = 32'h8220000;
      16521: inst = 32'h10408000;
      16522: inst = 32'hc4053ed;
      16523: inst = 32'h8220000;
      16524: inst = 32'h10408000;
      16525: inst = 32'hc4053ee;
      16526: inst = 32'h8220000;
      16527: inst = 32'h10408000;
      16528: inst = 32'hc4053ef;
      16529: inst = 32'h8220000;
      16530: inst = 32'h10408000;
      16531: inst = 32'hc4053f0;
      16532: inst = 32'h8220000;
      16533: inst = 32'h10408000;
      16534: inst = 32'hc4053f1;
      16535: inst = 32'h8220000;
      16536: inst = 32'h10408000;
      16537: inst = 32'hc4053f2;
      16538: inst = 32'h8220000;
      16539: inst = 32'h10408000;
      16540: inst = 32'hc4053f3;
      16541: inst = 32'h8220000;
      16542: inst = 32'h10408000;
      16543: inst = 32'hc4053f4;
      16544: inst = 32'h8220000;
      16545: inst = 32'h10408000;
      16546: inst = 32'hc4053f5;
      16547: inst = 32'h8220000;
      16548: inst = 32'h10408000;
      16549: inst = 32'hc405407;
      16550: inst = 32'h8220000;
      16551: inst = 32'h10408000;
      16552: inst = 32'hc405408;
      16553: inst = 32'h8220000;
      16554: inst = 32'h10408000;
      16555: inst = 32'hc405409;
      16556: inst = 32'h8220000;
      16557: inst = 32'h10408000;
      16558: inst = 32'hc40540a;
      16559: inst = 32'h8220000;
      16560: inst = 32'h10408000;
      16561: inst = 32'hc40540b;
      16562: inst = 32'h8220000;
      16563: inst = 32'h10408000;
      16564: inst = 32'hc40540c;
      16565: inst = 32'h8220000;
      16566: inst = 32'h10408000;
      16567: inst = 32'hc40540d;
      16568: inst = 32'h8220000;
      16569: inst = 32'h10408000;
      16570: inst = 32'hc40540e;
      16571: inst = 32'h8220000;
      16572: inst = 32'h10408000;
      16573: inst = 32'hc40540f;
      16574: inst = 32'h8220000;
      16575: inst = 32'h10408000;
      16576: inst = 32'hc405410;
      16577: inst = 32'h8220000;
      16578: inst = 32'h10408000;
      16579: inst = 32'hc405411;
      16580: inst = 32'h8220000;
      16581: inst = 32'h10408000;
      16582: inst = 32'hc405412;
      16583: inst = 32'h8220000;
      16584: inst = 32'h10408000;
      16585: inst = 32'hc405413;
      16586: inst = 32'h8220000;
      16587: inst = 32'h10408000;
      16588: inst = 32'hc405414;
      16589: inst = 32'h8220000;
      16590: inst = 32'h10408000;
      16591: inst = 32'hc405415;
      16592: inst = 32'h8220000;
      16593: inst = 32'h10408000;
      16594: inst = 32'hc405416;
      16595: inst = 32'h8220000;
      16596: inst = 32'h10408000;
      16597: inst = 32'hc405417;
      16598: inst = 32'h8220000;
      16599: inst = 32'h10408000;
      16600: inst = 32'hc405418;
      16601: inst = 32'h8220000;
      16602: inst = 32'h10408000;
      16603: inst = 32'hc405419;
      16604: inst = 32'h8220000;
      16605: inst = 32'h10408000;
      16606: inst = 32'hc40541a;
      16607: inst = 32'h8220000;
      16608: inst = 32'h10408000;
      16609: inst = 32'hc40541b;
      16610: inst = 32'h8220000;
      16611: inst = 32'h10408000;
      16612: inst = 32'hc40541c;
      16613: inst = 32'h8220000;
      16614: inst = 32'h10408000;
      16615: inst = 32'hc40541d;
      16616: inst = 32'h8220000;
      16617: inst = 32'h10408000;
      16618: inst = 32'hc40541e;
      16619: inst = 32'h8220000;
      16620: inst = 32'h10408000;
      16621: inst = 32'hc40541f;
      16622: inst = 32'h8220000;
      16623: inst = 32'h10408000;
      16624: inst = 32'hc405420;
      16625: inst = 32'h8220000;
      16626: inst = 32'h10408000;
      16627: inst = 32'hc405421;
      16628: inst = 32'h8220000;
      16629: inst = 32'h10408000;
      16630: inst = 32'hc405422;
      16631: inst = 32'h8220000;
      16632: inst = 32'h10408000;
      16633: inst = 32'hc405423;
      16634: inst = 32'h8220000;
      16635: inst = 32'h10408000;
      16636: inst = 32'hc405424;
      16637: inst = 32'h8220000;
      16638: inst = 32'h10408000;
      16639: inst = 32'hc405425;
      16640: inst = 32'h8220000;
      16641: inst = 32'h10408000;
      16642: inst = 32'hc405426;
      16643: inst = 32'h8220000;
      16644: inst = 32'h10408000;
      16645: inst = 32'hc405427;
      16646: inst = 32'h8220000;
      16647: inst = 32'h10408000;
      16648: inst = 32'hc405428;
      16649: inst = 32'h8220000;
      16650: inst = 32'h10408000;
      16651: inst = 32'hc405429;
      16652: inst = 32'h8220000;
      16653: inst = 32'h10408000;
      16654: inst = 32'hc40542a;
      16655: inst = 32'h8220000;
      16656: inst = 32'h10408000;
      16657: inst = 32'hc40542b;
      16658: inst = 32'h8220000;
      16659: inst = 32'h10408000;
      16660: inst = 32'hc40542c;
      16661: inst = 32'h8220000;
      16662: inst = 32'h10408000;
      16663: inst = 32'hc40542d;
      16664: inst = 32'h8220000;
      16665: inst = 32'h10408000;
      16666: inst = 32'hc40542e;
      16667: inst = 32'h8220000;
      16668: inst = 32'h10408000;
      16669: inst = 32'hc40542f;
      16670: inst = 32'h8220000;
      16671: inst = 32'h10408000;
      16672: inst = 32'hc405430;
      16673: inst = 32'h8220000;
      16674: inst = 32'h10408000;
      16675: inst = 32'hc405431;
      16676: inst = 32'h8220000;
      16677: inst = 32'h10408000;
      16678: inst = 32'hc405432;
      16679: inst = 32'h8220000;
      16680: inst = 32'h10408000;
      16681: inst = 32'hc405433;
      16682: inst = 32'h8220000;
      16683: inst = 32'h10408000;
      16684: inst = 32'hc405434;
      16685: inst = 32'h8220000;
      16686: inst = 32'h10408000;
      16687: inst = 32'hc405435;
      16688: inst = 32'h8220000;
      16689: inst = 32'h10408000;
      16690: inst = 32'hc405436;
      16691: inst = 32'h8220000;
      16692: inst = 32'h10408000;
      16693: inst = 32'hc405437;
      16694: inst = 32'h8220000;
      16695: inst = 32'h10408000;
      16696: inst = 32'hc405438;
      16697: inst = 32'h8220000;
      16698: inst = 32'h10408000;
      16699: inst = 32'hc40544a;
      16700: inst = 32'h8220000;
      16701: inst = 32'h10408000;
      16702: inst = 32'hc40544b;
      16703: inst = 32'h8220000;
      16704: inst = 32'h10408000;
      16705: inst = 32'hc40544c;
      16706: inst = 32'h8220000;
      16707: inst = 32'h10408000;
      16708: inst = 32'hc40544d;
      16709: inst = 32'h8220000;
      16710: inst = 32'h10408000;
      16711: inst = 32'hc40544e;
      16712: inst = 32'h8220000;
      16713: inst = 32'h10408000;
      16714: inst = 32'hc40544f;
      16715: inst = 32'h8220000;
      16716: inst = 32'h10408000;
      16717: inst = 32'hc405450;
      16718: inst = 32'h8220000;
      16719: inst = 32'h10408000;
      16720: inst = 32'hc405451;
      16721: inst = 32'h8220000;
      16722: inst = 32'h10408000;
      16723: inst = 32'hc405452;
      16724: inst = 32'h8220000;
      16725: inst = 32'h10408000;
      16726: inst = 32'hc405453;
      16727: inst = 32'h8220000;
      16728: inst = 32'h10408000;
      16729: inst = 32'hc405454;
      16730: inst = 32'h8220000;
      16731: inst = 32'h10408000;
      16732: inst = 32'hc405455;
      16733: inst = 32'h8220000;
      16734: inst = 32'h10408000;
      16735: inst = 32'hc405467;
      16736: inst = 32'h8220000;
      16737: inst = 32'h10408000;
      16738: inst = 32'hc405468;
      16739: inst = 32'h8220000;
      16740: inst = 32'h10408000;
      16741: inst = 32'hc405469;
      16742: inst = 32'h8220000;
      16743: inst = 32'h10408000;
      16744: inst = 32'hc40546a;
      16745: inst = 32'h8220000;
      16746: inst = 32'h10408000;
      16747: inst = 32'hc40546b;
      16748: inst = 32'h8220000;
      16749: inst = 32'h10408000;
      16750: inst = 32'hc40546c;
      16751: inst = 32'h8220000;
      16752: inst = 32'h10408000;
      16753: inst = 32'hc40546d;
      16754: inst = 32'h8220000;
      16755: inst = 32'h10408000;
      16756: inst = 32'hc40546e;
      16757: inst = 32'h8220000;
      16758: inst = 32'h10408000;
      16759: inst = 32'hc40546f;
      16760: inst = 32'h8220000;
      16761: inst = 32'h10408000;
      16762: inst = 32'hc405470;
      16763: inst = 32'h8220000;
      16764: inst = 32'h10408000;
      16765: inst = 32'hc405471;
      16766: inst = 32'h8220000;
      16767: inst = 32'h10408000;
      16768: inst = 32'hc405472;
      16769: inst = 32'h8220000;
      16770: inst = 32'h10408000;
      16771: inst = 32'hc405473;
      16772: inst = 32'h8220000;
      16773: inst = 32'h10408000;
      16774: inst = 32'hc405474;
      16775: inst = 32'h8220000;
      16776: inst = 32'h10408000;
      16777: inst = 32'hc405475;
      16778: inst = 32'h8220000;
      16779: inst = 32'h10408000;
      16780: inst = 32'hc405476;
      16781: inst = 32'h8220000;
      16782: inst = 32'h10408000;
      16783: inst = 32'hc405477;
      16784: inst = 32'h8220000;
      16785: inst = 32'h10408000;
      16786: inst = 32'hc405478;
      16787: inst = 32'h8220000;
      16788: inst = 32'h10408000;
      16789: inst = 32'hc405479;
      16790: inst = 32'h8220000;
      16791: inst = 32'h10408000;
      16792: inst = 32'hc40547a;
      16793: inst = 32'h8220000;
      16794: inst = 32'h10408000;
      16795: inst = 32'hc40547b;
      16796: inst = 32'h8220000;
      16797: inst = 32'h10408000;
      16798: inst = 32'hc40547c;
      16799: inst = 32'h8220000;
      16800: inst = 32'h10408000;
      16801: inst = 32'hc40547d;
      16802: inst = 32'h8220000;
      16803: inst = 32'h10408000;
      16804: inst = 32'hc40547e;
      16805: inst = 32'h8220000;
      16806: inst = 32'h10408000;
      16807: inst = 32'hc40547f;
      16808: inst = 32'h8220000;
      16809: inst = 32'h10408000;
      16810: inst = 32'hc405480;
      16811: inst = 32'h8220000;
      16812: inst = 32'h10408000;
      16813: inst = 32'hc405481;
      16814: inst = 32'h8220000;
      16815: inst = 32'h10408000;
      16816: inst = 32'hc405482;
      16817: inst = 32'h8220000;
      16818: inst = 32'h10408000;
      16819: inst = 32'hc405483;
      16820: inst = 32'h8220000;
      16821: inst = 32'h10408000;
      16822: inst = 32'hc405484;
      16823: inst = 32'h8220000;
      16824: inst = 32'h10408000;
      16825: inst = 32'hc405485;
      16826: inst = 32'h8220000;
      16827: inst = 32'h10408000;
      16828: inst = 32'hc405486;
      16829: inst = 32'h8220000;
      16830: inst = 32'h10408000;
      16831: inst = 32'hc405487;
      16832: inst = 32'h8220000;
      16833: inst = 32'h10408000;
      16834: inst = 32'hc405488;
      16835: inst = 32'h8220000;
      16836: inst = 32'h10408000;
      16837: inst = 32'hc405489;
      16838: inst = 32'h8220000;
      16839: inst = 32'h10408000;
      16840: inst = 32'hc40548a;
      16841: inst = 32'h8220000;
      16842: inst = 32'h10408000;
      16843: inst = 32'hc40548b;
      16844: inst = 32'h8220000;
      16845: inst = 32'h10408000;
      16846: inst = 32'hc40548c;
      16847: inst = 32'h8220000;
      16848: inst = 32'h10408000;
      16849: inst = 32'hc40548d;
      16850: inst = 32'h8220000;
      16851: inst = 32'h10408000;
      16852: inst = 32'hc40548e;
      16853: inst = 32'h8220000;
      16854: inst = 32'h10408000;
      16855: inst = 32'hc40548f;
      16856: inst = 32'h8220000;
      16857: inst = 32'h10408000;
      16858: inst = 32'hc405490;
      16859: inst = 32'h8220000;
      16860: inst = 32'h10408000;
      16861: inst = 32'hc405491;
      16862: inst = 32'h8220000;
      16863: inst = 32'h10408000;
      16864: inst = 32'hc405492;
      16865: inst = 32'h8220000;
      16866: inst = 32'h10408000;
      16867: inst = 32'hc405493;
      16868: inst = 32'h8220000;
      16869: inst = 32'h10408000;
      16870: inst = 32'hc405494;
      16871: inst = 32'h8220000;
      16872: inst = 32'h10408000;
      16873: inst = 32'hc405495;
      16874: inst = 32'h8220000;
      16875: inst = 32'h10408000;
      16876: inst = 32'hc405496;
      16877: inst = 32'h8220000;
      16878: inst = 32'h10408000;
      16879: inst = 32'hc405497;
      16880: inst = 32'h8220000;
      16881: inst = 32'h10408000;
      16882: inst = 32'hc4054aa;
      16883: inst = 32'h8220000;
      16884: inst = 32'h10408000;
      16885: inst = 32'hc4054ab;
      16886: inst = 32'h8220000;
      16887: inst = 32'h10408000;
      16888: inst = 32'hc4054ac;
      16889: inst = 32'h8220000;
      16890: inst = 32'h10408000;
      16891: inst = 32'hc4054ad;
      16892: inst = 32'h8220000;
      16893: inst = 32'h10408000;
      16894: inst = 32'hc4054ae;
      16895: inst = 32'h8220000;
      16896: inst = 32'h10408000;
      16897: inst = 32'hc4054af;
      16898: inst = 32'h8220000;
      16899: inst = 32'h10408000;
      16900: inst = 32'hc4054b0;
      16901: inst = 32'h8220000;
      16902: inst = 32'h10408000;
      16903: inst = 32'hc4054b1;
      16904: inst = 32'h8220000;
      16905: inst = 32'h10408000;
      16906: inst = 32'hc4054b2;
      16907: inst = 32'h8220000;
      16908: inst = 32'h10408000;
      16909: inst = 32'hc4054b3;
      16910: inst = 32'h8220000;
      16911: inst = 32'h10408000;
      16912: inst = 32'hc4054b4;
      16913: inst = 32'h8220000;
      16914: inst = 32'h10408000;
      16915: inst = 32'hc4054b5;
      16916: inst = 32'h8220000;
      16917: inst = 32'h10408000;
      16918: inst = 32'hc4054c8;
      16919: inst = 32'h8220000;
      16920: inst = 32'h10408000;
      16921: inst = 32'hc4054c9;
      16922: inst = 32'h8220000;
      16923: inst = 32'h10408000;
      16924: inst = 32'hc4054ca;
      16925: inst = 32'h8220000;
      16926: inst = 32'h10408000;
      16927: inst = 32'hc4054cb;
      16928: inst = 32'h8220000;
      16929: inst = 32'h10408000;
      16930: inst = 32'hc4054cc;
      16931: inst = 32'h8220000;
      16932: inst = 32'h10408000;
      16933: inst = 32'hc4054cd;
      16934: inst = 32'h8220000;
      16935: inst = 32'h10408000;
      16936: inst = 32'hc4054ce;
      16937: inst = 32'h8220000;
      16938: inst = 32'h10408000;
      16939: inst = 32'hc4054cf;
      16940: inst = 32'h8220000;
      16941: inst = 32'h10408000;
      16942: inst = 32'hc4054d0;
      16943: inst = 32'h8220000;
      16944: inst = 32'h10408000;
      16945: inst = 32'hc4054d1;
      16946: inst = 32'h8220000;
      16947: inst = 32'h10408000;
      16948: inst = 32'hc4054d2;
      16949: inst = 32'h8220000;
      16950: inst = 32'h10408000;
      16951: inst = 32'hc4054d3;
      16952: inst = 32'h8220000;
      16953: inst = 32'h10408000;
      16954: inst = 32'hc4054d4;
      16955: inst = 32'h8220000;
      16956: inst = 32'h10408000;
      16957: inst = 32'hc4054d5;
      16958: inst = 32'h8220000;
      16959: inst = 32'h10408000;
      16960: inst = 32'hc4054d6;
      16961: inst = 32'h8220000;
      16962: inst = 32'h10408000;
      16963: inst = 32'hc4054d7;
      16964: inst = 32'h8220000;
      16965: inst = 32'h10408000;
      16966: inst = 32'hc4054d8;
      16967: inst = 32'h8220000;
      16968: inst = 32'h10408000;
      16969: inst = 32'hc4054d9;
      16970: inst = 32'h8220000;
      16971: inst = 32'h10408000;
      16972: inst = 32'hc4054da;
      16973: inst = 32'h8220000;
      16974: inst = 32'h10408000;
      16975: inst = 32'hc4054db;
      16976: inst = 32'h8220000;
      16977: inst = 32'h10408000;
      16978: inst = 32'hc4054dc;
      16979: inst = 32'h8220000;
      16980: inst = 32'h10408000;
      16981: inst = 32'hc4054dd;
      16982: inst = 32'h8220000;
      16983: inst = 32'h10408000;
      16984: inst = 32'hc4054de;
      16985: inst = 32'h8220000;
      16986: inst = 32'h10408000;
      16987: inst = 32'hc4054df;
      16988: inst = 32'h8220000;
      16989: inst = 32'h10408000;
      16990: inst = 32'hc4054e0;
      16991: inst = 32'h8220000;
      16992: inst = 32'h10408000;
      16993: inst = 32'hc4054e1;
      16994: inst = 32'h8220000;
      16995: inst = 32'h10408000;
      16996: inst = 32'hc4054e2;
      16997: inst = 32'h8220000;
      16998: inst = 32'h10408000;
      16999: inst = 32'hc4054e3;
      17000: inst = 32'h8220000;
      17001: inst = 32'h10408000;
      17002: inst = 32'hc4054e4;
      17003: inst = 32'h8220000;
      17004: inst = 32'h10408000;
      17005: inst = 32'hc4054e5;
      17006: inst = 32'h8220000;
      17007: inst = 32'h10408000;
      17008: inst = 32'hc4054e6;
      17009: inst = 32'h8220000;
      17010: inst = 32'h10408000;
      17011: inst = 32'hc4054e7;
      17012: inst = 32'h8220000;
      17013: inst = 32'h10408000;
      17014: inst = 32'hc4054e8;
      17015: inst = 32'h8220000;
      17016: inst = 32'h10408000;
      17017: inst = 32'hc4054e9;
      17018: inst = 32'h8220000;
      17019: inst = 32'h10408000;
      17020: inst = 32'hc4054ea;
      17021: inst = 32'h8220000;
      17022: inst = 32'h10408000;
      17023: inst = 32'hc4054eb;
      17024: inst = 32'h8220000;
      17025: inst = 32'h10408000;
      17026: inst = 32'hc4054ec;
      17027: inst = 32'h8220000;
      17028: inst = 32'h10408000;
      17029: inst = 32'hc4054ed;
      17030: inst = 32'h8220000;
      17031: inst = 32'h10408000;
      17032: inst = 32'hc4054ee;
      17033: inst = 32'h8220000;
      17034: inst = 32'h10408000;
      17035: inst = 32'hc4054ef;
      17036: inst = 32'h8220000;
      17037: inst = 32'h10408000;
      17038: inst = 32'hc4054f0;
      17039: inst = 32'h8220000;
      17040: inst = 32'h10408000;
      17041: inst = 32'hc4054f1;
      17042: inst = 32'h8220000;
      17043: inst = 32'h10408000;
      17044: inst = 32'hc4054f2;
      17045: inst = 32'h8220000;
      17046: inst = 32'h10408000;
      17047: inst = 32'hc4054f3;
      17048: inst = 32'h8220000;
      17049: inst = 32'h10408000;
      17050: inst = 32'hc4054f4;
      17051: inst = 32'h8220000;
      17052: inst = 32'h10408000;
      17053: inst = 32'hc4054f5;
      17054: inst = 32'h8220000;
      17055: inst = 32'h10408000;
      17056: inst = 32'hc4054f6;
      17057: inst = 32'h8220000;
      17058: inst = 32'h10408000;
      17059: inst = 32'hc40550a;
      17060: inst = 32'h8220000;
      17061: inst = 32'h10408000;
      17062: inst = 32'hc40550b;
      17063: inst = 32'h8220000;
      17064: inst = 32'h10408000;
      17065: inst = 32'hc40550c;
      17066: inst = 32'h8220000;
      17067: inst = 32'h10408000;
      17068: inst = 32'hc40550d;
      17069: inst = 32'h8220000;
      17070: inst = 32'h10408000;
      17071: inst = 32'hc40550e;
      17072: inst = 32'h8220000;
      17073: inst = 32'h10408000;
      17074: inst = 32'hc40550f;
      17075: inst = 32'h8220000;
      17076: inst = 32'h10408000;
      17077: inst = 32'hc405510;
      17078: inst = 32'h8220000;
      17079: inst = 32'h10408000;
      17080: inst = 32'hc405511;
      17081: inst = 32'h8220000;
      17082: inst = 32'h10408000;
      17083: inst = 32'hc405512;
      17084: inst = 32'h8220000;
      17085: inst = 32'h10408000;
      17086: inst = 32'hc405513;
      17087: inst = 32'h8220000;
      17088: inst = 32'h10408000;
      17089: inst = 32'hc405514;
      17090: inst = 32'h8220000;
      17091: inst = 32'h10408000;
      17092: inst = 32'hc405515;
      17093: inst = 32'h8220000;
      17094: inst = 32'h10408000;
      17095: inst = 32'hc405529;
      17096: inst = 32'h8220000;
      17097: inst = 32'h10408000;
      17098: inst = 32'hc40552a;
      17099: inst = 32'h8220000;
      17100: inst = 32'h10408000;
      17101: inst = 32'hc40552b;
      17102: inst = 32'h8220000;
      17103: inst = 32'h10408000;
      17104: inst = 32'hc40552c;
      17105: inst = 32'h8220000;
      17106: inst = 32'h10408000;
      17107: inst = 32'hc40552d;
      17108: inst = 32'h8220000;
      17109: inst = 32'h10408000;
      17110: inst = 32'hc40552e;
      17111: inst = 32'h8220000;
      17112: inst = 32'h10408000;
      17113: inst = 32'hc40552f;
      17114: inst = 32'h8220000;
      17115: inst = 32'h10408000;
      17116: inst = 32'hc405530;
      17117: inst = 32'h8220000;
      17118: inst = 32'h10408000;
      17119: inst = 32'hc405531;
      17120: inst = 32'h8220000;
      17121: inst = 32'h10408000;
      17122: inst = 32'hc405532;
      17123: inst = 32'h8220000;
      17124: inst = 32'h10408000;
      17125: inst = 32'hc405533;
      17126: inst = 32'h8220000;
      17127: inst = 32'h10408000;
      17128: inst = 32'hc405534;
      17129: inst = 32'h8220000;
      17130: inst = 32'h10408000;
      17131: inst = 32'hc405535;
      17132: inst = 32'h8220000;
      17133: inst = 32'h10408000;
      17134: inst = 32'hc405536;
      17135: inst = 32'h8220000;
      17136: inst = 32'h10408000;
      17137: inst = 32'hc405537;
      17138: inst = 32'h8220000;
      17139: inst = 32'h10408000;
      17140: inst = 32'hc405538;
      17141: inst = 32'h8220000;
      17142: inst = 32'h10408000;
      17143: inst = 32'hc405539;
      17144: inst = 32'h8220000;
      17145: inst = 32'h10408000;
      17146: inst = 32'hc40553a;
      17147: inst = 32'h8220000;
      17148: inst = 32'h10408000;
      17149: inst = 32'hc40553b;
      17150: inst = 32'h8220000;
      17151: inst = 32'h10408000;
      17152: inst = 32'hc40553c;
      17153: inst = 32'h8220000;
      17154: inst = 32'h10408000;
      17155: inst = 32'hc40553d;
      17156: inst = 32'h8220000;
      17157: inst = 32'h10408000;
      17158: inst = 32'hc40553e;
      17159: inst = 32'h8220000;
      17160: inst = 32'h10408000;
      17161: inst = 32'hc40553f;
      17162: inst = 32'h8220000;
      17163: inst = 32'h10408000;
      17164: inst = 32'hc405540;
      17165: inst = 32'h8220000;
      17166: inst = 32'h10408000;
      17167: inst = 32'hc405541;
      17168: inst = 32'h8220000;
      17169: inst = 32'h10408000;
      17170: inst = 32'hc405542;
      17171: inst = 32'h8220000;
      17172: inst = 32'h10408000;
      17173: inst = 32'hc405543;
      17174: inst = 32'h8220000;
      17175: inst = 32'h10408000;
      17176: inst = 32'hc405544;
      17177: inst = 32'h8220000;
      17178: inst = 32'h10408000;
      17179: inst = 32'hc405545;
      17180: inst = 32'h8220000;
      17181: inst = 32'h10408000;
      17182: inst = 32'hc405546;
      17183: inst = 32'h8220000;
      17184: inst = 32'h10408000;
      17185: inst = 32'hc405547;
      17186: inst = 32'h8220000;
      17187: inst = 32'h10408000;
      17188: inst = 32'hc405548;
      17189: inst = 32'h8220000;
      17190: inst = 32'h10408000;
      17191: inst = 32'hc405549;
      17192: inst = 32'h8220000;
      17193: inst = 32'h10408000;
      17194: inst = 32'hc40554a;
      17195: inst = 32'h8220000;
      17196: inst = 32'h10408000;
      17197: inst = 32'hc40554b;
      17198: inst = 32'h8220000;
      17199: inst = 32'h10408000;
      17200: inst = 32'hc40554c;
      17201: inst = 32'h8220000;
      17202: inst = 32'h10408000;
      17203: inst = 32'hc40554d;
      17204: inst = 32'h8220000;
      17205: inst = 32'h10408000;
      17206: inst = 32'hc40554e;
      17207: inst = 32'h8220000;
      17208: inst = 32'h10408000;
      17209: inst = 32'hc40554f;
      17210: inst = 32'h8220000;
      17211: inst = 32'h10408000;
      17212: inst = 32'hc405550;
      17213: inst = 32'h8220000;
      17214: inst = 32'h10408000;
      17215: inst = 32'hc405551;
      17216: inst = 32'h8220000;
      17217: inst = 32'h10408000;
      17218: inst = 32'hc405552;
      17219: inst = 32'h8220000;
      17220: inst = 32'h10408000;
      17221: inst = 32'hc405553;
      17222: inst = 32'h8220000;
      17223: inst = 32'h10408000;
      17224: inst = 32'hc405554;
      17225: inst = 32'h8220000;
      17226: inst = 32'h10408000;
      17227: inst = 32'hc405555;
      17228: inst = 32'h8220000;
      17229: inst = 32'h10408000;
      17230: inst = 32'hc40556a;
      17231: inst = 32'h8220000;
      17232: inst = 32'h10408000;
      17233: inst = 32'hc40556b;
      17234: inst = 32'h8220000;
      17235: inst = 32'h10408000;
      17236: inst = 32'hc40556c;
      17237: inst = 32'h8220000;
      17238: inst = 32'h10408000;
      17239: inst = 32'hc40556d;
      17240: inst = 32'h8220000;
      17241: inst = 32'h10408000;
      17242: inst = 32'hc40556e;
      17243: inst = 32'h8220000;
      17244: inst = 32'h10408000;
      17245: inst = 32'hc40556f;
      17246: inst = 32'h8220000;
      17247: inst = 32'h10408000;
      17248: inst = 32'hc405570;
      17249: inst = 32'h8220000;
      17250: inst = 32'h10408000;
      17251: inst = 32'hc405571;
      17252: inst = 32'h8220000;
      17253: inst = 32'h10408000;
      17254: inst = 32'hc405572;
      17255: inst = 32'h8220000;
      17256: inst = 32'h10408000;
      17257: inst = 32'hc405573;
      17258: inst = 32'h8220000;
      17259: inst = 32'h10408000;
      17260: inst = 32'hc405574;
      17261: inst = 32'h8220000;
      17262: inst = 32'h10408000;
      17263: inst = 32'hc405575;
      17264: inst = 32'h8220000;
      17265: inst = 32'h10408000;
      17266: inst = 32'hc40558a;
      17267: inst = 32'h8220000;
      17268: inst = 32'h10408000;
      17269: inst = 32'hc40558b;
      17270: inst = 32'h8220000;
      17271: inst = 32'h10408000;
      17272: inst = 32'hc40558c;
      17273: inst = 32'h8220000;
      17274: inst = 32'h10408000;
      17275: inst = 32'hc40558d;
      17276: inst = 32'h8220000;
      17277: inst = 32'h10408000;
      17278: inst = 32'hc40558e;
      17279: inst = 32'h8220000;
      17280: inst = 32'h10408000;
      17281: inst = 32'hc40558f;
      17282: inst = 32'h8220000;
      17283: inst = 32'h10408000;
      17284: inst = 32'hc405590;
      17285: inst = 32'h8220000;
      17286: inst = 32'h10408000;
      17287: inst = 32'hc405591;
      17288: inst = 32'h8220000;
      17289: inst = 32'h10408000;
      17290: inst = 32'hc405592;
      17291: inst = 32'h8220000;
      17292: inst = 32'h10408000;
      17293: inst = 32'hc405593;
      17294: inst = 32'h8220000;
      17295: inst = 32'h10408000;
      17296: inst = 32'hc405594;
      17297: inst = 32'h8220000;
      17298: inst = 32'h10408000;
      17299: inst = 32'hc405595;
      17300: inst = 32'h8220000;
      17301: inst = 32'h10408000;
      17302: inst = 32'hc405596;
      17303: inst = 32'h8220000;
      17304: inst = 32'h10408000;
      17305: inst = 32'hc405597;
      17306: inst = 32'h8220000;
      17307: inst = 32'h10408000;
      17308: inst = 32'hc405598;
      17309: inst = 32'h8220000;
      17310: inst = 32'h10408000;
      17311: inst = 32'hc405599;
      17312: inst = 32'h8220000;
      17313: inst = 32'h10408000;
      17314: inst = 32'hc40559a;
      17315: inst = 32'h8220000;
      17316: inst = 32'h10408000;
      17317: inst = 32'hc40559b;
      17318: inst = 32'h8220000;
      17319: inst = 32'h10408000;
      17320: inst = 32'hc40559c;
      17321: inst = 32'h8220000;
      17322: inst = 32'h10408000;
      17323: inst = 32'hc40559d;
      17324: inst = 32'h8220000;
      17325: inst = 32'h10408000;
      17326: inst = 32'hc40559e;
      17327: inst = 32'h8220000;
      17328: inst = 32'h10408000;
      17329: inst = 32'hc40559f;
      17330: inst = 32'h8220000;
      17331: inst = 32'h10408000;
      17332: inst = 32'hc4055a0;
      17333: inst = 32'h8220000;
      17334: inst = 32'h10408000;
      17335: inst = 32'hc4055a1;
      17336: inst = 32'h8220000;
      17337: inst = 32'h10408000;
      17338: inst = 32'hc4055a2;
      17339: inst = 32'h8220000;
      17340: inst = 32'h10408000;
      17341: inst = 32'hc4055a3;
      17342: inst = 32'h8220000;
      17343: inst = 32'h10408000;
      17344: inst = 32'hc4055a4;
      17345: inst = 32'h8220000;
      17346: inst = 32'h10408000;
      17347: inst = 32'hc4055a5;
      17348: inst = 32'h8220000;
      17349: inst = 32'h10408000;
      17350: inst = 32'hc4055a6;
      17351: inst = 32'h8220000;
      17352: inst = 32'h10408000;
      17353: inst = 32'hc4055a7;
      17354: inst = 32'h8220000;
      17355: inst = 32'h10408000;
      17356: inst = 32'hc4055a8;
      17357: inst = 32'h8220000;
      17358: inst = 32'h10408000;
      17359: inst = 32'hc4055a9;
      17360: inst = 32'h8220000;
      17361: inst = 32'h10408000;
      17362: inst = 32'hc4055aa;
      17363: inst = 32'h8220000;
      17364: inst = 32'h10408000;
      17365: inst = 32'hc4055ab;
      17366: inst = 32'h8220000;
      17367: inst = 32'h10408000;
      17368: inst = 32'hc4055ac;
      17369: inst = 32'h8220000;
      17370: inst = 32'h10408000;
      17371: inst = 32'hc4055ad;
      17372: inst = 32'h8220000;
      17373: inst = 32'h10408000;
      17374: inst = 32'hc4055ae;
      17375: inst = 32'h8220000;
      17376: inst = 32'h10408000;
      17377: inst = 32'hc4055af;
      17378: inst = 32'h8220000;
      17379: inst = 32'h10408000;
      17380: inst = 32'hc4055b0;
      17381: inst = 32'h8220000;
      17382: inst = 32'h10408000;
      17383: inst = 32'hc4055b1;
      17384: inst = 32'h8220000;
      17385: inst = 32'h10408000;
      17386: inst = 32'hc4055b2;
      17387: inst = 32'h8220000;
      17388: inst = 32'h10408000;
      17389: inst = 32'hc4055b3;
      17390: inst = 32'h8220000;
      17391: inst = 32'h10408000;
      17392: inst = 32'hc4055b4;
      17393: inst = 32'h8220000;
      17394: inst = 32'h10408000;
      17395: inst = 32'hc4055ca;
      17396: inst = 32'h8220000;
      17397: inst = 32'h10408000;
      17398: inst = 32'hc4055cb;
      17399: inst = 32'h8220000;
      17400: inst = 32'h10408000;
      17401: inst = 32'hc4055cc;
      17402: inst = 32'h8220000;
      17403: inst = 32'h10408000;
      17404: inst = 32'hc4055cd;
      17405: inst = 32'h8220000;
      17406: inst = 32'h10408000;
      17407: inst = 32'hc4055ce;
      17408: inst = 32'h8220000;
      17409: inst = 32'h10408000;
      17410: inst = 32'hc4055cf;
      17411: inst = 32'h8220000;
      17412: inst = 32'h10408000;
      17413: inst = 32'hc4055d0;
      17414: inst = 32'h8220000;
      17415: inst = 32'h10408000;
      17416: inst = 32'hc4055d1;
      17417: inst = 32'h8220000;
      17418: inst = 32'h10408000;
      17419: inst = 32'hc4055d2;
      17420: inst = 32'h8220000;
      17421: inst = 32'h10408000;
      17422: inst = 32'hc4055d3;
      17423: inst = 32'h8220000;
      17424: inst = 32'h10408000;
      17425: inst = 32'hc4055d4;
      17426: inst = 32'h8220000;
      17427: inst = 32'h10408000;
      17428: inst = 32'hc4055d5;
      17429: inst = 32'h8220000;
      17430: inst = 32'h10408000;
      17431: inst = 32'hc4055eb;
      17432: inst = 32'h8220000;
      17433: inst = 32'h10408000;
      17434: inst = 32'hc4055ec;
      17435: inst = 32'h8220000;
      17436: inst = 32'h10408000;
      17437: inst = 32'hc4055ed;
      17438: inst = 32'h8220000;
      17439: inst = 32'h10408000;
      17440: inst = 32'hc4055ee;
      17441: inst = 32'h8220000;
      17442: inst = 32'h10408000;
      17443: inst = 32'hc4055ef;
      17444: inst = 32'h8220000;
      17445: inst = 32'h10408000;
      17446: inst = 32'hc4055f0;
      17447: inst = 32'h8220000;
      17448: inst = 32'h10408000;
      17449: inst = 32'hc4055f1;
      17450: inst = 32'h8220000;
      17451: inst = 32'h10408000;
      17452: inst = 32'hc4055f2;
      17453: inst = 32'h8220000;
      17454: inst = 32'h10408000;
      17455: inst = 32'hc4055f3;
      17456: inst = 32'h8220000;
      17457: inst = 32'h10408000;
      17458: inst = 32'hc4055f4;
      17459: inst = 32'h8220000;
      17460: inst = 32'h10408000;
      17461: inst = 32'hc4055f5;
      17462: inst = 32'h8220000;
      17463: inst = 32'h10408000;
      17464: inst = 32'hc4055f6;
      17465: inst = 32'h8220000;
      17466: inst = 32'h10408000;
      17467: inst = 32'hc4055f7;
      17468: inst = 32'h8220000;
      17469: inst = 32'h10408000;
      17470: inst = 32'hc4055f8;
      17471: inst = 32'h8220000;
      17472: inst = 32'h10408000;
      17473: inst = 32'hc4055f9;
      17474: inst = 32'h8220000;
      17475: inst = 32'h10408000;
      17476: inst = 32'hc4055fa;
      17477: inst = 32'h8220000;
      17478: inst = 32'h10408000;
      17479: inst = 32'hc4055fb;
      17480: inst = 32'h8220000;
      17481: inst = 32'h10408000;
      17482: inst = 32'hc4055fc;
      17483: inst = 32'h8220000;
      17484: inst = 32'h10408000;
      17485: inst = 32'hc4055fd;
      17486: inst = 32'h8220000;
      17487: inst = 32'h10408000;
      17488: inst = 32'hc4055fe;
      17489: inst = 32'h8220000;
      17490: inst = 32'h10408000;
      17491: inst = 32'hc4055ff;
      17492: inst = 32'h8220000;
      17493: inst = 32'h10408000;
      17494: inst = 32'hc405600;
      17495: inst = 32'h8220000;
      17496: inst = 32'h10408000;
      17497: inst = 32'hc405601;
      17498: inst = 32'h8220000;
      17499: inst = 32'h10408000;
      17500: inst = 32'hc405602;
      17501: inst = 32'h8220000;
      17502: inst = 32'h10408000;
      17503: inst = 32'hc405603;
      17504: inst = 32'h8220000;
      17505: inst = 32'h10408000;
      17506: inst = 32'hc405604;
      17507: inst = 32'h8220000;
      17508: inst = 32'h10408000;
      17509: inst = 32'hc405605;
      17510: inst = 32'h8220000;
      17511: inst = 32'h10408000;
      17512: inst = 32'hc405606;
      17513: inst = 32'h8220000;
      17514: inst = 32'h10408000;
      17515: inst = 32'hc405607;
      17516: inst = 32'h8220000;
      17517: inst = 32'h10408000;
      17518: inst = 32'hc405608;
      17519: inst = 32'h8220000;
      17520: inst = 32'h10408000;
      17521: inst = 32'hc405609;
      17522: inst = 32'h8220000;
      17523: inst = 32'h10408000;
      17524: inst = 32'hc40560a;
      17525: inst = 32'h8220000;
      17526: inst = 32'h10408000;
      17527: inst = 32'hc40560b;
      17528: inst = 32'h8220000;
      17529: inst = 32'h10408000;
      17530: inst = 32'hc40560c;
      17531: inst = 32'h8220000;
      17532: inst = 32'h10408000;
      17533: inst = 32'hc40560d;
      17534: inst = 32'h8220000;
      17535: inst = 32'h10408000;
      17536: inst = 32'hc40560e;
      17537: inst = 32'h8220000;
      17538: inst = 32'h10408000;
      17539: inst = 32'hc40560f;
      17540: inst = 32'h8220000;
      17541: inst = 32'h10408000;
      17542: inst = 32'hc405610;
      17543: inst = 32'h8220000;
      17544: inst = 32'h10408000;
      17545: inst = 32'hc405611;
      17546: inst = 32'h8220000;
      17547: inst = 32'h10408000;
      17548: inst = 32'hc405612;
      17549: inst = 32'h8220000;
      17550: inst = 32'h10408000;
      17551: inst = 32'hc405613;
      17552: inst = 32'h8220000;
      17553: inst = 32'h10408000;
      17554: inst = 32'hc405614;
      17555: inst = 32'h8220000;
      17556: inst = 32'h10408000;
      17557: inst = 32'hc40562a;
      17558: inst = 32'h8220000;
      17559: inst = 32'h10408000;
      17560: inst = 32'hc40562b;
      17561: inst = 32'h8220000;
      17562: inst = 32'h10408000;
      17563: inst = 32'hc40562c;
      17564: inst = 32'h8220000;
      17565: inst = 32'h10408000;
      17566: inst = 32'hc40562d;
      17567: inst = 32'h8220000;
      17568: inst = 32'h10408000;
      17569: inst = 32'hc40562e;
      17570: inst = 32'h8220000;
      17571: inst = 32'h10408000;
      17572: inst = 32'hc40562f;
      17573: inst = 32'h8220000;
      17574: inst = 32'h10408000;
      17575: inst = 32'hc405630;
      17576: inst = 32'h8220000;
      17577: inst = 32'h10408000;
      17578: inst = 32'hc405631;
      17579: inst = 32'h8220000;
      17580: inst = 32'h10408000;
      17581: inst = 32'hc405632;
      17582: inst = 32'h8220000;
      17583: inst = 32'h10408000;
      17584: inst = 32'hc405633;
      17585: inst = 32'h8220000;
      17586: inst = 32'h10408000;
      17587: inst = 32'hc405634;
      17588: inst = 32'h8220000;
      17589: inst = 32'h10408000;
      17590: inst = 32'hc405635;
      17591: inst = 32'h8220000;
      17592: inst = 32'h10408000;
      17593: inst = 32'hc40564b;
      17594: inst = 32'h8220000;
      17595: inst = 32'h10408000;
      17596: inst = 32'hc40564c;
      17597: inst = 32'h8220000;
      17598: inst = 32'h10408000;
      17599: inst = 32'hc40564d;
      17600: inst = 32'h8220000;
      17601: inst = 32'h10408000;
      17602: inst = 32'hc40564e;
      17603: inst = 32'h8220000;
      17604: inst = 32'h10408000;
      17605: inst = 32'hc40564f;
      17606: inst = 32'h8220000;
      17607: inst = 32'h10408000;
      17608: inst = 32'hc405650;
      17609: inst = 32'h8220000;
      17610: inst = 32'h10408000;
      17611: inst = 32'hc405651;
      17612: inst = 32'h8220000;
      17613: inst = 32'h10408000;
      17614: inst = 32'hc405652;
      17615: inst = 32'h8220000;
      17616: inst = 32'h10408000;
      17617: inst = 32'hc405653;
      17618: inst = 32'h8220000;
      17619: inst = 32'h10408000;
      17620: inst = 32'hc405654;
      17621: inst = 32'h8220000;
      17622: inst = 32'h10408000;
      17623: inst = 32'hc405655;
      17624: inst = 32'h8220000;
      17625: inst = 32'h10408000;
      17626: inst = 32'hc405656;
      17627: inst = 32'h8220000;
      17628: inst = 32'h10408000;
      17629: inst = 32'hc405657;
      17630: inst = 32'h8220000;
      17631: inst = 32'h10408000;
      17632: inst = 32'hc405658;
      17633: inst = 32'h8220000;
      17634: inst = 32'h10408000;
      17635: inst = 32'hc405659;
      17636: inst = 32'h8220000;
      17637: inst = 32'h10408000;
      17638: inst = 32'hc40565a;
      17639: inst = 32'h8220000;
      17640: inst = 32'h10408000;
      17641: inst = 32'hc40565b;
      17642: inst = 32'h8220000;
      17643: inst = 32'h10408000;
      17644: inst = 32'hc40565c;
      17645: inst = 32'h8220000;
      17646: inst = 32'h10408000;
      17647: inst = 32'hc40565d;
      17648: inst = 32'h8220000;
      17649: inst = 32'h10408000;
      17650: inst = 32'hc40565e;
      17651: inst = 32'h8220000;
      17652: inst = 32'h10408000;
      17653: inst = 32'hc40565f;
      17654: inst = 32'h8220000;
      17655: inst = 32'h10408000;
      17656: inst = 32'hc405660;
      17657: inst = 32'h8220000;
      17658: inst = 32'h10408000;
      17659: inst = 32'hc405661;
      17660: inst = 32'h8220000;
      17661: inst = 32'h10408000;
      17662: inst = 32'hc405662;
      17663: inst = 32'h8220000;
      17664: inst = 32'h10408000;
      17665: inst = 32'hc405663;
      17666: inst = 32'h8220000;
      17667: inst = 32'h10408000;
      17668: inst = 32'hc405664;
      17669: inst = 32'h8220000;
      17670: inst = 32'h10408000;
      17671: inst = 32'hc405665;
      17672: inst = 32'h8220000;
      17673: inst = 32'h10408000;
      17674: inst = 32'hc405666;
      17675: inst = 32'h8220000;
      17676: inst = 32'h10408000;
      17677: inst = 32'hc405667;
      17678: inst = 32'h8220000;
      17679: inst = 32'h10408000;
      17680: inst = 32'hc405668;
      17681: inst = 32'h8220000;
      17682: inst = 32'h10408000;
      17683: inst = 32'hc405669;
      17684: inst = 32'h8220000;
      17685: inst = 32'h10408000;
      17686: inst = 32'hc40566a;
      17687: inst = 32'h8220000;
      17688: inst = 32'h10408000;
      17689: inst = 32'hc40566b;
      17690: inst = 32'h8220000;
      17691: inst = 32'h10408000;
      17692: inst = 32'hc40566c;
      17693: inst = 32'h8220000;
      17694: inst = 32'h10408000;
      17695: inst = 32'hc40566d;
      17696: inst = 32'h8220000;
      17697: inst = 32'h10408000;
      17698: inst = 32'hc40566e;
      17699: inst = 32'h8220000;
      17700: inst = 32'h10408000;
      17701: inst = 32'hc40566f;
      17702: inst = 32'h8220000;
      17703: inst = 32'h10408000;
      17704: inst = 32'hc405670;
      17705: inst = 32'h8220000;
      17706: inst = 32'h10408000;
      17707: inst = 32'hc405671;
      17708: inst = 32'h8220000;
      17709: inst = 32'h10408000;
      17710: inst = 32'hc405672;
      17711: inst = 32'h8220000;
      17712: inst = 32'h10408000;
      17713: inst = 32'hc405673;
      17714: inst = 32'h8220000;
      17715: inst = 32'h10408000;
      17716: inst = 32'hc40568a;
      17717: inst = 32'h8220000;
      17718: inst = 32'h10408000;
      17719: inst = 32'hc40568b;
      17720: inst = 32'h8220000;
      17721: inst = 32'h10408000;
      17722: inst = 32'hc40568c;
      17723: inst = 32'h8220000;
      17724: inst = 32'h10408000;
      17725: inst = 32'hc40568d;
      17726: inst = 32'h8220000;
      17727: inst = 32'h10408000;
      17728: inst = 32'hc40568e;
      17729: inst = 32'h8220000;
      17730: inst = 32'h10408000;
      17731: inst = 32'hc40568f;
      17732: inst = 32'h8220000;
      17733: inst = 32'h10408000;
      17734: inst = 32'hc405690;
      17735: inst = 32'h8220000;
      17736: inst = 32'h10408000;
      17737: inst = 32'hc405691;
      17738: inst = 32'h8220000;
      17739: inst = 32'h10408000;
      17740: inst = 32'hc405692;
      17741: inst = 32'h8220000;
      17742: inst = 32'h10408000;
      17743: inst = 32'hc405693;
      17744: inst = 32'h8220000;
      17745: inst = 32'h10408000;
      17746: inst = 32'hc405694;
      17747: inst = 32'h8220000;
      17748: inst = 32'h10408000;
      17749: inst = 32'hc405695;
      17750: inst = 32'h8220000;
      17751: inst = 32'h10408000;
      17752: inst = 32'hc4056ac;
      17753: inst = 32'h8220000;
      17754: inst = 32'h10408000;
      17755: inst = 32'hc4056ad;
      17756: inst = 32'h8220000;
      17757: inst = 32'h10408000;
      17758: inst = 32'hc4056ae;
      17759: inst = 32'h8220000;
      17760: inst = 32'h10408000;
      17761: inst = 32'hc4056af;
      17762: inst = 32'h8220000;
      17763: inst = 32'h10408000;
      17764: inst = 32'hc4056b0;
      17765: inst = 32'h8220000;
      17766: inst = 32'h10408000;
      17767: inst = 32'hc4056b1;
      17768: inst = 32'h8220000;
      17769: inst = 32'h10408000;
      17770: inst = 32'hc4056b2;
      17771: inst = 32'h8220000;
      17772: inst = 32'h10408000;
      17773: inst = 32'hc4056b3;
      17774: inst = 32'h8220000;
      17775: inst = 32'h10408000;
      17776: inst = 32'hc4056b4;
      17777: inst = 32'h8220000;
      17778: inst = 32'h10408000;
      17779: inst = 32'hc4056b5;
      17780: inst = 32'h8220000;
      17781: inst = 32'h10408000;
      17782: inst = 32'hc4056b6;
      17783: inst = 32'h8220000;
      17784: inst = 32'h10408000;
      17785: inst = 32'hc4056b7;
      17786: inst = 32'h8220000;
      17787: inst = 32'h10408000;
      17788: inst = 32'hc4056b8;
      17789: inst = 32'h8220000;
      17790: inst = 32'h10408000;
      17791: inst = 32'hc4056b9;
      17792: inst = 32'h8220000;
      17793: inst = 32'h10408000;
      17794: inst = 32'hc4056ba;
      17795: inst = 32'h8220000;
      17796: inst = 32'h10408000;
      17797: inst = 32'hc4056bb;
      17798: inst = 32'h8220000;
      17799: inst = 32'h10408000;
      17800: inst = 32'hc4056bc;
      17801: inst = 32'h8220000;
      17802: inst = 32'h10408000;
      17803: inst = 32'hc4056bd;
      17804: inst = 32'h8220000;
      17805: inst = 32'h10408000;
      17806: inst = 32'hc4056be;
      17807: inst = 32'h8220000;
      17808: inst = 32'h10408000;
      17809: inst = 32'hc4056bf;
      17810: inst = 32'h8220000;
      17811: inst = 32'h10408000;
      17812: inst = 32'hc4056c0;
      17813: inst = 32'h8220000;
      17814: inst = 32'h10408000;
      17815: inst = 32'hc4056c1;
      17816: inst = 32'h8220000;
      17817: inst = 32'h10408000;
      17818: inst = 32'hc4056c2;
      17819: inst = 32'h8220000;
      17820: inst = 32'h10408000;
      17821: inst = 32'hc4056c3;
      17822: inst = 32'h8220000;
      17823: inst = 32'h10408000;
      17824: inst = 32'hc4056c4;
      17825: inst = 32'h8220000;
      17826: inst = 32'h10408000;
      17827: inst = 32'hc4056c5;
      17828: inst = 32'h8220000;
      17829: inst = 32'h10408000;
      17830: inst = 32'hc4056c6;
      17831: inst = 32'h8220000;
      17832: inst = 32'h10408000;
      17833: inst = 32'hc4056c7;
      17834: inst = 32'h8220000;
      17835: inst = 32'h10408000;
      17836: inst = 32'hc4056c8;
      17837: inst = 32'h8220000;
      17838: inst = 32'h10408000;
      17839: inst = 32'hc4056c9;
      17840: inst = 32'h8220000;
      17841: inst = 32'h10408000;
      17842: inst = 32'hc4056ca;
      17843: inst = 32'h8220000;
      17844: inst = 32'h10408000;
      17845: inst = 32'hc4056cb;
      17846: inst = 32'h8220000;
      17847: inst = 32'h10408000;
      17848: inst = 32'hc4056cc;
      17849: inst = 32'h8220000;
      17850: inst = 32'h10408000;
      17851: inst = 32'hc4056cd;
      17852: inst = 32'h8220000;
      17853: inst = 32'h10408000;
      17854: inst = 32'hc4056ce;
      17855: inst = 32'h8220000;
      17856: inst = 32'h10408000;
      17857: inst = 32'hc4056cf;
      17858: inst = 32'h8220000;
      17859: inst = 32'h10408000;
      17860: inst = 32'hc4056d0;
      17861: inst = 32'h8220000;
      17862: inst = 32'h10408000;
      17863: inst = 32'hc4056d1;
      17864: inst = 32'h8220000;
      17865: inst = 32'h10408000;
      17866: inst = 32'hc4056d2;
      17867: inst = 32'h8220000;
      17868: inst = 32'h10408000;
      17869: inst = 32'hc4056ea;
      17870: inst = 32'h8220000;
      17871: inst = 32'h10408000;
      17872: inst = 32'hc4056eb;
      17873: inst = 32'h8220000;
      17874: inst = 32'h10408000;
      17875: inst = 32'hc4056ec;
      17876: inst = 32'h8220000;
      17877: inst = 32'h10408000;
      17878: inst = 32'hc4056ed;
      17879: inst = 32'h8220000;
      17880: inst = 32'h10408000;
      17881: inst = 32'hc4056ee;
      17882: inst = 32'h8220000;
      17883: inst = 32'h10408000;
      17884: inst = 32'hc4056ef;
      17885: inst = 32'h8220000;
      17886: inst = 32'h10408000;
      17887: inst = 32'hc4056f0;
      17888: inst = 32'h8220000;
      17889: inst = 32'h10408000;
      17890: inst = 32'hc4056f1;
      17891: inst = 32'h8220000;
      17892: inst = 32'h10408000;
      17893: inst = 32'hc4056f2;
      17894: inst = 32'h8220000;
      17895: inst = 32'h10408000;
      17896: inst = 32'hc4056f3;
      17897: inst = 32'h8220000;
      17898: inst = 32'h10408000;
      17899: inst = 32'hc4056f4;
      17900: inst = 32'h8220000;
      17901: inst = 32'h10408000;
      17902: inst = 32'hc4056f5;
      17903: inst = 32'h8220000;
      17904: inst = 32'h10408000;
      17905: inst = 32'hc40570d;
      17906: inst = 32'h8220000;
      17907: inst = 32'h10408000;
      17908: inst = 32'hc40570e;
      17909: inst = 32'h8220000;
      17910: inst = 32'h10408000;
      17911: inst = 32'hc40570f;
      17912: inst = 32'h8220000;
      17913: inst = 32'h10408000;
      17914: inst = 32'hc405710;
      17915: inst = 32'h8220000;
      17916: inst = 32'h10408000;
      17917: inst = 32'hc405711;
      17918: inst = 32'h8220000;
      17919: inst = 32'h10408000;
      17920: inst = 32'hc405712;
      17921: inst = 32'h8220000;
      17922: inst = 32'h10408000;
      17923: inst = 32'hc405713;
      17924: inst = 32'h8220000;
      17925: inst = 32'h10408000;
      17926: inst = 32'hc405714;
      17927: inst = 32'h8220000;
      17928: inst = 32'h10408000;
      17929: inst = 32'hc405715;
      17930: inst = 32'h8220000;
      17931: inst = 32'h10408000;
      17932: inst = 32'hc405716;
      17933: inst = 32'h8220000;
      17934: inst = 32'h10408000;
      17935: inst = 32'hc405717;
      17936: inst = 32'h8220000;
      17937: inst = 32'h10408000;
      17938: inst = 32'hc405718;
      17939: inst = 32'h8220000;
      17940: inst = 32'h10408000;
      17941: inst = 32'hc405719;
      17942: inst = 32'h8220000;
      17943: inst = 32'h10408000;
      17944: inst = 32'hc40571a;
      17945: inst = 32'h8220000;
      17946: inst = 32'h10408000;
      17947: inst = 32'hc40571b;
      17948: inst = 32'h8220000;
      17949: inst = 32'h10408000;
      17950: inst = 32'hc40571c;
      17951: inst = 32'h8220000;
      17952: inst = 32'h10408000;
      17953: inst = 32'hc40571d;
      17954: inst = 32'h8220000;
      17955: inst = 32'h10408000;
      17956: inst = 32'hc40571e;
      17957: inst = 32'h8220000;
      17958: inst = 32'h10408000;
      17959: inst = 32'hc40571f;
      17960: inst = 32'h8220000;
      17961: inst = 32'h10408000;
      17962: inst = 32'hc405720;
      17963: inst = 32'h8220000;
      17964: inst = 32'h10408000;
      17965: inst = 32'hc405721;
      17966: inst = 32'h8220000;
      17967: inst = 32'h10408000;
      17968: inst = 32'hc405722;
      17969: inst = 32'h8220000;
      17970: inst = 32'h10408000;
      17971: inst = 32'hc405723;
      17972: inst = 32'h8220000;
      17973: inst = 32'h10408000;
      17974: inst = 32'hc405724;
      17975: inst = 32'h8220000;
      17976: inst = 32'h10408000;
      17977: inst = 32'hc405725;
      17978: inst = 32'h8220000;
      17979: inst = 32'h10408000;
      17980: inst = 32'hc405726;
      17981: inst = 32'h8220000;
      17982: inst = 32'h10408000;
      17983: inst = 32'hc405727;
      17984: inst = 32'h8220000;
      17985: inst = 32'h10408000;
      17986: inst = 32'hc405728;
      17987: inst = 32'h8220000;
      17988: inst = 32'h10408000;
      17989: inst = 32'hc405729;
      17990: inst = 32'h8220000;
      17991: inst = 32'h10408000;
      17992: inst = 32'hc40572a;
      17993: inst = 32'h8220000;
      17994: inst = 32'h10408000;
      17995: inst = 32'hc40572b;
      17996: inst = 32'h8220000;
      17997: inst = 32'h10408000;
      17998: inst = 32'hc40572c;
      17999: inst = 32'h8220000;
      18000: inst = 32'h10408000;
      18001: inst = 32'hc40572d;
      18002: inst = 32'h8220000;
      18003: inst = 32'h10408000;
      18004: inst = 32'hc40572e;
      18005: inst = 32'h8220000;
      18006: inst = 32'h10408000;
      18007: inst = 32'hc40572f;
      18008: inst = 32'h8220000;
      18009: inst = 32'h10408000;
      18010: inst = 32'hc405730;
      18011: inst = 32'h8220000;
      18012: inst = 32'h10408000;
      18013: inst = 32'hc405731;
      18014: inst = 32'h8220000;
      18015: inst = 32'h10408000;
      18016: inst = 32'hc40574a;
      18017: inst = 32'h8220000;
      18018: inst = 32'h10408000;
      18019: inst = 32'hc40574b;
      18020: inst = 32'h8220000;
      18021: inst = 32'h10408000;
      18022: inst = 32'hc40574c;
      18023: inst = 32'h8220000;
      18024: inst = 32'h10408000;
      18025: inst = 32'hc40574d;
      18026: inst = 32'h8220000;
      18027: inst = 32'h10408000;
      18028: inst = 32'hc40574e;
      18029: inst = 32'h8220000;
      18030: inst = 32'h10408000;
      18031: inst = 32'hc40574f;
      18032: inst = 32'h8220000;
      18033: inst = 32'h10408000;
      18034: inst = 32'hc405750;
      18035: inst = 32'h8220000;
      18036: inst = 32'h10408000;
      18037: inst = 32'hc405751;
      18038: inst = 32'h8220000;
      18039: inst = 32'h10408000;
      18040: inst = 32'hc405752;
      18041: inst = 32'h8220000;
      18042: inst = 32'h10408000;
      18043: inst = 32'hc405753;
      18044: inst = 32'h8220000;
      18045: inst = 32'h10408000;
      18046: inst = 32'hc405754;
      18047: inst = 32'h8220000;
      18048: inst = 32'h10408000;
      18049: inst = 32'hc405755;
      18050: inst = 32'h8220000;
      18051: inst = 32'h10408000;
      18052: inst = 32'hc40576e;
      18053: inst = 32'h8220000;
      18054: inst = 32'h10408000;
      18055: inst = 32'hc40576f;
      18056: inst = 32'h8220000;
      18057: inst = 32'h10408000;
      18058: inst = 32'hc405770;
      18059: inst = 32'h8220000;
      18060: inst = 32'h10408000;
      18061: inst = 32'hc405771;
      18062: inst = 32'h8220000;
      18063: inst = 32'h10408000;
      18064: inst = 32'hc405772;
      18065: inst = 32'h8220000;
      18066: inst = 32'h10408000;
      18067: inst = 32'hc405773;
      18068: inst = 32'h8220000;
      18069: inst = 32'h10408000;
      18070: inst = 32'hc405774;
      18071: inst = 32'h8220000;
      18072: inst = 32'h10408000;
      18073: inst = 32'hc405775;
      18074: inst = 32'h8220000;
      18075: inst = 32'h10408000;
      18076: inst = 32'hc405776;
      18077: inst = 32'h8220000;
      18078: inst = 32'h10408000;
      18079: inst = 32'hc405777;
      18080: inst = 32'h8220000;
      18081: inst = 32'h10408000;
      18082: inst = 32'hc405778;
      18083: inst = 32'h8220000;
      18084: inst = 32'h10408000;
      18085: inst = 32'hc405779;
      18086: inst = 32'h8220000;
      18087: inst = 32'h10408000;
      18088: inst = 32'hc40577a;
      18089: inst = 32'h8220000;
      18090: inst = 32'h10408000;
      18091: inst = 32'hc40577b;
      18092: inst = 32'h8220000;
      18093: inst = 32'h10408000;
      18094: inst = 32'hc40577c;
      18095: inst = 32'h8220000;
      18096: inst = 32'h10408000;
      18097: inst = 32'hc40577d;
      18098: inst = 32'h8220000;
      18099: inst = 32'h10408000;
      18100: inst = 32'hc40577e;
      18101: inst = 32'h8220000;
      18102: inst = 32'h10408000;
      18103: inst = 32'hc40577f;
      18104: inst = 32'h8220000;
      18105: inst = 32'h10408000;
      18106: inst = 32'hc405780;
      18107: inst = 32'h8220000;
      18108: inst = 32'h10408000;
      18109: inst = 32'hc405781;
      18110: inst = 32'h8220000;
      18111: inst = 32'h10408000;
      18112: inst = 32'hc405782;
      18113: inst = 32'h8220000;
      18114: inst = 32'h10408000;
      18115: inst = 32'hc405783;
      18116: inst = 32'h8220000;
      18117: inst = 32'h10408000;
      18118: inst = 32'hc405784;
      18119: inst = 32'h8220000;
      18120: inst = 32'h10408000;
      18121: inst = 32'hc405785;
      18122: inst = 32'h8220000;
      18123: inst = 32'h10408000;
      18124: inst = 32'hc405786;
      18125: inst = 32'h8220000;
      18126: inst = 32'h10408000;
      18127: inst = 32'hc405787;
      18128: inst = 32'h8220000;
      18129: inst = 32'h10408000;
      18130: inst = 32'hc405788;
      18131: inst = 32'h8220000;
      18132: inst = 32'h10408000;
      18133: inst = 32'hc405789;
      18134: inst = 32'h8220000;
      18135: inst = 32'h10408000;
      18136: inst = 32'hc40578a;
      18137: inst = 32'h8220000;
      18138: inst = 32'h10408000;
      18139: inst = 32'hc40578b;
      18140: inst = 32'h8220000;
      18141: inst = 32'h10408000;
      18142: inst = 32'hc40578c;
      18143: inst = 32'h8220000;
      18144: inst = 32'h10408000;
      18145: inst = 32'hc40578d;
      18146: inst = 32'h8220000;
      18147: inst = 32'h10408000;
      18148: inst = 32'hc40578e;
      18149: inst = 32'h8220000;
      18150: inst = 32'h10408000;
      18151: inst = 32'hc40578f;
      18152: inst = 32'h8220000;
      18153: inst = 32'h10408000;
      18154: inst = 32'hc405790;
      18155: inst = 32'h8220000;
      18156: inst = 32'h10408000;
      18157: inst = 32'hc405791;
      18158: inst = 32'h8220000;
      18159: inst = 32'h10408000;
      18160: inst = 32'hc4057aa;
      18161: inst = 32'h8220000;
      18162: inst = 32'h10408000;
      18163: inst = 32'hc4057ab;
      18164: inst = 32'h8220000;
      18165: inst = 32'h10408000;
      18166: inst = 32'hc4057ac;
      18167: inst = 32'h8220000;
      18168: inst = 32'h10408000;
      18169: inst = 32'hc4057ad;
      18170: inst = 32'h8220000;
      18171: inst = 32'h10408000;
      18172: inst = 32'hc4057ae;
      18173: inst = 32'h8220000;
      18174: inst = 32'h10408000;
      18175: inst = 32'hc4057af;
      18176: inst = 32'h8220000;
      18177: inst = 32'h10408000;
      18178: inst = 32'hc4057b0;
      18179: inst = 32'h8220000;
      18180: inst = 32'h10408000;
      18181: inst = 32'hc4057b1;
      18182: inst = 32'h8220000;
      18183: inst = 32'h10408000;
      18184: inst = 32'hc4057b2;
      18185: inst = 32'h8220000;
      18186: inst = 32'h10408000;
      18187: inst = 32'hc4057b3;
      18188: inst = 32'h8220000;
      18189: inst = 32'h10408000;
      18190: inst = 32'hc4057b4;
      18191: inst = 32'h8220000;
      18192: inst = 32'h10408000;
      18193: inst = 32'hc4057b5;
      18194: inst = 32'h8220000;
      18195: inst = 32'h10408000;
      18196: inst = 32'hc4057ce;
      18197: inst = 32'h8220000;
      18198: inst = 32'h10408000;
      18199: inst = 32'hc4057cf;
      18200: inst = 32'h8220000;
      18201: inst = 32'h10408000;
      18202: inst = 32'hc4057d0;
      18203: inst = 32'h8220000;
      18204: inst = 32'h10408000;
      18205: inst = 32'hc4057d1;
      18206: inst = 32'h8220000;
      18207: inst = 32'h10408000;
      18208: inst = 32'hc4057d2;
      18209: inst = 32'h8220000;
      18210: inst = 32'h10408000;
      18211: inst = 32'hc4057d3;
      18212: inst = 32'h8220000;
      18213: inst = 32'h10408000;
      18214: inst = 32'hc4057d4;
      18215: inst = 32'h8220000;
      18216: inst = 32'h10408000;
      18217: inst = 32'hc4057d5;
      18218: inst = 32'h8220000;
      18219: inst = 32'h10408000;
      18220: inst = 32'hc4057d6;
      18221: inst = 32'h8220000;
      18222: inst = 32'h10408000;
      18223: inst = 32'hc4057d7;
      18224: inst = 32'h8220000;
      18225: inst = 32'h10408000;
      18226: inst = 32'hc4057d8;
      18227: inst = 32'h8220000;
      18228: inst = 32'h10408000;
      18229: inst = 32'hc4057d9;
      18230: inst = 32'h8220000;
      18231: inst = 32'h10408000;
      18232: inst = 32'hc4057da;
      18233: inst = 32'h8220000;
      18234: inst = 32'h10408000;
      18235: inst = 32'hc4057db;
      18236: inst = 32'h8220000;
      18237: inst = 32'h10408000;
      18238: inst = 32'hc4057dc;
      18239: inst = 32'h8220000;
      18240: inst = 32'h10408000;
      18241: inst = 32'hc4057dd;
      18242: inst = 32'h8220000;
      18243: inst = 32'h10408000;
      18244: inst = 32'hc4057de;
      18245: inst = 32'h8220000;
      18246: inst = 32'h10408000;
      18247: inst = 32'hc4057df;
      18248: inst = 32'h8220000;
      18249: inst = 32'hc207bd0;
      18250: inst = 32'h10408000;
      18251: inst = 32'hc40531b;
      18252: inst = 32'h8220000;
      18253: inst = 32'h10408000;
      18254: inst = 32'hc405344;
      18255: inst = 32'h8220000;
      18256: inst = 32'hc207bcf;
      18257: inst = 32'h10408000;
      18258: inst = 32'hc405321;
      18259: inst = 32'h8220000;
      18260: inst = 32'h10408000;
      18261: inst = 32'hc40533e;
      18262: inst = 32'h8220000;
      18263: inst = 32'h10408000;
      18264: inst = 32'hc405381;
      18265: inst = 32'h8220000;
      18266: inst = 32'h10408000;
      18267: inst = 32'hc40539e;
      18268: inst = 32'h8220000;
      18269: inst = 32'h10408000;
      18270: inst = 32'hc4053e1;
      18271: inst = 32'h8220000;
      18272: inst = 32'h10408000;
      18273: inst = 32'hc4053fe;
      18274: inst = 32'h8220000;
      18275: inst = 32'h10408000;
      18276: inst = 32'hc405441;
      18277: inst = 32'h8220000;
      18278: inst = 32'h10408000;
      18279: inst = 32'hc405448;
      18280: inst = 32'h8220000;
      18281: inst = 32'h10408000;
      18282: inst = 32'hc405457;
      18283: inst = 32'h8220000;
      18284: inst = 32'h10408000;
      18285: inst = 32'hc40545e;
      18286: inst = 32'h8220000;
      18287: inst = 32'h10408000;
      18288: inst = 32'hc405501;
      18289: inst = 32'h8220000;
      18290: inst = 32'h10408000;
      18291: inst = 32'hc40551e;
      18292: inst = 32'h8220000;
      18293: inst = 32'h10408000;
      18294: inst = 32'hc405561;
      18295: inst = 32'h8220000;
      18296: inst = 32'h10408000;
      18297: inst = 32'hc40557e;
      18298: inst = 32'h8220000;
      18299: inst = 32'h10408000;
      18300: inst = 32'hc4055b9;
      18301: inst = 32'h8220000;
      18302: inst = 32'h10408000;
      18303: inst = 32'hc4055c1;
      18304: inst = 32'h8220000;
      18305: inst = 32'h10408000;
      18306: inst = 32'hc4055de;
      18307: inst = 32'h8220000;
      18308: inst = 32'h10408000;
      18309: inst = 32'hc4055e6;
      18310: inst = 32'h8220000;
      18311: inst = 32'h10408000;
      18312: inst = 32'hc40561e;
      18313: inst = 32'h8220000;
      18314: inst = 32'h10408000;
      18315: inst = 32'hc405621;
      18316: inst = 32'h8220000;
      18317: inst = 32'h10408000;
      18318: inst = 32'hc40563e;
      18319: inst = 32'h8220000;
      18320: inst = 32'h10408000;
      18321: inst = 32'hc405641;
      18322: inst = 32'h8220000;
      18323: inst = 32'h10408000;
      18324: inst = 32'hc405681;
      18325: inst = 32'h8220000;
      18326: inst = 32'h10408000;
      18327: inst = 32'hc405698;
      18328: inst = 32'h8220000;
      18329: inst = 32'h10408000;
      18330: inst = 32'hc40569e;
      18331: inst = 32'h8220000;
      18332: inst = 32'h10408000;
      18333: inst = 32'hc4056e1;
      18334: inst = 32'h8220000;
      18335: inst = 32'h10408000;
      18336: inst = 32'hc4056fe;
      18337: inst = 32'h8220000;
      18338: inst = 32'hc207390;
      18339: inst = 32'h10408000;
      18340: inst = 32'hc40537a;
      18341: inst = 32'h8220000;
      18342: inst = 32'h10408000;
      18343: inst = 32'hc4053a5;
      18344: inst = 32'h8220000;
      18345: inst = 32'hc2052aa;
      18346: inst = 32'h10408000;
      18347: inst = 32'hc405389;
      18348: inst = 32'h8220000;
      18349: inst = 32'h10408000;
      18350: inst = 32'hc405396;
      18351: inst = 32'h8220000;
      18352: inst = 32'h10408000;
      18353: inst = 32'hc4054fb;
      18354: inst = 32'h8220000;
      18355: inst = 32'h10408000;
      18356: inst = 32'hc405503;
      18357: inst = 32'h8220000;
      18358: inst = 32'h10408000;
      18359: inst = 32'hc40551c;
      18360: inst = 32'h8220000;
      18361: inst = 32'h10408000;
      18362: inst = 32'hc405524;
      18363: inst = 32'h8220000;
      18364: inst = 32'h10408000;
      18365: inst = 32'hc4055c8;
      18366: inst = 32'h8220000;
      18367: inst = 32'h10408000;
      18368: inst = 32'hc4055d7;
      18369: inst = 32'h8220000;
      18370: inst = 32'h10408000;
      18371: inst = 32'hc405619;
      18372: inst = 32'h8220000;
      18373: inst = 32'h10408000;
      18374: inst = 32'hc405622;
      18375: inst = 32'h8220000;
      18376: inst = 32'h10408000;
      18377: inst = 32'hc40563d;
      18378: inst = 32'h8220000;
      18379: inst = 32'h10408000;
      18380: inst = 32'hc405646;
      18381: inst = 32'h8220000;
      18382: inst = 32'hc206b70;
      18383: inst = 32'h10408000;
      18384: inst = 32'hc4053d9;
      18385: inst = 32'h8220000;
      18386: inst = 32'h10408000;
      18387: inst = 32'hc405406;
      18388: inst = 32'h8220000;
      18389: inst = 32'h10408000;
      18390: inst = 32'hc405556;
      18391: inst = 32'h8220000;
      18392: inst = 32'h10408000;
      18393: inst = 32'hc405589;
      18394: inst = 32'h8220000;
      18395: inst = 32'h10408000;
      18396: inst = 32'hc4055b5;
      18397: inst = 32'h8220000;
      18398: inst = 32'h10408000;
      18399: inst = 32'hc4055ea;
      18400: inst = 32'h8220000;
      18401: inst = 32'h10408000;
      18402: inst = 32'hc405732;
      18403: inst = 32'h8220000;
      18404: inst = 32'h10408000;
      18405: inst = 32'hc40576d;
      18406: inst = 32'h8220000;
      18407: inst = 32'hc20736e;
      18408: inst = 32'h10408000;
      18409: inst = 32'hc4053e0;
      18410: inst = 32'h8220000;
      18411: inst = 32'h10408000;
      18412: inst = 32'hc4053ff;
      18413: inst = 32'h8220000;
      18414: inst = 32'hc205aaa;
      18415: inst = 32'h10408000;
      18416: inst = 32'hc4053e4;
      18417: inst = 32'h8220000;
      18418: inst = 32'h10408000;
      18419: inst = 32'hc4053fb;
      18420: inst = 32'h8220000;
      18421: inst = 32'hc208431;
      18422: inst = 32'h10408000;
      18423: inst = 32'hc4053e8;
      18424: inst = 32'h8220000;
      18425: inst = 32'h10408000;
      18426: inst = 32'hc4053f7;
      18427: inst = 32'h8220000;
      18428: inst = 32'h10408000;
      18429: inst = 32'hc405439;
      18430: inst = 32'h8220000;
      18431: inst = 32'h10408000;
      18432: inst = 32'hc405466;
      18433: inst = 32'h8220000;
      18434: inst = 32'h10408000;
      18435: inst = 32'hc4055b6;
      18436: inst = 32'h8220000;
      18437: inst = 32'h10408000;
      18438: inst = 32'hc4055e9;
      18439: inst = 32'h8220000;
      18440: inst = 32'h10408000;
      18441: inst = 32'hc405733;
      18442: inst = 32'h8220000;
      18443: inst = 32'h10408000;
      18444: inst = 32'hc40576c;
      18445: inst = 32'h8220000;
      18446: inst = 32'hc206b4d;
      18447: inst = 32'h10408000;
      18448: inst = 32'hc40543c;
      18449: inst = 32'h8220000;
      18450: inst = 32'h10408000;
      18451: inst = 32'hc405444;
      18452: inst = 32'h8220000;
      18453: inst = 32'h10408000;
      18454: inst = 32'hc40545b;
      18455: inst = 32'h8220000;
      18456: inst = 32'h10408000;
      18457: inst = 32'hc405463;
      18458: inst = 32'h8220000;
      18459: inst = 32'h10408000;
      18460: inst = 32'hc405563;
      18461: inst = 32'h8220000;
      18462: inst = 32'h10408000;
      18463: inst = 32'hc40557c;
      18464: inst = 32'h8220000;
      18465: inst = 32'h10408000;
      18466: inst = 32'hc405682;
      18467: inst = 32'h8220000;
      18468: inst = 32'h10408000;
      18469: inst = 32'hc40569d;
      18470: inst = 32'h8220000;
      18471: inst = 32'hc208430;
      18472: inst = 32'h10408000;
      18473: inst = 32'hc405440;
      18474: inst = 32'h8220000;
      18475: inst = 32'h10408000;
      18476: inst = 32'hc40545f;
      18477: inst = 32'h8220000;
      18478: inst = 32'hc207bf1;
      18479: inst = 32'h10408000;
      18480: inst = 32'hc405498;
      18481: inst = 32'h8220000;
      18482: inst = 32'h10408000;
      18483: inst = 32'hc4054c7;
      18484: inst = 32'h8220000;
      18485: inst = 32'h10408000;
      18486: inst = 32'hc405615;
      18487: inst = 32'h8220000;
      18488: inst = 32'h10408000;
      18489: inst = 32'hc40564a;
      18490: inst = 32'h8220000;
      18491: inst = 32'hc207bef;
      18492: inst = 32'h10408000;
      18493: inst = 32'hc40549b;
      18494: inst = 32'h8220000;
      18495: inst = 32'h10408000;
      18496: inst = 32'hc4054c4;
      18497: inst = 32'h8220000;
      18498: inst = 32'h10408000;
      18499: inst = 32'hc405687;
      18500: inst = 32'h8220000;
      18501: inst = 32'h10408000;
      18502: inst = 32'hc4056e2;
      18503: inst = 32'h8220000;
      18504: inst = 32'h10408000;
      18505: inst = 32'hc4056fd;
      18506: inst = 32'h8220000;
      18507: inst = 32'hc205aeb;
      18508: inst = 32'h10408000;
      18509: inst = 32'hc40549f;
      18510: inst = 32'h8220000;
      18511: inst = 32'h10408000;
      18512: inst = 32'hc4054c0;
      18513: inst = 32'h8220000;
      18514: inst = 32'hc206b6e;
      18515: inst = 32'h10408000;
      18516: inst = 32'hc4054a8;
      18517: inst = 32'h8220000;
      18518: inst = 32'h10408000;
      18519: inst = 32'hc4054b7;
      18520: inst = 32'h8220000;
      18521: inst = 32'h10408000;
      18522: inst = 32'hc4056e7;
      18523: inst = 32'h8220000;
      18524: inst = 32'h10408000;
      18525: inst = 32'hc4056f8;
      18526: inst = 32'h8220000;
      18527: inst = 32'hc2073b0;
      18528: inst = 32'h10408000;
      18529: inst = 32'hc4054f7;
      18530: inst = 32'h8220000;
      18531: inst = 32'h10408000;
      18532: inst = 32'hc405528;
      18533: inst = 32'h8220000;
      18534: inst = 32'h10408000;
      18535: inst = 32'hc405674;
      18536: inst = 32'h8220000;
      18537: inst = 32'h10408000;
      18538: inst = 32'hc4056ab;
      18539: inst = 32'h8220000;
      18540: inst = 32'hc2073ae;
      18541: inst = 32'h10408000;
      18542: inst = 32'hc4054ff;
      18543: inst = 32'h8220000;
      18544: inst = 32'h10408000;
      18545: inst = 32'hc405520;
      18546: inst = 32'h8220000;
      18547: inst = 32'hc20632d;
      18548: inst = 32'h10408000;
      18549: inst = 32'hc405508;
      18550: inst = 32'h8220000;
      18551: inst = 32'h10408000;
      18552: inst = 32'hc405517;
      18553: inst = 32'h8220000;
      18554: inst = 32'h10408000;
      18555: inst = 32'hc405747;
      18556: inst = 32'h8220000;
      18557: inst = 32'h10408000;
      18558: inst = 32'hc405758;
      18559: inst = 32'h8220000;
      18560: inst = 32'hc206b2d;
      18561: inst = 32'h10408000;
      18562: inst = 32'hc40555a;
      18563: inst = 32'h8220000;
      18564: inst = 32'h10408000;
      18565: inst = 32'hc405585;
      18566: inst = 32'h8220000;
      18567: inst = 32'hc20630c;
      18568: inst = 32'h10408000;
      18569: inst = 32'hc4055be;
      18570: inst = 32'h8220000;
      18571: inst = 32'h10408000;
      18572: inst = 32'hc4055e1;
      18573: inst = 32'h8220000;
      18574: inst = 32'h10408000;
      18575: inst = 32'hc405678;
      18576: inst = 32'h8220000;
      18577: inst = 32'hc20632c;
      18578: inst = 32'h10408000;
      18579: inst = 32'hc4056a7;
      18580: inst = 32'h8220000;
      18581: inst = 32'hc206b90;
      18582: inst = 32'h10408000;
      18583: inst = 32'hc4056d3;
      18584: inst = 32'h8220000;
      18585: inst = 32'h10408000;
      18586: inst = 32'hc40570c;
      18587: inst = 32'h8220000;
      18588: inst = 32'hc207c11;
      18589: inst = 32'h10408000;
      18590: inst = 32'hc405792;
      18591: inst = 32'h8220000;
      18592: inst = 32'h10408000;
      18593: inst = 32'hc4057cd;
      18594: inst = 32'h8220000;
      18595: inst = 32'h58000000;
      18596: inst = 32'hc20ea25;
      18597: inst = 32'h10408000;
      18598: inst = 32'hc40464d;
      18599: inst = 32'h8220000;
      18600: inst = 32'h10408000;
      18601: inst = 32'hc40464e;
      18602: inst = 32'h8220000;
      18603: inst = 32'h10408000;
      18604: inst = 32'hc40464f;
      18605: inst = 32'h8220000;
      18606: inst = 32'h10408000;
      18607: inst = 32'hc404650;
      18608: inst = 32'h8220000;
      18609: inst = 32'h10408000;
      18610: inst = 32'hc404651;
      18611: inst = 32'h8220000;
      18612: inst = 32'h10408000;
      18613: inst = 32'hc404652;
      18614: inst = 32'h8220000;
      18615: inst = 32'h10408000;
      18616: inst = 32'hc404653;
      18617: inst = 32'h8220000;
      18618: inst = 32'h10408000;
      18619: inst = 32'hc404654;
      18620: inst = 32'h8220000;
      18621: inst = 32'h10408000;
      18622: inst = 32'hc404655;
      18623: inst = 32'h8220000;
      18624: inst = 32'h10408000;
      18625: inst = 32'hc404659;
      18626: inst = 32'h8220000;
      18627: inst = 32'h10408000;
      18628: inst = 32'hc40465a;
      18629: inst = 32'h8220000;
      18630: inst = 32'h10408000;
      18631: inst = 32'hc40465b;
      18632: inst = 32'h8220000;
      18633: inst = 32'h10408000;
      18634: inst = 32'hc40465c;
      18635: inst = 32'h8220000;
      18636: inst = 32'h10408000;
      18637: inst = 32'hc40465d;
      18638: inst = 32'h8220000;
      18639: inst = 32'h10408000;
      18640: inst = 32'hc40465e;
      18641: inst = 32'h8220000;
      18642: inst = 32'h10408000;
      18643: inst = 32'hc40465f;
      18644: inst = 32'h8220000;
      18645: inst = 32'h10408000;
      18646: inst = 32'hc404660;
      18647: inst = 32'h8220000;
      18648: inst = 32'h10408000;
      18649: inst = 32'hc404661;
      18650: inst = 32'h8220000;
      18651: inst = 32'h10408000;
      18652: inst = 32'hc404663;
      18653: inst = 32'h8220000;
      18654: inst = 32'h10408000;
      18655: inst = 32'hc404664;
      18656: inst = 32'h8220000;
      18657: inst = 32'h10408000;
      18658: inst = 32'hc404665;
      18659: inst = 32'h8220000;
      18660: inst = 32'h10408000;
      18661: inst = 32'hc404666;
      18662: inst = 32'h8220000;
      18663: inst = 32'h10408000;
      18664: inst = 32'hc404667;
      18665: inst = 32'h8220000;
      18666: inst = 32'h10408000;
      18667: inst = 32'hc404668;
      18668: inst = 32'h8220000;
      18669: inst = 32'h10408000;
      18670: inst = 32'hc404669;
      18671: inst = 32'h8220000;
      18672: inst = 32'h10408000;
      18673: inst = 32'hc40466a;
      18674: inst = 32'h8220000;
      18675: inst = 32'h10408000;
      18676: inst = 32'hc40466b;
      18677: inst = 32'h8220000;
      18678: inst = 32'h10408000;
      18679: inst = 32'hc404671;
      18680: inst = 32'h8220000;
      18681: inst = 32'h10408000;
      18682: inst = 32'hc404672;
      18683: inst = 32'h8220000;
      18684: inst = 32'h10408000;
      18685: inst = 32'hc404673;
      18686: inst = 32'h8220000;
      18687: inst = 32'h10408000;
      18688: inst = 32'hc404674;
      18689: inst = 32'h8220000;
      18690: inst = 32'h10408000;
      18691: inst = 32'hc404675;
      18692: inst = 32'h8220000;
      18693: inst = 32'h10408000;
      18694: inst = 32'hc404676;
      18695: inst = 32'h8220000;
      18696: inst = 32'h10408000;
      18697: inst = 32'hc404677;
      18698: inst = 32'h8220000;
      18699: inst = 32'h10408000;
      18700: inst = 32'hc404678;
      18701: inst = 32'h8220000;
      18702: inst = 32'h10408000;
      18703: inst = 32'hc404679;
      18704: inst = 32'h8220000;
      18705: inst = 32'h10408000;
      18706: inst = 32'hc40467c;
      18707: inst = 32'h8220000;
      18708: inst = 32'h10408000;
      18709: inst = 32'hc40467d;
      18710: inst = 32'h8220000;
      18711: inst = 32'h10408000;
      18712: inst = 32'hc40467e;
      18713: inst = 32'h8220000;
      18714: inst = 32'h10408000;
      18715: inst = 32'hc40467f;
      18716: inst = 32'h8220000;
      18717: inst = 32'h10408000;
      18718: inst = 32'hc404680;
      18719: inst = 32'h8220000;
      18720: inst = 32'h10408000;
      18721: inst = 32'hc404681;
      18722: inst = 32'h8220000;
      18723: inst = 32'h10408000;
      18724: inst = 32'hc404682;
      18725: inst = 32'h8220000;
      18726: inst = 32'h10408000;
      18727: inst = 32'hc404683;
      18728: inst = 32'h8220000;
      18729: inst = 32'h10408000;
      18730: inst = 32'hc404684;
      18731: inst = 32'h8220000;
      18732: inst = 32'h10408000;
      18733: inst = 32'hc404685;
      18734: inst = 32'h8220000;
      18735: inst = 32'h10408000;
      18736: inst = 32'hc40468b;
      18737: inst = 32'h8220000;
      18738: inst = 32'h10408000;
      18739: inst = 32'hc40468c;
      18740: inst = 32'h8220000;
      18741: inst = 32'h10408000;
      18742: inst = 32'hc40468d;
      18743: inst = 32'h8220000;
      18744: inst = 32'h10408000;
      18745: inst = 32'hc40468e;
      18746: inst = 32'h8220000;
      18747: inst = 32'h10408000;
      18748: inst = 32'hc40468f;
      18749: inst = 32'h8220000;
      18750: inst = 32'h10408000;
      18751: inst = 32'hc404690;
      18752: inst = 32'h8220000;
      18753: inst = 32'h10408000;
      18754: inst = 32'hc404691;
      18755: inst = 32'h8220000;
      18756: inst = 32'h10408000;
      18757: inst = 32'hc404692;
      18758: inst = 32'h8220000;
      18759: inst = 32'h10408000;
      18760: inst = 32'hc404693;
      18761: inst = 32'h8220000;
      18762: inst = 32'h10408000;
      18763: inst = 32'hc4046ac;
      18764: inst = 32'h8220000;
      18765: inst = 32'h10408000;
      18766: inst = 32'hc4046ad;
      18767: inst = 32'h8220000;
      18768: inst = 32'h10408000;
      18769: inst = 32'hc4046ae;
      18770: inst = 32'h8220000;
      18771: inst = 32'h10408000;
      18772: inst = 32'hc4046af;
      18773: inst = 32'h8220000;
      18774: inst = 32'h10408000;
      18775: inst = 32'hc4046b0;
      18776: inst = 32'h8220000;
      18777: inst = 32'h10408000;
      18778: inst = 32'hc4046b1;
      18779: inst = 32'h8220000;
      18780: inst = 32'h10408000;
      18781: inst = 32'hc4046b2;
      18782: inst = 32'h8220000;
      18783: inst = 32'h10408000;
      18784: inst = 32'hc4046b3;
      18785: inst = 32'h8220000;
      18786: inst = 32'h10408000;
      18787: inst = 32'hc4046b4;
      18788: inst = 32'h8220000;
      18789: inst = 32'h10408000;
      18790: inst = 32'hc4046b5;
      18791: inst = 32'h8220000;
      18792: inst = 32'h10408000;
      18793: inst = 32'hc4046b8;
      18794: inst = 32'h8220000;
      18795: inst = 32'h10408000;
      18796: inst = 32'hc4046b9;
      18797: inst = 32'h8220000;
      18798: inst = 32'h10408000;
      18799: inst = 32'hc4046ba;
      18800: inst = 32'h8220000;
      18801: inst = 32'h10408000;
      18802: inst = 32'hc4046bb;
      18803: inst = 32'h8220000;
      18804: inst = 32'h10408000;
      18805: inst = 32'hc4046bc;
      18806: inst = 32'h8220000;
      18807: inst = 32'h10408000;
      18808: inst = 32'hc4046bd;
      18809: inst = 32'h8220000;
      18810: inst = 32'h10408000;
      18811: inst = 32'hc4046be;
      18812: inst = 32'h8220000;
      18813: inst = 32'h10408000;
      18814: inst = 32'hc4046bf;
      18815: inst = 32'h8220000;
      18816: inst = 32'h10408000;
      18817: inst = 32'hc4046c0;
      18818: inst = 32'h8220000;
      18819: inst = 32'h10408000;
      18820: inst = 32'hc4046c1;
      18821: inst = 32'h8220000;
      18822: inst = 32'h10408000;
      18823: inst = 32'hc4046c3;
      18824: inst = 32'h8220000;
      18825: inst = 32'h10408000;
      18826: inst = 32'hc4046c4;
      18827: inst = 32'h8220000;
      18828: inst = 32'h10408000;
      18829: inst = 32'hc4046c5;
      18830: inst = 32'h8220000;
      18831: inst = 32'h10408000;
      18832: inst = 32'hc4046c6;
      18833: inst = 32'h8220000;
      18834: inst = 32'h10408000;
      18835: inst = 32'hc4046c7;
      18836: inst = 32'h8220000;
      18837: inst = 32'h10408000;
      18838: inst = 32'hc4046c8;
      18839: inst = 32'h8220000;
      18840: inst = 32'h10408000;
      18841: inst = 32'hc4046c9;
      18842: inst = 32'h8220000;
      18843: inst = 32'h10408000;
      18844: inst = 32'hc4046ca;
      18845: inst = 32'h8220000;
      18846: inst = 32'h10408000;
      18847: inst = 32'hc4046cb;
      18848: inst = 32'h8220000;
      18849: inst = 32'h10408000;
      18850: inst = 32'hc4046d0;
      18851: inst = 32'h8220000;
      18852: inst = 32'h10408000;
      18853: inst = 32'hc4046d1;
      18854: inst = 32'h8220000;
      18855: inst = 32'h10408000;
      18856: inst = 32'hc4046d2;
      18857: inst = 32'h8220000;
      18858: inst = 32'h10408000;
      18859: inst = 32'hc4046d3;
      18860: inst = 32'h8220000;
      18861: inst = 32'h10408000;
      18862: inst = 32'hc4046d4;
      18863: inst = 32'h8220000;
      18864: inst = 32'h10408000;
      18865: inst = 32'hc4046d5;
      18866: inst = 32'h8220000;
      18867: inst = 32'h10408000;
      18868: inst = 32'hc4046d6;
      18869: inst = 32'h8220000;
      18870: inst = 32'h10408000;
      18871: inst = 32'hc4046d7;
      18872: inst = 32'h8220000;
      18873: inst = 32'h10408000;
      18874: inst = 32'hc4046d8;
      18875: inst = 32'h8220000;
      18876: inst = 32'h10408000;
      18877: inst = 32'hc4046da;
      18878: inst = 32'h8220000;
      18879: inst = 32'h10408000;
      18880: inst = 32'hc4046dc;
      18881: inst = 32'h8220000;
      18882: inst = 32'h10408000;
      18883: inst = 32'hc4046dd;
      18884: inst = 32'h8220000;
      18885: inst = 32'h10408000;
      18886: inst = 32'hc4046de;
      18887: inst = 32'h8220000;
      18888: inst = 32'h10408000;
      18889: inst = 32'hc4046df;
      18890: inst = 32'h8220000;
      18891: inst = 32'h10408000;
      18892: inst = 32'hc4046e0;
      18893: inst = 32'h8220000;
      18894: inst = 32'h10408000;
      18895: inst = 32'hc4046e1;
      18896: inst = 32'h8220000;
      18897: inst = 32'h10408000;
      18898: inst = 32'hc4046e2;
      18899: inst = 32'h8220000;
      18900: inst = 32'h10408000;
      18901: inst = 32'hc4046e3;
      18902: inst = 32'h8220000;
      18903: inst = 32'h10408000;
      18904: inst = 32'hc4046e4;
      18905: inst = 32'h8220000;
      18906: inst = 32'h10408000;
      18907: inst = 32'hc4046e5;
      18908: inst = 32'h8220000;
      18909: inst = 32'h10408000;
      18910: inst = 32'hc4046ea;
      18911: inst = 32'h8220000;
      18912: inst = 32'h10408000;
      18913: inst = 32'hc4046eb;
      18914: inst = 32'h8220000;
      18915: inst = 32'h10408000;
      18916: inst = 32'hc4046ec;
      18917: inst = 32'h8220000;
      18918: inst = 32'h10408000;
      18919: inst = 32'hc4046ed;
      18920: inst = 32'h8220000;
      18921: inst = 32'h10408000;
      18922: inst = 32'hc4046ee;
      18923: inst = 32'h8220000;
      18924: inst = 32'h10408000;
      18925: inst = 32'hc4046ef;
      18926: inst = 32'h8220000;
      18927: inst = 32'h10408000;
      18928: inst = 32'hc4046f0;
      18929: inst = 32'h8220000;
      18930: inst = 32'h10408000;
      18931: inst = 32'hc4046f1;
      18932: inst = 32'h8220000;
      18933: inst = 32'h10408000;
      18934: inst = 32'hc4046f2;
      18935: inst = 32'h8220000;
      18936: inst = 32'h10408000;
      18937: inst = 32'hc4046f3;
      18938: inst = 32'h8220000;
      18939: inst = 32'h10408000;
      18940: inst = 32'hc40470b;
      18941: inst = 32'h8220000;
      18942: inst = 32'h10408000;
      18943: inst = 32'hc40470c;
      18944: inst = 32'h8220000;
      18945: inst = 32'h10408000;
      18946: inst = 32'hc40470d;
      18947: inst = 32'h8220000;
      18948: inst = 32'h10408000;
      18949: inst = 32'hc404717;
      18950: inst = 32'h8220000;
      18951: inst = 32'h10408000;
      18952: inst = 32'hc404718;
      18953: inst = 32'h8220000;
      18954: inst = 32'h10408000;
      18955: inst = 32'hc404719;
      18956: inst = 32'h8220000;
      18957: inst = 32'h10408000;
      18958: inst = 32'hc404728;
      18959: inst = 32'h8220000;
      18960: inst = 32'h10408000;
      18961: inst = 32'hc404729;
      18962: inst = 32'h8220000;
      18963: inst = 32'h10408000;
      18964: inst = 32'hc40472a;
      18965: inst = 32'h8220000;
      18966: inst = 32'h10408000;
      18967: inst = 32'hc40472b;
      18968: inst = 32'h8220000;
      18969: inst = 32'h10408000;
      18970: inst = 32'hc404730;
      18971: inst = 32'h8220000;
      18972: inst = 32'h10408000;
      18973: inst = 32'hc404731;
      18974: inst = 32'h8220000;
      18975: inst = 32'h10408000;
      18976: inst = 32'hc404735;
      18977: inst = 32'h8220000;
      18978: inst = 32'h10408000;
      18979: inst = 32'hc404736;
      18980: inst = 32'h8220000;
      18981: inst = 32'h10408000;
      18982: inst = 32'hc404737;
      18983: inst = 32'h8220000;
      18984: inst = 32'h10408000;
      18985: inst = 32'hc404739;
      18986: inst = 32'h8220000;
      18987: inst = 32'h10408000;
      18988: inst = 32'hc40473a;
      18989: inst = 32'h8220000;
      18990: inst = 32'h10408000;
      18991: inst = 32'hc404742;
      18992: inst = 32'h8220000;
      18993: inst = 32'h10408000;
      18994: inst = 32'hc404743;
      18995: inst = 32'h8220000;
      18996: inst = 32'h10408000;
      18997: inst = 32'hc404744;
      18998: inst = 32'h8220000;
      18999: inst = 32'h10408000;
      19000: inst = 32'hc404745;
      19001: inst = 32'h8220000;
      19002: inst = 32'h10408000;
      19003: inst = 32'hc404749;
      19004: inst = 32'h8220000;
      19005: inst = 32'h10408000;
      19006: inst = 32'hc40474a;
      19007: inst = 32'h8220000;
      19008: inst = 32'h10408000;
      19009: inst = 32'hc40474b;
      19010: inst = 32'h8220000;
      19011: inst = 32'h10408000;
      19012: inst = 32'hc40476b;
      19013: inst = 32'h8220000;
      19014: inst = 32'h10408000;
      19015: inst = 32'hc40476c;
      19016: inst = 32'h8220000;
      19017: inst = 32'h10408000;
      19018: inst = 32'hc404777;
      19019: inst = 32'h8220000;
      19020: inst = 32'h10408000;
      19021: inst = 32'hc404778;
      19022: inst = 32'h8220000;
      19023: inst = 32'h10408000;
      19024: inst = 32'hc404788;
      19025: inst = 32'h8220000;
      19026: inst = 32'h10408000;
      19027: inst = 32'hc404789;
      19028: inst = 32'h8220000;
      19029: inst = 32'h10408000;
      19030: inst = 32'hc40478a;
      19031: inst = 32'h8220000;
      19032: inst = 32'h10408000;
      19033: inst = 32'hc404790;
      19034: inst = 32'h8220000;
      19035: inst = 32'h10408000;
      19036: inst = 32'hc404791;
      19037: inst = 32'h8220000;
      19038: inst = 32'h10408000;
      19039: inst = 32'hc404795;
      19040: inst = 32'h8220000;
      19041: inst = 32'h10408000;
      19042: inst = 32'hc404799;
      19043: inst = 32'h8220000;
      19044: inst = 32'h10408000;
      19045: inst = 32'hc40479a;
      19046: inst = 32'h8220000;
      19047: inst = 32'h10408000;
      19048: inst = 32'hc4047a2;
      19049: inst = 32'h8220000;
      19050: inst = 32'h10408000;
      19051: inst = 32'hc4047a3;
      19052: inst = 32'h8220000;
      19053: inst = 32'h10408000;
      19054: inst = 32'hc4047a4;
      19055: inst = 32'h8220000;
      19056: inst = 32'h10408000;
      19057: inst = 32'hc4047a9;
      19058: inst = 32'h8220000;
      19059: inst = 32'h10408000;
      19060: inst = 32'hc4047aa;
      19061: inst = 32'h8220000;
      19062: inst = 32'h10408000;
      19063: inst = 32'hc4047cb;
      19064: inst = 32'h8220000;
      19065: inst = 32'h10408000;
      19066: inst = 32'hc4047cc;
      19067: inst = 32'h8220000;
      19068: inst = 32'h10408000;
      19069: inst = 32'hc4047ce;
      19070: inst = 32'h8220000;
      19071: inst = 32'h10408000;
      19072: inst = 32'hc4047cf;
      19073: inst = 32'h8220000;
      19074: inst = 32'h10408000;
      19075: inst = 32'hc4047d0;
      19076: inst = 32'h8220000;
      19077: inst = 32'h10408000;
      19078: inst = 32'hc4047d1;
      19079: inst = 32'h8220000;
      19080: inst = 32'h10408000;
      19081: inst = 32'hc4047d2;
      19082: inst = 32'h8220000;
      19083: inst = 32'h10408000;
      19084: inst = 32'hc4047d7;
      19085: inst = 32'h8220000;
      19086: inst = 32'h10408000;
      19087: inst = 32'hc4047d8;
      19088: inst = 32'h8220000;
      19089: inst = 32'h10408000;
      19090: inst = 32'hc4047da;
      19091: inst = 32'h8220000;
      19092: inst = 32'h10408000;
      19093: inst = 32'hc4047db;
      19094: inst = 32'h8220000;
      19095: inst = 32'h10408000;
      19096: inst = 32'hc4047dc;
      19097: inst = 32'h8220000;
      19098: inst = 32'h10408000;
      19099: inst = 32'hc4047dd;
      19100: inst = 32'h8220000;
      19101: inst = 32'h10408000;
      19102: inst = 32'hc4047de;
      19103: inst = 32'h8220000;
      19104: inst = 32'h10408000;
      19105: inst = 32'hc4047e7;
      19106: inst = 32'h8220000;
      19107: inst = 32'h10408000;
      19108: inst = 32'hc4047e8;
      19109: inst = 32'h8220000;
      19110: inst = 32'h10408000;
      19111: inst = 32'hc4047e9;
      19112: inst = 32'h8220000;
      19113: inst = 32'h10408000;
      19114: inst = 32'hc4047f0;
      19115: inst = 32'h8220000;
      19116: inst = 32'h10408000;
      19117: inst = 32'hc4047f1;
      19118: inst = 32'h8220000;
      19119: inst = 32'h10408000;
      19120: inst = 32'hc4047f9;
      19121: inst = 32'h8220000;
      19122: inst = 32'h10408000;
      19123: inst = 32'hc4047fa;
      19124: inst = 32'h8220000;
      19125: inst = 32'h10408000;
      19126: inst = 32'hc404800;
      19127: inst = 32'h8220000;
      19128: inst = 32'h10408000;
      19129: inst = 32'hc404801;
      19130: inst = 32'h8220000;
      19131: inst = 32'h10408000;
      19132: inst = 32'hc404802;
      19133: inst = 32'h8220000;
      19134: inst = 32'h10408000;
      19135: inst = 32'hc404803;
      19136: inst = 32'h8220000;
      19137: inst = 32'h10408000;
      19138: inst = 32'hc404809;
      19139: inst = 32'h8220000;
      19140: inst = 32'h10408000;
      19141: inst = 32'hc40480a;
      19142: inst = 32'h8220000;
      19143: inst = 32'h10408000;
      19144: inst = 32'hc40480c;
      19145: inst = 32'h8220000;
      19146: inst = 32'h10408000;
      19147: inst = 32'hc40480d;
      19148: inst = 32'h8220000;
      19149: inst = 32'h10408000;
      19150: inst = 32'hc40480e;
      19151: inst = 32'h8220000;
      19152: inst = 32'h10408000;
      19153: inst = 32'hc40480f;
      19154: inst = 32'h8220000;
      19155: inst = 32'h10408000;
      19156: inst = 32'hc404810;
      19157: inst = 32'h8220000;
      19158: inst = 32'h10408000;
      19159: inst = 32'hc404811;
      19160: inst = 32'h8220000;
      19161: inst = 32'h10408000;
      19162: inst = 32'hc40482b;
      19163: inst = 32'h8220000;
      19164: inst = 32'h10408000;
      19165: inst = 32'hc40482c;
      19166: inst = 32'h8220000;
      19167: inst = 32'h10408000;
      19168: inst = 32'hc40482e;
      19169: inst = 32'h8220000;
      19170: inst = 32'h10408000;
      19171: inst = 32'hc40482f;
      19172: inst = 32'h8220000;
      19173: inst = 32'h10408000;
      19174: inst = 32'hc404830;
      19175: inst = 32'h8220000;
      19176: inst = 32'h10408000;
      19177: inst = 32'hc404831;
      19178: inst = 32'h8220000;
      19179: inst = 32'h10408000;
      19180: inst = 32'hc404832;
      19181: inst = 32'h8220000;
      19182: inst = 32'h10408000;
      19183: inst = 32'hc404837;
      19184: inst = 32'h8220000;
      19185: inst = 32'h10408000;
      19186: inst = 32'hc404838;
      19187: inst = 32'h8220000;
      19188: inst = 32'h10408000;
      19189: inst = 32'hc40483a;
      19190: inst = 32'h8220000;
      19191: inst = 32'h10408000;
      19192: inst = 32'hc40483b;
      19193: inst = 32'h8220000;
      19194: inst = 32'h10408000;
      19195: inst = 32'hc40483c;
      19196: inst = 32'h8220000;
      19197: inst = 32'h10408000;
      19198: inst = 32'hc40483d;
      19199: inst = 32'h8220000;
      19200: inst = 32'h10408000;
      19201: inst = 32'hc40483e;
      19202: inst = 32'h8220000;
      19203: inst = 32'h10408000;
      19204: inst = 32'hc404846;
      19205: inst = 32'h8220000;
      19206: inst = 32'h10408000;
      19207: inst = 32'hc404847;
      19208: inst = 32'h8220000;
      19209: inst = 32'h10408000;
      19210: inst = 32'hc404848;
      19211: inst = 32'h8220000;
      19212: inst = 32'h10408000;
      19213: inst = 32'hc404850;
      19214: inst = 32'h8220000;
      19215: inst = 32'h10408000;
      19216: inst = 32'hc404851;
      19217: inst = 32'h8220000;
      19218: inst = 32'h10408000;
      19219: inst = 32'hc404859;
      19220: inst = 32'h8220000;
      19221: inst = 32'h10408000;
      19222: inst = 32'hc40485a;
      19223: inst = 32'h8220000;
      19224: inst = 32'h10408000;
      19225: inst = 32'hc40485f;
      19226: inst = 32'h8220000;
      19227: inst = 32'h10408000;
      19228: inst = 32'hc404860;
      19229: inst = 32'h8220000;
      19230: inst = 32'h10408000;
      19231: inst = 32'hc404861;
      19232: inst = 32'h8220000;
      19233: inst = 32'h10408000;
      19234: inst = 32'hc404862;
      19235: inst = 32'h8220000;
      19236: inst = 32'h10408000;
      19237: inst = 32'hc404869;
      19238: inst = 32'h8220000;
      19239: inst = 32'h10408000;
      19240: inst = 32'hc40486a;
      19241: inst = 32'h8220000;
      19242: inst = 32'h10408000;
      19243: inst = 32'hc40486c;
      19244: inst = 32'h8220000;
      19245: inst = 32'h10408000;
      19246: inst = 32'hc40486d;
      19247: inst = 32'h8220000;
      19248: inst = 32'h10408000;
      19249: inst = 32'hc40486e;
      19250: inst = 32'h8220000;
      19251: inst = 32'h10408000;
      19252: inst = 32'hc40486f;
      19253: inst = 32'h8220000;
      19254: inst = 32'h10408000;
      19255: inst = 32'hc404870;
      19256: inst = 32'h8220000;
      19257: inst = 32'h10408000;
      19258: inst = 32'hc404871;
      19259: inst = 32'h8220000;
      19260: inst = 32'h10408000;
      19261: inst = 32'hc404872;
      19262: inst = 32'h8220000;
      19263: inst = 32'h10408000;
      19264: inst = 32'hc40488b;
      19265: inst = 32'h8220000;
      19266: inst = 32'h10408000;
      19267: inst = 32'hc40488c;
      19268: inst = 32'h8220000;
      19269: inst = 32'h10408000;
      19270: inst = 32'hc404897;
      19271: inst = 32'h8220000;
      19272: inst = 32'h10408000;
      19273: inst = 32'hc404898;
      19274: inst = 32'h8220000;
      19275: inst = 32'h10408000;
      19276: inst = 32'hc4048a6;
      19277: inst = 32'h8220000;
      19278: inst = 32'h10408000;
      19279: inst = 32'hc4048b0;
      19280: inst = 32'h8220000;
      19281: inst = 32'h10408000;
      19282: inst = 32'hc4048b1;
      19283: inst = 32'h8220000;
      19284: inst = 32'h10408000;
      19285: inst = 32'hc4048b4;
      19286: inst = 32'h8220000;
      19287: inst = 32'h10408000;
      19288: inst = 32'hc4048b5;
      19289: inst = 32'h8220000;
      19290: inst = 32'h10408000;
      19291: inst = 32'hc4048b9;
      19292: inst = 32'h8220000;
      19293: inst = 32'h10408000;
      19294: inst = 32'hc4048ba;
      19295: inst = 32'h8220000;
      19296: inst = 32'h10408000;
      19297: inst = 32'hc4048bf;
      19298: inst = 32'h8220000;
      19299: inst = 32'h10408000;
      19300: inst = 32'hc4048c9;
      19301: inst = 32'h8220000;
      19302: inst = 32'h10408000;
      19303: inst = 32'hc4048ca;
      19304: inst = 32'h8220000;
      19305: inst = 32'h10408000;
      19306: inst = 32'hc4048d1;
      19307: inst = 32'h8220000;
      19308: inst = 32'h10408000;
      19309: inst = 32'hc4048d2;
      19310: inst = 32'h8220000;
      19311: inst = 32'h10408000;
      19312: inst = 32'hc4048d3;
      19313: inst = 32'h8220000;
      19314: inst = 32'h10408000;
      19315: inst = 32'hc4048eb;
      19316: inst = 32'h8220000;
      19317: inst = 32'h10408000;
      19318: inst = 32'hc4048ec;
      19319: inst = 32'h8220000;
      19320: inst = 32'h10408000;
      19321: inst = 32'hc4048ed;
      19322: inst = 32'h8220000;
      19323: inst = 32'h10408000;
      19324: inst = 32'hc4048ee;
      19325: inst = 32'h8220000;
      19326: inst = 32'h10408000;
      19327: inst = 32'hc4048ef;
      19328: inst = 32'h8220000;
      19329: inst = 32'h10408000;
      19330: inst = 32'hc4048f0;
      19331: inst = 32'h8220000;
      19332: inst = 32'h10408000;
      19333: inst = 32'hc4048f1;
      19334: inst = 32'h8220000;
      19335: inst = 32'h10408000;
      19336: inst = 32'hc4048f2;
      19337: inst = 32'h8220000;
      19338: inst = 32'h10408000;
      19339: inst = 32'hc4048f3;
      19340: inst = 32'h8220000;
      19341: inst = 32'h10408000;
      19342: inst = 32'hc4048f4;
      19343: inst = 32'h8220000;
      19344: inst = 32'h10408000;
      19345: inst = 32'hc4048f5;
      19346: inst = 32'h8220000;
      19347: inst = 32'h10408000;
      19348: inst = 32'hc4048f7;
      19349: inst = 32'h8220000;
      19350: inst = 32'h10408000;
      19351: inst = 32'hc4048f8;
      19352: inst = 32'h8220000;
      19353: inst = 32'h10408000;
      19354: inst = 32'hc4048f9;
      19355: inst = 32'h8220000;
      19356: inst = 32'h10408000;
      19357: inst = 32'hc4048fa;
      19358: inst = 32'h8220000;
      19359: inst = 32'h10408000;
      19360: inst = 32'hc4048fb;
      19361: inst = 32'h8220000;
      19362: inst = 32'h10408000;
      19363: inst = 32'hc4048fc;
      19364: inst = 32'h8220000;
      19365: inst = 32'h10408000;
      19366: inst = 32'hc4048fd;
      19367: inst = 32'h8220000;
      19368: inst = 32'h10408000;
      19369: inst = 32'hc4048fe;
      19370: inst = 32'h8220000;
      19371: inst = 32'h10408000;
      19372: inst = 32'hc4048ff;
      19373: inst = 32'h8220000;
      19374: inst = 32'h10408000;
      19375: inst = 32'hc404900;
      19376: inst = 32'h8220000;
      19377: inst = 32'h10408000;
      19378: inst = 32'hc404901;
      19379: inst = 32'h8220000;
      19380: inst = 32'h10408000;
      19381: inst = 32'hc404904;
      19382: inst = 32'h8220000;
      19383: inst = 32'h10408000;
      19384: inst = 32'hc404905;
      19385: inst = 32'h8220000;
      19386: inst = 32'h10408000;
      19387: inst = 32'hc404906;
      19388: inst = 32'h8220000;
      19389: inst = 32'h10408000;
      19390: inst = 32'hc404907;
      19391: inst = 32'h8220000;
      19392: inst = 32'h10408000;
      19393: inst = 32'hc404908;
      19394: inst = 32'h8220000;
      19395: inst = 32'h10408000;
      19396: inst = 32'hc404909;
      19397: inst = 32'h8220000;
      19398: inst = 32'h10408000;
      19399: inst = 32'hc40490a;
      19400: inst = 32'h8220000;
      19401: inst = 32'h10408000;
      19402: inst = 32'hc40490b;
      19403: inst = 32'h8220000;
      19404: inst = 32'h10408000;
      19405: inst = 32'hc40490c;
      19406: inst = 32'h8220000;
      19407: inst = 32'h10408000;
      19408: inst = 32'hc40490d;
      19409: inst = 32'h8220000;
      19410: inst = 32'h10408000;
      19411: inst = 32'hc404910;
      19412: inst = 32'h8220000;
      19413: inst = 32'h10408000;
      19414: inst = 32'hc404911;
      19415: inst = 32'h8220000;
      19416: inst = 32'h10408000;
      19417: inst = 32'hc404912;
      19418: inst = 32'h8220000;
      19419: inst = 32'h10408000;
      19420: inst = 32'hc404913;
      19421: inst = 32'h8220000;
      19422: inst = 32'h10408000;
      19423: inst = 32'hc404914;
      19424: inst = 32'h8220000;
      19425: inst = 32'h10408000;
      19426: inst = 32'hc404915;
      19427: inst = 32'h8220000;
      19428: inst = 32'h10408000;
      19429: inst = 32'hc404916;
      19430: inst = 32'h8220000;
      19431: inst = 32'h10408000;
      19432: inst = 32'hc404917;
      19433: inst = 32'h8220000;
      19434: inst = 32'h10408000;
      19435: inst = 32'hc404918;
      19436: inst = 32'h8220000;
      19437: inst = 32'h10408000;
      19438: inst = 32'hc404919;
      19439: inst = 32'h8220000;
      19440: inst = 32'h10408000;
      19441: inst = 32'hc40491a;
      19442: inst = 32'h8220000;
      19443: inst = 32'h10408000;
      19444: inst = 32'hc40491e;
      19445: inst = 32'h8220000;
      19446: inst = 32'h10408000;
      19447: inst = 32'hc40491f;
      19448: inst = 32'h8220000;
      19449: inst = 32'h10408000;
      19450: inst = 32'hc404920;
      19451: inst = 32'h8220000;
      19452: inst = 32'h10408000;
      19453: inst = 32'hc404921;
      19454: inst = 32'h8220000;
      19455: inst = 32'h10408000;
      19456: inst = 32'hc404922;
      19457: inst = 32'h8220000;
      19458: inst = 32'h10408000;
      19459: inst = 32'hc404923;
      19460: inst = 32'h8220000;
      19461: inst = 32'h10408000;
      19462: inst = 32'hc404924;
      19463: inst = 32'h8220000;
      19464: inst = 32'h10408000;
      19465: inst = 32'hc404925;
      19466: inst = 32'h8220000;
      19467: inst = 32'h10408000;
      19468: inst = 32'hc404926;
      19469: inst = 32'h8220000;
      19470: inst = 32'h10408000;
      19471: inst = 32'hc404927;
      19472: inst = 32'h8220000;
      19473: inst = 32'h10408000;
      19474: inst = 32'hc404929;
      19475: inst = 32'h8220000;
      19476: inst = 32'h10408000;
      19477: inst = 32'hc40492a;
      19478: inst = 32'h8220000;
      19479: inst = 32'h10408000;
      19480: inst = 32'hc40492b;
      19481: inst = 32'h8220000;
      19482: inst = 32'h10408000;
      19483: inst = 32'hc40492c;
      19484: inst = 32'h8220000;
      19485: inst = 32'h10408000;
      19486: inst = 32'hc40492d;
      19487: inst = 32'h8220000;
      19488: inst = 32'h10408000;
      19489: inst = 32'hc40492e;
      19490: inst = 32'h8220000;
      19491: inst = 32'h10408000;
      19492: inst = 32'hc40492f;
      19493: inst = 32'h8220000;
      19494: inst = 32'h10408000;
      19495: inst = 32'hc404930;
      19496: inst = 32'h8220000;
      19497: inst = 32'h10408000;
      19498: inst = 32'hc404931;
      19499: inst = 32'h8220000;
      19500: inst = 32'h10408000;
      19501: inst = 32'hc404932;
      19502: inst = 32'h8220000;
      19503: inst = 32'h10408000;
      19504: inst = 32'hc404933;
      19505: inst = 32'h8220000;
      19506: inst = 32'h10408000;
      19507: inst = 32'hc40494b;
      19508: inst = 32'h8220000;
      19509: inst = 32'h10408000;
      19510: inst = 32'hc40494c;
      19511: inst = 32'h8220000;
      19512: inst = 32'h10408000;
      19513: inst = 32'hc40494d;
      19514: inst = 32'h8220000;
      19515: inst = 32'h10408000;
      19516: inst = 32'hc40494e;
      19517: inst = 32'h8220000;
      19518: inst = 32'h10408000;
      19519: inst = 32'hc40494f;
      19520: inst = 32'h8220000;
      19521: inst = 32'h10408000;
      19522: inst = 32'hc404950;
      19523: inst = 32'h8220000;
      19524: inst = 32'h10408000;
      19525: inst = 32'hc404951;
      19526: inst = 32'h8220000;
      19527: inst = 32'h10408000;
      19528: inst = 32'hc404952;
      19529: inst = 32'h8220000;
      19530: inst = 32'h10408000;
      19531: inst = 32'hc404953;
      19532: inst = 32'h8220000;
      19533: inst = 32'h10408000;
      19534: inst = 32'hc404954;
      19535: inst = 32'h8220000;
      19536: inst = 32'h10408000;
      19537: inst = 32'hc404957;
      19538: inst = 32'h8220000;
      19539: inst = 32'h10408000;
      19540: inst = 32'hc404958;
      19541: inst = 32'h8220000;
      19542: inst = 32'h10408000;
      19543: inst = 32'hc404959;
      19544: inst = 32'h8220000;
      19545: inst = 32'h10408000;
      19546: inst = 32'hc40495a;
      19547: inst = 32'h8220000;
      19548: inst = 32'h10408000;
      19549: inst = 32'hc40495b;
      19550: inst = 32'h8220000;
      19551: inst = 32'h10408000;
      19552: inst = 32'hc40495c;
      19553: inst = 32'h8220000;
      19554: inst = 32'h10408000;
      19555: inst = 32'hc40495d;
      19556: inst = 32'h8220000;
      19557: inst = 32'h10408000;
      19558: inst = 32'hc40495e;
      19559: inst = 32'h8220000;
      19560: inst = 32'h10408000;
      19561: inst = 32'hc40495f;
      19562: inst = 32'h8220000;
      19563: inst = 32'h10408000;
      19564: inst = 32'hc404960;
      19565: inst = 32'h8220000;
      19566: inst = 32'h10408000;
      19567: inst = 32'hc404961;
      19568: inst = 32'h8220000;
      19569: inst = 32'h10408000;
      19570: inst = 32'hc404963;
      19571: inst = 32'h8220000;
      19572: inst = 32'h10408000;
      19573: inst = 32'hc404964;
      19574: inst = 32'h8220000;
      19575: inst = 32'h10408000;
      19576: inst = 32'hc404965;
      19577: inst = 32'h8220000;
      19578: inst = 32'h10408000;
      19579: inst = 32'hc404966;
      19580: inst = 32'h8220000;
      19581: inst = 32'h10408000;
      19582: inst = 32'hc404967;
      19583: inst = 32'h8220000;
      19584: inst = 32'h10408000;
      19585: inst = 32'hc404968;
      19586: inst = 32'h8220000;
      19587: inst = 32'h10408000;
      19588: inst = 32'hc404969;
      19589: inst = 32'h8220000;
      19590: inst = 32'h10408000;
      19591: inst = 32'hc40496a;
      19592: inst = 32'h8220000;
      19593: inst = 32'h10408000;
      19594: inst = 32'hc40496b;
      19595: inst = 32'h8220000;
      19596: inst = 32'h10408000;
      19597: inst = 32'hc40496c;
      19598: inst = 32'h8220000;
      19599: inst = 32'h10408000;
      19600: inst = 32'hc40496d;
      19601: inst = 32'h8220000;
      19602: inst = 32'h10408000;
      19603: inst = 32'hc404970;
      19604: inst = 32'h8220000;
      19605: inst = 32'h10408000;
      19606: inst = 32'hc404971;
      19607: inst = 32'h8220000;
      19608: inst = 32'h10408000;
      19609: inst = 32'hc404972;
      19610: inst = 32'h8220000;
      19611: inst = 32'h10408000;
      19612: inst = 32'hc404973;
      19613: inst = 32'h8220000;
      19614: inst = 32'h10408000;
      19615: inst = 32'hc404974;
      19616: inst = 32'h8220000;
      19617: inst = 32'h10408000;
      19618: inst = 32'hc404975;
      19619: inst = 32'h8220000;
      19620: inst = 32'h10408000;
      19621: inst = 32'hc404976;
      19622: inst = 32'h8220000;
      19623: inst = 32'h10408000;
      19624: inst = 32'hc404977;
      19625: inst = 32'h8220000;
      19626: inst = 32'h10408000;
      19627: inst = 32'hc404978;
      19628: inst = 32'h8220000;
      19629: inst = 32'h10408000;
      19630: inst = 32'hc404979;
      19631: inst = 32'h8220000;
      19632: inst = 32'h10408000;
      19633: inst = 32'hc40497d;
      19634: inst = 32'h8220000;
      19635: inst = 32'h10408000;
      19636: inst = 32'hc40497e;
      19637: inst = 32'h8220000;
      19638: inst = 32'h10408000;
      19639: inst = 32'hc40497f;
      19640: inst = 32'h8220000;
      19641: inst = 32'h10408000;
      19642: inst = 32'hc404980;
      19643: inst = 32'h8220000;
      19644: inst = 32'h10408000;
      19645: inst = 32'hc404981;
      19646: inst = 32'h8220000;
      19647: inst = 32'h10408000;
      19648: inst = 32'hc404982;
      19649: inst = 32'h8220000;
      19650: inst = 32'h10408000;
      19651: inst = 32'hc404983;
      19652: inst = 32'h8220000;
      19653: inst = 32'h10408000;
      19654: inst = 32'hc404984;
      19655: inst = 32'h8220000;
      19656: inst = 32'h10408000;
      19657: inst = 32'hc404985;
      19658: inst = 32'h8220000;
      19659: inst = 32'h10408000;
      19660: inst = 32'hc404986;
      19661: inst = 32'h8220000;
      19662: inst = 32'h10408000;
      19663: inst = 32'hc404987;
      19664: inst = 32'h8220000;
      19665: inst = 32'h10408000;
      19666: inst = 32'hc404989;
      19667: inst = 32'h8220000;
      19668: inst = 32'h10408000;
      19669: inst = 32'hc40498a;
      19670: inst = 32'h8220000;
      19671: inst = 32'h10408000;
      19672: inst = 32'hc40498b;
      19673: inst = 32'h8220000;
      19674: inst = 32'h10408000;
      19675: inst = 32'hc40498c;
      19676: inst = 32'h8220000;
      19677: inst = 32'h10408000;
      19678: inst = 32'hc40498d;
      19679: inst = 32'h8220000;
      19680: inst = 32'h10408000;
      19681: inst = 32'hc40498e;
      19682: inst = 32'h8220000;
      19683: inst = 32'h10408000;
      19684: inst = 32'hc40498f;
      19685: inst = 32'h8220000;
      19686: inst = 32'h10408000;
      19687: inst = 32'hc404990;
      19688: inst = 32'h8220000;
      19689: inst = 32'h10408000;
      19690: inst = 32'hc404991;
      19691: inst = 32'h8220000;
      19692: inst = 32'h10408000;
      19693: inst = 32'hc404992;
      19694: inst = 32'h8220000;
      19695: inst = 32'h10408000;
      19696: inst = 32'hc404993;
      19697: inst = 32'h8220000;
      19698: inst = 32'h10408000;
      19699: inst = 32'hc404dcd;
      19700: inst = 32'h8220000;
      19701: inst = 32'h10408000;
      19702: inst = 32'hc404dce;
      19703: inst = 32'h8220000;
      19704: inst = 32'h10408000;
      19705: inst = 32'hc404dcf;
      19706: inst = 32'h8220000;
      19707: inst = 32'h10408000;
      19708: inst = 32'hc404dd0;
      19709: inst = 32'h8220000;
      19710: inst = 32'h10408000;
      19711: inst = 32'hc404dd1;
      19712: inst = 32'h8220000;
      19713: inst = 32'h10408000;
      19714: inst = 32'hc404dd2;
      19715: inst = 32'h8220000;
      19716: inst = 32'h10408000;
      19717: inst = 32'hc404dd3;
      19718: inst = 32'h8220000;
      19719: inst = 32'h10408000;
      19720: inst = 32'hc404dd4;
      19721: inst = 32'h8220000;
      19722: inst = 32'h10408000;
      19723: inst = 32'hc404dd5;
      19724: inst = 32'h8220000;
      19725: inst = 32'h10408000;
      19726: inst = 32'hc404dd7;
      19727: inst = 32'h8220000;
      19728: inst = 32'h10408000;
      19729: inst = 32'hc404dd8;
      19730: inst = 32'h8220000;
      19731: inst = 32'h10408000;
      19732: inst = 32'hc404dd9;
      19733: inst = 32'h8220000;
      19734: inst = 32'h10408000;
      19735: inst = 32'hc404dda;
      19736: inst = 32'h8220000;
      19737: inst = 32'h10408000;
      19738: inst = 32'hc404ddb;
      19739: inst = 32'h8220000;
      19740: inst = 32'h10408000;
      19741: inst = 32'hc404ddc;
      19742: inst = 32'h8220000;
      19743: inst = 32'h10408000;
      19744: inst = 32'hc404ddd;
      19745: inst = 32'h8220000;
      19746: inst = 32'h10408000;
      19747: inst = 32'hc404dde;
      19748: inst = 32'h8220000;
      19749: inst = 32'h10408000;
      19750: inst = 32'hc404ddf;
      19751: inst = 32'h8220000;
      19752: inst = 32'h10408000;
      19753: inst = 32'hc404de0;
      19754: inst = 32'h8220000;
      19755: inst = 32'h10408000;
      19756: inst = 32'hc404de1;
      19757: inst = 32'h8220000;
      19758: inst = 32'h10408000;
      19759: inst = 32'hc404de2;
      19760: inst = 32'h8220000;
      19761: inst = 32'h10408000;
      19762: inst = 32'hc404de4;
      19763: inst = 32'h8220000;
      19764: inst = 32'h10408000;
      19765: inst = 32'hc404de5;
      19766: inst = 32'h8220000;
      19767: inst = 32'h10408000;
      19768: inst = 32'hc404de6;
      19769: inst = 32'h8220000;
      19770: inst = 32'h10408000;
      19771: inst = 32'hc404de7;
      19772: inst = 32'h8220000;
      19773: inst = 32'h10408000;
      19774: inst = 32'hc404de8;
      19775: inst = 32'h8220000;
      19776: inst = 32'h10408000;
      19777: inst = 32'hc404de9;
      19778: inst = 32'h8220000;
      19779: inst = 32'h10408000;
      19780: inst = 32'hc404dea;
      19781: inst = 32'h8220000;
      19782: inst = 32'h10408000;
      19783: inst = 32'hc404deb;
      19784: inst = 32'h8220000;
      19785: inst = 32'h10408000;
      19786: inst = 32'hc404dec;
      19787: inst = 32'h8220000;
      19788: inst = 32'h10408000;
      19789: inst = 32'hc404ded;
      19790: inst = 32'h8220000;
      19791: inst = 32'h10408000;
      19792: inst = 32'hc404df0;
      19793: inst = 32'h8220000;
      19794: inst = 32'h10408000;
      19795: inst = 32'hc404df1;
      19796: inst = 32'h8220000;
      19797: inst = 32'h10408000;
      19798: inst = 32'hc404df2;
      19799: inst = 32'h8220000;
      19800: inst = 32'h10408000;
      19801: inst = 32'hc404dfc;
      19802: inst = 32'h8220000;
      19803: inst = 32'h10408000;
      19804: inst = 32'hc404dfd;
      19805: inst = 32'h8220000;
      19806: inst = 32'h10408000;
      19807: inst = 32'hc404dfe;
      19808: inst = 32'h8220000;
      19809: inst = 32'h10408000;
      19810: inst = 32'hc404dff;
      19811: inst = 32'h8220000;
      19812: inst = 32'h10408000;
      19813: inst = 32'hc404e00;
      19814: inst = 32'h8220000;
      19815: inst = 32'h10408000;
      19816: inst = 32'hc404e01;
      19817: inst = 32'h8220000;
      19818: inst = 32'h10408000;
      19819: inst = 32'hc404e02;
      19820: inst = 32'h8220000;
      19821: inst = 32'h10408000;
      19822: inst = 32'hc404e03;
      19823: inst = 32'h8220000;
      19824: inst = 32'h10408000;
      19825: inst = 32'hc404e04;
      19826: inst = 32'h8220000;
      19827: inst = 32'h10408000;
      19828: inst = 32'hc404e05;
      19829: inst = 32'h8220000;
      19830: inst = 32'h10408000;
      19831: inst = 32'hc404e06;
      19832: inst = 32'h8220000;
      19833: inst = 32'h10408000;
      19834: inst = 32'hc404e07;
      19835: inst = 32'h8220000;
      19836: inst = 32'h10408000;
      19837: inst = 32'hc404e0b;
      19838: inst = 32'h8220000;
      19839: inst = 32'h10408000;
      19840: inst = 32'hc404e0c;
      19841: inst = 32'h8220000;
      19842: inst = 32'h10408000;
      19843: inst = 32'hc404e0d;
      19844: inst = 32'h8220000;
      19845: inst = 32'h10408000;
      19846: inst = 32'hc404e0e;
      19847: inst = 32'h8220000;
      19848: inst = 32'h10408000;
      19849: inst = 32'hc404e0f;
      19850: inst = 32'h8220000;
      19851: inst = 32'h10408000;
      19852: inst = 32'hc404e10;
      19853: inst = 32'h8220000;
      19854: inst = 32'h10408000;
      19855: inst = 32'hc404e11;
      19856: inst = 32'h8220000;
      19857: inst = 32'h10408000;
      19858: inst = 32'hc404e12;
      19859: inst = 32'h8220000;
      19860: inst = 32'h10408000;
      19861: inst = 32'hc404e13;
      19862: inst = 32'h8220000;
      19863: inst = 32'h10408000;
      19864: inst = 32'hc404e2c;
      19865: inst = 32'h8220000;
      19866: inst = 32'h10408000;
      19867: inst = 32'hc404e2d;
      19868: inst = 32'h8220000;
      19869: inst = 32'h10408000;
      19870: inst = 32'hc404e2e;
      19871: inst = 32'h8220000;
      19872: inst = 32'h10408000;
      19873: inst = 32'hc404e2f;
      19874: inst = 32'h8220000;
      19875: inst = 32'h10408000;
      19876: inst = 32'hc404e30;
      19877: inst = 32'h8220000;
      19878: inst = 32'h10408000;
      19879: inst = 32'hc404e31;
      19880: inst = 32'h8220000;
      19881: inst = 32'h10408000;
      19882: inst = 32'hc404e32;
      19883: inst = 32'h8220000;
      19884: inst = 32'h10408000;
      19885: inst = 32'hc404e33;
      19886: inst = 32'h8220000;
      19887: inst = 32'h10408000;
      19888: inst = 32'hc404e34;
      19889: inst = 32'h8220000;
      19890: inst = 32'h10408000;
      19891: inst = 32'hc404e35;
      19892: inst = 32'h8220000;
      19893: inst = 32'h10408000;
      19894: inst = 32'hc404e38;
      19895: inst = 32'h8220000;
      19896: inst = 32'h10408000;
      19897: inst = 32'hc404e39;
      19898: inst = 32'h8220000;
      19899: inst = 32'h10408000;
      19900: inst = 32'hc404e3a;
      19901: inst = 32'h8220000;
      19902: inst = 32'h10408000;
      19903: inst = 32'hc404e3b;
      19904: inst = 32'h8220000;
      19905: inst = 32'h10408000;
      19906: inst = 32'hc404e3c;
      19907: inst = 32'h8220000;
      19908: inst = 32'h10408000;
      19909: inst = 32'hc404e3d;
      19910: inst = 32'h8220000;
      19911: inst = 32'h10408000;
      19912: inst = 32'hc404e3e;
      19913: inst = 32'h8220000;
      19914: inst = 32'h10408000;
      19915: inst = 32'hc404e3f;
      19916: inst = 32'h8220000;
      19917: inst = 32'h10408000;
      19918: inst = 32'hc404e40;
      19919: inst = 32'h8220000;
      19920: inst = 32'h10408000;
      19921: inst = 32'hc404e41;
      19922: inst = 32'h8220000;
      19923: inst = 32'h10408000;
      19924: inst = 32'hc404e42;
      19925: inst = 32'h8220000;
      19926: inst = 32'h10408000;
      19927: inst = 32'hc404e44;
      19928: inst = 32'h8220000;
      19929: inst = 32'h10408000;
      19930: inst = 32'hc404e45;
      19931: inst = 32'h8220000;
      19932: inst = 32'h10408000;
      19933: inst = 32'hc404e46;
      19934: inst = 32'h8220000;
      19935: inst = 32'h10408000;
      19936: inst = 32'hc404e47;
      19937: inst = 32'h8220000;
      19938: inst = 32'h10408000;
      19939: inst = 32'hc404e48;
      19940: inst = 32'h8220000;
      19941: inst = 32'h10408000;
      19942: inst = 32'hc404e49;
      19943: inst = 32'h8220000;
      19944: inst = 32'h10408000;
      19945: inst = 32'hc404e4a;
      19946: inst = 32'h8220000;
      19947: inst = 32'h10408000;
      19948: inst = 32'hc404e4b;
      19949: inst = 32'h8220000;
      19950: inst = 32'h10408000;
      19951: inst = 32'hc404e4c;
      19952: inst = 32'h8220000;
      19953: inst = 32'h10408000;
      19954: inst = 32'hc404e4d;
      19955: inst = 32'h8220000;
      19956: inst = 32'h10408000;
      19957: inst = 32'hc404e50;
      19958: inst = 32'h8220000;
      19959: inst = 32'h10408000;
      19960: inst = 32'hc404e51;
      19961: inst = 32'h8220000;
      19962: inst = 32'h10408000;
      19963: inst = 32'hc404e52;
      19964: inst = 32'h8220000;
      19965: inst = 32'h10408000;
      19966: inst = 32'hc404e53;
      19967: inst = 32'h8220000;
      19968: inst = 32'h10408000;
      19969: inst = 32'hc404e5c;
      19970: inst = 32'h8220000;
      19971: inst = 32'h10408000;
      19972: inst = 32'hc404e5d;
      19973: inst = 32'h8220000;
      19974: inst = 32'h10408000;
      19975: inst = 32'hc404e5e;
      19976: inst = 32'h8220000;
      19977: inst = 32'h10408000;
      19978: inst = 32'hc404e5f;
      19979: inst = 32'h8220000;
      19980: inst = 32'h10408000;
      19981: inst = 32'hc404e60;
      19982: inst = 32'h8220000;
      19983: inst = 32'h10408000;
      19984: inst = 32'hc404e61;
      19985: inst = 32'h8220000;
      19986: inst = 32'h10408000;
      19987: inst = 32'hc404e62;
      19988: inst = 32'h8220000;
      19989: inst = 32'h10408000;
      19990: inst = 32'hc404e63;
      19991: inst = 32'h8220000;
      19992: inst = 32'h10408000;
      19993: inst = 32'hc404e64;
      19994: inst = 32'h8220000;
      19995: inst = 32'h10408000;
      19996: inst = 32'hc404e65;
      19997: inst = 32'h8220000;
      19998: inst = 32'h10408000;
      19999: inst = 32'hc404e66;
      20000: inst = 32'h8220000;
      20001: inst = 32'h10408000;
      20002: inst = 32'hc404e6a;
      20003: inst = 32'h8220000;
      20004: inst = 32'h10408000;
      20005: inst = 32'hc404e6b;
      20006: inst = 32'h8220000;
      20007: inst = 32'h10408000;
      20008: inst = 32'hc404e6c;
      20009: inst = 32'h8220000;
      20010: inst = 32'h10408000;
      20011: inst = 32'hc404e6d;
      20012: inst = 32'h8220000;
      20013: inst = 32'h10408000;
      20014: inst = 32'hc404e6e;
      20015: inst = 32'h8220000;
      20016: inst = 32'h10408000;
      20017: inst = 32'hc404e6f;
      20018: inst = 32'h8220000;
      20019: inst = 32'h10408000;
      20020: inst = 32'hc404e70;
      20021: inst = 32'h8220000;
      20022: inst = 32'h10408000;
      20023: inst = 32'hc404e71;
      20024: inst = 32'h8220000;
      20025: inst = 32'h10408000;
      20026: inst = 32'hc404e72;
      20027: inst = 32'h8220000;
      20028: inst = 32'h10408000;
      20029: inst = 32'hc404e73;
      20030: inst = 32'h8220000;
      20031: inst = 32'h10408000;
      20032: inst = 32'hc404e8b;
      20033: inst = 32'h8220000;
      20034: inst = 32'h10408000;
      20035: inst = 32'hc404e8c;
      20036: inst = 32'h8220000;
      20037: inst = 32'h10408000;
      20038: inst = 32'hc404e8d;
      20039: inst = 32'h8220000;
      20040: inst = 32'h10408000;
      20041: inst = 32'hc404e99;
      20042: inst = 32'h8220000;
      20043: inst = 32'h10408000;
      20044: inst = 32'hc404e9a;
      20045: inst = 32'h8220000;
      20046: inst = 32'h10408000;
      20047: inst = 32'hc404e9b;
      20048: inst = 32'h8220000;
      20049: inst = 32'h10408000;
      20050: inst = 32'hc404e9c;
      20051: inst = 32'h8220000;
      20052: inst = 32'h10408000;
      20053: inst = 32'hc404ea4;
      20054: inst = 32'h8220000;
      20055: inst = 32'h10408000;
      20056: inst = 32'hc404ea5;
      20057: inst = 32'h8220000;
      20058: inst = 32'h10408000;
      20059: inst = 32'hc404eac;
      20060: inst = 32'h8220000;
      20061: inst = 32'h10408000;
      20062: inst = 32'hc404ead;
      20063: inst = 32'h8220000;
      20064: inst = 32'h10408000;
      20065: inst = 32'hc404eb0;
      20066: inst = 32'h8220000;
      20067: inst = 32'h10408000;
      20068: inst = 32'hc404eb1;
      20069: inst = 32'h8220000;
      20070: inst = 32'h10408000;
      20071: inst = 32'hc404eb2;
      20072: inst = 32'h8220000;
      20073: inst = 32'h10408000;
      20074: inst = 32'hc404eb3;
      20075: inst = 32'h8220000;
      20076: inst = 32'h10408000;
      20077: inst = 32'hc404eb4;
      20078: inst = 32'h8220000;
      20079: inst = 32'h10408000;
      20080: inst = 32'hc404ebc;
      20081: inst = 32'h8220000;
      20082: inst = 32'h10408000;
      20083: inst = 32'hc404ebd;
      20084: inst = 32'h8220000;
      20085: inst = 32'h10408000;
      20086: inst = 32'hc404ec2;
      20087: inst = 32'h8220000;
      20088: inst = 32'h10408000;
      20089: inst = 32'hc404ec3;
      20090: inst = 32'h8220000;
      20091: inst = 32'h10408000;
      20092: inst = 32'hc404ec4;
      20093: inst = 32'h8220000;
      20094: inst = 32'h10408000;
      20095: inst = 32'hc404ec5;
      20096: inst = 32'h8220000;
      20097: inst = 32'h10408000;
      20098: inst = 32'hc404ec9;
      20099: inst = 32'h8220000;
      20100: inst = 32'h10408000;
      20101: inst = 32'hc404eca;
      20102: inst = 32'h8220000;
      20103: inst = 32'h10408000;
      20104: inst = 32'hc404eeb;
      20105: inst = 32'h8220000;
      20106: inst = 32'h10408000;
      20107: inst = 32'hc404eec;
      20108: inst = 32'h8220000;
      20109: inst = 32'h10408000;
      20110: inst = 32'hc404efa;
      20111: inst = 32'h8220000;
      20112: inst = 32'h10408000;
      20113: inst = 32'hc404efb;
      20114: inst = 32'h8220000;
      20115: inst = 32'h10408000;
      20116: inst = 32'hc404efc;
      20117: inst = 32'h8220000;
      20118: inst = 32'h10408000;
      20119: inst = 32'hc404f04;
      20120: inst = 32'h8220000;
      20121: inst = 32'h10408000;
      20122: inst = 32'hc404f05;
      20123: inst = 32'h8220000;
      20124: inst = 32'h10408000;
      20125: inst = 32'hc404f0c;
      20126: inst = 32'h8220000;
      20127: inst = 32'h10408000;
      20128: inst = 32'hc404f0d;
      20129: inst = 32'h8220000;
      20130: inst = 32'h10408000;
      20131: inst = 32'hc404f10;
      20132: inst = 32'h8220000;
      20133: inst = 32'h10408000;
      20134: inst = 32'hc404f12;
      20135: inst = 32'h8220000;
      20136: inst = 32'h10408000;
      20137: inst = 32'hc404f13;
      20138: inst = 32'h8220000;
      20139: inst = 32'h10408000;
      20140: inst = 32'hc404f14;
      20141: inst = 32'h8220000;
      20142: inst = 32'h10408000;
      20143: inst = 32'hc404f15;
      20144: inst = 32'h8220000;
      20145: inst = 32'h10408000;
      20146: inst = 32'hc404f1c;
      20147: inst = 32'h8220000;
      20148: inst = 32'h10408000;
      20149: inst = 32'hc404f1d;
      20150: inst = 32'h8220000;
      20151: inst = 32'h10408000;
      20152: inst = 32'hc404f22;
      20153: inst = 32'h8220000;
      20154: inst = 32'h10408000;
      20155: inst = 32'hc404f23;
      20156: inst = 32'h8220000;
      20157: inst = 32'h10408000;
      20158: inst = 32'hc404f24;
      20159: inst = 32'h8220000;
      20160: inst = 32'h10408000;
      20161: inst = 32'hc404f29;
      20162: inst = 32'h8220000;
      20163: inst = 32'h10408000;
      20164: inst = 32'hc404f2a;
      20165: inst = 32'h8220000;
      20166: inst = 32'h10408000;
      20167: inst = 32'hc404f4b;
      20168: inst = 32'h8220000;
      20169: inst = 32'h10408000;
      20170: inst = 32'hc404f4c;
      20171: inst = 32'h8220000;
      20172: inst = 32'h10408000;
      20173: inst = 32'hc404f4e;
      20174: inst = 32'h8220000;
      20175: inst = 32'h10408000;
      20176: inst = 32'hc404f4f;
      20177: inst = 32'h8220000;
      20178: inst = 32'h10408000;
      20179: inst = 32'hc404f50;
      20180: inst = 32'h8220000;
      20181: inst = 32'h10408000;
      20182: inst = 32'hc404f51;
      20183: inst = 32'h8220000;
      20184: inst = 32'h10408000;
      20185: inst = 32'hc404f52;
      20186: inst = 32'h8220000;
      20187: inst = 32'h10408000;
      20188: inst = 32'hc404f5b;
      20189: inst = 32'h8220000;
      20190: inst = 32'h10408000;
      20191: inst = 32'hc404f5c;
      20192: inst = 32'h8220000;
      20193: inst = 32'h10408000;
      20194: inst = 32'hc404f5d;
      20195: inst = 32'h8220000;
      20196: inst = 32'h10408000;
      20197: inst = 32'hc404f64;
      20198: inst = 32'h8220000;
      20199: inst = 32'h10408000;
      20200: inst = 32'hc404f65;
      20201: inst = 32'h8220000;
      20202: inst = 32'h10408000;
      20203: inst = 32'hc404f6c;
      20204: inst = 32'h8220000;
      20205: inst = 32'h10408000;
      20206: inst = 32'hc404f70;
      20207: inst = 32'h8220000;
      20208: inst = 32'h10408000;
      20209: inst = 32'hc404f71;
      20210: inst = 32'h8220000;
      20211: inst = 32'h10408000;
      20212: inst = 32'hc404f72;
      20213: inst = 32'h8220000;
      20214: inst = 32'h10408000;
      20215: inst = 32'hc404f73;
      20216: inst = 32'h8220000;
      20217: inst = 32'h10408000;
      20218: inst = 32'hc404f74;
      20219: inst = 32'h8220000;
      20220: inst = 32'h10408000;
      20221: inst = 32'hc404f75;
      20222: inst = 32'h8220000;
      20223: inst = 32'h10408000;
      20224: inst = 32'hc404f76;
      20225: inst = 32'h8220000;
      20226: inst = 32'h10408000;
      20227: inst = 32'hc404f7c;
      20228: inst = 32'h8220000;
      20229: inst = 32'h10408000;
      20230: inst = 32'hc404f7d;
      20231: inst = 32'h8220000;
      20232: inst = 32'h10408000;
      20233: inst = 32'hc404f7f;
      20234: inst = 32'h8220000;
      20235: inst = 32'h10408000;
      20236: inst = 32'hc404f80;
      20237: inst = 32'h8220000;
      20238: inst = 32'h10408000;
      20239: inst = 32'hc404f81;
      20240: inst = 32'h8220000;
      20241: inst = 32'h10408000;
      20242: inst = 32'hc404f82;
      20243: inst = 32'h8220000;
      20244: inst = 32'h10408000;
      20245: inst = 32'hc404f83;
      20246: inst = 32'h8220000;
      20247: inst = 32'h10408000;
      20248: inst = 32'hc404f89;
      20249: inst = 32'h8220000;
      20250: inst = 32'h10408000;
      20251: inst = 32'hc404f8a;
      20252: inst = 32'h8220000;
      20253: inst = 32'h10408000;
      20254: inst = 32'hc404f8c;
      20255: inst = 32'h8220000;
      20256: inst = 32'h10408000;
      20257: inst = 32'hc404f8d;
      20258: inst = 32'h8220000;
      20259: inst = 32'h10408000;
      20260: inst = 32'hc404f8e;
      20261: inst = 32'h8220000;
      20262: inst = 32'h10408000;
      20263: inst = 32'hc404f8f;
      20264: inst = 32'h8220000;
      20265: inst = 32'h10408000;
      20266: inst = 32'hc404f90;
      20267: inst = 32'h8220000;
      20268: inst = 32'h10408000;
      20269: inst = 32'hc404fab;
      20270: inst = 32'h8220000;
      20271: inst = 32'h10408000;
      20272: inst = 32'hc404fac;
      20273: inst = 32'h8220000;
      20274: inst = 32'h10408000;
      20275: inst = 32'hc404fae;
      20276: inst = 32'h8220000;
      20277: inst = 32'h10408000;
      20278: inst = 32'hc404faf;
      20279: inst = 32'h8220000;
      20280: inst = 32'h10408000;
      20281: inst = 32'hc404fb0;
      20282: inst = 32'h8220000;
      20283: inst = 32'h10408000;
      20284: inst = 32'hc404fb1;
      20285: inst = 32'h8220000;
      20286: inst = 32'h10408000;
      20287: inst = 32'hc404fb2;
      20288: inst = 32'h8220000;
      20289: inst = 32'h10408000;
      20290: inst = 32'hc404fbc;
      20291: inst = 32'h8220000;
      20292: inst = 32'h10408000;
      20293: inst = 32'hc404fbd;
      20294: inst = 32'h8220000;
      20295: inst = 32'h10408000;
      20296: inst = 32'hc404fbe;
      20297: inst = 32'h8220000;
      20298: inst = 32'h10408000;
      20299: inst = 32'hc404fc4;
      20300: inst = 32'h8220000;
      20301: inst = 32'h10408000;
      20302: inst = 32'hc404fc5;
      20303: inst = 32'h8220000;
      20304: inst = 32'h10408000;
      20305: inst = 32'hc404fd0;
      20306: inst = 32'h8220000;
      20307: inst = 32'h10408000;
      20308: inst = 32'hc404fd1;
      20309: inst = 32'h8220000;
      20310: inst = 32'h10408000;
      20311: inst = 32'hc404fd2;
      20312: inst = 32'h8220000;
      20313: inst = 32'h10408000;
      20314: inst = 32'hc404fd4;
      20315: inst = 32'h8220000;
      20316: inst = 32'h10408000;
      20317: inst = 32'hc404fd5;
      20318: inst = 32'h8220000;
      20319: inst = 32'h10408000;
      20320: inst = 32'hc404fd6;
      20321: inst = 32'h8220000;
      20322: inst = 32'h10408000;
      20323: inst = 32'hc404fd7;
      20324: inst = 32'h8220000;
      20325: inst = 32'h10408000;
      20326: inst = 32'hc404fdc;
      20327: inst = 32'h8220000;
      20328: inst = 32'h10408000;
      20329: inst = 32'hc404fdd;
      20330: inst = 32'h8220000;
      20331: inst = 32'h10408000;
      20332: inst = 32'hc404fdf;
      20333: inst = 32'h8220000;
      20334: inst = 32'h10408000;
      20335: inst = 32'hc404fe0;
      20336: inst = 32'h8220000;
      20337: inst = 32'h10408000;
      20338: inst = 32'hc404fe1;
      20339: inst = 32'h8220000;
      20340: inst = 32'h10408000;
      20341: inst = 32'hc404fe2;
      20342: inst = 32'h8220000;
      20343: inst = 32'h10408000;
      20344: inst = 32'hc404fe9;
      20345: inst = 32'h8220000;
      20346: inst = 32'h10408000;
      20347: inst = 32'hc404fea;
      20348: inst = 32'h8220000;
      20349: inst = 32'h10408000;
      20350: inst = 32'hc404fec;
      20351: inst = 32'h8220000;
      20352: inst = 32'h10408000;
      20353: inst = 32'hc404fed;
      20354: inst = 32'h8220000;
      20355: inst = 32'h10408000;
      20356: inst = 32'hc404fee;
      20357: inst = 32'h8220000;
      20358: inst = 32'h10408000;
      20359: inst = 32'hc404fef;
      20360: inst = 32'h8220000;
      20361: inst = 32'h10408000;
      20362: inst = 32'hc404ff0;
      20363: inst = 32'h8220000;
      20364: inst = 32'h10408000;
      20365: inst = 32'hc40500b;
      20366: inst = 32'h8220000;
      20367: inst = 32'h10408000;
      20368: inst = 32'hc40500c;
      20369: inst = 32'h8220000;
      20370: inst = 32'h10408000;
      20371: inst = 32'hc40501d;
      20372: inst = 32'h8220000;
      20373: inst = 32'h10408000;
      20374: inst = 32'hc40501e;
      20375: inst = 32'h8220000;
      20376: inst = 32'h10408000;
      20377: inst = 32'hc40501f;
      20378: inst = 32'h8220000;
      20379: inst = 32'h10408000;
      20380: inst = 32'hc405024;
      20381: inst = 32'h8220000;
      20382: inst = 32'h10408000;
      20383: inst = 32'hc405025;
      20384: inst = 32'h8220000;
      20385: inst = 32'h10408000;
      20386: inst = 32'hc405030;
      20387: inst = 32'h8220000;
      20388: inst = 32'h10408000;
      20389: inst = 32'hc405031;
      20390: inst = 32'h8220000;
      20391: inst = 32'h10408000;
      20392: inst = 32'hc405032;
      20393: inst = 32'h8220000;
      20394: inst = 32'h10408000;
      20395: inst = 32'hc405033;
      20396: inst = 32'h8220000;
      20397: inst = 32'h10408000;
      20398: inst = 32'hc405034;
      20399: inst = 32'h8220000;
      20400: inst = 32'h10408000;
      20401: inst = 32'hc405035;
      20402: inst = 32'h8220000;
      20403: inst = 32'h10408000;
      20404: inst = 32'hc405036;
      20405: inst = 32'h8220000;
      20406: inst = 32'h10408000;
      20407: inst = 32'hc405037;
      20408: inst = 32'h8220000;
      20409: inst = 32'h10408000;
      20410: inst = 32'hc405038;
      20411: inst = 32'h8220000;
      20412: inst = 32'h10408000;
      20413: inst = 32'hc40503c;
      20414: inst = 32'h8220000;
      20415: inst = 32'h10408000;
      20416: inst = 32'hc40503d;
      20417: inst = 32'h8220000;
      20418: inst = 32'h10408000;
      20419: inst = 32'hc405049;
      20420: inst = 32'h8220000;
      20421: inst = 32'h10408000;
      20422: inst = 32'hc40504a;
      20423: inst = 32'h8220000;
      20424: inst = 32'h10408000;
      20425: inst = 32'hc40506b;
      20426: inst = 32'h8220000;
      20427: inst = 32'h10408000;
      20428: inst = 32'hc40506c;
      20429: inst = 32'h8220000;
      20430: inst = 32'h10408000;
      20431: inst = 32'hc40506d;
      20432: inst = 32'h8220000;
      20433: inst = 32'h10408000;
      20434: inst = 32'hc40506e;
      20435: inst = 32'h8220000;
      20436: inst = 32'h10408000;
      20437: inst = 32'hc40506f;
      20438: inst = 32'h8220000;
      20439: inst = 32'h10408000;
      20440: inst = 32'hc405070;
      20441: inst = 32'h8220000;
      20442: inst = 32'h10408000;
      20443: inst = 32'hc405071;
      20444: inst = 32'h8220000;
      20445: inst = 32'h10408000;
      20446: inst = 32'hc405072;
      20447: inst = 32'h8220000;
      20448: inst = 32'h10408000;
      20449: inst = 32'hc405073;
      20450: inst = 32'h8220000;
      20451: inst = 32'h10408000;
      20452: inst = 32'hc405074;
      20453: inst = 32'h8220000;
      20454: inst = 32'h10408000;
      20455: inst = 32'hc405075;
      20456: inst = 32'h8220000;
      20457: inst = 32'h10408000;
      20458: inst = 32'hc405077;
      20459: inst = 32'h8220000;
      20460: inst = 32'h10408000;
      20461: inst = 32'hc405078;
      20462: inst = 32'h8220000;
      20463: inst = 32'h10408000;
      20464: inst = 32'hc405079;
      20465: inst = 32'h8220000;
      20466: inst = 32'h10408000;
      20467: inst = 32'hc40507a;
      20468: inst = 32'h8220000;
      20469: inst = 32'h10408000;
      20470: inst = 32'hc40507b;
      20471: inst = 32'h8220000;
      20472: inst = 32'h10408000;
      20473: inst = 32'hc40507c;
      20474: inst = 32'h8220000;
      20475: inst = 32'h10408000;
      20476: inst = 32'hc40507d;
      20477: inst = 32'h8220000;
      20478: inst = 32'h10408000;
      20479: inst = 32'hc40507e;
      20480: inst = 32'h8220000;
      20481: inst = 32'h10408000;
      20482: inst = 32'hc40507f;
      20483: inst = 32'h8220000;
      20484: inst = 32'h10408000;
      20485: inst = 32'hc405080;
      20486: inst = 32'h8220000;
      20487: inst = 32'h10408000;
      20488: inst = 32'hc405084;
      20489: inst = 32'h8220000;
      20490: inst = 32'h10408000;
      20491: inst = 32'hc405085;
      20492: inst = 32'h8220000;
      20493: inst = 32'h10408000;
      20494: inst = 32'hc405086;
      20495: inst = 32'h8220000;
      20496: inst = 32'h10408000;
      20497: inst = 32'hc405087;
      20498: inst = 32'h8220000;
      20499: inst = 32'h10408000;
      20500: inst = 32'hc405088;
      20501: inst = 32'h8220000;
      20502: inst = 32'h10408000;
      20503: inst = 32'hc405089;
      20504: inst = 32'h8220000;
      20505: inst = 32'h10408000;
      20506: inst = 32'hc40508a;
      20507: inst = 32'h8220000;
      20508: inst = 32'h10408000;
      20509: inst = 32'hc40508b;
      20510: inst = 32'h8220000;
      20511: inst = 32'h10408000;
      20512: inst = 32'hc40508c;
      20513: inst = 32'h8220000;
      20514: inst = 32'h10408000;
      20515: inst = 32'hc40508d;
      20516: inst = 32'h8220000;
      20517: inst = 32'h10408000;
      20518: inst = 32'hc405090;
      20519: inst = 32'h8220000;
      20520: inst = 32'h10408000;
      20521: inst = 32'hc405091;
      20522: inst = 32'h8220000;
      20523: inst = 32'h10408000;
      20524: inst = 32'hc405096;
      20525: inst = 32'h8220000;
      20526: inst = 32'h10408000;
      20527: inst = 32'hc405097;
      20528: inst = 32'h8220000;
      20529: inst = 32'h10408000;
      20530: inst = 32'hc405098;
      20531: inst = 32'h8220000;
      20532: inst = 32'h10408000;
      20533: inst = 32'hc405099;
      20534: inst = 32'h8220000;
      20535: inst = 32'h10408000;
      20536: inst = 32'hc40509c;
      20537: inst = 32'h8220000;
      20538: inst = 32'h10408000;
      20539: inst = 32'hc40509d;
      20540: inst = 32'h8220000;
      20541: inst = 32'h10408000;
      20542: inst = 32'hc4050a9;
      20543: inst = 32'h8220000;
      20544: inst = 32'h10408000;
      20545: inst = 32'hc4050aa;
      20546: inst = 32'h8220000;
      20547: inst = 32'h10408000;
      20548: inst = 32'hc4050ab;
      20549: inst = 32'h8220000;
      20550: inst = 32'h10408000;
      20551: inst = 32'hc4050ac;
      20552: inst = 32'h8220000;
      20553: inst = 32'h10408000;
      20554: inst = 32'hc4050ad;
      20555: inst = 32'h8220000;
      20556: inst = 32'h10408000;
      20557: inst = 32'hc4050ae;
      20558: inst = 32'h8220000;
      20559: inst = 32'h10408000;
      20560: inst = 32'hc4050af;
      20561: inst = 32'h8220000;
      20562: inst = 32'h10408000;
      20563: inst = 32'hc4050b0;
      20564: inst = 32'h8220000;
      20565: inst = 32'h10408000;
      20566: inst = 32'hc4050b1;
      20567: inst = 32'h8220000;
      20568: inst = 32'h10408000;
      20569: inst = 32'hc4050b2;
      20570: inst = 32'h8220000;
      20571: inst = 32'h10408000;
      20572: inst = 32'hc4050b3;
      20573: inst = 32'h8220000;
      20574: inst = 32'h10408000;
      20575: inst = 32'hc4050cb;
      20576: inst = 32'h8220000;
      20577: inst = 32'h10408000;
      20578: inst = 32'hc4050cc;
      20579: inst = 32'h8220000;
      20580: inst = 32'h10408000;
      20581: inst = 32'hc4050cd;
      20582: inst = 32'h8220000;
      20583: inst = 32'h10408000;
      20584: inst = 32'hc4050ce;
      20585: inst = 32'h8220000;
      20586: inst = 32'h10408000;
      20587: inst = 32'hc4050cf;
      20588: inst = 32'h8220000;
      20589: inst = 32'h10408000;
      20590: inst = 32'hc4050d0;
      20591: inst = 32'h8220000;
      20592: inst = 32'h10408000;
      20593: inst = 32'hc4050d1;
      20594: inst = 32'h8220000;
      20595: inst = 32'h10408000;
      20596: inst = 32'hc4050d2;
      20597: inst = 32'h8220000;
      20598: inst = 32'h10408000;
      20599: inst = 32'hc4050d3;
      20600: inst = 32'h8220000;
      20601: inst = 32'h10408000;
      20602: inst = 32'hc4050d4;
      20603: inst = 32'h8220000;
      20604: inst = 32'h10408000;
      20605: inst = 32'hc4050d7;
      20606: inst = 32'h8220000;
      20607: inst = 32'h10408000;
      20608: inst = 32'hc4050d8;
      20609: inst = 32'h8220000;
      20610: inst = 32'h10408000;
      20611: inst = 32'hc4050d9;
      20612: inst = 32'h8220000;
      20613: inst = 32'h10408000;
      20614: inst = 32'hc4050da;
      20615: inst = 32'h8220000;
      20616: inst = 32'h10408000;
      20617: inst = 32'hc4050db;
      20618: inst = 32'h8220000;
      20619: inst = 32'h10408000;
      20620: inst = 32'hc4050dc;
      20621: inst = 32'h8220000;
      20622: inst = 32'h10408000;
      20623: inst = 32'hc4050dd;
      20624: inst = 32'h8220000;
      20625: inst = 32'h10408000;
      20626: inst = 32'hc4050de;
      20627: inst = 32'h8220000;
      20628: inst = 32'h10408000;
      20629: inst = 32'hc4050df;
      20630: inst = 32'h8220000;
      20631: inst = 32'h10408000;
      20632: inst = 32'hc4050e0;
      20633: inst = 32'h8220000;
      20634: inst = 32'h10408000;
      20635: inst = 32'hc4050e1;
      20636: inst = 32'h8220000;
      20637: inst = 32'h10408000;
      20638: inst = 32'hc4050e5;
      20639: inst = 32'h8220000;
      20640: inst = 32'h10408000;
      20641: inst = 32'hc4050e6;
      20642: inst = 32'h8220000;
      20643: inst = 32'h10408000;
      20644: inst = 32'hc4050e7;
      20645: inst = 32'h8220000;
      20646: inst = 32'h10408000;
      20647: inst = 32'hc4050e8;
      20648: inst = 32'h8220000;
      20649: inst = 32'h10408000;
      20650: inst = 32'hc4050e9;
      20651: inst = 32'h8220000;
      20652: inst = 32'h10408000;
      20653: inst = 32'hc4050ea;
      20654: inst = 32'h8220000;
      20655: inst = 32'h10408000;
      20656: inst = 32'hc4050eb;
      20657: inst = 32'h8220000;
      20658: inst = 32'h10408000;
      20659: inst = 32'hc4050ec;
      20660: inst = 32'h8220000;
      20661: inst = 32'h10408000;
      20662: inst = 32'hc4050ed;
      20663: inst = 32'h8220000;
      20664: inst = 32'h10408000;
      20665: inst = 32'hc4050f0;
      20666: inst = 32'h8220000;
      20667: inst = 32'h10408000;
      20668: inst = 32'hc4050f1;
      20669: inst = 32'h8220000;
      20670: inst = 32'h10408000;
      20671: inst = 32'hc4050f6;
      20672: inst = 32'h8220000;
      20673: inst = 32'h10408000;
      20674: inst = 32'hc4050f7;
      20675: inst = 32'h8220000;
      20676: inst = 32'h10408000;
      20677: inst = 32'hc4050f8;
      20678: inst = 32'h8220000;
      20679: inst = 32'h10408000;
      20680: inst = 32'hc4050f9;
      20681: inst = 32'h8220000;
      20682: inst = 32'h10408000;
      20683: inst = 32'hc4050fa;
      20684: inst = 32'h8220000;
      20685: inst = 32'h10408000;
      20686: inst = 32'hc4050fc;
      20687: inst = 32'h8220000;
      20688: inst = 32'h10408000;
      20689: inst = 32'hc4050fd;
      20690: inst = 32'h8220000;
      20691: inst = 32'h10408000;
      20692: inst = 32'hc405109;
      20693: inst = 32'h8220000;
      20694: inst = 32'h10408000;
      20695: inst = 32'hc40510a;
      20696: inst = 32'h8220000;
      20697: inst = 32'h10408000;
      20698: inst = 32'hc40510b;
      20699: inst = 32'h8220000;
      20700: inst = 32'h10408000;
      20701: inst = 32'hc40510c;
      20702: inst = 32'h8220000;
      20703: inst = 32'h10408000;
      20704: inst = 32'hc40510d;
      20705: inst = 32'h8220000;
      20706: inst = 32'h10408000;
      20707: inst = 32'hc40510e;
      20708: inst = 32'h8220000;
      20709: inst = 32'h10408000;
      20710: inst = 32'hc40510f;
      20711: inst = 32'h8220000;
      20712: inst = 32'h10408000;
      20713: inst = 32'hc405110;
      20714: inst = 32'h8220000;
      20715: inst = 32'h10408000;
      20716: inst = 32'hc405111;
      20717: inst = 32'h8220000;
      20718: inst = 32'h10408000;
      20719: inst = 32'hc405112;
      20720: inst = 32'h8220000;
      20721: inst = 32'h10408000;
      20722: inst = 32'hc405113;
      20723: inst = 32'h8220000;
      20724: inst = 32'h58000000;
      20725: inst = 32'hc20529c;
      20726: inst = 32'h10408000;
      20727: inst = 32'hc404224;
      20728: inst = 32'h8220000;
      20729: inst = 32'h10408000;
      20730: inst = 32'hc404225;
      20731: inst = 32'h8220000;
      20732: inst = 32'h10408000;
      20733: inst = 32'hc404226;
      20734: inst = 32'h8220000;
      20735: inst = 32'h10408000;
      20736: inst = 32'hc404227;
      20737: inst = 32'h8220000;
      20738: inst = 32'h10408000;
      20739: inst = 32'hc404228;
      20740: inst = 32'h8220000;
      20741: inst = 32'h10408000;
      20742: inst = 32'hc404229;
      20743: inst = 32'h8220000;
      20744: inst = 32'h10408000;
      20745: inst = 32'hc40422a;
      20746: inst = 32'h8220000;
      20747: inst = 32'h10408000;
      20748: inst = 32'hc40422b;
      20749: inst = 32'h8220000;
      20750: inst = 32'h10408000;
      20751: inst = 32'hc40422c;
      20752: inst = 32'h8220000;
      20753: inst = 32'h10408000;
      20754: inst = 32'hc40422d;
      20755: inst = 32'h8220000;
      20756: inst = 32'h10408000;
      20757: inst = 32'hc40422e;
      20758: inst = 32'h8220000;
      20759: inst = 32'h10408000;
      20760: inst = 32'hc40422f;
      20761: inst = 32'h8220000;
      20762: inst = 32'h10408000;
      20763: inst = 32'hc404230;
      20764: inst = 32'h8220000;
      20765: inst = 32'h10408000;
      20766: inst = 32'hc404231;
      20767: inst = 32'h8220000;
      20768: inst = 32'h10408000;
      20769: inst = 32'hc404232;
      20770: inst = 32'h8220000;
      20771: inst = 32'h10408000;
      20772: inst = 32'hc404233;
      20773: inst = 32'h8220000;
      20774: inst = 32'h10408000;
      20775: inst = 32'hc404234;
      20776: inst = 32'h8220000;
      20777: inst = 32'h10408000;
      20778: inst = 32'hc404235;
      20779: inst = 32'h8220000;
      20780: inst = 32'h10408000;
      20781: inst = 32'hc404236;
      20782: inst = 32'h8220000;
      20783: inst = 32'h10408000;
      20784: inst = 32'hc404237;
      20785: inst = 32'h8220000;
      20786: inst = 32'h10408000;
      20787: inst = 32'hc404238;
      20788: inst = 32'h8220000;
      20789: inst = 32'h10408000;
      20790: inst = 32'hc404239;
      20791: inst = 32'h8220000;
      20792: inst = 32'h10408000;
      20793: inst = 32'hc40423a;
      20794: inst = 32'h8220000;
      20795: inst = 32'h10408000;
      20796: inst = 32'hc40423b;
      20797: inst = 32'h8220000;
      20798: inst = 32'h10408000;
      20799: inst = 32'hc40423c;
      20800: inst = 32'h8220000;
      20801: inst = 32'h10408000;
      20802: inst = 32'hc40423d;
      20803: inst = 32'h8220000;
      20804: inst = 32'h10408000;
      20805: inst = 32'hc40423e;
      20806: inst = 32'h8220000;
      20807: inst = 32'h10408000;
      20808: inst = 32'hc40423f;
      20809: inst = 32'h8220000;
      20810: inst = 32'h10408000;
      20811: inst = 32'hc404240;
      20812: inst = 32'h8220000;
      20813: inst = 32'h10408000;
      20814: inst = 32'hc404241;
      20815: inst = 32'h8220000;
      20816: inst = 32'h10408000;
      20817: inst = 32'hc404242;
      20818: inst = 32'h8220000;
      20819: inst = 32'h10408000;
      20820: inst = 32'hc404243;
      20821: inst = 32'h8220000;
      20822: inst = 32'h10408000;
      20823: inst = 32'hc404244;
      20824: inst = 32'h8220000;
      20825: inst = 32'h10408000;
      20826: inst = 32'hc404245;
      20827: inst = 32'h8220000;
      20828: inst = 32'h10408000;
      20829: inst = 32'hc404246;
      20830: inst = 32'h8220000;
      20831: inst = 32'h10408000;
      20832: inst = 32'hc404247;
      20833: inst = 32'h8220000;
      20834: inst = 32'h10408000;
      20835: inst = 32'hc404248;
      20836: inst = 32'h8220000;
      20837: inst = 32'h10408000;
      20838: inst = 32'hc404249;
      20839: inst = 32'h8220000;
      20840: inst = 32'h10408000;
      20841: inst = 32'hc40424a;
      20842: inst = 32'h8220000;
      20843: inst = 32'h10408000;
      20844: inst = 32'hc40424b;
      20845: inst = 32'h8220000;
      20846: inst = 32'h10408000;
      20847: inst = 32'hc40424c;
      20848: inst = 32'h8220000;
      20849: inst = 32'h10408000;
      20850: inst = 32'hc40424d;
      20851: inst = 32'h8220000;
      20852: inst = 32'h10408000;
      20853: inst = 32'hc40424e;
      20854: inst = 32'h8220000;
      20855: inst = 32'h10408000;
      20856: inst = 32'hc40424f;
      20857: inst = 32'h8220000;
      20858: inst = 32'h10408000;
      20859: inst = 32'hc404250;
      20860: inst = 32'h8220000;
      20861: inst = 32'h10408000;
      20862: inst = 32'hc404251;
      20863: inst = 32'h8220000;
      20864: inst = 32'h10408000;
      20865: inst = 32'hc404252;
      20866: inst = 32'h8220000;
      20867: inst = 32'h10408000;
      20868: inst = 32'hc404253;
      20869: inst = 32'h8220000;
      20870: inst = 32'h10408000;
      20871: inst = 32'hc404254;
      20872: inst = 32'h8220000;
      20873: inst = 32'h10408000;
      20874: inst = 32'hc404255;
      20875: inst = 32'h8220000;
      20876: inst = 32'h10408000;
      20877: inst = 32'hc404256;
      20878: inst = 32'h8220000;
      20879: inst = 32'h10408000;
      20880: inst = 32'hc404257;
      20881: inst = 32'h8220000;
      20882: inst = 32'h10408000;
      20883: inst = 32'hc404258;
      20884: inst = 32'h8220000;
      20885: inst = 32'h10408000;
      20886: inst = 32'hc404259;
      20887: inst = 32'h8220000;
      20888: inst = 32'h10408000;
      20889: inst = 32'hc40425a;
      20890: inst = 32'h8220000;
      20891: inst = 32'h10408000;
      20892: inst = 32'hc40425b;
      20893: inst = 32'h8220000;
      20894: inst = 32'h10408000;
      20895: inst = 32'hc40425c;
      20896: inst = 32'h8220000;
      20897: inst = 32'h10408000;
      20898: inst = 32'hc40425d;
      20899: inst = 32'h8220000;
      20900: inst = 32'h10408000;
      20901: inst = 32'hc40425e;
      20902: inst = 32'h8220000;
      20903: inst = 32'h10408000;
      20904: inst = 32'hc40425f;
      20905: inst = 32'h8220000;
      20906: inst = 32'h10408000;
      20907: inst = 32'hc404260;
      20908: inst = 32'h8220000;
      20909: inst = 32'h10408000;
      20910: inst = 32'hc404261;
      20911: inst = 32'h8220000;
      20912: inst = 32'h10408000;
      20913: inst = 32'hc404262;
      20914: inst = 32'h8220000;
      20915: inst = 32'h10408000;
      20916: inst = 32'hc404263;
      20917: inst = 32'h8220000;
      20918: inst = 32'h10408000;
      20919: inst = 32'hc404264;
      20920: inst = 32'h8220000;
      20921: inst = 32'h10408000;
      20922: inst = 32'hc404265;
      20923: inst = 32'h8220000;
      20924: inst = 32'h10408000;
      20925: inst = 32'hc404266;
      20926: inst = 32'h8220000;
      20927: inst = 32'h10408000;
      20928: inst = 32'hc404267;
      20929: inst = 32'h8220000;
      20930: inst = 32'h10408000;
      20931: inst = 32'hc404268;
      20932: inst = 32'h8220000;
      20933: inst = 32'h10408000;
      20934: inst = 32'hc404269;
      20935: inst = 32'h8220000;
      20936: inst = 32'h10408000;
      20937: inst = 32'hc40426a;
      20938: inst = 32'h8220000;
      20939: inst = 32'h10408000;
      20940: inst = 32'hc40426b;
      20941: inst = 32'h8220000;
      20942: inst = 32'h10408000;
      20943: inst = 32'hc40426c;
      20944: inst = 32'h8220000;
      20945: inst = 32'h10408000;
      20946: inst = 32'hc40426d;
      20947: inst = 32'h8220000;
      20948: inst = 32'h10408000;
      20949: inst = 32'hc40426e;
      20950: inst = 32'h8220000;
      20951: inst = 32'h10408000;
      20952: inst = 32'hc40426f;
      20953: inst = 32'h8220000;
      20954: inst = 32'h10408000;
      20955: inst = 32'hc404270;
      20956: inst = 32'h8220000;
      20957: inst = 32'h10408000;
      20958: inst = 32'hc404271;
      20959: inst = 32'h8220000;
      20960: inst = 32'h10408000;
      20961: inst = 32'hc404272;
      20962: inst = 32'h8220000;
      20963: inst = 32'h10408000;
      20964: inst = 32'hc404273;
      20965: inst = 32'h8220000;
      20966: inst = 32'h10408000;
      20967: inst = 32'hc404274;
      20968: inst = 32'h8220000;
      20969: inst = 32'h10408000;
      20970: inst = 32'hc404275;
      20971: inst = 32'h8220000;
      20972: inst = 32'h10408000;
      20973: inst = 32'hc404276;
      20974: inst = 32'h8220000;
      20975: inst = 32'h10408000;
      20976: inst = 32'hc404277;
      20977: inst = 32'h8220000;
      20978: inst = 32'h10408000;
      20979: inst = 32'hc404278;
      20980: inst = 32'h8220000;
      20981: inst = 32'h10408000;
      20982: inst = 32'hc404279;
      20983: inst = 32'h8220000;
      20984: inst = 32'h10408000;
      20985: inst = 32'hc40427a;
      20986: inst = 32'h8220000;
      20987: inst = 32'h10408000;
      20988: inst = 32'hc40427b;
      20989: inst = 32'h8220000;
      20990: inst = 32'h10408000;
      20991: inst = 32'hc404284;
      20992: inst = 32'h8220000;
      20993: inst = 32'h10408000;
      20994: inst = 32'hc404285;
      20995: inst = 32'h8220000;
      20996: inst = 32'h10408000;
      20997: inst = 32'hc404286;
      20998: inst = 32'h8220000;
      20999: inst = 32'h10408000;
      21000: inst = 32'hc404287;
      21001: inst = 32'h8220000;
      21002: inst = 32'h10408000;
      21003: inst = 32'hc404288;
      21004: inst = 32'h8220000;
      21005: inst = 32'h10408000;
      21006: inst = 32'hc404289;
      21007: inst = 32'h8220000;
      21008: inst = 32'h10408000;
      21009: inst = 32'hc40428a;
      21010: inst = 32'h8220000;
      21011: inst = 32'h10408000;
      21012: inst = 32'hc40428b;
      21013: inst = 32'h8220000;
      21014: inst = 32'h10408000;
      21015: inst = 32'hc40428c;
      21016: inst = 32'h8220000;
      21017: inst = 32'h10408000;
      21018: inst = 32'hc40428d;
      21019: inst = 32'h8220000;
      21020: inst = 32'h10408000;
      21021: inst = 32'hc40428e;
      21022: inst = 32'h8220000;
      21023: inst = 32'h10408000;
      21024: inst = 32'hc40428f;
      21025: inst = 32'h8220000;
      21026: inst = 32'h10408000;
      21027: inst = 32'hc404290;
      21028: inst = 32'h8220000;
      21029: inst = 32'h10408000;
      21030: inst = 32'hc404291;
      21031: inst = 32'h8220000;
      21032: inst = 32'h10408000;
      21033: inst = 32'hc404292;
      21034: inst = 32'h8220000;
      21035: inst = 32'h10408000;
      21036: inst = 32'hc404293;
      21037: inst = 32'h8220000;
      21038: inst = 32'h10408000;
      21039: inst = 32'hc404294;
      21040: inst = 32'h8220000;
      21041: inst = 32'h10408000;
      21042: inst = 32'hc404295;
      21043: inst = 32'h8220000;
      21044: inst = 32'h10408000;
      21045: inst = 32'hc404296;
      21046: inst = 32'h8220000;
      21047: inst = 32'h10408000;
      21048: inst = 32'hc404297;
      21049: inst = 32'h8220000;
      21050: inst = 32'h10408000;
      21051: inst = 32'hc404298;
      21052: inst = 32'h8220000;
      21053: inst = 32'h10408000;
      21054: inst = 32'hc404299;
      21055: inst = 32'h8220000;
      21056: inst = 32'h10408000;
      21057: inst = 32'hc40429a;
      21058: inst = 32'h8220000;
      21059: inst = 32'h10408000;
      21060: inst = 32'hc40429b;
      21061: inst = 32'h8220000;
      21062: inst = 32'h10408000;
      21063: inst = 32'hc40429c;
      21064: inst = 32'h8220000;
      21065: inst = 32'h10408000;
      21066: inst = 32'hc40429d;
      21067: inst = 32'h8220000;
      21068: inst = 32'h10408000;
      21069: inst = 32'hc40429e;
      21070: inst = 32'h8220000;
      21071: inst = 32'h10408000;
      21072: inst = 32'hc40429f;
      21073: inst = 32'h8220000;
      21074: inst = 32'h10408000;
      21075: inst = 32'hc4042a0;
      21076: inst = 32'h8220000;
      21077: inst = 32'h10408000;
      21078: inst = 32'hc4042a1;
      21079: inst = 32'h8220000;
      21080: inst = 32'h10408000;
      21081: inst = 32'hc4042a2;
      21082: inst = 32'h8220000;
      21083: inst = 32'h10408000;
      21084: inst = 32'hc4042a3;
      21085: inst = 32'h8220000;
      21086: inst = 32'h10408000;
      21087: inst = 32'hc4042a4;
      21088: inst = 32'h8220000;
      21089: inst = 32'h10408000;
      21090: inst = 32'hc4042a5;
      21091: inst = 32'h8220000;
      21092: inst = 32'h10408000;
      21093: inst = 32'hc4042a6;
      21094: inst = 32'h8220000;
      21095: inst = 32'h10408000;
      21096: inst = 32'hc4042a7;
      21097: inst = 32'h8220000;
      21098: inst = 32'h10408000;
      21099: inst = 32'hc4042a8;
      21100: inst = 32'h8220000;
      21101: inst = 32'h10408000;
      21102: inst = 32'hc4042a9;
      21103: inst = 32'h8220000;
      21104: inst = 32'h10408000;
      21105: inst = 32'hc4042aa;
      21106: inst = 32'h8220000;
      21107: inst = 32'h10408000;
      21108: inst = 32'hc4042ab;
      21109: inst = 32'h8220000;
      21110: inst = 32'h10408000;
      21111: inst = 32'hc4042ac;
      21112: inst = 32'h8220000;
      21113: inst = 32'h10408000;
      21114: inst = 32'hc4042ad;
      21115: inst = 32'h8220000;
      21116: inst = 32'h10408000;
      21117: inst = 32'hc4042ae;
      21118: inst = 32'h8220000;
      21119: inst = 32'h10408000;
      21120: inst = 32'hc4042af;
      21121: inst = 32'h8220000;
      21122: inst = 32'h10408000;
      21123: inst = 32'hc4042b0;
      21124: inst = 32'h8220000;
      21125: inst = 32'h10408000;
      21126: inst = 32'hc4042b1;
      21127: inst = 32'h8220000;
      21128: inst = 32'h10408000;
      21129: inst = 32'hc4042b2;
      21130: inst = 32'h8220000;
      21131: inst = 32'h10408000;
      21132: inst = 32'hc4042b3;
      21133: inst = 32'h8220000;
      21134: inst = 32'h10408000;
      21135: inst = 32'hc4042b4;
      21136: inst = 32'h8220000;
      21137: inst = 32'h10408000;
      21138: inst = 32'hc4042b5;
      21139: inst = 32'h8220000;
      21140: inst = 32'h10408000;
      21141: inst = 32'hc4042b6;
      21142: inst = 32'h8220000;
      21143: inst = 32'h10408000;
      21144: inst = 32'hc4042b7;
      21145: inst = 32'h8220000;
      21146: inst = 32'h10408000;
      21147: inst = 32'hc4042b8;
      21148: inst = 32'h8220000;
      21149: inst = 32'h10408000;
      21150: inst = 32'hc4042b9;
      21151: inst = 32'h8220000;
      21152: inst = 32'h10408000;
      21153: inst = 32'hc4042ba;
      21154: inst = 32'h8220000;
      21155: inst = 32'h10408000;
      21156: inst = 32'hc4042bb;
      21157: inst = 32'h8220000;
      21158: inst = 32'h10408000;
      21159: inst = 32'hc4042bc;
      21160: inst = 32'h8220000;
      21161: inst = 32'h10408000;
      21162: inst = 32'hc4042bd;
      21163: inst = 32'h8220000;
      21164: inst = 32'h10408000;
      21165: inst = 32'hc4042be;
      21166: inst = 32'h8220000;
      21167: inst = 32'h10408000;
      21168: inst = 32'hc4042bf;
      21169: inst = 32'h8220000;
      21170: inst = 32'h10408000;
      21171: inst = 32'hc4042c0;
      21172: inst = 32'h8220000;
      21173: inst = 32'h10408000;
      21174: inst = 32'hc4042c1;
      21175: inst = 32'h8220000;
      21176: inst = 32'h10408000;
      21177: inst = 32'hc4042c2;
      21178: inst = 32'h8220000;
      21179: inst = 32'h10408000;
      21180: inst = 32'hc4042c3;
      21181: inst = 32'h8220000;
      21182: inst = 32'h10408000;
      21183: inst = 32'hc4042c4;
      21184: inst = 32'h8220000;
      21185: inst = 32'h10408000;
      21186: inst = 32'hc4042c5;
      21187: inst = 32'h8220000;
      21188: inst = 32'h10408000;
      21189: inst = 32'hc4042c6;
      21190: inst = 32'h8220000;
      21191: inst = 32'h10408000;
      21192: inst = 32'hc4042c7;
      21193: inst = 32'h8220000;
      21194: inst = 32'h10408000;
      21195: inst = 32'hc4042c8;
      21196: inst = 32'h8220000;
      21197: inst = 32'h10408000;
      21198: inst = 32'hc4042c9;
      21199: inst = 32'h8220000;
      21200: inst = 32'h10408000;
      21201: inst = 32'hc4042ca;
      21202: inst = 32'h8220000;
      21203: inst = 32'h10408000;
      21204: inst = 32'hc4042cb;
      21205: inst = 32'h8220000;
      21206: inst = 32'h10408000;
      21207: inst = 32'hc4042cc;
      21208: inst = 32'h8220000;
      21209: inst = 32'h10408000;
      21210: inst = 32'hc4042cd;
      21211: inst = 32'h8220000;
      21212: inst = 32'h10408000;
      21213: inst = 32'hc4042ce;
      21214: inst = 32'h8220000;
      21215: inst = 32'h10408000;
      21216: inst = 32'hc4042cf;
      21217: inst = 32'h8220000;
      21218: inst = 32'h10408000;
      21219: inst = 32'hc4042d0;
      21220: inst = 32'h8220000;
      21221: inst = 32'h10408000;
      21222: inst = 32'hc4042d1;
      21223: inst = 32'h8220000;
      21224: inst = 32'h10408000;
      21225: inst = 32'hc4042d2;
      21226: inst = 32'h8220000;
      21227: inst = 32'h10408000;
      21228: inst = 32'hc4042d3;
      21229: inst = 32'h8220000;
      21230: inst = 32'h10408000;
      21231: inst = 32'hc4042d4;
      21232: inst = 32'h8220000;
      21233: inst = 32'h10408000;
      21234: inst = 32'hc4042d5;
      21235: inst = 32'h8220000;
      21236: inst = 32'h10408000;
      21237: inst = 32'hc4042d6;
      21238: inst = 32'h8220000;
      21239: inst = 32'h10408000;
      21240: inst = 32'hc4042d7;
      21241: inst = 32'h8220000;
      21242: inst = 32'h10408000;
      21243: inst = 32'hc4042d8;
      21244: inst = 32'h8220000;
      21245: inst = 32'h10408000;
      21246: inst = 32'hc4042d9;
      21247: inst = 32'h8220000;
      21248: inst = 32'h10408000;
      21249: inst = 32'hc4042da;
      21250: inst = 32'h8220000;
      21251: inst = 32'h10408000;
      21252: inst = 32'hc4042db;
      21253: inst = 32'h8220000;
      21254: inst = 32'h10408000;
      21255: inst = 32'hc4042e4;
      21256: inst = 32'h8220000;
      21257: inst = 32'h10408000;
      21258: inst = 32'hc4042e5;
      21259: inst = 32'h8220000;
      21260: inst = 32'h10408000;
      21261: inst = 32'hc4042e6;
      21262: inst = 32'h8220000;
      21263: inst = 32'h10408000;
      21264: inst = 32'hc404339;
      21265: inst = 32'h8220000;
      21266: inst = 32'h10408000;
      21267: inst = 32'hc40433a;
      21268: inst = 32'h8220000;
      21269: inst = 32'h10408000;
      21270: inst = 32'hc40433b;
      21271: inst = 32'h8220000;
      21272: inst = 32'h10408000;
      21273: inst = 32'hc404344;
      21274: inst = 32'h8220000;
      21275: inst = 32'h10408000;
      21276: inst = 32'hc404345;
      21277: inst = 32'h8220000;
      21278: inst = 32'h10408000;
      21279: inst = 32'hc40439a;
      21280: inst = 32'h8220000;
      21281: inst = 32'h10408000;
      21282: inst = 32'hc40439b;
      21283: inst = 32'h8220000;
      21284: inst = 32'h10408000;
      21285: inst = 32'hc4043a4;
      21286: inst = 32'h8220000;
      21287: inst = 32'h10408000;
      21288: inst = 32'hc4043a5;
      21289: inst = 32'h8220000;
      21290: inst = 32'h10408000;
      21291: inst = 32'hc4043fa;
      21292: inst = 32'h8220000;
      21293: inst = 32'h10408000;
      21294: inst = 32'hc4043fb;
      21295: inst = 32'h8220000;
      21296: inst = 32'h10408000;
      21297: inst = 32'hc404404;
      21298: inst = 32'h8220000;
      21299: inst = 32'h10408000;
      21300: inst = 32'hc404405;
      21301: inst = 32'h8220000;
      21302: inst = 32'h10408000;
      21303: inst = 32'hc40445a;
      21304: inst = 32'h8220000;
      21305: inst = 32'h10408000;
      21306: inst = 32'hc40445b;
      21307: inst = 32'h8220000;
      21308: inst = 32'h10408000;
      21309: inst = 32'hc404464;
      21310: inst = 32'h8220000;
      21311: inst = 32'h10408000;
      21312: inst = 32'hc404465;
      21313: inst = 32'h8220000;
      21314: inst = 32'h10408000;
      21315: inst = 32'hc4044ba;
      21316: inst = 32'h8220000;
      21317: inst = 32'h10408000;
      21318: inst = 32'hc4044bb;
      21319: inst = 32'h8220000;
      21320: inst = 32'h10408000;
      21321: inst = 32'hc4044c4;
      21322: inst = 32'h8220000;
      21323: inst = 32'h10408000;
      21324: inst = 32'hc4044c5;
      21325: inst = 32'h8220000;
      21326: inst = 32'h10408000;
      21327: inst = 32'hc40451a;
      21328: inst = 32'h8220000;
      21329: inst = 32'h10408000;
      21330: inst = 32'hc40451b;
      21331: inst = 32'h8220000;
      21332: inst = 32'h10408000;
      21333: inst = 32'hc404524;
      21334: inst = 32'h8220000;
      21335: inst = 32'h10408000;
      21336: inst = 32'hc404525;
      21337: inst = 32'h8220000;
      21338: inst = 32'h10408000;
      21339: inst = 32'hc40457a;
      21340: inst = 32'h8220000;
      21341: inst = 32'h10408000;
      21342: inst = 32'hc40457b;
      21343: inst = 32'h8220000;
      21344: inst = 32'h10408000;
      21345: inst = 32'hc404584;
      21346: inst = 32'h8220000;
      21347: inst = 32'h10408000;
      21348: inst = 32'hc404585;
      21349: inst = 32'h8220000;
      21350: inst = 32'h10408000;
      21351: inst = 32'hc4045da;
      21352: inst = 32'h8220000;
      21353: inst = 32'h10408000;
      21354: inst = 32'hc4045db;
      21355: inst = 32'h8220000;
      21356: inst = 32'h10408000;
      21357: inst = 32'hc4045e4;
      21358: inst = 32'h8220000;
      21359: inst = 32'h10408000;
      21360: inst = 32'hc4045e5;
      21361: inst = 32'h8220000;
      21362: inst = 32'h10408000;
      21363: inst = 32'hc40463a;
      21364: inst = 32'h8220000;
      21365: inst = 32'h10408000;
      21366: inst = 32'hc40463b;
      21367: inst = 32'h8220000;
      21368: inst = 32'h10408000;
      21369: inst = 32'hc404644;
      21370: inst = 32'h8220000;
      21371: inst = 32'h10408000;
      21372: inst = 32'hc404645;
      21373: inst = 32'h8220000;
      21374: inst = 32'h10408000;
      21375: inst = 32'hc40469a;
      21376: inst = 32'h8220000;
      21377: inst = 32'h10408000;
      21378: inst = 32'hc40469b;
      21379: inst = 32'h8220000;
      21380: inst = 32'h10408000;
      21381: inst = 32'hc4046a4;
      21382: inst = 32'h8220000;
      21383: inst = 32'h10408000;
      21384: inst = 32'hc4046a5;
      21385: inst = 32'h8220000;
      21386: inst = 32'h10408000;
      21387: inst = 32'hc4046fa;
      21388: inst = 32'h8220000;
      21389: inst = 32'h10408000;
      21390: inst = 32'hc4046fb;
      21391: inst = 32'h8220000;
      21392: inst = 32'h10408000;
      21393: inst = 32'hc404704;
      21394: inst = 32'h8220000;
      21395: inst = 32'h10408000;
      21396: inst = 32'hc404705;
      21397: inst = 32'h8220000;
      21398: inst = 32'h10408000;
      21399: inst = 32'hc40475a;
      21400: inst = 32'h8220000;
      21401: inst = 32'h10408000;
      21402: inst = 32'hc40475b;
      21403: inst = 32'h8220000;
      21404: inst = 32'h10408000;
      21405: inst = 32'hc404764;
      21406: inst = 32'h8220000;
      21407: inst = 32'h10408000;
      21408: inst = 32'hc404765;
      21409: inst = 32'h8220000;
      21410: inst = 32'h10408000;
      21411: inst = 32'hc4047ba;
      21412: inst = 32'h8220000;
      21413: inst = 32'h10408000;
      21414: inst = 32'hc4047bb;
      21415: inst = 32'h8220000;
      21416: inst = 32'h10408000;
      21417: inst = 32'hc4047c4;
      21418: inst = 32'h8220000;
      21419: inst = 32'h10408000;
      21420: inst = 32'hc4047c5;
      21421: inst = 32'h8220000;
      21422: inst = 32'h10408000;
      21423: inst = 32'hc40481a;
      21424: inst = 32'h8220000;
      21425: inst = 32'h10408000;
      21426: inst = 32'hc40481b;
      21427: inst = 32'h8220000;
      21428: inst = 32'h10408000;
      21429: inst = 32'hc404824;
      21430: inst = 32'h8220000;
      21431: inst = 32'h10408000;
      21432: inst = 32'hc404825;
      21433: inst = 32'h8220000;
      21434: inst = 32'h10408000;
      21435: inst = 32'hc40487a;
      21436: inst = 32'h8220000;
      21437: inst = 32'h10408000;
      21438: inst = 32'hc40487b;
      21439: inst = 32'h8220000;
      21440: inst = 32'h10408000;
      21441: inst = 32'hc404884;
      21442: inst = 32'h8220000;
      21443: inst = 32'h10408000;
      21444: inst = 32'hc404885;
      21445: inst = 32'h8220000;
      21446: inst = 32'h10408000;
      21447: inst = 32'hc4048da;
      21448: inst = 32'h8220000;
      21449: inst = 32'h10408000;
      21450: inst = 32'hc4048db;
      21451: inst = 32'h8220000;
      21452: inst = 32'h10408000;
      21453: inst = 32'hc4048e4;
      21454: inst = 32'h8220000;
      21455: inst = 32'h10408000;
      21456: inst = 32'hc4048e5;
      21457: inst = 32'h8220000;
      21458: inst = 32'h10408000;
      21459: inst = 32'hc40493a;
      21460: inst = 32'h8220000;
      21461: inst = 32'h10408000;
      21462: inst = 32'hc40493b;
      21463: inst = 32'h8220000;
      21464: inst = 32'h10408000;
      21465: inst = 32'hc404944;
      21466: inst = 32'h8220000;
      21467: inst = 32'h10408000;
      21468: inst = 32'hc404945;
      21469: inst = 32'h8220000;
      21470: inst = 32'h10408000;
      21471: inst = 32'hc40499a;
      21472: inst = 32'h8220000;
      21473: inst = 32'h10408000;
      21474: inst = 32'hc40499b;
      21475: inst = 32'h8220000;
      21476: inst = 32'h10408000;
      21477: inst = 32'hc4049a4;
      21478: inst = 32'h8220000;
      21479: inst = 32'h10408000;
      21480: inst = 32'hc4049a5;
      21481: inst = 32'h8220000;
      21482: inst = 32'h10408000;
      21483: inst = 32'hc4049fa;
      21484: inst = 32'h8220000;
      21485: inst = 32'h10408000;
      21486: inst = 32'hc4049fb;
      21487: inst = 32'h8220000;
      21488: inst = 32'h10408000;
      21489: inst = 32'hc404a04;
      21490: inst = 32'h8220000;
      21491: inst = 32'h10408000;
      21492: inst = 32'hc404a05;
      21493: inst = 32'h8220000;
      21494: inst = 32'h10408000;
      21495: inst = 32'hc404a5a;
      21496: inst = 32'h8220000;
      21497: inst = 32'h10408000;
      21498: inst = 32'hc404a5b;
      21499: inst = 32'h8220000;
      21500: inst = 32'h10408000;
      21501: inst = 32'hc404a64;
      21502: inst = 32'h8220000;
      21503: inst = 32'h10408000;
      21504: inst = 32'hc404a65;
      21505: inst = 32'h8220000;
      21506: inst = 32'h10408000;
      21507: inst = 32'hc404aba;
      21508: inst = 32'h8220000;
      21509: inst = 32'h10408000;
      21510: inst = 32'hc404abb;
      21511: inst = 32'h8220000;
      21512: inst = 32'h10408000;
      21513: inst = 32'hc404ac4;
      21514: inst = 32'h8220000;
      21515: inst = 32'h10408000;
      21516: inst = 32'hc404ac5;
      21517: inst = 32'h8220000;
      21518: inst = 32'h10408000;
      21519: inst = 32'hc404b1a;
      21520: inst = 32'h8220000;
      21521: inst = 32'h10408000;
      21522: inst = 32'hc404b1b;
      21523: inst = 32'h8220000;
      21524: inst = 32'h10408000;
      21525: inst = 32'hc404b24;
      21526: inst = 32'h8220000;
      21527: inst = 32'h10408000;
      21528: inst = 32'hc404b25;
      21529: inst = 32'h8220000;
      21530: inst = 32'h10408000;
      21531: inst = 32'hc404b7a;
      21532: inst = 32'h8220000;
      21533: inst = 32'h10408000;
      21534: inst = 32'hc404b7b;
      21535: inst = 32'h8220000;
      21536: inst = 32'h10408000;
      21537: inst = 32'hc404b84;
      21538: inst = 32'h8220000;
      21539: inst = 32'h10408000;
      21540: inst = 32'hc404b85;
      21541: inst = 32'h8220000;
      21542: inst = 32'h10408000;
      21543: inst = 32'hc404bda;
      21544: inst = 32'h8220000;
      21545: inst = 32'h10408000;
      21546: inst = 32'hc404bdb;
      21547: inst = 32'h8220000;
      21548: inst = 32'h10408000;
      21549: inst = 32'hc404be4;
      21550: inst = 32'h8220000;
      21551: inst = 32'h10408000;
      21552: inst = 32'hc404be5;
      21553: inst = 32'h8220000;
      21554: inst = 32'h10408000;
      21555: inst = 32'hc404c3a;
      21556: inst = 32'h8220000;
      21557: inst = 32'h10408000;
      21558: inst = 32'hc404c3b;
      21559: inst = 32'h8220000;
      21560: inst = 32'h10408000;
      21561: inst = 32'hc404c44;
      21562: inst = 32'h8220000;
      21563: inst = 32'h10408000;
      21564: inst = 32'hc404c45;
      21565: inst = 32'h8220000;
      21566: inst = 32'h10408000;
      21567: inst = 32'hc404c9a;
      21568: inst = 32'h8220000;
      21569: inst = 32'h10408000;
      21570: inst = 32'hc404c9b;
      21571: inst = 32'h8220000;
      21572: inst = 32'h10408000;
      21573: inst = 32'hc404ca4;
      21574: inst = 32'h8220000;
      21575: inst = 32'h10408000;
      21576: inst = 32'hc404ca5;
      21577: inst = 32'h8220000;
      21578: inst = 32'h10408000;
      21579: inst = 32'hc404cfa;
      21580: inst = 32'h8220000;
      21581: inst = 32'h10408000;
      21582: inst = 32'hc404cfb;
      21583: inst = 32'h8220000;
      21584: inst = 32'h10408000;
      21585: inst = 32'hc404d04;
      21586: inst = 32'h8220000;
      21587: inst = 32'h10408000;
      21588: inst = 32'hc404d05;
      21589: inst = 32'h8220000;
      21590: inst = 32'h10408000;
      21591: inst = 32'hc404d5a;
      21592: inst = 32'h8220000;
      21593: inst = 32'h10408000;
      21594: inst = 32'hc404d5b;
      21595: inst = 32'h8220000;
      21596: inst = 32'h10408000;
      21597: inst = 32'hc404d64;
      21598: inst = 32'h8220000;
      21599: inst = 32'h10408000;
      21600: inst = 32'hc404d65;
      21601: inst = 32'h8220000;
      21602: inst = 32'h10408000;
      21603: inst = 32'hc404dba;
      21604: inst = 32'h8220000;
      21605: inst = 32'h10408000;
      21606: inst = 32'hc404dbb;
      21607: inst = 32'h8220000;
      21608: inst = 32'h10408000;
      21609: inst = 32'hc404dc4;
      21610: inst = 32'h8220000;
      21611: inst = 32'h10408000;
      21612: inst = 32'hc404dc5;
      21613: inst = 32'h8220000;
      21614: inst = 32'h10408000;
      21615: inst = 32'hc404e1a;
      21616: inst = 32'h8220000;
      21617: inst = 32'h10408000;
      21618: inst = 32'hc404e1b;
      21619: inst = 32'h8220000;
      21620: inst = 32'h10408000;
      21621: inst = 32'hc404e24;
      21622: inst = 32'h8220000;
      21623: inst = 32'h10408000;
      21624: inst = 32'hc404e25;
      21625: inst = 32'h8220000;
      21626: inst = 32'h10408000;
      21627: inst = 32'hc404e7a;
      21628: inst = 32'h8220000;
      21629: inst = 32'h10408000;
      21630: inst = 32'hc404e7b;
      21631: inst = 32'h8220000;
      21632: inst = 32'h10408000;
      21633: inst = 32'hc404e84;
      21634: inst = 32'h8220000;
      21635: inst = 32'h10408000;
      21636: inst = 32'hc404e85;
      21637: inst = 32'h8220000;
      21638: inst = 32'h10408000;
      21639: inst = 32'hc404eda;
      21640: inst = 32'h8220000;
      21641: inst = 32'h10408000;
      21642: inst = 32'hc404edb;
      21643: inst = 32'h8220000;
      21644: inst = 32'h10408000;
      21645: inst = 32'hc404ee4;
      21646: inst = 32'h8220000;
      21647: inst = 32'h10408000;
      21648: inst = 32'hc404ee5;
      21649: inst = 32'h8220000;
      21650: inst = 32'h10408000;
      21651: inst = 32'hc404f3a;
      21652: inst = 32'h8220000;
      21653: inst = 32'h10408000;
      21654: inst = 32'hc404f3b;
      21655: inst = 32'h8220000;
      21656: inst = 32'h10408000;
      21657: inst = 32'hc404f44;
      21658: inst = 32'h8220000;
      21659: inst = 32'h10408000;
      21660: inst = 32'hc404f45;
      21661: inst = 32'h8220000;
      21662: inst = 32'h10408000;
      21663: inst = 32'hc404f9a;
      21664: inst = 32'h8220000;
      21665: inst = 32'h10408000;
      21666: inst = 32'hc404f9b;
      21667: inst = 32'h8220000;
      21668: inst = 32'h10408000;
      21669: inst = 32'hc404fa4;
      21670: inst = 32'h8220000;
      21671: inst = 32'h10408000;
      21672: inst = 32'hc404fa5;
      21673: inst = 32'h8220000;
      21674: inst = 32'h10408000;
      21675: inst = 32'hc404ffa;
      21676: inst = 32'h8220000;
      21677: inst = 32'h10408000;
      21678: inst = 32'hc404ffb;
      21679: inst = 32'h8220000;
      21680: inst = 32'h10408000;
      21681: inst = 32'hc405004;
      21682: inst = 32'h8220000;
      21683: inst = 32'h10408000;
      21684: inst = 32'hc405005;
      21685: inst = 32'h8220000;
      21686: inst = 32'h10408000;
      21687: inst = 32'hc40505a;
      21688: inst = 32'h8220000;
      21689: inst = 32'h10408000;
      21690: inst = 32'hc40505b;
      21691: inst = 32'h8220000;
      21692: inst = 32'h10408000;
      21693: inst = 32'hc405064;
      21694: inst = 32'h8220000;
      21695: inst = 32'h10408000;
      21696: inst = 32'hc405065;
      21697: inst = 32'h8220000;
      21698: inst = 32'h10408000;
      21699: inst = 32'hc4050ba;
      21700: inst = 32'h8220000;
      21701: inst = 32'h10408000;
      21702: inst = 32'hc4050bb;
      21703: inst = 32'h8220000;
      21704: inst = 32'h10408000;
      21705: inst = 32'hc4050c4;
      21706: inst = 32'h8220000;
      21707: inst = 32'h10408000;
      21708: inst = 32'hc4050c5;
      21709: inst = 32'h8220000;
      21710: inst = 32'h10408000;
      21711: inst = 32'hc40511a;
      21712: inst = 32'h8220000;
      21713: inst = 32'h10408000;
      21714: inst = 32'hc40511b;
      21715: inst = 32'h8220000;
      21716: inst = 32'h10408000;
      21717: inst = 32'hc405124;
      21718: inst = 32'h8220000;
      21719: inst = 32'h10408000;
      21720: inst = 32'hc405125;
      21721: inst = 32'h8220000;
      21722: inst = 32'h10408000;
      21723: inst = 32'hc40517a;
      21724: inst = 32'h8220000;
      21725: inst = 32'h10408000;
      21726: inst = 32'hc40517b;
      21727: inst = 32'h8220000;
      21728: inst = 32'h10408000;
      21729: inst = 32'hc405184;
      21730: inst = 32'h8220000;
      21731: inst = 32'h10408000;
      21732: inst = 32'hc405185;
      21733: inst = 32'h8220000;
      21734: inst = 32'h10408000;
      21735: inst = 32'hc4051da;
      21736: inst = 32'h8220000;
      21737: inst = 32'h10408000;
      21738: inst = 32'hc4051db;
      21739: inst = 32'h8220000;
      21740: inst = 32'h10408000;
      21741: inst = 32'hc4051e4;
      21742: inst = 32'h8220000;
      21743: inst = 32'h10408000;
      21744: inst = 32'hc4051e5;
      21745: inst = 32'h8220000;
      21746: inst = 32'h10408000;
      21747: inst = 32'hc40523a;
      21748: inst = 32'h8220000;
      21749: inst = 32'h10408000;
      21750: inst = 32'hc40523b;
      21751: inst = 32'h8220000;
      21752: inst = 32'h10408000;
      21753: inst = 32'hc405244;
      21754: inst = 32'h8220000;
      21755: inst = 32'h10408000;
      21756: inst = 32'hc405245;
      21757: inst = 32'h8220000;
      21758: inst = 32'h10408000;
      21759: inst = 32'hc40529a;
      21760: inst = 32'h8220000;
      21761: inst = 32'h10408000;
      21762: inst = 32'hc40529b;
      21763: inst = 32'h8220000;
      21764: inst = 32'h10408000;
      21765: inst = 32'hc4052a4;
      21766: inst = 32'h8220000;
      21767: inst = 32'h10408000;
      21768: inst = 32'hc4052a5;
      21769: inst = 32'h8220000;
      21770: inst = 32'h10408000;
      21771: inst = 32'hc4052fa;
      21772: inst = 32'h8220000;
      21773: inst = 32'h10408000;
      21774: inst = 32'hc4052fb;
      21775: inst = 32'h8220000;
      21776: inst = 32'h10408000;
      21777: inst = 32'hc405304;
      21778: inst = 32'h8220000;
      21779: inst = 32'h10408000;
      21780: inst = 32'hc405305;
      21781: inst = 32'h8220000;
      21782: inst = 32'h10408000;
      21783: inst = 32'hc40535a;
      21784: inst = 32'h8220000;
      21785: inst = 32'h10408000;
      21786: inst = 32'hc40535b;
      21787: inst = 32'h8220000;
      21788: inst = 32'h10408000;
      21789: inst = 32'hc405364;
      21790: inst = 32'h8220000;
      21791: inst = 32'h10408000;
      21792: inst = 32'hc405365;
      21793: inst = 32'h8220000;
      21794: inst = 32'h10408000;
      21795: inst = 32'hc4053ba;
      21796: inst = 32'h8220000;
      21797: inst = 32'h10408000;
      21798: inst = 32'hc4053bb;
      21799: inst = 32'h8220000;
      21800: inst = 32'h10408000;
      21801: inst = 32'hc4053c4;
      21802: inst = 32'h8220000;
      21803: inst = 32'h10408000;
      21804: inst = 32'hc4053c5;
      21805: inst = 32'h8220000;
      21806: inst = 32'h10408000;
      21807: inst = 32'hc40541a;
      21808: inst = 32'h8220000;
      21809: inst = 32'h10408000;
      21810: inst = 32'hc40541b;
      21811: inst = 32'h8220000;
      21812: inst = 32'h10408000;
      21813: inst = 32'hc405424;
      21814: inst = 32'h8220000;
      21815: inst = 32'h10408000;
      21816: inst = 32'hc405425;
      21817: inst = 32'h8220000;
      21818: inst = 32'h10408000;
      21819: inst = 32'hc405426;
      21820: inst = 32'h8220000;
      21821: inst = 32'h10408000;
      21822: inst = 32'hc405479;
      21823: inst = 32'h8220000;
      21824: inst = 32'h10408000;
      21825: inst = 32'hc40547a;
      21826: inst = 32'h8220000;
      21827: inst = 32'h10408000;
      21828: inst = 32'hc40547b;
      21829: inst = 32'h8220000;
      21830: inst = 32'h10408000;
      21831: inst = 32'hc405484;
      21832: inst = 32'h8220000;
      21833: inst = 32'h10408000;
      21834: inst = 32'hc405485;
      21835: inst = 32'h8220000;
      21836: inst = 32'h10408000;
      21837: inst = 32'hc405486;
      21838: inst = 32'h8220000;
      21839: inst = 32'h10408000;
      21840: inst = 32'hc405487;
      21841: inst = 32'h8220000;
      21842: inst = 32'h10408000;
      21843: inst = 32'hc405488;
      21844: inst = 32'h8220000;
      21845: inst = 32'h10408000;
      21846: inst = 32'hc405489;
      21847: inst = 32'h8220000;
      21848: inst = 32'h10408000;
      21849: inst = 32'hc40548a;
      21850: inst = 32'h8220000;
      21851: inst = 32'h10408000;
      21852: inst = 32'hc40548b;
      21853: inst = 32'h8220000;
      21854: inst = 32'h10408000;
      21855: inst = 32'hc40548c;
      21856: inst = 32'h8220000;
      21857: inst = 32'h10408000;
      21858: inst = 32'hc40548d;
      21859: inst = 32'h8220000;
      21860: inst = 32'h10408000;
      21861: inst = 32'hc40548e;
      21862: inst = 32'h8220000;
      21863: inst = 32'h10408000;
      21864: inst = 32'hc40548f;
      21865: inst = 32'h8220000;
      21866: inst = 32'h10408000;
      21867: inst = 32'hc405490;
      21868: inst = 32'h8220000;
      21869: inst = 32'h10408000;
      21870: inst = 32'hc405491;
      21871: inst = 32'h8220000;
      21872: inst = 32'h10408000;
      21873: inst = 32'hc405492;
      21874: inst = 32'h8220000;
      21875: inst = 32'h10408000;
      21876: inst = 32'hc405493;
      21877: inst = 32'h8220000;
      21878: inst = 32'h10408000;
      21879: inst = 32'hc405494;
      21880: inst = 32'h8220000;
      21881: inst = 32'h10408000;
      21882: inst = 32'hc405495;
      21883: inst = 32'h8220000;
      21884: inst = 32'h10408000;
      21885: inst = 32'hc405496;
      21886: inst = 32'h8220000;
      21887: inst = 32'h10408000;
      21888: inst = 32'hc405497;
      21889: inst = 32'h8220000;
      21890: inst = 32'h10408000;
      21891: inst = 32'hc405498;
      21892: inst = 32'h8220000;
      21893: inst = 32'h10408000;
      21894: inst = 32'hc405499;
      21895: inst = 32'h8220000;
      21896: inst = 32'h10408000;
      21897: inst = 32'hc40549a;
      21898: inst = 32'h8220000;
      21899: inst = 32'h10408000;
      21900: inst = 32'hc40549b;
      21901: inst = 32'h8220000;
      21902: inst = 32'h10408000;
      21903: inst = 32'hc40549c;
      21904: inst = 32'h8220000;
      21905: inst = 32'h10408000;
      21906: inst = 32'hc40549d;
      21907: inst = 32'h8220000;
      21908: inst = 32'h10408000;
      21909: inst = 32'hc40549e;
      21910: inst = 32'h8220000;
      21911: inst = 32'h10408000;
      21912: inst = 32'hc40549f;
      21913: inst = 32'h8220000;
      21914: inst = 32'h10408000;
      21915: inst = 32'hc4054a0;
      21916: inst = 32'h8220000;
      21917: inst = 32'h10408000;
      21918: inst = 32'hc4054a1;
      21919: inst = 32'h8220000;
      21920: inst = 32'h10408000;
      21921: inst = 32'hc4054a2;
      21922: inst = 32'h8220000;
      21923: inst = 32'h10408000;
      21924: inst = 32'hc4054a3;
      21925: inst = 32'h8220000;
      21926: inst = 32'h10408000;
      21927: inst = 32'hc4054a4;
      21928: inst = 32'h8220000;
      21929: inst = 32'h10408000;
      21930: inst = 32'hc4054a5;
      21931: inst = 32'h8220000;
      21932: inst = 32'h10408000;
      21933: inst = 32'hc4054a6;
      21934: inst = 32'h8220000;
      21935: inst = 32'h10408000;
      21936: inst = 32'hc4054a7;
      21937: inst = 32'h8220000;
      21938: inst = 32'h10408000;
      21939: inst = 32'hc4054a8;
      21940: inst = 32'h8220000;
      21941: inst = 32'h10408000;
      21942: inst = 32'hc4054a9;
      21943: inst = 32'h8220000;
      21944: inst = 32'h10408000;
      21945: inst = 32'hc4054aa;
      21946: inst = 32'h8220000;
      21947: inst = 32'h10408000;
      21948: inst = 32'hc4054ab;
      21949: inst = 32'h8220000;
      21950: inst = 32'h10408000;
      21951: inst = 32'hc4054ac;
      21952: inst = 32'h8220000;
      21953: inst = 32'h10408000;
      21954: inst = 32'hc4054ad;
      21955: inst = 32'h8220000;
      21956: inst = 32'h10408000;
      21957: inst = 32'hc4054ae;
      21958: inst = 32'h8220000;
      21959: inst = 32'h10408000;
      21960: inst = 32'hc4054af;
      21961: inst = 32'h8220000;
      21962: inst = 32'h10408000;
      21963: inst = 32'hc4054b0;
      21964: inst = 32'h8220000;
      21965: inst = 32'h10408000;
      21966: inst = 32'hc4054b1;
      21967: inst = 32'h8220000;
      21968: inst = 32'h10408000;
      21969: inst = 32'hc4054b2;
      21970: inst = 32'h8220000;
      21971: inst = 32'h10408000;
      21972: inst = 32'hc4054b3;
      21973: inst = 32'h8220000;
      21974: inst = 32'h10408000;
      21975: inst = 32'hc4054b4;
      21976: inst = 32'h8220000;
      21977: inst = 32'h10408000;
      21978: inst = 32'hc4054b5;
      21979: inst = 32'h8220000;
      21980: inst = 32'h10408000;
      21981: inst = 32'hc4054b6;
      21982: inst = 32'h8220000;
      21983: inst = 32'h10408000;
      21984: inst = 32'hc4054b7;
      21985: inst = 32'h8220000;
      21986: inst = 32'h10408000;
      21987: inst = 32'hc4054b8;
      21988: inst = 32'h8220000;
      21989: inst = 32'h10408000;
      21990: inst = 32'hc4054b9;
      21991: inst = 32'h8220000;
      21992: inst = 32'h10408000;
      21993: inst = 32'hc4054ba;
      21994: inst = 32'h8220000;
      21995: inst = 32'h10408000;
      21996: inst = 32'hc4054bb;
      21997: inst = 32'h8220000;
      21998: inst = 32'h10408000;
      21999: inst = 32'hc4054bc;
      22000: inst = 32'h8220000;
      22001: inst = 32'h10408000;
      22002: inst = 32'hc4054bd;
      22003: inst = 32'h8220000;
      22004: inst = 32'h10408000;
      22005: inst = 32'hc4054be;
      22006: inst = 32'h8220000;
      22007: inst = 32'h10408000;
      22008: inst = 32'hc4054bf;
      22009: inst = 32'h8220000;
      22010: inst = 32'h10408000;
      22011: inst = 32'hc4054c0;
      22012: inst = 32'h8220000;
      22013: inst = 32'h10408000;
      22014: inst = 32'hc4054c1;
      22015: inst = 32'h8220000;
      22016: inst = 32'h10408000;
      22017: inst = 32'hc4054c2;
      22018: inst = 32'h8220000;
      22019: inst = 32'h10408000;
      22020: inst = 32'hc4054c3;
      22021: inst = 32'h8220000;
      22022: inst = 32'h10408000;
      22023: inst = 32'hc4054c4;
      22024: inst = 32'h8220000;
      22025: inst = 32'h10408000;
      22026: inst = 32'hc4054c5;
      22027: inst = 32'h8220000;
      22028: inst = 32'h10408000;
      22029: inst = 32'hc4054c6;
      22030: inst = 32'h8220000;
      22031: inst = 32'h10408000;
      22032: inst = 32'hc4054c7;
      22033: inst = 32'h8220000;
      22034: inst = 32'h10408000;
      22035: inst = 32'hc4054c8;
      22036: inst = 32'h8220000;
      22037: inst = 32'h10408000;
      22038: inst = 32'hc4054c9;
      22039: inst = 32'h8220000;
      22040: inst = 32'h10408000;
      22041: inst = 32'hc4054ca;
      22042: inst = 32'h8220000;
      22043: inst = 32'h10408000;
      22044: inst = 32'hc4054cb;
      22045: inst = 32'h8220000;
      22046: inst = 32'h10408000;
      22047: inst = 32'hc4054cc;
      22048: inst = 32'h8220000;
      22049: inst = 32'h10408000;
      22050: inst = 32'hc4054cd;
      22051: inst = 32'h8220000;
      22052: inst = 32'h10408000;
      22053: inst = 32'hc4054ce;
      22054: inst = 32'h8220000;
      22055: inst = 32'h10408000;
      22056: inst = 32'hc4054cf;
      22057: inst = 32'h8220000;
      22058: inst = 32'h10408000;
      22059: inst = 32'hc4054d0;
      22060: inst = 32'h8220000;
      22061: inst = 32'h10408000;
      22062: inst = 32'hc4054d1;
      22063: inst = 32'h8220000;
      22064: inst = 32'h10408000;
      22065: inst = 32'hc4054d2;
      22066: inst = 32'h8220000;
      22067: inst = 32'h10408000;
      22068: inst = 32'hc4054d3;
      22069: inst = 32'h8220000;
      22070: inst = 32'h10408000;
      22071: inst = 32'hc4054d4;
      22072: inst = 32'h8220000;
      22073: inst = 32'h10408000;
      22074: inst = 32'hc4054d5;
      22075: inst = 32'h8220000;
      22076: inst = 32'h10408000;
      22077: inst = 32'hc4054d6;
      22078: inst = 32'h8220000;
      22079: inst = 32'h10408000;
      22080: inst = 32'hc4054d7;
      22081: inst = 32'h8220000;
      22082: inst = 32'h10408000;
      22083: inst = 32'hc4054d8;
      22084: inst = 32'h8220000;
      22085: inst = 32'h10408000;
      22086: inst = 32'hc4054d9;
      22087: inst = 32'h8220000;
      22088: inst = 32'h10408000;
      22089: inst = 32'hc4054da;
      22090: inst = 32'h8220000;
      22091: inst = 32'h10408000;
      22092: inst = 32'hc4054db;
      22093: inst = 32'h8220000;
      22094: inst = 32'h10408000;
      22095: inst = 32'hc4054e4;
      22096: inst = 32'h8220000;
      22097: inst = 32'h10408000;
      22098: inst = 32'hc4054e5;
      22099: inst = 32'h8220000;
      22100: inst = 32'h10408000;
      22101: inst = 32'hc4054e6;
      22102: inst = 32'h8220000;
      22103: inst = 32'h10408000;
      22104: inst = 32'hc4054e7;
      22105: inst = 32'h8220000;
      22106: inst = 32'h10408000;
      22107: inst = 32'hc4054e8;
      22108: inst = 32'h8220000;
      22109: inst = 32'h10408000;
      22110: inst = 32'hc4054e9;
      22111: inst = 32'h8220000;
      22112: inst = 32'h10408000;
      22113: inst = 32'hc4054ea;
      22114: inst = 32'h8220000;
      22115: inst = 32'h10408000;
      22116: inst = 32'hc4054eb;
      22117: inst = 32'h8220000;
      22118: inst = 32'h10408000;
      22119: inst = 32'hc4054ec;
      22120: inst = 32'h8220000;
      22121: inst = 32'h10408000;
      22122: inst = 32'hc4054ed;
      22123: inst = 32'h8220000;
      22124: inst = 32'h10408000;
      22125: inst = 32'hc4054ee;
      22126: inst = 32'h8220000;
      22127: inst = 32'h10408000;
      22128: inst = 32'hc4054ef;
      22129: inst = 32'h8220000;
      22130: inst = 32'h10408000;
      22131: inst = 32'hc4054f0;
      22132: inst = 32'h8220000;
      22133: inst = 32'h10408000;
      22134: inst = 32'hc4054f1;
      22135: inst = 32'h8220000;
      22136: inst = 32'h10408000;
      22137: inst = 32'hc4054f2;
      22138: inst = 32'h8220000;
      22139: inst = 32'h10408000;
      22140: inst = 32'hc4054f3;
      22141: inst = 32'h8220000;
      22142: inst = 32'h10408000;
      22143: inst = 32'hc4054f4;
      22144: inst = 32'h8220000;
      22145: inst = 32'h10408000;
      22146: inst = 32'hc4054f5;
      22147: inst = 32'h8220000;
      22148: inst = 32'h10408000;
      22149: inst = 32'hc4054f6;
      22150: inst = 32'h8220000;
      22151: inst = 32'h10408000;
      22152: inst = 32'hc4054f7;
      22153: inst = 32'h8220000;
      22154: inst = 32'h10408000;
      22155: inst = 32'hc4054f8;
      22156: inst = 32'h8220000;
      22157: inst = 32'h10408000;
      22158: inst = 32'hc4054f9;
      22159: inst = 32'h8220000;
      22160: inst = 32'h10408000;
      22161: inst = 32'hc4054fa;
      22162: inst = 32'h8220000;
      22163: inst = 32'h10408000;
      22164: inst = 32'hc4054fb;
      22165: inst = 32'h8220000;
      22166: inst = 32'h10408000;
      22167: inst = 32'hc4054fc;
      22168: inst = 32'h8220000;
      22169: inst = 32'h10408000;
      22170: inst = 32'hc4054fd;
      22171: inst = 32'h8220000;
      22172: inst = 32'h10408000;
      22173: inst = 32'hc4054fe;
      22174: inst = 32'h8220000;
      22175: inst = 32'h10408000;
      22176: inst = 32'hc4054ff;
      22177: inst = 32'h8220000;
      22178: inst = 32'h10408000;
      22179: inst = 32'hc405500;
      22180: inst = 32'h8220000;
      22181: inst = 32'h10408000;
      22182: inst = 32'hc405501;
      22183: inst = 32'h8220000;
      22184: inst = 32'h10408000;
      22185: inst = 32'hc405502;
      22186: inst = 32'h8220000;
      22187: inst = 32'h10408000;
      22188: inst = 32'hc405503;
      22189: inst = 32'h8220000;
      22190: inst = 32'h10408000;
      22191: inst = 32'hc405504;
      22192: inst = 32'h8220000;
      22193: inst = 32'h10408000;
      22194: inst = 32'hc405505;
      22195: inst = 32'h8220000;
      22196: inst = 32'h10408000;
      22197: inst = 32'hc405506;
      22198: inst = 32'h8220000;
      22199: inst = 32'h10408000;
      22200: inst = 32'hc405507;
      22201: inst = 32'h8220000;
      22202: inst = 32'h10408000;
      22203: inst = 32'hc405508;
      22204: inst = 32'h8220000;
      22205: inst = 32'h10408000;
      22206: inst = 32'hc405509;
      22207: inst = 32'h8220000;
      22208: inst = 32'h10408000;
      22209: inst = 32'hc40550a;
      22210: inst = 32'h8220000;
      22211: inst = 32'h10408000;
      22212: inst = 32'hc40550b;
      22213: inst = 32'h8220000;
      22214: inst = 32'h10408000;
      22215: inst = 32'hc40550c;
      22216: inst = 32'h8220000;
      22217: inst = 32'h10408000;
      22218: inst = 32'hc40550d;
      22219: inst = 32'h8220000;
      22220: inst = 32'h10408000;
      22221: inst = 32'hc40550e;
      22222: inst = 32'h8220000;
      22223: inst = 32'h10408000;
      22224: inst = 32'hc40550f;
      22225: inst = 32'h8220000;
      22226: inst = 32'h10408000;
      22227: inst = 32'hc405510;
      22228: inst = 32'h8220000;
      22229: inst = 32'h10408000;
      22230: inst = 32'hc405511;
      22231: inst = 32'h8220000;
      22232: inst = 32'h10408000;
      22233: inst = 32'hc405512;
      22234: inst = 32'h8220000;
      22235: inst = 32'h10408000;
      22236: inst = 32'hc405513;
      22237: inst = 32'h8220000;
      22238: inst = 32'h10408000;
      22239: inst = 32'hc405514;
      22240: inst = 32'h8220000;
      22241: inst = 32'h10408000;
      22242: inst = 32'hc405515;
      22243: inst = 32'h8220000;
      22244: inst = 32'h10408000;
      22245: inst = 32'hc405516;
      22246: inst = 32'h8220000;
      22247: inst = 32'h10408000;
      22248: inst = 32'hc405517;
      22249: inst = 32'h8220000;
      22250: inst = 32'h10408000;
      22251: inst = 32'hc405518;
      22252: inst = 32'h8220000;
      22253: inst = 32'h10408000;
      22254: inst = 32'hc405519;
      22255: inst = 32'h8220000;
      22256: inst = 32'h10408000;
      22257: inst = 32'hc40551a;
      22258: inst = 32'h8220000;
      22259: inst = 32'h10408000;
      22260: inst = 32'hc40551b;
      22261: inst = 32'h8220000;
      22262: inst = 32'h10408000;
      22263: inst = 32'hc40551c;
      22264: inst = 32'h8220000;
      22265: inst = 32'h10408000;
      22266: inst = 32'hc40551d;
      22267: inst = 32'h8220000;
      22268: inst = 32'h10408000;
      22269: inst = 32'hc40551e;
      22270: inst = 32'h8220000;
      22271: inst = 32'h10408000;
      22272: inst = 32'hc40551f;
      22273: inst = 32'h8220000;
      22274: inst = 32'h10408000;
      22275: inst = 32'hc405520;
      22276: inst = 32'h8220000;
      22277: inst = 32'h10408000;
      22278: inst = 32'hc405521;
      22279: inst = 32'h8220000;
      22280: inst = 32'h10408000;
      22281: inst = 32'hc405522;
      22282: inst = 32'h8220000;
      22283: inst = 32'h10408000;
      22284: inst = 32'hc405523;
      22285: inst = 32'h8220000;
      22286: inst = 32'h10408000;
      22287: inst = 32'hc405524;
      22288: inst = 32'h8220000;
      22289: inst = 32'h10408000;
      22290: inst = 32'hc405525;
      22291: inst = 32'h8220000;
      22292: inst = 32'h10408000;
      22293: inst = 32'hc405526;
      22294: inst = 32'h8220000;
      22295: inst = 32'h10408000;
      22296: inst = 32'hc405527;
      22297: inst = 32'h8220000;
      22298: inst = 32'h10408000;
      22299: inst = 32'hc405528;
      22300: inst = 32'h8220000;
      22301: inst = 32'h10408000;
      22302: inst = 32'hc405529;
      22303: inst = 32'h8220000;
      22304: inst = 32'h10408000;
      22305: inst = 32'hc40552a;
      22306: inst = 32'h8220000;
      22307: inst = 32'h10408000;
      22308: inst = 32'hc40552b;
      22309: inst = 32'h8220000;
      22310: inst = 32'h10408000;
      22311: inst = 32'hc40552c;
      22312: inst = 32'h8220000;
      22313: inst = 32'h10408000;
      22314: inst = 32'hc40552d;
      22315: inst = 32'h8220000;
      22316: inst = 32'h10408000;
      22317: inst = 32'hc40552e;
      22318: inst = 32'h8220000;
      22319: inst = 32'h10408000;
      22320: inst = 32'hc40552f;
      22321: inst = 32'h8220000;
      22322: inst = 32'h10408000;
      22323: inst = 32'hc405530;
      22324: inst = 32'h8220000;
      22325: inst = 32'h10408000;
      22326: inst = 32'hc405531;
      22327: inst = 32'h8220000;
      22328: inst = 32'h10408000;
      22329: inst = 32'hc405532;
      22330: inst = 32'h8220000;
      22331: inst = 32'h10408000;
      22332: inst = 32'hc405533;
      22333: inst = 32'h8220000;
      22334: inst = 32'h10408000;
      22335: inst = 32'hc405534;
      22336: inst = 32'h8220000;
      22337: inst = 32'h10408000;
      22338: inst = 32'hc405535;
      22339: inst = 32'h8220000;
      22340: inst = 32'h10408000;
      22341: inst = 32'hc405536;
      22342: inst = 32'h8220000;
      22343: inst = 32'h10408000;
      22344: inst = 32'hc405537;
      22345: inst = 32'h8220000;
      22346: inst = 32'h10408000;
      22347: inst = 32'hc405538;
      22348: inst = 32'h8220000;
      22349: inst = 32'h10408000;
      22350: inst = 32'hc405539;
      22351: inst = 32'h8220000;
      22352: inst = 32'h10408000;
      22353: inst = 32'hc40553a;
      22354: inst = 32'h8220000;
      22355: inst = 32'h10408000;
      22356: inst = 32'hc40553b;
      22357: inst = 32'h8220000;
      22358: inst = 32'hc204a7a;
      22359: inst = 32'h10408000;
      22360: inst = 32'hc4042e7;
      22361: inst = 32'h8220000;
      22362: inst = 32'h10408000;
      22363: inst = 32'hc404338;
      22364: inst = 32'h8220000;
      22365: inst = 32'h10408000;
      22366: inst = 32'hc404346;
      22367: inst = 32'h8220000;
      22368: inst = 32'h10408000;
      22369: inst = 32'hc404399;
      22370: inst = 32'h8220000;
      22371: inst = 32'h10408000;
      22372: inst = 32'hc4053c6;
      22373: inst = 32'h8220000;
      22374: inst = 32'h10408000;
      22375: inst = 32'hc405419;
      22376: inst = 32'h8220000;
      22377: inst = 32'h10408000;
      22378: inst = 32'hc405427;
      22379: inst = 32'h8220000;
      22380: inst = 32'h10408000;
      22381: inst = 32'hc405478;
      22382: inst = 32'h8220000;
      22383: inst = 32'hc20294f;
      22384: inst = 32'h10408000;
      22385: inst = 32'hc4042e8;
      22386: inst = 32'h8220000;
      22387: inst = 32'h10408000;
      22388: inst = 32'hc404337;
      22389: inst = 32'h8220000;
      22390: inst = 32'h10408000;
      22391: inst = 32'hc405428;
      22392: inst = 32'h8220000;
      22393: inst = 32'h10408000;
      22394: inst = 32'hc405477;
      22395: inst = 32'h8220000;
      22396: inst = 32'hc20210b;
      22397: inst = 32'h10408000;
      22398: inst = 32'hc4042e9;
      22399: inst = 32'h8220000;
      22400: inst = 32'h10408000;
      22401: inst = 32'hc4042ea;
      22402: inst = 32'h8220000;
      22403: inst = 32'h10408000;
      22404: inst = 32'hc4042eb;
      22405: inst = 32'h8220000;
      22406: inst = 32'h10408000;
      22407: inst = 32'hc4042ec;
      22408: inst = 32'h8220000;
      22409: inst = 32'h10408000;
      22410: inst = 32'hc4042ed;
      22411: inst = 32'h8220000;
      22412: inst = 32'h10408000;
      22413: inst = 32'hc4042ee;
      22414: inst = 32'h8220000;
      22415: inst = 32'h10408000;
      22416: inst = 32'hc4042ef;
      22417: inst = 32'h8220000;
      22418: inst = 32'h10408000;
      22419: inst = 32'hc4042f0;
      22420: inst = 32'h8220000;
      22421: inst = 32'h10408000;
      22422: inst = 32'hc4042f1;
      22423: inst = 32'h8220000;
      22424: inst = 32'h10408000;
      22425: inst = 32'hc4042f2;
      22426: inst = 32'h8220000;
      22427: inst = 32'h10408000;
      22428: inst = 32'hc4042f3;
      22429: inst = 32'h8220000;
      22430: inst = 32'h10408000;
      22431: inst = 32'hc4042f4;
      22432: inst = 32'h8220000;
      22433: inst = 32'h10408000;
      22434: inst = 32'hc4042f5;
      22435: inst = 32'h8220000;
      22436: inst = 32'h10408000;
      22437: inst = 32'hc4042f6;
      22438: inst = 32'h8220000;
      22439: inst = 32'h10408000;
      22440: inst = 32'hc4042f7;
      22441: inst = 32'h8220000;
      22442: inst = 32'h10408000;
      22443: inst = 32'hc4042f8;
      22444: inst = 32'h8220000;
      22445: inst = 32'h10408000;
      22446: inst = 32'hc4042f9;
      22447: inst = 32'h8220000;
      22448: inst = 32'h10408000;
      22449: inst = 32'hc4042fa;
      22450: inst = 32'h8220000;
      22451: inst = 32'h10408000;
      22452: inst = 32'hc4042fb;
      22453: inst = 32'h8220000;
      22454: inst = 32'h10408000;
      22455: inst = 32'hc4042fc;
      22456: inst = 32'h8220000;
      22457: inst = 32'h10408000;
      22458: inst = 32'hc4042fd;
      22459: inst = 32'h8220000;
      22460: inst = 32'h10408000;
      22461: inst = 32'hc4042fe;
      22462: inst = 32'h8220000;
      22463: inst = 32'h10408000;
      22464: inst = 32'hc4042ff;
      22465: inst = 32'h8220000;
      22466: inst = 32'h10408000;
      22467: inst = 32'hc404300;
      22468: inst = 32'h8220000;
      22469: inst = 32'h10408000;
      22470: inst = 32'hc404301;
      22471: inst = 32'h8220000;
      22472: inst = 32'h10408000;
      22473: inst = 32'hc404302;
      22474: inst = 32'h8220000;
      22475: inst = 32'h10408000;
      22476: inst = 32'hc404303;
      22477: inst = 32'h8220000;
      22478: inst = 32'h10408000;
      22479: inst = 32'hc404304;
      22480: inst = 32'h8220000;
      22481: inst = 32'h10408000;
      22482: inst = 32'hc404305;
      22483: inst = 32'h8220000;
      22484: inst = 32'h10408000;
      22485: inst = 32'hc404306;
      22486: inst = 32'h8220000;
      22487: inst = 32'h10408000;
      22488: inst = 32'hc404307;
      22489: inst = 32'h8220000;
      22490: inst = 32'h10408000;
      22491: inst = 32'hc404308;
      22492: inst = 32'h8220000;
      22493: inst = 32'h10408000;
      22494: inst = 32'hc404309;
      22495: inst = 32'h8220000;
      22496: inst = 32'h10408000;
      22497: inst = 32'hc40430a;
      22498: inst = 32'h8220000;
      22499: inst = 32'h10408000;
      22500: inst = 32'hc40430b;
      22501: inst = 32'h8220000;
      22502: inst = 32'h10408000;
      22503: inst = 32'hc40430c;
      22504: inst = 32'h8220000;
      22505: inst = 32'h10408000;
      22506: inst = 32'hc40430d;
      22507: inst = 32'h8220000;
      22508: inst = 32'h10408000;
      22509: inst = 32'hc40430e;
      22510: inst = 32'h8220000;
      22511: inst = 32'h10408000;
      22512: inst = 32'hc40430f;
      22513: inst = 32'h8220000;
      22514: inst = 32'h10408000;
      22515: inst = 32'hc404310;
      22516: inst = 32'h8220000;
      22517: inst = 32'h10408000;
      22518: inst = 32'hc404311;
      22519: inst = 32'h8220000;
      22520: inst = 32'h10408000;
      22521: inst = 32'hc404312;
      22522: inst = 32'h8220000;
      22523: inst = 32'h10408000;
      22524: inst = 32'hc404313;
      22525: inst = 32'h8220000;
      22526: inst = 32'h10408000;
      22527: inst = 32'hc404314;
      22528: inst = 32'h8220000;
      22529: inst = 32'h10408000;
      22530: inst = 32'hc404315;
      22531: inst = 32'h8220000;
      22532: inst = 32'h10408000;
      22533: inst = 32'hc404316;
      22534: inst = 32'h8220000;
      22535: inst = 32'h10408000;
      22536: inst = 32'hc404317;
      22537: inst = 32'h8220000;
      22538: inst = 32'h10408000;
      22539: inst = 32'hc404318;
      22540: inst = 32'h8220000;
      22541: inst = 32'h10408000;
      22542: inst = 32'hc404319;
      22543: inst = 32'h8220000;
      22544: inst = 32'h10408000;
      22545: inst = 32'hc40431a;
      22546: inst = 32'h8220000;
      22547: inst = 32'h10408000;
      22548: inst = 32'hc40431b;
      22549: inst = 32'h8220000;
      22550: inst = 32'h10408000;
      22551: inst = 32'hc40431c;
      22552: inst = 32'h8220000;
      22553: inst = 32'h10408000;
      22554: inst = 32'hc40431d;
      22555: inst = 32'h8220000;
      22556: inst = 32'h10408000;
      22557: inst = 32'hc40431e;
      22558: inst = 32'h8220000;
      22559: inst = 32'h10408000;
      22560: inst = 32'hc40431f;
      22561: inst = 32'h8220000;
      22562: inst = 32'h10408000;
      22563: inst = 32'hc404320;
      22564: inst = 32'h8220000;
      22565: inst = 32'h10408000;
      22566: inst = 32'hc404321;
      22567: inst = 32'h8220000;
      22568: inst = 32'h10408000;
      22569: inst = 32'hc404322;
      22570: inst = 32'h8220000;
      22571: inst = 32'h10408000;
      22572: inst = 32'hc404323;
      22573: inst = 32'h8220000;
      22574: inst = 32'h10408000;
      22575: inst = 32'hc404324;
      22576: inst = 32'h8220000;
      22577: inst = 32'h10408000;
      22578: inst = 32'hc404325;
      22579: inst = 32'h8220000;
      22580: inst = 32'h10408000;
      22581: inst = 32'hc404326;
      22582: inst = 32'h8220000;
      22583: inst = 32'h10408000;
      22584: inst = 32'hc404327;
      22585: inst = 32'h8220000;
      22586: inst = 32'h10408000;
      22587: inst = 32'hc404328;
      22588: inst = 32'h8220000;
      22589: inst = 32'h10408000;
      22590: inst = 32'hc404329;
      22591: inst = 32'h8220000;
      22592: inst = 32'h10408000;
      22593: inst = 32'hc40432a;
      22594: inst = 32'h8220000;
      22595: inst = 32'h10408000;
      22596: inst = 32'hc40432b;
      22597: inst = 32'h8220000;
      22598: inst = 32'h10408000;
      22599: inst = 32'hc40432c;
      22600: inst = 32'h8220000;
      22601: inst = 32'h10408000;
      22602: inst = 32'hc40432d;
      22603: inst = 32'h8220000;
      22604: inst = 32'h10408000;
      22605: inst = 32'hc40432e;
      22606: inst = 32'h8220000;
      22607: inst = 32'h10408000;
      22608: inst = 32'hc40432f;
      22609: inst = 32'h8220000;
      22610: inst = 32'h10408000;
      22611: inst = 32'hc404330;
      22612: inst = 32'h8220000;
      22613: inst = 32'h10408000;
      22614: inst = 32'hc404331;
      22615: inst = 32'h8220000;
      22616: inst = 32'h10408000;
      22617: inst = 32'hc404332;
      22618: inst = 32'h8220000;
      22619: inst = 32'h10408000;
      22620: inst = 32'hc404333;
      22621: inst = 32'h8220000;
      22622: inst = 32'h10408000;
      22623: inst = 32'hc404334;
      22624: inst = 32'h8220000;
      22625: inst = 32'h10408000;
      22626: inst = 32'hc404335;
      22627: inst = 32'h8220000;
      22628: inst = 32'h10408000;
      22629: inst = 32'hc404336;
      22630: inst = 32'h8220000;
      22631: inst = 32'h10408000;
      22632: inst = 32'hc405429;
      22633: inst = 32'h8220000;
      22634: inst = 32'h10408000;
      22635: inst = 32'hc40542a;
      22636: inst = 32'h8220000;
      22637: inst = 32'h10408000;
      22638: inst = 32'hc40542b;
      22639: inst = 32'h8220000;
      22640: inst = 32'h10408000;
      22641: inst = 32'hc40542c;
      22642: inst = 32'h8220000;
      22643: inst = 32'h10408000;
      22644: inst = 32'hc40542d;
      22645: inst = 32'h8220000;
      22646: inst = 32'h10408000;
      22647: inst = 32'hc40542e;
      22648: inst = 32'h8220000;
      22649: inst = 32'h10408000;
      22650: inst = 32'hc40542f;
      22651: inst = 32'h8220000;
      22652: inst = 32'h10408000;
      22653: inst = 32'hc405430;
      22654: inst = 32'h8220000;
      22655: inst = 32'h10408000;
      22656: inst = 32'hc405431;
      22657: inst = 32'h8220000;
      22658: inst = 32'h10408000;
      22659: inst = 32'hc405432;
      22660: inst = 32'h8220000;
      22661: inst = 32'h10408000;
      22662: inst = 32'hc405433;
      22663: inst = 32'h8220000;
      22664: inst = 32'h10408000;
      22665: inst = 32'hc405434;
      22666: inst = 32'h8220000;
      22667: inst = 32'h10408000;
      22668: inst = 32'hc405435;
      22669: inst = 32'h8220000;
      22670: inst = 32'h10408000;
      22671: inst = 32'hc405436;
      22672: inst = 32'h8220000;
      22673: inst = 32'h10408000;
      22674: inst = 32'hc405437;
      22675: inst = 32'h8220000;
      22676: inst = 32'h10408000;
      22677: inst = 32'hc405438;
      22678: inst = 32'h8220000;
      22679: inst = 32'h10408000;
      22680: inst = 32'hc405439;
      22681: inst = 32'h8220000;
      22682: inst = 32'h10408000;
      22683: inst = 32'hc40543a;
      22684: inst = 32'h8220000;
      22685: inst = 32'h10408000;
      22686: inst = 32'hc40543b;
      22687: inst = 32'h8220000;
      22688: inst = 32'h10408000;
      22689: inst = 32'hc40543c;
      22690: inst = 32'h8220000;
      22691: inst = 32'h10408000;
      22692: inst = 32'hc40543d;
      22693: inst = 32'h8220000;
      22694: inst = 32'h10408000;
      22695: inst = 32'hc40543e;
      22696: inst = 32'h8220000;
      22697: inst = 32'h10408000;
      22698: inst = 32'hc40543f;
      22699: inst = 32'h8220000;
      22700: inst = 32'h10408000;
      22701: inst = 32'hc405440;
      22702: inst = 32'h8220000;
      22703: inst = 32'h10408000;
      22704: inst = 32'hc405441;
      22705: inst = 32'h8220000;
      22706: inst = 32'h10408000;
      22707: inst = 32'hc405442;
      22708: inst = 32'h8220000;
      22709: inst = 32'h10408000;
      22710: inst = 32'hc405443;
      22711: inst = 32'h8220000;
      22712: inst = 32'h10408000;
      22713: inst = 32'hc405444;
      22714: inst = 32'h8220000;
      22715: inst = 32'h10408000;
      22716: inst = 32'hc405445;
      22717: inst = 32'h8220000;
      22718: inst = 32'h10408000;
      22719: inst = 32'hc405446;
      22720: inst = 32'h8220000;
      22721: inst = 32'h10408000;
      22722: inst = 32'hc405447;
      22723: inst = 32'h8220000;
      22724: inst = 32'h10408000;
      22725: inst = 32'hc405448;
      22726: inst = 32'h8220000;
      22727: inst = 32'h10408000;
      22728: inst = 32'hc405449;
      22729: inst = 32'h8220000;
      22730: inst = 32'h10408000;
      22731: inst = 32'hc40544a;
      22732: inst = 32'h8220000;
      22733: inst = 32'h10408000;
      22734: inst = 32'hc40544b;
      22735: inst = 32'h8220000;
      22736: inst = 32'h10408000;
      22737: inst = 32'hc40544c;
      22738: inst = 32'h8220000;
      22739: inst = 32'h10408000;
      22740: inst = 32'hc40544d;
      22741: inst = 32'h8220000;
      22742: inst = 32'h10408000;
      22743: inst = 32'hc40544e;
      22744: inst = 32'h8220000;
      22745: inst = 32'h10408000;
      22746: inst = 32'hc40544f;
      22747: inst = 32'h8220000;
      22748: inst = 32'h10408000;
      22749: inst = 32'hc405450;
      22750: inst = 32'h8220000;
      22751: inst = 32'h10408000;
      22752: inst = 32'hc405451;
      22753: inst = 32'h8220000;
      22754: inst = 32'h10408000;
      22755: inst = 32'hc405452;
      22756: inst = 32'h8220000;
      22757: inst = 32'h10408000;
      22758: inst = 32'hc405453;
      22759: inst = 32'h8220000;
      22760: inst = 32'h10408000;
      22761: inst = 32'hc405454;
      22762: inst = 32'h8220000;
      22763: inst = 32'h10408000;
      22764: inst = 32'hc405455;
      22765: inst = 32'h8220000;
      22766: inst = 32'h10408000;
      22767: inst = 32'hc405456;
      22768: inst = 32'h8220000;
      22769: inst = 32'h10408000;
      22770: inst = 32'hc405457;
      22771: inst = 32'h8220000;
      22772: inst = 32'h10408000;
      22773: inst = 32'hc405458;
      22774: inst = 32'h8220000;
      22775: inst = 32'h10408000;
      22776: inst = 32'hc405459;
      22777: inst = 32'h8220000;
      22778: inst = 32'h10408000;
      22779: inst = 32'hc40545a;
      22780: inst = 32'h8220000;
      22781: inst = 32'h10408000;
      22782: inst = 32'hc40545b;
      22783: inst = 32'h8220000;
      22784: inst = 32'h10408000;
      22785: inst = 32'hc40545c;
      22786: inst = 32'h8220000;
      22787: inst = 32'h10408000;
      22788: inst = 32'hc40545d;
      22789: inst = 32'h8220000;
      22790: inst = 32'h10408000;
      22791: inst = 32'hc40545e;
      22792: inst = 32'h8220000;
      22793: inst = 32'h10408000;
      22794: inst = 32'hc40545f;
      22795: inst = 32'h8220000;
      22796: inst = 32'h10408000;
      22797: inst = 32'hc405460;
      22798: inst = 32'h8220000;
      22799: inst = 32'h10408000;
      22800: inst = 32'hc405461;
      22801: inst = 32'h8220000;
      22802: inst = 32'h10408000;
      22803: inst = 32'hc405462;
      22804: inst = 32'h8220000;
      22805: inst = 32'h10408000;
      22806: inst = 32'hc405463;
      22807: inst = 32'h8220000;
      22808: inst = 32'h10408000;
      22809: inst = 32'hc405464;
      22810: inst = 32'h8220000;
      22811: inst = 32'h10408000;
      22812: inst = 32'hc405465;
      22813: inst = 32'h8220000;
      22814: inst = 32'h10408000;
      22815: inst = 32'hc405466;
      22816: inst = 32'h8220000;
      22817: inst = 32'h10408000;
      22818: inst = 32'hc405467;
      22819: inst = 32'h8220000;
      22820: inst = 32'h10408000;
      22821: inst = 32'hc405468;
      22822: inst = 32'h8220000;
      22823: inst = 32'h10408000;
      22824: inst = 32'hc405469;
      22825: inst = 32'h8220000;
      22826: inst = 32'h10408000;
      22827: inst = 32'hc40546a;
      22828: inst = 32'h8220000;
      22829: inst = 32'h10408000;
      22830: inst = 32'hc40546b;
      22831: inst = 32'h8220000;
      22832: inst = 32'h10408000;
      22833: inst = 32'hc40546c;
      22834: inst = 32'h8220000;
      22835: inst = 32'h10408000;
      22836: inst = 32'hc40546d;
      22837: inst = 32'h8220000;
      22838: inst = 32'h10408000;
      22839: inst = 32'hc40546e;
      22840: inst = 32'h8220000;
      22841: inst = 32'h10408000;
      22842: inst = 32'hc40546f;
      22843: inst = 32'h8220000;
      22844: inst = 32'h10408000;
      22845: inst = 32'hc405470;
      22846: inst = 32'h8220000;
      22847: inst = 32'h10408000;
      22848: inst = 32'hc405471;
      22849: inst = 32'h8220000;
      22850: inst = 32'h10408000;
      22851: inst = 32'hc405472;
      22852: inst = 32'h8220000;
      22853: inst = 32'h10408000;
      22854: inst = 32'hc405473;
      22855: inst = 32'h8220000;
      22856: inst = 32'h10408000;
      22857: inst = 32'hc405474;
      22858: inst = 32'h8220000;
      22859: inst = 32'h10408000;
      22860: inst = 32'hc405475;
      22861: inst = 32'h8220000;
      22862: inst = 32'h10408000;
      22863: inst = 32'hc405476;
      22864: inst = 32'h8220000;
      22865: inst = 32'hc200864;
      22866: inst = 32'h10408000;
      22867: inst = 32'hc404347;
      22868: inst = 32'h8220000;
      22869: inst = 32'h10408000;
      22870: inst = 32'hc404398;
      22871: inst = 32'h8220000;
      22872: inst = 32'h10408000;
      22873: inst = 32'hc4053c7;
      22874: inst = 32'h8220000;
      22875: inst = 32'h10408000;
      22876: inst = 32'hc405418;
      22877: inst = 32'h8220000;
      22878: inst = 32'hc20294e;
      22879: inst = 32'h10408000;
      22880: inst = 32'hc4043a6;
      22881: inst = 32'h8220000;
      22882: inst = 32'h10408000;
      22883: inst = 32'hc4043f9;
      22884: inst = 32'h8220000;
      22885: inst = 32'h10408000;
      22886: inst = 32'hc405366;
      22887: inst = 32'h8220000;
      22888: inst = 32'h10408000;
      22889: inst = 32'hc4053b9;
      22890: inst = 32'h8220000;
      22891: inst = 32'hc2018ea;
      22892: inst = 32'h10408000;
      22893: inst = 32'hc404406;
      22894: inst = 32'h8220000;
      22895: inst = 32'h10408000;
      22896: inst = 32'hc404459;
      22897: inst = 32'h8220000;
      22898: inst = 32'h10408000;
      22899: inst = 32'hc404466;
      22900: inst = 32'h8220000;
      22901: inst = 32'h10408000;
      22902: inst = 32'hc4044b9;
      22903: inst = 32'h8220000;
      22904: inst = 32'h10408000;
      22905: inst = 32'hc4044c6;
      22906: inst = 32'h8220000;
      22907: inst = 32'h10408000;
      22908: inst = 32'hc404519;
      22909: inst = 32'h8220000;
      22910: inst = 32'h10408000;
      22911: inst = 32'hc404526;
      22912: inst = 32'h8220000;
      22913: inst = 32'h10408000;
      22914: inst = 32'hc404579;
      22915: inst = 32'h8220000;
      22916: inst = 32'h10408000;
      22917: inst = 32'hc404586;
      22918: inst = 32'h8220000;
      22919: inst = 32'h10408000;
      22920: inst = 32'hc4045d9;
      22921: inst = 32'h8220000;
      22922: inst = 32'h10408000;
      22923: inst = 32'hc4045e6;
      22924: inst = 32'h8220000;
      22925: inst = 32'h10408000;
      22926: inst = 32'hc404639;
      22927: inst = 32'h8220000;
      22928: inst = 32'h10408000;
      22929: inst = 32'hc404646;
      22930: inst = 32'h8220000;
      22931: inst = 32'h10408000;
      22932: inst = 32'hc404699;
      22933: inst = 32'h8220000;
      22934: inst = 32'h10408000;
      22935: inst = 32'hc4046a6;
      22936: inst = 32'h8220000;
      22937: inst = 32'h10408000;
      22938: inst = 32'hc4046f9;
      22939: inst = 32'h8220000;
      22940: inst = 32'h10408000;
      22941: inst = 32'hc404706;
      22942: inst = 32'h8220000;
      22943: inst = 32'h10408000;
      22944: inst = 32'hc404759;
      22945: inst = 32'h8220000;
      22946: inst = 32'h10408000;
      22947: inst = 32'hc404766;
      22948: inst = 32'h8220000;
      22949: inst = 32'h10408000;
      22950: inst = 32'hc4047b9;
      22951: inst = 32'h8220000;
      22952: inst = 32'h10408000;
      22953: inst = 32'hc4047c6;
      22954: inst = 32'h8220000;
      22955: inst = 32'h10408000;
      22956: inst = 32'hc404819;
      22957: inst = 32'h8220000;
      22958: inst = 32'h10408000;
      22959: inst = 32'hc404826;
      22960: inst = 32'h8220000;
      22961: inst = 32'h10408000;
      22962: inst = 32'hc404879;
      22963: inst = 32'h8220000;
      22964: inst = 32'h10408000;
      22965: inst = 32'hc404886;
      22966: inst = 32'h8220000;
      22967: inst = 32'h10408000;
      22968: inst = 32'hc4048d9;
      22969: inst = 32'h8220000;
      22970: inst = 32'h10408000;
      22971: inst = 32'hc4048e6;
      22972: inst = 32'h8220000;
      22973: inst = 32'h10408000;
      22974: inst = 32'hc404939;
      22975: inst = 32'h8220000;
      22976: inst = 32'h10408000;
      22977: inst = 32'hc404946;
      22978: inst = 32'h8220000;
      22979: inst = 32'h10408000;
      22980: inst = 32'hc404999;
      22981: inst = 32'h8220000;
      22982: inst = 32'h10408000;
      22983: inst = 32'hc4049a6;
      22984: inst = 32'h8220000;
      22985: inst = 32'h10408000;
      22986: inst = 32'hc4049f9;
      22987: inst = 32'h8220000;
      22988: inst = 32'h10408000;
      22989: inst = 32'hc404a06;
      22990: inst = 32'h8220000;
      22991: inst = 32'h10408000;
      22992: inst = 32'hc404a59;
      22993: inst = 32'h8220000;
      22994: inst = 32'h10408000;
      22995: inst = 32'hc404a66;
      22996: inst = 32'h8220000;
      22997: inst = 32'h10408000;
      22998: inst = 32'hc404ab9;
      22999: inst = 32'h8220000;
      23000: inst = 32'h10408000;
      23001: inst = 32'hc404ac6;
      23002: inst = 32'h8220000;
      23003: inst = 32'h10408000;
      23004: inst = 32'hc404b19;
      23005: inst = 32'h8220000;
      23006: inst = 32'h10408000;
      23007: inst = 32'hc404b26;
      23008: inst = 32'h8220000;
      23009: inst = 32'h10408000;
      23010: inst = 32'hc404b79;
      23011: inst = 32'h8220000;
      23012: inst = 32'h10408000;
      23013: inst = 32'hc404b86;
      23014: inst = 32'h8220000;
      23015: inst = 32'h10408000;
      23016: inst = 32'hc404bd9;
      23017: inst = 32'h8220000;
      23018: inst = 32'h10408000;
      23019: inst = 32'hc404be6;
      23020: inst = 32'h8220000;
      23021: inst = 32'h10408000;
      23022: inst = 32'hc404c39;
      23023: inst = 32'h8220000;
      23024: inst = 32'h10408000;
      23025: inst = 32'hc404c46;
      23026: inst = 32'h8220000;
      23027: inst = 32'h10408000;
      23028: inst = 32'hc404c99;
      23029: inst = 32'h8220000;
      23030: inst = 32'h10408000;
      23031: inst = 32'hc404ca6;
      23032: inst = 32'h8220000;
      23033: inst = 32'h10408000;
      23034: inst = 32'hc404cf9;
      23035: inst = 32'h8220000;
      23036: inst = 32'h10408000;
      23037: inst = 32'hc404d06;
      23038: inst = 32'h8220000;
      23039: inst = 32'h10408000;
      23040: inst = 32'hc404d59;
      23041: inst = 32'h8220000;
      23042: inst = 32'h10408000;
      23043: inst = 32'hc404d66;
      23044: inst = 32'h8220000;
      23045: inst = 32'h10408000;
      23046: inst = 32'hc404db9;
      23047: inst = 32'h8220000;
      23048: inst = 32'h10408000;
      23049: inst = 32'hc404dc6;
      23050: inst = 32'h8220000;
      23051: inst = 32'h10408000;
      23052: inst = 32'hc404e19;
      23053: inst = 32'h8220000;
      23054: inst = 32'h10408000;
      23055: inst = 32'hc404e26;
      23056: inst = 32'h8220000;
      23057: inst = 32'h10408000;
      23058: inst = 32'hc404e79;
      23059: inst = 32'h8220000;
      23060: inst = 32'h10408000;
      23061: inst = 32'hc404e86;
      23062: inst = 32'h8220000;
      23063: inst = 32'h10408000;
      23064: inst = 32'hc404ed9;
      23065: inst = 32'h8220000;
      23066: inst = 32'h10408000;
      23067: inst = 32'hc404ee6;
      23068: inst = 32'h8220000;
      23069: inst = 32'h10408000;
      23070: inst = 32'hc404f39;
      23071: inst = 32'h8220000;
      23072: inst = 32'h10408000;
      23073: inst = 32'hc404f46;
      23074: inst = 32'h8220000;
      23075: inst = 32'h10408000;
      23076: inst = 32'hc404f99;
      23077: inst = 32'h8220000;
      23078: inst = 32'h10408000;
      23079: inst = 32'hc404fa6;
      23080: inst = 32'h8220000;
      23081: inst = 32'h10408000;
      23082: inst = 32'hc404ff9;
      23083: inst = 32'h8220000;
      23084: inst = 32'h10408000;
      23085: inst = 32'hc405006;
      23086: inst = 32'h8220000;
      23087: inst = 32'h10408000;
      23088: inst = 32'hc405059;
      23089: inst = 32'h8220000;
      23090: inst = 32'h10408000;
      23091: inst = 32'hc405066;
      23092: inst = 32'h8220000;
      23093: inst = 32'h10408000;
      23094: inst = 32'hc4050b9;
      23095: inst = 32'h8220000;
      23096: inst = 32'h10408000;
      23097: inst = 32'hc4050c6;
      23098: inst = 32'h8220000;
      23099: inst = 32'h10408000;
      23100: inst = 32'hc405119;
      23101: inst = 32'h8220000;
      23102: inst = 32'h10408000;
      23103: inst = 32'hc405126;
      23104: inst = 32'h8220000;
      23105: inst = 32'h10408000;
      23106: inst = 32'hc405179;
      23107: inst = 32'h8220000;
      23108: inst = 32'h10408000;
      23109: inst = 32'hc405186;
      23110: inst = 32'h8220000;
      23111: inst = 32'h10408000;
      23112: inst = 32'hc4051d9;
      23113: inst = 32'h8220000;
      23114: inst = 32'h10408000;
      23115: inst = 32'hc4051e6;
      23116: inst = 32'h8220000;
      23117: inst = 32'h10408000;
      23118: inst = 32'hc405239;
      23119: inst = 32'h8220000;
      23120: inst = 32'h10408000;
      23121: inst = 32'hc405246;
      23122: inst = 32'h8220000;
      23123: inst = 32'h10408000;
      23124: inst = 32'hc405299;
      23125: inst = 32'h8220000;
      23126: inst = 32'h10408000;
      23127: inst = 32'hc4052a6;
      23128: inst = 32'h8220000;
      23129: inst = 32'h10408000;
      23130: inst = 32'hc4052f9;
      23131: inst = 32'h8220000;
      23132: inst = 32'h10408000;
      23133: inst = 32'hc405306;
      23134: inst = 32'h8220000;
      23135: inst = 32'h10408000;
      23136: inst = 32'hc405359;
      23137: inst = 32'h8220000;
      23138: inst = 32'hc206b4d;
      23139: inst = 32'h10408000;
      23140: inst = 32'hc40464e;
      23141: inst = 32'h8220000;
      23142: inst = 32'h10408000;
      23143: inst = 32'hc404690;
      23144: inst = 32'h8220000;
      23145: inst = 32'h10408000;
      23146: inst = 32'hc4046ae;
      23147: inst = 32'h8220000;
      23148: inst = 32'h10408000;
      23149: inst = 32'hc4046f0;
      23150: inst = 32'h8220000;
      23151: inst = 32'h10408000;
      23152: inst = 32'hc4047d3;
      23153: inst = 32'h8220000;
      23154: inst = 32'h10408000;
      23155: inst = 32'hc4047dd;
      23156: inst = 32'h8220000;
      23157: inst = 32'h10408000;
      23158: inst = 32'hc404800;
      23159: inst = 32'h8220000;
      23160: inst = 32'h10408000;
      23161: inst = 32'hc40483a;
      23162: inst = 32'h8220000;
      23163: inst = 32'h10408000;
      23164: inst = 32'hc40485d;
      23165: inst = 32'h8220000;
      23166: inst = 32'h10408000;
      23167: inst = 32'hc4049b8;
      23168: inst = 32'h8220000;
      23169: inst = 32'h10408000;
      23170: inst = 32'hc4049c7;
      23171: inst = 32'h8220000;
      23172: inst = 32'h10408000;
      23173: inst = 32'hc4049e5;
      23174: inst = 32'h8220000;
      23175: inst = 32'h10408000;
      23176: inst = 32'hc4049f0;
      23177: inst = 32'h8220000;
      23178: inst = 32'h10408000;
      23179: inst = 32'hc404cb1;
      23180: inst = 32'h8220000;
      23181: inst = 32'h10408000;
      23182: inst = 32'hc404cf2;
      23183: inst = 32'h8220000;
      23184: inst = 32'h10408000;
      23185: inst = 32'hc404dda;
      23186: inst = 32'h8220000;
      23187: inst = 32'h10408000;
      23188: inst = 32'hc404e5c;
      23189: inst = 32'h8220000;
      23190: inst = 32'h10408000;
      23191: inst = 32'hc404e6b;
      23192: inst = 32'h8220000;
      23193: inst = 32'h10408000;
      23194: inst = 32'hc404e96;
      23195: inst = 32'h8220000;
      23196: inst = 32'h10408000;
      23197: inst = 32'hc404eaf;
      23198: inst = 32'h8220000;
      23199: inst = 32'h10408000;
      23200: inst = 32'hc404fb6;
      23201: inst = 32'h8220000;
      23202: inst = 32'h10408000;
      23203: inst = 32'hc404fcf;
      23204: inst = 32'h8220000;
      23205: inst = 32'h10408000;
      23206: inst = 32'hc40501a;
      23207: inst = 32'h8220000;
      23208: inst = 32'hc20ad55;
      23209: inst = 32'h10408000;
      23210: inst = 32'hc40464f;
      23211: inst = 32'h8220000;
      23212: inst = 32'h10408000;
      23213: inst = 32'hc404692;
      23214: inst = 32'h8220000;
      23215: inst = 32'h10408000;
      23216: inst = 32'hc404809;
      23217: inst = 32'h8220000;
      23218: inst = 32'h10408000;
      23219: inst = 32'hc40483d;
      23220: inst = 32'h8220000;
      23221: inst = 32'h10408000;
      23222: inst = 32'hc404860;
      23223: inst = 32'h8220000;
      23224: inst = 32'h10408000;
      23225: inst = 32'hc404e58;
      23226: inst = 32'h8220000;
      23227: inst = 32'h10408000;
      23228: inst = 32'hc404e59;
      23229: inst = 32'h8220000;
      23230: inst = 32'h10408000;
      23231: inst = 32'hc404e67;
      23232: inst = 32'h8220000;
      23233: inst = 32'h10408000;
      23234: inst = 32'hc404e68;
      23235: inst = 32'h8220000;
      23236: inst = 32'h10408000;
      23237: inst = 32'hc404f19;
      23238: inst = 32'h8220000;
      23239: inst = 32'h10408000;
      23240: inst = 32'hc404f28;
      23241: inst = 32'h8220000;
      23242: inst = 32'h10408000;
      23243: inst = 32'hc404f4f;
      23244: inst = 32'h8220000;
      23245: inst = 32'h10408000;
      23246: inst = 32'hc404fc3;
      23247: inst = 32'h8220000;
      23248: inst = 32'h10408000;
      23249: inst = 32'hc404fcd;
      23250: inst = 32'h8220000;
      23251: inst = 32'h10408000;
      23252: inst = 32'hc404fe1;
      23253: inst = 32'h8220000;
      23254: inst = 32'h10408000;
      23255: inst = 32'hc404ff0;
      23256: inst = 32'h8220000;
      23257: inst = 32'h10408000;
      23258: inst = 32'hc40500e;
      23259: inst = 32'h8220000;
      23260: inst = 32'h10408000;
      23261: inst = 32'hc405054;
      23262: inst = 32'h8220000;
      23263: inst = 32'hc202124;
      23264: inst = 32'h10408000;
      23265: inst = 32'hc404650;
      23266: inst = 32'h8220000;
      23267: inst = 32'h10408000;
      23268: inst = 32'hc404772;
      23269: inst = 32'h8220000;
      23270: inst = 32'h10408000;
      23271: inst = 32'hc40477a;
      23272: inst = 32'h8220000;
      23273: inst = 32'h10408000;
      23274: inst = 32'hc40478b;
      23275: inst = 32'h8220000;
      23276: inst = 32'h10408000;
      23277: inst = 32'hc404793;
      23278: inst = 32'h8220000;
      23279: inst = 32'h10408000;
      23280: inst = 32'hc404795;
      23281: inst = 32'h8220000;
      23282: inst = 32'h10408000;
      23283: inst = 32'hc40479a;
      23284: inst = 32'h8220000;
      23285: inst = 32'h10408000;
      23286: inst = 32'hc40479d;
      23287: inst = 32'h8220000;
      23288: inst = 32'h10408000;
      23289: inst = 32'hc4047ae;
      23290: inst = 32'h8220000;
      23291: inst = 32'h10408000;
      23292: inst = 32'hc404847;
      23293: inst = 32'h8220000;
      23294: inst = 32'h10408000;
      23295: inst = 32'hc404971;
      23296: inst = 32'h8220000;
      23297: inst = 32'h10408000;
      23298: inst = 32'hc40498a;
      23299: inst = 32'h8220000;
      23300: inst = 32'h10408000;
      23301: inst = 32'hc404a10;
      23302: inst = 32'h8220000;
      23303: inst = 32'h10408000;
      23304: inst = 32'hc404a18;
      23305: inst = 32'h8220000;
      23306: inst = 32'h10408000;
      23307: inst = 32'hc404a35;
      23308: inst = 32'h8220000;
      23309: inst = 32'h10408000;
      23310: inst = 32'hc404a3b;
      23311: inst = 32'h8220000;
      23312: inst = 32'h10408000;
      23313: inst = 32'hc404a45;
      23314: inst = 32'h8220000;
      23315: inst = 32'h10408000;
      23316: inst = 32'hc404a50;
      23317: inst = 32'h8220000;
      23318: inst = 32'h10408000;
      23319: inst = 32'hc404d21;
      23320: inst = 32'h8220000;
      23321: inst = 32'h10408000;
      23322: inst = 32'hc404d2b;
      23323: inst = 32'h8220000;
      23324: inst = 32'h10408000;
      23325: inst = 32'hc404d3f;
      23326: inst = 32'h8220000;
      23327: inst = 32'h10408000;
      23328: inst = 32'hc404d44;
      23329: inst = 32'h8220000;
      23330: inst = 32'h10408000;
      23331: inst = 32'hc404dcc;
      23332: inst = 32'h8220000;
      23333: inst = 32'h10408000;
      23334: inst = 32'hc404dcf;
      23335: inst = 32'h8220000;
      23336: inst = 32'h10408000;
      23337: inst = 32'hc404dd6;
      23338: inst = 32'h8220000;
      23339: inst = 32'h10408000;
      23340: inst = 32'hc404def;
      23341: inst = 32'h8220000;
      23342: inst = 32'h10408000;
      23343: inst = 32'hc404e98;
      23344: inst = 32'h8220000;
      23345: inst = 32'h10408000;
      23346: inst = 32'hc404eb1;
      23347: inst = 32'h8220000;
      23348: inst = 32'h10408000;
      23349: inst = 32'hc404fac;
      23350: inst = 32'h8220000;
      23351: inst = 32'h10408000;
      23352: inst = 32'hc404fb8;
      23353: inst = 32'h8220000;
      23354: inst = 32'h10408000;
      23355: inst = 32'hc404fd1;
      23356: inst = 32'h8220000;
      23357: inst = 32'h10408000;
      23358: inst = 32'hc404fd3;
      23359: inst = 32'h8220000;
      23360: inst = 32'h10408000;
      23361: inst = 32'hc40506b;
      23362: inst = 32'h8220000;
      23363: inst = 32'h10408000;
      23364: inst = 32'hc405076;
      23365: inst = 32'h8220000;
      23366: inst = 32'h10408000;
      23367: inst = 32'hc405078;
      23368: inst = 32'h8220000;
      23369: inst = 32'h10408000;
      23370: inst = 32'hc405081;
      23371: inst = 32'h8220000;
      23372: inst = 32'h10408000;
      23373: inst = 32'hc40508b;
      23374: inst = 32'h8220000;
      23375: inst = 32'h10408000;
      23376: inst = 32'hc40508f;
      23377: inst = 32'h8220000;
      23378: inst = 32'h10408000;
      23379: inst = 32'hc405091;
      23380: inst = 32'h8220000;
      23381: inst = 32'h10408000;
      23382: inst = 32'hc40509f;
      23383: inst = 32'h8220000;
      23384: inst = 32'h10408000;
      23385: inst = 32'hc4050a4;
      23386: inst = 32'h8220000;
      23387: inst = 32'h10408000;
      23388: inst = 32'hc4050ad;
      23389: inst = 32'h8220000;
      23390: inst = 32'hc209cf3;
      23391: inst = 32'h10408000;
      23392: inst = 32'hc404691;
      23393: inst = 32'h8220000;
      23394: inst = 32'h10408000;
      23395: inst = 32'hc4046f1;
      23396: inst = 32'h8220000;
      23397: inst = 32'h10408000;
      23398: inst = 32'hc404715;
      23399: inst = 32'h8220000;
      23400: inst = 32'h10408000;
      23401: inst = 32'hc404716;
      23402: inst = 32'h8220000;
      23403: inst = 32'h10408000;
      23404: inst = 32'hc404724;
      23405: inst = 32'h8220000;
      23406: inst = 32'h10408000;
      23407: inst = 32'hc404725;
      23408: inst = 32'h8220000;
      23409: inst = 32'h10408000;
      23410: inst = 32'hc404742;
      23411: inst = 32'h8220000;
      23412: inst = 32'h10408000;
      23413: inst = 32'hc404743;
      23414: inst = 32'h8220000;
      23415: inst = 32'h10408000;
      23416: inst = 32'hc404776;
      23417: inst = 32'h8220000;
      23418: inst = 32'h10408000;
      23419: inst = 32'hc404785;
      23420: inst = 32'h8220000;
      23421: inst = 32'h10408000;
      23422: inst = 32'hc4047a3;
      23423: inst = 32'h8220000;
      23424: inst = 32'h10408000;
      23425: inst = 32'hc4047d4;
      23426: inst = 32'h8220000;
      23427: inst = 32'h10408000;
      23428: inst = 32'hc4047d7;
      23429: inst = 32'h8220000;
      23430: inst = 32'h10408000;
      23431: inst = 32'hc4047db;
      23432: inst = 32'h8220000;
      23433: inst = 32'h10408000;
      23434: inst = 32'hc4047e3;
      23435: inst = 32'h8220000;
      23436: inst = 32'h10408000;
      23437: inst = 32'hc4047e6;
      23438: inst = 32'h8220000;
      23439: inst = 32'h10408000;
      23440: inst = 32'hc4047ea;
      23441: inst = 32'h8220000;
      23442: inst = 32'h10408000;
      23443: inst = 32'hc4047f4;
      23444: inst = 32'h8220000;
      23445: inst = 32'h10408000;
      23446: inst = 32'hc4047f9;
      23447: inst = 32'h8220000;
      23448: inst = 32'h10408000;
      23449: inst = 32'hc4047fe;
      23450: inst = 32'h8220000;
      23451: inst = 32'h10408000;
      23452: inst = 32'hc404801;
      23453: inst = 32'h8220000;
      23454: inst = 32'h10408000;
      23455: inst = 32'hc404804;
      23456: inst = 32'h8220000;
      23457: inst = 32'h10408000;
      23458: inst = 32'hc404806;
      23459: inst = 32'h8220000;
      23460: inst = 32'h10408000;
      23461: inst = 32'hc404808;
      23462: inst = 32'h8220000;
      23463: inst = 32'h10408000;
      23464: inst = 32'hc40480d;
      23465: inst = 32'h8220000;
      23466: inst = 32'h10408000;
      23467: inst = 32'hc404836;
      23468: inst = 32'h8220000;
      23469: inst = 32'h10408000;
      23470: inst = 32'hc40483c;
      23471: inst = 32'h8220000;
      23472: inst = 32'h10408000;
      23473: inst = 32'hc404845;
      23474: inst = 32'h8220000;
      23475: inst = 32'h10408000;
      23476: inst = 32'hc404856;
      23477: inst = 32'h8220000;
      23478: inst = 32'h10408000;
      23479: inst = 32'hc40485f;
      23480: inst = 32'h8220000;
      23481: inst = 32'h10408000;
      23482: inst = 32'hc404863;
      23483: inst = 32'h8220000;
      23484: inst = 32'h10408000;
      23485: inst = 32'hc40486a;
      23486: inst = 32'h8220000;
      23487: inst = 32'h10408000;
      23488: inst = 32'hc404896;
      23489: inst = 32'h8220000;
      23490: inst = 32'h10408000;
      23491: inst = 32'hc40489c;
      23492: inst = 32'h8220000;
      23493: inst = 32'h10408000;
      23494: inst = 32'hc4048a5;
      23495: inst = 32'h8220000;
      23496: inst = 32'h10408000;
      23497: inst = 32'hc4048bf;
      23498: inst = 32'h8220000;
      23499: inst = 32'h10408000;
      23500: inst = 32'hc4048c3;
      23501: inst = 32'h8220000;
      23502: inst = 32'h10408000;
      23503: inst = 32'hc4048f6;
      23504: inst = 32'h8220000;
      23505: inst = 32'h10408000;
      23506: inst = 32'hc4048fc;
      23507: inst = 32'h8220000;
      23508: inst = 32'h10408000;
      23509: inst = 32'hc404905;
      23510: inst = 32'h8220000;
      23511: inst = 32'h10408000;
      23512: inst = 32'hc40491f;
      23513: inst = 32'h8220000;
      23514: inst = 32'h10408000;
      23515: inst = 32'hc404923;
      23516: inst = 32'h8220000;
      23517: inst = 32'h10408000;
      23518: inst = 32'hc404956;
      23519: inst = 32'h8220000;
      23520: inst = 32'h10408000;
      23521: inst = 32'hc404958;
      23522: inst = 32'h8220000;
      23523: inst = 32'h10408000;
      23524: inst = 32'hc40495c;
      23525: inst = 32'h8220000;
      23526: inst = 32'h10408000;
      23527: inst = 32'hc404965;
      23528: inst = 32'h8220000;
      23529: inst = 32'h10408000;
      23530: inst = 32'hc404967;
      23531: inst = 32'h8220000;
      23532: inst = 32'h10408000;
      23533: inst = 32'hc404976;
      23534: inst = 32'h8220000;
      23535: inst = 32'h10408000;
      23536: inst = 32'hc40497f;
      23537: inst = 32'h8220000;
      23538: inst = 32'h10408000;
      23539: inst = 32'hc404983;
      23540: inst = 32'h8220000;
      23541: inst = 32'h10408000;
      23542: inst = 32'hc404985;
      23543: inst = 32'h8220000;
      23544: inst = 32'h10408000;
      23545: inst = 32'hc4049b1;
      23546: inst = 32'h8220000;
      23547: inst = 32'h10408000;
      23548: inst = 32'hc4049b5;
      23549: inst = 32'h8220000;
      23550: inst = 32'h10408000;
      23551: inst = 32'hc4049ba;
      23552: inst = 32'h8220000;
      23553: inst = 32'h10408000;
      23554: inst = 32'hc4049c4;
      23555: inst = 32'h8220000;
      23556: inst = 32'h10408000;
      23557: inst = 32'hc4049ca;
      23558: inst = 32'h8220000;
      23559: inst = 32'h10408000;
      23560: inst = 32'hc4049d4;
      23561: inst = 32'h8220000;
      23562: inst = 32'h10408000;
      23563: inst = 32'hc4049d9;
      23564: inst = 32'h8220000;
      23565: inst = 32'h10408000;
      23566: inst = 32'hc4049dd;
      23567: inst = 32'h8220000;
      23568: inst = 32'h10408000;
      23569: inst = 32'hc4049e2;
      23570: inst = 32'h8220000;
      23571: inst = 32'h10408000;
      23572: inst = 32'hc4049e6;
      23573: inst = 32'h8220000;
      23574: inst = 32'h10408000;
      23575: inst = 32'hc4049e8;
      23576: inst = 32'h8220000;
      23577: inst = 32'h10408000;
      23578: inst = 32'hc4049ed;
      23579: inst = 32'h8220000;
      23580: inst = 32'h10408000;
      23581: inst = 32'hc4049f1;
      23582: inst = 32'h8220000;
      23583: inst = 32'h10408000;
      23584: inst = 32'hc4049f3;
      23585: inst = 32'h8220000;
      23586: inst = 32'h10408000;
      23587: inst = 32'hc404cb0;
      23588: inst = 32'h8220000;
      23589: inst = 32'h10408000;
      23590: inst = 32'hc404cf1;
      23591: inst = 32'h8220000;
      23592: inst = 32'h10408000;
      23593: inst = 32'hc404d11;
      23594: inst = 32'h8220000;
      23595: inst = 32'h10408000;
      23596: inst = 32'hc404d52;
      23597: inst = 32'h8220000;
      23598: inst = 32'h10408000;
      23599: inst = 32'hc404d71;
      23600: inst = 32'h8220000;
      23601: inst = 32'h10408000;
      23602: inst = 32'hc404db2;
      23603: inst = 32'h8220000;
      23604: inst = 32'h10408000;
      23605: inst = 32'hc404dd1;
      23606: inst = 32'h8220000;
      23607: inst = 32'h10408000;
      23608: inst = 32'hc404e12;
      23609: inst = 32'h8220000;
      23610: inst = 32'h10408000;
      23611: inst = 32'hc404e2d;
      23612: inst = 32'h8220000;
      23613: inst = 32'h10408000;
      23614: inst = 32'hc404e34;
      23615: inst = 32'h8220000;
      23616: inst = 32'h10408000;
      23617: inst = 32'hc404e37;
      23618: inst = 32'h8220000;
      23619: inst = 32'h10408000;
      23620: inst = 32'hc404e39;
      23621: inst = 32'h8220000;
      23622: inst = 32'h10408000;
      23623: inst = 32'hc404e3b;
      23624: inst = 32'h8220000;
      23625: inst = 32'h10408000;
      23626: inst = 32'hc404e3d;
      23627: inst = 32'h8220000;
      23628: inst = 32'h10408000;
      23629: inst = 32'hc404e42;
      23630: inst = 32'h8220000;
      23631: inst = 32'h10408000;
      23632: inst = 32'hc404e4c;
      23633: inst = 32'h8220000;
      23634: inst = 32'h10408000;
      23635: inst = 32'hc404e50;
      23636: inst = 32'h8220000;
      23637: inst = 32'h10408000;
      23638: inst = 32'hc404e5a;
      23639: inst = 32'h8220000;
      23640: inst = 32'h10408000;
      23641: inst = 32'hc404e60;
      23642: inst = 32'h8220000;
      23643: inst = 32'h10408000;
      23644: inst = 32'hc404e65;
      23645: inst = 32'h8220000;
      23646: inst = 32'h10408000;
      23647: inst = 32'hc404e69;
      23648: inst = 32'h8220000;
      23649: inst = 32'h10408000;
      23650: inst = 32'hc404e6e;
      23651: inst = 32'h8220000;
      23652: inst = 32'h10408000;
      23653: inst = 32'hc404e70;
      23654: inst = 32'h8220000;
      23655: inst = 32'h10408000;
      23656: inst = 32'hc404e72;
      23657: inst = 32'h8220000;
      23658: inst = 32'h10408000;
      23659: inst = 32'hc404e75;
      23660: inst = 32'h8220000;
      23661: inst = 32'h10408000;
      23662: inst = 32'hc404e8b;
      23663: inst = 32'h8220000;
      23664: inst = 32'h10408000;
      23665: inst = 32'hc404e8c;
      23666: inst = 32'h8220000;
      23667: inst = 32'h10408000;
      23668: inst = 32'hc404e91;
      23669: inst = 32'h8220000;
      23670: inst = 32'h10408000;
      23671: inst = 32'hc404e9b;
      23672: inst = 32'h8220000;
      23673: inst = 32'h10408000;
      23674: inst = 32'hc404ea0;
      23675: inst = 32'h8220000;
      23676: inst = 32'h10408000;
      23677: inst = 32'hc404eaa;
      23678: inst = 32'h8220000;
      23679: inst = 32'h10408000;
      23680: inst = 32'hc404ebb;
      23681: inst = 32'h8220000;
      23682: inst = 32'h10408000;
      23683: inst = 32'hc404ebe;
      23684: inst = 32'h8220000;
      23685: inst = 32'h10408000;
      23686: inst = 32'hc404ec3;
      23687: inst = 32'h8220000;
      23688: inst = 32'h10408000;
      23689: inst = 32'hc404eca;
      23690: inst = 32'h8220000;
      23691: inst = 32'h10408000;
      23692: inst = 32'hc404ecd;
      23693: inst = 32'h8220000;
      23694: inst = 32'h10408000;
      23695: inst = 32'hc404ed2;
      23696: inst = 32'h8220000;
      23697: inst = 32'h10408000;
      23698: inst = 32'hc404ed3;
      23699: inst = 32'h8220000;
      23700: inst = 32'h10408000;
      23701: inst = 32'hc404ed4;
      23702: inst = 32'h8220000;
      23703: inst = 32'h10408000;
      23704: inst = 32'hc404ef1;
      23705: inst = 32'h8220000;
      23706: inst = 32'h10408000;
      23707: inst = 32'hc404efb;
      23708: inst = 32'h8220000;
      23709: inst = 32'h10408000;
      23710: inst = 32'hc404f00;
      23711: inst = 32'h8220000;
      23712: inst = 32'h10408000;
      23713: inst = 32'hc404f0a;
      23714: inst = 32'h8220000;
      23715: inst = 32'h10408000;
      23716: inst = 32'hc404f1e;
      23717: inst = 32'h8220000;
      23718: inst = 32'h10408000;
      23719: inst = 32'hc404f23;
      23720: inst = 32'h8220000;
      23721: inst = 32'h10408000;
      23722: inst = 32'hc404f4d;
      23723: inst = 32'h8220000;
      23724: inst = 32'h10408000;
      23725: inst = 32'hc404f51;
      23726: inst = 32'h8220000;
      23727: inst = 32'h10408000;
      23728: inst = 32'hc404f5b;
      23729: inst = 32'h8220000;
      23730: inst = 32'h10408000;
      23731: inst = 32'hc404f60;
      23732: inst = 32'h8220000;
      23733: inst = 32'h10408000;
      23734: inst = 32'hc404f6a;
      23735: inst = 32'h8220000;
      23736: inst = 32'h10408000;
      23737: inst = 32'hc404f7b;
      23738: inst = 32'h8220000;
      23739: inst = 32'h10408000;
      23740: inst = 32'hc404f7e;
      23741: inst = 32'h8220000;
      23742: inst = 32'h10408000;
      23743: inst = 32'hc404f83;
      23744: inst = 32'h8220000;
      23745: inst = 32'h10408000;
      23746: inst = 32'hc404f8a;
      23747: inst = 32'h8220000;
      23748: inst = 32'h10408000;
      23749: inst = 32'hc404f93;
      23750: inst = 32'h8220000;
      23751: inst = 32'h10408000;
      23752: inst = 32'hc404fb1;
      23753: inst = 32'h8220000;
      23754: inst = 32'h10408000;
      23755: inst = 32'hc404fbb;
      23756: inst = 32'h8220000;
      23757: inst = 32'h10408000;
      23758: inst = 32'hc404fbd;
      23759: inst = 32'h8220000;
      23760: inst = 32'h10408000;
      23761: inst = 32'hc404fc0;
      23762: inst = 32'h8220000;
      23763: inst = 32'h10408000;
      23764: inst = 32'hc404fca;
      23765: inst = 32'h8220000;
      23766: inst = 32'h10408000;
      23767: inst = 32'hc404fdb;
      23768: inst = 32'h8220000;
      23769: inst = 32'h10408000;
      23770: inst = 32'hc404fde;
      23771: inst = 32'h8220000;
      23772: inst = 32'h10408000;
      23773: inst = 32'hc404fe3;
      23774: inst = 32'h8220000;
      23775: inst = 32'h10408000;
      23776: inst = 32'hc404fea;
      23777: inst = 32'h8220000;
      23778: inst = 32'h10408000;
      23779: inst = 32'hc404ff2;
      23780: inst = 32'h8220000;
      23781: inst = 32'h10408000;
      23782: inst = 32'hc40500d;
      23783: inst = 32'h8220000;
      23784: inst = 32'h10408000;
      23785: inst = 32'hc40500f;
      23786: inst = 32'h8220000;
      23787: inst = 32'h10408000;
      23788: inst = 32'hc405013;
      23789: inst = 32'h8220000;
      23790: inst = 32'h10408000;
      23791: inst = 32'hc405017;
      23792: inst = 32'h8220000;
      23793: inst = 32'h10408000;
      23794: inst = 32'hc405023;
      23795: inst = 32'h8220000;
      23796: inst = 32'h10408000;
      23797: inst = 32'hc40502d;
      23798: inst = 32'h8220000;
      23799: inst = 32'h10408000;
      23800: inst = 32'hc405030;
      23801: inst = 32'h8220000;
      23802: inst = 32'h10408000;
      23803: inst = 32'hc40503a;
      23804: inst = 32'h8220000;
      23805: inst = 32'h10408000;
      23806: inst = 32'hc40503d;
      23807: inst = 32'h8220000;
      23808: inst = 32'h10408000;
      23809: inst = 32'hc405041;
      23810: inst = 32'h8220000;
      23811: inst = 32'h10408000;
      23812: inst = 32'hc405046;
      23813: inst = 32'h8220000;
      23814: inst = 32'h10408000;
      23815: inst = 32'hc405049;
      23816: inst = 32'h8220000;
      23817: inst = 32'h10408000;
      23818: inst = 32'hc40504c;
      23819: inst = 32'h8220000;
      23820: inst = 32'h10408000;
      23821: inst = 32'hc40504e;
      23822: inst = 32'h8220000;
      23823: inst = 32'hc20f7be;
      23824: inst = 32'h10408000;
      23825: inst = 32'hc4046af;
      23826: inst = 32'h8220000;
      23827: inst = 32'h10408000;
      23828: inst = 32'hc4046f2;
      23829: inst = 32'h8220000;
      23830: inst = 32'h10408000;
      23831: inst = 32'hc40470f;
      23832: inst = 32'h8220000;
      23833: inst = 32'h10408000;
      23834: inst = 32'hc404752;
      23835: inst = 32'h8220000;
      23836: inst = 32'h10408000;
      23837: inst = 32'hc40476f;
      23838: inst = 32'h8220000;
      23839: inst = 32'h10408000;
      23840: inst = 32'hc4047b2;
      23841: inst = 32'h8220000;
      23842: inst = 32'h10408000;
      23843: inst = 32'hc4047cf;
      23844: inst = 32'h8220000;
      23845: inst = 32'h10408000;
      23846: inst = 32'hc4047d9;
      23847: inst = 32'h8220000;
      23848: inst = 32'h10408000;
      23849: inst = 32'hc4047fc;
      23850: inst = 32'h8220000;
      23851: inst = 32'h10408000;
      23852: inst = 32'hc404807;
      23853: inst = 32'h8220000;
      23854: inst = 32'h10408000;
      23855: inst = 32'hc40480a;
      23856: inst = 32'h8220000;
      23857: inst = 32'h10408000;
      23858: inst = 32'hc404812;
      23859: inst = 32'h8220000;
      23860: inst = 32'h10408000;
      23861: inst = 32'hc40482f;
      23862: inst = 32'h8220000;
      23863: inst = 32'h10408000;
      23864: inst = 32'hc404839;
      23865: inst = 32'h8220000;
      23866: inst = 32'h10408000;
      23867: inst = 32'hc40485c;
      23868: inst = 32'h8220000;
      23869: inst = 32'h10408000;
      23870: inst = 32'hc404867;
      23871: inst = 32'h8220000;
      23872: inst = 32'h10408000;
      23873: inst = 32'hc404872;
      23874: inst = 32'h8220000;
      23875: inst = 32'h10408000;
      23876: inst = 32'hc40488f;
      23877: inst = 32'h8220000;
      23878: inst = 32'h10408000;
      23879: inst = 32'hc404893;
      23880: inst = 32'h8220000;
      23881: inst = 32'h10408000;
      23882: inst = 32'hc404899;
      23883: inst = 32'h8220000;
      23884: inst = 32'h10408000;
      23885: inst = 32'hc4048ac;
      23886: inst = 32'h8220000;
      23887: inst = 32'h10408000;
      23888: inst = 32'hc4048b2;
      23889: inst = 32'h8220000;
      23890: inst = 32'h10408000;
      23891: inst = 32'hc4048bb;
      23892: inst = 32'h8220000;
      23893: inst = 32'h10408000;
      23894: inst = 32'hc4048bc;
      23895: inst = 32'h8220000;
      23896: inst = 32'h10408000;
      23897: inst = 32'hc4048c7;
      23898: inst = 32'h8220000;
      23899: inst = 32'h10408000;
      23900: inst = 32'hc4048cf;
      23901: inst = 32'h8220000;
      23902: inst = 32'h10408000;
      23903: inst = 32'hc4048d2;
      23904: inst = 32'h8220000;
      23905: inst = 32'h10408000;
      23906: inst = 32'hc4048ef;
      23907: inst = 32'h8220000;
      23908: inst = 32'h10408000;
      23909: inst = 32'hc4048f3;
      23910: inst = 32'h8220000;
      23911: inst = 32'h10408000;
      23912: inst = 32'hc4048f9;
      23913: inst = 32'h8220000;
      23914: inst = 32'h10408000;
      23915: inst = 32'hc40490c;
      23916: inst = 32'h8220000;
      23917: inst = 32'h10408000;
      23918: inst = 32'hc404912;
      23919: inst = 32'h8220000;
      23920: inst = 32'h10408000;
      23921: inst = 32'hc40491b;
      23922: inst = 32'h8220000;
      23923: inst = 32'h10408000;
      23924: inst = 32'hc40491c;
      23925: inst = 32'h8220000;
      23926: inst = 32'h10408000;
      23927: inst = 32'hc404927;
      23928: inst = 32'h8220000;
      23929: inst = 32'h10408000;
      23930: inst = 32'hc40492f;
      23931: inst = 32'h8220000;
      23932: inst = 32'h10408000;
      23933: inst = 32'hc404932;
      23934: inst = 32'h8220000;
      23935: inst = 32'h10408000;
      23936: inst = 32'hc40494f;
      23937: inst = 32'h8220000;
      23938: inst = 32'h10408000;
      23939: inst = 32'hc404959;
      23940: inst = 32'h8220000;
      23941: inst = 32'h10408000;
      23942: inst = 32'hc404972;
      23943: inst = 32'h8220000;
      23944: inst = 32'h10408000;
      23945: inst = 32'hc40497c;
      23946: inst = 32'h8220000;
      23947: inst = 32'h10408000;
      23948: inst = 32'hc404987;
      23949: inst = 32'h8220000;
      23950: inst = 32'h10408000;
      23951: inst = 32'hc404992;
      23952: inst = 32'h8220000;
      23953: inst = 32'h10408000;
      23954: inst = 32'hc4049b9;
      23955: inst = 32'h8220000;
      23956: inst = 32'h10408000;
      23957: inst = 32'hc4049dc;
      23958: inst = 32'h8220000;
      23959: inst = 32'h10408000;
      23960: inst = 32'hc4049e7;
      23961: inst = 32'h8220000;
      23962: inst = 32'h10408000;
      23963: inst = 32'hc4049f2;
      23964: inst = 32'h8220000;
      23965: inst = 32'h10408000;
      23966: inst = 32'hc404e74;
      23967: inst = 32'h8220000;
      23968: inst = 32'h10408000;
      23969: inst = 32'hc404ef4;
      23970: inst = 32'h8220000;
      23971: inst = 32'h10408000;
      23972: inst = 32'hc404ef5;
      23973: inst = 32'h8220000;
      23974: inst = 32'h10408000;
      23975: inst = 32'hc404ef9;
      23976: inst = 32'h8220000;
      23977: inst = 32'h10408000;
      23978: inst = 32'hc404f0e;
      23979: inst = 32'h8220000;
      23980: inst = 32'h10408000;
      23981: inst = 32'hc404f12;
      23982: inst = 32'h8220000;
      23983: inst = 32'h10408000;
      23984: inst = 32'hc404f2c;
      23985: inst = 32'h8220000;
      23986: inst = 32'h10408000;
      23987: inst = 32'hc404f33;
      23988: inst = 32'h8220000;
      23989: inst = 32'h10408000;
      23990: inst = 32'hc404f54;
      23991: inst = 32'h8220000;
      23992: inst = 32'h10408000;
      23993: inst = 32'hc404f59;
      23994: inst = 32'h8220000;
      23995: inst = 32'h10408000;
      23996: inst = 32'hc404f72;
      23997: inst = 32'h8220000;
      23998: inst = 32'h10408000;
      23999: inst = 32'hc404f8c;
      24000: inst = 32'h8220000;
      24001: inst = 32'h10408000;
      24002: inst = 32'hc404fb4;
      24003: inst = 32'h8220000;
      24004: inst = 32'h10408000;
      24005: inst = 32'hc404fb9;
      24006: inst = 32'h8220000;
      24007: inst = 32'h10408000;
      24008: inst = 32'hc404fd2;
      24009: inst = 32'h8220000;
      24010: inst = 32'h10408000;
      24011: inst = 32'hc404fd8;
      24012: inst = 32'h8220000;
      24013: inst = 32'h10408000;
      24014: inst = 32'hc404fe7;
      24015: inst = 32'h8220000;
      24016: inst = 32'h10408000;
      24017: inst = 32'hc405014;
      24018: inst = 32'h8220000;
      24019: inst = 32'hc205acb;
      24020: inst = 32'h10408000;
      24021: inst = 32'hc4046b0;
      24022: inst = 32'h8220000;
      24023: inst = 32'h10408000;
      24024: inst = 32'hc404710;
      24025: inst = 32'h8220000;
      24026: inst = 32'h10408000;
      24027: inst = 32'hc404751;
      24028: inst = 32'h8220000;
      24029: inst = 32'h10408000;
      24030: inst = 32'hc404770;
      24031: inst = 32'h8220000;
      24032: inst = 32'h10408000;
      24033: inst = 32'hc404771;
      24034: inst = 32'h8220000;
      24035: inst = 32'h10408000;
      24036: inst = 32'hc404774;
      24037: inst = 32'h8220000;
      24038: inst = 32'h10408000;
      24039: inst = 32'hc404777;
      24040: inst = 32'h8220000;
      24041: inst = 32'h10408000;
      24042: inst = 32'hc40477b;
      24043: inst = 32'h8220000;
      24044: inst = 32'h10408000;
      24045: inst = 32'hc404783;
      24046: inst = 32'h8220000;
      24047: inst = 32'h10408000;
      24048: inst = 32'hc404786;
      24049: inst = 32'h8220000;
      24050: inst = 32'h10408000;
      24051: inst = 32'hc40478a;
      24052: inst = 32'h8220000;
      24053: inst = 32'h10408000;
      24054: inst = 32'hc404794;
      24055: inst = 32'h8220000;
      24056: inst = 32'h10408000;
      24057: inst = 32'hc404799;
      24058: inst = 32'h8220000;
      24059: inst = 32'h10408000;
      24060: inst = 32'hc40479e;
      24061: inst = 32'h8220000;
      24062: inst = 32'h10408000;
      24063: inst = 32'hc4047a1;
      24064: inst = 32'h8220000;
      24065: inst = 32'h10408000;
      24066: inst = 32'hc4047a4;
      24067: inst = 32'h8220000;
      24068: inst = 32'h10408000;
      24069: inst = 32'hc4047a6;
      24070: inst = 32'h8220000;
      24071: inst = 32'h10408000;
      24072: inst = 32'hc4047a9;
      24073: inst = 32'h8220000;
      24074: inst = 32'h10408000;
      24075: inst = 32'hc4047ad;
      24076: inst = 32'h8220000;
      24077: inst = 32'h10408000;
      24078: inst = 32'hc4047b1;
      24079: inst = 32'h8220000;
      24080: inst = 32'h10408000;
      24081: inst = 32'hc4047f6;
      24082: inst = 32'h8220000;
      24083: inst = 32'h10408000;
      24084: inst = 32'hc404811;
      24085: inst = 32'h8220000;
      24086: inst = 32'h10408000;
      24087: inst = 32'hc404853;
      24088: inst = 32'h8220000;
      24089: inst = 32'h10408000;
      24090: inst = 32'hc404866;
      24091: inst = 32'h8220000;
      24092: inst = 32'h10408000;
      24093: inst = 32'hc404871;
      24094: inst = 32'h8220000;
      24095: inst = 32'h10408000;
      24096: inst = 32'hc404890;
      24097: inst = 32'h8220000;
      24098: inst = 32'h10408000;
      24099: inst = 32'hc404892;
      24100: inst = 32'h8220000;
      24101: inst = 32'h10408000;
      24102: inst = 32'hc40489a;
      24103: inst = 32'h8220000;
      24104: inst = 32'h10408000;
      24105: inst = 32'hc4048ab;
      24106: inst = 32'h8220000;
      24107: inst = 32'h10408000;
      24108: inst = 32'hc4048b1;
      24109: inst = 32'h8220000;
      24110: inst = 32'h10408000;
      24111: inst = 32'hc4048ba;
      24112: inst = 32'h8220000;
      24113: inst = 32'h10408000;
      24114: inst = 32'hc4048bd;
      24115: inst = 32'h8220000;
      24116: inst = 32'h10408000;
      24117: inst = 32'hc4048c6;
      24118: inst = 32'h8220000;
      24119: inst = 32'h10408000;
      24120: inst = 32'hc4048ce;
      24121: inst = 32'h8220000;
      24122: inst = 32'h10408000;
      24123: inst = 32'hc4048d1;
      24124: inst = 32'h8220000;
      24125: inst = 32'h10408000;
      24126: inst = 32'hc4048f0;
      24127: inst = 32'h8220000;
      24128: inst = 32'h10408000;
      24129: inst = 32'hc4048f2;
      24130: inst = 32'h8220000;
      24131: inst = 32'h10408000;
      24132: inst = 32'hc4048fa;
      24133: inst = 32'h8220000;
      24134: inst = 32'h10408000;
      24135: inst = 32'hc40490b;
      24136: inst = 32'h8220000;
      24137: inst = 32'h10408000;
      24138: inst = 32'hc404911;
      24139: inst = 32'h8220000;
      24140: inst = 32'h10408000;
      24141: inst = 32'hc40491a;
      24142: inst = 32'h8220000;
      24143: inst = 32'h10408000;
      24144: inst = 32'hc40491d;
      24145: inst = 32'h8220000;
      24146: inst = 32'h10408000;
      24147: inst = 32'hc404926;
      24148: inst = 32'h8220000;
      24149: inst = 32'h10408000;
      24150: inst = 32'hc40492e;
      24151: inst = 32'h8220000;
      24152: inst = 32'h10408000;
      24153: inst = 32'hc404931;
      24154: inst = 32'h8220000;
      24155: inst = 32'h10408000;
      24156: inst = 32'hc404950;
      24157: inst = 32'h8220000;
      24158: inst = 32'h10408000;
      24159: inst = 32'hc40495a;
      24160: inst = 32'h8220000;
      24161: inst = 32'h10408000;
      24162: inst = 32'hc40497d;
      24163: inst = 32'h8220000;
      24164: inst = 32'h10408000;
      24165: inst = 32'hc404986;
      24166: inst = 32'h8220000;
      24167: inst = 32'h10408000;
      24168: inst = 32'hc404991;
      24169: inst = 32'h8220000;
      24170: inst = 32'h10408000;
      24171: inst = 32'hc404a11;
      24172: inst = 32'h8220000;
      24173: inst = 32'h10408000;
      24174: inst = 32'hc404a19;
      24175: inst = 32'h8220000;
      24176: inst = 32'h10408000;
      24177: inst = 32'hc404a1c;
      24178: inst = 32'h8220000;
      24179: inst = 32'h10408000;
      24180: inst = 32'hc404a1d;
      24181: inst = 32'h8220000;
      24182: inst = 32'h10408000;
      24183: inst = 32'hc404a2a;
      24184: inst = 32'h8220000;
      24185: inst = 32'h10408000;
      24186: inst = 32'hc404a34;
      24187: inst = 32'h8220000;
      24188: inst = 32'h10408000;
      24189: inst = 32'hc404a39;
      24190: inst = 32'h8220000;
      24191: inst = 32'h10408000;
      24192: inst = 32'hc404a3c;
      24193: inst = 32'h8220000;
      24194: inst = 32'h10408000;
      24195: inst = 32'hc404a3f;
      24196: inst = 32'h8220000;
      24197: inst = 32'h10408000;
      24198: inst = 32'hc404a40;
      24199: inst = 32'h8220000;
      24200: inst = 32'h10408000;
      24201: inst = 32'hc404a46;
      24202: inst = 32'h8220000;
      24203: inst = 32'h10408000;
      24204: inst = 32'hc404a47;
      24205: inst = 32'h8220000;
      24206: inst = 32'h10408000;
      24207: inst = 32'hc404a48;
      24208: inst = 32'h8220000;
      24209: inst = 32'h10408000;
      24210: inst = 32'hc404a4d;
      24211: inst = 32'h8220000;
      24212: inst = 32'h10408000;
      24213: inst = 32'hc404a51;
      24214: inst = 32'h8220000;
      24215: inst = 32'h10408000;
      24216: inst = 32'hc404a52;
      24217: inst = 32'h8220000;
      24218: inst = 32'h10408000;
      24219: inst = 32'hc404a53;
      24220: inst = 32'h8220000;
      24221: inst = 32'h10408000;
      24222: inst = 32'hc404d80;
      24223: inst = 32'h8220000;
      24224: inst = 32'h10408000;
      24225: inst = 32'hc404d8a;
      24226: inst = 32'h8220000;
      24227: inst = 32'h10408000;
      24228: inst = 32'hc404d9e;
      24229: inst = 32'h8220000;
      24230: inst = 32'h10408000;
      24231: inst = 32'hc404da3;
      24232: inst = 32'h8220000;
      24233: inst = 32'h10408000;
      24234: inst = 32'hc404dcd;
      24235: inst = 32'h8220000;
      24236: inst = 32'h10408000;
      24237: inst = 32'hc404dd2;
      24238: inst = 32'h8220000;
      24239: inst = 32'h10408000;
      24240: inst = 32'hc404dd3;
      24241: inst = 32'h8220000;
      24242: inst = 32'h10408000;
      24243: inst = 32'hc404dd7;
      24244: inst = 32'h8220000;
      24245: inst = 32'h10408000;
      24246: inst = 32'hc404dde;
      24247: inst = 32'h8220000;
      24248: inst = 32'h10408000;
      24249: inst = 32'hc404de2;
      24250: inst = 32'h8220000;
      24251: inst = 32'h10408000;
      24252: inst = 32'hc404dec;
      24253: inst = 32'h8220000;
      24254: inst = 32'h10408000;
      24255: inst = 32'hc404df0;
      24256: inst = 32'h8220000;
      24257: inst = 32'h10408000;
      24258: inst = 32'hc404dfa;
      24259: inst = 32'h8220000;
      24260: inst = 32'h10408000;
      24261: inst = 32'hc404e00;
      24262: inst = 32'h8220000;
      24263: inst = 32'h10408000;
      24264: inst = 32'hc404e05;
      24265: inst = 32'h8220000;
      24266: inst = 32'h10408000;
      24267: inst = 32'hc404e09;
      24268: inst = 32'h8220000;
      24269: inst = 32'h10408000;
      24270: inst = 32'hc404e0e;
      24271: inst = 32'h8220000;
      24272: inst = 32'h10408000;
      24273: inst = 32'hc404e14;
      24274: inst = 32'h8220000;
      24275: inst = 32'h10408000;
      24276: inst = 32'hc404e15;
      24277: inst = 32'h8220000;
      24278: inst = 32'h10408000;
      24279: inst = 32'hc404e93;
      24280: inst = 32'h8220000;
      24281: inst = 32'h10408000;
      24282: inst = 32'hc404e9d;
      24283: inst = 32'h8220000;
      24284: inst = 32'h10408000;
      24285: inst = 32'hc404eb9;
      24286: inst = 32'h8220000;
      24287: inst = 32'h10408000;
      24288: inst = 32'hc404ec8;
      24289: inst = 32'h8220000;
      24290: inst = 32'h10408000;
      24291: inst = 32'hc404ef3;
      24292: inst = 32'h8220000;
      24293: inst = 32'h10408000;
      24294: inst = 32'hc404efd;
      24295: inst = 32'h8220000;
      24296: inst = 32'h10408000;
      24297: inst = 32'hc404f13;
      24298: inst = 32'h8220000;
      24299: inst = 32'h10408000;
      24300: inst = 32'hc404f2d;
      24301: inst = 32'h8220000;
      24302: inst = 32'h10408000;
      24303: inst = 32'hc404f53;
      24304: inst = 32'h8220000;
      24305: inst = 32'h10408000;
      24306: inst = 32'hc404f5d;
      24307: inst = 32'h8220000;
      24308: inst = 32'h10408000;
      24309: inst = 32'hc404f73;
      24310: inst = 32'h8220000;
      24311: inst = 32'h10408000;
      24312: inst = 32'hc404f8d;
      24313: inst = 32'h8220000;
      24314: inst = 32'h10408000;
      24315: inst = 32'hc404fb3;
      24316: inst = 32'h8220000;
      24317: inst = 32'h10408000;
      24318: inst = 32'hc404fd7;
      24319: inst = 32'h8220000;
      24320: inst = 32'h10408000;
      24321: inst = 32'hc404fdd;
      24322: inst = 32'h8220000;
      24323: inst = 32'h10408000;
      24324: inst = 32'hc405020;
      24325: inst = 32'h8220000;
      24326: inst = 32'h10408000;
      24327: inst = 32'hc40502a;
      24328: inst = 32'h8220000;
      24329: inst = 32'h10408000;
      24330: inst = 32'hc40503e;
      24331: inst = 32'h8220000;
      24332: inst = 32'h10408000;
      24333: inst = 32'hc405043;
      24334: inst = 32'h8220000;
      24335: inst = 32'h10408000;
      24336: inst = 32'hc40506d;
      24337: inst = 32'h8220000;
      24338: inst = 32'h10408000;
      24339: inst = 32'hc405070;
      24340: inst = 32'h8220000;
      24341: inst = 32'h10408000;
      24342: inst = 32'hc405071;
      24343: inst = 32'h8220000;
      24344: inst = 32'h10408000;
      24345: inst = 32'hc405074;
      24346: inst = 32'h8220000;
      24347: inst = 32'h10408000;
      24348: inst = 32'hc405077;
      24349: inst = 32'h8220000;
      24350: inst = 32'h10408000;
      24351: inst = 32'hc40507c;
      24352: inst = 32'h8220000;
      24353: inst = 32'h10408000;
      24354: inst = 32'hc405082;
      24355: inst = 32'h8220000;
      24356: inst = 32'h10408000;
      24357: inst = 32'hc40508c;
      24358: inst = 32'h8220000;
      24359: inst = 32'h10408000;
      24360: inst = 32'hc405090;
      24361: inst = 32'h8220000;
      24362: inst = 32'h10408000;
      24363: inst = 32'hc405099;
      24364: inst = 32'h8220000;
      24365: inst = 32'h10408000;
      24366: inst = 32'hc40509c;
      24367: inst = 32'h8220000;
      24368: inst = 32'h10408000;
      24369: inst = 32'hc4050a0;
      24370: inst = 32'h8220000;
      24371: inst = 32'h10408000;
      24372: inst = 32'hc4050a5;
      24373: inst = 32'h8220000;
      24374: inst = 32'h10408000;
      24375: inst = 32'hc4050a8;
      24376: inst = 32'h8220000;
      24377: inst = 32'h10408000;
      24378: inst = 32'hc4050ab;
      24379: inst = 32'h8220000;
      24380: inst = 32'h10408000;
      24381: inst = 32'hc4050ae;
      24382: inst = 32'h8220000;
      24383: inst = 32'h10408000;
      24384: inst = 32'hc4050b1;
      24385: inst = 32'h8220000;
      24386: inst = 32'h10408000;
      24387: inst = 32'hc4050b2;
      24388: inst = 32'h8220000;
      24389: inst = 32'h10408000;
      24390: inst = 32'hc4050b5;
      24391: inst = 32'h8220000;
      24392: inst = 32'hc20defb;
      24393: inst = 32'h10408000;
      24394: inst = 32'hc404775;
      24395: inst = 32'h8220000;
      24396: inst = 32'h10408000;
      24397: inst = 32'hc404784;
      24398: inst = 32'h8220000;
      24399: inst = 32'h10408000;
      24400: inst = 32'hc4047a2;
      24401: inst = 32'h8220000;
      24402: inst = 32'h10408000;
      24403: inst = 32'hc4047d2;
      24404: inst = 32'h8220000;
      24405: inst = 32'h10408000;
      24406: inst = 32'hc4047d5;
      24407: inst = 32'h8220000;
      24408: inst = 32'h10408000;
      24409: inst = 32'hc4047e4;
      24410: inst = 32'h8220000;
      24411: inst = 32'h10408000;
      24412: inst = 32'hc4047eb;
      24413: inst = 32'h8220000;
      24414: inst = 32'h10408000;
      24415: inst = 32'hc4047fa;
      24416: inst = 32'h8220000;
      24417: inst = 32'h10408000;
      24418: inst = 32'hc404802;
      24419: inst = 32'h8220000;
      24420: inst = 32'h10408000;
      24421: inst = 32'hc40480e;
      24422: inst = 32'h8220000;
      24423: inst = 32'h10408000;
      24424: inst = 32'hc404833;
      24425: inst = 32'h8220000;
      24426: inst = 32'h10408000;
      24427: inst = 32'hc40496c;
      24428: inst = 32'h8220000;
      24429: inst = 32'h10408000;
      24430: inst = 32'hc40497b;
      24431: inst = 32'h8220000;
      24432: inst = 32'h10408000;
      24433: inst = 32'hc40498f;
      24434: inst = 32'h8220000;
      24435: inst = 32'h10408000;
      24436: inst = 32'hc4049af;
      24437: inst = 32'h8220000;
      24438: inst = 32'h10408000;
      24439: inst = 32'hc4049b6;
      24440: inst = 32'h8220000;
      24441: inst = 32'h10408000;
      24442: inst = 32'hc4049bd;
      24443: inst = 32'h8220000;
      24444: inst = 32'h10408000;
      24445: inst = 32'hc4049c5;
      24446: inst = 32'h8220000;
      24447: inst = 32'h10408000;
      24448: inst = 32'hc4049d3;
      24449: inst = 32'h8220000;
      24450: inst = 32'h10408000;
      24451: inst = 32'hc4049e0;
      24452: inst = 32'h8220000;
      24453: inst = 32'h10408000;
      24454: inst = 32'hc4049e3;
      24455: inst = 32'h8220000;
      24456: inst = 32'h10408000;
      24457: inst = 32'hc404d10;
      24458: inst = 32'h8220000;
      24459: inst = 32'h10408000;
      24460: inst = 32'hc404d51;
      24461: inst = 32'h8220000;
      24462: inst = 32'h10408000;
      24463: inst = 32'hc404e31;
      24464: inst = 32'h8220000;
      24465: inst = 32'h10408000;
      24466: inst = 32'hc404e3a;
      24467: inst = 32'h8220000;
      24468: inst = 32'h10408000;
      24469: inst = 32'hc404e41;
      24470: inst = 32'h8220000;
      24471: inst = 32'h10408000;
      24472: inst = 32'hc404e4b;
      24473: inst = 32'h8220000;
      24474: inst = 32'h10408000;
      24475: inst = 32'hc404e5f;
      24476: inst = 32'h8220000;
      24477: inst = 32'h10408000;
      24478: inst = 32'hc404e64;
      24479: inst = 32'h8220000;
      24480: inst = 32'h10408000;
      24481: inst = 32'hc404e94;
      24482: inst = 32'h8220000;
      24483: inst = 32'h10408000;
      24484: inst = 32'hc404e95;
      24485: inst = 32'h8220000;
      24486: inst = 32'h10408000;
      24487: inst = 32'hc404e99;
      24488: inst = 32'h8220000;
      24489: inst = 32'h10408000;
      24490: inst = 32'hc404eae;
      24491: inst = 32'h8220000;
      24492: inst = 32'h10408000;
      24493: inst = 32'hc404eb2;
      24494: inst = 32'h8220000;
      24495: inst = 32'h10408000;
      24496: inst = 32'hc404f4e;
      24497: inst = 32'h8220000;
      24498: inst = 32'h10408000;
      24499: inst = 32'hc404fb5;
      24500: inst = 32'h8220000;
      24501: inst = 32'h10408000;
      24502: inst = 32'hc404fce;
      24503: inst = 32'h8220000;
      24504: inst = 32'h10408000;
      24505: inst = 32'hc405010;
      24506: inst = 32'h8220000;
      24507: inst = 32'h10408000;
      24508: inst = 32'hc40504d;
      24509: inst = 32'h8220000;
      24510: inst = 32'h10408000;
      24511: inst = 32'hc405051;
      24512: inst = 32'h8220000;
      24513: inst = 32'hc207bef;
      24514: inst = 32'h10408000;
      24515: inst = 32'hc404779;
      24516: inst = 32'h8220000;
      24517: inst = 32'h10408000;
      24518: inst = 32'hc40479c;
      24519: inst = 32'h8220000;
      24520: inst = 32'h10408000;
      24521: inst = 32'hc4047e8;
      24522: inst = 32'h8220000;
      24523: inst = 32'h10408000;
      24524: inst = 32'hc4047f2;
      24525: inst = 32'h8220000;
      24526: inst = 32'h10408000;
      24527: inst = 32'hc4047f7;
      24528: inst = 32'h8220000;
      24529: inst = 32'h10408000;
      24530: inst = 32'hc40480b;
      24531: inst = 32'h8220000;
      24532: inst = 32'h10408000;
      24533: inst = 32'hc404830;
      24534: inst = 32'h8220000;
      24535: inst = 32'h10408000;
      24536: inst = 32'hc40484b;
      24537: inst = 32'h8220000;
      24538: inst = 32'h10408000;
      24539: inst = 32'hc40485a;
      24540: inst = 32'h8220000;
      24541: inst = 32'h10408000;
      24542: inst = 32'hc40486e;
      24543: inst = 32'h8220000;
      24544: inst = 32'h10408000;
      24545: inst = 32'hc40496b;
      24546: inst = 32'h8220000;
      24547: inst = 32'h10408000;
      24548: inst = 32'hc40497a;
      24549: inst = 32'h8220000;
      24550: inst = 32'h10408000;
      24551: inst = 32'hc40498e;
      24552: inst = 32'h8220000;
      24553: inst = 32'h10408000;
      24554: inst = 32'hc4049c8;
      24555: inst = 32'h8220000;
      24556: inst = 32'h10408000;
      24557: inst = 32'hc4049d2;
      24558: inst = 32'h8220000;
      24559: inst = 32'h10408000;
      24560: inst = 32'hc4049d7;
      24561: inst = 32'h8220000;
      24562: inst = 32'h10408000;
      24563: inst = 32'hc4049eb;
      24564: inst = 32'h8220000;
      24565: inst = 32'h10408000;
      24566: inst = 32'hc404e52;
      24567: inst = 32'h8220000;
      24568: inst = 32'h10408000;
      24569: inst = 32'hc404eee;
      24570: inst = 32'h8220000;
      24571: inst = 32'h10408000;
      24572: inst = 32'hc404ff5;
      24573: inst = 32'h8220000;
      24574: inst = 32'h10408000;
      24575: inst = 32'hc405019;
      24576: inst = 32'h8220000;
      24577: inst = 32'h10408000;
      24578: inst = 32'hc40501f;
      24579: inst = 32'h8220000;
      24580: inst = 32'h10408000;
      24581: inst = 32'hc405032;
      24582: inst = 32'h8220000;
      24583: inst = 32'h10408000;
      24584: inst = 32'hc405050;
      24585: inst = 32'h8220000;
      24586: inst = 32'hc204208;
      24587: inst = 32'h10408000;
      24588: inst = 32'hc40477c;
      24589: inst = 32'h8220000;
      24590: inst = 32'h10408000;
      24591: inst = 32'hc404789;
      24592: inst = 32'h8220000;
      24593: inst = 32'h10408000;
      24594: inst = 32'hc404798;
      24595: inst = 32'h8220000;
      24596: inst = 32'h10408000;
      24597: inst = 32'hc40479f;
      24598: inst = 32'h8220000;
      24599: inst = 32'h10408000;
      24600: inst = 32'hc4047aa;
      24601: inst = 32'h8220000;
      24602: inst = 32'h10408000;
      24603: inst = 32'hc4047ac;
      24604: inst = 32'h8220000;
      24605: inst = 32'h10408000;
      24606: inst = 32'hc4047d8;
      24607: inst = 32'h8220000;
      24608: inst = 32'h10408000;
      24609: inst = 32'hc4047ec;
      24610: inst = 32'h8220000;
      24611: inst = 32'h10408000;
      24612: inst = 32'hc4047fb;
      24613: inst = 32'h8220000;
      24614: inst = 32'h10408000;
      24615: inst = 32'hc404805;
      24616: inst = 32'h8220000;
      24617: inst = 32'h10408000;
      24618: inst = 32'hc40480f;
      24619: inst = 32'h8220000;
      24620: inst = 32'h10408000;
      24621: inst = 32'hc404973;
      24622: inst = 32'h8220000;
      24623: inst = 32'h10408000;
      24624: inst = 32'hc4049b3;
      24625: inst = 32'h8220000;
      24626: inst = 32'h10408000;
      24627: inst = 32'hc4049cc;
      24628: inst = 32'h8220000;
      24629: inst = 32'h10408000;
      24630: inst = 32'hc4049d6;
      24631: inst = 32'h8220000;
      24632: inst = 32'h10408000;
      24633: inst = 32'hc4049e9;
      24634: inst = 32'h8220000;
      24635: inst = 32'h10408000;
      24636: inst = 32'hc4049ef;
      24637: inst = 32'h8220000;
      24638: inst = 32'h10408000;
      24639: inst = 32'hc4049f4;
      24640: inst = 32'h8220000;
      24641: inst = 32'h10408000;
      24642: inst = 32'hc404a16;
      24643: inst = 32'h8220000;
      24644: inst = 32'h10408000;
      24645: inst = 32'hc404a17;
      24646: inst = 32'h8220000;
      24647: inst = 32'h10408000;
      24648: inst = 32'hc404a1a;
      24649: inst = 32'h8220000;
      24650: inst = 32'h10408000;
      24651: inst = 32'hc404a25;
      24652: inst = 32'h8220000;
      24653: inst = 32'h10408000;
      24654: inst = 32'hc404a26;
      24655: inst = 32'h8220000;
      24656: inst = 32'h10408000;
      24657: inst = 32'hc404a29;
      24658: inst = 32'h8220000;
      24659: inst = 32'h10408000;
      24660: inst = 32'hc404a33;
      24661: inst = 32'h8220000;
      24662: inst = 32'h10408000;
      24663: inst = 32'hc404a38;
      24664: inst = 32'h8220000;
      24665: inst = 32'h10408000;
      24666: inst = 32'hc404a3d;
      24667: inst = 32'h8220000;
      24668: inst = 32'h10408000;
      24669: inst = 32'hc404a43;
      24670: inst = 32'h8220000;
      24671: inst = 32'h10408000;
      24672: inst = 32'hc404a44;
      24673: inst = 32'h8220000;
      24674: inst = 32'h10408000;
      24675: inst = 32'hc404a4c;
      24676: inst = 32'h8220000;
      24677: inst = 32'h10408000;
      24678: inst = 32'hc404caf;
      24679: inst = 32'h8220000;
      24680: inst = 32'h10408000;
      24681: inst = 32'hc404cf0;
      24682: inst = 32'h8220000;
      24683: inst = 32'h10408000;
      24684: inst = 32'hc404d0f;
      24685: inst = 32'h8220000;
      24686: inst = 32'h10408000;
      24687: inst = 32'hc404d50;
      24688: inst = 32'h8220000;
      24689: inst = 32'h10408000;
      24690: inst = 32'hc404dce;
      24691: inst = 32'h8220000;
      24692: inst = 32'h10408000;
      24693: inst = 32'hc404dd8;
      24694: inst = 32'h8220000;
      24695: inst = 32'h10408000;
      24696: inst = 32'hc404ddb;
      24697: inst = 32'h8220000;
      24698: inst = 32'h10408000;
      24699: inst = 32'hc404ddd;
      24700: inst = 32'h8220000;
      24701: inst = 32'h10408000;
      24702: inst = 32'hc404ddf;
      24703: inst = 32'h8220000;
      24704: inst = 32'h10408000;
      24705: inst = 32'hc404de9;
      24706: inst = 32'h8220000;
      24707: inst = 32'h10408000;
      24708: inst = 32'hc404df1;
      24709: inst = 32'h8220000;
      24710: inst = 32'h10408000;
      24711: inst = 32'hc404df9;
      24712: inst = 32'h8220000;
      24713: inst = 32'h10408000;
      24714: inst = 32'hc404dfb;
      24715: inst = 32'h8220000;
      24716: inst = 32'h10408000;
      24717: inst = 32'hc404dfd;
      24718: inst = 32'h8220000;
      24719: inst = 32'h10408000;
      24720: inst = 32'hc404e02;
      24721: inst = 32'h8220000;
      24722: inst = 32'h10408000;
      24723: inst = 32'hc404e08;
      24724: inst = 32'h8220000;
      24725: inst = 32'h10408000;
      24726: inst = 32'hc404e0a;
      24727: inst = 32'h8220000;
      24728: inst = 32'h10408000;
      24729: inst = 32'hc404e0f;
      24730: inst = 32'h8220000;
      24731: inst = 32'h10408000;
      24732: inst = 32'hc404e2b;
      24733: inst = 32'h8220000;
      24734: inst = 32'h10408000;
      24735: inst = 32'hc404e35;
      24736: inst = 32'h8220000;
      24737: inst = 32'h10408000;
      24738: inst = 32'hc404e43;
      24739: inst = 32'h8220000;
      24740: inst = 32'h10408000;
      24741: inst = 32'hc404e4d;
      24742: inst = 32'h8220000;
      24743: inst = 32'h10408000;
      24744: inst = 32'hc404e4e;
      24745: inst = 32'h8220000;
      24746: inst = 32'h10408000;
      24747: inst = 32'hc404e61;
      24748: inst = 32'h8220000;
      24749: inst = 32'h10408000;
      24750: inst = 32'hc404e66;
      24751: inst = 32'h8220000;
      24752: inst = 32'h10408000;
      24753: inst = 32'hc404e6c;
      24754: inst = 32'h8220000;
      24755: inst = 32'h10408000;
      24756: inst = 32'hc404e73;
      24757: inst = 32'h8220000;
      24758: inst = 32'h10408000;
      24759: inst = 32'hc404eeb;
      24760: inst = 32'h8220000;
      24761: inst = 32'h10408000;
      24762: inst = 32'hc404f0d;
      24763: inst = 32'h8220000;
      24764: inst = 32'h10408000;
      24765: inst = 32'hc404f18;
      24766: inst = 32'h8220000;
      24767: inst = 32'h10408000;
      24768: inst = 32'hc404f27;
      24769: inst = 32'h8220000;
      24770: inst = 32'h10408000;
      24771: inst = 32'hc404f34;
      24772: inst = 32'h8220000;
      24773: inst = 32'h10408000;
      24774: inst = 32'hc404f6d;
      24775: inst = 32'h8220000;
      24776: inst = 32'h10408000;
      24777: inst = 32'hc405015;
      24778: inst = 32'h8220000;
      24779: inst = 32'h10408000;
      24780: inst = 32'hc40502e;
      24781: inst = 32'h8220000;
      24782: inst = 32'h10408000;
      24783: inst = 32'hc405056;
      24784: inst = 32'h8220000;
      24785: inst = 32'h10408000;
      24786: inst = 32'hc40506e;
      24787: inst = 32'h8220000;
      24788: inst = 32'h10408000;
      24789: inst = 32'hc405073;
      24790: inst = 32'h8220000;
      24791: inst = 32'h10408000;
      24792: inst = 32'hc40507b;
      24793: inst = 32'h8220000;
      24794: inst = 32'h10408000;
      24795: inst = 32'hc40509a;
      24796: inst = 32'h8220000;
      24797: inst = 32'h10408000;
      24798: inst = 32'hc4050a9;
      24799: inst = 32'h8220000;
      24800: inst = 32'h10408000;
      24801: inst = 32'hc4050af;
      24802: inst = 32'h8220000;
      24803: inst = 32'h10408000;
      24804: inst = 32'hc4050b4;
      24805: inst = 32'h8220000;
      24806: inst = 32'hc208c71;
      24807: inst = 32'h10408000;
      24808: inst = 32'hc4047a7;
      24809: inst = 32'h8220000;
      24810: inst = 32'h10408000;
      24811: inst = 32'hc404832;
      24812: inst = 32'h8220000;
      24813: inst = 32'h10408000;
      24814: inst = 32'hc404868;
      24815: inst = 32'h8220000;
      24816: inst = 32'h10408000;
      24817: inst = 32'hc4048a7;
      24818: inst = 32'h8220000;
      24819: inst = 32'h10408000;
      24820: inst = 32'hc4048b6;
      24821: inst = 32'h8220000;
      24822: inst = 32'h10408000;
      24823: inst = 32'hc4048ca;
      24824: inst = 32'h8220000;
      24825: inst = 32'h10408000;
      24826: inst = 32'hc404907;
      24827: inst = 32'h8220000;
      24828: inst = 32'h10408000;
      24829: inst = 32'hc404916;
      24830: inst = 32'h8220000;
      24831: inst = 32'h10408000;
      24832: inst = 32'hc40492a;
      24833: inst = 32'h8220000;
      24834: inst = 32'h10408000;
      24835: inst = 32'hc404952;
      24836: inst = 32'h8220000;
      24837: inst = 32'h10408000;
      24838: inst = 32'hc4049db;
      24839: inst = 32'h8220000;
      24840: inst = 32'h10408000;
      24841: inst = 32'hc404e3f;
      24842: inst = 32'h8220000;
      24843: inst = 32'h10408000;
      24844: inst = 32'hc404e49;
      24845: inst = 32'h8220000;
      24846: inst = 32'h10408000;
      24847: inst = 32'hc404e5d;
      24848: inst = 32'h8220000;
      24849: inst = 32'h10408000;
      24850: inst = 32'hc404e62;
      24851: inst = 32'h8220000;
      24852: inst = 32'h10408000;
      24853: inst = 32'hc404ecf;
      24854: inst = 32'h8220000;
      24855: inst = 32'h10408000;
      24856: inst = 32'hc404f79;
      24857: inst = 32'h8220000;
      24858: inst = 32'h10408000;
      24859: inst = 32'hc404f88;
      24860: inst = 32'h8220000;
      24861: inst = 32'h10408000;
      24862: inst = 32'hc404fed;
      24863: inst = 32'h8220000;
      24864: inst = 32'hc20d69a;
      24865: inst = 32'h10408000;
      24866: inst = 32'hc4047d0;
      24867: inst = 32'h8220000;
      24868: inst = 32'h10408000;
      24869: inst = 32'hc4047da;
      24870: inst = 32'h8220000;
      24871: inst = 32'h10408000;
      24872: inst = 32'hc4047f5;
      24873: inst = 32'h8220000;
      24874: inst = 32'h10408000;
      24875: inst = 32'hc4047fd;
      24876: inst = 32'h8220000;
      24877: inst = 32'h10408000;
      24878: inst = 32'hc4048a8;
      24879: inst = 32'h8220000;
      24880: inst = 32'h10408000;
      24881: inst = 32'hc4048b7;
      24882: inst = 32'h8220000;
      24883: inst = 32'h10408000;
      24884: inst = 32'hc4048cb;
      24885: inst = 32'h8220000;
      24886: inst = 32'h10408000;
      24887: inst = 32'hc404953;
      24888: inst = 32'h8220000;
      24889: inst = 32'h10408000;
      24890: inst = 32'hc4049b2;
      24891: inst = 32'h8220000;
      24892: inst = 32'h10408000;
      24893: inst = 32'hc4049cb;
      24894: inst = 32'h8220000;
      24895: inst = 32'h10408000;
      24896: inst = 32'hc4049da;
      24897: inst = 32'h8220000;
      24898: inst = 32'h10408000;
      24899: inst = 32'hc4049ee;
      24900: inst = 32'h8220000;
      24901: inst = 32'h10408000;
      24902: inst = 32'hc404e33;
      24903: inst = 32'h8220000;
      24904: inst = 32'h10408000;
      24905: inst = 32'hc404e36;
      24906: inst = 32'h8220000;
      24907: inst = 32'h10408000;
      24908: inst = 32'hc404e38;
      24909: inst = 32'h8220000;
      24910: inst = 32'h10408000;
      24911: inst = 32'hc404e4f;
      24912: inst = 32'h8220000;
      24913: inst = 32'h10408000;
      24914: inst = 32'hc404e51;
      24915: inst = 32'h8220000;
      24916: inst = 32'h10408000;
      24917: inst = 32'hc404e5b;
      24918: inst = 32'h8220000;
      24919: inst = 32'h10408000;
      24920: inst = 32'hc404e6a;
      24921: inst = 32'h8220000;
      24922: inst = 32'h10408000;
      24923: inst = 32'hc404e6d;
      24924: inst = 32'h8220000;
      24925: inst = 32'h10408000;
      24926: inst = 32'hc404eed;
      24927: inst = 32'h8220000;
      24928: inst = 32'h10408000;
      24929: inst = 32'hc404efa;
      24930: inst = 32'h8220000;
      24931: inst = 32'h10408000;
      24932: inst = 32'hc404f1a;
      24933: inst = 32'h8220000;
      24934: inst = 32'h10408000;
      24935: inst = 32'hc404f1b;
      24936: inst = 32'h8220000;
      24937: inst = 32'h10408000;
      24938: inst = 32'hc404f29;
      24939: inst = 32'h8220000;
      24940: inst = 32'h10408000;
      24941: inst = 32'hc404f2a;
      24942: inst = 32'h8220000;
      24943: inst = 32'h10408000;
      24944: inst = 32'hc404f5a;
      24945: inst = 32'h8220000;
      24946: inst = 32'h10408000;
      24947: inst = 32'hc404fba;
      24948: inst = 32'h8220000;
      24949: inst = 32'h10408000;
      24950: inst = 32'hc404fe6;
      24951: inst = 32'h8220000;
      24952: inst = 32'h10408000;
      24953: inst = 32'hc40500c;
      24954: inst = 32'h8220000;
      24955: inst = 32'h10408000;
      24956: inst = 32'hc405038;
      24957: inst = 32'h8220000;
      24958: inst = 32'h10408000;
      24959: inst = 32'hc40503b;
      24960: inst = 32'h8220000;
      24961: inst = 32'h10408000;
      24962: inst = 32'hc405047;
      24963: inst = 32'h8220000;
      24964: inst = 32'h10408000;
      24965: inst = 32'hc40504a;
      24966: inst = 32'h8220000;
      24967: inst = 32'hc20bdd7;
      24968: inst = 32'h10408000;
      24969: inst = 32'hc4047d1;
      24970: inst = 32'h8220000;
      24971: inst = 32'h10408000;
      24972: inst = 32'hc4047d6;
      24973: inst = 32'h8220000;
      24974: inst = 32'h10408000;
      24975: inst = 32'hc4047e5;
      24976: inst = 32'h8220000;
      24977: inst = 32'h10408000;
      24978: inst = 32'hc404803;
      24979: inst = 32'h8220000;
      24980: inst = 32'h10408000;
      24981: inst = 32'hc404855;
      24982: inst = 32'h8220000;
      24983: inst = 32'h10408000;
      24984: inst = 32'hc4049c9;
      24985: inst = 32'h8220000;
      24986: inst = 32'h10408000;
      24987: inst = 32'hc4049d8;
      24988: inst = 32'h8220000;
      24989: inst = 32'h10408000;
      24990: inst = 32'hc4049ec;
      24991: inst = 32'h8220000;
      24992: inst = 32'h10408000;
      24993: inst = 32'hc404de0;
      24994: inst = 32'h8220000;
      24995: inst = 32'h10408000;
      24996: inst = 32'hc404dea;
      24997: inst = 32'h8220000;
      24998: inst = 32'h10408000;
      24999: inst = 32'hc404dfe;
      25000: inst = 32'h8220000;
      25001: inst = 32'h10408000;
      25002: inst = 32'hc404e03;
      25003: inst = 32'h8220000;
      25004: inst = 32'h10408000;
      25005: inst = 32'hc404e2c;
      25006: inst = 32'h8220000;
      25007: inst = 32'h10408000;
      25008: inst = 32'hc404e2e;
      25009: inst = 32'h8220000;
      25010: inst = 32'h10408000;
      25011: inst = 32'hc404e32;
      25012: inst = 32'h8220000;
      25013: inst = 32'h10408000;
      25014: inst = 32'hc404e40;
      25015: inst = 32'h8220000;
      25016: inst = 32'h10408000;
      25017: inst = 32'hc404e4a;
      25018: inst = 32'h8220000;
      25019: inst = 32'h10408000;
      25020: inst = 32'hc404e5e;
      25021: inst = 32'h8220000;
      25022: inst = 32'h10408000;
      25023: inst = 32'hc404e63;
      25024: inst = 32'h8220000;
      25025: inst = 32'h10408000;
      25026: inst = 32'hc404e6f;
      25027: inst = 32'h8220000;
      25028: inst = 32'h10408000;
      25029: inst = 32'hc404e8f;
      25030: inst = 32'h8220000;
      25031: inst = 32'h10408000;
      25032: inst = 32'hc404ed0;
      25033: inst = 32'h8220000;
      25034: inst = 32'h10408000;
      25035: inst = 32'hc404fab;
      25036: inst = 32'h8220000;
      25037: inst = 32'h10408000;
      25038: inst = 32'hc405039;
      25039: inst = 32'h8220000;
      25040: inst = 32'h10408000;
      25041: inst = 32'hc405048;
      25042: inst = 32'h8220000;
      25043: inst = 32'h10408000;
      25044: inst = 32'hc40504f;
      25045: inst = 32'h8220000;
      25046: inst = 32'hc20ef5d;
      25047: inst = 32'h10408000;
      25048: inst = 32'hc4047dc;
      25049: inst = 32'h8220000;
      25050: inst = 32'h10408000;
      25051: inst = 32'hc4047ff;
      25052: inst = 32'h8220000;
      25053: inst = 32'h10408000;
      25054: inst = 32'hc404848;
      25055: inst = 32'h8220000;
      25056: inst = 32'h10408000;
      25057: inst = 32'hc404852;
      25058: inst = 32'h8220000;
      25059: inst = 32'h10408000;
      25060: inst = 32'hc404857;
      25061: inst = 32'h8220000;
      25062: inst = 32'h10408000;
      25063: inst = 32'hc40486b;
      25064: inst = 32'h8220000;
      25065: inst = 32'h10408000;
      25066: inst = 32'hc404968;
      25067: inst = 32'h8220000;
      25068: inst = 32'h10408000;
      25069: inst = 32'hc404977;
      25070: inst = 32'h8220000;
      25071: inst = 32'h10408000;
      25072: inst = 32'hc40498b;
      25073: inst = 32'h8220000;
      25074: inst = 32'h10408000;
      25075: inst = 32'hc404eec;
      25076: inst = 32'h8220000;
      25077: inst = 32'h10408000;
      25078: inst = 32'hc404f55;
      25079: inst = 32'h8220000;
      25080: inst = 32'h10408000;
      25081: inst = 32'hc404f6e;
      25082: inst = 32'h8220000;
      25083: inst = 32'h10408000;
      25084: inst = 32'hc404f78;
      25085: inst = 32'h8220000;
      25086: inst = 32'h10408000;
      25087: inst = 32'hc404f87;
      25088: inst = 32'h8220000;
      25089: inst = 32'h10408000;
      25090: inst = 32'hc404faf;
      25091: inst = 32'h8220000;
      25092: inst = 32'h10408000;
      25093: inst = 32'hc404ff4;
      25094: inst = 32'h8220000;
      25095: inst = 32'h10408000;
      25096: inst = 32'hc40501b;
      25097: inst = 32'h8220000;
      25098: inst = 32'h10408000;
      25099: inst = 32'hc40501e;
      25100: inst = 32'h8220000;
      25101: inst = 32'h10408000;
      25102: inst = 32'hc405021;
      25103: inst = 32'h8220000;
      25104: inst = 32'h10408000;
      25105: inst = 32'hc40502b;
      25106: inst = 32'h8220000;
      25107: inst = 32'h10408000;
      25108: inst = 32'hc40503c;
      25109: inst = 32'h8220000;
      25110: inst = 32'h10408000;
      25111: inst = 32'hc40503f;
      25112: inst = 32'h8220000;
      25113: inst = 32'h10408000;
      25114: inst = 32'hc405044;
      25115: inst = 32'h8220000;
      25116: inst = 32'h10408000;
      25117: inst = 32'hc40504b;
      25118: inst = 32'h8220000;
      25119: inst = 32'h10408000;
      25120: inst = 32'hc405055;
      25121: inst = 32'h8220000;
      25122: inst = 32'hc20c638;
      25123: inst = 32'h10408000;
      25124: inst = 32'hc4047e9;
      25125: inst = 32'h8220000;
      25126: inst = 32'h10408000;
      25127: inst = 32'hc4047f3;
      25128: inst = 32'h8220000;
      25129: inst = 32'h10408000;
      25130: inst = 32'hc4047f8;
      25131: inst = 32'h8220000;
      25132: inst = 32'h10408000;
      25133: inst = 32'hc40480c;
      25134: inst = 32'h8220000;
      25135: inst = 32'h10408000;
      25136: inst = 32'hc404835;
      25137: inst = 32'h8220000;
      25138: inst = 32'h10408000;
      25139: inst = 32'hc404844;
      25140: inst = 32'h8220000;
      25141: inst = 32'h10408000;
      25142: inst = 32'hc40484c;
      25143: inst = 32'h8220000;
      25144: inst = 32'h10408000;
      25145: inst = 32'hc40485b;
      25146: inst = 32'h8220000;
      25147: inst = 32'h10408000;
      25148: inst = 32'hc404862;
      25149: inst = 32'h8220000;
      25150: inst = 32'h10408000;
      25151: inst = 32'hc40486f;
      25152: inst = 32'h8220000;
      25153: inst = 32'h10408000;
      25154: inst = 32'hc404895;
      25155: inst = 32'h8220000;
      25156: inst = 32'h10408000;
      25157: inst = 32'hc40489d;
      25158: inst = 32'h8220000;
      25159: inst = 32'h10408000;
      25160: inst = 32'hc4048a4;
      25161: inst = 32'h8220000;
      25162: inst = 32'h10408000;
      25163: inst = 32'hc4048c0;
      25164: inst = 32'h8220000;
      25165: inst = 32'h10408000;
      25166: inst = 32'hc4048c2;
      25167: inst = 32'h8220000;
      25168: inst = 32'h10408000;
      25169: inst = 32'hc4048f5;
      25170: inst = 32'h8220000;
      25171: inst = 32'h10408000;
      25172: inst = 32'hc4048fd;
      25173: inst = 32'h8220000;
      25174: inst = 32'h10408000;
      25175: inst = 32'hc404904;
      25176: inst = 32'h8220000;
      25177: inst = 32'h10408000;
      25178: inst = 32'hc404908;
      25179: inst = 32'h8220000;
      25180: inst = 32'h10408000;
      25181: inst = 32'hc404917;
      25182: inst = 32'h8220000;
      25183: inst = 32'h10408000;
      25184: inst = 32'hc404920;
      25185: inst = 32'h8220000;
      25186: inst = 32'h10408000;
      25187: inst = 32'hc404922;
      25188: inst = 32'h8220000;
      25189: inst = 32'h10408000;
      25190: inst = 32'hc40492b;
      25191: inst = 32'h8220000;
      25192: inst = 32'h10408000;
      25193: inst = 32'hc404955;
      25194: inst = 32'h8220000;
      25195: inst = 32'h10408000;
      25196: inst = 32'hc40495d;
      25197: inst = 32'h8220000;
      25198: inst = 32'h10408000;
      25199: inst = 32'hc404964;
      25200: inst = 32'h8220000;
      25201: inst = 32'h10408000;
      25202: inst = 32'hc404980;
      25203: inst = 32'h8220000;
      25204: inst = 32'h10408000;
      25205: inst = 32'hc404982;
      25206: inst = 32'h8220000;
      25207: inst = 32'h10408000;
      25208: inst = 32'hc4049b0;
      25209: inst = 32'h8220000;
      25210: inst = 32'h10408000;
      25211: inst = 32'hc4049b7;
      25212: inst = 32'h8220000;
      25213: inst = 32'h10408000;
      25214: inst = 32'hc4049bc;
      25215: inst = 32'h8220000;
      25216: inst = 32'h10408000;
      25217: inst = 32'hc4049c6;
      25218: inst = 32'h8220000;
      25219: inst = 32'h10408000;
      25220: inst = 32'hc4049d5;
      25221: inst = 32'h8220000;
      25222: inst = 32'h10408000;
      25223: inst = 32'hc4049df;
      25224: inst = 32'h8220000;
      25225: inst = 32'h10408000;
      25226: inst = 32'hc4049e4;
      25227: inst = 32'h8220000;
      25228: inst = 32'h10408000;
      25229: inst = 32'hc404d70;
      25230: inst = 32'h8220000;
      25231: inst = 32'h10408000;
      25232: inst = 32'hc404d81;
      25233: inst = 32'h8220000;
      25234: inst = 32'h10408000;
      25235: inst = 32'hc404d8b;
      25236: inst = 32'h8220000;
      25237: inst = 32'h10408000;
      25238: inst = 32'hc404d9f;
      25239: inst = 32'h8220000;
      25240: inst = 32'h10408000;
      25241: inst = 32'hc404da4;
      25242: inst = 32'h8220000;
      25243: inst = 32'h10408000;
      25244: inst = 32'hc404db1;
      25245: inst = 32'h8220000;
      25246: inst = 32'h10408000;
      25247: inst = 32'hc404dd0;
      25248: inst = 32'h8220000;
      25249: inst = 32'h10408000;
      25250: inst = 32'hc404de1;
      25251: inst = 32'h8220000;
      25252: inst = 32'h10408000;
      25253: inst = 32'hc404deb;
      25254: inst = 32'h8220000;
      25255: inst = 32'h10408000;
      25256: inst = 32'hc404dff;
      25257: inst = 32'h8220000;
      25258: inst = 32'h10408000;
      25259: inst = 32'hc404e04;
      25260: inst = 32'h8220000;
      25261: inst = 32'h10408000;
      25262: inst = 32'hc404e11;
      25263: inst = 32'h8220000;
      25264: inst = 32'h10408000;
      25265: inst = 32'hc404e2f;
      25266: inst = 32'h8220000;
      25267: inst = 32'h10408000;
      25268: inst = 32'hc404e30;
      25269: inst = 32'h8220000;
      25270: inst = 32'h10408000;
      25271: inst = 32'hc404e3e;
      25272: inst = 32'h8220000;
      25273: inst = 32'h10408000;
      25274: inst = 32'hc404e71;
      25275: inst = 32'h8220000;
      25276: inst = 32'h10408000;
      25277: inst = 32'hc404e90;
      25278: inst = 32'h8220000;
      25279: inst = 32'h10408000;
      25280: inst = 32'hc404e9a;
      25281: inst = 32'h8220000;
      25282: inst = 32'h10408000;
      25283: inst = 32'hc404e9e;
      25284: inst = 32'h8220000;
      25285: inst = 32'h10408000;
      25286: inst = 32'hc404ea1;
      25287: inst = 32'h8220000;
      25288: inst = 32'h10408000;
      25289: inst = 32'hc404eab;
      25290: inst = 32'h8220000;
      25291: inst = 32'h10408000;
      25292: inst = 32'hc404eb8;
      25293: inst = 32'h8220000;
      25294: inst = 32'h10408000;
      25295: inst = 32'hc404ebc;
      25296: inst = 32'h8220000;
      25297: inst = 32'h10408000;
      25298: inst = 32'hc404ebf;
      25299: inst = 32'h8220000;
      25300: inst = 32'h10408000;
      25301: inst = 32'hc404ec4;
      25302: inst = 32'h8220000;
      25303: inst = 32'h10408000;
      25304: inst = 32'hc404ec7;
      25305: inst = 32'h8220000;
      25306: inst = 32'h10408000;
      25307: inst = 32'hc404ecb;
      25308: inst = 32'h8220000;
      25309: inst = 32'h10408000;
      25310: inst = 32'hc404ecc;
      25311: inst = 32'h8220000;
      25312: inst = 32'h10408000;
      25313: inst = 32'hc404ed1;
      25314: inst = 32'h8220000;
      25315: inst = 32'h10408000;
      25316: inst = 32'hc404ef0;
      25317: inst = 32'h8220000;
      25318: inst = 32'h10408000;
      25319: inst = 32'hc404efe;
      25320: inst = 32'h8220000;
      25321: inst = 32'h10408000;
      25322: inst = 32'hc404f01;
      25323: inst = 32'h8220000;
      25324: inst = 32'h10408000;
      25325: inst = 32'hc404f0b;
      25326: inst = 32'h8220000;
      25327: inst = 32'h10408000;
      25328: inst = 32'hc404f1c;
      25329: inst = 32'h8220000;
      25330: inst = 32'h10408000;
      25331: inst = 32'hc404f1f;
      25332: inst = 32'h8220000;
      25333: inst = 32'h10408000;
      25334: inst = 32'hc404f24;
      25335: inst = 32'h8220000;
      25336: inst = 32'h10408000;
      25337: inst = 32'hc404f2b;
      25338: inst = 32'h8220000;
      25339: inst = 32'h10408000;
      25340: inst = 32'hc404f31;
      25341: inst = 32'h8220000;
      25342: inst = 32'h10408000;
      25343: inst = 32'hc404f32;
      25344: inst = 32'h8220000;
      25345: inst = 32'h10408000;
      25346: inst = 32'hc404f50;
      25347: inst = 32'h8220000;
      25348: inst = 32'h10408000;
      25349: inst = 32'hc404f5e;
      25350: inst = 32'h8220000;
      25351: inst = 32'h10408000;
      25352: inst = 32'hc404f61;
      25353: inst = 32'h8220000;
      25354: inst = 32'h10408000;
      25355: inst = 32'hc404f6b;
      25356: inst = 32'h8220000;
      25357: inst = 32'h10408000;
      25358: inst = 32'hc404f7c;
      25359: inst = 32'h8220000;
      25360: inst = 32'h10408000;
      25361: inst = 32'hc404f7f;
      25362: inst = 32'h8220000;
      25363: inst = 32'h10408000;
      25364: inst = 32'hc404f84;
      25365: inst = 32'h8220000;
      25366: inst = 32'h10408000;
      25367: inst = 32'hc404f8b;
      25368: inst = 32'h8220000;
      25369: inst = 32'h10408000;
      25370: inst = 32'hc404f91;
      25371: inst = 32'h8220000;
      25372: inst = 32'h10408000;
      25373: inst = 32'hc404f92;
      25374: inst = 32'h8220000;
      25375: inst = 32'h10408000;
      25376: inst = 32'hc404f94;
      25377: inst = 32'h8220000;
      25378: inst = 32'h10408000;
      25379: inst = 32'hc404fb0;
      25380: inst = 32'h8220000;
      25381: inst = 32'h10408000;
      25382: inst = 32'hc404fbe;
      25383: inst = 32'h8220000;
      25384: inst = 32'h10408000;
      25385: inst = 32'hc404fc1;
      25386: inst = 32'h8220000;
      25387: inst = 32'h10408000;
      25388: inst = 32'hc404fcb;
      25389: inst = 32'h8220000;
      25390: inst = 32'h10408000;
      25391: inst = 32'hc404fdc;
      25392: inst = 32'h8220000;
      25393: inst = 32'h10408000;
      25394: inst = 32'hc404fdf;
      25395: inst = 32'h8220000;
      25396: inst = 32'h10408000;
      25397: inst = 32'hc404fe4;
      25398: inst = 32'h8220000;
      25399: inst = 32'h10408000;
      25400: inst = 32'hc404feb;
      25401: inst = 32'h8220000;
      25402: inst = 32'h10408000;
      25403: inst = 32'hc404ff1;
      25404: inst = 32'h8220000;
      25405: inst = 32'h10408000;
      25406: inst = 32'hc40500b;
      25407: inst = 32'h8220000;
      25408: inst = 32'h10408000;
      25409: inst = 32'hc405011;
      25410: inst = 32'h8220000;
      25411: inst = 32'h10408000;
      25412: inst = 32'hc405016;
      25413: inst = 32'h8220000;
      25414: inst = 32'h10408000;
      25415: inst = 32'hc405018;
      25416: inst = 32'h8220000;
      25417: inst = 32'h10408000;
      25418: inst = 32'hc40501c;
      25419: inst = 32'h8220000;
      25420: inst = 32'h10408000;
      25421: inst = 32'hc40501d;
      25422: inst = 32'h8220000;
      25423: inst = 32'h10408000;
      25424: inst = 32'hc405022;
      25425: inst = 32'h8220000;
      25426: inst = 32'h10408000;
      25427: inst = 32'hc40502c;
      25428: inst = 32'h8220000;
      25429: inst = 32'h10408000;
      25430: inst = 32'hc40502f;
      25431: inst = 32'h8220000;
      25432: inst = 32'h10408000;
      25433: inst = 32'hc405031;
      25434: inst = 32'h8220000;
      25435: inst = 32'h10408000;
      25436: inst = 32'hc405040;
      25437: inst = 32'h8220000;
      25438: inst = 32'h10408000;
      25439: inst = 32'hc405045;
      25440: inst = 32'h8220000;
      25441: inst = 32'h10408000;
      25442: inst = 32'hc405052;
      25443: inst = 32'h8220000;
      25444: inst = 32'hc20ffff;
      25445: inst = 32'h10408000;
      25446: inst = 32'hc404fec;
      25447: inst = 32'h8220000;
      25448: inst = 32'h58000000;
      25449: inst = 32'h13e0ffff;
      25450: inst = 32'h13e00000;
      25451: inst = 32'hfe06380;
      25452: inst = 32'h5be00000;
      25453: inst = 32'h13e0ffff;
      25454: inst = 32'h13e00000;
      25455: inst = 32'hfe06529;
      25456: inst = 32'h5be00000;
      25457: inst = 32'h13e0ffff;
      25458: inst = 32'h13e00000;
      25459: inst = 32'hfe06529;
      25460: inst = 32'h5be00000;
      25461: inst = 32'h13e0ffff;
      25462: inst = 32'h13e00000;
      25463: inst = 32'hfe06454;
      25464: inst = 32'h5be00000;
      25465: inst = 32'h13e0ffff;
      25466: inst = 32'h13e00000;
      25467: inst = 32'hfe06454;
      25468: inst = 32'h5be00000;
      25469: inst = 32'h13e00000;
      25470: inst = 32'hfe06380;
      25471: inst = 32'h5be00000;
      25472: inst = 32'hc60f4ce;
      25473: inst = 32'h10408000;
      25474: inst = 32'hc404a8c;
      25475: inst = 32'h8620000;
      25476: inst = 32'h10408000;
      25477: inst = 32'hc404a8d;
      25478: inst = 32'h8620000;
      25479: inst = 32'h10408000;
      25480: inst = 32'hc404a8e;
      25481: inst = 32'h8620000;
      25482: inst = 32'h10408000;
      25483: inst = 32'hc404a8f;
      25484: inst = 32'h8620000;
      25485: inst = 32'h10408000;
      25486: inst = 32'hc404a90;
      25487: inst = 32'h8620000;
      25488: inst = 32'h10408000;
      25489: inst = 32'hc404a91;
      25490: inst = 32'h8620000;
      25491: inst = 32'h10408000;
      25492: inst = 32'hc404a92;
      25493: inst = 32'h8620000;
      25494: inst = 32'h10408000;
      25495: inst = 32'hc404a93;
      25496: inst = 32'h8620000;
      25497: inst = 32'h10408000;
      25498: inst = 32'hc404aec;
      25499: inst = 32'h8620000;
      25500: inst = 32'h10408000;
      25501: inst = 32'hc404aee;
      25502: inst = 32'h8620000;
      25503: inst = 32'h10408000;
      25504: inst = 32'hc404aef;
      25505: inst = 32'h8620000;
      25506: inst = 32'h10408000;
      25507: inst = 32'hc404af0;
      25508: inst = 32'h8620000;
      25509: inst = 32'h10408000;
      25510: inst = 32'hc404af1;
      25511: inst = 32'h8620000;
      25512: inst = 32'h10408000;
      25513: inst = 32'hc404af3;
      25514: inst = 32'h8620000;
      25515: inst = 32'h10408000;
      25516: inst = 32'hc404b4c;
      25517: inst = 32'h8620000;
      25518: inst = 32'h10408000;
      25519: inst = 32'hc404b4e;
      25520: inst = 32'h8620000;
      25521: inst = 32'h10408000;
      25522: inst = 32'hc404b4f;
      25523: inst = 32'h8620000;
      25524: inst = 32'h10408000;
      25525: inst = 32'hc404b50;
      25526: inst = 32'h8620000;
      25527: inst = 32'h10408000;
      25528: inst = 32'hc404b51;
      25529: inst = 32'h8620000;
      25530: inst = 32'h10408000;
      25531: inst = 32'hc404b53;
      25532: inst = 32'h8620000;
      25533: inst = 32'h10408000;
      25534: inst = 32'hc404bac;
      25535: inst = 32'h8620000;
      25536: inst = 32'h10408000;
      25537: inst = 32'hc404bad;
      25538: inst = 32'h8620000;
      25539: inst = 32'h10408000;
      25540: inst = 32'hc404bae;
      25541: inst = 32'h8620000;
      25542: inst = 32'h10408000;
      25543: inst = 32'hc404baf;
      25544: inst = 32'h8620000;
      25545: inst = 32'h10408000;
      25546: inst = 32'hc404bb0;
      25547: inst = 32'h8620000;
      25548: inst = 32'h10408000;
      25549: inst = 32'hc404bb1;
      25550: inst = 32'h8620000;
      25551: inst = 32'h10408000;
      25552: inst = 32'hc404bb2;
      25553: inst = 32'h8620000;
      25554: inst = 32'h10408000;
      25555: inst = 32'hc404bb3;
      25556: inst = 32'h8620000;
      25557: inst = 32'h10408000;
      25558: inst = 32'hc404c0c;
      25559: inst = 32'h8620000;
      25560: inst = 32'h10408000;
      25561: inst = 32'hc404c0d;
      25562: inst = 32'h8620000;
      25563: inst = 32'h10408000;
      25564: inst = 32'hc404c0e;
      25565: inst = 32'h8620000;
      25566: inst = 32'h10408000;
      25567: inst = 32'hc404c0f;
      25568: inst = 32'h8620000;
      25569: inst = 32'h10408000;
      25570: inst = 32'hc404c10;
      25571: inst = 32'h8620000;
      25572: inst = 32'h10408000;
      25573: inst = 32'hc404c11;
      25574: inst = 32'h8620000;
      25575: inst = 32'h10408000;
      25576: inst = 32'hc404c12;
      25577: inst = 32'h8620000;
      25578: inst = 32'h10408000;
      25579: inst = 32'hc404c13;
      25580: inst = 32'h8620000;
      25581: inst = 32'h10408000;
      25582: inst = 32'hc404ccb;
      25583: inst = 32'h8620000;
      25584: inst = 32'h10408000;
      25585: inst = 32'hc404ccc;
      25586: inst = 32'h8620000;
      25587: inst = 32'h10408000;
      25588: inst = 32'hc404cd3;
      25589: inst = 32'h8620000;
      25590: inst = 32'h10408000;
      25591: inst = 32'hc404cd4;
      25592: inst = 32'h8620000;
      25593: inst = 32'h10408000;
      25594: inst = 32'hc404e4e;
      25595: inst = 32'h8620000;
      25596: inst = 32'h10408000;
      25597: inst = 32'hc404e51;
      25598: inst = 32'h8620000;
      25599: inst = 32'hc607800;
      25600: inst = 32'h10408000;
      25601: inst = 32'hc404c6d;
      25602: inst = 32'h8620000;
      25603: inst = 32'h10408000;
      25604: inst = 32'hc404c6e;
      25605: inst = 32'h8620000;
      25606: inst = 32'h10408000;
      25607: inst = 32'hc404c71;
      25608: inst = 32'h8620000;
      25609: inst = 32'h10408000;
      25610: inst = 32'hc404c72;
      25611: inst = 32'h8620000;
      25612: inst = 32'hc60a000;
      25613: inst = 32'h10408000;
      25614: inst = 32'hc404c6f;
      25615: inst = 32'h8620000;
      25616: inst = 32'h10408000;
      25617: inst = 32'hc404c70;
      25618: inst = 32'h8620000;
      25619: inst = 32'h10408000;
      25620: inst = 32'hc404ccd;
      25621: inst = 32'h8620000;
      25622: inst = 32'h10408000;
      25623: inst = 32'hc404cce;
      25624: inst = 32'h8620000;
      25625: inst = 32'h10408000;
      25626: inst = 32'hc404ccf;
      25627: inst = 32'h8620000;
      25628: inst = 32'h10408000;
      25629: inst = 32'hc404cd0;
      25630: inst = 32'h8620000;
      25631: inst = 32'h10408000;
      25632: inst = 32'hc404cd1;
      25633: inst = 32'h8620000;
      25634: inst = 32'h10408000;
      25635: inst = 32'hc404cd2;
      25636: inst = 32'h8620000;
      25637: inst = 32'h10408000;
      25638: inst = 32'hc404d2d;
      25639: inst = 32'h8620000;
      25640: inst = 32'h10408000;
      25641: inst = 32'hc404d2e;
      25642: inst = 32'h8620000;
      25643: inst = 32'h10408000;
      25644: inst = 32'hc404d2f;
      25645: inst = 32'h8620000;
      25646: inst = 32'h10408000;
      25647: inst = 32'hc404d30;
      25648: inst = 32'h8620000;
      25649: inst = 32'h10408000;
      25650: inst = 32'hc404d31;
      25651: inst = 32'h8620000;
      25652: inst = 32'h10408000;
      25653: inst = 32'hc404d32;
      25654: inst = 32'h8620000;
      25655: inst = 32'hc6010ac;
      25656: inst = 32'h10408000;
      25657: inst = 32'hc404d8d;
      25658: inst = 32'h8620000;
      25659: inst = 32'h10408000;
      25660: inst = 32'hc404d8e;
      25661: inst = 32'h8620000;
      25662: inst = 32'h10408000;
      25663: inst = 32'hc404d8f;
      25664: inst = 32'h8620000;
      25665: inst = 32'h10408000;
      25666: inst = 32'hc404d90;
      25667: inst = 32'h8620000;
      25668: inst = 32'h10408000;
      25669: inst = 32'hc404d91;
      25670: inst = 32'h8620000;
      25671: inst = 32'h10408000;
      25672: inst = 32'hc404d92;
      25673: inst = 32'h8620000;
      25674: inst = 32'hc60d42c;
      25675: inst = 32'h10408000;
      25676: inst = 32'hc404dee;
      25677: inst = 32'h8620000;
      25678: inst = 32'h10408000;
      25679: inst = 32'hc404df1;
      25680: inst = 32'h8620000;
      25681: inst = 32'h13e00000;
      25682: inst = 32'hfe065fe;
      25683: inst = 32'h5be00000;
      25684: inst = 32'hc60d42c;
      25685: inst = 32'h10408000;
      25686: inst = 32'hc404a8d;
      25687: inst = 32'h8620000;
      25688: inst = 32'h10408000;
      25689: inst = 32'hc404a8e;
      25690: inst = 32'h8620000;
      25691: inst = 32'h10408000;
      25692: inst = 32'hc404a8f;
      25693: inst = 32'h8620000;
      25694: inst = 32'h10408000;
      25695: inst = 32'hc404a90;
      25696: inst = 32'h8620000;
      25697: inst = 32'h10408000;
      25698: inst = 32'hc404a91;
      25699: inst = 32'h8620000;
      25700: inst = 32'h10408000;
      25701: inst = 32'hc404a92;
      25702: inst = 32'h8620000;
      25703: inst = 32'h10408000;
      25704: inst = 32'hc404a93;
      25705: inst = 32'h8620000;
      25706: inst = 32'h10408000;
      25707: inst = 32'hc404a94;
      25708: inst = 32'h8620000;
      25709: inst = 32'h10408000;
      25710: inst = 32'hc404bad;
      25711: inst = 32'h8620000;
      25712: inst = 32'h10408000;
      25713: inst = 32'hc404c0d;
      25714: inst = 32'h8620000;
      25715: inst = 32'h10408000;
      25716: inst = 32'hc404dee;
      25717: inst = 32'h8620000;
      25718: inst = 32'h10408000;
      25719: inst = 32'hc404df1;
      25720: inst = 32'h8620000;
      25721: inst = 32'hc60f4ce;
      25722: inst = 32'h10408000;
      25723: inst = 32'hc404aec;
      25724: inst = 32'h8620000;
      25725: inst = 32'h10408000;
      25726: inst = 32'hc404aed;
      25727: inst = 32'h8620000;
      25728: inst = 32'h10408000;
      25729: inst = 32'hc404aee;
      25730: inst = 32'h8620000;
      25731: inst = 32'h10408000;
      25732: inst = 32'hc404aef;
      25733: inst = 32'h8620000;
      25734: inst = 32'h10408000;
      25735: inst = 32'hc404af0;
      25736: inst = 32'h8620000;
      25737: inst = 32'h10408000;
      25738: inst = 32'hc404af1;
      25739: inst = 32'h8620000;
      25740: inst = 32'h10408000;
      25741: inst = 32'hc404af2;
      25742: inst = 32'h8620000;
      25743: inst = 32'h10408000;
      25744: inst = 32'hc404af4;
      25745: inst = 32'h8620000;
      25746: inst = 32'h10408000;
      25747: inst = 32'hc404b4c;
      25748: inst = 32'h8620000;
      25749: inst = 32'h10408000;
      25750: inst = 32'hc404b4d;
      25751: inst = 32'h8620000;
      25752: inst = 32'h10408000;
      25753: inst = 32'hc404b4e;
      25754: inst = 32'h8620000;
      25755: inst = 32'h10408000;
      25756: inst = 32'hc404b4f;
      25757: inst = 32'h8620000;
      25758: inst = 32'h10408000;
      25759: inst = 32'hc404b50;
      25760: inst = 32'h8620000;
      25761: inst = 32'h10408000;
      25762: inst = 32'hc404b51;
      25763: inst = 32'h8620000;
      25764: inst = 32'h10408000;
      25765: inst = 32'hc404b52;
      25766: inst = 32'h8620000;
      25767: inst = 32'h10408000;
      25768: inst = 32'hc404b54;
      25769: inst = 32'h8620000;
      25770: inst = 32'h10408000;
      25771: inst = 32'hc404bae;
      25772: inst = 32'h8620000;
      25773: inst = 32'h10408000;
      25774: inst = 32'hc404baf;
      25775: inst = 32'h8620000;
      25776: inst = 32'h10408000;
      25777: inst = 32'hc404bb0;
      25778: inst = 32'h8620000;
      25779: inst = 32'h10408000;
      25780: inst = 32'hc404bb1;
      25781: inst = 32'h8620000;
      25782: inst = 32'h10408000;
      25783: inst = 32'hc404bb2;
      25784: inst = 32'h8620000;
      25785: inst = 32'h10408000;
      25786: inst = 32'hc404bb3;
      25787: inst = 32'h8620000;
      25788: inst = 32'h10408000;
      25789: inst = 32'hc404bb4;
      25790: inst = 32'h8620000;
      25791: inst = 32'h10408000;
      25792: inst = 32'hc404c0e;
      25793: inst = 32'h8620000;
      25794: inst = 32'h10408000;
      25795: inst = 32'hc404c0f;
      25796: inst = 32'h8620000;
      25797: inst = 32'h10408000;
      25798: inst = 32'hc404c10;
      25799: inst = 32'h8620000;
      25800: inst = 32'h10408000;
      25801: inst = 32'hc404c11;
      25802: inst = 32'h8620000;
      25803: inst = 32'h10408000;
      25804: inst = 32'hc404c12;
      25805: inst = 32'h8620000;
      25806: inst = 32'h10408000;
      25807: inst = 32'hc404c13;
      25808: inst = 32'h8620000;
      25809: inst = 32'h10408000;
      25810: inst = 32'hc404c14;
      25811: inst = 32'h8620000;
      25812: inst = 32'h10408000;
      25813: inst = 32'hc404ccf;
      25814: inst = 32'h8620000;
      25815: inst = 32'hc607841;
      25816: inst = 32'h10408000;
      25817: inst = 32'hc404c6d;
      25818: inst = 32'h8620000;
      25819: inst = 32'h10408000;
      25820: inst = 32'hc404ccd;
      25821: inst = 32'h8620000;
      25822: inst = 32'hc60a000;
      25823: inst = 32'h10408000;
      25824: inst = 32'hc404c6e;
      25825: inst = 32'h8620000;
      25826: inst = 32'h10408000;
      25827: inst = 32'hc404c6f;
      25828: inst = 32'h8620000;
      25829: inst = 32'h10408000;
      25830: inst = 32'hc404c70;
      25831: inst = 32'h8620000;
      25832: inst = 32'h10408000;
      25833: inst = 32'hc404c71;
      25834: inst = 32'h8620000;
      25835: inst = 32'h10408000;
      25836: inst = 32'hc404c72;
      25837: inst = 32'h8620000;
      25838: inst = 32'h10408000;
      25839: inst = 32'hc404cce;
      25840: inst = 32'h8620000;
      25841: inst = 32'h10408000;
      25842: inst = 32'hc404cd0;
      25843: inst = 32'h8620000;
      25844: inst = 32'h10408000;
      25845: inst = 32'hc404cd1;
      25846: inst = 32'h8620000;
      25847: inst = 32'h10408000;
      25848: inst = 32'hc404cd2;
      25849: inst = 32'h8620000;
      25850: inst = 32'h10408000;
      25851: inst = 32'hc404d2d;
      25852: inst = 32'h8620000;
      25853: inst = 32'h10408000;
      25854: inst = 32'hc404d2e;
      25855: inst = 32'h8620000;
      25856: inst = 32'h10408000;
      25857: inst = 32'hc404d2f;
      25858: inst = 32'h8620000;
      25859: inst = 32'h10408000;
      25860: inst = 32'hc404d30;
      25861: inst = 32'h8620000;
      25862: inst = 32'h10408000;
      25863: inst = 32'hc404d31;
      25864: inst = 32'h8620000;
      25865: inst = 32'h10408000;
      25866: inst = 32'hc404d32;
      25867: inst = 32'h8620000;
      25868: inst = 32'hc6010ac;
      25869: inst = 32'h10408000;
      25870: inst = 32'hc404d8d;
      25871: inst = 32'h8620000;
      25872: inst = 32'h10408000;
      25873: inst = 32'hc404d8e;
      25874: inst = 32'h8620000;
      25875: inst = 32'h10408000;
      25876: inst = 32'hc404d8f;
      25877: inst = 32'h8620000;
      25878: inst = 32'h10408000;
      25879: inst = 32'hc404d90;
      25880: inst = 32'h8620000;
      25881: inst = 32'h10408000;
      25882: inst = 32'hc404d91;
      25883: inst = 32'h8620000;
      25884: inst = 32'h10408000;
      25885: inst = 32'hc404d92;
      25886: inst = 32'h8620000;
      25887: inst = 32'h13e0ffff;
      25888: inst = 32'h13e00000;
      25889: inst = 32'hfe06526;
      25890: inst = 32'h5be00000;
      25891: inst = 32'h13e00000;
      25892: inst = 32'hfe065fe;
      25893: inst = 32'h5be00000;
      25894: inst = 32'h13e00000;
      25895: inst = 32'hfe065fe;
      25896: inst = 32'h5be00000;
      25897: inst = 32'hc60d42c;
      25898: inst = 32'h10408000;
      25899: inst = 32'hc404ae9;
      25900: inst = 32'h8620000;
      25901: inst = 32'h10408000;
      25902: inst = 32'hc404ae8;
      25903: inst = 32'h8620000;
      25904: inst = 32'h10408000;
      25905: inst = 32'hc404ae7;
      25906: inst = 32'h8620000;
      25907: inst = 32'h10408000;
      25908: inst = 32'hc404ae6;
      25909: inst = 32'h8620000;
      25910: inst = 32'h10408000;
      25911: inst = 32'hc404ae5;
      25912: inst = 32'h8620000;
      25913: inst = 32'h10408000;
      25914: inst = 32'hc404ae4;
      25915: inst = 32'h8620000;
      25916: inst = 32'h10408000;
      25917: inst = 32'hc404ae3;
      25918: inst = 32'h8620000;
      25919: inst = 32'h10408000;
      25920: inst = 32'hc404ae2;
      25921: inst = 32'h8620000;
      25922: inst = 32'h10408000;
      25923: inst = 32'hc404c09;
      25924: inst = 32'h8620000;
      25925: inst = 32'h10408000;
      25926: inst = 32'hc404c69;
      25927: inst = 32'h8620000;
      25928: inst = 32'h10408000;
      25929: inst = 32'hc404e48;
      25930: inst = 32'h8620000;
      25931: inst = 32'h10408000;
      25932: inst = 32'hc404e45;
      25933: inst = 32'h8620000;
      25934: inst = 32'hc60f4ce;
      25935: inst = 32'h10408000;
      25936: inst = 32'hc404b4a;
      25937: inst = 32'h8620000;
      25938: inst = 32'h10408000;
      25939: inst = 32'hc404b49;
      25940: inst = 32'h8620000;
      25941: inst = 32'h10408000;
      25942: inst = 32'hc404b48;
      25943: inst = 32'h8620000;
      25944: inst = 32'h10408000;
      25945: inst = 32'hc404b47;
      25946: inst = 32'h8620000;
      25947: inst = 32'h10408000;
      25948: inst = 32'hc404b46;
      25949: inst = 32'h8620000;
      25950: inst = 32'h10408000;
      25951: inst = 32'hc404b45;
      25952: inst = 32'h8620000;
      25953: inst = 32'h10408000;
      25954: inst = 32'hc404b44;
      25955: inst = 32'h8620000;
      25956: inst = 32'h10408000;
      25957: inst = 32'hc404b42;
      25958: inst = 32'h8620000;
      25959: inst = 32'h10408000;
      25960: inst = 32'hc404baa;
      25961: inst = 32'h8620000;
      25962: inst = 32'h10408000;
      25963: inst = 32'hc404ba9;
      25964: inst = 32'h8620000;
      25965: inst = 32'h10408000;
      25966: inst = 32'hc404ba8;
      25967: inst = 32'h8620000;
      25968: inst = 32'h10408000;
      25969: inst = 32'hc404ba7;
      25970: inst = 32'h8620000;
      25971: inst = 32'h10408000;
      25972: inst = 32'hc404ba6;
      25973: inst = 32'h8620000;
      25974: inst = 32'h10408000;
      25975: inst = 32'hc404ba5;
      25976: inst = 32'h8620000;
      25977: inst = 32'h10408000;
      25978: inst = 32'hc404ba4;
      25979: inst = 32'h8620000;
      25980: inst = 32'h10408000;
      25981: inst = 32'hc404ba2;
      25982: inst = 32'h8620000;
      25983: inst = 32'h10408000;
      25984: inst = 32'hc404c08;
      25985: inst = 32'h8620000;
      25986: inst = 32'h10408000;
      25987: inst = 32'hc404c07;
      25988: inst = 32'h8620000;
      25989: inst = 32'h10408000;
      25990: inst = 32'hc404c06;
      25991: inst = 32'h8620000;
      25992: inst = 32'h10408000;
      25993: inst = 32'hc404c05;
      25994: inst = 32'h8620000;
      25995: inst = 32'h10408000;
      25996: inst = 32'hc404c04;
      25997: inst = 32'h8620000;
      25998: inst = 32'h10408000;
      25999: inst = 32'hc404c03;
      26000: inst = 32'h8620000;
      26001: inst = 32'h10408000;
      26002: inst = 32'hc404c02;
      26003: inst = 32'h8620000;
      26004: inst = 32'h10408000;
      26005: inst = 32'hc404c68;
      26006: inst = 32'h8620000;
      26007: inst = 32'h10408000;
      26008: inst = 32'hc404c67;
      26009: inst = 32'h8620000;
      26010: inst = 32'h10408000;
      26011: inst = 32'hc404c66;
      26012: inst = 32'h8620000;
      26013: inst = 32'h10408000;
      26014: inst = 32'hc404c65;
      26015: inst = 32'h8620000;
      26016: inst = 32'h10408000;
      26017: inst = 32'hc404c64;
      26018: inst = 32'h8620000;
      26019: inst = 32'h10408000;
      26020: inst = 32'hc404c63;
      26021: inst = 32'h8620000;
      26022: inst = 32'h10408000;
      26023: inst = 32'hc404c62;
      26024: inst = 32'h8620000;
      26025: inst = 32'h10408000;
      26026: inst = 32'hc404d27;
      26027: inst = 32'h8620000;
      26028: inst = 32'hc607841;
      26029: inst = 32'h10408000;
      26030: inst = 32'hc404cc9;
      26031: inst = 32'h8620000;
      26032: inst = 32'h10408000;
      26033: inst = 32'hc404d29;
      26034: inst = 32'h8620000;
      26035: inst = 32'hc60a000;
      26036: inst = 32'h10408000;
      26037: inst = 32'hc404cc8;
      26038: inst = 32'h8620000;
      26039: inst = 32'h10408000;
      26040: inst = 32'hc404cc7;
      26041: inst = 32'h8620000;
      26042: inst = 32'h10408000;
      26043: inst = 32'hc404cc6;
      26044: inst = 32'h8620000;
      26045: inst = 32'h10408000;
      26046: inst = 32'hc404cc5;
      26047: inst = 32'h8620000;
      26048: inst = 32'h10408000;
      26049: inst = 32'hc404cc4;
      26050: inst = 32'h8620000;
      26051: inst = 32'h10408000;
      26052: inst = 32'hc404d28;
      26053: inst = 32'h8620000;
      26054: inst = 32'h10408000;
      26055: inst = 32'hc404d26;
      26056: inst = 32'h8620000;
      26057: inst = 32'h10408000;
      26058: inst = 32'hc404d25;
      26059: inst = 32'h8620000;
      26060: inst = 32'h10408000;
      26061: inst = 32'hc404d24;
      26062: inst = 32'h8620000;
      26063: inst = 32'h10408000;
      26064: inst = 32'hc404d89;
      26065: inst = 32'h8620000;
      26066: inst = 32'h10408000;
      26067: inst = 32'hc404d88;
      26068: inst = 32'h8620000;
      26069: inst = 32'h10408000;
      26070: inst = 32'hc404d87;
      26071: inst = 32'h8620000;
      26072: inst = 32'h10408000;
      26073: inst = 32'hc404d86;
      26074: inst = 32'h8620000;
      26075: inst = 32'h10408000;
      26076: inst = 32'hc404d85;
      26077: inst = 32'h8620000;
      26078: inst = 32'h10408000;
      26079: inst = 32'hc404d84;
      26080: inst = 32'h8620000;
      26081: inst = 32'hc6010ac;
      26082: inst = 32'h10408000;
      26083: inst = 32'hc404de9;
      26084: inst = 32'h8620000;
      26085: inst = 32'h10408000;
      26086: inst = 32'hc404de8;
      26087: inst = 32'h8620000;
      26088: inst = 32'h10408000;
      26089: inst = 32'hc404de7;
      26090: inst = 32'h8620000;
      26091: inst = 32'h10408000;
      26092: inst = 32'hc404de6;
      26093: inst = 32'h8620000;
      26094: inst = 32'h10408000;
      26095: inst = 32'hc404de5;
      26096: inst = 32'h8620000;
      26097: inst = 32'h10408000;
      26098: inst = 32'hc404de4;
      26099: inst = 32'h8620000;
      26100: inst = 32'h13e0ffff;
      26101: inst = 32'h13e00000;
      26102: inst = 32'hfe065fb;
      26103: inst = 32'h5be00000;
      26104: inst = 32'h13e00000;
      26105: inst = 32'hfe065fe;
      26106: inst = 32'h5be00000;
      26107: inst = 32'h13e00000;
      26108: inst = 32'hfe065fe;
      26109: inst = 32'h5be00000;
      26110: inst = 32'h58000000;
      26111: inst = 32'h10408000;
      26112: inst = 32'hc400002;
      26113: inst = 32'h4420000;
      26114: inst = 32'h10600000;
      26115: inst = 32'hc600010;
      26116: inst = 32'h38421800;
      26117: inst = 32'h4042000f;
      26118: inst = 32'h1c40000f;
      26119: inst = 32'h58000000;
      26120: inst = 32'h58200000;
    endcase
  end
endmodule
